module basic_2500_25000_3000_25_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_246,In_251);
or U1 (N_1,In_1441,In_2244);
xnor U2 (N_2,In_1083,In_1114);
nand U3 (N_3,In_906,In_419);
nor U4 (N_4,In_1995,In_816);
nor U5 (N_5,In_2124,In_607);
nand U6 (N_6,In_2145,In_1798);
nor U7 (N_7,In_548,In_431);
xor U8 (N_8,In_2243,In_294);
and U9 (N_9,In_943,In_498);
and U10 (N_10,In_503,In_1291);
xor U11 (N_11,In_412,In_2090);
and U12 (N_12,In_689,In_1195);
nor U13 (N_13,In_38,In_2371);
and U14 (N_14,In_1575,In_1813);
nor U15 (N_15,In_1430,In_651);
nor U16 (N_16,In_2466,In_1850);
nor U17 (N_17,In_1810,In_2429);
and U18 (N_18,In_2203,In_111);
xor U19 (N_19,In_197,In_552);
nor U20 (N_20,In_1647,In_2011);
nand U21 (N_21,In_2322,In_541);
nor U22 (N_22,In_2006,In_142);
xor U23 (N_23,In_2084,In_1416);
nor U24 (N_24,In_183,In_1775);
or U25 (N_25,In_585,In_2072);
nor U26 (N_26,In_430,In_1363);
and U27 (N_27,In_528,In_1700);
xnor U28 (N_28,In_1477,In_190);
nand U29 (N_29,In_1787,In_2037);
xor U30 (N_30,In_1208,In_1838);
and U31 (N_31,In_2337,In_1953);
and U32 (N_32,In_1497,In_32);
or U33 (N_33,In_290,In_165);
or U34 (N_34,In_817,In_1827);
nand U35 (N_35,In_2059,In_1724);
nand U36 (N_36,In_923,In_2030);
nand U37 (N_37,In_1256,In_286);
xnor U38 (N_38,In_1920,In_156);
nor U39 (N_39,In_2320,In_1734);
xnor U40 (N_40,In_314,In_268);
and U41 (N_41,In_2132,In_166);
nor U42 (N_42,In_1158,In_2123);
nand U43 (N_43,In_2,In_473);
nor U44 (N_44,In_643,In_2001);
xnor U45 (N_45,In_1139,In_2015);
nand U46 (N_46,In_935,In_465);
nor U47 (N_47,In_729,In_2456);
and U48 (N_48,In_2373,In_1316);
nand U49 (N_49,In_1938,In_949);
and U50 (N_50,In_1485,In_1402);
xnor U51 (N_51,In_1797,In_136);
nand U52 (N_52,In_1173,In_168);
and U53 (N_53,In_2185,In_445);
or U54 (N_54,In_2038,In_233);
xnor U55 (N_55,In_1310,In_1180);
nand U56 (N_56,In_653,In_495);
and U57 (N_57,In_1157,In_1899);
xor U58 (N_58,In_1740,In_561);
xor U59 (N_59,In_1333,In_2008);
nand U60 (N_60,In_2089,In_728);
nor U61 (N_61,In_2211,In_2433);
and U62 (N_62,In_1522,In_2193);
or U63 (N_63,In_471,In_65);
nor U64 (N_64,In_1183,In_411);
and U65 (N_65,In_1892,In_87);
nand U66 (N_66,In_123,In_491);
nand U67 (N_67,In_1220,In_2122);
nor U68 (N_68,In_364,In_1624);
nand U69 (N_69,In_2188,In_570);
xor U70 (N_70,In_2171,In_2368);
xnor U71 (N_71,In_407,In_738);
and U72 (N_72,In_1891,In_776);
or U73 (N_73,In_1658,In_2233);
and U74 (N_74,In_1293,In_72);
nand U75 (N_75,In_1414,In_203);
or U76 (N_76,In_383,In_571);
xor U77 (N_77,In_1520,In_1983);
or U78 (N_78,In_1109,In_1517);
or U79 (N_79,In_686,In_5);
nor U80 (N_80,In_12,In_959);
and U81 (N_81,In_1088,In_226);
or U82 (N_82,In_2436,In_1613);
and U83 (N_83,In_2170,In_103);
or U84 (N_84,In_456,In_596);
and U85 (N_85,In_14,In_1851);
and U86 (N_86,In_1006,In_1816);
nand U87 (N_87,In_1901,In_2022);
xor U88 (N_88,In_1202,In_750);
nor U89 (N_89,In_2146,In_2131);
nand U90 (N_90,In_2109,In_615);
or U91 (N_91,In_1991,In_146);
xnor U92 (N_92,In_1136,In_786);
or U93 (N_93,In_2063,In_1011);
or U94 (N_94,In_2444,In_67);
or U95 (N_95,In_2409,In_1253);
or U96 (N_96,In_1128,In_1799);
or U97 (N_97,In_1100,In_618);
and U98 (N_98,In_800,In_2181);
or U99 (N_99,In_721,In_267);
xor U100 (N_100,In_1640,In_1345);
nor U101 (N_101,In_2484,In_1019);
and U102 (N_102,In_1969,In_1324);
and U103 (N_103,In_1067,In_2443);
nor U104 (N_104,In_892,In_870);
nand U105 (N_105,In_1272,In_1886);
and U106 (N_106,In_112,In_1672);
nand U107 (N_107,In_1465,In_444);
nor U108 (N_108,In_1980,In_1584);
nand U109 (N_109,In_1265,In_2350);
xnor U110 (N_110,In_133,In_809);
nand U111 (N_111,In_2182,In_1817);
or U112 (N_112,In_170,In_89);
and U113 (N_113,In_1839,In_1944);
nand U114 (N_114,In_2199,In_2302);
or U115 (N_115,In_1808,In_296);
or U116 (N_116,In_1752,In_1794);
nand U117 (N_117,In_1326,In_390);
and U118 (N_118,In_1359,In_2414);
nor U119 (N_119,In_1247,In_752);
or U120 (N_120,In_2078,In_512);
and U121 (N_121,In_1962,In_1832);
or U122 (N_122,In_231,In_1713);
nand U123 (N_123,In_1072,In_2025);
or U124 (N_124,In_1726,In_1244);
nand U125 (N_125,In_2057,In_19);
or U126 (N_126,In_864,In_1870);
xnor U127 (N_127,In_2021,In_2246);
nand U128 (N_128,In_159,In_1593);
nor U129 (N_129,In_104,In_1421);
nand U130 (N_130,In_2305,In_118);
nand U131 (N_131,In_1046,In_536);
and U132 (N_132,In_2100,In_1668);
nor U133 (N_133,In_455,In_1388);
nor U134 (N_134,In_1468,In_458);
nor U135 (N_135,In_1720,In_2391);
or U136 (N_136,In_303,In_2134);
nand U137 (N_137,In_534,In_780);
xor U138 (N_138,In_779,In_815);
nand U139 (N_139,In_692,In_626);
and U140 (N_140,In_256,In_2272);
or U141 (N_141,In_356,In_1507);
and U142 (N_142,In_1677,In_119);
and U143 (N_143,In_1286,In_460);
or U144 (N_144,In_2197,In_2251);
nand U145 (N_145,In_485,In_2164);
and U146 (N_146,In_1634,In_1274);
and U147 (N_147,In_253,In_1262);
nor U148 (N_148,In_1612,In_1177);
or U149 (N_149,In_1340,In_590);
nor U150 (N_150,In_1225,In_1214);
nand U151 (N_151,In_249,In_1091);
or U152 (N_152,In_2394,In_82);
nor U153 (N_153,In_1488,In_1943);
or U154 (N_154,In_154,In_2329);
or U155 (N_155,In_898,In_223);
nor U156 (N_156,In_746,In_1629);
and U157 (N_157,In_2256,In_1048);
nand U158 (N_158,In_813,In_2447);
or U159 (N_159,In_1496,In_241);
and U160 (N_160,In_1346,In_1308);
nor U161 (N_161,In_1967,In_574);
nand U162 (N_162,In_436,In_1552);
nand U163 (N_163,In_1864,In_848);
and U164 (N_164,In_1550,In_1765);
nand U165 (N_165,In_261,In_1207);
xnor U166 (N_166,In_1948,In_2195);
nor U167 (N_167,In_369,In_913);
or U168 (N_168,In_794,In_1628);
and U169 (N_169,In_1354,In_1319);
xnor U170 (N_170,In_164,In_69);
and U171 (N_171,In_1108,In_91);
or U172 (N_172,In_986,In_10);
nor U173 (N_173,In_2288,In_175);
nor U174 (N_174,In_1130,In_1587);
or U175 (N_175,In_2128,In_2151);
xnor U176 (N_176,In_2293,In_631);
nand U177 (N_177,In_519,In_228);
or U178 (N_178,In_2055,In_796);
or U179 (N_179,In_857,In_1877);
nand U180 (N_180,In_215,In_2376);
nand U181 (N_181,In_2052,In_1396);
and U182 (N_182,In_127,In_956);
xor U183 (N_183,In_1945,In_2228);
nor U184 (N_184,In_1446,In_1600);
or U185 (N_185,In_1674,In_374);
xor U186 (N_186,In_1410,In_1954);
xor U187 (N_187,In_1859,In_1748);
nor U188 (N_188,In_106,In_1737);
nor U189 (N_189,In_23,In_1411);
nand U190 (N_190,In_1486,In_524);
nand U191 (N_191,In_2277,In_1524);
or U192 (N_192,In_1979,In_821);
nor U193 (N_193,In_1175,In_1408);
xnor U194 (N_194,In_218,In_1074);
nor U195 (N_195,In_274,In_844);
or U196 (N_196,In_2278,In_1518);
nand U197 (N_197,In_860,In_1124);
or U198 (N_198,In_2377,In_2083);
xor U199 (N_199,In_375,In_2452);
or U200 (N_200,In_696,In_2460);
or U201 (N_201,In_1289,In_1106);
xor U202 (N_202,In_1875,In_143);
or U203 (N_203,In_1435,In_772);
and U204 (N_204,In_1656,In_426);
nand U205 (N_205,In_1662,In_845);
or U206 (N_206,In_1768,In_2117);
or U207 (N_207,In_377,In_505);
nor U208 (N_208,In_1878,In_1467);
and U209 (N_209,In_1927,In_1125);
nor U210 (N_210,In_351,In_598);
or U211 (N_211,In_1131,In_1523);
nor U212 (N_212,In_1546,In_1320);
xnor U213 (N_213,In_2381,In_70);
and U214 (N_214,In_2494,In_2470);
nor U215 (N_215,In_646,In_824);
xor U216 (N_216,In_1189,In_1163);
nor U217 (N_217,In_791,In_157);
and U218 (N_218,In_2156,In_874);
nor U219 (N_219,In_2121,In_348);
or U220 (N_220,In_1348,In_1578);
nand U221 (N_221,In_1454,In_2372);
nor U222 (N_222,In_988,In_397);
nand U223 (N_223,In_2398,In_2060);
and U224 (N_224,In_1260,In_2374);
or U225 (N_225,In_1843,In_1494);
or U226 (N_226,In_2205,In_2370);
or U227 (N_227,In_1044,In_1473);
nand U228 (N_228,In_318,In_808);
nand U229 (N_229,In_2492,In_1182);
and U230 (N_230,In_248,In_1423);
nand U231 (N_231,In_1258,In_939);
nand U232 (N_232,In_184,In_773);
nor U233 (N_233,In_202,In_1480);
nor U234 (N_234,In_2094,In_176);
xnor U235 (N_235,In_2343,In_526);
nor U236 (N_236,In_575,In_2497);
xnor U237 (N_237,In_2112,In_468);
nor U238 (N_238,In_1929,In_1982);
and U239 (N_239,In_1322,In_1660);
nor U240 (N_240,In_555,In_214);
and U241 (N_241,In_99,In_2073);
and U242 (N_242,In_662,In_2058);
nor U243 (N_243,In_2104,In_1919);
and U244 (N_244,In_2077,In_459);
xnor U245 (N_245,In_350,In_167);
nor U246 (N_246,In_2441,In_1950);
nand U247 (N_247,In_1916,In_1167);
or U248 (N_248,In_2189,In_151);
or U249 (N_249,In_1984,In_990);
nand U250 (N_250,In_991,In_1707);
nor U251 (N_251,In_1837,In_2388);
nand U252 (N_252,In_305,In_636);
xor U253 (N_253,In_2066,In_843);
xor U254 (N_254,In_1470,In_35);
nand U255 (N_255,In_1392,In_1655);
or U256 (N_256,In_915,In_47);
xnor U257 (N_257,In_1543,In_1830);
xnor U258 (N_258,In_1528,In_881);
nor U259 (N_259,In_1554,In_1825);
nand U260 (N_260,In_819,In_1921);
nand U261 (N_261,In_1669,In_889);
nor U262 (N_262,In_1042,In_2389);
nor U263 (N_263,In_1299,In_987);
and U264 (N_264,In_442,In_1013);
and U265 (N_265,In_1425,In_464);
and U266 (N_266,In_885,In_404);
and U267 (N_267,In_288,In_1712);
nor U268 (N_268,In_677,In_358);
nand U269 (N_269,In_114,In_625);
xnor U270 (N_270,In_567,In_2431);
or U271 (N_271,In_622,In_2312);
or U272 (N_272,In_1598,In_2029);
and U273 (N_273,In_2307,In_1907);
xnor U274 (N_274,In_1696,In_1164);
xnor U275 (N_275,In_1273,In_1458);
and U276 (N_276,In_1012,In_1084);
and U277 (N_277,In_2331,In_1498);
or U278 (N_278,In_2005,In_532);
xnor U279 (N_279,In_80,In_833);
or U280 (N_280,In_583,In_1481);
or U281 (N_281,In_74,In_1478);
xor U282 (N_282,In_593,In_985);
and U283 (N_283,In_1888,In_2369);
xor U284 (N_284,In_1802,In_2014);
nor U285 (N_285,In_2040,In_1255);
nor U286 (N_286,In_1024,In_1034);
or U287 (N_287,In_483,In_1197);
xnor U288 (N_288,In_1039,In_806);
nor U289 (N_289,In_1357,In_487);
xor U290 (N_290,In_605,In_1460);
nor U291 (N_291,In_1176,In_1156);
and U292 (N_292,In_2098,In_1236);
and U293 (N_293,In_588,In_982);
or U294 (N_294,In_1705,In_1592);
and U295 (N_295,In_448,In_2150);
and U296 (N_296,In_679,In_1860);
or U297 (N_297,In_1235,In_797);
or U298 (N_298,In_1956,In_2129);
and U299 (N_299,In_266,In_171);
and U300 (N_300,In_2476,In_116);
nand U301 (N_301,In_878,In_2355);
or U302 (N_302,In_2438,In_1519);
nor U303 (N_303,In_153,In_531);
nor U304 (N_304,In_716,In_763);
nand U305 (N_305,In_362,In_1026);
or U306 (N_306,In_2314,In_11);
or U307 (N_307,In_2324,In_335);
nand U308 (N_308,In_2088,In_1788);
xnor U309 (N_309,In_467,In_1332);
nand U310 (N_310,In_1051,In_1449);
or U311 (N_311,In_1654,In_2126);
and U312 (N_312,In_393,In_2190);
xor U313 (N_313,In_1409,In_1107);
nor U314 (N_314,In_258,In_1190);
xor U315 (N_315,In_2400,In_387);
xor U316 (N_316,In_178,In_90);
nor U317 (N_317,In_1532,In_1703);
nand U318 (N_318,In_1213,In_937);
and U319 (N_319,In_2280,In_392);
nand U320 (N_320,In_649,In_1922);
and U321 (N_321,In_1635,In_403);
and U322 (N_322,In_1290,In_1772);
and U323 (N_323,In_997,In_370);
nand U324 (N_324,In_940,In_1254);
nor U325 (N_325,In_149,In_2289);
nor U326 (N_326,In_556,In_970);
and U327 (N_327,In_658,In_2475);
xnor U328 (N_328,In_2119,In_1725);
or U329 (N_329,In_1504,In_737);
nand U330 (N_330,In_2493,In_659);
nor U331 (N_331,In_690,In_788);
xnor U332 (N_332,In_135,In_1355);
or U333 (N_333,In_1501,In_1721);
nor U334 (N_334,In_782,In_2327);
or U335 (N_335,In_1054,In_757);
and U336 (N_336,In_1942,In_616);
or U337 (N_337,In_1469,In_688);
and U338 (N_338,In_1148,In_1426);
nand U339 (N_339,In_1372,In_2264);
xnor U340 (N_340,In_51,In_2361);
nor U341 (N_341,In_2483,In_989);
nand U342 (N_342,In_862,In_1579);
nor U343 (N_343,In_1229,In_1754);
xnor U344 (N_344,In_1495,In_1599);
nand U345 (N_345,In_1377,In_1898);
nand U346 (N_346,In_1933,In_1362);
and U347 (N_347,In_1018,In_875);
or U348 (N_348,In_2294,In_2056);
nor U349 (N_349,In_319,In_1951);
xor U350 (N_350,In_46,In_179);
nand U351 (N_351,In_1476,In_841);
nand U352 (N_352,In_1219,In_1037);
xor U353 (N_353,In_1249,In_128);
nand U354 (N_354,In_193,In_2212);
or U355 (N_355,In_1492,In_1147);
xnor U356 (N_356,In_617,In_1076);
nor U357 (N_357,In_191,In_2292);
xor U358 (N_358,In_1344,In_1815);
or U359 (N_359,In_2044,In_909);
or U360 (N_360,In_2136,In_1077);
nand U361 (N_361,In_2408,In_1230);
nor U362 (N_362,In_324,In_2255);
or U363 (N_363,In_1152,In_1323);
xor U364 (N_364,In_1420,In_384);
nand U365 (N_365,In_840,In_944);
and U366 (N_366,In_2419,In_1267);
or U367 (N_367,In_2249,In_1116);
nor U368 (N_368,In_1089,In_1706);
nand U369 (N_369,In_667,In_914);
xor U370 (N_370,In_1664,In_1111);
or U371 (N_371,In_654,In_2477);
or U372 (N_372,In_2236,In_490);
or U373 (N_373,In_2213,In_1840);
or U374 (N_374,In_1560,In_447);
or U375 (N_375,In_601,In_1279);
and U376 (N_376,In_2157,In_1149);
or U377 (N_377,In_1889,In_2219);
xnor U378 (N_378,In_2092,In_417);
and U379 (N_379,In_921,In_731);
nand U380 (N_380,In_1561,In_1678);
or U381 (N_381,In_742,In_2340);
nor U382 (N_382,In_2403,In_60);
xor U383 (N_383,In_1973,In_2216);
and U384 (N_384,In_141,In_26);
or U385 (N_385,In_2323,In_2245);
nand U386 (N_386,In_2455,In_2375);
and U387 (N_387,In_2160,In_767);
or U388 (N_388,In_229,In_1146);
nand U389 (N_389,In_1911,In_199);
nor U390 (N_390,In_814,In_1031);
or U391 (N_391,In_2478,In_2379);
nand U392 (N_392,In_420,In_735);
or U393 (N_393,In_2486,In_352);
or U394 (N_394,In_1017,In_1895);
or U395 (N_395,In_1620,In_2267);
and U396 (N_396,In_1849,In_276);
nand U397 (N_397,In_748,In_1555);
and U398 (N_398,In_507,In_105);
nor U399 (N_399,In_2107,In_993);
nor U400 (N_400,In_357,In_1387);
xor U401 (N_401,In_2163,In_2495);
and U402 (N_402,In_2306,In_323);
xnor U403 (N_403,In_754,In_1763);
nor U404 (N_404,In_409,In_2465);
and U405 (N_405,In_934,In_1580);
xnor U406 (N_406,In_1661,In_1221);
nand U407 (N_407,In_68,In_1440);
nand U408 (N_408,In_1766,In_185);
xnor U409 (N_409,In_2259,In_482);
nand U410 (N_410,In_2162,In_2062);
nor U411 (N_411,In_832,In_2106);
xor U412 (N_412,In_1761,In_1779);
nor U413 (N_413,In_1193,In_1959);
or U414 (N_414,In_2242,In_2127);
nor U415 (N_415,In_1646,In_2018);
nor U416 (N_416,In_573,In_488);
nand U417 (N_417,In_926,In_492);
xor U418 (N_418,In_1746,In_1785);
or U419 (N_419,In_945,In_1399);
nor U420 (N_420,In_1756,In_1665);
nand U421 (N_421,In_1893,In_1404);
nand U422 (N_422,In_1744,In_2023);
xor U423 (N_423,In_1003,In_1904);
xor U424 (N_424,In_922,In_1818);
xnor U425 (N_425,In_1949,In_1004);
and U426 (N_426,In_500,In_2087);
or U427 (N_427,In_1294,In_938);
and U428 (N_428,In_770,In_2054);
nor U429 (N_429,In_978,In_1887);
nand U430 (N_430,In_1010,In_852);
xor U431 (N_431,In_1287,In_1852);
xnor U432 (N_432,In_701,In_299);
xnor U433 (N_433,In_2168,In_602);
nor U434 (N_434,In_1800,In_927);
nand U435 (N_435,In_1078,In_1227);
xnor U436 (N_436,In_2009,In_1671);
nand U437 (N_437,In_1179,In_315);
or U438 (N_438,In_1917,In_1814);
xnor U439 (N_439,In_3,In_2184);
nand U440 (N_440,In_1924,In_2224);
and U441 (N_441,In_2393,In_2165);
nand U442 (N_442,In_1753,In_341);
and U443 (N_443,In_671,In_186);
or U444 (N_444,In_1226,In_1269);
and U445 (N_445,In_1276,In_1419);
and U446 (N_446,In_2366,In_1585);
xor U447 (N_447,In_1448,In_1104);
xnor U448 (N_448,In_2206,In_401);
and U449 (N_449,In_1978,In_463);
xor U450 (N_450,In_1591,In_1187);
nand U451 (N_451,In_976,In_1038);
or U452 (N_452,In_1015,In_962);
nor U453 (N_453,In_744,In_1701);
and U454 (N_454,In_2413,In_1025);
or U455 (N_455,In_1375,In_830);
and U456 (N_456,In_1994,In_423);
xnor U457 (N_457,In_869,In_1963);
or U458 (N_458,In_1988,In_2392);
nand U459 (N_459,In_916,In_1456);
or U460 (N_460,In_2308,In_1536);
or U461 (N_461,In_1977,In_2420);
xnor U462 (N_462,In_272,In_254);
or U463 (N_463,In_1563,In_1021);
nor U464 (N_464,In_1621,In_1383);
and U465 (N_465,In_2296,In_2003);
xor U466 (N_466,In_2461,In_1397);
nand U467 (N_467,In_331,In_2095);
xnor U468 (N_468,In_73,In_1191);
nor U469 (N_469,In_1045,In_784);
xor U470 (N_470,In_1394,In_908);
nor U471 (N_471,In_180,In_563);
or U472 (N_472,In_858,In_1606);
nor U473 (N_473,In_1718,In_297);
or U474 (N_474,In_515,In_1594);
nor U475 (N_475,In_1196,In_2238);
or U476 (N_476,In_353,In_477);
or U477 (N_477,In_525,In_879);
nor U478 (N_478,In_1069,In_1464);
xor U479 (N_479,In_230,In_514);
and U480 (N_480,In_155,In_2020);
or U481 (N_481,In_2035,In_1502);
and U482 (N_482,In_504,In_1301);
or U483 (N_483,In_1568,In_1861);
nand U484 (N_484,In_1940,In_1424);
nor U485 (N_485,In_257,In_1443);
nand U486 (N_486,In_1902,In_568);
nand U487 (N_487,In_196,In_2489);
nand U488 (N_488,In_790,In_29);
xnor U489 (N_489,In_1288,In_306);
and U490 (N_490,In_1846,In_21);
and U491 (N_491,In_714,In_506);
or U492 (N_492,In_1801,In_842);
and U493 (N_493,In_542,In_1261);
nor U494 (N_494,In_182,In_1442);
xor U495 (N_495,In_64,In_1343);
nand U496 (N_496,In_1341,In_1311);
xnor U497 (N_497,In_1831,In_1459);
or U498 (N_498,In_2342,In_2004);
nor U499 (N_499,In_2177,In_1514);
and U500 (N_500,In_405,In_1466);
xnor U501 (N_501,In_97,In_2075);
or U502 (N_502,In_325,In_1393);
nor U503 (N_503,In_371,In_1493);
nand U504 (N_504,In_2458,In_386);
nor U505 (N_505,In_2354,In_1023);
nor U506 (N_506,In_2446,In_1565);
and U507 (N_507,In_2139,In_2265);
or U508 (N_508,In_309,In_117);
xnor U509 (N_509,In_1728,In_1047);
nor U510 (N_510,In_295,In_2103);
nand U511 (N_511,In_1542,In_826);
xor U512 (N_512,In_2260,In_1926);
xnor U513 (N_513,In_243,In_422);
and U514 (N_514,In_227,In_2232);
xor U515 (N_515,In_1162,In_2387);
nand U516 (N_516,In_208,In_2442);
xor U517 (N_517,In_1049,In_2031);
nand U518 (N_518,In_928,In_494);
xor U519 (N_519,In_2462,In_640);
and U520 (N_520,In_917,In_544);
nand U521 (N_521,In_1437,In_2194);
nor U522 (N_522,In_1650,In_216);
xor U523 (N_523,In_967,In_478);
nor U524 (N_524,In_1014,In_2286);
nand U525 (N_525,In_560,In_1704);
xor U526 (N_526,In_726,In_785);
and U527 (N_527,In_1248,In_207);
or U528 (N_528,In_756,In_893);
nor U529 (N_529,In_1822,In_1548);
nand U530 (N_530,In_1989,In_1540);
and U531 (N_531,In_2417,In_547);
or U532 (N_532,In_326,In_1491);
nor U533 (N_533,In_802,In_1836);
and U534 (N_534,In_1095,In_687);
nand U535 (N_535,In_2347,In_224);
xor U536 (N_536,In_1259,In_2336);
nor U537 (N_537,In_76,In_2352);
and U538 (N_538,In_2247,In_2315);
nor U539 (N_539,In_1958,In_1867);
and U540 (N_540,In_1129,In_741);
xor U541 (N_541,In_2013,In_1667);
xor U542 (N_542,In_1809,In_2027);
or U543 (N_543,In_2469,In_1622);
nor U544 (N_544,In_1562,In_234);
xnor U545 (N_545,In_1185,In_1856);
and U546 (N_546,In_2330,In_1337);
nor U547 (N_547,In_1525,In_664);
nor U548 (N_548,In_521,In_1747);
xnor U549 (N_549,In_1303,In_1834);
or U550 (N_550,In_1807,In_1215);
or U551 (N_551,In_2108,In_1334);
nor U552 (N_552,In_1615,In_2344);
nor U553 (N_553,In_2445,In_1688);
nor U554 (N_554,In_1643,In_545);
xnor U555 (N_555,In_699,In_1285);
or U556 (N_556,In_1796,In_2421);
or U557 (N_557,In_213,In_537);
nor U558 (N_558,In_1068,In_432);
and U559 (N_559,In_433,In_2479);
and U560 (N_560,In_961,In_1367);
or U561 (N_561,In_413,In_1854);
nor U562 (N_562,In_2099,In_2217);
or U563 (N_563,In_520,In_656);
and U564 (N_564,In_1342,In_1602);
nand U565 (N_565,In_1113,In_700);
and U566 (N_566,In_1365,In_1586);
nand U567 (N_567,In_867,In_2353);
nor U568 (N_568,In_49,In_553);
nor U569 (N_569,In_2356,In_1406);
and U570 (N_570,In_1858,In_1842);
or U571 (N_571,In_1738,In_781);
nand U572 (N_572,In_2069,In_1739);
nand U573 (N_573,In_2214,In_2430);
nand U574 (N_574,In_2042,In_807);
nand U575 (N_575,In_1166,In_2328);
xor U576 (N_576,In_1745,In_1900);
xor U577 (N_577,In_1064,In_438);
nand U578 (N_578,In_1509,In_502);
xor U579 (N_579,In_691,In_2457);
or U580 (N_580,In_2363,In_1691);
xnor U581 (N_581,In_2333,In_2153);
and U582 (N_582,In_1243,In_1931);
nor U583 (N_583,In_670,In_2178);
and U584 (N_584,In_1511,In_2076);
nor U585 (N_585,In_695,In_2482);
nor U586 (N_586,In_895,In_96);
xnor U587 (N_587,In_1237,In_57);
nor U588 (N_588,In_195,In_1429);
or U589 (N_589,In_1936,In_1595);
nor U590 (N_590,In_1092,In_1648);
nand U591 (N_591,In_328,In_727);
and U592 (N_592,In_1263,In_2276);
and U593 (N_593,In_2454,In_1475);
xor U594 (N_594,In_1389,In_1063);
nand U595 (N_595,In_2273,In_1144);
or U596 (N_596,In_2406,In_1118);
and U597 (N_597,In_1251,In_883);
nor U598 (N_598,In_609,In_1376);
and U599 (N_599,In_2326,In_134);
and U600 (N_600,In_1829,In_457);
and U601 (N_601,In_2176,In_1928);
nor U602 (N_602,In_551,In_1804);
nand U603 (N_603,In_920,In_2180);
and U604 (N_604,In_912,In_206);
nand U605 (N_605,In_903,In_1431);
or U606 (N_606,In_1264,In_1823);
nand U607 (N_607,In_8,In_1329);
nand U608 (N_608,In_1769,In_1645);
or U609 (N_609,In_1325,In_932);
nand U610 (N_610,In_783,In_1022);
nand U611 (N_611,In_408,In_395);
and U612 (N_612,In_2048,In_977);
nor U613 (N_613,In_2226,In_1056);
nor U614 (N_614,In_2474,In_1360);
xnor U615 (N_615,In_372,In_584);
nor U616 (N_616,In_416,In_345);
nor U617 (N_617,In_774,In_1137);
xnor U618 (N_618,In_132,In_1266);
and U619 (N_619,In_344,In_421);
nor U620 (N_620,In_1352,In_1217);
nor U621 (N_621,In_2196,In_1783);
or U622 (N_622,In_628,In_1422);
xor U623 (N_623,In_2110,In_1857);
nor U624 (N_624,In_308,In_733);
or U625 (N_625,In_1890,In_1719);
and U626 (N_626,In_242,In_668);
xor U627 (N_627,In_2316,In_1702);
nand U628 (N_628,In_1110,In_676);
or U629 (N_629,In_2167,In_337);
nand U630 (N_630,In_188,In_84);
and U631 (N_631,In_1998,In_110);
nand U632 (N_632,In_367,In_623);
nand U633 (N_633,In_595,In_1134);
nor U634 (N_634,In_169,In_1597);
nand U635 (N_635,In_1427,In_1304);
nor U636 (N_636,In_1708,In_650);
nand U637 (N_637,In_890,In_1181);
and U638 (N_638,In_918,In_311);
or U639 (N_639,In_680,In_2471);
and U640 (N_640,In_675,In_666);
xor U641 (N_641,In_284,In_313);
xor U642 (N_642,In_2270,In_265);
or U643 (N_643,In_277,In_1053);
or U644 (N_644,In_131,In_1793);
nand U645 (N_645,In_298,In_1627);
nor U646 (N_646,In_1512,In_720);
xor U647 (N_647,In_1307,In_1371);
nor U648 (N_648,In_2348,In_1663);
nor U649 (N_649,In_354,In_282);
or U650 (N_650,In_148,In_1234);
or U651 (N_651,In_1418,In_1675);
xor U652 (N_652,In_378,In_388);
or U653 (N_653,In_1617,In_302);
xor U654 (N_654,In_2291,In_1228);
and U655 (N_655,In_1882,In_1690);
nor U656 (N_656,In_174,In_2472);
and U657 (N_657,In_511,In_334);
and U658 (N_658,In_713,In_2487);
nor U659 (N_659,In_2240,In_517);
or U660 (N_660,In_1611,In_1642);
or U661 (N_661,In_1727,In_1242);
or U662 (N_662,In_2459,In_1847);
or U663 (N_663,In_1596,In_58);
xnor U664 (N_664,In_1052,In_1370);
xor U665 (N_665,In_48,In_2252);
or U666 (N_666,In_1709,In_107);
or U667 (N_667,In_1302,In_1576);
and U668 (N_668,In_2271,In_24);
nand U669 (N_669,In_376,In_1161);
and U670 (N_670,In_373,In_2235);
nor U671 (N_671,In_1194,In_1641);
and U672 (N_672,In_569,In_1897);
xnor U673 (N_673,In_28,In_919);
and U674 (N_674,In_1281,In_1059);
xnor U675 (N_675,In_1760,In_1820);
nand U676 (N_676,In_2120,In_150);
nor U677 (N_677,In_1687,In_1484);
nor U678 (N_678,In_238,In_2362);
nand U679 (N_679,In_2318,In_1623);
or U680 (N_680,In_1805,In_2485);
or U681 (N_681,In_59,In_2017);
and U682 (N_682,In_2097,In_722);
and U683 (N_683,In_2116,In_759);
nand U684 (N_684,In_2125,In_2105);
and U685 (N_685,In_672,In_1444);
nand U686 (N_686,In_1246,In_1450);
or U687 (N_687,In_1101,In_2341);
or U688 (N_688,In_942,In_1366);
and U689 (N_689,In_1122,In_831);
and U690 (N_690,In_891,In_732);
nand U691 (N_691,In_1071,In_361);
nor U692 (N_692,In_1349,In_1682);
nor U693 (N_693,In_2423,In_1210);
xnor U694 (N_694,In_1997,In_52);
xnor U695 (N_695,In_1380,In_1417);
or U696 (N_696,In_1698,In_2229);
nand U697 (N_697,In_2222,In_454);
or U698 (N_698,In_2453,In_2439);
nor U699 (N_699,In_2173,In_627);
xnor U700 (N_700,In_2133,In_1506);
and U701 (N_701,In_866,In_1780);
and U702 (N_702,In_522,In_2378);
or U703 (N_703,In_1201,In_724);
nand U704 (N_704,In_566,In_854);
or U705 (N_705,In_270,In_663);
nor U706 (N_706,In_1335,In_1205);
xnor U707 (N_707,In_888,In_108);
nor U708 (N_708,In_992,In_1020);
nand U709 (N_709,In_1445,In_2425);
nand U710 (N_710,In_453,In_639);
or U711 (N_711,In_321,In_2186);
and U712 (N_712,In_1903,In_75);
nand U713 (N_713,In_1755,In_2281);
and U714 (N_714,In_1451,In_37);
and U715 (N_715,In_2448,In_1065);
xnor U716 (N_716,In_2287,In_262);
nand U717 (N_717,In_1123,In_619);
nand U718 (N_718,In_1941,In_414);
and U719 (N_719,In_449,In_1913);
xor U720 (N_720,In_2297,In_882);
and U721 (N_721,In_2338,In_851);
xnor U722 (N_722,In_865,In_34);
xor U723 (N_723,In_122,In_1534);
nand U724 (N_724,In_1240,In_947);
xnor U725 (N_725,In_1970,In_475);
and U726 (N_726,In_1035,In_1633);
or U727 (N_727,In_589,In_222);
nand U728 (N_728,In_880,In_172);
nand U729 (N_729,In_92,In_572);
and U730 (N_730,In_1996,In_98);
nand U731 (N_731,In_1614,In_530);
or U732 (N_732,In_1767,In_2405);
and U733 (N_733,In_538,In_1117);
and U734 (N_734,In_236,In_793);
and U735 (N_735,In_2093,In_513);
and U736 (N_736,In_1499,In_1577);
nand U737 (N_737,In_1364,In_2074);
nand U738 (N_738,In_829,In_204);
or U739 (N_739,In_2274,In_810);
and U740 (N_740,In_264,In_894);
and U741 (N_741,In_1438,In_1694);
nand U742 (N_742,In_201,In_768);
and U743 (N_743,In_1103,In_428);
and U744 (N_744,In_734,In_884);
xnor U745 (N_745,In_1239,In_979);
xnor U746 (N_746,In_33,In_958);
and U747 (N_747,In_836,In_1043);
nor U748 (N_748,In_2138,In_2113);
nand U749 (N_749,In_901,In_693);
xor U750 (N_750,In_245,In_2434);
nor U751 (N_751,In_644,In_685);
or U752 (N_752,In_2283,In_2385);
nor U753 (N_753,In_7,In_2158);
and U754 (N_754,In_896,In_1005);
and U755 (N_755,In_486,In_2351);
nand U756 (N_756,In_1203,In_220);
and U757 (N_757,In_2192,In_93);
and U758 (N_758,In_1717,In_1680);
or U759 (N_759,In_1073,In_2473);
nor U760 (N_760,In_1759,In_45);
nand U761 (N_761,In_1058,In_771);
nand U762 (N_762,In_1573,In_1385);
nand U763 (N_763,In_861,In_899);
xnor U764 (N_764,In_173,In_820);
nand U765 (N_765,In_1777,In_418);
nor U766 (N_766,In_973,In_145);
or U767 (N_767,In_493,In_22);
and U768 (N_768,In_260,In_2187);
and U769 (N_769,In_966,In_291);
xnor U770 (N_770,In_1403,In_1601);
or U771 (N_771,In_1905,In_1439);
or U772 (N_772,In_529,In_1508);
xor U773 (N_773,In_725,In_630);
and U774 (N_774,In_6,In_1915);
nand U775 (N_775,In_1165,In_1126);
or U776 (N_776,In_2467,In_332);
and U777 (N_777,In_360,In_1541);
xnor U778 (N_778,In_2335,In_1075);
nand U779 (N_779,In_1297,In_124);
and U780 (N_780,In_31,In_1918);
and U781 (N_781,In_1009,In_2464);
nor U782 (N_782,In_1127,In_1758);
or U783 (N_783,In_1955,In_1711);
or U784 (N_784,In_1869,In_9);
and U785 (N_785,In_1676,In_2135);
and U786 (N_786,In_2039,In_489);
xnor U787 (N_787,In_130,In_2221);
xnor U788 (N_788,In_330,In_1199);
nor U789 (N_789,In_1061,In_316);
nand U790 (N_790,In_285,In_579);
and U791 (N_791,In_1331,In_834);
or U792 (N_792,In_2068,In_2012);
and U793 (N_793,In_446,In_1781);
nor U794 (N_794,In_971,In_1786);
or U795 (N_795,In_641,In_1863);
nand U796 (N_796,In_484,In_2435);
nor U797 (N_797,In_496,In_327);
nand U798 (N_798,In_1681,In_610);
and U799 (N_799,In_1007,In_1521);
nand U800 (N_800,In_948,In_129);
nand U801 (N_801,In_1732,In_1742);
xnor U802 (N_802,In_240,In_1689);
or U803 (N_803,In_710,In_2401);
or U804 (N_804,In_2064,In_1551);
or U805 (N_805,In_795,In_398);
and U806 (N_806,In_2141,In_2261);
and U807 (N_807,In_1280,In_95);
xnor U808 (N_808,In_1605,In_876);
or U809 (N_809,In_805,In_1378);
and U810 (N_810,In_1588,In_289);
and U811 (N_811,In_1966,In_1218);
xor U812 (N_812,In_1729,In_1821);
nor U813 (N_813,In_766,In_2026);
nand U814 (N_814,In_1774,In_981);
nor U815 (N_815,In_499,In_307);
and U816 (N_816,In_705,In_1209);
nand U817 (N_817,In_1200,In_77);
or U818 (N_818,In_924,In_2300);
nor U819 (N_819,In_2339,In_1057);
and U820 (N_820,In_2349,In_789);
xor U821 (N_821,In_1666,In_564);
nor U822 (N_822,In_1300,In_1872);
nor U823 (N_823,In_2313,In_1224);
and U824 (N_824,In_822,In_1313);
xnor U825 (N_825,In_1268,In_1170);
nand U826 (N_826,In_210,In_539);
xnor U827 (N_827,In_1041,In_1939);
nor U828 (N_828,In_1330,In_2191);
or U829 (N_829,In_2140,In_1539);
nor U830 (N_830,In_2395,In_846);
nor U831 (N_831,In_61,In_1699);
nand U832 (N_832,In_15,In_1960);
or U833 (N_833,In_147,In_1604);
xor U834 (N_834,In_2225,In_582);
nor U835 (N_835,In_1008,In_681);
xor U836 (N_836,In_1413,In_2301);
and U837 (N_837,In_349,In_969);
or U838 (N_838,In_1743,In_642);
xnor U839 (N_839,In_2114,In_2016);
nor U840 (N_840,In_2215,In_391);
nand U841 (N_841,In_1673,In_336);
xor U842 (N_842,In_718,In_1638);
xnor U843 (N_843,In_647,In_2000);
and U844 (N_844,In_271,In_877);
nor U845 (N_845,In_435,In_162);
or U846 (N_846,In_2045,In_706);
nor U847 (N_847,In_953,In_1462);
nor U848 (N_848,In_2468,In_1692);
or U849 (N_849,In_86,In_1603);
or U850 (N_850,In_1407,In_79);
xnor U851 (N_851,In_1790,In_1657);
nor U852 (N_852,In_2346,In_2161);
or U853 (N_853,In_1885,In_632);
and U854 (N_854,In_1145,In_2290);
nor U855 (N_855,In_2262,In_2299);
nand U856 (N_856,In_925,In_2390);
xnor U857 (N_857,In_683,In_755);
nand U858 (N_858,In_1992,In_2411);
xnor U859 (N_859,In_964,In_219);
xor U860 (N_860,In_1453,In_339);
nand U861 (N_861,In_871,In_329);
or U862 (N_862,In_2410,In_2269);
xnor U863 (N_863,In_1975,In_1472);
and U864 (N_864,In_1947,In_2085);
nand U865 (N_865,In_1571,In_2295);
nor U866 (N_866,In_1029,In_2426);
or U867 (N_867,In_1186,In_2399);
and U868 (N_868,In_1327,In_17);
nand U869 (N_869,In_980,In_762);
and U870 (N_870,In_1296,In_1062);
nor U871 (N_871,In_1,In_2147);
or U872 (N_872,In_581,In_1222);
nor U873 (N_873,In_1770,In_974);
xnor U874 (N_874,In_2263,In_587);
nand U875 (N_875,In_1981,In_1590);
xor U876 (N_876,In_1537,In_381);
xnor U877 (N_877,In_44,In_1559);
and U878 (N_878,In_2081,In_1487);
or U879 (N_879,In_1844,In_1993);
nand U880 (N_880,In_1060,In_36);
xnor U881 (N_881,In_1490,In_1516);
nor U882 (N_882,In_63,In_1723);
or U883 (N_883,In_469,In_900);
nand U884 (N_884,In_53,In_745);
nor U885 (N_885,In_1401,In_40);
nand U886 (N_886,In_2179,In_2144);
and U887 (N_887,In_1474,In_472);
nand U888 (N_888,In_1686,In_540);
nor U889 (N_889,In_1792,In_1632);
nand U890 (N_890,In_2234,In_2220);
xor U891 (N_891,In_217,In_2266);
xor U892 (N_892,In_1538,In_479);
nand U893 (N_893,In_1455,In_1652);
nor U894 (N_894,In_2154,In_1154);
or U895 (N_895,In_269,In_527);
nand U896 (N_896,In_1278,In_255);
nor U897 (N_897,In_71,In_804);
nor U898 (N_898,In_2051,In_2449);
xnor U899 (N_899,In_439,In_760);
xor U900 (N_900,In_205,In_1277);
or U901 (N_901,In_2496,In_25);
xnor U902 (N_902,In_719,In_678);
xnor U903 (N_903,In_2364,In_2480);
or U904 (N_904,In_2428,In_1835);
nand U905 (N_905,In_778,In_1500);
nand U906 (N_906,In_2298,In_279);
xnor U907 (N_907,In_1353,In_2137);
or U908 (N_908,In_614,In_41);
nand U909 (N_909,In_1855,In_209);
xor U910 (N_910,In_1986,In_1976);
nor U911 (N_911,In_835,In_232);
or U912 (N_912,In_798,In_1232);
xnor U913 (N_913,In_624,In_1102);
xor U914 (N_914,In_1381,In_152);
nand U915 (N_915,In_968,In_1143);
nand U916 (N_916,In_2010,In_2258);
nand U917 (N_917,In_1391,In_1971);
and U918 (N_918,In_1896,In_437);
or U919 (N_919,In_1631,In_1873);
and U920 (N_920,In_1305,In_1862);
xor U921 (N_921,In_825,In_2002);
and U922 (N_922,In_1174,In_27);
nor U923 (N_923,In_2257,In_1027);
and U924 (N_924,In_1544,In_2007);
nand U925 (N_925,In_1618,In_863);
nor U926 (N_926,In_1270,In_1384);
nor U927 (N_927,In_2386,In_1853);
nor U928 (N_928,In_1211,In_424);
and U929 (N_929,In_1306,In_211);
nor U930 (N_930,In_501,In_1099);
nand U931 (N_931,In_1985,In_1298);
nor U932 (N_932,In_1168,In_902);
xor U933 (N_933,In_1828,In_1819);
nor U934 (N_934,In_965,In_2082);
nor U935 (N_935,In_247,In_954);
or U936 (N_936,In_1395,In_2463);
xor U937 (N_937,In_1876,In_56);
nor U938 (N_938,In_586,In_1447);
nor U939 (N_939,In_1716,In_1433);
or U940 (N_940,In_2209,In_1762);
nand U941 (N_941,In_78,In_1112);
and U942 (N_942,In_1098,In_1040);
and U943 (N_943,In_194,In_1625);
nand U944 (N_944,In_1379,In_765);
and U945 (N_945,In_1564,In_694);
or U946 (N_946,In_1339,In_1070);
xor U947 (N_947,In_281,In_2345);
and U948 (N_948,In_2067,In_594);
and U949 (N_949,In_275,In_2079);
and U950 (N_950,In_1894,In_2143);
and U951 (N_951,In_160,In_1811);
nor U952 (N_952,In_897,In_2332);
and U953 (N_953,In_2032,In_708);
and U954 (N_954,In_1382,In_1275);
nand U955 (N_955,In_1999,In_775);
or U956 (N_956,In_2481,In_2241);
and U957 (N_957,In_1080,In_2237);
or U958 (N_958,In_1778,In_333);
or U959 (N_959,In_2357,In_1284);
nand U960 (N_960,In_818,In_1990);
and U961 (N_961,In_1549,In_1909);
and U962 (N_962,In_1529,In_1086);
or U963 (N_963,In_604,In_1198);
xnor U964 (N_964,In_2159,In_304);
xnor U965 (N_965,In_2041,In_273);
nor U966 (N_966,In_1865,In_2321);
xnor U967 (N_967,In_753,In_1567);
and U968 (N_968,In_198,In_1935);
or U969 (N_969,In_1482,In_1463);
and U970 (N_970,In_730,In_221);
xnor U971 (N_971,In_648,In_1081);
nand U972 (N_972,In_1093,In_1257);
and U973 (N_973,In_481,In_704);
nor U974 (N_974,In_2282,In_2118);
and U975 (N_975,In_1231,In_559);
nand U976 (N_976,In_109,In_2275);
nor U977 (N_977,In_535,In_975);
nor U978 (N_978,In_100,In_451);
nand U979 (N_979,In_1570,In_2450);
xor U980 (N_980,In_1581,In_1368);
nor U981 (N_981,In_1771,In_994);
nand U982 (N_982,In_363,In_2200);
nand U983 (N_983,In_1252,In_2284);
nand U984 (N_984,In_707,In_399);
or U985 (N_985,In_2210,In_929);
or U986 (N_986,In_950,In_43);
nand U987 (N_987,In_66,In_1957);
xnor U988 (N_988,In_2169,In_1659);
xnor U989 (N_989,In_1937,In_983);
and U990 (N_990,In_612,In_963);
nand U991 (N_991,In_1171,In_1925);
or U992 (N_992,In_508,In_936);
xnor U993 (N_993,In_1361,In_88);
and U994 (N_994,In_2404,In_2365);
and U995 (N_995,In_1569,In_2397);
nand U996 (N_996,In_252,In_1097);
nand U997 (N_997,In_137,In_1881);
and U998 (N_998,In_1159,In_2053);
xor U999 (N_999,In_1964,In_736);
nand U1000 (N_1000,In_1557,In_711);
nor U1001 (N_1001,In_102,N_790);
nor U1002 (N_1002,In_1216,N_891);
nor U1003 (N_1003,N_888,In_674);
xor U1004 (N_1004,N_627,N_844);
or U1005 (N_1005,N_682,In_237);
and U1006 (N_1006,N_921,In_1153);
nand U1007 (N_1007,In_1558,N_135);
nor U1008 (N_1008,In_434,N_856);
or U1009 (N_1009,N_278,In_850);
nor U1010 (N_1010,N_807,N_557);
or U1011 (N_1011,N_541,N_897);
nor U1012 (N_1012,N_20,N_865);
nand U1013 (N_1013,N_753,N_591);
or U1014 (N_1014,N_518,N_637);
and U1015 (N_1015,In_1693,N_235);
or U1016 (N_1016,N_901,In_2311);
nor U1017 (N_1017,N_512,N_568);
and U1018 (N_1018,In_39,N_368);
xor U1019 (N_1019,N_130,N_413);
nand U1020 (N_1020,N_266,N_519);
nand U1021 (N_1021,N_462,N_800);
nand U1022 (N_1022,N_401,In_2065);
nor U1023 (N_1023,N_230,In_1722);
and U1024 (N_1024,N_767,N_970);
xnor U1025 (N_1025,In_402,In_1952);
or U1026 (N_1026,N_661,N_454);
xnor U1027 (N_1027,In_1965,N_995);
nand U1028 (N_1028,In_1733,N_62);
or U1029 (N_1029,N_811,N_678);
or U1030 (N_1030,N_525,N_314);
nor U1031 (N_1031,In_1050,In_2096);
and U1032 (N_1032,N_595,N_110);
xor U1033 (N_1033,In_1282,N_876);
nand U1034 (N_1034,N_23,N_480);
and U1035 (N_1035,N_258,In_740);
and U1036 (N_1036,N_468,In_638);
and U1037 (N_1037,In_558,N_744);
nor U1038 (N_1038,N_319,In_657);
xor U1039 (N_1039,N_727,In_849);
nand U1040 (N_1040,N_990,N_172);
xnor U1041 (N_1041,In_2091,In_2416);
nand U1042 (N_1042,N_108,N_329);
and U1043 (N_1043,N_4,N_833);
or U1044 (N_1044,In_1336,In_1547);
nand U1045 (N_1045,In_474,N_118);
or U1046 (N_1046,N_296,In_715);
and U1047 (N_1047,In_1736,N_26);
nand U1048 (N_1048,N_563,N_375);
nor U1049 (N_1049,N_244,N_789);
xor U1050 (N_1050,N_411,N_404);
xor U1051 (N_1051,N_30,N_873);
xor U1052 (N_1052,N_983,N_919);
and U1053 (N_1053,N_660,N_492);
nor U1054 (N_1054,In_1776,N_645);
nand U1055 (N_1055,N_561,N_605);
or U1056 (N_1056,In_1731,N_904);
and U1057 (N_1057,In_905,N_654);
and U1058 (N_1058,In_2149,In_1879);
nand U1059 (N_1059,N_500,N_201);
nand U1060 (N_1060,In_263,N_261);
or U1061 (N_1061,N_379,N_636);
nand U1062 (N_1062,N_128,N_883);
nand U1063 (N_1063,N_633,In_2028);
or U1064 (N_1064,In_278,N_885);
and U1065 (N_1065,In_0,N_305);
nand U1066 (N_1066,N_526,N_43);
xnor U1067 (N_1067,N_403,N_792);
and U1068 (N_1068,N_194,N_506);
and U1069 (N_1069,In_340,N_465);
nand U1070 (N_1070,N_24,In_1206);
and U1071 (N_1071,N_966,N_320);
nor U1072 (N_1072,N_618,N_560);
nor U1073 (N_1073,N_182,N_592);
or U1074 (N_1074,N_334,N_125);
nor U1075 (N_1075,N_298,In_62);
and U1076 (N_1076,N_429,In_347);
xnor U1077 (N_1077,N_324,N_700);
nand U1078 (N_1078,N_330,In_293);
or U1079 (N_1079,N_126,N_156);
xnor U1080 (N_1080,N_672,N_945);
nor U1081 (N_1081,N_496,In_2359);
or U1082 (N_1082,N_339,N_708);
or U1083 (N_1083,N_40,N_632);
nor U1084 (N_1084,N_940,N_750);
nor U1085 (N_1085,In_1826,In_2402);
and U1086 (N_1086,In_2268,N_388);
xnor U1087 (N_1087,N_609,N_655);
or U1088 (N_1088,In_2427,In_2360);
nand U1089 (N_1089,In_2036,In_1489);
xor U1090 (N_1090,In_189,N_279);
xnor U1091 (N_1091,N_529,N_674);
and U1092 (N_1092,N_651,N_692);
nand U1093 (N_1093,N_662,N_896);
and U1094 (N_1094,N_70,In_1651);
and U1095 (N_1095,In_1784,N_284);
or U1096 (N_1096,In_2499,N_817);
and U1097 (N_1097,N_819,In_565);
nor U1098 (N_1098,N_579,N_853);
or U1099 (N_1099,N_89,N_276);
or U1100 (N_1100,N_694,N_987);
nor U1101 (N_1101,N_504,N_162);
or U1102 (N_1102,In_600,N_301);
nor U1103 (N_1103,N_198,In_1609);
nand U1104 (N_1104,N_25,N_340);
nand U1105 (N_1105,N_976,N_48);
or U1106 (N_1106,N_470,In_322);
xnor U1107 (N_1107,N_378,N_313);
xor U1108 (N_1108,In_1135,N_345);
nand U1109 (N_1109,N_963,N_136);
and U1110 (N_1110,N_810,N_769);
xnor U1111 (N_1111,In_2239,N_507);
nor U1112 (N_1112,In_1923,N_559);
nor U1113 (N_1113,In_1079,In_1373);
nand U1114 (N_1114,N_912,N_606);
or U1115 (N_1115,N_780,N_881);
nor U1116 (N_1116,N_17,In_2111);
or U1117 (N_1117,N_497,In_1974);
nand U1118 (N_1118,N_782,N_797);
xnor U1119 (N_1119,N_836,N_570);
nand U1120 (N_1120,N_95,In_1812);
xnor U1121 (N_1121,N_300,N_240);
nor U1122 (N_1122,In_140,N_624);
nor U1123 (N_1123,N_15,In_1192);
xor U1124 (N_1124,N_845,N_505);
nand U1125 (N_1125,In_1094,N_285);
or U1126 (N_1126,N_770,In_904);
and U1127 (N_1127,N_486,N_181);
and U1128 (N_1128,N_688,N_806);
nor U1129 (N_1129,In_2198,N_850);
or U1130 (N_1130,In_2382,N_978);
nand U1131 (N_1131,N_848,In_1412);
nand U1132 (N_1132,N_151,N_446);
nand U1133 (N_1133,In_2130,In_1803);
and U1134 (N_1134,In_2325,N_835);
or U1135 (N_1135,N_880,N_170);
nor U1136 (N_1136,N_716,In_2207);
and U1137 (N_1137,N_996,In_310);
xor U1138 (N_1138,N_50,In_910);
nand U1139 (N_1139,N_527,N_703);
or U1140 (N_1140,In_2488,N_22);
nand U1141 (N_1141,In_1369,In_2142);
xor U1142 (N_1142,In_1841,In_1710);
nor U1143 (N_1143,N_635,In_1434);
xnor U1144 (N_1144,N_90,N_709);
nor U1145 (N_1145,N_416,In_933);
or U1146 (N_1146,In_1795,In_2407);
xor U1147 (N_1147,N_47,N_977);
nand U1148 (N_1148,In_839,N_209);
or U1149 (N_1149,N_696,N_701);
or U1150 (N_1150,In_599,In_81);
or U1151 (N_1151,N_517,N_450);
and U1152 (N_1152,N_31,N_88);
and U1153 (N_1153,N_357,N_493);
nor U1154 (N_1154,N_351,In_2231);
nand U1155 (N_1155,N_473,N_422);
xnor U1156 (N_1156,N_5,N_402);
and U1157 (N_1157,In_554,In_2155);
and U1158 (N_1158,N_166,In_292);
and U1159 (N_1159,N_653,N_268);
and U1160 (N_1160,In_801,N_697);
nor U1161 (N_1161,N_426,N_399);
nand U1162 (N_1162,N_167,N_575);
nand U1163 (N_1163,In_1314,N_537);
nor U1164 (N_1164,N_812,In_382);
xor U1165 (N_1165,N_36,N_202);
nor U1166 (N_1166,In_637,N_316);
or U1167 (N_1167,N_659,N_61);
or U1168 (N_1168,In_2152,N_117);
nor U1169 (N_1169,N_231,In_121);
and U1170 (N_1170,N_488,N_720);
xor U1171 (N_1171,N_628,In_54);
nor U1172 (N_1172,N_347,In_2047);
nor U1173 (N_1173,N_225,N_93);
xor U1174 (N_1174,N_864,N_287);
nand U1175 (N_1175,N_951,N_142);
xnor U1176 (N_1176,N_207,N_430);
xor U1177 (N_1177,N_299,N_155);
nand U1178 (N_1178,N_91,N_359);
nor U1179 (N_1179,N_362,N_304);
or U1180 (N_1180,N_915,N_262);
xor U1181 (N_1181,N_482,In_1415);
nand U1182 (N_1182,N_171,In_250);
xnor U1183 (N_1183,In_930,In_1160);
nor U1184 (N_1184,N_216,N_926);
and U1185 (N_1185,N_221,N_754);
nand U1186 (N_1186,N_373,In_1142);
nor U1187 (N_1187,N_523,N_736);
and U1188 (N_1188,N_86,In_406);
or U1189 (N_1189,N_867,In_1607);
or U1190 (N_1190,N_711,N_639);
and U1191 (N_1191,N_327,N_311);
nand U1192 (N_1192,In_1347,N_157);
or U1193 (N_1193,N_874,In_1582);
nand U1194 (N_1194,N_94,In_1987);
or U1195 (N_1195,N_342,In_1589);
xnor U1196 (N_1196,In_1946,In_317);
or U1197 (N_1197,N_478,N_842);
xnor U1198 (N_1198,N_431,N_796);
nand U1199 (N_1199,N_228,N_690);
xor U1200 (N_1200,N_710,N_163);
nor U1201 (N_1201,In_239,N_712);
or U1202 (N_1202,N_719,N_116);
or U1203 (N_1203,N_409,N_617);
nand U1204 (N_1204,N_747,N_589);
and U1205 (N_1205,N_944,In_1505);
xnor U1206 (N_1206,N_365,N_367);
xor U1207 (N_1207,N_161,N_755);
nor U1208 (N_1208,N_18,N_177);
nand U1209 (N_1209,In_2033,N_0);
nand U1210 (N_1210,N_81,In_1105);
nor U1211 (N_1211,N_799,N_732);
or U1212 (N_1212,In_2490,N_415);
nand U1213 (N_1213,N_728,In_139);
or U1214 (N_1214,In_2412,In_2384);
nor U1215 (N_1215,N_100,N_994);
and U1216 (N_1216,N_918,In_1910);
xnor U1217 (N_1217,In_1150,N_997);
and U1218 (N_1218,N_457,In_1695);
and U1219 (N_1219,N_964,N_937);
xor U1220 (N_1220,N_626,N_286);
nand U1221 (N_1221,In_1241,N_607);
or U1222 (N_1222,In_577,In_1250);
or U1223 (N_1223,In_461,In_2046);
and U1224 (N_1224,N_993,In_1356);
nor U1225 (N_1225,N_691,N_869);
nor U1226 (N_1226,N_543,N_369);
nor U1227 (N_1227,N_585,N_818);
and U1228 (N_1228,N_272,In_2174);
nand U1229 (N_1229,N_393,N_603);
xnor U1230 (N_1230,In_995,N_449);
or U1231 (N_1231,In_1028,N_913);
or U1232 (N_1232,N_364,In_1644);
nand U1233 (N_1233,In_645,N_890);
nand U1234 (N_1234,N_290,N_948);
xnor U1235 (N_1235,N_785,N_586);
nand U1236 (N_1236,In_192,In_280);
or U1237 (N_1237,In_2422,In_1866);
nor U1238 (N_1238,N_427,In_1583);
xnor U1239 (N_1239,In_633,N_2);
xnor U1240 (N_1240,N_600,In_749);
and U1241 (N_1241,N_707,N_619);
xnor U1242 (N_1242,N_148,In_951);
nor U1243 (N_1243,In_621,In_2317);
nand U1244 (N_1244,In_1741,In_346);
or U1245 (N_1245,N_571,N_562);
nand U1246 (N_1246,In_855,In_946);
nand U1247 (N_1247,In_2358,N_650);
nor U1248 (N_1248,N_631,In_343);
and U1249 (N_1249,N_573,N_693);
and U1250 (N_1250,N_21,N_992);
nor U1251 (N_1251,N_882,In_2218);
and U1252 (N_1252,In_2248,N_494);
nor U1253 (N_1253,N_657,N_787);
xor U1254 (N_1254,N_9,In_1871);
and U1255 (N_1255,In_955,In_320);
xor U1256 (N_1256,N_933,In_138);
and U1257 (N_1257,N_957,N_795);
xor U1258 (N_1258,In_669,N_137);
nor U1259 (N_1259,N_676,In_608);
and U1260 (N_1260,N_434,N_82);
xor U1261 (N_1261,N_621,N_67);
and U1262 (N_1262,N_140,N_777);
or U1263 (N_1263,In_1036,In_466);
and U1264 (N_1264,In_859,In_2071);
xor U1265 (N_1265,N_699,In_476);
nand U1266 (N_1266,N_28,N_695);
or U1267 (N_1267,In_1848,In_1608);
nand U1268 (N_1268,In_1880,N_16);
nand U1269 (N_1269,N_932,N_341);
xnor U1270 (N_1270,In_200,In_868);
or U1271 (N_1271,N_555,N_574);
or U1272 (N_1272,In_1271,N_802);
or U1273 (N_1273,In_1515,In_429);
or U1274 (N_1274,N_849,N_54);
nand U1275 (N_1275,N_12,In_1121);
nand U1276 (N_1276,In_1789,In_394);
xor U1277 (N_1277,N_510,N_927);
or U1278 (N_1278,N_337,N_294);
xor U1279 (N_1279,In_1883,N_255);
xnor U1280 (N_1280,In_2383,In_1833);
nand U1281 (N_1281,N_804,N_303);
nand U1282 (N_1282,In_2424,N_269);
nand U1283 (N_1283,N_721,In_126);
xor U1284 (N_1284,N_545,N_476);
xor U1285 (N_1285,In_799,N_752);
or U1286 (N_1286,N_98,In_2183);
nor U1287 (N_1287,N_121,N_929);
nor U1288 (N_1288,In_1572,N_950);
nand U1289 (N_1289,N_96,N_58);
or U1290 (N_1290,N_200,N_165);
nand U1291 (N_1291,N_734,N_217);
nand U1292 (N_1292,In_1315,N_490);
xnor U1293 (N_1293,N_863,N_946);
or U1294 (N_1294,N_936,N_572);
or U1295 (N_1295,N_238,N_291);
nand U1296 (N_1296,N_213,N_312);
nor U1297 (N_1297,In_576,N_798);
or U1298 (N_1298,In_761,N_514);
or U1299 (N_1299,N_197,N_613);
or U1300 (N_1300,N_513,N_698);
nand U1301 (N_1301,N_870,N_39);
or U1302 (N_1302,In_1119,N_872);
xor U1303 (N_1303,N_566,N_19);
nand U1304 (N_1304,N_593,N_421);
xnor U1305 (N_1305,N_596,N_689);
and U1306 (N_1306,N_743,In_812);
and U1307 (N_1307,N_778,N_159);
nand U1308 (N_1308,In_2309,N_467);
nand U1309 (N_1309,In_2437,In_1972);
xnor U1310 (N_1310,N_243,N_899);
and U1311 (N_1311,In_591,In_2019);
nand U1312 (N_1312,N_952,N_361);
or U1313 (N_1313,N_920,In_1749);
xnor U1314 (N_1314,In_30,In_1141);
or U1315 (N_1315,N_939,N_111);
nand U1316 (N_1316,In_960,N_60);
xor U1317 (N_1317,N_986,N_14);
and U1318 (N_1318,In_1318,N_544);
nand U1319 (N_1319,In_462,N_99);
xor U1320 (N_1320,In_1630,N_71);
nor U1321 (N_1321,In_1531,N_671);
and U1322 (N_1322,In_380,N_644);
and U1323 (N_1323,In_1556,N_847);
or U1324 (N_1324,N_590,N_828);
or U1325 (N_1325,N_335,N_214);
nand U1326 (N_1326,N_717,N_179);
or U1327 (N_1327,N_975,In_1626);
xnor U1328 (N_1328,N_775,N_914);
or U1329 (N_1329,N_332,In_523);
nor U1330 (N_1330,N_532,In_2396);
nand U1331 (N_1331,N_190,In_634);
nand U1332 (N_1332,In_385,N_158);
and U1333 (N_1333,N_348,In_1714);
or U1334 (N_1334,N_793,N_400);
nor U1335 (N_1335,N_75,In_1283);
or U1336 (N_1336,N_229,N_134);
and U1337 (N_1337,N_569,In_872);
nor U1338 (N_1338,N_471,N_124);
or U1339 (N_1339,In_1757,N_176);
or U1340 (N_1340,N_540,N_178);
nor U1341 (N_1341,In_1824,In_629);
and U1342 (N_1342,N_281,In_1566);
nand U1343 (N_1343,In_827,N_938);
nand U1344 (N_1344,In_562,N_396);
nand U1345 (N_1345,In_2043,In_1132);
nand U1346 (N_1346,In_873,In_1120);
or U1347 (N_1347,N_212,N_909);
and U1348 (N_1348,In_1479,N_251);
xnor U1349 (N_1349,N_3,In_312);
and U1350 (N_1350,N_681,N_664);
and U1351 (N_1351,N_702,N_270);
xor U1352 (N_1352,In_1653,N_822);
or U1353 (N_1353,N_538,N_398);
xor U1354 (N_1354,N_346,N_580);
nor U1355 (N_1355,N_11,N_855);
or U1356 (N_1356,N_192,In_811);
nor U1357 (N_1357,N_455,In_1204);
or U1358 (N_1358,N_677,N_784);
nand U1359 (N_1359,N_981,In_941);
nor U1360 (N_1360,N_508,N_680);
or U1361 (N_1361,In_1968,N_223);
or U1362 (N_1362,In_655,N_826);
xor U1363 (N_1363,N_109,In_1471);
xor U1364 (N_1364,In_1553,N_612);
nor U1365 (N_1365,N_491,N_218);
nand U1366 (N_1366,N_406,N_634);
xnor U1367 (N_1367,N_961,In_2208);
and U1368 (N_1368,N_683,N_308);
xor U1369 (N_1369,In_838,N_168);
or U1370 (N_1370,In_546,In_1533);
nand U1371 (N_1371,In_1773,In_1390);
and U1372 (N_1372,N_420,N_353);
xor U1373 (N_1373,N_239,N_382);
or U1374 (N_1374,N_955,In_2451);
nor U1375 (N_1375,N_935,N_999);
xnor U1376 (N_1376,In_712,N_153);
or U1377 (N_1377,In_300,N_760);
and U1378 (N_1378,N_588,N_419);
and U1379 (N_1379,N_295,N_412);
nand U1380 (N_1380,In_1398,N_911);
nand U1381 (N_1381,In_1405,N_271);
and U1382 (N_1382,N_943,In_1133);
or U1383 (N_1383,N_601,N_722);
nand U1384 (N_1384,N_57,N_791);
or U1385 (N_1385,N_174,N_843);
and U1386 (N_1386,In_698,In_787);
and U1387 (N_1387,N_587,In_2034);
nand U1388 (N_1388,In_1155,N_437);
nand U1389 (N_1389,In_1764,In_792);
nor U1390 (N_1390,N_112,N_73);
and U1391 (N_1391,In_2201,N_499);
nand U1392 (N_1392,N_37,N_428);
nand U1393 (N_1393,In_1172,In_18);
and U1394 (N_1394,N_803,In_2250);
xnor U1395 (N_1395,N_852,N_831);
nor U1396 (N_1396,In_1115,N_448);
nor U1397 (N_1397,N_38,In_42);
and U1398 (N_1398,N_851,N_495);
nor U1399 (N_1399,N_355,In_497);
and U1400 (N_1400,N_289,N_610);
or U1401 (N_1401,In_1140,In_823);
xor U1402 (N_1402,In_1912,N_321);
xnor U1403 (N_1403,N_27,In_1527);
xnor U1404 (N_1404,In_2254,In_1461);
xor U1405 (N_1405,In_1874,In_758);
xnor U1406 (N_1406,In_550,N_139);
nand U1407 (N_1407,In_803,N_718);
or U1408 (N_1408,N_854,N_264);
xor U1409 (N_1409,In_702,N_907);
xnor U1410 (N_1410,N_141,N_199);
xnor U1411 (N_1411,N_418,N_928);
and U1412 (N_1412,In_2101,N_887);
xor U1413 (N_1413,N_878,N_840);
nand U1414 (N_1414,N_42,N_224);
and U1415 (N_1415,N_147,In_1309);
nor U1416 (N_1416,N_673,In_1317);
nor U1417 (N_1417,In_828,N_438);
or U1418 (N_1418,In_1884,N_834);
or U1419 (N_1419,N_175,N_931);
xnor U1420 (N_1420,N_889,N_539);
and U1421 (N_1421,In_50,N_759);
nor U1422 (N_1422,N_577,N_83);
nand U1423 (N_1423,N_80,N_528);
nand U1424 (N_1424,In_2304,N_247);
nor U1425 (N_1425,N_389,In_1530);
nor U1426 (N_1426,In_181,In_1386);
nor U1427 (N_1427,In_396,N_556);
nand U1428 (N_1428,In_703,In_2415);
and U1429 (N_1429,N_530,N_275);
nand U1430 (N_1430,N_248,N_253);
nand U1431 (N_1431,N_667,In_452);
nand U1432 (N_1432,In_427,In_673);
nor U1433 (N_1433,N_726,N_805);
xnor U1434 (N_1434,N_705,N_184);
nor U1435 (N_1435,N_485,N_594);
xor U1436 (N_1436,In_518,N_622);
xor U1437 (N_1437,N_511,N_860);
or U1438 (N_1438,In_1670,N_646);
and U1439 (N_1439,In_1649,N_922);
xor U1440 (N_1440,N_129,N_971);
nand U1441 (N_1441,N_322,N_267);
and U1442 (N_1442,N_443,N_547);
nor U1443 (N_1443,N_232,N_598);
and U1444 (N_1444,In_543,In_1914);
xnor U1445 (N_1445,In_1292,In_1735);
xor U1446 (N_1446,N_452,N_105);
or U1447 (N_1447,N_503,In_235);
nor U1448 (N_1448,In_1791,N_392);
nand U1449 (N_1449,N_871,In_578);
xor U1450 (N_1450,In_177,N_858);
and U1451 (N_1451,N_783,N_64);
or U1452 (N_1452,N_991,In_684);
xor U1453 (N_1453,In_2310,N_808);
nor U1454 (N_1454,N_260,N_830);
nor U1455 (N_1455,N_735,N_445);
or U1456 (N_1456,In_1358,N_10);
nand U1457 (N_1457,N_788,N_820);
or U1458 (N_1458,N_256,N_730);
xnor U1459 (N_1459,N_669,In_101);
and U1460 (N_1460,N_832,In_907);
or U1461 (N_1461,N_466,N_829);
or U1462 (N_1462,In_1683,N_567);
nand U1463 (N_1463,In_1428,In_611);
and U1464 (N_1464,N_280,N_8);
xor U1465 (N_1465,N_620,In_1033);
and U1466 (N_1466,In_415,In_2050);
or U1467 (N_1467,N_502,In_125);
xnor U1468 (N_1468,N_114,N_647);
xnor U1469 (N_1469,N_704,N_461);
and U1470 (N_1470,N_824,N_46);
xor U1471 (N_1471,In_342,In_887);
xor U1472 (N_1472,N_293,In_1312);
nand U1473 (N_1473,N_953,N_917);
or U1474 (N_1474,In_723,N_738);
or U1475 (N_1475,N_87,N_962);
or U1476 (N_1476,In_743,N_522);
nor U1477 (N_1477,In_1932,In_379);
or U1478 (N_1478,In_1350,N_7);
nor U1479 (N_1479,In_999,N_906);
and U1480 (N_1480,In_1338,N_273);
xnor U1481 (N_1481,In_1930,N_297);
and U1482 (N_1482,In_1016,N_552);
and U1483 (N_1483,N_424,N_998);
xor U1484 (N_1484,In_1934,In_510);
or U1485 (N_1485,N_183,N_63);
and U1486 (N_1486,N_186,N_751);
nor U1487 (N_1487,N_436,In_2380);
xor U1488 (N_1488,In_1436,N_742);
or U1489 (N_1489,In_1503,N_959);
xnor U1490 (N_1490,N_154,N_447);
xor U1491 (N_1491,In_1138,N_241);
or U1492 (N_1492,N_469,N_180);
and U1493 (N_1493,N_45,N_122);
nor U1494 (N_1494,In_1151,N_144);
or U1495 (N_1495,N_942,N_59);
and U1496 (N_1496,N_684,In_697);
nand U1497 (N_1497,N_766,N_435);
or U1498 (N_1498,N_219,N_638);
and U1499 (N_1499,N_282,N_456);
or U1500 (N_1500,N_553,N_69);
xnor U1501 (N_1501,N_227,In_440);
xor U1502 (N_1502,N_685,N_827);
nor U1503 (N_1503,N_772,N_648);
xor U1504 (N_1504,N_371,N_226);
nor U1505 (N_1505,N_894,N_516);
or U1506 (N_1506,In_16,N_756);
or U1507 (N_1507,In_1610,N_85);
nor U1508 (N_1508,N_97,In_470);
xor U1509 (N_1509,N_924,N_774);
xnor U1510 (N_1510,N_947,N_386);
or U1511 (N_1511,N_823,N_484);
xor U1512 (N_1512,N_895,In_400);
or U1513 (N_1513,N_551,N_686);
xor U1514 (N_1514,N_614,N_602);
nor U1515 (N_1515,In_1055,In_777);
nand U1516 (N_1516,In_1002,N_576);
nand U1517 (N_1517,N_210,In_1782);
and U1518 (N_1518,N_123,In_2172);
or U1519 (N_1519,In_998,In_603);
nand U1520 (N_1520,N_724,In_635);
or U1521 (N_1521,In_83,N_414);
xor U1522 (N_1522,N_193,N_1);
nand U1523 (N_1523,In_2102,N_862);
and U1524 (N_1524,N_444,N_509);
xnor U1525 (N_1525,N_363,In_747);
or U1526 (N_1526,In_158,N_250);
and U1527 (N_1527,N_344,N_127);
xor U1528 (N_1528,N_611,N_625);
or U1529 (N_1529,In_592,In_957);
nor U1530 (N_1530,N_548,In_597);
xnor U1531 (N_1531,N_908,N_733);
nand U1532 (N_1532,In_606,N_41);
xor U1533 (N_1533,N_374,N_13);
nand U1534 (N_1534,In_853,In_1295);
and U1535 (N_1535,N_149,N_6);
xor U1536 (N_1536,In_1030,In_2319);
and U1537 (N_1537,N_809,N_630);
nand U1538 (N_1538,N_879,N_326);
nor U1539 (N_1539,N_546,N_934);
or U1540 (N_1540,In_366,N_930);
or U1541 (N_1541,In_1452,N_816);
nand U1542 (N_1542,In_2432,N_839);
nand U1543 (N_1543,N_453,In_1845);
xor U1544 (N_1544,In_2115,N_323);
nand U1545 (N_1545,N_211,N_658);
nand U1546 (N_1546,In_2334,In_301);
nand U1547 (N_1547,In_1636,N_338);
or U1548 (N_1548,N_115,N_582);
or U1549 (N_1549,N_318,N_259);
or U1550 (N_1550,In_717,In_2061);
or U1551 (N_1551,N_973,N_150);
or U1552 (N_1552,N_536,N_336);
nor U1553 (N_1553,In_212,N_520);
xnor U1554 (N_1554,N_615,In_1032);
or U1555 (N_1555,N_665,N_533);
nand U1556 (N_1556,N_395,In_682);
or U1557 (N_1557,N_66,In_2070);
or U1558 (N_1558,In_480,In_163);
or U1559 (N_1559,N_670,N_283);
and U1560 (N_1560,In_1639,N_35);
and U1561 (N_1561,N_106,N_203);
nand U1562 (N_1562,N_643,N_394);
nor U1563 (N_1563,In_2175,N_425);
nor U1564 (N_1564,In_13,In_1684);
nand U1565 (N_1565,In_225,N_958);
and U1566 (N_1566,In_1751,In_613);
nand U1567 (N_1567,In_2285,In_2498);
xor U1568 (N_1568,In_359,N_196);
and U1569 (N_1569,N_846,N_234);
nor U1570 (N_1570,N_49,In_1178);
or U1571 (N_1571,N_898,In_161);
nor U1572 (N_1572,N_739,In_1906);
nand U1573 (N_1573,N_352,N_145);
nor U1574 (N_1574,N_813,N_220);
nor U1575 (N_1575,In_533,In_847);
xnor U1576 (N_1576,N_309,N_185);
and U1577 (N_1577,N_474,N_965);
nor U1578 (N_1578,In_1457,N_206);
or U1579 (N_1579,N_310,N_55);
nand U1580 (N_1580,In_1697,N_815);
xor U1581 (N_1581,N_152,In_355);
and U1582 (N_1582,In_368,N_746);
xnor U1583 (N_1583,N_941,In_972);
nor U1584 (N_1584,N_679,In_1679);
nand U1585 (N_1585,In_580,N_472);
xor U1586 (N_1586,In_2253,N_460);
xor U1587 (N_1587,N_745,N_34);
and U1588 (N_1588,In_287,N_169);
and U1589 (N_1589,In_509,In_931);
nand U1590 (N_1590,N_838,N_902);
nor U1591 (N_1591,N_479,N_903);
or U1592 (N_1592,N_408,N_758);
and U1593 (N_1593,N_113,N_53);
and U1594 (N_1594,N_663,In_144);
nor U1595 (N_1595,In_1223,N_354);
xor U1596 (N_1596,N_417,N_980);
or U1597 (N_1597,In_1574,N_246);
and U1598 (N_1598,N_988,In_1212);
nand U1599 (N_1599,N_133,In_1432);
nand U1600 (N_1600,N_236,In_952);
nor U1601 (N_1601,In_389,N_954);
nor U1602 (N_1602,N_349,N_102);
nor U1603 (N_1603,In_751,N_265);
xor U1604 (N_1604,N_749,N_328);
and U1605 (N_1605,N_101,N_498);
xnor U1606 (N_1606,In_1619,N_967);
and U1607 (N_1607,N_565,N_549);
nand U1608 (N_1608,N_410,N_441);
xor U1609 (N_1609,N_208,N_877);
and U1610 (N_1610,N_252,N_825);
xnor U1611 (N_1611,In_1085,N_771);
nor U1612 (N_1612,N_857,In_2227);
nor U1613 (N_1613,In_516,In_709);
nor U1614 (N_1614,N_188,N_288);
xnor U1615 (N_1615,In_1090,N_731);
xnor U1616 (N_1616,In_450,N_979);
and U1617 (N_1617,N_173,N_531);
xor U1618 (N_1618,N_583,N_306);
and U1619 (N_1619,N_866,N_376);
and U1620 (N_1620,N_925,N_761);
nand U1621 (N_1621,N_432,In_443);
xnor U1622 (N_1622,N_315,In_557);
and U1623 (N_1623,N_187,N_765);
nand U1624 (N_1624,N_68,In_1000);
xor U1625 (N_1625,N_558,N_103);
or U1626 (N_1626,N_956,N_554);
xnor U1627 (N_1627,N_652,In_20);
nand U1628 (N_1628,N_343,N_76);
or U1629 (N_1629,N_52,In_2279);
xnor U1630 (N_1630,N_960,In_94);
nor U1631 (N_1631,In_1526,N_263);
nor U1632 (N_1632,N_56,N_892);
nor U1633 (N_1633,In_984,In_244);
nor U1634 (N_1634,N_706,N_143);
xor U1635 (N_1635,N_464,N_249);
or U1636 (N_1636,In_283,N_762);
and U1637 (N_1637,N_542,N_477);
xnor U1638 (N_1638,In_1908,N_292);
xnor U1639 (N_1639,N_779,N_74);
and U1640 (N_1640,N_277,N_515);
or U1641 (N_1641,N_77,In_410);
and U1642 (N_1642,In_1961,N_675);
and U1643 (N_1643,N_741,N_385);
or U1644 (N_1644,N_668,In_2166);
and U1645 (N_1645,In_911,N_475);
and U1646 (N_1646,N_764,In_55);
nor U1647 (N_1647,N_160,N_215);
xor U1648 (N_1648,N_302,In_665);
nor U1649 (N_1649,In_113,N_985);
nor U1650 (N_1650,In_2418,N_968);
and U1651 (N_1651,N_146,In_338);
nor U1652 (N_1652,N_687,N_245);
nor U1653 (N_1653,N_274,In_856);
xnor U1654 (N_1654,N_642,N_821);
xnor U1655 (N_1655,N_459,N_905);
xnor U1656 (N_1656,N_768,N_974);
and U1657 (N_1657,N_360,N_381);
nor U1658 (N_1658,N_715,N_32);
nor U1659 (N_1659,In_2204,N_725);
nand U1660 (N_1660,N_358,N_900);
or U1661 (N_1661,N_623,In_85);
and U1662 (N_1662,N_550,In_2491);
nor U1663 (N_1663,N_205,N_489);
or U1664 (N_1664,N_483,N_781);
nand U1665 (N_1665,N_923,N_372);
and U1666 (N_1666,N_984,In_1184);
xnor U1667 (N_1667,N_104,N_597);
or U1668 (N_1668,N_317,N_629);
or U1669 (N_1669,N_723,In_1321);
xnor U1670 (N_1670,N_189,N_640);
or U1671 (N_1671,In_661,N_501);
and U1672 (N_1672,In_441,N_407);
xnor U1673 (N_1673,N_79,In_1001);
or U1674 (N_1674,N_578,N_729);
nor U1675 (N_1675,N_786,N_439);
or U1676 (N_1676,In_1245,In_2230);
nand U1677 (N_1677,N_307,N_33);
xor U1678 (N_1678,N_72,In_187);
nor U1679 (N_1679,In_1082,In_2440);
xnor U1680 (N_1680,N_748,N_969);
nor U1681 (N_1681,N_132,N_814);
nand U1682 (N_1682,N_195,In_1096);
and U1683 (N_1683,In_996,In_1750);
nor U1684 (N_1684,In_1513,N_331);
or U1685 (N_1685,In_1238,N_366);
nor U1686 (N_1686,N_29,N_383);
and U1687 (N_1687,N_656,In_2024);
and U1688 (N_1688,N_972,In_1545);
xnor U1689 (N_1689,N_390,N_801);
nand U1690 (N_1690,N_458,N_191);
nand U1691 (N_1691,N_604,N_616);
nand U1692 (N_1692,In_425,In_120);
and U1693 (N_1693,In_365,In_837);
and U1694 (N_1694,In_1400,In_1868);
xor U1695 (N_1695,In_1510,In_1169);
and U1696 (N_1696,N_92,N_666);
nor U1697 (N_1697,N_325,N_773);
and U1698 (N_1698,N_237,In_1715);
nor U1699 (N_1699,In_115,In_2367);
and U1700 (N_1700,N_776,N_442);
nor U1701 (N_1701,N_916,In_2148);
and U1702 (N_1702,In_1087,In_1188);
nand U1703 (N_1703,N_44,N_204);
or U1704 (N_1704,N_599,N_451);
xnor U1705 (N_1705,N_982,In_2202);
nor U1706 (N_1706,N_841,N_763);
or U1707 (N_1707,N_254,N_584);
or U1708 (N_1708,In_739,In_2303);
xor U1709 (N_1709,N_440,N_910);
and U1710 (N_1710,N_138,In_549);
or U1711 (N_1711,N_222,N_463);
and U1712 (N_1712,N_164,In_660);
nand U1713 (N_1713,N_740,N_405);
nand U1714 (N_1714,N_884,N_131);
or U1715 (N_1715,In_1535,N_257);
xnor U1716 (N_1716,In_1637,N_649);
and U1717 (N_1717,N_356,In_1233);
xor U1718 (N_1718,N_868,N_608);
or U1719 (N_1719,N_886,N_534);
nor U1720 (N_1720,N_242,In_1351);
and U1721 (N_1721,N_65,In_259);
or U1722 (N_1722,N_859,N_119);
or U1723 (N_1723,In_1066,In_1806);
xnor U1724 (N_1724,N_949,N_794);
xnor U1725 (N_1725,In_620,N_387);
xnor U1726 (N_1726,N_233,N_333);
or U1727 (N_1727,N_893,N_875);
or U1728 (N_1728,N_84,N_989);
xor U1729 (N_1729,N_350,N_713);
xnor U1730 (N_1730,In_2223,N_120);
nand U1731 (N_1731,N_397,N_521);
xnor U1732 (N_1732,N_535,N_737);
nand U1733 (N_1733,In_886,N_78);
or U1734 (N_1734,N_641,In_1374);
and U1735 (N_1735,N_714,N_423);
xnor U1736 (N_1736,N_581,N_107);
or U1737 (N_1737,In_1730,N_51);
or U1738 (N_1738,In_2049,N_524);
xor U1739 (N_1739,In_2086,N_384);
nor U1740 (N_1740,N_837,In_2080);
nor U1741 (N_1741,N_487,N_380);
nand U1742 (N_1742,In_652,N_861);
xor U1743 (N_1743,In_4,In_1483);
nand U1744 (N_1744,N_481,N_370);
or U1745 (N_1745,N_757,In_769);
nand U1746 (N_1746,N_377,In_1328);
nand U1747 (N_1747,N_433,In_1685);
and U1748 (N_1748,N_391,In_1616);
nor U1749 (N_1749,In_764,N_564);
or U1750 (N_1750,N_131,N_814);
and U1751 (N_1751,N_154,In_102);
xor U1752 (N_1752,N_159,N_552);
nand U1753 (N_1753,In_1866,N_646);
or U1754 (N_1754,N_902,N_243);
xor U1755 (N_1755,N_783,N_444);
nand U1756 (N_1756,N_779,N_879);
nor U1757 (N_1757,N_532,N_909);
nand U1758 (N_1758,In_239,N_996);
nor U1759 (N_1759,N_266,In_2218);
or U1760 (N_1760,N_784,N_348);
nand U1761 (N_1761,N_617,N_916);
or U1762 (N_1762,In_2382,In_1582);
nand U1763 (N_1763,In_577,N_656);
or U1764 (N_1764,N_474,N_174);
nand U1765 (N_1765,N_936,N_952);
and U1766 (N_1766,N_293,N_960);
or U1767 (N_1767,N_895,N_474);
nand U1768 (N_1768,N_504,N_937);
and U1769 (N_1769,N_223,N_420);
nand U1770 (N_1770,N_488,N_987);
and U1771 (N_1771,In_1757,In_1515);
nand U1772 (N_1772,N_335,In_2142);
nor U1773 (N_1773,N_16,N_914);
nor U1774 (N_1774,N_820,N_903);
nor U1775 (N_1775,N_806,In_2130);
xor U1776 (N_1776,N_745,N_872);
xor U1777 (N_1777,N_251,In_1412);
and U1778 (N_1778,N_804,In_1751);
nor U1779 (N_1779,In_225,N_781);
or U1780 (N_1780,N_848,N_970);
nand U1781 (N_1781,In_1483,In_300);
xor U1782 (N_1782,N_402,N_835);
and U1783 (N_1783,In_2279,In_709);
nor U1784 (N_1784,N_411,N_740);
nor U1785 (N_1785,N_956,N_899);
xor U1786 (N_1786,N_719,N_578);
xnor U1787 (N_1787,N_633,N_309);
and U1788 (N_1788,N_107,In_1908);
nor U1789 (N_1789,In_557,N_127);
xnor U1790 (N_1790,N_431,N_407);
or U1791 (N_1791,In_1776,In_1153);
nand U1792 (N_1792,In_717,N_219);
nand U1793 (N_1793,N_224,In_1649);
or U1794 (N_1794,N_581,In_907);
nor U1795 (N_1795,In_1685,N_173);
nor U1796 (N_1796,In_702,N_985);
and U1797 (N_1797,N_620,In_1952);
or U1798 (N_1798,In_1055,N_916);
xor U1799 (N_1799,N_287,In_1412);
or U1800 (N_1800,N_842,N_220);
nand U1801 (N_1801,N_327,N_371);
nand U1802 (N_1802,N_74,In_1557);
xor U1803 (N_1803,N_411,In_2309);
nand U1804 (N_1804,N_728,N_280);
xnor U1805 (N_1805,N_870,In_2319);
xor U1806 (N_1806,N_343,N_220);
and U1807 (N_1807,N_547,N_858);
and U1808 (N_1808,In_126,N_938);
nor U1809 (N_1809,N_824,N_404);
nand U1810 (N_1810,N_937,In_2202);
xor U1811 (N_1811,N_65,N_431);
nor U1812 (N_1812,In_2227,N_366);
and U1813 (N_1813,In_1094,N_136);
and U1814 (N_1814,N_363,In_657);
nand U1815 (N_1815,N_554,N_378);
xnor U1816 (N_1816,N_105,N_652);
nand U1817 (N_1817,N_658,N_646);
or U1818 (N_1818,N_163,In_1412);
xor U1819 (N_1819,N_313,N_743);
or U1820 (N_1820,N_316,In_2499);
or U1821 (N_1821,In_394,In_955);
or U1822 (N_1822,N_110,N_852);
or U1823 (N_1823,In_847,N_706);
nand U1824 (N_1824,N_767,N_163);
nor U1825 (N_1825,N_289,N_683);
xnor U1826 (N_1826,N_991,In_2498);
nor U1827 (N_1827,N_6,N_474);
nand U1828 (N_1828,N_417,N_501);
or U1829 (N_1829,In_1358,In_603);
or U1830 (N_1830,In_597,N_467);
xor U1831 (N_1831,In_1115,N_552);
xor U1832 (N_1832,N_631,N_947);
and U1833 (N_1833,In_712,In_400);
or U1834 (N_1834,N_182,N_101);
and U1835 (N_1835,N_560,N_94);
or U1836 (N_1836,In_1773,N_368);
or U1837 (N_1837,N_366,In_1735);
or U1838 (N_1838,In_578,N_902);
or U1839 (N_1839,N_315,In_42);
or U1840 (N_1840,N_368,N_713);
or U1841 (N_1841,N_508,N_736);
and U1842 (N_1842,N_44,N_839);
or U1843 (N_1843,N_451,N_542);
and U1844 (N_1844,N_807,In_1515);
nor U1845 (N_1845,In_2166,N_398);
nor U1846 (N_1846,N_164,N_381);
or U1847 (N_1847,In_1282,In_715);
nor U1848 (N_1848,In_887,In_855);
and U1849 (N_1849,In_380,N_962);
or U1850 (N_1850,N_143,N_430);
xnor U1851 (N_1851,In_787,In_1636);
or U1852 (N_1852,N_640,In_382);
and U1853 (N_1853,In_1292,N_901);
and U1854 (N_1854,In_1530,N_332);
nand U1855 (N_1855,In_1968,N_33);
or U1856 (N_1856,N_193,In_2309);
xnor U1857 (N_1857,In_697,N_620);
xor U1858 (N_1858,In_50,N_575);
or U1859 (N_1859,In_1241,N_456);
xnor U1860 (N_1860,N_80,N_550);
xnor U1861 (N_1861,In_1735,N_82);
and U1862 (N_1862,N_456,In_338);
or U1863 (N_1863,N_540,In_1946);
or U1864 (N_1864,N_143,N_497);
or U1865 (N_1865,N_6,N_680);
and U1866 (N_1866,In_2034,N_432);
xnor U1867 (N_1867,In_177,N_787);
or U1868 (N_1868,In_2248,In_1733);
xor U1869 (N_1869,N_496,N_961);
and U1870 (N_1870,N_214,N_48);
and U1871 (N_1871,In_85,In_2086);
and U1872 (N_1872,N_899,N_303);
and U1873 (N_1873,In_1347,In_2440);
xor U1874 (N_1874,N_730,N_527);
nand U1875 (N_1875,N_605,In_2047);
and U1876 (N_1876,In_410,In_1216);
xnor U1877 (N_1877,N_893,N_507);
nor U1878 (N_1878,In_342,N_951);
nand U1879 (N_1879,N_237,N_111);
and U1880 (N_1880,In_1295,In_2142);
xnor U1881 (N_1881,N_889,In_1946);
or U1882 (N_1882,In_1619,N_893);
and U1883 (N_1883,N_876,In_1120);
nor U1884 (N_1884,N_865,N_236);
or U1885 (N_1885,In_2024,N_74);
or U1886 (N_1886,In_2248,N_866);
nor U1887 (N_1887,In_237,N_513);
and U1888 (N_1888,N_622,N_636);
or U1889 (N_1889,N_833,In_812);
nor U1890 (N_1890,In_1722,N_604);
xor U1891 (N_1891,In_1412,In_1016);
and U1892 (N_1892,In_470,N_332);
or U1893 (N_1893,In_340,N_839);
nand U1894 (N_1894,In_2227,N_996);
and U1895 (N_1895,N_230,N_621);
and U1896 (N_1896,N_622,N_272);
nor U1897 (N_1897,In_2050,In_868);
nor U1898 (N_1898,N_777,N_484);
xnor U1899 (N_1899,In_1141,In_1884);
xnor U1900 (N_1900,N_663,N_625);
nor U1901 (N_1901,N_975,In_645);
xnor U1902 (N_1902,N_535,In_1961);
and U1903 (N_1903,N_0,N_561);
or U1904 (N_1904,N_174,N_957);
xor U1905 (N_1905,N_227,In_2424);
and U1906 (N_1906,In_1142,N_447);
nor U1907 (N_1907,N_982,In_1282);
or U1908 (N_1908,N_499,N_794);
nand U1909 (N_1909,In_322,N_316);
nor U1910 (N_1910,N_260,In_2101);
nand U1911 (N_1911,In_1824,N_935);
xor U1912 (N_1912,N_677,In_1238);
nand U1913 (N_1913,N_12,N_436);
and U1914 (N_1914,N_654,In_312);
nor U1915 (N_1915,N_976,N_442);
nand U1916 (N_1916,In_474,N_910);
nand U1917 (N_1917,In_1833,N_87);
xor U1918 (N_1918,In_1188,In_2043);
xor U1919 (N_1919,N_202,In_957);
nand U1920 (N_1920,N_80,N_197);
or U1921 (N_1921,N_919,N_152);
xor U1922 (N_1922,N_995,N_383);
xor U1923 (N_1923,N_43,N_483);
or U1924 (N_1924,N_315,In_717);
nand U1925 (N_1925,N_674,In_120);
nand U1926 (N_1926,N_321,N_544);
and U1927 (N_1927,In_1782,N_641);
xnor U1928 (N_1928,N_529,N_61);
xnor U1929 (N_1929,N_737,In_853);
nor U1930 (N_1930,In_2111,N_798);
or U1931 (N_1931,N_929,N_624);
nor U1932 (N_1932,N_366,N_1);
and U1933 (N_1933,N_67,In_886);
nand U1934 (N_1934,N_80,In_910);
nor U1935 (N_1935,N_470,N_329);
nand U1936 (N_1936,In_1934,N_882);
nor U1937 (N_1937,N_812,N_668);
xnor U1938 (N_1938,N_552,In_872);
or U1939 (N_1939,N_638,N_500);
nor U1940 (N_1940,N_178,N_99);
nor U1941 (N_1941,In_50,In_599);
and U1942 (N_1942,N_806,N_520);
and U1943 (N_1943,N_503,N_288);
or U1944 (N_1944,In_1670,In_972);
and U1945 (N_1945,N_487,N_475);
xor U1946 (N_1946,In_368,N_384);
or U1947 (N_1947,In_292,N_458);
and U1948 (N_1948,N_651,N_261);
nand U1949 (N_1949,N_31,In_1282);
nand U1950 (N_1950,N_58,N_389);
xnor U1951 (N_1951,N_791,N_513);
or U1952 (N_1952,N_946,In_278);
or U1953 (N_1953,N_117,In_827);
nor U1954 (N_1954,N_451,N_12);
or U1955 (N_1955,N_308,In_1002);
nand U1956 (N_1956,N_845,In_1428);
or U1957 (N_1957,In_287,In_42);
or U1958 (N_1958,N_375,N_859);
and U1959 (N_1959,In_2115,N_424);
xnor U1960 (N_1960,N_135,N_522);
nand U1961 (N_1961,N_374,N_277);
nand U1962 (N_1962,In_2437,N_992);
nor U1963 (N_1963,N_276,N_521);
nand U1964 (N_1964,N_526,N_823);
and U1965 (N_1965,N_517,N_762);
or U1966 (N_1966,In_1946,In_998);
nor U1967 (N_1967,N_708,In_1140);
nor U1968 (N_1968,In_702,N_459);
and U1969 (N_1969,In_474,In_2451);
or U1970 (N_1970,N_25,N_961);
nand U1971 (N_1971,In_400,N_344);
or U1972 (N_1972,In_1639,N_689);
xnor U1973 (N_1973,N_660,N_706);
nand U1974 (N_1974,N_721,N_211);
nand U1975 (N_1975,N_8,N_621);
nand U1976 (N_1976,In_81,N_650);
xnor U1977 (N_1977,N_883,In_2319);
xor U1978 (N_1978,N_678,N_168);
nor U1979 (N_1979,N_448,In_1910);
or U1980 (N_1980,N_48,In_1292);
and U1981 (N_1981,N_522,In_1066);
xor U1982 (N_1982,N_660,N_289);
xor U1983 (N_1983,In_1204,N_845);
nand U1984 (N_1984,N_928,In_1178);
or U1985 (N_1985,N_326,In_1153);
and U1986 (N_1986,N_990,N_528);
nand U1987 (N_1987,In_1373,In_613);
nor U1988 (N_1988,N_282,N_468);
nand U1989 (N_1989,N_243,N_183);
nor U1990 (N_1990,N_5,N_346);
or U1991 (N_1991,In_2383,N_616);
nor U1992 (N_1992,N_818,N_815);
xor U1993 (N_1993,N_322,In_1751);
xnor U1994 (N_1994,N_563,N_227);
nand U1995 (N_1995,In_470,N_704);
and U1996 (N_1996,N_756,N_723);
and U1997 (N_1997,In_2268,In_1608);
or U1998 (N_1998,N_140,In_702);
nand U1999 (N_1999,N_460,N_377);
nor U2000 (N_2000,N_1751,N_1792);
nor U2001 (N_2001,N_1173,N_1222);
xnor U2002 (N_2002,N_1512,N_1265);
and U2003 (N_2003,N_1073,N_1533);
nand U2004 (N_2004,N_1897,N_1353);
or U2005 (N_2005,N_1221,N_1345);
and U2006 (N_2006,N_1266,N_1016);
and U2007 (N_2007,N_1707,N_1996);
and U2008 (N_2008,N_1796,N_1167);
xnor U2009 (N_2009,N_1777,N_1291);
or U2010 (N_2010,N_1184,N_1986);
or U2011 (N_2011,N_1971,N_1021);
and U2012 (N_2012,N_1463,N_1113);
nand U2013 (N_2013,N_1629,N_1185);
nand U2014 (N_2014,N_1779,N_1709);
xor U2015 (N_2015,N_1359,N_1428);
nor U2016 (N_2016,N_1789,N_1880);
or U2017 (N_2017,N_1338,N_1166);
xnor U2018 (N_2018,N_1117,N_1708);
and U2019 (N_2019,N_1325,N_1989);
xnor U2020 (N_2020,N_1961,N_1775);
or U2021 (N_2021,N_1169,N_1432);
nor U2022 (N_2022,N_1627,N_1981);
nor U2023 (N_2023,N_1928,N_1774);
nor U2024 (N_2024,N_1664,N_1451);
xor U2025 (N_2025,N_1028,N_1488);
or U2026 (N_2026,N_1066,N_1308);
and U2027 (N_2027,N_1519,N_1870);
xor U2028 (N_2028,N_1554,N_1137);
nor U2029 (N_2029,N_1223,N_1980);
xnor U2030 (N_2030,N_1203,N_1361);
or U2031 (N_2031,N_1835,N_1483);
nand U2032 (N_2032,N_1450,N_1903);
nor U2033 (N_2033,N_1301,N_1472);
and U2034 (N_2034,N_1955,N_1697);
or U2035 (N_2035,N_1430,N_1857);
or U2036 (N_2036,N_1381,N_1245);
nand U2037 (N_2037,N_1691,N_1085);
nand U2038 (N_2038,N_1926,N_1787);
nor U2039 (N_2039,N_1452,N_1677);
nor U2040 (N_2040,N_1878,N_1150);
nor U2041 (N_2041,N_1761,N_1500);
xor U2042 (N_2042,N_1283,N_1997);
and U2043 (N_2043,N_1635,N_1410);
nand U2044 (N_2044,N_1847,N_1657);
xor U2045 (N_2045,N_1929,N_1667);
nand U2046 (N_2046,N_1760,N_1622);
nand U2047 (N_2047,N_1863,N_1319);
nand U2048 (N_2048,N_1302,N_1471);
xor U2049 (N_2049,N_1019,N_1322);
nor U2050 (N_2050,N_1142,N_1972);
nor U2051 (N_2051,N_1174,N_1820);
nand U2052 (N_2052,N_1672,N_1965);
or U2053 (N_2053,N_1236,N_1172);
nor U2054 (N_2054,N_1018,N_1321);
xor U2055 (N_2055,N_1821,N_1932);
nor U2056 (N_2056,N_1403,N_1521);
and U2057 (N_2057,N_1589,N_1966);
nand U2058 (N_2058,N_1230,N_1548);
nor U2059 (N_2059,N_1815,N_1336);
nor U2060 (N_2060,N_1138,N_1890);
nor U2061 (N_2061,N_1412,N_1682);
or U2062 (N_2062,N_1746,N_1941);
nor U2063 (N_2063,N_1942,N_1023);
and U2064 (N_2064,N_1656,N_1839);
xnor U2065 (N_2065,N_1573,N_1426);
or U2066 (N_2066,N_1703,N_1700);
nand U2067 (N_2067,N_1770,N_1836);
nor U2068 (N_2068,N_1045,N_1509);
or U2069 (N_2069,N_1343,N_1904);
and U2070 (N_2070,N_1603,N_1183);
or U2071 (N_2071,N_1048,N_1017);
xnor U2072 (N_2072,N_1163,N_1597);
or U2073 (N_2073,N_1885,N_1197);
nand U2074 (N_2074,N_1837,N_1952);
and U2075 (N_2075,N_1742,N_1541);
nor U2076 (N_2076,N_1539,N_1634);
or U2077 (N_2077,N_1768,N_1022);
nand U2078 (N_2078,N_1038,N_1907);
nand U2079 (N_2079,N_1094,N_1103);
or U2080 (N_2080,N_1131,N_1323);
nand U2081 (N_2081,N_1642,N_1532);
xor U2082 (N_2082,N_1062,N_1758);
or U2083 (N_2083,N_1944,N_1069);
or U2084 (N_2084,N_1369,N_1258);
xnor U2085 (N_2085,N_1335,N_1604);
nor U2086 (N_2086,N_1171,N_1090);
nor U2087 (N_2087,N_1508,N_1195);
nor U2088 (N_2088,N_1581,N_1606);
or U2089 (N_2089,N_1477,N_1724);
xnor U2090 (N_2090,N_1311,N_1752);
and U2091 (N_2091,N_1162,N_1010);
and U2092 (N_2092,N_1395,N_1374);
or U2093 (N_2093,N_1825,N_1389);
or U2094 (N_2094,N_1438,N_1262);
nor U2095 (N_2095,N_1177,N_1578);
nor U2096 (N_2096,N_1347,N_1498);
xnor U2097 (N_2097,N_1371,N_1119);
nand U2098 (N_2098,N_1782,N_1909);
or U2099 (N_2099,N_1273,N_1349);
or U2100 (N_2100,N_1009,N_1666);
nor U2101 (N_2101,N_1553,N_1831);
or U2102 (N_2102,N_1118,N_1812);
nand U2103 (N_2103,N_1688,N_1020);
nand U2104 (N_2104,N_1189,N_1620);
xor U2105 (N_2105,N_1940,N_1895);
xor U2106 (N_2106,N_1702,N_1765);
nor U2107 (N_2107,N_1797,N_1008);
and U2108 (N_2108,N_1566,N_1753);
and U2109 (N_2109,N_1954,N_1088);
nand U2110 (N_2110,N_1816,N_1969);
nand U2111 (N_2111,N_1133,N_1535);
nand U2112 (N_2112,N_1784,N_1605);
nor U2113 (N_2113,N_1851,N_1274);
nand U2114 (N_2114,N_1084,N_1098);
nor U2115 (N_2115,N_1795,N_1234);
xnor U2116 (N_2116,N_1511,N_1300);
xnor U2117 (N_2117,N_1208,N_1675);
nor U2118 (N_2118,N_1344,N_1694);
and U2119 (N_2119,N_1687,N_1292);
and U2120 (N_2120,N_1998,N_1264);
or U2121 (N_2121,N_1780,N_1003);
nor U2122 (N_2122,N_1276,N_1995);
and U2123 (N_2123,N_1176,N_1976);
xor U2124 (N_2124,N_1872,N_1446);
nand U2125 (N_2125,N_1316,N_1609);
xor U2126 (N_2126,N_1729,N_1107);
and U2127 (N_2127,N_1644,N_1306);
nand U2128 (N_2128,N_1447,N_1143);
nor U2129 (N_2129,N_1502,N_1803);
or U2130 (N_2130,N_1778,N_1884);
nor U2131 (N_2131,N_1757,N_1407);
and U2132 (N_2132,N_1528,N_1585);
nor U2133 (N_2133,N_1899,N_1728);
xnor U2134 (N_2134,N_1396,N_1948);
nor U2135 (N_2135,N_1975,N_1394);
nor U2136 (N_2136,N_1806,N_1617);
or U2137 (N_2137,N_1469,N_1994);
nand U2138 (N_2138,N_1937,N_1791);
nand U2139 (N_2139,N_1382,N_1399);
nand U2140 (N_2140,N_1494,N_1492);
nor U2141 (N_2141,N_1040,N_1035);
xor U2142 (N_2142,N_1091,N_1120);
xor U2143 (N_2143,N_1482,N_1141);
nand U2144 (N_2144,N_1653,N_1550);
and U2145 (N_2145,N_1648,N_1848);
nor U2146 (N_2146,N_1525,N_1484);
and U2147 (N_2147,N_1736,N_1582);
nand U2148 (N_2148,N_1786,N_1641);
xnor U2149 (N_2149,N_1351,N_1953);
nand U2150 (N_2150,N_1727,N_1425);
nand U2151 (N_2151,N_1423,N_1254);
nor U2152 (N_2152,N_1661,N_1717);
and U2153 (N_2153,N_1920,N_1852);
or U2154 (N_2154,N_1612,N_1523);
nand U2155 (N_2155,N_1756,N_1096);
nand U2156 (N_2156,N_1411,N_1075);
and U2157 (N_2157,N_1862,N_1845);
or U2158 (N_2158,N_1649,N_1520);
and U2159 (N_2159,N_1468,N_1654);
xnor U2160 (N_2160,N_1284,N_1346);
xnor U2161 (N_2161,N_1486,N_1571);
xor U2162 (N_2162,N_1211,N_1050);
nor U2163 (N_2163,N_1012,N_1310);
nor U2164 (N_2164,N_1507,N_1695);
nand U2165 (N_2165,N_1684,N_1487);
and U2166 (N_2166,N_1652,N_1813);
xor U2167 (N_2167,N_1330,N_1655);
nor U2168 (N_2168,N_1456,N_1187);
nand U2169 (N_2169,N_1755,N_1636);
or U2170 (N_2170,N_1122,N_1248);
nand U2171 (N_2171,N_1748,N_1945);
nand U2172 (N_2172,N_1930,N_1561);
nor U2173 (N_2173,N_1854,N_1326);
xor U2174 (N_2174,N_1624,N_1810);
nand U2175 (N_2175,N_1489,N_1046);
xor U2176 (N_2176,N_1646,N_1591);
or U2177 (N_2177,N_1136,N_1056);
and U2178 (N_2178,N_1415,N_1917);
nand U2179 (N_2179,N_1065,N_1357);
or U2180 (N_2180,N_1332,N_1607);
nand U2181 (N_2181,N_1424,N_1720);
nand U2182 (N_2182,N_1828,N_1239);
nand U2183 (N_2183,N_1387,N_1296);
nand U2184 (N_2184,N_1275,N_1315);
xnor U2185 (N_2185,N_1252,N_1112);
nand U2186 (N_2186,N_1470,N_1567);
xor U2187 (N_2187,N_1776,N_1946);
nand U2188 (N_2188,N_1280,N_1632);
nand U2189 (N_2189,N_1421,N_1958);
xor U2190 (N_2190,N_1750,N_1026);
and U2191 (N_2191,N_1517,N_1647);
or U2192 (N_2192,N_1706,N_1988);
nor U2193 (N_2193,N_1053,N_1157);
nand U2194 (N_2194,N_1401,N_1538);
or U2195 (N_2195,N_1933,N_1598);
or U2196 (N_2196,N_1095,N_1373);
or U2197 (N_2197,N_1216,N_1071);
nand U2198 (N_2198,N_1840,N_1715);
nand U2199 (N_2199,N_1288,N_1874);
or U2200 (N_2200,N_1237,N_1043);
nor U2201 (N_2201,N_1414,N_1584);
xnor U2202 (N_2202,N_1984,N_1429);
nand U2203 (N_2203,N_1910,N_1537);
or U2204 (N_2204,N_1923,N_1179);
nand U2205 (N_2205,N_1089,N_1466);
nor U2206 (N_2206,N_1377,N_1145);
nor U2207 (N_2207,N_1514,N_1147);
and U2208 (N_2208,N_1983,N_1207);
and U2209 (N_2209,N_1467,N_1362);
nor U2210 (N_2210,N_1490,N_1723);
and U2211 (N_2211,N_1229,N_1444);
nor U2212 (N_2212,N_1549,N_1305);
nand U2213 (N_2213,N_1979,N_1586);
or U2214 (N_2214,N_1670,N_1331);
nand U2215 (N_2215,N_1406,N_1194);
or U2216 (N_2216,N_1455,N_1398);
nand U2217 (N_2217,N_1294,N_1327);
or U2218 (N_2218,N_1564,N_1059);
and U2219 (N_2219,N_1767,N_1485);
and U2220 (N_2220,N_1210,N_1834);
xor U2221 (N_2221,N_1154,N_1613);
xor U2222 (N_2222,N_1730,N_1417);
or U2223 (N_2223,N_1151,N_1633);
nor U2224 (N_2224,N_1693,N_1741);
nand U2225 (N_2225,N_1201,N_1731);
and U2226 (N_2226,N_1393,N_1220);
or U2227 (N_2227,N_1449,N_1832);
xor U2228 (N_2228,N_1156,N_1200);
nand U2229 (N_2229,N_1384,N_1978);
xnor U2230 (N_2230,N_1843,N_1547);
and U2231 (N_2231,N_1552,N_1555);
or U2232 (N_2232,N_1722,N_1130);
and U2233 (N_2233,N_1129,N_1376);
or U2234 (N_2234,N_1039,N_1850);
and U2235 (N_2235,N_1918,N_1745);
nand U2236 (N_2236,N_1320,N_1557);
nand U2237 (N_2237,N_1186,N_1427);
xor U2238 (N_2238,N_1146,N_1947);
nand U2239 (N_2239,N_1800,N_1809);
xor U2240 (N_2240,N_1999,N_1608);
nor U2241 (N_2241,N_1256,N_1811);
nor U2242 (N_2242,N_1808,N_1788);
nand U2243 (N_2243,N_1052,N_1665);
and U2244 (N_2244,N_1830,N_1799);
or U2245 (N_2245,N_1710,N_1372);
nor U2246 (N_2246,N_1974,N_1576);
and U2247 (N_2247,N_1977,N_1842);
xor U2248 (N_2248,N_1737,N_1562);
or U2249 (N_2249,N_1199,N_1299);
nand U2250 (N_2250,N_1272,N_1864);
nor U2251 (N_2251,N_1902,N_1716);
or U2252 (N_2252,N_1559,N_1970);
nor U2253 (N_2253,N_1445,N_1202);
nor U2254 (N_2254,N_1919,N_1893);
nor U2255 (N_2255,N_1312,N_1712);
nor U2256 (N_2256,N_1668,N_1527);
nand U2257 (N_2257,N_1060,N_1504);
nand U2258 (N_2258,N_1224,N_1270);
or U2259 (N_2259,N_1630,N_1366);
or U2260 (N_2260,N_1253,N_1459);
xor U2261 (N_2261,N_1798,N_1277);
or U2262 (N_2262,N_1123,N_1911);
or U2263 (N_2263,N_1287,N_1804);
nor U2264 (N_2264,N_1900,N_1858);
nor U2265 (N_2265,N_1105,N_1704);
or U2266 (N_2266,N_1198,N_1121);
nand U2267 (N_2267,N_1987,N_1883);
and U2268 (N_2268,N_1114,N_1214);
nand U2269 (N_2269,N_1570,N_1462);
and U2270 (N_2270,N_1152,N_1031);
nor U2271 (N_2271,N_1409,N_1061);
xnor U2272 (N_2272,N_1626,N_1558);
or U2273 (N_2273,N_1030,N_1099);
xor U2274 (N_2274,N_1908,N_1378);
xor U2275 (N_2275,N_1293,N_1602);
or U2276 (N_2276,N_1610,N_1307);
or U2277 (N_2277,N_1771,N_1478);
xnor U2278 (N_2278,N_1713,N_1676);
and U2279 (N_2279,N_1473,N_1298);
and U2280 (N_2280,N_1826,N_1140);
xnor U2281 (N_2281,N_1587,N_1260);
xor U2282 (N_2282,N_1279,N_1155);
or U2283 (N_2283,N_1457,N_1696);
xnor U2284 (N_2284,N_1259,N_1574);
xor U2285 (N_2285,N_1464,N_1901);
nand U2286 (N_2286,N_1711,N_1355);
nand U2287 (N_2287,N_1419,N_1583);
xor U2288 (N_2288,N_1364,N_1191);
nand U2289 (N_2289,N_1556,N_1628);
and U2290 (N_2290,N_1093,N_1081);
or U2291 (N_2291,N_1663,N_1499);
or U2292 (N_2292,N_1599,N_1615);
or U2293 (N_2293,N_1125,N_1437);
or U2294 (N_2294,N_1973,N_1493);
xor U2295 (N_2295,N_1960,N_1681);
nand U2296 (N_2296,N_1754,N_1116);
and U2297 (N_2297,N_1241,N_1460);
nand U2298 (N_2298,N_1744,N_1442);
nor U2299 (N_2299,N_1070,N_1660);
nand U2300 (N_2300,N_1268,N_1416);
nand U2301 (N_2301,N_1213,N_1188);
or U2302 (N_2302,N_1049,N_1160);
or U2303 (N_2303,N_1422,N_1859);
and U2304 (N_2304,N_1856,N_1443);
or U2305 (N_2305,N_1178,N_1985);
and U2306 (N_2306,N_1014,N_1651);
and U2307 (N_2307,N_1855,N_1013);
nor U2308 (N_2308,N_1501,N_1454);
xor U2309 (N_2309,N_1064,N_1108);
nand U2310 (N_2310,N_1165,N_1569);
xor U2311 (N_2311,N_1993,N_1029);
nor U2312 (N_2312,N_1801,N_1645);
nand U2313 (N_2313,N_1982,N_1936);
xor U2314 (N_2314,N_1882,N_1408);
and U2315 (N_2315,N_1110,N_1916);
nand U2316 (N_2316,N_1225,N_1530);
or U2317 (N_2317,N_1853,N_1869);
and U2318 (N_2318,N_1625,N_1565);
nand U2319 (N_2319,N_1402,N_1139);
or U2320 (N_2320,N_1363,N_1314);
or U2321 (N_2321,N_1204,N_1790);
nor U2322 (N_2322,N_1898,N_1631);
nor U2323 (N_2323,N_1431,N_1887);
xor U2324 (N_2324,N_1518,N_1540);
nand U2325 (N_2325,N_1531,N_1873);
nand U2326 (N_2326,N_1912,N_1124);
xor U2327 (N_2327,N_1235,N_1699);
or U2328 (N_2328,N_1005,N_1563);
and U2329 (N_2329,N_1934,N_1285);
xor U2330 (N_2330,N_1297,N_1689);
and U2331 (N_2331,N_1168,N_1618);
or U2332 (N_2332,N_1823,N_1218);
or U2333 (N_2333,N_1659,N_1818);
or U2334 (N_2334,N_1196,N_1243);
nand U2335 (N_2335,N_1180,N_1405);
nor U2336 (N_2336,N_1611,N_1833);
nand U2337 (N_2337,N_1082,N_1546);
nand U2338 (N_2338,N_1764,N_1006);
and U2339 (N_2339,N_1956,N_1888);
xor U2340 (N_2340,N_1434,N_1205);
nor U2341 (N_2341,N_1106,N_1719);
nor U2342 (N_2342,N_1568,N_1244);
or U2343 (N_2343,N_1192,N_1058);
nand U2344 (N_2344,N_1705,N_1718);
or U2345 (N_2345,N_1922,N_1925);
and U2346 (N_2346,N_1905,N_1865);
or U2347 (N_2347,N_1435,N_1304);
nor U2348 (N_2348,N_1824,N_1232);
or U2349 (N_2349,N_1251,N_1068);
nor U2350 (N_2350,N_1324,N_1233);
nand U2351 (N_2351,N_1889,N_1219);
and U2352 (N_2352,N_1250,N_1759);
xnor U2353 (N_2353,N_1404,N_1924);
xnor U2354 (N_2354,N_1128,N_1935);
xnor U2355 (N_2355,N_1242,N_1092);
xor U2356 (N_2356,N_1126,N_1102);
nand U2357 (N_2357,N_1158,N_1441);
or U2358 (N_2358,N_1481,N_1807);
xnor U2359 (N_2359,N_1590,N_1572);
and U2360 (N_2360,N_1866,N_1181);
nor U2361 (N_2361,N_1747,N_1101);
and U2362 (N_2362,N_1593,N_1333);
nand U2363 (N_2363,N_1032,N_1391);
nand U2364 (N_2364,N_1001,N_1650);
nand U2365 (N_2365,N_1033,N_1621);
and U2366 (N_2366,N_1024,N_1475);
nor U2367 (N_2367,N_1733,N_1877);
and U2368 (N_2368,N_1692,N_1785);
and U2369 (N_2369,N_1240,N_1354);
and U2370 (N_2370,N_1115,N_1577);
or U2371 (N_2371,N_1734,N_1849);
or U2372 (N_2372,N_1543,N_1871);
or U2373 (N_2373,N_1397,N_1080);
xor U2374 (N_2374,N_1257,N_1943);
xnor U2375 (N_2375,N_1261,N_1164);
nor U2376 (N_2376,N_1515,N_1673);
xor U2377 (N_2377,N_1783,N_1968);
nand U2378 (N_2378,N_1057,N_1674);
or U2379 (N_2379,N_1614,N_1992);
nor U2380 (N_2380,N_1418,N_1350);
nor U2381 (N_2381,N_1051,N_1465);
nand U2382 (N_2382,N_1356,N_1328);
xor U2383 (N_2383,N_1303,N_1149);
nor U2384 (N_2384,N_1671,N_1891);
nand U2385 (N_2385,N_1819,N_1588);
nor U2386 (N_2386,N_1762,N_1639);
or U2387 (N_2387,N_1111,N_1949);
nand U2388 (N_2388,N_1063,N_1440);
nor U2389 (N_2389,N_1109,N_1036);
nand U2390 (N_2390,N_1217,N_1286);
nand U2391 (N_2391,N_1662,N_1370);
nand U2392 (N_2392,N_1025,N_1913);
xor U2393 (N_2393,N_1579,N_1915);
nand U2394 (N_2394,N_1011,N_1383);
and U2395 (N_2395,N_1506,N_1860);
and U2396 (N_2396,N_1749,N_1476);
and U2397 (N_2397,N_1153,N_1295);
or U2398 (N_2398,N_1726,N_1193);
nand U2399 (N_2399,N_1772,N_1209);
or U2400 (N_2400,N_1439,N_1781);
and U2401 (N_2401,N_1074,N_1990);
xnor U2402 (N_2402,N_1215,N_1551);
nand U2403 (N_2403,N_1067,N_1829);
or U2404 (N_2404,N_1247,N_1773);
and U2405 (N_2405,N_1365,N_1002);
and U2406 (N_2406,N_1991,N_1339);
xor U2407 (N_2407,N_1950,N_1802);
or U2408 (N_2408,N_1433,N_1846);
and U2409 (N_2409,N_1963,N_1448);
or U2410 (N_2410,N_1458,N_1015);
or U2411 (N_2411,N_1267,N_1278);
nand U2412 (N_2412,N_1637,N_1461);
nor U2413 (N_2413,N_1479,N_1600);
and U2414 (N_2414,N_1097,N_1685);
and U2415 (N_2415,N_1896,N_1875);
and U2416 (N_2416,N_1714,N_1739);
and U2417 (N_2417,N_1669,N_1868);
nand U2418 (N_2418,N_1255,N_1725);
nand U2419 (N_2419,N_1643,N_1545);
and U2420 (N_2420,N_1436,N_1938);
and U2421 (N_2421,N_1161,N_1000);
xor U2422 (N_2422,N_1601,N_1794);
nand U2423 (N_2423,N_1309,N_1341);
nand U2424 (N_2424,N_1827,N_1480);
nor U2425 (N_2425,N_1496,N_1360);
and U2426 (N_2426,N_1249,N_1078);
or U2427 (N_2427,N_1886,N_1542);
or U2428 (N_2428,N_1281,N_1732);
xor U2429 (N_2429,N_1861,N_1054);
and U2430 (N_2430,N_1740,N_1595);
nand U2431 (N_2431,N_1334,N_1317);
nand U2432 (N_2432,N_1290,N_1379);
xor U2433 (N_2433,N_1453,N_1190);
and U2434 (N_2434,N_1269,N_1516);
xor U2435 (N_2435,N_1623,N_1505);
xor U2436 (N_2436,N_1495,N_1701);
nand U2437 (N_2437,N_1616,N_1939);
nand U2438 (N_2438,N_1282,N_1735);
and U2439 (N_2439,N_1678,N_1104);
nand U2440 (N_2440,N_1544,N_1522);
or U2441 (N_2441,N_1738,N_1263);
and U2442 (N_2442,N_1144,N_1763);
xnor U2443 (N_2443,N_1079,N_1148);
nor U2444 (N_2444,N_1077,N_1159);
and U2445 (N_2445,N_1367,N_1822);
nor U2446 (N_2446,N_1175,N_1640);
nand U2447 (N_2447,N_1037,N_1951);
and U2448 (N_2448,N_1076,N_1580);
nor U2449 (N_2449,N_1385,N_1841);
xnor U2450 (N_2450,N_1047,N_1340);
nor U2451 (N_2451,N_1683,N_1231);
nor U2452 (N_2452,N_1817,N_1375);
xnor U2453 (N_2453,N_1690,N_1289);
nand U2454 (N_2454,N_1358,N_1793);
or U2455 (N_2455,N_1814,N_1238);
xnor U2456 (N_2456,N_1135,N_1127);
nand U2457 (N_2457,N_1007,N_1894);
or U2458 (N_2458,N_1004,N_1368);
nand U2459 (N_2459,N_1348,N_1967);
or U2460 (N_2460,N_1041,N_1083);
or U2461 (N_2461,N_1380,N_1638);
nor U2462 (N_2462,N_1914,N_1413);
nor U2463 (N_2463,N_1892,N_1686);
nand U2464 (N_2464,N_1619,N_1931);
and U2465 (N_2465,N_1536,N_1927);
nand U2466 (N_2466,N_1027,N_1921);
xor U2467 (N_2467,N_1227,N_1679);
or U2468 (N_2468,N_1534,N_1743);
nor U2469 (N_2469,N_1698,N_1087);
nand U2470 (N_2470,N_1529,N_1964);
or U2471 (N_2471,N_1560,N_1876);
nor U2472 (N_2472,N_1805,N_1503);
and U2473 (N_2473,N_1170,N_1838);
or U2474 (N_2474,N_1766,N_1132);
nand U2475 (N_2475,N_1034,N_1271);
xor U2476 (N_2476,N_1228,N_1881);
nand U2477 (N_2477,N_1400,N_1246);
or U2478 (N_2478,N_1182,N_1134);
and U2479 (N_2479,N_1721,N_1044);
nor U2480 (N_2480,N_1526,N_1212);
nand U2481 (N_2481,N_1962,N_1072);
nand U2482 (N_2482,N_1352,N_1906);
or U2483 (N_2483,N_1491,N_1769);
nor U2484 (N_2484,N_1313,N_1844);
and U2485 (N_2485,N_1879,N_1392);
xnor U2486 (N_2486,N_1592,N_1510);
nand U2487 (N_2487,N_1100,N_1206);
nor U2488 (N_2488,N_1329,N_1594);
and U2489 (N_2489,N_1680,N_1042);
xnor U2490 (N_2490,N_1658,N_1342);
and U2491 (N_2491,N_1957,N_1388);
nand U2492 (N_2492,N_1337,N_1474);
nor U2493 (N_2493,N_1867,N_1390);
nor U2494 (N_2494,N_1497,N_1596);
and U2495 (N_2495,N_1959,N_1420);
nor U2496 (N_2496,N_1318,N_1575);
and U2497 (N_2497,N_1226,N_1086);
nor U2498 (N_2498,N_1055,N_1513);
xor U2499 (N_2499,N_1386,N_1524);
or U2500 (N_2500,N_1274,N_1742);
xnor U2501 (N_2501,N_1788,N_1146);
xor U2502 (N_2502,N_1883,N_1518);
nand U2503 (N_2503,N_1798,N_1841);
xnor U2504 (N_2504,N_1524,N_1265);
xnor U2505 (N_2505,N_1211,N_1527);
nor U2506 (N_2506,N_1207,N_1852);
or U2507 (N_2507,N_1799,N_1211);
and U2508 (N_2508,N_1063,N_1023);
xnor U2509 (N_2509,N_1040,N_1558);
nand U2510 (N_2510,N_1725,N_1371);
nand U2511 (N_2511,N_1239,N_1684);
nand U2512 (N_2512,N_1573,N_1325);
nand U2513 (N_2513,N_1076,N_1706);
nor U2514 (N_2514,N_1785,N_1870);
and U2515 (N_2515,N_1596,N_1269);
and U2516 (N_2516,N_1594,N_1448);
nand U2517 (N_2517,N_1278,N_1245);
xnor U2518 (N_2518,N_1232,N_1999);
nor U2519 (N_2519,N_1034,N_1333);
xor U2520 (N_2520,N_1688,N_1278);
nand U2521 (N_2521,N_1407,N_1608);
nand U2522 (N_2522,N_1521,N_1606);
nor U2523 (N_2523,N_1221,N_1522);
nand U2524 (N_2524,N_1167,N_1605);
nand U2525 (N_2525,N_1954,N_1556);
and U2526 (N_2526,N_1115,N_1280);
nand U2527 (N_2527,N_1802,N_1179);
or U2528 (N_2528,N_1836,N_1511);
xor U2529 (N_2529,N_1811,N_1662);
xor U2530 (N_2530,N_1274,N_1582);
and U2531 (N_2531,N_1674,N_1374);
nor U2532 (N_2532,N_1866,N_1807);
and U2533 (N_2533,N_1364,N_1394);
nor U2534 (N_2534,N_1914,N_1796);
and U2535 (N_2535,N_1799,N_1420);
nor U2536 (N_2536,N_1802,N_1986);
or U2537 (N_2537,N_1762,N_1356);
nor U2538 (N_2538,N_1791,N_1680);
nor U2539 (N_2539,N_1114,N_1799);
xor U2540 (N_2540,N_1632,N_1410);
xor U2541 (N_2541,N_1083,N_1489);
nor U2542 (N_2542,N_1559,N_1869);
nor U2543 (N_2543,N_1807,N_1082);
nor U2544 (N_2544,N_1214,N_1750);
or U2545 (N_2545,N_1098,N_1460);
nand U2546 (N_2546,N_1827,N_1553);
xnor U2547 (N_2547,N_1608,N_1652);
or U2548 (N_2548,N_1922,N_1695);
nand U2549 (N_2549,N_1135,N_1701);
or U2550 (N_2550,N_1893,N_1084);
and U2551 (N_2551,N_1809,N_1504);
xnor U2552 (N_2552,N_1858,N_1757);
xnor U2553 (N_2553,N_1890,N_1772);
xnor U2554 (N_2554,N_1884,N_1496);
nor U2555 (N_2555,N_1658,N_1244);
and U2556 (N_2556,N_1795,N_1350);
or U2557 (N_2557,N_1186,N_1982);
xnor U2558 (N_2558,N_1870,N_1321);
nor U2559 (N_2559,N_1035,N_1297);
and U2560 (N_2560,N_1829,N_1293);
and U2561 (N_2561,N_1571,N_1529);
or U2562 (N_2562,N_1981,N_1397);
nand U2563 (N_2563,N_1591,N_1513);
nor U2564 (N_2564,N_1858,N_1206);
nor U2565 (N_2565,N_1572,N_1283);
nor U2566 (N_2566,N_1233,N_1890);
nor U2567 (N_2567,N_1498,N_1322);
or U2568 (N_2568,N_1008,N_1633);
or U2569 (N_2569,N_1856,N_1265);
and U2570 (N_2570,N_1316,N_1431);
nor U2571 (N_2571,N_1006,N_1685);
and U2572 (N_2572,N_1725,N_1080);
nand U2573 (N_2573,N_1313,N_1416);
or U2574 (N_2574,N_1956,N_1488);
and U2575 (N_2575,N_1746,N_1211);
or U2576 (N_2576,N_1476,N_1260);
xor U2577 (N_2577,N_1288,N_1320);
nand U2578 (N_2578,N_1565,N_1618);
and U2579 (N_2579,N_1377,N_1498);
nor U2580 (N_2580,N_1719,N_1556);
nand U2581 (N_2581,N_1343,N_1760);
and U2582 (N_2582,N_1141,N_1496);
xor U2583 (N_2583,N_1884,N_1053);
nand U2584 (N_2584,N_1190,N_1469);
xnor U2585 (N_2585,N_1102,N_1115);
nand U2586 (N_2586,N_1275,N_1051);
and U2587 (N_2587,N_1685,N_1606);
xnor U2588 (N_2588,N_1925,N_1250);
and U2589 (N_2589,N_1778,N_1542);
nor U2590 (N_2590,N_1066,N_1499);
nand U2591 (N_2591,N_1979,N_1165);
nor U2592 (N_2592,N_1502,N_1883);
xor U2593 (N_2593,N_1856,N_1864);
or U2594 (N_2594,N_1917,N_1867);
or U2595 (N_2595,N_1344,N_1134);
nand U2596 (N_2596,N_1795,N_1308);
xnor U2597 (N_2597,N_1976,N_1335);
nand U2598 (N_2598,N_1792,N_1198);
xnor U2599 (N_2599,N_1630,N_1347);
or U2600 (N_2600,N_1016,N_1353);
or U2601 (N_2601,N_1721,N_1851);
and U2602 (N_2602,N_1833,N_1943);
or U2603 (N_2603,N_1912,N_1919);
xor U2604 (N_2604,N_1323,N_1108);
and U2605 (N_2605,N_1245,N_1959);
nand U2606 (N_2606,N_1244,N_1990);
xnor U2607 (N_2607,N_1652,N_1950);
nand U2608 (N_2608,N_1218,N_1454);
nand U2609 (N_2609,N_1444,N_1271);
or U2610 (N_2610,N_1950,N_1795);
nor U2611 (N_2611,N_1574,N_1606);
or U2612 (N_2612,N_1793,N_1907);
nor U2613 (N_2613,N_1083,N_1001);
or U2614 (N_2614,N_1459,N_1645);
nor U2615 (N_2615,N_1883,N_1723);
and U2616 (N_2616,N_1565,N_1059);
and U2617 (N_2617,N_1702,N_1927);
and U2618 (N_2618,N_1681,N_1782);
and U2619 (N_2619,N_1245,N_1939);
xor U2620 (N_2620,N_1414,N_1530);
nor U2621 (N_2621,N_1743,N_1829);
nand U2622 (N_2622,N_1739,N_1801);
or U2623 (N_2623,N_1611,N_1012);
and U2624 (N_2624,N_1363,N_1649);
and U2625 (N_2625,N_1129,N_1573);
nand U2626 (N_2626,N_1772,N_1451);
and U2627 (N_2627,N_1747,N_1335);
xnor U2628 (N_2628,N_1516,N_1696);
nand U2629 (N_2629,N_1422,N_1297);
and U2630 (N_2630,N_1730,N_1186);
or U2631 (N_2631,N_1263,N_1488);
or U2632 (N_2632,N_1375,N_1299);
nor U2633 (N_2633,N_1034,N_1010);
or U2634 (N_2634,N_1972,N_1080);
xor U2635 (N_2635,N_1875,N_1563);
or U2636 (N_2636,N_1092,N_1195);
nand U2637 (N_2637,N_1035,N_1782);
nor U2638 (N_2638,N_1749,N_1059);
nor U2639 (N_2639,N_1494,N_1411);
nor U2640 (N_2640,N_1945,N_1900);
xnor U2641 (N_2641,N_1345,N_1227);
nand U2642 (N_2642,N_1139,N_1526);
xor U2643 (N_2643,N_1971,N_1423);
or U2644 (N_2644,N_1261,N_1319);
nor U2645 (N_2645,N_1500,N_1180);
or U2646 (N_2646,N_1548,N_1132);
nor U2647 (N_2647,N_1488,N_1431);
nor U2648 (N_2648,N_1545,N_1100);
or U2649 (N_2649,N_1783,N_1592);
nor U2650 (N_2650,N_1827,N_1375);
nor U2651 (N_2651,N_1866,N_1736);
or U2652 (N_2652,N_1170,N_1322);
xnor U2653 (N_2653,N_1847,N_1004);
or U2654 (N_2654,N_1477,N_1009);
xnor U2655 (N_2655,N_1452,N_1783);
xor U2656 (N_2656,N_1671,N_1343);
or U2657 (N_2657,N_1215,N_1091);
nand U2658 (N_2658,N_1475,N_1984);
or U2659 (N_2659,N_1143,N_1401);
or U2660 (N_2660,N_1177,N_1203);
or U2661 (N_2661,N_1886,N_1984);
and U2662 (N_2662,N_1693,N_1091);
or U2663 (N_2663,N_1835,N_1228);
xor U2664 (N_2664,N_1144,N_1336);
nand U2665 (N_2665,N_1559,N_1491);
or U2666 (N_2666,N_1011,N_1935);
or U2667 (N_2667,N_1834,N_1882);
nor U2668 (N_2668,N_1471,N_1831);
nor U2669 (N_2669,N_1401,N_1877);
nor U2670 (N_2670,N_1958,N_1866);
nand U2671 (N_2671,N_1130,N_1557);
and U2672 (N_2672,N_1310,N_1991);
or U2673 (N_2673,N_1289,N_1712);
nand U2674 (N_2674,N_1046,N_1457);
xnor U2675 (N_2675,N_1251,N_1633);
xor U2676 (N_2676,N_1707,N_1607);
nand U2677 (N_2677,N_1753,N_1708);
nor U2678 (N_2678,N_1602,N_1491);
nor U2679 (N_2679,N_1235,N_1132);
and U2680 (N_2680,N_1352,N_1182);
or U2681 (N_2681,N_1839,N_1579);
or U2682 (N_2682,N_1187,N_1607);
nor U2683 (N_2683,N_1761,N_1860);
and U2684 (N_2684,N_1760,N_1810);
xnor U2685 (N_2685,N_1076,N_1826);
and U2686 (N_2686,N_1512,N_1732);
nand U2687 (N_2687,N_1272,N_1896);
nand U2688 (N_2688,N_1410,N_1840);
nand U2689 (N_2689,N_1554,N_1363);
xnor U2690 (N_2690,N_1310,N_1177);
xnor U2691 (N_2691,N_1229,N_1302);
nor U2692 (N_2692,N_1896,N_1596);
and U2693 (N_2693,N_1503,N_1717);
xor U2694 (N_2694,N_1601,N_1579);
or U2695 (N_2695,N_1678,N_1203);
and U2696 (N_2696,N_1818,N_1316);
and U2697 (N_2697,N_1605,N_1259);
nand U2698 (N_2698,N_1574,N_1298);
xor U2699 (N_2699,N_1543,N_1619);
and U2700 (N_2700,N_1123,N_1925);
nand U2701 (N_2701,N_1809,N_1064);
nand U2702 (N_2702,N_1805,N_1217);
nand U2703 (N_2703,N_1226,N_1584);
xnor U2704 (N_2704,N_1677,N_1393);
nor U2705 (N_2705,N_1545,N_1638);
nand U2706 (N_2706,N_1322,N_1774);
and U2707 (N_2707,N_1587,N_1479);
and U2708 (N_2708,N_1980,N_1043);
nand U2709 (N_2709,N_1556,N_1623);
or U2710 (N_2710,N_1330,N_1906);
nor U2711 (N_2711,N_1885,N_1698);
or U2712 (N_2712,N_1590,N_1638);
nor U2713 (N_2713,N_1744,N_1474);
nor U2714 (N_2714,N_1315,N_1355);
and U2715 (N_2715,N_1630,N_1442);
xor U2716 (N_2716,N_1176,N_1140);
or U2717 (N_2717,N_1642,N_1892);
or U2718 (N_2718,N_1480,N_1996);
and U2719 (N_2719,N_1005,N_1169);
or U2720 (N_2720,N_1877,N_1659);
and U2721 (N_2721,N_1695,N_1049);
xnor U2722 (N_2722,N_1873,N_1470);
or U2723 (N_2723,N_1784,N_1254);
and U2724 (N_2724,N_1671,N_1449);
xnor U2725 (N_2725,N_1221,N_1514);
or U2726 (N_2726,N_1935,N_1066);
nand U2727 (N_2727,N_1831,N_1502);
and U2728 (N_2728,N_1161,N_1891);
xor U2729 (N_2729,N_1139,N_1129);
nand U2730 (N_2730,N_1699,N_1384);
or U2731 (N_2731,N_1031,N_1564);
nor U2732 (N_2732,N_1474,N_1662);
nand U2733 (N_2733,N_1310,N_1740);
nand U2734 (N_2734,N_1806,N_1308);
nand U2735 (N_2735,N_1352,N_1677);
xor U2736 (N_2736,N_1323,N_1687);
or U2737 (N_2737,N_1082,N_1898);
and U2738 (N_2738,N_1535,N_1387);
and U2739 (N_2739,N_1810,N_1520);
xor U2740 (N_2740,N_1426,N_1654);
or U2741 (N_2741,N_1527,N_1333);
and U2742 (N_2742,N_1128,N_1247);
nand U2743 (N_2743,N_1830,N_1563);
or U2744 (N_2744,N_1258,N_1811);
nor U2745 (N_2745,N_1377,N_1171);
and U2746 (N_2746,N_1258,N_1558);
xor U2747 (N_2747,N_1316,N_1653);
nor U2748 (N_2748,N_1840,N_1719);
or U2749 (N_2749,N_1775,N_1216);
and U2750 (N_2750,N_1180,N_1621);
and U2751 (N_2751,N_1903,N_1275);
nor U2752 (N_2752,N_1787,N_1863);
nand U2753 (N_2753,N_1790,N_1967);
xnor U2754 (N_2754,N_1869,N_1702);
nor U2755 (N_2755,N_1440,N_1569);
xor U2756 (N_2756,N_1188,N_1864);
and U2757 (N_2757,N_1497,N_1817);
and U2758 (N_2758,N_1339,N_1978);
nand U2759 (N_2759,N_1509,N_1696);
nand U2760 (N_2760,N_1575,N_1573);
and U2761 (N_2761,N_1805,N_1414);
and U2762 (N_2762,N_1546,N_1090);
xnor U2763 (N_2763,N_1728,N_1715);
nor U2764 (N_2764,N_1669,N_1217);
xnor U2765 (N_2765,N_1159,N_1029);
or U2766 (N_2766,N_1733,N_1466);
nand U2767 (N_2767,N_1259,N_1374);
xnor U2768 (N_2768,N_1226,N_1625);
and U2769 (N_2769,N_1973,N_1007);
and U2770 (N_2770,N_1942,N_1893);
and U2771 (N_2771,N_1046,N_1226);
xor U2772 (N_2772,N_1365,N_1452);
nor U2773 (N_2773,N_1001,N_1438);
xor U2774 (N_2774,N_1534,N_1720);
nor U2775 (N_2775,N_1687,N_1243);
and U2776 (N_2776,N_1625,N_1129);
nand U2777 (N_2777,N_1560,N_1545);
and U2778 (N_2778,N_1870,N_1875);
and U2779 (N_2779,N_1781,N_1729);
nand U2780 (N_2780,N_1717,N_1066);
nor U2781 (N_2781,N_1156,N_1538);
and U2782 (N_2782,N_1391,N_1116);
or U2783 (N_2783,N_1242,N_1411);
xnor U2784 (N_2784,N_1413,N_1767);
and U2785 (N_2785,N_1415,N_1977);
nand U2786 (N_2786,N_1868,N_1029);
and U2787 (N_2787,N_1806,N_1932);
or U2788 (N_2788,N_1127,N_1669);
nand U2789 (N_2789,N_1154,N_1874);
nand U2790 (N_2790,N_1600,N_1468);
nor U2791 (N_2791,N_1430,N_1196);
or U2792 (N_2792,N_1831,N_1346);
nor U2793 (N_2793,N_1556,N_1098);
nor U2794 (N_2794,N_1082,N_1170);
and U2795 (N_2795,N_1742,N_1316);
and U2796 (N_2796,N_1933,N_1416);
and U2797 (N_2797,N_1023,N_1171);
nand U2798 (N_2798,N_1207,N_1307);
xnor U2799 (N_2799,N_1420,N_1070);
nor U2800 (N_2800,N_1092,N_1869);
or U2801 (N_2801,N_1032,N_1553);
nand U2802 (N_2802,N_1847,N_1660);
nor U2803 (N_2803,N_1324,N_1849);
nand U2804 (N_2804,N_1406,N_1690);
and U2805 (N_2805,N_1199,N_1584);
nand U2806 (N_2806,N_1421,N_1531);
nor U2807 (N_2807,N_1020,N_1327);
or U2808 (N_2808,N_1184,N_1625);
nor U2809 (N_2809,N_1578,N_1598);
xor U2810 (N_2810,N_1189,N_1719);
and U2811 (N_2811,N_1020,N_1083);
nor U2812 (N_2812,N_1297,N_1303);
nor U2813 (N_2813,N_1036,N_1928);
nand U2814 (N_2814,N_1011,N_1449);
or U2815 (N_2815,N_1498,N_1878);
nand U2816 (N_2816,N_1908,N_1438);
xor U2817 (N_2817,N_1080,N_1991);
nor U2818 (N_2818,N_1728,N_1414);
and U2819 (N_2819,N_1918,N_1975);
or U2820 (N_2820,N_1132,N_1901);
nor U2821 (N_2821,N_1765,N_1873);
nor U2822 (N_2822,N_1304,N_1798);
nand U2823 (N_2823,N_1885,N_1171);
and U2824 (N_2824,N_1876,N_1648);
xor U2825 (N_2825,N_1155,N_1163);
nand U2826 (N_2826,N_1357,N_1353);
or U2827 (N_2827,N_1436,N_1129);
xor U2828 (N_2828,N_1064,N_1953);
and U2829 (N_2829,N_1812,N_1570);
nand U2830 (N_2830,N_1042,N_1155);
xor U2831 (N_2831,N_1306,N_1682);
and U2832 (N_2832,N_1964,N_1899);
nor U2833 (N_2833,N_1068,N_1107);
nand U2834 (N_2834,N_1962,N_1280);
or U2835 (N_2835,N_1913,N_1146);
xor U2836 (N_2836,N_1718,N_1083);
and U2837 (N_2837,N_1298,N_1139);
nand U2838 (N_2838,N_1824,N_1208);
nor U2839 (N_2839,N_1472,N_1758);
and U2840 (N_2840,N_1765,N_1704);
xnor U2841 (N_2841,N_1282,N_1276);
or U2842 (N_2842,N_1067,N_1942);
xnor U2843 (N_2843,N_1345,N_1139);
nor U2844 (N_2844,N_1056,N_1157);
nor U2845 (N_2845,N_1290,N_1749);
and U2846 (N_2846,N_1716,N_1270);
or U2847 (N_2847,N_1611,N_1951);
and U2848 (N_2848,N_1111,N_1940);
nor U2849 (N_2849,N_1771,N_1952);
and U2850 (N_2850,N_1086,N_1344);
nand U2851 (N_2851,N_1658,N_1914);
nand U2852 (N_2852,N_1939,N_1532);
nand U2853 (N_2853,N_1411,N_1515);
and U2854 (N_2854,N_1947,N_1244);
and U2855 (N_2855,N_1553,N_1093);
nand U2856 (N_2856,N_1981,N_1307);
xnor U2857 (N_2857,N_1352,N_1854);
nor U2858 (N_2858,N_1699,N_1224);
xnor U2859 (N_2859,N_1647,N_1937);
or U2860 (N_2860,N_1653,N_1807);
or U2861 (N_2861,N_1014,N_1116);
xnor U2862 (N_2862,N_1240,N_1567);
or U2863 (N_2863,N_1492,N_1654);
and U2864 (N_2864,N_1664,N_1093);
and U2865 (N_2865,N_1430,N_1152);
nand U2866 (N_2866,N_1750,N_1565);
nor U2867 (N_2867,N_1749,N_1200);
xnor U2868 (N_2868,N_1828,N_1118);
xnor U2869 (N_2869,N_1684,N_1598);
nor U2870 (N_2870,N_1450,N_1520);
and U2871 (N_2871,N_1944,N_1537);
nor U2872 (N_2872,N_1753,N_1435);
nand U2873 (N_2873,N_1130,N_1952);
nand U2874 (N_2874,N_1933,N_1571);
or U2875 (N_2875,N_1836,N_1359);
nand U2876 (N_2876,N_1576,N_1966);
xnor U2877 (N_2877,N_1780,N_1982);
or U2878 (N_2878,N_1819,N_1788);
and U2879 (N_2879,N_1453,N_1027);
xnor U2880 (N_2880,N_1406,N_1669);
nor U2881 (N_2881,N_1397,N_1729);
nand U2882 (N_2882,N_1158,N_1932);
or U2883 (N_2883,N_1349,N_1666);
nand U2884 (N_2884,N_1756,N_1118);
or U2885 (N_2885,N_1259,N_1828);
nor U2886 (N_2886,N_1883,N_1378);
and U2887 (N_2887,N_1959,N_1545);
nand U2888 (N_2888,N_1455,N_1839);
and U2889 (N_2889,N_1292,N_1720);
and U2890 (N_2890,N_1286,N_1083);
nor U2891 (N_2891,N_1560,N_1526);
nand U2892 (N_2892,N_1322,N_1629);
nor U2893 (N_2893,N_1387,N_1020);
xnor U2894 (N_2894,N_1490,N_1407);
nand U2895 (N_2895,N_1294,N_1804);
xnor U2896 (N_2896,N_1527,N_1471);
nor U2897 (N_2897,N_1697,N_1373);
or U2898 (N_2898,N_1176,N_1142);
nor U2899 (N_2899,N_1404,N_1490);
or U2900 (N_2900,N_1181,N_1861);
or U2901 (N_2901,N_1286,N_1521);
xnor U2902 (N_2902,N_1024,N_1546);
or U2903 (N_2903,N_1430,N_1001);
xor U2904 (N_2904,N_1674,N_1488);
and U2905 (N_2905,N_1477,N_1277);
and U2906 (N_2906,N_1412,N_1401);
or U2907 (N_2907,N_1812,N_1344);
and U2908 (N_2908,N_1907,N_1705);
nand U2909 (N_2909,N_1124,N_1323);
xnor U2910 (N_2910,N_1503,N_1495);
and U2911 (N_2911,N_1058,N_1580);
and U2912 (N_2912,N_1976,N_1726);
and U2913 (N_2913,N_1534,N_1189);
nor U2914 (N_2914,N_1584,N_1964);
xnor U2915 (N_2915,N_1503,N_1834);
nand U2916 (N_2916,N_1476,N_1123);
or U2917 (N_2917,N_1918,N_1464);
nor U2918 (N_2918,N_1722,N_1910);
nand U2919 (N_2919,N_1314,N_1464);
nand U2920 (N_2920,N_1932,N_1419);
or U2921 (N_2921,N_1183,N_1237);
and U2922 (N_2922,N_1648,N_1612);
or U2923 (N_2923,N_1158,N_1014);
and U2924 (N_2924,N_1415,N_1292);
and U2925 (N_2925,N_1165,N_1106);
nand U2926 (N_2926,N_1813,N_1182);
or U2927 (N_2927,N_1810,N_1440);
nand U2928 (N_2928,N_1647,N_1173);
or U2929 (N_2929,N_1081,N_1842);
and U2930 (N_2930,N_1462,N_1958);
nor U2931 (N_2931,N_1121,N_1702);
nor U2932 (N_2932,N_1149,N_1123);
nand U2933 (N_2933,N_1365,N_1380);
xnor U2934 (N_2934,N_1795,N_1739);
nor U2935 (N_2935,N_1677,N_1149);
and U2936 (N_2936,N_1521,N_1682);
nand U2937 (N_2937,N_1855,N_1199);
and U2938 (N_2938,N_1844,N_1398);
nor U2939 (N_2939,N_1386,N_1606);
nor U2940 (N_2940,N_1036,N_1857);
nor U2941 (N_2941,N_1505,N_1388);
and U2942 (N_2942,N_1976,N_1105);
or U2943 (N_2943,N_1266,N_1742);
xnor U2944 (N_2944,N_1175,N_1229);
nor U2945 (N_2945,N_1468,N_1583);
xor U2946 (N_2946,N_1825,N_1158);
or U2947 (N_2947,N_1291,N_1249);
nor U2948 (N_2948,N_1194,N_1637);
and U2949 (N_2949,N_1033,N_1255);
xnor U2950 (N_2950,N_1972,N_1063);
xnor U2951 (N_2951,N_1284,N_1363);
nand U2952 (N_2952,N_1277,N_1043);
nand U2953 (N_2953,N_1389,N_1999);
nor U2954 (N_2954,N_1832,N_1837);
or U2955 (N_2955,N_1955,N_1887);
nor U2956 (N_2956,N_1423,N_1860);
nor U2957 (N_2957,N_1878,N_1018);
xor U2958 (N_2958,N_1580,N_1335);
or U2959 (N_2959,N_1501,N_1108);
and U2960 (N_2960,N_1938,N_1482);
and U2961 (N_2961,N_1522,N_1437);
nand U2962 (N_2962,N_1195,N_1024);
or U2963 (N_2963,N_1156,N_1325);
xor U2964 (N_2964,N_1655,N_1521);
xnor U2965 (N_2965,N_1408,N_1923);
nor U2966 (N_2966,N_1066,N_1923);
nand U2967 (N_2967,N_1117,N_1455);
or U2968 (N_2968,N_1680,N_1692);
nor U2969 (N_2969,N_1859,N_1482);
nand U2970 (N_2970,N_1810,N_1144);
and U2971 (N_2971,N_1539,N_1974);
xnor U2972 (N_2972,N_1806,N_1671);
xnor U2973 (N_2973,N_1725,N_1977);
nand U2974 (N_2974,N_1691,N_1976);
xor U2975 (N_2975,N_1596,N_1918);
and U2976 (N_2976,N_1234,N_1363);
nor U2977 (N_2977,N_1885,N_1358);
xor U2978 (N_2978,N_1582,N_1677);
and U2979 (N_2979,N_1284,N_1373);
nor U2980 (N_2980,N_1797,N_1251);
nand U2981 (N_2981,N_1673,N_1728);
and U2982 (N_2982,N_1920,N_1530);
or U2983 (N_2983,N_1410,N_1847);
or U2984 (N_2984,N_1018,N_1488);
and U2985 (N_2985,N_1194,N_1473);
nor U2986 (N_2986,N_1018,N_1326);
and U2987 (N_2987,N_1376,N_1062);
or U2988 (N_2988,N_1058,N_1134);
nand U2989 (N_2989,N_1923,N_1761);
xor U2990 (N_2990,N_1503,N_1482);
or U2991 (N_2991,N_1761,N_1541);
nand U2992 (N_2992,N_1830,N_1831);
nor U2993 (N_2993,N_1938,N_1143);
or U2994 (N_2994,N_1642,N_1778);
and U2995 (N_2995,N_1133,N_1344);
nor U2996 (N_2996,N_1139,N_1754);
nand U2997 (N_2997,N_1862,N_1950);
nand U2998 (N_2998,N_1153,N_1480);
nor U2999 (N_2999,N_1266,N_1141);
nand U3000 (N_3000,N_2534,N_2494);
nor U3001 (N_3001,N_2116,N_2679);
xor U3002 (N_3002,N_2815,N_2895);
or U3003 (N_3003,N_2404,N_2170);
or U3004 (N_3004,N_2532,N_2673);
nor U3005 (N_3005,N_2977,N_2531);
nor U3006 (N_3006,N_2466,N_2102);
or U3007 (N_3007,N_2600,N_2659);
and U3008 (N_3008,N_2546,N_2749);
nand U3009 (N_3009,N_2829,N_2548);
nor U3010 (N_3010,N_2806,N_2143);
or U3011 (N_3011,N_2629,N_2223);
or U3012 (N_3012,N_2471,N_2952);
nand U3013 (N_3013,N_2052,N_2825);
or U3014 (N_3014,N_2293,N_2299);
xnor U3015 (N_3015,N_2908,N_2281);
nand U3016 (N_3016,N_2300,N_2707);
nor U3017 (N_3017,N_2058,N_2426);
nor U3018 (N_3018,N_2236,N_2942);
nor U3019 (N_3019,N_2918,N_2044);
xor U3020 (N_3020,N_2482,N_2190);
or U3021 (N_3021,N_2203,N_2919);
nor U3022 (N_3022,N_2779,N_2422);
nand U3023 (N_3023,N_2269,N_2944);
nand U3024 (N_3024,N_2148,N_2138);
nor U3025 (N_3025,N_2978,N_2872);
nor U3026 (N_3026,N_2561,N_2086);
xnor U3027 (N_3027,N_2569,N_2354);
xor U3028 (N_3028,N_2960,N_2664);
xnor U3029 (N_3029,N_2896,N_2674);
and U3030 (N_3030,N_2245,N_2683);
xor U3031 (N_3031,N_2722,N_2270);
and U3032 (N_3032,N_2807,N_2405);
nand U3033 (N_3033,N_2400,N_2470);
or U3034 (N_3034,N_2828,N_2322);
nand U3035 (N_3035,N_2831,N_2994);
nor U3036 (N_3036,N_2115,N_2154);
and U3037 (N_3037,N_2634,N_2278);
and U3038 (N_3038,N_2816,N_2981);
nor U3039 (N_3039,N_2196,N_2976);
or U3040 (N_3040,N_2018,N_2056);
nor U3041 (N_3041,N_2847,N_2456);
and U3042 (N_3042,N_2624,N_2262);
and U3043 (N_3043,N_2787,N_2947);
nor U3044 (N_3044,N_2802,N_2121);
xor U3045 (N_3045,N_2195,N_2067);
nor U3046 (N_3046,N_2810,N_2536);
nor U3047 (N_3047,N_2805,N_2938);
nor U3048 (N_3048,N_2134,N_2343);
or U3049 (N_3049,N_2392,N_2220);
nand U3050 (N_3050,N_2845,N_2497);
nor U3051 (N_3051,N_2479,N_2450);
nor U3052 (N_3052,N_2601,N_2793);
nor U3053 (N_3053,N_2508,N_2698);
nand U3054 (N_3054,N_2791,N_2920);
xnor U3055 (N_3055,N_2595,N_2326);
or U3056 (N_3056,N_2417,N_2019);
nor U3057 (N_3057,N_2886,N_2352);
nor U3058 (N_3058,N_2016,N_2999);
xor U3059 (N_3059,N_2525,N_2452);
nor U3060 (N_3060,N_2499,N_2204);
and U3061 (N_3061,N_2515,N_2898);
nor U3062 (N_3062,N_2715,N_2020);
and U3063 (N_3063,N_2335,N_2611);
xnor U3064 (N_3064,N_2453,N_2260);
xor U3065 (N_3065,N_2932,N_2321);
or U3066 (N_3066,N_2647,N_2975);
nand U3067 (N_3067,N_2788,N_2137);
nand U3068 (N_3068,N_2147,N_2306);
nand U3069 (N_3069,N_2033,N_2133);
xnor U3070 (N_3070,N_2751,N_2042);
nand U3071 (N_3071,N_2481,N_2703);
xnor U3072 (N_3072,N_2850,N_2357);
or U3073 (N_3073,N_2192,N_2748);
nor U3074 (N_3074,N_2583,N_2053);
or U3075 (N_3075,N_2129,N_2030);
or U3076 (N_3076,N_2239,N_2567);
and U3077 (N_3077,N_2199,N_2012);
or U3078 (N_3078,N_2238,N_2750);
nor U3079 (N_3079,N_2607,N_2724);
and U3080 (N_3080,N_2465,N_2159);
nand U3081 (N_3081,N_2063,N_2535);
and U3082 (N_3082,N_2693,N_2430);
nor U3083 (N_3083,N_2903,N_2819);
nor U3084 (N_3084,N_2930,N_2101);
or U3085 (N_3085,N_2440,N_2575);
nand U3086 (N_3086,N_2565,N_2760);
or U3087 (N_3087,N_2311,N_2165);
nor U3088 (N_3088,N_2141,N_2467);
or U3089 (N_3089,N_2710,N_2506);
or U3090 (N_3090,N_2527,N_2718);
xnor U3091 (N_3091,N_2074,N_2295);
nand U3092 (N_3092,N_2432,N_2388);
and U3093 (N_3093,N_2226,N_2686);
xnor U3094 (N_3094,N_2604,N_2231);
nor U3095 (N_3095,N_2857,N_2860);
xnor U3096 (N_3096,N_2741,N_2248);
or U3097 (N_3097,N_2498,N_2089);
nand U3098 (N_3098,N_2969,N_2539);
or U3099 (N_3099,N_2706,N_2312);
nand U3100 (N_3100,N_2491,N_2655);
and U3101 (N_3101,N_2980,N_2642);
nor U3102 (N_3102,N_2556,N_2717);
xnor U3103 (N_3103,N_2317,N_2474);
nand U3104 (N_3104,N_2237,N_2837);
xor U3105 (N_3105,N_2692,N_2729);
xor U3106 (N_3106,N_2639,N_2576);
or U3107 (N_3107,N_2761,N_2219);
and U3108 (N_3108,N_2200,N_2080);
nand U3109 (N_3109,N_2992,N_2325);
nand U3110 (N_3110,N_2475,N_2571);
nand U3111 (N_3111,N_2855,N_2023);
nor U3112 (N_3112,N_2586,N_2946);
nor U3113 (N_3113,N_2821,N_2669);
and U3114 (N_3114,N_2330,N_2924);
or U3115 (N_3115,N_2570,N_2684);
nand U3116 (N_3116,N_2566,N_2769);
or U3117 (N_3117,N_2770,N_2716);
xnor U3118 (N_3118,N_2983,N_2344);
and U3119 (N_3119,N_2839,N_2910);
or U3120 (N_3120,N_2727,N_2774);
xor U3121 (N_3121,N_2222,N_2229);
or U3122 (N_3122,N_2383,N_2504);
and U3123 (N_3123,N_2112,N_2078);
and U3124 (N_3124,N_2447,N_2364);
nor U3125 (N_3125,N_2830,N_2146);
and U3126 (N_3126,N_2641,N_2161);
xnor U3127 (N_3127,N_2778,N_2500);
xnor U3128 (N_3128,N_2909,N_2984);
nor U3129 (N_3129,N_2652,N_2153);
nand U3130 (N_3130,N_2290,N_2336);
and U3131 (N_3131,N_2657,N_2179);
nand U3132 (N_3132,N_2926,N_2893);
and U3133 (N_3133,N_2851,N_2766);
nand U3134 (N_3134,N_2773,N_2109);
nor U3135 (N_3135,N_2676,N_2472);
and U3136 (N_3136,N_2826,N_2093);
nor U3137 (N_3137,N_2462,N_2796);
and U3138 (N_3138,N_2419,N_2970);
nand U3139 (N_3139,N_2987,N_2218);
and U3140 (N_3140,N_2890,N_2785);
xnor U3141 (N_3141,N_2743,N_2072);
nand U3142 (N_3142,N_2734,N_2823);
or U3143 (N_3143,N_2907,N_2927);
or U3144 (N_3144,N_2603,N_2360);
nor U3145 (N_3145,N_2243,N_2911);
or U3146 (N_3146,N_2297,N_2764);
and U3147 (N_3147,N_2635,N_2398);
or U3148 (N_3148,N_2117,N_2084);
nor U3149 (N_3149,N_2097,N_2241);
xnor U3150 (N_3150,N_2746,N_2547);
xnor U3151 (N_3151,N_2233,N_2616);
and U3152 (N_3152,N_2509,N_2054);
and U3153 (N_3153,N_2041,N_2458);
nand U3154 (N_3154,N_2198,N_2666);
and U3155 (N_3155,N_2971,N_2363);
nor U3156 (N_3156,N_2412,N_2661);
nand U3157 (N_3157,N_2221,N_2224);
and U3158 (N_3158,N_2866,N_2160);
nand U3159 (N_3159,N_2202,N_2988);
xnor U3160 (N_3160,N_2242,N_2800);
nor U3161 (N_3161,N_2542,N_2162);
nand U3162 (N_3162,N_2521,N_2653);
or U3163 (N_3163,N_2613,N_2838);
or U3164 (N_3164,N_2768,N_2172);
and U3165 (N_3165,N_2913,N_2522);
or U3166 (N_3166,N_2956,N_2714);
nor U3167 (N_3167,N_2752,N_2758);
and U3168 (N_3168,N_2277,N_2985);
xnor U3169 (N_3169,N_2377,N_2777);
or U3170 (N_3170,N_2094,N_2873);
and U3171 (N_3171,N_2756,N_2891);
xnor U3172 (N_3172,N_2959,N_2549);
and U3173 (N_3173,N_2687,N_2541);
nand U3174 (N_3174,N_2520,N_2079);
nand U3175 (N_3175,N_2010,N_2348);
and U3176 (N_3176,N_2071,N_2875);
xor U3177 (N_3177,N_2393,N_2407);
or U3178 (N_3178,N_2609,N_2197);
nor U3179 (N_3179,N_2883,N_2037);
nor U3180 (N_3180,N_2767,N_2399);
xnor U3181 (N_3181,N_2713,N_2022);
nor U3182 (N_3182,N_2083,N_2708);
xor U3183 (N_3183,N_2511,N_2662);
nor U3184 (N_3184,N_2411,N_2776);
or U3185 (N_3185,N_2421,N_2418);
or U3186 (N_3186,N_2107,N_2914);
or U3187 (N_3187,N_2711,N_2606);
and U3188 (N_3188,N_2637,N_2897);
xor U3189 (N_3189,N_2283,N_2077);
nand U3190 (N_3190,N_2289,N_2617);
xor U3191 (N_3191,N_2332,N_2867);
xnor U3192 (N_3192,N_2291,N_2486);
xor U3193 (N_3193,N_2665,N_2904);
nor U3194 (N_3194,N_2763,N_2982);
or U3195 (N_3195,N_2518,N_2061);
xor U3196 (N_3196,N_2303,N_2285);
or U3197 (N_3197,N_2186,N_2414);
and U3198 (N_3198,N_2574,N_2091);
or U3199 (N_3199,N_2730,N_2582);
or U3200 (N_3200,N_2870,N_2517);
nor U3201 (N_3201,N_2279,N_2436);
xnor U3202 (N_3202,N_2113,N_2118);
nand U3203 (N_3203,N_2028,N_2869);
nor U3204 (N_3204,N_2728,N_2205);
xor U3205 (N_3205,N_2699,N_2468);
xor U3206 (N_3206,N_2187,N_2055);
nor U3207 (N_3207,N_2599,N_2428);
xnor U3208 (N_3208,N_2085,N_2382);
xor U3209 (N_3209,N_2409,N_2573);
nor U3210 (N_3210,N_2214,N_2130);
or U3211 (N_3211,N_2865,N_2258);
nor U3212 (N_3212,N_2502,N_2394);
xnor U3213 (N_3213,N_2705,N_2308);
nor U3214 (N_3214,N_2098,N_2167);
and U3215 (N_3215,N_2431,N_2358);
nor U3216 (N_3216,N_2709,N_2644);
or U3217 (N_3217,N_2524,N_2043);
nand U3218 (N_3218,N_2965,N_2658);
nor U3219 (N_3219,N_2680,N_2026);
xor U3220 (N_3220,N_2798,N_2366);
and U3221 (N_3221,N_2783,N_2164);
nor U3222 (N_3222,N_2885,N_2862);
xor U3223 (N_3223,N_2068,N_2349);
and U3224 (N_3224,N_2045,N_2048);
xor U3225 (N_3225,N_2073,N_2145);
and U3226 (N_3226,N_2100,N_2027);
nand U3227 (N_3227,N_2671,N_2941);
or U3228 (N_3228,N_2381,N_2631);
or U3229 (N_3229,N_2670,N_2998);
nand U3230 (N_3230,N_2681,N_2024);
nand U3231 (N_3231,N_2577,N_2917);
xor U3232 (N_3232,N_2545,N_2070);
nand U3233 (N_3233,N_2782,N_2081);
xnor U3234 (N_3234,N_2386,N_2902);
nor U3235 (N_3235,N_2943,N_2700);
xor U3236 (N_3236,N_2150,N_2212);
xor U3237 (N_3237,N_2841,N_2046);
nor U3238 (N_3238,N_2808,N_2822);
and U3239 (N_3239,N_2813,N_2678);
or U3240 (N_3240,N_2844,N_2995);
nor U3241 (N_3241,N_2209,N_2090);
nand U3242 (N_3242,N_2612,N_2721);
xnor U3243 (N_3243,N_2302,N_2744);
or U3244 (N_3244,N_2039,N_2811);
and U3245 (N_3245,N_2395,N_2255);
nor U3246 (N_3246,N_2923,N_2110);
nor U3247 (N_3247,N_2413,N_2415);
or U3248 (N_3248,N_2305,N_2244);
nand U3249 (N_3249,N_2435,N_2194);
xnor U3250 (N_3250,N_2921,N_2859);
nor U3251 (N_3251,N_2126,N_2925);
xnor U3252 (N_3252,N_2256,N_2848);
nand U3253 (N_3253,N_2207,N_2530);
or U3254 (N_3254,N_2120,N_2775);
nand U3255 (N_3255,N_2350,N_2286);
xnor U3256 (N_3256,N_2342,N_2814);
and U3257 (N_3257,N_2799,N_2628);
nor U3258 (N_3258,N_2257,N_2972);
xor U3259 (N_3259,N_2476,N_2391);
nand U3260 (N_3260,N_2210,N_2062);
nor U3261 (N_3261,N_2996,N_2442);
and U3262 (N_3262,N_2108,N_2296);
xor U3263 (N_3263,N_2585,N_2533);
nand U3264 (N_3264,N_2501,N_2884);
xor U3265 (N_3265,N_2333,N_2832);
xnor U3266 (N_3266,N_2614,N_2651);
and U3267 (N_3267,N_2217,N_2955);
and U3268 (N_3268,N_2177,N_2967);
nor U3269 (N_3269,N_2341,N_2590);
or U3270 (N_3270,N_2185,N_2092);
or U3271 (N_3271,N_2310,N_2964);
and U3272 (N_3272,N_2438,N_2630);
and U3273 (N_3273,N_2201,N_2408);
and U3274 (N_3274,N_2123,N_2000);
xor U3275 (N_3275,N_2275,N_2818);
or U3276 (N_3276,N_2294,N_2578);
xnor U3277 (N_3277,N_2892,N_2228);
nand U3278 (N_3278,N_2009,N_2958);
xnor U3279 (N_3279,N_2781,N_2842);
nand U3280 (N_3280,N_2166,N_2211);
and U3281 (N_3281,N_2564,N_2880);
nor U3282 (N_3282,N_2227,N_2608);
or U3283 (N_3283,N_2368,N_2650);
nor U3284 (N_3284,N_2874,N_2329);
nor U3285 (N_3285,N_2712,N_2929);
nand U3286 (N_3286,N_2966,N_2347);
or U3287 (N_3287,N_2151,N_2789);
nor U3288 (N_3288,N_2663,N_2261);
nand U3289 (N_3289,N_2206,N_2621);
nor U3290 (N_3290,N_2933,N_2922);
and U3291 (N_3291,N_2240,N_2552);
and U3292 (N_3292,N_2375,N_2493);
nand U3293 (N_3293,N_2455,N_2139);
or U3294 (N_3294,N_2991,N_2304);
or U3295 (N_3295,N_2719,N_2581);
or U3296 (N_3296,N_2979,N_2973);
xnor U3297 (N_3297,N_2370,N_2274);
xnor U3298 (N_3298,N_2250,N_2373);
xnor U3299 (N_3299,N_2060,N_2340);
xnor U3300 (N_3300,N_2230,N_2132);
or U3301 (N_3301,N_2036,N_2439);
nor U3302 (N_3302,N_2843,N_2131);
nand U3303 (N_3303,N_2178,N_2812);
nand U3304 (N_3304,N_2423,N_2868);
and U3305 (N_3305,N_2954,N_2646);
and U3306 (N_3306,N_2588,N_2265);
or U3307 (N_3307,N_2881,N_2849);
and U3308 (N_3308,N_2754,N_2735);
xnor U3309 (N_3309,N_2945,N_2272);
xor U3310 (N_3310,N_2739,N_2801);
nand U3311 (N_3311,N_2753,N_2013);
xor U3312 (N_3312,N_2402,N_2319);
nand U3313 (N_3313,N_2794,N_2594);
xor U3314 (N_3314,N_2840,N_2096);
xor U3315 (N_3315,N_2864,N_2856);
or U3316 (N_3316,N_2015,N_2526);
nor U3317 (N_3317,N_2353,N_2136);
nand U3318 (N_3318,N_2733,N_2915);
or U3319 (N_3319,N_2732,N_2605);
or U3320 (N_3320,N_2029,N_2280);
xnor U3321 (N_3321,N_2620,N_2731);
or U3322 (N_3322,N_2682,N_2528);
and U3323 (N_3323,N_2276,N_2420);
xnor U3324 (N_3324,N_2047,N_2636);
and U3325 (N_3325,N_2384,N_2064);
nor U3326 (N_3326,N_2858,N_2899);
nor U3327 (N_3327,N_2017,N_2745);
xor U3328 (N_3328,N_2820,N_2189);
or U3329 (N_3329,N_2809,N_2490);
or U3330 (N_3330,N_2580,N_2579);
or U3331 (N_3331,N_2460,N_2057);
or U3332 (N_3332,N_2505,N_2403);
xnor U3333 (N_3333,N_2378,N_2372);
nor U3334 (N_3334,N_2066,N_2193);
and U3335 (N_3335,N_2355,N_2318);
and U3336 (N_3336,N_2689,N_2558);
nand U3337 (N_3337,N_2263,N_2288);
xnor U3338 (N_3338,N_2327,N_2495);
xnor U3339 (N_3339,N_2448,N_2292);
xor U3340 (N_3340,N_2759,N_2677);
xnor U3341 (N_3341,N_2804,N_2485);
nand U3342 (N_3342,N_2551,N_2633);
nand U3343 (N_3343,N_2792,N_2598);
xnor U3344 (N_3344,N_2174,N_2704);
nor U3345 (N_3345,N_2443,N_2050);
nor U3346 (N_3346,N_2688,N_2592);
and U3347 (N_3347,N_2171,N_2181);
nor U3348 (N_3348,N_2152,N_2338);
nand U3349 (N_3349,N_2668,N_2445);
nand U3350 (N_3350,N_2254,N_2496);
or U3351 (N_3351,N_2374,N_2401);
and U3352 (N_3352,N_2544,N_2345);
or U3353 (N_3353,N_2114,N_2213);
xnor U3354 (N_3354,N_2622,N_2519);
nand U3355 (N_3355,N_2314,N_2259);
nor U3356 (N_3356,N_2315,N_2961);
nand U3357 (N_3357,N_2584,N_2572);
and U3358 (N_3358,N_2597,N_2088);
nand U3359 (N_3359,N_2540,N_2111);
xnor U3360 (N_3360,N_2901,N_2183);
nand U3361 (N_3361,N_2948,N_2216);
or U3362 (N_3362,N_2287,N_2461);
and U3363 (N_3363,N_2361,N_2469);
nand U3364 (N_3364,N_2833,N_2747);
nor U3365 (N_3365,N_2169,N_2429);
and U3366 (N_3366,N_2021,N_2514);
and U3367 (N_3367,N_2626,N_2695);
or U3368 (N_3368,N_2191,N_2997);
nor U3369 (N_3369,N_2034,N_2182);
nor U3370 (N_3370,N_2334,N_2007);
and U3371 (N_3371,N_2173,N_2852);
nor U3372 (N_3372,N_2691,N_2433);
and U3373 (N_3373,N_2035,N_2434);
and U3374 (N_3374,N_2477,N_2284);
xnor U3375 (N_3375,N_2484,N_2784);
and U3376 (N_3376,N_2742,N_2723);
or U3377 (N_3377,N_2672,N_2268);
or U3378 (N_3378,N_2425,N_2974);
and U3379 (N_3379,N_2105,N_2158);
xnor U3380 (N_3380,N_2615,N_2876);
nand U3381 (N_3381,N_2369,N_2135);
or U3382 (N_3382,N_2008,N_2301);
nand U3383 (N_3383,N_2376,N_2738);
nand U3384 (N_3384,N_2627,N_2990);
nor U3385 (N_3385,N_2643,N_2038);
nor U3386 (N_3386,N_2379,N_2632);
nor U3387 (N_3387,N_2963,N_2937);
xor U3388 (N_3388,N_2444,N_2264);
xnor U3389 (N_3389,N_2790,N_2025);
xnor U3390 (N_3390,N_2266,N_2957);
xnor U3391 (N_3391,N_2331,N_2095);
nand U3392 (N_3392,N_2451,N_2441);
nand U3393 (N_3393,N_2503,N_2916);
or U3394 (N_3394,N_2313,N_2877);
nand U3395 (N_3395,N_2690,N_2140);
and U3396 (N_3396,N_2675,N_2654);
xor U3397 (N_3397,N_2619,N_2473);
and U3398 (N_3398,N_2065,N_2529);
nor U3399 (N_3399,N_2625,N_2523);
and U3400 (N_3400,N_2596,N_2168);
xnor U3401 (N_3401,N_2051,N_2762);
and U3402 (N_3402,N_2853,N_2246);
xor U3403 (N_3403,N_2765,N_2737);
xor U3404 (N_3404,N_2049,N_2149);
or U3405 (N_3405,N_2568,N_2871);
xnor U3406 (N_3406,N_2492,N_2934);
xor U3407 (N_3407,N_2755,N_2188);
nor U3408 (N_3408,N_2390,N_2396);
xor U3409 (N_3409,N_2176,N_2128);
nand U3410 (N_3410,N_2235,N_2795);
nand U3411 (N_3411,N_2253,N_2771);
nor U3412 (N_3412,N_2273,N_2488);
nor U3413 (N_3413,N_2968,N_2487);
xnor U3414 (N_3414,N_2427,N_2082);
or U3415 (N_3415,N_2252,N_2559);
nand U3416 (N_3416,N_2157,N_2513);
xor U3417 (N_3417,N_2075,N_2457);
nor U3418 (N_3418,N_2483,N_2339);
nand U3419 (N_3419,N_2316,N_2180);
nand U3420 (N_3420,N_2410,N_2175);
or U3421 (N_3421,N_2900,N_2122);
and U3422 (N_3422,N_2725,N_2824);
and U3423 (N_3423,N_2538,N_2562);
xnor U3424 (N_3424,N_2645,N_2602);
xor U3425 (N_3425,N_2772,N_2298);
nor U3426 (N_3426,N_2359,N_2702);
xor U3427 (N_3427,N_2649,N_2424);
nor U3428 (N_3428,N_2014,N_2463);
nand U3429 (N_3429,N_2416,N_2104);
nand U3430 (N_3430,N_2356,N_2454);
or U3431 (N_3431,N_2863,N_2726);
nor U3432 (N_3432,N_2163,N_2587);
nand U3433 (N_3433,N_2685,N_2124);
nand U3434 (N_3434,N_2593,N_2931);
xnor U3435 (N_3435,N_2701,N_2406);
nor U3436 (N_3436,N_2640,N_2003);
and U3437 (N_3437,N_2951,N_2371);
nor U3438 (N_3438,N_2879,N_2786);
and U3439 (N_3439,N_2106,N_2251);
nand U3440 (N_3440,N_2127,N_2510);
nand U3441 (N_3441,N_2385,N_2362);
or U3442 (N_3442,N_2489,N_2367);
and U3443 (N_3443,N_2119,N_2512);
or U3444 (N_3444,N_2365,N_2537);
nor U3445 (N_3445,N_2249,N_2660);
nand U3446 (N_3446,N_2397,N_2940);
or U3447 (N_3447,N_2797,N_2480);
or U3448 (N_3448,N_2834,N_2953);
xor U3449 (N_3449,N_2835,N_2610);
or U3450 (N_3450,N_2803,N_2031);
and U3451 (N_3451,N_2667,N_2032);
nor U3452 (N_3452,N_2912,N_2889);
nor U3453 (N_3453,N_2069,N_2320);
nor U3454 (N_3454,N_2950,N_2648);
nand U3455 (N_3455,N_2271,N_2516);
nor U3456 (N_3456,N_2696,N_2697);
and U3457 (N_3457,N_2328,N_2142);
nor U3458 (N_3458,N_2215,N_2346);
nand U3459 (N_3459,N_2888,N_2155);
and U3460 (N_3460,N_2076,N_2861);
and U3461 (N_3461,N_2004,N_2905);
nor U3462 (N_3462,N_2935,N_2001);
nand U3463 (N_3463,N_2459,N_2543);
nor U3464 (N_3464,N_2591,N_2232);
nor U3465 (N_3465,N_2894,N_2618);
and U3466 (N_3466,N_2507,N_2555);
or U3467 (N_3467,N_2740,N_2234);
nand U3468 (N_3468,N_2993,N_2125);
nor U3469 (N_3469,N_2208,N_2817);
nor U3470 (N_3470,N_2040,N_2656);
nand U3471 (N_3471,N_2059,N_2309);
nand U3472 (N_3472,N_2846,N_2560);
or U3473 (N_3473,N_2736,N_2389);
or U3474 (N_3474,N_2836,N_2557);
nand U3475 (N_3475,N_2184,N_2247);
xor U3476 (N_3476,N_2553,N_2225);
and U3477 (N_3477,N_2156,N_2387);
or U3478 (N_3478,N_2323,N_2906);
nor U3479 (N_3479,N_2554,N_2854);
and U3480 (N_3480,N_2936,N_2337);
and U3481 (N_3481,N_2589,N_2437);
or U3482 (N_3482,N_2011,N_2478);
nor U3483 (N_3483,N_2962,N_2757);
nor U3484 (N_3484,N_2720,N_2986);
or U3485 (N_3485,N_2694,N_2638);
nand U3486 (N_3486,N_2887,N_2006);
and U3487 (N_3487,N_2282,N_2780);
and U3488 (N_3488,N_2563,N_2103);
nor U3489 (N_3489,N_2550,N_2324);
or U3490 (N_3490,N_2449,N_2351);
or U3491 (N_3491,N_2882,N_2827);
xnor U3492 (N_3492,N_2446,N_2380);
xnor U3493 (N_3493,N_2144,N_2878);
xnor U3494 (N_3494,N_2099,N_2939);
xnor U3495 (N_3495,N_2623,N_2464);
or U3496 (N_3496,N_2267,N_2989);
xor U3497 (N_3497,N_2002,N_2005);
and U3498 (N_3498,N_2087,N_2949);
nor U3499 (N_3499,N_2928,N_2307);
nor U3500 (N_3500,N_2032,N_2525);
nor U3501 (N_3501,N_2378,N_2311);
xnor U3502 (N_3502,N_2588,N_2765);
and U3503 (N_3503,N_2767,N_2671);
or U3504 (N_3504,N_2831,N_2763);
and U3505 (N_3505,N_2885,N_2927);
nand U3506 (N_3506,N_2026,N_2476);
or U3507 (N_3507,N_2857,N_2383);
nor U3508 (N_3508,N_2153,N_2494);
or U3509 (N_3509,N_2348,N_2236);
nand U3510 (N_3510,N_2621,N_2425);
nand U3511 (N_3511,N_2535,N_2686);
nand U3512 (N_3512,N_2913,N_2827);
nand U3513 (N_3513,N_2600,N_2090);
nor U3514 (N_3514,N_2154,N_2100);
and U3515 (N_3515,N_2863,N_2355);
and U3516 (N_3516,N_2084,N_2879);
xor U3517 (N_3517,N_2688,N_2414);
xor U3518 (N_3518,N_2600,N_2310);
xnor U3519 (N_3519,N_2080,N_2674);
and U3520 (N_3520,N_2183,N_2363);
and U3521 (N_3521,N_2236,N_2870);
or U3522 (N_3522,N_2688,N_2845);
and U3523 (N_3523,N_2232,N_2298);
nand U3524 (N_3524,N_2254,N_2740);
or U3525 (N_3525,N_2616,N_2986);
nand U3526 (N_3526,N_2230,N_2176);
nand U3527 (N_3527,N_2464,N_2922);
nand U3528 (N_3528,N_2263,N_2633);
or U3529 (N_3529,N_2235,N_2968);
or U3530 (N_3530,N_2045,N_2415);
or U3531 (N_3531,N_2759,N_2451);
xnor U3532 (N_3532,N_2577,N_2767);
and U3533 (N_3533,N_2099,N_2363);
nand U3534 (N_3534,N_2334,N_2842);
xnor U3535 (N_3535,N_2987,N_2571);
nor U3536 (N_3536,N_2677,N_2673);
xor U3537 (N_3537,N_2164,N_2547);
nor U3538 (N_3538,N_2741,N_2414);
and U3539 (N_3539,N_2062,N_2545);
or U3540 (N_3540,N_2944,N_2208);
xor U3541 (N_3541,N_2712,N_2622);
or U3542 (N_3542,N_2635,N_2340);
or U3543 (N_3543,N_2213,N_2705);
nand U3544 (N_3544,N_2780,N_2510);
or U3545 (N_3545,N_2145,N_2619);
or U3546 (N_3546,N_2061,N_2366);
nand U3547 (N_3547,N_2261,N_2596);
and U3548 (N_3548,N_2561,N_2305);
nor U3549 (N_3549,N_2289,N_2194);
nor U3550 (N_3550,N_2811,N_2441);
or U3551 (N_3551,N_2283,N_2523);
and U3552 (N_3552,N_2633,N_2251);
nor U3553 (N_3553,N_2916,N_2470);
xor U3554 (N_3554,N_2528,N_2315);
xor U3555 (N_3555,N_2746,N_2662);
xnor U3556 (N_3556,N_2807,N_2467);
or U3557 (N_3557,N_2476,N_2444);
nor U3558 (N_3558,N_2683,N_2851);
and U3559 (N_3559,N_2273,N_2549);
nor U3560 (N_3560,N_2070,N_2072);
xnor U3561 (N_3561,N_2674,N_2669);
and U3562 (N_3562,N_2397,N_2959);
nand U3563 (N_3563,N_2684,N_2643);
xnor U3564 (N_3564,N_2472,N_2090);
and U3565 (N_3565,N_2558,N_2764);
or U3566 (N_3566,N_2804,N_2208);
nand U3567 (N_3567,N_2914,N_2275);
and U3568 (N_3568,N_2018,N_2638);
nand U3569 (N_3569,N_2471,N_2898);
and U3570 (N_3570,N_2791,N_2440);
nor U3571 (N_3571,N_2671,N_2528);
and U3572 (N_3572,N_2757,N_2304);
nor U3573 (N_3573,N_2999,N_2973);
nor U3574 (N_3574,N_2501,N_2403);
or U3575 (N_3575,N_2790,N_2583);
and U3576 (N_3576,N_2039,N_2179);
nor U3577 (N_3577,N_2728,N_2967);
nor U3578 (N_3578,N_2457,N_2115);
and U3579 (N_3579,N_2907,N_2292);
xor U3580 (N_3580,N_2573,N_2939);
nand U3581 (N_3581,N_2335,N_2317);
nand U3582 (N_3582,N_2776,N_2490);
or U3583 (N_3583,N_2378,N_2273);
or U3584 (N_3584,N_2146,N_2495);
and U3585 (N_3585,N_2366,N_2833);
and U3586 (N_3586,N_2599,N_2038);
and U3587 (N_3587,N_2564,N_2023);
nor U3588 (N_3588,N_2025,N_2859);
and U3589 (N_3589,N_2628,N_2817);
nor U3590 (N_3590,N_2168,N_2002);
xnor U3591 (N_3591,N_2388,N_2858);
and U3592 (N_3592,N_2198,N_2392);
nand U3593 (N_3593,N_2979,N_2330);
and U3594 (N_3594,N_2203,N_2437);
and U3595 (N_3595,N_2463,N_2221);
and U3596 (N_3596,N_2478,N_2198);
xnor U3597 (N_3597,N_2162,N_2666);
nor U3598 (N_3598,N_2488,N_2189);
nor U3599 (N_3599,N_2328,N_2876);
and U3600 (N_3600,N_2049,N_2770);
nand U3601 (N_3601,N_2635,N_2248);
nand U3602 (N_3602,N_2025,N_2378);
xnor U3603 (N_3603,N_2888,N_2201);
nand U3604 (N_3604,N_2485,N_2438);
nor U3605 (N_3605,N_2893,N_2002);
or U3606 (N_3606,N_2898,N_2712);
nand U3607 (N_3607,N_2365,N_2504);
or U3608 (N_3608,N_2599,N_2176);
nand U3609 (N_3609,N_2387,N_2191);
nor U3610 (N_3610,N_2528,N_2362);
nor U3611 (N_3611,N_2434,N_2438);
nor U3612 (N_3612,N_2819,N_2972);
and U3613 (N_3613,N_2809,N_2205);
or U3614 (N_3614,N_2140,N_2829);
and U3615 (N_3615,N_2421,N_2286);
nand U3616 (N_3616,N_2452,N_2791);
nor U3617 (N_3617,N_2794,N_2078);
and U3618 (N_3618,N_2243,N_2121);
xnor U3619 (N_3619,N_2786,N_2611);
nand U3620 (N_3620,N_2918,N_2398);
nor U3621 (N_3621,N_2155,N_2392);
and U3622 (N_3622,N_2014,N_2521);
xnor U3623 (N_3623,N_2327,N_2416);
xnor U3624 (N_3624,N_2624,N_2661);
or U3625 (N_3625,N_2105,N_2568);
nand U3626 (N_3626,N_2088,N_2380);
or U3627 (N_3627,N_2988,N_2915);
or U3628 (N_3628,N_2697,N_2348);
xnor U3629 (N_3629,N_2093,N_2019);
xor U3630 (N_3630,N_2134,N_2169);
nand U3631 (N_3631,N_2204,N_2136);
nor U3632 (N_3632,N_2156,N_2964);
or U3633 (N_3633,N_2866,N_2932);
and U3634 (N_3634,N_2397,N_2400);
nor U3635 (N_3635,N_2734,N_2097);
nor U3636 (N_3636,N_2145,N_2391);
and U3637 (N_3637,N_2002,N_2804);
xor U3638 (N_3638,N_2177,N_2048);
xor U3639 (N_3639,N_2487,N_2316);
nand U3640 (N_3640,N_2895,N_2124);
xor U3641 (N_3641,N_2747,N_2332);
or U3642 (N_3642,N_2513,N_2250);
nor U3643 (N_3643,N_2948,N_2145);
nand U3644 (N_3644,N_2911,N_2313);
nor U3645 (N_3645,N_2932,N_2410);
and U3646 (N_3646,N_2207,N_2811);
or U3647 (N_3647,N_2928,N_2748);
nand U3648 (N_3648,N_2187,N_2904);
nand U3649 (N_3649,N_2627,N_2304);
or U3650 (N_3650,N_2963,N_2135);
xnor U3651 (N_3651,N_2720,N_2687);
nor U3652 (N_3652,N_2452,N_2953);
xnor U3653 (N_3653,N_2416,N_2065);
xor U3654 (N_3654,N_2651,N_2412);
xnor U3655 (N_3655,N_2518,N_2363);
nor U3656 (N_3656,N_2774,N_2953);
nand U3657 (N_3657,N_2960,N_2128);
or U3658 (N_3658,N_2553,N_2802);
nor U3659 (N_3659,N_2129,N_2211);
nand U3660 (N_3660,N_2073,N_2911);
and U3661 (N_3661,N_2713,N_2673);
nand U3662 (N_3662,N_2072,N_2103);
and U3663 (N_3663,N_2700,N_2218);
nor U3664 (N_3664,N_2529,N_2116);
nand U3665 (N_3665,N_2737,N_2746);
or U3666 (N_3666,N_2587,N_2497);
or U3667 (N_3667,N_2975,N_2805);
and U3668 (N_3668,N_2734,N_2631);
nor U3669 (N_3669,N_2573,N_2980);
or U3670 (N_3670,N_2557,N_2130);
and U3671 (N_3671,N_2149,N_2836);
and U3672 (N_3672,N_2520,N_2387);
and U3673 (N_3673,N_2153,N_2977);
xor U3674 (N_3674,N_2170,N_2683);
xnor U3675 (N_3675,N_2303,N_2641);
xor U3676 (N_3676,N_2145,N_2613);
xnor U3677 (N_3677,N_2076,N_2088);
xor U3678 (N_3678,N_2734,N_2971);
and U3679 (N_3679,N_2340,N_2044);
or U3680 (N_3680,N_2739,N_2135);
xor U3681 (N_3681,N_2467,N_2913);
and U3682 (N_3682,N_2962,N_2450);
nand U3683 (N_3683,N_2815,N_2135);
nor U3684 (N_3684,N_2064,N_2428);
xor U3685 (N_3685,N_2661,N_2897);
or U3686 (N_3686,N_2938,N_2046);
xnor U3687 (N_3687,N_2209,N_2156);
nand U3688 (N_3688,N_2215,N_2754);
nor U3689 (N_3689,N_2661,N_2640);
nand U3690 (N_3690,N_2176,N_2588);
or U3691 (N_3691,N_2700,N_2573);
or U3692 (N_3692,N_2556,N_2485);
nand U3693 (N_3693,N_2969,N_2597);
or U3694 (N_3694,N_2429,N_2068);
and U3695 (N_3695,N_2656,N_2041);
nor U3696 (N_3696,N_2008,N_2501);
nand U3697 (N_3697,N_2230,N_2120);
xnor U3698 (N_3698,N_2507,N_2249);
nand U3699 (N_3699,N_2723,N_2943);
nor U3700 (N_3700,N_2364,N_2867);
and U3701 (N_3701,N_2392,N_2729);
and U3702 (N_3702,N_2133,N_2355);
nor U3703 (N_3703,N_2401,N_2762);
nor U3704 (N_3704,N_2447,N_2616);
or U3705 (N_3705,N_2656,N_2086);
nor U3706 (N_3706,N_2330,N_2037);
nand U3707 (N_3707,N_2633,N_2689);
or U3708 (N_3708,N_2720,N_2071);
nand U3709 (N_3709,N_2553,N_2676);
nand U3710 (N_3710,N_2152,N_2336);
or U3711 (N_3711,N_2632,N_2837);
xor U3712 (N_3712,N_2386,N_2760);
nor U3713 (N_3713,N_2533,N_2947);
and U3714 (N_3714,N_2975,N_2061);
xnor U3715 (N_3715,N_2617,N_2787);
and U3716 (N_3716,N_2694,N_2705);
and U3717 (N_3717,N_2735,N_2425);
xnor U3718 (N_3718,N_2657,N_2101);
and U3719 (N_3719,N_2978,N_2107);
and U3720 (N_3720,N_2768,N_2616);
xor U3721 (N_3721,N_2414,N_2449);
and U3722 (N_3722,N_2061,N_2004);
or U3723 (N_3723,N_2879,N_2070);
nor U3724 (N_3724,N_2780,N_2328);
nor U3725 (N_3725,N_2501,N_2835);
nand U3726 (N_3726,N_2341,N_2296);
nor U3727 (N_3727,N_2038,N_2125);
xnor U3728 (N_3728,N_2476,N_2901);
nor U3729 (N_3729,N_2437,N_2527);
and U3730 (N_3730,N_2142,N_2677);
and U3731 (N_3731,N_2320,N_2034);
nor U3732 (N_3732,N_2083,N_2227);
nor U3733 (N_3733,N_2524,N_2513);
or U3734 (N_3734,N_2501,N_2648);
xor U3735 (N_3735,N_2576,N_2199);
nand U3736 (N_3736,N_2945,N_2086);
nor U3737 (N_3737,N_2963,N_2380);
or U3738 (N_3738,N_2030,N_2344);
or U3739 (N_3739,N_2378,N_2633);
or U3740 (N_3740,N_2043,N_2760);
xnor U3741 (N_3741,N_2618,N_2109);
nand U3742 (N_3742,N_2837,N_2067);
nand U3743 (N_3743,N_2367,N_2990);
xor U3744 (N_3744,N_2030,N_2131);
xor U3745 (N_3745,N_2172,N_2791);
nor U3746 (N_3746,N_2018,N_2103);
and U3747 (N_3747,N_2559,N_2601);
and U3748 (N_3748,N_2456,N_2243);
nand U3749 (N_3749,N_2345,N_2704);
nor U3750 (N_3750,N_2708,N_2407);
nor U3751 (N_3751,N_2515,N_2762);
and U3752 (N_3752,N_2163,N_2899);
xnor U3753 (N_3753,N_2909,N_2345);
nand U3754 (N_3754,N_2034,N_2860);
xnor U3755 (N_3755,N_2407,N_2279);
or U3756 (N_3756,N_2280,N_2210);
nor U3757 (N_3757,N_2340,N_2326);
or U3758 (N_3758,N_2470,N_2150);
xnor U3759 (N_3759,N_2927,N_2520);
nand U3760 (N_3760,N_2105,N_2374);
xor U3761 (N_3761,N_2759,N_2326);
nand U3762 (N_3762,N_2377,N_2003);
nor U3763 (N_3763,N_2650,N_2325);
xor U3764 (N_3764,N_2675,N_2371);
or U3765 (N_3765,N_2707,N_2865);
nand U3766 (N_3766,N_2942,N_2860);
and U3767 (N_3767,N_2858,N_2397);
and U3768 (N_3768,N_2576,N_2009);
and U3769 (N_3769,N_2628,N_2239);
xor U3770 (N_3770,N_2985,N_2576);
nor U3771 (N_3771,N_2750,N_2807);
xnor U3772 (N_3772,N_2007,N_2066);
and U3773 (N_3773,N_2475,N_2696);
nand U3774 (N_3774,N_2758,N_2173);
xor U3775 (N_3775,N_2788,N_2854);
and U3776 (N_3776,N_2286,N_2646);
or U3777 (N_3777,N_2865,N_2445);
xor U3778 (N_3778,N_2303,N_2500);
and U3779 (N_3779,N_2864,N_2832);
or U3780 (N_3780,N_2156,N_2612);
xnor U3781 (N_3781,N_2658,N_2942);
or U3782 (N_3782,N_2987,N_2057);
xnor U3783 (N_3783,N_2199,N_2475);
or U3784 (N_3784,N_2415,N_2933);
nor U3785 (N_3785,N_2803,N_2804);
nor U3786 (N_3786,N_2232,N_2633);
nand U3787 (N_3787,N_2465,N_2114);
xor U3788 (N_3788,N_2905,N_2632);
nor U3789 (N_3789,N_2040,N_2089);
nor U3790 (N_3790,N_2240,N_2924);
xnor U3791 (N_3791,N_2623,N_2714);
xnor U3792 (N_3792,N_2804,N_2211);
and U3793 (N_3793,N_2441,N_2053);
nor U3794 (N_3794,N_2531,N_2631);
and U3795 (N_3795,N_2543,N_2927);
nor U3796 (N_3796,N_2718,N_2232);
nor U3797 (N_3797,N_2016,N_2037);
xnor U3798 (N_3798,N_2425,N_2333);
or U3799 (N_3799,N_2975,N_2319);
or U3800 (N_3800,N_2461,N_2337);
nand U3801 (N_3801,N_2062,N_2535);
nand U3802 (N_3802,N_2039,N_2816);
nor U3803 (N_3803,N_2354,N_2595);
and U3804 (N_3804,N_2228,N_2355);
and U3805 (N_3805,N_2472,N_2396);
and U3806 (N_3806,N_2571,N_2748);
and U3807 (N_3807,N_2857,N_2786);
xnor U3808 (N_3808,N_2173,N_2637);
and U3809 (N_3809,N_2944,N_2878);
and U3810 (N_3810,N_2741,N_2116);
or U3811 (N_3811,N_2899,N_2130);
and U3812 (N_3812,N_2216,N_2123);
and U3813 (N_3813,N_2905,N_2612);
and U3814 (N_3814,N_2421,N_2881);
and U3815 (N_3815,N_2736,N_2353);
and U3816 (N_3816,N_2494,N_2285);
nor U3817 (N_3817,N_2628,N_2245);
xnor U3818 (N_3818,N_2795,N_2063);
nor U3819 (N_3819,N_2884,N_2294);
or U3820 (N_3820,N_2008,N_2451);
or U3821 (N_3821,N_2534,N_2638);
and U3822 (N_3822,N_2530,N_2861);
and U3823 (N_3823,N_2164,N_2304);
nor U3824 (N_3824,N_2054,N_2095);
nand U3825 (N_3825,N_2025,N_2312);
or U3826 (N_3826,N_2556,N_2971);
or U3827 (N_3827,N_2395,N_2770);
xnor U3828 (N_3828,N_2878,N_2909);
and U3829 (N_3829,N_2215,N_2048);
nand U3830 (N_3830,N_2659,N_2731);
nor U3831 (N_3831,N_2730,N_2294);
or U3832 (N_3832,N_2170,N_2359);
and U3833 (N_3833,N_2185,N_2021);
nand U3834 (N_3834,N_2615,N_2118);
nand U3835 (N_3835,N_2377,N_2750);
or U3836 (N_3836,N_2511,N_2604);
nand U3837 (N_3837,N_2590,N_2406);
or U3838 (N_3838,N_2429,N_2989);
nor U3839 (N_3839,N_2343,N_2268);
and U3840 (N_3840,N_2561,N_2549);
and U3841 (N_3841,N_2841,N_2973);
and U3842 (N_3842,N_2862,N_2872);
or U3843 (N_3843,N_2053,N_2415);
or U3844 (N_3844,N_2015,N_2478);
and U3845 (N_3845,N_2254,N_2412);
nor U3846 (N_3846,N_2776,N_2511);
and U3847 (N_3847,N_2421,N_2556);
xor U3848 (N_3848,N_2122,N_2563);
xnor U3849 (N_3849,N_2573,N_2067);
or U3850 (N_3850,N_2268,N_2190);
and U3851 (N_3851,N_2173,N_2610);
nor U3852 (N_3852,N_2091,N_2757);
nor U3853 (N_3853,N_2170,N_2234);
nand U3854 (N_3854,N_2028,N_2490);
nand U3855 (N_3855,N_2720,N_2666);
nand U3856 (N_3856,N_2807,N_2552);
and U3857 (N_3857,N_2733,N_2772);
nand U3858 (N_3858,N_2881,N_2197);
or U3859 (N_3859,N_2999,N_2997);
or U3860 (N_3860,N_2629,N_2646);
nand U3861 (N_3861,N_2690,N_2116);
and U3862 (N_3862,N_2318,N_2842);
nand U3863 (N_3863,N_2932,N_2533);
xor U3864 (N_3864,N_2637,N_2959);
or U3865 (N_3865,N_2743,N_2720);
or U3866 (N_3866,N_2247,N_2870);
or U3867 (N_3867,N_2980,N_2918);
xnor U3868 (N_3868,N_2344,N_2730);
xnor U3869 (N_3869,N_2787,N_2682);
or U3870 (N_3870,N_2678,N_2972);
and U3871 (N_3871,N_2584,N_2354);
nor U3872 (N_3872,N_2283,N_2250);
nor U3873 (N_3873,N_2213,N_2431);
or U3874 (N_3874,N_2164,N_2488);
xor U3875 (N_3875,N_2773,N_2305);
and U3876 (N_3876,N_2384,N_2093);
and U3877 (N_3877,N_2868,N_2531);
nor U3878 (N_3878,N_2224,N_2792);
nor U3879 (N_3879,N_2606,N_2285);
and U3880 (N_3880,N_2167,N_2210);
and U3881 (N_3881,N_2041,N_2951);
nor U3882 (N_3882,N_2254,N_2045);
xor U3883 (N_3883,N_2378,N_2987);
and U3884 (N_3884,N_2237,N_2403);
nor U3885 (N_3885,N_2148,N_2875);
xnor U3886 (N_3886,N_2666,N_2388);
nand U3887 (N_3887,N_2209,N_2862);
xor U3888 (N_3888,N_2384,N_2131);
nor U3889 (N_3889,N_2036,N_2552);
nor U3890 (N_3890,N_2706,N_2118);
and U3891 (N_3891,N_2851,N_2049);
xor U3892 (N_3892,N_2003,N_2443);
xnor U3893 (N_3893,N_2999,N_2048);
nor U3894 (N_3894,N_2774,N_2612);
and U3895 (N_3895,N_2446,N_2011);
nand U3896 (N_3896,N_2985,N_2684);
nor U3897 (N_3897,N_2185,N_2539);
xnor U3898 (N_3898,N_2701,N_2005);
and U3899 (N_3899,N_2924,N_2651);
xnor U3900 (N_3900,N_2830,N_2362);
or U3901 (N_3901,N_2340,N_2597);
or U3902 (N_3902,N_2265,N_2236);
xnor U3903 (N_3903,N_2075,N_2956);
or U3904 (N_3904,N_2321,N_2243);
nand U3905 (N_3905,N_2105,N_2775);
nand U3906 (N_3906,N_2124,N_2235);
or U3907 (N_3907,N_2520,N_2114);
nand U3908 (N_3908,N_2116,N_2308);
nand U3909 (N_3909,N_2467,N_2097);
and U3910 (N_3910,N_2241,N_2832);
and U3911 (N_3911,N_2517,N_2978);
xor U3912 (N_3912,N_2792,N_2042);
xor U3913 (N_3913,N_2665,N_2415);
xnor U3914 (N_3914,N_2505,N_2224);
or U3915 (N_3915,N_2233,N_2683);
or U3916 (N_3916,N_2721,N_2269);
or U3917 (N_3917,N_2293,N_2166);
and U3918 (N_3918,N_2596,N_2271);
and U3919 (N_3919,N_2572,N_2583);
nor U3920 (N_3920,N_2026,N_2944);
nand U3921 (N_3921,N_2562,N_2565);
xnor U3922 (N_3922,N_2398,N_2949);
and U3923 (N_3923,N_2207,N_2650);
nor U3924 (N_3924,N_2395,N_2830);
nand U3925 (N_3925,N_2326,N_2852);
nor U3926 (N_3926,N_2672,N_2694);
and U3927 (N_3927,N_2765,N_2888);
nor U3928 (N_3928,N_2139,N_2655);
nand U3929 (N_3929,N_2083,N_2358);
nor U3930 (N_3930,N_2203,N_2789);
nor U3931 (N_3931,N_2304,N_2558);
xor U3932 (N_3932,N_2292,N_2763);
nand U3933 (N_3933,N_2206,N_2115);
or U3934 (N_3934,N_2538,N_2073);
or U3935 (N_3935,N_2019,N_2897);
nand U3936 (N_3936,N_2517,N_2421);
or U3937 (N_3937,N_2715,N_2718);
nand U3938 (N_3938,N_2488,N_2493);
and U3939 (N_3939,N_2756,N_2584);
and U3940 (N_3940,N_2491,N_2227);
or U3941 (N_3941,N_2302,N_2433);
nor U3942 (N_3942,N_2751,N_2814);
nor U3943 (N_3943,N_2809,N_2730);
xor U3944 (N_3944,N_2727,N_2843);
nor U3945 (N_3945,N_2730,N_2506);
nand U3946 (N_3946,N_2650,N_2871);
and U3947 (N_3947,N_2635,N_2690);
xor U3948 (N_3948,N_2744,N_2935);
nand U3949 (N_3949,N_2277,N_2456);
xnor U3950 (N_3950,N_2935,N_2391);
xnor U3951 (N_3951,N_2277,N_2664);
nor U3952 (N_3952,N_2160,N_2337);
or U3953 (N_3953,N_2314,N_2762);
or U3954 (N_3954,N_2683,N_2601);
and U3955 (N_3955,N_2572,N_2524);
or U3956 (N_3956,N_2448,N_2665);
or U3957 (N_3957,N_2266,N_2007);
xnor U3958 (N_3958,N_2626,N_2968);
and U3959 (N_3959,N_2665,N_2427);
nand U3960 (N_3960,N_2696,N_2340);
and U3961 (N_3961,N_2570,N_2659);
nand U3962 (N_3962,N_2728,N_2746);
nand U3963 (N_3963,N_2706,N_2212);
or U3964 (N_3964,N_2881,N_2406);
or U3965 (N_3965,N_2873,N_2262);
nand U3966 (N_3966,N_2771,N_2599);
nand U3967 (N_3967,N_2781,N_2409);
nand U3968 (N_3968,N_2134,N_2540);
nand U3969 (N_3969,N_2518,N_2110);
nand U3970 (N_3970,N_2657,N_2131);
nand U3971 (N_3971,N_2488,N_2755);
or U3972 (N_3972,N_2067,N_2562);
nor U3973 (N_3973,N_2440,N_2862);
nand U3974 (N_3974,N_2671,N_2050);
xor U3975 (N_3975,N_2065,N_2248);
nor U3976 (N_3976,N_2148,N_2656);
or U3977 (N_3977,N_2721,N_2506);
nand U3978 (N_3978,N_2858,N_2704);
xnor U3979 (N_3979,N_2991,N_2639);
and U3980 (N_3980,N_2056,N_2142);
and U3981 (N_3981,N_2395,N_2784);
and U3982 (N_3982,N_2114,N_2210);
xnor U3983 (N_3983,N_2707,N_2705);
xnor U3984 (N_3984,N_2748,N_2009);
xor U3985 (N_3985,N_2089,N_2379);
or U3986 (N_3986,N_2534,N_2000);
xnor U3987 (N_3987,N_2850,N_2102);
and U3988 (N_3988,N_2417,N_2716);
nor U3989 (N_3989,N_2501,N_2498);
nor U3990 (N_3990,N_2003,N_2273);
nand U3991 (N_3991,N_2576,N_2395);
nor U3992 (N_3992,N_2260,N_2593);
and U3993 (N_3993,N_2527,N_2602);
and U3994 (N_3994,N_2322,N_2342);
nor U3995 (N_3995,N_2382,N_2948);
xor U3996 (N_3996,N_2246,N_2905);
xnor U3997 (N_3997,N_2261,N_2053);
and U3998 (N_3998,N_2766,N_2679);
nand U3999 (N_3999,N_2925,N_2439);
nand U4000 (N_4000,N_3127,N_3000);
nor U4001 (N_4001,N_3905,N_3172);
nand U4002 (N_4002,N_3886,N_3403);
nor U4003 (N_4003,N_3453,N_3089);
nor U4004 (N_4004,N_3246,N_3238);
nor U4005 (N_4005,N_3558,N_3445);
nor U4006 (N_4006,N_3166,N_3845);
and U4007 (N_4007,N_3601,N_3695);
or U4008 (N_4008,N_3686,N_3224);
nand U4009 (N_4009,N_3211,N_3998);
or U4010 (N_4010,N_3449,N_3337);
and U4011 (N_4011,N_3621,N_3259);
and U4012 (N_4012,N_3634,N_3201);
nand U4013 (N_4013,N_3703,N_3240);
nor U4014 (N_4014,N_3554,N_3305);
xor U4015 (N_4015,N_3606,N_3414);
and U4016 (N_4016,N_3884,N_3515);
and U4017 (N_4017,N_3043,N_3516);
or U4018 (N_4018,N_3815,N_3080);
xnor U4019 (N_4019,N_3039,N_3219);
and U4020 (N_4020,N_3985,N_3233);
nand U4021 (N_4021,N_3207,N_3848);
or U4022 (N_4022,N_3145,N_3605);
nand U4023 (N_4023,N_3744,N_3077);
nand U4024 (N_4024,N_3252,N_3951);
or U4025 (N_4025,N_3781,N_3035);
and U4026 (N_4026,N_3796,N_3106);
xnor U4027 (N_4027,N_3272,N_3274);
or U4028 (N_4028,N_3447,N_3939);
xnor U4029 (N_4029,N_3673,N_3231);
xor U4030 (N_4030,N_3922,N_3596);
or U4031 (N_4031,N_3283,N_3868);
and U4032 (N_4032,N_3338,N_3756);
or U4033 (N_4033,N_3739,N_3003);
or U4034 (N_4034,N_3661,N_3121);
and U4035 (N_4035,N_3674,N_3830);
or U4036 (N_4036,N_3365,N_3698);
xnor U4037 (N_4037,N_3766,N_3617);
nand U4038 (N_4038,N_3431,N_3385);
nor U4039 (N_4039,N_3426,N_3742);
or U4040 (N_4040,N_3086,N_3390);
and U4041 (N_4041,N_3051,N_3986);
xor U4042 (N_4042,N_3457,N_3740);
nand U4043 (N_4043,N_3297,N_3943);
and U4044 (N_4044,N_3346,N_3169);
xor U4045 (N_4045,N_3441,N_3876);
nor U4046 (N_4046,N_3637,N_3239);
and U4047 (N_4047,N_3576,N_3570);
xnor U4048 (N_4048,N_3652,N_3225);
or U4049 (N_4049,N_3456,N_3693);
or U4050 (N_4050,N_3021,N_3977);
or U4051 (N_4051,N_3679,N_3372);
xnor U4052 (N_4052,N_3728,N_3310);
or U4053 (N_4053,N_3108,N_3509);
xnor U4054 (N_4054,N_3993,N_3340);
nor U4055 (N_4055,N_3521,N_3389);
or U4056 (N_4056,N_3140,N_3858);
nor U4057 (N_4057,N_3263,N_3490);
nor U4058 (N_4058,N_3037,N_3780);
nor U4059 (N_4059,N_3997,N_3746);
nor U4060 (N_4060,N_3005,N_3591);
nor U4061 (N_4061,N_3782,N_3170);
nand U4062 (N_4062,N_3134,N_3292);
nand U4063 (N_4063,N_3113,N_3123);
nor U4064 (N_4064,N_3324,N_3339);
nand U4065 (N_4065,N_3421,N_3991);
xor U4066 (N_4066,N_3460,N_3241);
nand U4067 (N_4067,N_3598,N_3212);
or U4068 (N_4068,N_3408,N_3306);
nor U4069 (N_4069,N_3869,N_3588);
nor U4070 (N_4070,N_3811,N_3709);
xnor U4071 (N_4071,N_3304,N_3342);
and U4072 (N_4072,N_3485,N_3178);
xor U4073 (N_4073,N_3633,N_3446);
nand U4074 (N_4074,N_3575,N_3741);
xor U4075 (N_4075,N_3569,N_3094);
nand U4076 (N_4076,N_3941,N_3293);
xor U4077 (N_4077,N_3085,N_3931);
and U4078 (N_4078,N_3062,N_3948);
xnor U4079 (N_4079,N_3850,N_3102);
xor U4080 (N_4080,N_3187,N_3434);
and U4081 (N_4081,N_3567,N_3197);
nand U4082 (N_4082,N_3041,N_3415);
nor U4083 (N_4083,N_3139,N_3291);
nand U4084 (N_4084,N_3579,N_3797);
nand U4085 (N_4085,N_3683,N_3608);
xnor U4086 (N_4086,N_3377,N_3029);
nand U4087 (N_4087,N_3896,N_3440);
xor U4088 (N_4088,N_3120,N_3573);
and U4089 (N_4089,N_3607,N_3542);
or U4090 (N_4090,N_3995,N_3894);
and U4091 (N_4091,N_3510,N_3543);
nand U4092 (N_4092,N_3836,N_3935);
xor U4093 (N_4093,N_3594,N_3158);
nand U4094 (N_4094,N_3787,N_3639);
and U4095 (N_4095,N_3331,N_3568);
nand U4096 (N_4096,N_3507,N_3032);
nor U4097 (N_4097,N_3899,N_3553);
nand U4098 (N_4098,N_3915,N_3027);
xnor U4099 (N_4099,N_3437,N_3433);
nand U4100 (N_4100,N_3128,N_3196);
nand U4101 (N_4101,N_3467,N_3511);
xnor U4102 (N_4102,N_3857,N_3821);
or U4103 (N_4103,N_3011,N_3073);
xor U4104 (N_4104,N_3273,N_3056);
and U4105 (N_4105,N_3798,N_3046);
nand U4106 (N_4106,N_3940,N_3171);
nand U4107 (N_4107,N_3435,N_3716);
and U4108 (N_4108,N_3154,N_3028);
nand U4109 (N_4109,N_3471,N_3363);
nor U4110 (N_4110,N_3767,N_3982);
and U4111 (N_4111,N_3557,N_3720);
xor U4112 (N_4112,N_3959,N_3413);
nor U4113 (N_4113,N_3548,N_3450);
or U4114 (N_4114,N_3812,N_3373);
and U4115 (N_4115,N_3146,N_3612);
xnor U4116 (N_4116,N_3919,N_3049);
or U4117 (N_4117,N_3451,N_3153);
nand U4118 (N_4118,N_3105,N_3249);
or U4119 (N_4119,N_3026,N_3148);
nor U4120 (N_4120,N_3384,N_3820);
or U4121 (N_4121,N_3984,N_3700);
or U4122 (N_4122,N_3934,N_3795);
or U4123 (N_4123,N_3161,N_3816);
xnor U4124 (N_4124,N_3779,N_3945);
nor U4125 (N_4125,N_3929,N_3132);
and U4126 (N_4126,N_3595,N_3719);
nor U4127 (N_4127,N_3404,N_3459);
nor U4128 (N_4128,N_3793,N_3859);
xnor U4129 (N_4129,N_3743,N_3523);
nor U4130 (N_4130,N_3974,N_3937);
or U4131 (N_4131,N_3824,N_3671);
nor U4132 (N_4132,N_3953,N_3495);
nand U4133 (N_4133,N_3186,N_3764);
nand U4134 (N_4134,N_3354,N_3770);
or U4135 (N_4135,N_3417,N_3602);
and U4136 (N_4136,N_3429,N_3109);
nand U4137 (N_4137,N_3494,N_3090);
or U4138 (N_4138,N_3358,N_3823);
or U4139 (N_4139,N_3177,N_3466);
and U4140 (N_4140,N_3017,N_3091);
or U4141 (N_4141,N_3060,N_3866);
nor U4142 (N_4142,N_3498,N_3670);
and U4143 (N_4143,N_3651,N_3057);
or U4144 (N_4144,N_3957,N_3748);
nand U4145 (N_4145,N_3111,N_3278);
and U4146 (N_4146,N_3001,N_3343);
or U4147 (N_4147,N_3375,N_3650);
and U4148 (N_4148,N_3654,N_3009);
xor U4149 (N_4149,N_3980,N_3462);
nor U4150 (N_4150,N_3938,N_3103);
or U4151 (N_4151,N_3101,N_3374);
and U4152 (N_4152,N_3334,N_3712);
xnor U4153 (N_4153,N_3152,N_3402);
nor U4154 (N_4154,N_3505,N_3512);
xor U4155 (N_4155,N_3890,N_3540);
or U4156 (N_4156,N_3662,N_3299);
and U4157 (N_4157,N_3463,N_3862);
and U4158 (N_4158,N_3844,N_3150);
nand U4159 (N_4159,N_3735,N_3578);
and U4160 (N_4160,N_3107,N_3873);
or U4161 (N_4161,N_3618,N_3174);
xor U4162 (N_4162,N_3175,N_3646);
nand U4163 (N_4163,N_3678,N_3410);
xnor U4164 (N_4164,N_3914,N_3318);
or U4165 (N_4165,N_3465,N_3100);
nand U4166 (N_4166,N_3478,N_3015);
and U4167 (N_4167,N_3666,N_3788);
nor U4168 (N_4168,N_3183,N_3371);
xor U4169 (N_4169,N_3789,N_3800);
nor U4170 (N_4170,N_3794,N_3849);
and U4171 (N_4171,N_3279,N_3475);
nand U4172 (N_4172,N_3059,N_3874);
nor U4173 (N_4173,N_3379,N_3627);
xnor U4174 (N_4174,N_3226,N_3296);
nand U4175 (N_4175,N_3638,N_3260);
or U4176 (N_4176,N_3353,N_3040);
nor U4177 (N_4177,N_3427,N_3772);
and U4178 (N_4178,N_3572,N_3600);
and U4179 (N_4179,N_3277,N_3968);
nand U4180 (N_4180,N_3909,N_3069);
nor U4181 (N_4181,N_3286,N_3738);
nor U4182 (N_4182,N_3988,N_3355);
nor U4183 (N_4183,N_3645,N_3122);
nor U4184 (N_4184,N_3078,N_3571);
nand U4185 (N_4185,N_3904,N_3492);
nand U4186 (N_4186,N_3526,N_3084);
xnor U4187 (N_4187,N_3685,N_3513);
xor U4188 (N_4188,N_3883,N_3269);
nor U4189 (N_4189,N_3368,N_3133);
nor U4190 (N_4190,N_3087,N_3870);
or U4191 (N_4191,N_3393,N_3932);
and U4192 (N_4192,N_3416,N_3762);
nand U4193 (N_4193,N_3903,N_3577);
or U4194 (N_4194,N_3411,N_3332);
xor U4195 (N_4195,N_3229,N_3765);
or U4196 (N_4196,N_3658,N_3834);
nand U4197 (N_4197,N_3706,N_3865);
or U4198 (N_4198,N_3315,N_3692);
nand U4199 (N_4199,N_3665,N_3649);
xor U4200 (N_4200,N_3232,N_3036);
or U4201 (N_4201,N_3684,N_3852);
and U4202 (N_4202,N_3129,N_3344);
or U4203 (N_4203,N_3616,N_3659);
and U4204 (N_4204,N_3395,N_3587);
and U4205 (N_4205,N_3841,N_3137);
nor U4206 (N_4206,N_3159,N_3614);
and U4207 (N_4207,N_3061,N_3644);
and U4208 (N_4208,N_3267,N_3620);
nor U4209 (N_4209,N_3290,N_3911);
xor U4210 (N_4210,N_3536,N_3847);
nand U4211 (N_4211,N_3992,N_3892);
and U4212 (N_4212,N_3973,N_3407);
or U4213 (N_4213,N_3777,N_3387);
and U4214 (N_4214,N_3042,N_3615);
or U4215 (N_4215,N_3258,N_3335);
and U4216 (N_4216,N_3330,N_3047);
and U4217 (N_4217,N_3244,N_3484);
or U4218 (N_4218,N_3877,N_3966);
and U4219 (N_4219,N_3609,N_3535);
nand U4220 (N_4220,N_3173,N_3967);
xnor U4221 (N_4221,N_3574,N_3033);
xnor U4222 (N_4222,N_3981,N_3603);
or U4223 (N_4223,N_3625,N_3264);
xnor U4224 (N_4224,N_3491,N_3923);
or U4225 (N_4225,N_3710,N_3584);
or U4226 (N_4226,N_3217,N_3308);
nor U4227 (N_4227,N_3209,N_3970);
or U4228 (N_4228,N_3301,N_3480);
nand U4229 (N_4229,N_3829,N_3176);
and U4230 (N_4230,N_3030,N_3486);
and U4231 (N_4231,N_3112,N_3696);
or U4232 (N_4232,N_3619,N_3546);
xnor U4233 (N_4233,N_3020,N_3541);
and U4234 (N_4234,N_3382,N_3717);
nor U4235 (N_4235,N_3640,N_3641);
xor U4236 (N_4236,N_3708,N_3452);
nor U4237 (N_4237,N_3302,N_3157);
and U4238 (N_4238,N_3955,N_3882);
and U4239 (N_4239,N_3819,N_3549);
nand U4240 (N_4240,N_3432,N_3851);
nor U4241 (N_4241,N_3499,N_3255);
xor U4242 (N_4242,N_3702,N_3326);
xnor U4243 (N_4243,N_3628,N_3223);
nor U4244 (N_4244,N_3200,N_3400);
nor U4245 (N_4245,N_3281,N_3097);
nor U4246 (N_4246,N_3329,N_3804);
nand U4247 (N_4247,N_3555,N_3624);
xor U4248 (N_4248,N_3726,N_3864);
or U4249 (N_4249,N_3531,N_3235);
nand U4250 (N_4250,N_3520,N_3551);
xnor U4251 (N_4251,N_3333,N_3018);
nor U4252 (N_4252,N_3220,N_3533);
and U4253 (N_4253,N_3908,N_3420);
nor U4254 (N_4254,N_3597,N_3253);
and U4255 (N_4255,N_3162,N_3774);
nor U4256 (N_4256,N_3814,N_3856);
and U4257 (N_4257,N_3356,N_3715);
and U4258 (N_4258,N_3117,N_3733);
nor U4259 (N_4259,N_3885,N_3916);
or U4260 (N_4260,N_3629,N_3002);
nor U4261 (N_4261,N_3773,N_3527);
nor U4262 (N_4262,N_3803,N_3325);
nor U4263 (N_4263,N_3544,N_3401);
nor U4264 (N_4264,N_3663,N_3736);
nor U4265 (N_4265,N_3843,N_3730);
xor U4266 (N_4266,N_3156,N_3359);
nand U4267 (N_4267,N_3810,N_3270);
and U4268 (N_4268,N_3257,N_3063);
or U4269 (N_4269,N_3960,N_3718);
or U4270 (N_4270,N_3163,N_3345);
xnor U4271 (N_4271,N_3230,N_3054);
nand U4272 (N_4272,N_3783,N_3454);
xnor U4273 (N_4273,N_3635,N_3282);
xor U4274 (N_4274,N_3838,N_3376);
xnor U4275 (N_4275,N_3759,N_3522);
nand U4276 (N_4276,N_3048,N_3912);
and U4277 (N_4277,N_3469,N_3473);
nand U4278 (N_4278,N_3023,N_3118);
nand U4279 (N_4279,N_3626,N_3083);
or U4280 (N_4280,N_3755,N_3822);
and U4281 (N_4281,N_3221,N_3058);
nand U4282 (N_4282,N_3754,N_3688);
nand U4283 (N_4283,N_3502,N_3479);
nor U4284 (N_4284,N_3381,N_3248);
xor U4285 (N_4285,N_3312,N_3422);
xor U4286 (N_4286,N_3289,N_3236);
xor U4287 (N_4287,N_3461,N_3095);
and U4288 (N_4288,N_3202,N_3802);
nand U4289 (N_4289,N_3562,N_3776);
or U4290 (N_4290,N_3317,N_3439);
and U4291 (N_4291,N_3074,N_3907);
and U4292 (N_4292,N_3623,N_3070);
nor U4293 (N_4293,N_3950,N_3016);
and U4294 (N_4294,N_3891,N_3768);
or U4295 (N_4295,N_3954,N_3831);
xnor U4296 (N_4296,N_3725,N_3604);
nand U4297 (N_4297,N_3983,N_3455);
nor U4298 (N_4298,N_3487,N_3825);
nand U4299 (N_4299,N_3927,N_3593);
nand U4300 (N_4300,N_3581,N_3357);
or U4301 (N_4301,N_3917,N_3989);
and U4302 (N_4302,N_3632,N_3999);
and U4303 (N_4303,N_3947,N_3131);
and U4304 (N_4304,N_3737,N_3251);
nand U4305 (N_4305,N_3871,N_3622);
nand U4306 (N_4306,N_3280,N_3364);
nor U4307 (N_4307,N_3500,N_3067);
or U4308 (N_4308,N_3323,N_3470);
xnor U4309 (N_4309,N_3068,N_3181);
or U4310 (N_4310,N_3321,N_3933);
and U4311 (N_4311,N_3294,N_3946);
and U4312 (N_4312,N_3972,N_3468);
nand U4313 (N_4313,N_3206,N_3750);
nor U4314 (N_4314,N_3517,N_3397);
xnor U4315 (N_4315,N_3930,N_3707);
and U4316 (N_4316,N_3012,N_3504);
nand U4317 (N_4317,N_3889,N_3965);
xnor U4318 (N_4318,N_3918,N_3749);
and U4319 (N_4319,N_3832,N_3563);
and U4320 (N_4320,N_3566,N_3518);
nand U4321 (N_4321,N_3116,N_3093);
xnor U4322 (N_4322,N_3860,N_3184);
nand U4323 (N_4323,N_3295,N_3099);
nand U4324 (N_4324,N_3758,N_3045);
nor U4325 (N_4325,N_3014,N_3271);
nor U4326 (N_4326,N_3556,N_3669);
nor U4327 (N_4327,N_3436,N_3753);
nor U4328 (N_4328,N_3818,N_3066);
nor U4329 (N_4329,N_3921,N_3214);
and U4330 (N_4330,N_3147,N_3472);
nand U4331 (N_4331,N_3428,N_3006);
nand U4332 (N_4332,N_3423,N_3010);
nor U4333 (N_4333,N_3004,N_3705);
nor U4334 (N_4334,N_3360,N_3532);
xor U4335 (N_4335,N_3496,N_3583);
or U4336 (N_4336,N_3243,N_3052);
and U4337 (N_4337,N_3901,N_3963);
nand U4338 (N_4338,N_3443,N_3138);
and U4339 (N_4339,N_3550,N_3867);
nor U4340 (N_4340,N_3007,N_3840);
nand U4341 (N_4341,N_3350,N_3714);
and U4342 (N_4342,N_3198,N_3367);
xor U4343 (N_4343,N_3880,N_3194);
and U4344 (N_4344,N_3846,N_3881);
nand U4345 (N_4345,N_3370,N_3298);
and U4346 (N_4346,N_3668,N_3419);
xnor U4347 (N_4347,N_3261,N_3320);
or U4348 (N_4348,N_3613,N_3114);
and U4349 (N_4349,N_3722,N_3193);
and U4350 (N_4350,N_3971,N_3474);
nand U4351 (N_4351,N_3477,N_3180);
nor U4352 (N_4352,N_3388,N_3547);
or U4353 (N_4353,N_3994,N_3792);
xnor U4354 (N_4354,N_3529,N_3514);
or U4355 (N_4355,N_3893,N_3817);
nand U4356 (N_4356,N_3481,N_3534);
and U4357 (N_4357,N_3254,N_3341);
nor U4358 (N_4358,N_3208,N_3978);
nand U4359 (N_4359,N_3352,N_3394);
or U4360 (N_4360,N_3386,N_3675);
nand U4361 (N_4361,N_3348,N_3697);
nand U4362 (N_4362,N_3655,N_3444);
or U4363 (N_4363,N_3813,N_3242);
nand U4364 (N_4364,N_3322,N_3210);
nand U4365 (N_4365,N_3676,N_3539);
or U4366 (N_4366,N_3050,N_3942);
or U4367 (N_4367,N_3380,N_3961);
nor U4368 (N_4368,N_3694,N_3053);
nor U4369 (N_4369,N_3237,N_3245);
or U4370 (N_4370,N_3537,N_3808);
xnor U4371 (N_4371,N_3672,N_3366);
nor U4372 (N_4372,N_3732,N_3319);
xnor U4373 (N_4373,N_3250,N_3424);
and U4374 (N_4374,N_3936,N_3895);
or U4375 (N_4375,N_3476,N_3731);
or U4376 (N_4376,N_3786,N_3647);
nor U4377 (N_4377,N_3228,N_3227);
and U4378 (N_4378,N_3412,N_3124);
or U4379 (N_4379,N_3975,N_3913);
or U4380 (N_4380,N_3837,N_3826);
or U4381 (N_4381,N_3727,N_3369);
xor U4382 (N_4382,N_3448,N_3530);
and U4383 (N_4383,N_3336,N_3398);
xnor U4384 (N_4384,N_3488,N_3660);
and U4385 (N_4385,N_3098,N_3506);
xor U4386 (N_4386,N_3680,N_3378);
nand U4387 (N_4387,N_3979,N_3524);
nand U4388 (N_4388,N_3144,N_3164);
nor U4389 (N_4389,N_3835,N_3853);
nand U4390 (N_4390,N_3022,N_3580);
nand U4391 (N_4391,N_3642,N_3656);
nor U4392 (N_4392,N_3136,N_3110);
or U4393 (N_4393,N_3809,N_3778);
nor U4394 (N_4394,N_3256,N_3019);
xor U4395 (N_4395,N_3179,N_3976);
nor U4396 (N_4396,N_3215,N_3126);
nand U4397 (N_4397,N_3664,N_3842);
and U4398 (N_4398,N_3752,N_3438);
or U4399 (N_4399,N_3160,N_3760);
nor U4400 (N_4400,N_3590,N_3805);
nor U4401 (N_4401,N_3082,N_3682);
and U4402 (N_4402,N_3631,N_3956);
and U4403 (N_4403,N_3503,N_3216);
xnor U4404 (N_4404,N_3268,N_3285);
xnor U4405 (N_4405,N_3119,N_3205);
xor U4406 (N_4406,N_3801,N_3065);
nor U4407 (N_4407,N_3872,N_3888);
nand U4408 (N_4408,N_3088,N_3025);
nand U4409 (N_4409,N_3863,N_3189);
nand U4410 (N_4410,N_3724,N_3721);
and U4411 (N_4411,N_3704,N_3799);
xnor U4412 (N_4412,N_3687,N_3168);
or U4413 (N_4413,N_3875,N_3636);
or U4414 (N_4414,N_3031,N_3906);
and U4415 (N_4415,N_3926,N_3653);
xnor U4416 (N_4416,N_3962,N_3833);
and U4417 (N_4417,N_3489,N_3072);
nor U4418 (N_4418,N_3564,N_3952);
xor U4419 (N_4419,N_3151,N_3910);
nand U4420 (N_4420,N_3565,N_3141);
xnor U4421 (N_4421,N_3828,N_3545);
or U4422 (N_4422,N_3185,N_3222);
nor U4423 (N_4423,N_3648,N_3044);
nor U4424 (N_4424,N_3076,N_3711);
or U4425 (N_4425,N_3213,N_3839);
or U4426 (N_4426,N_3897,N_3483);
nor U4427 (N_4427,N_3898,N_3677);
nand U4428 (N_4428,N_3347,N_3288);
nand U4429 (N_4429,N_3482,N_3008);
or U4430 (N_4430,N_3525,N_3855);
and U4431 (N_4431,N_3405,N_3024);
or U4432 (N_4432,N_3155,N_3199);
nor U4433 (N_4433,N_3757,N_3130);
nand U4434 (N_4434,N_3262,N_3311);
nor U4435 (N_4435,N_3309,N_3092);
and U4436 (N_4436,N_3081,N_3561);
nor U4437 (N_4437,N_3807,N_3806);
nor U4438 (N_4438,N_3191,N_3790);
or U4439 (N_4439,N_3681,N_3508);
or U4440 (N_4440,N_3643,N_3079);
and U4441 (N_4441,N_3610,N_3391);
and U4442 (N_4442,N_3300,N_3861);
and U4443 (N_4443,N_3854,N_3075);
or U4444 (N_4444,N_3188,N_3038);
xor U4445 (N_4445,N_3538,N_3878);
xor U4446 (N_4446,N_3589,N_3713);
and U4447 (N_4447,N_3418,N_3497);
or U4448 (N_4448,N_3701,N_3275);
nand U4449 (N_4449,N_3314,N_3396);
xnor U4450 (N_4450,N_3071,N_3192);
or U4451 (N_4451,N_3519,N_3691);
nor U4452 (N_4452,N_3990,N_3969);
nand U4453 (N_4453,N_3723,N_3925);
xor U4454 (N_4454,N_3392,N_3287);
xor U4455 (N_4455,N_3442,N_3464);
nor U4456 (N_4456,N_3265,N_3409);
and U4457 (N_4457,N_3689,N_3747);
xor U4458 (N_4458,N_3690,N_3055);
or U4459 (N_4459,N_3064,N_3611);
or U4460 (N_4460,N_3734,N_3552);
xnor U4461 (N_4461,N_3328,N_3182);
or U4462 (N_4462,N_3887,N_3430);
nor U4463 (N_4463,N_3924,N_3203);
xnor U4464 (N_4464,N_3351,N_3195);
and U4465 (N_4465,N_3987,N_3582);
or U4466 (N_4466,N_3327,N_3900);
nor U4467 (N_4467,N_3667,N_3425);
or U4468 (N_4468,N_3125,N_3528);
or U4469 (N_4469,N_3218,N_3303);
nand U4470 (N_4470,N_3458,N_3775);
nor U4471 (N_4471,N_3559,N_3096);
nor U4472 (N_4472,N_3399,N_3592);
and U4473 (N_4473,N_3266,N_3585);
nor U4474 (N_4474,N_3958,N_3729);
nand U4475 (N_4475,N_3104,N_3165);
nor U4476 (N_4476,N_3284,N_3190);
nand U4477 (N_4477,N_3313,N_3204);
nor U4478 (N_4478,N_3234,N_3383);
nor U4479 (N_4479,N_3920,N_3362);
nor U4480 (N_4480,N_3143,N_3879);
nor U4481 (N_4481,N_3167,N_3247);
and U4482 (N_4482,N_3784,N_3630);
and U4483 (N_4483,N_3034,N_3785);
and U4484 (N_4484,N_3827,N_3996);
and U4485 (N_4485,N_3599,N_3769);
xor U4486 (N_4486,N_3902,N_3501);
nand U4487 (N_4487,N_3771,N_3751);
and U4488 (N_4488,N_3949,N_3149);
xnor U4489 (N_4489,N_3560,N_3349);
nand U4490 (N_4490,N_3493,N_3791);
xor U4491 (N_4491,N_3115,N_3361);
nand U4492 (N_4492,N_3944,N_3013);
nor U4493 (N_4493,N_3316,N_3142);
nand U4494 (N_4494,N_3586,N_3699);
nand U4495 (N_4495,N_3657,N_3135);
nor U4496 (N_4496,N_3307,N_3763);
xor U4497 (N_4497,N_3761,N_3745);
nand U4498 (N_4498,N_3964,N_3928);
xor U4499 (N_4499,N_3406,N_3276);
nor U4500 (N_4500,N_3381,N_3688);
nor U4501 (N_4501,N_3469,N_3446);
or U4502 (N_4502,N_3564,N_3004);
nand U4503 (N_4503,N_3315,N_3533);
nand U4504 (N_4504,N_3617,N_3410);
nand U4505 (N_4505,N_3047,N_3269);
and U4506 (N_4506,N_3159,N_3245);
and U4507 (N_4507,N_3488,N_3826);
or U4508 (N_4508,N_3047,N_3310);
xnor U4509 (N_4509,N_3451,N_3434);
or U4510 (N_4510,N_3368,N_3839);
or U4511 (N_4511,N_3444,N_3692);
and U4512 (N_4512,N_3733,N_3748);
and U4513 (N_4513,N_3520,N_3120);
and U4514 (N_4514,N_3716,N_3338);
xnor U4515 (N_4515,N_3840,N_3635);
nor U4516 (N_4516,N_3067,N_3591);
xnor U4517 (N_4517,N_3404,N_3331);
nand U4518 (N_4518,N_3950,N_3174);
and U4519 (N_4519,N_3513,N_3408);
and U4520 (N_4520,N_3353,N_3684);
nor U4521 (N_4521,N_3215,N_3842);
or U4522 (N_4522,N_3484,N_3175);
nand U4523 (N_4523,N_3630,N_3418);
and U4524 (N_4524,N_3394,N_3557);
or U4525 (N_4525,N_3882,N_3208);
or U4526 (N_4526,N_3513,N_3352);
nand U4527 (N_4527,N_3449,N_3871);
and U4528 (N_4528,N_3566,N_3801);
or U4529 (N_4529,N_3434,N_3306);
nor U4530 (N_4530,N_3323,N_3381);
and U4531 (N_4531,N_3542,N_3437);
and U4532 (N_4532,N_3734,N_3987);
nor U4533 (N_4533,N_3371,N_3562);
and U4534 (N_4534,N_3072,N_3321);
nand U4535 (N_4535,N_3243,N_3897);
and U4536 (N_4536,N_3630,N_3668);
or U4537 (N_4537,N_3576,N_3223);
and U4538 (N_4538,N_3472,N_3687);
xor U4539 (N_4539,N_3630,N_3605);
xor U4540 (N_4540,N_3905,N_3590);
nand U4541 (N_4541,N_3005,N_3960);
and U4542 (N_4542,N_3429,N_3655);
and U4543 (N_4543,N_3615,N_3028);
nor U4544 (N_4544,N_3109,N_3092);
nand U4545 (N_4545,N_3694,N_3582);
xor U4546 (N_4546,N_3169,N_3356);
and U4547 (N_4547,N_3253,N_3478);
and U4548 (N_4548,N_3090,N_3966);
or U4549 (N_4549,N_3824,N_3758);
and U4550 (N_4550,N_3303,N_3161);
xnor U4551 (N_4551,N_3841,N_3377);
nand U4552 (N_4552,N_3447,N_3039);
or U4553 (N_4553,N_3242,N_3358);
xnor U4554 (N_4554,N_3384,N_3590);
xnor U4555 (N_4555,N_3245,N_3098);
xnor U4556 (N_4556,N_3427,N_3807);
nor U4557 (N_4557,N_3895,N_3344);
nand U4558 (N_4558,N_3108,N_3508);
xnor U4559 (N_4559,N_3275,N_3603);
xnor U4560 (N_4560,N_3799,N_3632);
xor U4561 (N_4561,N_3481,N_3309);
xnor U4562 (N_4562,N_3226,N_3332);
nand U4563 (N_4563,N_3940,N_3395);
xor U4564 (N_4564,N_3979,N_3731);
or U4565 (N_4565,N_3401,N_3758);
nand U4566 (N_4566,N_3099,N_3984);
nor U4567 (N_4567,N_3891,N_3942);
nor U4568 (N_4568,N_3086,N_3403);
xnor U4569 (N_4569,N_3490,N_3179);
and U4570 (N_4570,N_3369,N_3405);
xnor U4571 (N_4571,N_3515,N_3038);
and U4572 (N_4572,N_3647,N_3258);
xor U4573 (N_4573,N_3043,N_3283);
xor U4574 (N_4574,N_3546,N_3209);
or U4575 (N_4575,N_3846,N_3951);
xor U4576 (N_4576,N_3636,N_3714);
and U4577 (N_4577,N_3658,N_3286);
and U4578 (N_4578,N_3929,N_3782);
or U4579 (N_4579,N_3025,N_3800);
xnor U4580 (N_4580,N_3056,N_3482);
xnor U4581 (N_4581,N_3649,N_3644);
and U4582 (N_4582,N_3995,N_3545);
nand U4583 (N_4583,N_3113,N_3995);
and U4584 (N_4584,N_3382,N_3926);
nand U4585 (N_4585,N_3301,N_3583);
xor U4586 (N_4586,N_3166,N_3799);
nor U4587 (N_4587,N_3014,N_3016);
or U4588 (N_4588,N_3176,N_3809);
and U4589 (N_4589,N_3027,N_3795);
or U4590 (N_4590,N_3137,N_3410);
xor U4591 (N_4591,N_3047,N_3654);
nor U4592 (N_4592,N_3606,N_3532);
nand U4593 (N_4593,N_3501,N_3391);
nand U4594 (N_4594,N_3675,N_3357);
xor U4595 (N_4595,N_3587,N_3531);
nand U4596 (N_4596,N_3699,N_3351);
nor U4597 (N_4597,N_3749,N_3233);
nand U4598 (N_4598,N_3554,N_3803);
nor U4599 (N_4599,N_3333,N_3190);
xnor U4600 (N_4600,N_3661,N_3961);
or U4601 (N_4601,N_3916,N_3115);
nor U4602 (N_4602,N_3831,N_3128);
or U4603 (N_4603,N_3316,N_3642);
xor U4604 (N_4604,N_3873,N_3298);
xnor U4605 (N_4605,N_3744,N_3034);
nor U4606 (N_4606,N_3202,N_3375);
nand U4607 (N_4607,N_3924,N_3137);
and U4608 (N_4608,N_3673,N_3377);
xnor U4609 (N_4609,N_3936,N_3354);
nor U4610 (N_4610,N_3349,N_3028);
nand U4611 (N_4611,N_3667,N_3558);
xnor U4612 (N_4612,N_3747,N_3109);
and U4613 (N_4613,N_3254,N_3672);
nand U4614 (N_4614,N_3630,N_3131);
nor U4615 (N_4615,N_3604,N_3368);
or U4616 (N_4616,N_3541,N_3799);
and U4617 (N_4617,N_3347,N_3400);
and U4618 (N_4618,N_3983,N_3441);
nor U4619 (N_4619,N_3384,N_3799);
nand U4620 (N_4620,N_3725,N_3625);
and U4621 (N_4621,N_3311,N_3154);
xor U4622 (N_4622,N_3429,N_3048);
or U4623 (N_4623,N_3794,N_3345);
nand U4624 (N_4624,N_3547,N_3024);
or U4625 (N_4625,N_3383,N_3730);
and U4626 (N_4626,N_3363,N_3731);
and U4627 (N_4627,N_3894,N_3746);
nand U4628 (N_4628,N_3746,N_3772);
nand U4629 (N_4629,N_3696,N_3228);
nor U4630 (N_4630,N_3427,N_3317);
xor U4631 (N_4631,N_3437,N_3219);
and U4632 (N_4632,N_3945,N_3314);
nand U4633 (N_4633,N_3847,N_3676);
xor U4634 (N_4634,N_3895,N_3995);
xor U4635 (N_4635,N_3992,N_3466);
nand U4636 (N_4636,N_3076,N_3751);
nor U4637 (N_4637,N_3046,N_3815);
or U4638 (N_4638,N_3767,N_3460);
and U4639 (N_4639,N_3080,N_3024);
xor U4640 (N_4640,N_3062,N_3830);
and U4641 (N_4641,N_3920,N_3935);
nand U4642 (N_4642,N_3380,N_3661);
xor U4643 (N_4643,N_3501,N_3730);
xnor U4644 (N_4644,N_3657,N_3379);
and U4645 (N_4645,N_3971,N_3215);
or U4646 (N_4646,N_3935,N_3191);
nor U4647 (N_4647,N_3639,N_3129);
nor U4648 (N_4648,N_3023,N_3620);
nand U4649 (N_4649,N_3153,N_3901);
xor U4650 (N_4650,N_3061,N_3815);
nor U4651 (N_4651,N_3968,N_3315);
and U4652 (N_4652,N_3689,N_3559);
or U4653 (N_4653,N_3268,N_3110);
or U4654 (N_4654,N_3404,N_3186);
nor U4655 (N_4655,N_3686,N_3735);
or U4656 (N_4656,N_3214,N_3593);
and U4657 (N_4657,N_3782,N_3445);
and U4658 (N_4658,N_3415,N_3625);
nand U4659 (N_4659,N_3601,N_3770);
nor U4660 (N_4660,N_3966,N_3899);
or U4661 (N_4661,N_3208,N_3458);
xnor U4662 (N_4662,N_3836,N_3195);
nor U4663 (N_4663,N_3709,N_3571);
or U4664 (N_4664,N_3715,N_3981);
or U4665 (N_4665,N_3748,N_3717);
nand U4666 (N_4666,N_3899,N_3472);
and U4667 (N_4667,N_3874,N_3794);
xor U4668 (N_4668,N_3401,N_3034);
nor U4669 (N_4669,N_3975,N_3815);
and U4670 (N_4670,N_3531,N_3644);
xnor U4671 (N_4671,N_3416,N_3149);
or U4672 (N_4672,N_3525,N_3334);
and U4673 (N_4673,N_3465,N_3640);
nand U4674 (N_4674,N_3015,N_3232);
nand U4675 (N_4675,N_3413,N_3000);
or U4676 (N_4676,N_3732,N_3567);
nor U4677 (N_4677,N_3989,N_3893);
nor U4678 (N_4678,N_3871,N_3548);
nand U4679 (N_4679,N_3169,N_3479);
and U4680 (N_4680,N_3368,N_3081);
nor U4681 (N_4681,N_3906,N_3959);
nand U4682 (N_4682,N_3580,N_3570);
or U4683 (N_4683,N_3449,N_3737);
or U4684 (N_4684,N_3514,N_3100);
and U4685 (N_4685,N_3160,N_3047);
or U4686 (N_4686,N_3842,N_3849);
or U4687 (N_4687,N_3050,N_3888);
xnor U4688 (N_4688,N_3574,N_3267);
nor U4689 (N_4689,N_3860,N_3983);
nor U4690 (N_4690,N_3718,N_3851);
and U4691 (N_4691,N_3630,N_3694);
nand U4692 (N_4692,N_3561,N_3825);
or U4693 (N_4693,N_3201,N_3166);
xnor U4694 (N_4694,N_3777,N_3991);
nor U4695 (N_4695,N_3207,N_3018);
nand U4696 (N_4696,N_3212,N_3637);
nand U4697 (N_4697,N_3868,N_3377);
nand U4698 (N_4698,N_3253,N_3833);
xor U4699 (N_4699,N_3947,N_3758);
nand U4700 (N_4700,N_3177,N_3678);
and U4701 (N_4701,N_3358,N_3436);
and U4702 (N_4702,N_3493,N_3603);
nand U4703 (N_4703,N_3007,N_3272);
nand U4704 (N_4704,N_3189,N_3162);
and U4705 (N_4705,N_3685,N_3096);
nand U4706 (N_4706,N_3139,N_3421);
or U4707 (N_4707,N_3995,N_3035);
nor U4708 (N_4708,N_3176,N_3668);
nor U4709 (N_4709,N_3529,N_3247);
xnor U4710 (N_4710,N_3685,N_3406);
and U4711 (N_4711,N_3835,N_3124);
xor U4712 (N_4712,N_3686,N_3900);
or U4713 (N_4713,N_3963,N_3900);
or U4714 (N_4714,N_3227,N_3026);
or U4715 (N_4715,N_3579,N_3280);
nor U4716 (N_4716,N_3760,N_3046);
nand U4717 (N_4717,N_3308,N_3271);
nor U4718 (N_4718,N_3261,N_3546);
and U4719 (N_4719,N_3867,N_3521);
nand U4720 (N_4720,N_3612,N_3338);
nand U4721 (N_4721,N_3833,N_3907);
and U4722 (N_4722,N_3192,N_3113);
nor U4723 (N_4723,N_3933,N_3368);
and U4724 (N_4724,N_3185,N_3029);
nand U4725 (N_4725,N_3253,N_3665);
xor U4726 (N_4726,N_3380,N_3558);
nand U4727 (N_4727,N_3025,N_3640);
xor U4728 (N_4728,N_3499,N_3612);
or U4729 (N_4729,N_3693,N_3227);
nor U4730 (N_4730,N_3523,N_3924);
nand U4731 (N_4731,N_3237,N_3999);
xor U4732 (N_4732,N_3134,N_3271);
nor U4733 (N_4733,N_3751,N_3175);
xor U4734 (N_4734,N_3764,N_3035);
or U4735 (N_4735,N_3186,N_3834);
or U4736 (N_4736,N_3139,N_3916);
and U4737 (N_4737,N_3877,N_3085);
or U4738 (N_4738,N_3538,N_3326);
nor U4739 (N_4739,N_3409,N_3353);
and U4740 (N_4740,N_3578,N_3440);
or U4741 (N_4741,N_3201,N_3171);
and U4742 (N_4742,N_3597,N_3005);
xnor U4743 (N_4743,N_3253,N_3338);
and U4744 (N_4744,N_3579,N_3051);
or U4745 (N_4745,N_3960,N_3401);
xor U4746 (N_4746,N_3975,N_3605);
nand U4747 (N_4747,N_3406,N_3254);
and U4748 (N_4748,N_3033,N_3021);
xor U4749 (N_4749,N_3943,N_3485);
nor U4750 (N_4750,N_3853,N_3891);
xnor U4751 (N_4751,N_3833,N_3611);
or U4752 (N_4752,N_3597,N_3965);
nor U4753 (N_4753,N_3853,N_3223);
nor U4754 (N_4754,N_3089,N_3872);
nand U4755 (N_4755,N_3573,N_3206);
nand U4756 (N_4756,N_3512,N_3145);
or U4757 (N_4757,N_3147,N_3592);
nor U4758 (N_4758,N_3786,N_3492);
or U4759 (N_4759,N_3041,N_3624);
xnor U4760 (N_4760,N_3190,N_3219);
nor U4761 (N_4761,N_3253,N_3844);
nand U4762 (N_4762,N_3385,N_3433);
and U4763 (N_4763,N_3910,N_3478);
nand U4764 (N_4764,N_3941,N_3674);
and U4765 (N_4765,N_3621,N_3607);
nand U4766 (N_4766,N_3979,N_3077);
xor U4767 (N_4767,N_3584,N_3618);
nor U4768 (N_4768,N_3255,N_3367);
xnor U4769 (N_4769,N_3678,N_3164);
or U4770 (N_4770,N_3304,N_3325);
nand U4771 (N_4771,N_3247,N_3932);
nand U4772 (N_4772,N_3294,N_3196);
and U4773 (N_4773,N_3880,N_3146);
nor U4774 (N_4774,N_3583,N_3806);
or U4775 (N_4775,N_3760,N_3389);
nand U4776 (N_4776,N_3757,N_3758);
nor U4777 (N_4777,N_3364,N_3626);
and U4778 (N_4778,N_3883,N_3188);
xnor U4779 (N_4779,N_3412,N_3070);
and U4780 (N_4780,N_3054,N_3126);
nor U4781 (N_4781,N_3145,N_3771);
and U4782 (N_4782,N_3844,N_3885);
nand U4783 (N_4783,N_3184,N_3805);
and U4784 (N_4784,N_3998,N_3668);
xnor U4785 (N_4785,N_3369,N_3973);
xnor U4786 (N_4786,N_3990,N_3518);
or U4787 (N_4787,N_3159,N_3168);
xnor U4788 (N_4788,N_3100,N_3961);
or U4789 (N_4789,N_3620,N_3817);
xor U4790 (N_4790,N_3325,N_3197);
nor U4791 (N_4791,N_3128,N_3204);
xor U4792 (N_4792,N_3854,N_3664);
xnor U4793 (N_4793,N_3885,N_3328);
nand U4794 (N_4794,N_3510,N_3431);
and U4795 (N_4795,N_3620,N_3870);
or U4796 (N_4796,N_3963,N_3467);
or U4797 (N_4797,N_3890,N_3409);
or U4798 (N_4798,N_3170,N_3440);
nor U4799 (N_4799,N_3503,N_3272);
and U4800 (N_4800,N_3897,N_3303);
nor U4801 (N_4801,N_3537,N_3639);
nor U4802 (N_4802,N_3093,N_3440);
nand U4803 (N_4803,N_3401,N_3143);
nand U4804 (N_4804,N_3160,N_3361);
nand U4805 (N_4805,N_3292,N_3070);
and U4806 (N_4806,N_3240,N_3145);
nand U4807 (N_4807,N_3766,N_3812);
or U4808 (N_4808,N_3033,N_3326);
and U4809 (N_4809,N_3736,N_3333);
nor U4810 (N_4810,N_3534,N_3253);
and U4811 (N_4811,N_3431,N_3961);
or U4812 (N_4812,N_3326,N_3866);
xor U4813 (N_4813,N_3858,N_3068);
nor U4814 (N_4814,N_3996,N_3587);
xor U4815 (N_4815,N_3145,N_3044);
or U4816 (N_4816,N_3264,N_3935);
nand U4817 (N_4817,N_3013,N_3353);
xor U4818 (N_4818,N_3717,N_3517);
xor U4819 (N_4819,N_3009,N_3121);
and U4820 (N_4820,N_3934,N_3404);
xnor U4821 (N_4821,N_3337,N_3585);
and U4822 (N_4822,N_3640,N_3441);
xor U4823 (N_4823,N_3991,N_3196);
xnor U4824 (N_4824,N_3689,N_3564);
nor U4825 (N_4825,N_3614,N_3097);
nor U4826 (N_4826,N_3292,N_3466);
nor U4827 (N_4827,N_3634,N_3830);
and U4828 (N_4828,N_3757,N_3023);
nand U4829 (N_4829,N_3006,N_3032);
nand U4830 (N_4830,N_3107,N_3411);
nor U4831 (N_4831,N_3325,N_3378);
nor U4832 (N_4832,N_3409,N_3217);
xnor U4833 (N_4833,N_3262,N_3071);
and U4834 (N_4834,N_3223,N_3424);
nor U4835 (N_4835,N_3011,N_3516);
xnor U4836 (N_4836,N_3568,N_3006);
nor U4837 (N_4837,N_3588,N_3849);
or U4838 (N_4838,N_3953,N_3526);
or U4839 (N_4839,N_3988,N_3418);
or U4840 (N_4840,N_3044,N_3055);
nor U4841 (N_4841,N_3202,N_3304);
nand U4842 (N_4842,N_3364,N_3547);
nand U4843 (N_4843,N_3577,N_3429);
or U4844 (N_4844,N_3541,N_3588);
and U4845 (N_4845,N_3488,N_3029);
nor U4846 (N_4846,N_3734,N_3613);
nand U4847 (N_4847,N_3384,N_3385);
and U4848 (N_4848,N_3638,N_3404);
and U4849 (N_4849,N_3673,N_3527);
or U4850 (N_4850,N_3298,N_3108);
nor U4851 (N_4851,N_3599,N_3679);
nor U4852 (N_4852,N_3464,N_3975);
xnor U4853 (N_4853,N_3894,N_3252);
and U4854 (N_4854,N_3426,N_3853);
xnor U4855 (N_4855,N_3176,N_3458);
or U4856 (N_4856,N_3005,N_3883);
and U4857 (N_4857,N_3347,N_3685);
or U4858 (N_4858,N_3218,N_3022);
nor U4859 (N_4859,N_3294,N_3571);
or U4860 (N_4860,N_3021,N_3214);
nand U4861 (N_4861,N_3811,N_3588);
nor U4862 (N_4862,N_3215,N_3008);
and U4863 (N_4863,N_3938,N_3939);
and U4864 (N_4864,N_3269,N_3037);
xnor U4865 (N_4865,N_3574,N_3891);
or U4866 (N_4866,N_3507,N_3439);
or U4867 (N_4867,N_3542,N_3827);
nand U4868 (N_4868,N_3375,N_3769);
or U4869 (N_4869,N_3215,N_3774);
or U4870 (N_4870,N_3225,N_3025);
nand U4871 (N_4871,N_3479,N_3528);
and U4872 (N_4872,N_3476,N_3630);
nor U4873 (N_4873,N_3229,N_3364);
and U4874 (N_4874,N_3448,N_3618);
nand U4875 (N_4875,N_3988,N_3780);
nand U4876 (N_4876,N_3812,N_3304);
and U4877 (N_4877,N_3593,N_3471);
nor U4878 (N_4878,N_3862,N_3517);
nand U4879 (N_4879,N_3470,N_3268);
nand U4880 (N_4880,N_3189,N_3656);
and U4881 (N_4881,N_3104,N_3636);
xor U4882 (N_4882,N_3065,N_3125);
nand U4883 (N_4883,N_3372,N_3084);
nand U4884 (N_4884,N_3566,N_3305);
nor U4885 (N_4885,N_3050,N_3943);
nand U4886 (N_4886,N_3334,N_3495);
or U4887 (N_4887,N_3820,N_3127);
nand U4888 (N_4888,N_3367,N_3568);
or U4889 (N_4889,N_3218,N_3302);
xnor U4890 (N_4890,N_3191,N_3757);
nand U4891 (N_4891,N_3045,N_3173);
nor U4892 (N_4892,N_3189,N_3499);
nand U4893 (N_4893,N_3225,N_3527);
and U4894 (N_4894,N_3929,N_3843);
nor U4895 (N_4895,N_3647,N_3280);
nor U4896 (N_4896,N_3988,N_3860);
nor U4897 (N_4897,N_3168,N_3366);
nand U4898 (N_4898,N_3770,N_3625);
xor U4899 (N_4899,N_3604,N_3689);
xor U4900 (N_4900,N_3664,N_3700);
nor U4901 (N_4901,N_3739,N_3495);
nand U4902 (N_4902,N_3282,N_3598);
and U4903 (N_4903,N_3095,N_3707);
and U4904 (N_4904,N_3376,N_3016);
nand U4905 (N_4905,N_3157,N_3442);
nor U4906 (N_4906,N_3592,N_3813);
nand U4907 (N_4907,N_3743,N_3067);
or U4908 (N_4908,N_3488,N_3722);
nand U4909 (N_4909,N_3173,N_3092);
or U4910 (N_4910,N_3060,N_3133);
and U4911 (N_4911,N_3783,N_3199);
or U4912 (N_4912,N_3789,N_3730);
nand U4913 (N_4913,N_3749,N_3994);
xnor U4914 (N_4914,N_3563,N_3204);
xnor U4915 (N_4915,N_3829,N_3044);
nor U4916 (N_4916,N_3997,N_3119);
nand U4917 (N_4917,N_3940,N_3481);
and U4918 (N_4918,N_3272,N_3052);
nand U4919 (N_4919,N_3124,N_3431);
nor U4920 (N_4920,N_3766,N_3734);
xnor U4921 (N_4921,N_3918,N_3919);
nand U4922 (N_4922,N_3233,N_3759);
nand U4923 (N_4923,N_3209,N_3560);
xor U4924 (N_4924,N_3506,N_3422);
xor U4925 (N_4925,N_3825,N_3164);
or U4926 (N_4926,N_3914,N_3398);
and U4927 (N_4927,N_3003,N_3892);
xor U4928 (N_4928,N_3070,N_3154);
or U4929 (N_4929,N_3486,N_3284);
nand U4930 (N_4930,N_3941,N_3655);
and U4931 (N_4931,N_3547,N_3811);
nor U4932 (N_4932,N_3910,N_3105);
xor U4933 (N_4933,N_3843,N_3031);
nand U4934 (N_4934,N_3690,N_3593);
nand U4935 (N_4935,N_3855,N_3450);
nand U4936 (N_4936,N_3181,N_3361);
and U4937 (N_4937,N_3499,N_3706);
nand U4938 (N_4938,N_3705,N_3582);
or U4939 (N_4939,N_3787,N_3494);
xnor U4940 (N_4940,N_3654,N_3508);
or U4941 (N_4941,N_3508,N_3020);
or U4942 (N_4942,N_3121,N_3543);
nor U4943 (N_4943,N_3875,N_3526);
or U4944 (N_4944,N_3332,N_3231);
and U4945 (N_4945,N_3068,N_3619);
or U4946 (N_4946,N_3050,N_3000);
or U4947 (N_4947,N_3505,N_3267);
and U4948 (N_4948,N_3879,N_3768);
and U4949 (N_4949,N_3135,N_3636);
and U4950 (N_4950,N_3495,N_3962);
or U4951 (N_4951,N_3062,N_3489);
xor U4952 (N_4952,N_3010,N_3848);
xnor U4953 (N_4953,N_3001,N_3250);
nor U4954 (N_4954,N_3105,N_3440);
and U4955 (N_4955,N_3165,N_3483);
xor U4956 (N_4956,N_3229,N_3332);
and U4957 (N_4957,N_3871,N_3284);
nand U4958 (N_4958,N_3141,N_3825);
nand U4959 (N_4959,N_3420,N_3271);
or U4960 (N_4960,N_3162,N_3629);
nor U4961 (N_4961,N_3894,N_3418);
nand U4962 (N_4962,N_3660,N_3066);
xor U4963 (N_4963,N_3043,N_3493);
nor U4964 (N_4964,N_3397,N_3858);
xnor U4965 (N_4965,N_3728,N_3689);
xnor U4966 (N_4966,N_3477,N_3201);
and U4967 (N_4967,N_3106,N_3984);
xor U4968 (N_4968,N_3984,N_3428);
xor U4969 (N_4969,N_3684,N_3670);
nor U4970 (N_4970,N_3135,N_3433);
nor U4971 (N_4971,N_3100,N_3822);
nor U4972 (N_4972,N_3020,N_3315);
or U4973 (N_4973,N_3113,N_3863);
or U4974 (N_4974,N_3800,N_3153);
nand U4975 (N_4975,N_3336,N_3326);
and U4976 (N_4976,N_3588,N_3752);
nand U4977 (N_4977,N_3379,N_3531);
and U4978 (N_4978,N_3455,N_3028);
or U4979 (N_4979,N_3701,N_3416);
nand U4980 (N_4980,N_3940,N_3470);
or U4981 (N_4981,N_3201,N_3190);
and U4982 (N_4982,N_3606,N_3004);
or U4983 (N_4983,N_3413,N_3277);
xnor U4984 (N_4984,N_3988,N_3808);
or U4985 (N_4985,N_3036,N_3045);
nand U4986 (N_4986,N_3926,N_3373);
nand U4987 (N_4987,N_3488,N_3709);
xnor U4988 (N_4988,N_3248,N_3514);
xnor U4989 (N_4989,N_3188,N_3900);
or U4990 (N_4990,N_3977,N_3586);
nor U4991 (N_4991,N_3805,N_3067);
nand U4992 (N_4992,N_3414,N_3173);
xnor U4993 (N_4993,N_3493,N_3064);
or U4994 (N_4994,N_3126,N_3712);
xnor U4995 (N_4995,N_3019,N_3652);
or U4996 (N_4996,N_3110,N_3943);
nor U4997 (N_4997,N_3607,N_3063);
or U4998 (N_4998,N_3457,N_3861);
or U4999 (N_4999,N_3736,N_3826);
and U5000 (N_5000,N_4953,N_4891);
xnor U5001 (N_5001,N_4734,N_4050);
or U5002 (N_5002,N_4958,N_4048);
nor U5003 (N_5003,N_4866,N_4034);
nand U5004 (N_5004,N_4922,N_4004);
nand U5005 (N_5005,N_4143,N_4523);
xor U5006 (N_5006,N_4077,N_4967);
or U5007 (N_5007,N_4805,N_4752);
nand U5008 (N_5008,N_4309,N_4457);
or U5009 (N_5009,N_4336,N_4913);
or U5010 (N_5010,N_4701,N_4296);
nand U5011 (N_5011,N_4237,N_4773);
nor U5012 (N_5012,N_4769,N_4152);
xor U5013 (N_5013,N_4522,N_4629);
nor U5014 (N_5014,N_4973,N_4311);
nor U5015 (N_5015,N_4101,N_4995);
nor U5016 (N_5016,N_4212,N_4455);
xor U5017 (N_5017,N_4096,N_4124);
or U5018 (N_5018,N_4492,N_4470);
nor U5019 (N_5019,N_4510,N_4855);
nor U5020 (N_5020,N_4424,N_4809);
nor U5021 (N_5021,N_4007,N_4924);
xnor U5022 (N_5022,N_4477,N_4733);
nor U5023 (N_5023,N_4329,N_4977);
or U5024 (N_5024,N_4692,N_4886);
nand U5025 (N_5025,N_4756,N_4109);
nand U5026 (N_5026,N_4850,N_4175);
nor U5027 (N_5027,N_4353,N_4873);
nor U5028 (N_5028,N_4919,N_4060);
xor U5029 (N_5029,N_4578,N_4279);
nand U5030 (N_5030,N_4009,N_4204);
nand U5031 (N_5031,N_4509,N_4154);
and U5032 (N_5032,N_4747,N_4673);
nand U5033 (N_5033,N_4577,N_4306);
and U5034 (N_5034,N_4003,N_4650);
and U5035 (N_5035,N_4189,N_4615);
and U5036 (N_5036,N_4349,N_4384);
or U5037 (N_5037,N_4616,N_4837);
xnor U5038 (N_5038,N_4020,N_4851);
nand U5039 (N_5039,N_4759,N_4861);
and U5040 (N_5040,N_4671,N_4555);
and U5041 (N_5041,N_4064,N_4902);
nand U5042 (N_5042,N_4637,N_4613);
nand U5043 (N_5043,N_4153,N_4651);
or U5044 (N_5044,N_4184,N_4411);
nor U5045 (N_5045,N_4036,N_4225);
nor U5046 (N_5046,N_4920,N_4592);
nor U5047 (N_5047,N_4600,N_4707);
xor U5048 (N_5048,N_4682,N_4749);
nand U5049 (N_5049,N_4952,N_4361);
xnor U5050 (N_5050,N_4617,N_4541);
and U5051 (N_5051,N_4945,N_4338);
xor U5052 (N_5052,N_4303,N_4795);
xnor U5053 (N_5053,N_4081,N_4086);
or U5054 (N_5054,N_4818,N_4243);
nand U5055 (N_5055,N_4657,N_4833);
nand U5056 (N_5056,N_4224,N_4151);
and U5057 (N_5057,N_4943,N_4743);
nor U5058 (N_5058,N_4423,N_4986);
nor U5059 (N_5059,N_4881,N_4126);
nor U5060 (N_5060,N_4827,N_4915);
nand U5061 (N_5061,N_4770,N_4999);
or U5062 (N_5062,N_4929,N_4275);
nor U5063 (N_5063,N_4174,N_4794);
and U5064 (N_5064,N_4413,N_4829);
or U5065 (N_5065,N_4519,N_4343);
xor U5066 (N_5066,N_4711,N_4565);
xnor U5067 (N_5067,N_4830,N_4567);
nor U5068 (N_5068,N_4216,N_4508);
nor U5069 (N_5069,N_4543,N_4108);
xnor U5070 (N_5070,N_4382,N_4043);
nor U5071 (N_5071,N_4217,N_4718);
nor U5072 (N_5072,N_4813,N_4713);
or U5073 (N_5073,N_4019,N_4140);
and U5074 (N_5074,N_4193,N_4067);
or U5075 (N_5075,N_4878,N_4319);
nor U5076 (N_5076,N_4339,N_4645);
and U5077 (N_5077,N_4488,N_4797);
nor U5078 (N_5078,N_4038,N_4787);
nor U5079 (N_5079,N_4497,N_4642);
nor U5080 (N_5080,N_4901,N_4116);
xor U5081 (N_5081,N_4894,N_4857);
xnor U5082 (N_5082,N_4808,N_4277);
xor U5083 (N_5083,N_4027,N_4199);
nor U5084 (N_5084,N_4241,N_4934);
or U5085 (N_5085,N_4580,N_4087);
and U5086 (N_5086,N_4513,N_4284);
xor U5087 (N_5087,N_4438,N_4793);
nand U5088 (N_5088,N_4149,N_4935);
nand U5089 (N_5089,N_4334,N_4897);
nand U5090 (N_5090,N_4791,N_4993);
xnor U5091 (N_5091,N_4156,N_4778);
xnor U5092 (N_5092,N_4378,N_4582);
nand U5093 (N_5093,N_4176,N_4363);
xor U5094 (N_5094,N_4469,N_4017);
and U5095 (N_5095,N_4210,N_4679);
xnor U5096 (N_5096,N_4643,N_4820);
nor U5097 (N_5097,N_4804,N_4233);
nand U5098 (N_5098,N_4505,N_4232);
nor U5099 (N_5099,N_4005,N_4664);
nor U5100 (N_5100,N_4404,N_4948);
or U5101 (N_5101,N_4992,N_4052);
nor U5102 (N_5102,N_4507,N_4668);
or U5103 (N_5103,N_4843,N_4723);
nor U5104 (N_5104,N_4099,N_4313);
xnor U5105 (N_5105,N_4214,N_4937);
or U5106 (N_5106,N_4991,N_4148);
nor U5107 (N_5107,N_4355,N_4435);
nand U5108 (N_5108,N_4010,N_4364);
or U5109 (N_5109,N_4622,N_4185);
and U5110 (N_5110,N_4905,N_4740);
nor U5111 (N_5111,N_4766,N_4211);
and U5112 (N_5112,N_4688,N_4448);
nand U5113 (N_5113,N_4301,N_4796);
nand U5114 (N_5114,N_4655,N_4244);
and U5115 (N_5115,N_4842,N_4587);
nand U5116 (N_5116,N_4234,N_4367);
xor U5117 (N_5117,N_4408,N_4480);
nand U5118 (N_5118,N_4856,N_4771);
xnor U5119 (N_5119,N_4253,N_4931);
nor U5120 (N_5120,N_4160,N_4951);
xnor U5121 (N_5121,N_4606,N_4443);
nor U5122 (N_5122,N_4459,N_4100);
and U5123 (N_5123,N_4485,N_4240);
nand U5124 (N_5124,N_4235,N_4647);
nor U5125 (N_5125,N_4489,N_4868);
xor U5126 (N_5126,N_4517,N_4976);
and U5127 (N_5127,N_4325,N_4884);
or U5128 (N_5128,N_4854,N_4465);
and U5129 (N_5129,N_4798,N_4468);
xor U5130 (N_5130,N_4910,N_4428);
nand U5131 (N_5131,N_4129,N_4558);
xnor U5132 (N_5132,N_4903,N_4520);
nand U5133 (N_5133,N_4088,N_4663);
nand U5134 (N_5134,N_4144,N_4526);
xor U5135 (N_5135,N_4907,N_4104);
or U5136 (N_5136,N_4012,N_4524);
xor U5137 (N_5137,N_4464,N_4693);
xor U5138 (N_5138,N_4627,N_4539);
and U5139 (N_5139,N_4248,N_4178);
xnor U5140 (N_5140,N_4134,N_4848);
or U5141 (N_5141,N_4708,N_4705);
nand U5142 (N_5142,N_4187,N_4201);
nor U5143 (N_5143,N_4603,N_4841);
xnor U5144 (N_5144,N_4453,N_4754);
nor U5145 (N_5145,N_4638,N_4990);
or U5146 (N_5146,N_4365,N_4849);
or U5147 (N_5147,N_4700,N_4936);
and U5148 (N_5148,N_4712,N_4724);
xor U5149 (N_5149,N_4197,N_4258);
or U5150 (N_5150,N_4389,N_4691);
nand U5151 (N_5151,N_4345,N_4097);
or U5152 (N_5152,N_4699,N_4062);
nand U5153 (N_5153,N_4553,N_4788);
nand U5154 (N_5154,N_4521,N_4230);
and U5155 (N_5155,N_4737,N_4816);
nor U5156 (N_5156,N_4022,N_4231);
nand U5157 (N_5157,N_4481,N_4511);
and U5158 (N_5158,N_4860,N_4800);
or U5159 (N_5159,N_4262,N_4698);
or U5160 (N_5160,N_4653,N_4584);
nor U5161 (N_5161,N_4912,N_4709);
nand U5162 (N_5162,N_4792,N_4661);
nand U5163 (N_5163,N_4888,N_4568);
and U5164 (N_5164,N_4098,N_4726);
nor U5165 (N_5165,N_4786,N_4023);
xnor U5166 (N_5166,N_4076,N_4107);
xnor U5167 (N_5167,N_4066,N_4678);
xor U5168 (N_5168,N_4503,N_4748);
and U5169 (N_5169,N_4859,N_4342);
nand U5170 (N_5170,N_4205,N_4347);
and U5171 (N_5171,N_4422,N_4035);
and U5172 (N_5172,N_4670,N_4562);
nor U5173 (N_5173,N_4269,N_4890);
or U5174 (N_5174,N_4400,N_4581);
nand U5175 (N_5175,N_4839,N_4351);
or U5176 (N_5176,N_4121,N_4242);
xnor U5177 (N_5177,N_4760,N_4321);
or U5178 (N_5178,N_4728,N_4433);
nand U5179 (N_5179,N_4458,N_4652);
xnor U5180 (N_5180,N_4406,N_4304);
and U5181 (N_5181,N_4872,N_4028);
nand U5182 (N_5182,N_4405,N_4179);
nor U5183 (N_5183,N_4730,N_4495);
nand U5184 (N_5184,N_4180,N_4956);
xor U5185 (N_5185,N_4376,N_4278);
and U5186 (N_5186,N_4904,N_4844);
nor U5187 (N_5187,N_4683,N_4672);
nor U5188 (N_5188,N_4011,N_4646);
nand U5189 (N_5189,N_4970,N_4569);
or U5190 (N_5190,N_4989,N_4288);
nor U5191 (N_5191,N_4649,N_4535);
nor U5192 (N_5192,N_4331,N_4068);
or U5193 (N_5193,N_4946,N_4835);
or U5194 (N_5194,N_4467,N_4601);
nand U5195 (N_5195,N_4123,N_4282);
or U5196 (N_5196,N_4021,N_4291);
or U5197 (N_5197,N_4360,N_4083);
xor U5198 (N_5198,N_4255,N_4366);
nand U5199 (N_5199,N_4206,N_4430);
and U5200 (N_5200,N_4554,N_4263);
nor U5201 (N_5201,N_4298,N_4694);
nor U5202 (N_5202,N_4598,N_4681);
nor U5203 (N_5203,N_4528,N_4120);
nor U5204 (N_5204,N_4978,N_4559);
nor U5205 (N_5205,N_4172,N_4261);
and U5206 (N_5206,N_4130,N_4452);
nor U5207 (N_5207,N_4460,N_4239);
xor U5208 (N_5208,N_4611,N_4782);
and U5209 (N_5209,N_4079,N_4350);
nand U5210 (N_5210,N_4219,N_4473);
nor U5211 (N_5211,N_4359,N_4624);
nand U5212 (N_5212,N_4984,N_4639);
nor U5213 (N_5213,N_4665,N_4641);
nor U5214 (N_5214,N_4354,N_4719);
xor U5215 (N_5215,N_4714,N_4001);
xnor U5216 (N_5216,N_4985,N_4292);
nor U5217 (N_5217,N_4783,N_4092);
and U5218 (N_5218,N_4802,N_4466);
nand U5219 (N_5219,N_4625,N_4768);
or U5220 (N_5220,N_4078,N_4871);
xor U5221 (N_5221,N_4784,N_4572);
nor U5222 (N_5222,N_4640,N_4266);
nand U5223 (N_5223,N_4479,N_4105);
and U5224 (N_5224,N_4832,N_4727);
nand U5225 (N_5225,N_4826,N_4863);
nor U5226 (N_5226,N_4227,N_4744);
nand U5227 (N_5227,N_4381,N_4139);
or U5228 (N_5228,N_4751,N_4290);
and U5229 (N_5229,N_4772,N_4316);
xnor U5230 (N_5230,N_4941,N_4514);
or U5231 (N_5231,N_4142,N_4373);
and U5232 (N_5232,N_4811,N_4371);
and U5233 (N_5233,N_4735,N_4732);
nor U5234 (N_5234,N_4044,N_4516);
xnor U5235 (N_5235,N_4383,N_4075);
or U5236 (N_5236,N_4051,N_4574);
nor U5237 (N_5237,N_4324,N_4446);
xor U5238 (N_5238,N_4182,N_4566);
xor U5239 (N_5239,N_4379,N_4536);
nor U5240 (N_5240,N_4504,N_4780);
xor U5241 (N_5241,N_4057,N_4352);
nor U5242 (N_5242,N_4071,N_4385);
or U5243 (N_5243,N_4715,N_4660);
or U5244 (N_5244,N_4779,N_4300);
nor U5245 (N_5245,N_4529,N_4229);
xor U5246 (N_5246,N_4630,N_4418);
xnor U5247 (N_5247,N_4621,N_4133);
or U5248 (N_5248,N_4445,N_4801);
xnor U5249 (N_5249,N_4082,N_4447);
and U5250 (N_5250,N_4138,N_4059);
or U5251 (N_5251,N_4375,N_4131);
nand U5252 (N_5252,N_4450,N_4765);
nor U5253 (N_5253,N_4401,N_4703);
or U5254 (N_5254,N_4965,N_4061);
xor U5255 (N_5255,N_4073,N_4542);
or U5256 (N_5256,N_4315,N_4979);
and U5257 (N_5257,N_4106,N_4150);
and U5258 (N_5258,N_4158,N_4393);
and U5259 (N_5259,N_4456,N_4686);
xor U5260 (N_5260,N_4250,N_4357);
or U5261 (N_5261,N_4103,N_4675);
and U5262 (N_5262,N_4968,N_4918);
nor U5263 (N_5263,N_4631,N_4215);
or U5264 (N_5264,N_4746,N_4065);
nand U5265 (N_5265,N_4525,N_4824);
nand U5266 (N_5266,N_4398,N_4272);
xnor U5267 (N_5267,N_4380,N_4619);
or U5268 (N_5268,N_4238,N_4560);
nand U5269 (N_5269,N_4896,N_4926);
nor U5270 (N_5270,N_4940,N_4397);
nor U5271 (N_5271,N_4432,N_4648);
nor U5272 (N_5272,N_4399,N_4895);
nor U5273 (N_5273,N_4596,N_4392);
or U5274 (N_5274,N_4425,N_4122);
and U5275 (N_5275,N_4114,N_4685);
nor U5276 (N_5276,N_4717,N_4125);
nor U5277 (N_5277,N_4169,N_4825);
and U5278 (N_5278,N_4259,N_4982);
and U5279 (N_5279,N_4320,N_4420);
nand U5280 (N_5280,N_4449,N_4145);
and U5281 (N_5281,N_4203,N_4222);
xnor U5282 (N_5282,N_4118,N_4763);
nand U5283 (N_5283,N_4191,N_4720);
and U5284 (N_5284,N_4932,N_4869);
nor U5285 (N_5285,N_4190,N_4200);
or U5286 (N_5286,N_4476,N_4207);
nand U5287 (N_5287,N_4531,N_4341);
xor U5288 (N_5288,N_4530,N_4218);
and U5289 (N_5289,N_4595,N_4370);
nand U5290 (N_5290,N_4757,N_4274);
or U5291 (N_5291,N_4112,N_4745);
and U5292 (N_5292,N_4161,N_4391);
xnor U5293 (N_5293,N_4170,N_4208);
nor U5294 (N_5294,N_4486,N_4593);
nand U5295 (N_5295,N_4533,N_4494);
nand U5296 (N_5296,N_4113,N_4271);
xnor U5297 (N_5297,N_4484,N_4308);
nor U5298 (N_5298,N_4602,N_4966);
and U5299 (N_5299,N_4534,N_4729);
and U5300 (N_5300,N_4573,N_4579);
xor U5301 (N_5301,N_4908,N_4047);
and U5302 (N_5302,N_4472,N_4295);
nor U5303 (N_5303,N_4268,N_4846);
and U5304 (N_5304,N_4039,N_4944);
or U5305 (N_5305,N_4556,N_4527);
and U5306 (N_5306,N_4273,N_4662);
nor U5307 (N_5307,N_4564,N_4666);
xnor U5308 (N_5308,N_4736,N_4018);
xnor U5309 (N_5309,N_4141,N_4257);
and U5310 (N_5310,N_4583,N_4847);
nand U5311 (N_5311,N_4789,N_4988);
xnor U5312 (N_5312,N_4998,N_4026);
nor U5313 (N_5313,N_4997,N_4454);
and U5314 (N_5314,N_4680,N_4249);
nand U5315 (N_5315,N_4594,N_4429);
and U5316 (N_5316,N_4867,N_4500);
and U5317 (N_5317,N_4314,N_4310);
and U5318 (N_5318,N_4858,N_4089);
or U5319 (N_5319,N_4753,N_4323);
or U5320 (N_5320,N_4307,N_4000);
xor U5321 (N_5321,N_4202,N_4159);
nor U5322 (N_5322,N_4407,N_4147);
or U5323 (N_5323,N_4676,N_4821);
nand U5324 (N_5324,N_4247,N_4815);
xnor U5325 (N_5325,N_4403,N_4585);
nand U5326 (N_5326,N_4644,N_4550);
nand U5327 (N_5327,N_4845,N_4911);
and U5328 (N_5328,N_4111,N_4030);
or U5329 (N_5329,N_4416,N_4546);
and U5330 (N_5330,N_4634,N_4410);
and U5331 (N_5331,N_4725,N_4938);
or U5332 (N_5332,N_4590,N_4136);
or U5333 (N_5333,N_4177,N_4132);
and U5334 (N_5334,N_4223,N_4862);
nor U5335 (N_5335,N_4803,N_4168);
nor U5336 (N_5336,N_4927,N_4195);
nor U5337 (N_5337,N_4474,N_4939);
xnor U5338 (N_5338,N_4194,N_4612);
xnor U5339 (N_5339,N_4289,N_4914);
xor U5340 (N_5340,N_4610,N_4015);
or U5341 (N_5341,N_4540,N_4591);
and U5342 (N_5342,N_4337,N_4006);
nand U5343 (N_5343,N_4971,N_4762);
xnor U5344 (N_5344,N_4186,N_4016);
nor U5345 (N_5345,N_4969,N_4409);
and U5346 (N_5346,N_4776,N_4014);
nand U5347 (N_5347,N_4807,N_4117);
nor U5348 (N_5348,N_4395,N_4276);
nor U5349 (N_5349,N_4374,N_4388);
nor U5350 (N_5350,N_4689,N_4983);
and U5351 (N_5351,N_4876,N_4575);
or U5352 (N_5352,N_4942,N_4426);
nand U5353 (N_5353,N_4002,N_4716);
nand U5354 (N_5354,N_4742,N_4302);
nand U5355 (N_5355,N_4346,N_4236);
and U5356 (N_5356,N_4532,N_4974);
nand U5357 (N_5357,N_4695,N_4930);
or U5358 (N_5358,N_4055,N_4690);
xnor U5359 (N_5359,N_4348,N_4963);
and U5360 (N_5360,N_4221,N_4155);
nand U5361 (N_5361,N_4961,N_4632);
nand U5362 (N_5362,N_4072,N_4260);
or U5363 (N_5363,N_4491,N_4264);
nor U5364 (N_5364,N_4928,N_4070);
nor U5365 (N_5365,N_4333,N_4777);
nand U5366 (N_5366,N_4741,N_4879);
or U5367 (N_5367,N_4127,N_4386);
nor U5368 (N_5368,N_4933,N_4687);
and U5369 (N_5369,N_4317,N_4252);
and U5370 (N_5370,N_4722,N_4128);
nand U5371 (N_5371,N_4571,N_4774);
nand U5372 (N_5372,N_4318,N_4515);
nor U5373 (N_5373,N_4220,N_4164);
and U5374 (N_5374,N_4623,N_4885);
nor U5375 (N_5375,N_4335,N_4604);
nor U5376 (N_5376,N_4436,N_4823);
and U5377 (N_5377,N_4498,N_4954);
nand U5378 (N_5378,N_4656,N_4074);
xor U5379 (N_5379,N_4041,N_4293);
and U5380 (N_5380,N_4487,N_4909);
nand U5381 (N_5381,N_4659,N_4029);
nor U5382 (N_5382,N_4865,N_4955);
nor U5383 (N_5383,N_4758,N_4483);
nand U5384 (N_5384,N_4586,N_4957);
or U5385 (N_5385,N_4674,N_4167);
or U5386 (N_5386,N_4084,N_4281);
and U5387 (N_5387,N_4166,N_4297);
and U5388 (N_5388,N_4790,N_4892);
and U5389 (N_5389,N_4462,N_4045);
or U5390 (N_5390,N_4058,N_4040);
and U5391 (N_5391,N_4704,N_4093);
and U5392 (N_5392,N_4056,N_4923);
nand U5393 (N_5393,N_4960,N_4549);
nand U5394 (N_5394,N_4270,N_4327);
and U5395 (N_5395,N_4090,N_4738);
xor U5396 (N_5396,N_4377,N_4980);
nor U5397 (N_5397,N_4192,N_4094);
or U5398 (N_5398,N_4607,N_4209);
nor U5399 (N_5399,N_4570,N_4358);
or U5400 (N_5400,N_4119,N_4431);
xnor U5401 (N_5401,N_4024,N_4173);
nand U5402 (N_5402,N_4852,N_4667);
nand U5403 (N_5403,N_4394,N_4654);
nand U5404 (N_5404,N_4135,N_4755);
xor U5405 (N_5405,N_4981,N_4390);
nand U5406 (N_5406,N_4563,N_4506);
nor U5407 (N_5407,N_4947,N_4283);
nand U5408 (N_5408,N_4697,N_4183);
nor U5409 (N_5409,N_4775,N_4677);
xor U5410 (N_5410,N_4949,N_4095);
nand U5411 (N_5411,N_4490,N_4332);
or U5412 (N_5412,N_4893,N_4840);
and U5413 (N_5413,N_4702,N_4165);
xnor U5414 (N_5414,N_4870,N_4254);
and U5415 (N_5415,N_4146,N_4972);
and U5416 (N_5416,N_4368,N_4496);
or U5417 (N_5417,N_4764,N_4372);
nor U5418 (N_5418,N_4557,N_4538);
or U5419 (N_5419,N_4356,N_4620);
xor U5420 (N_5420,N_4157,N_4493);
xnor U5421 (N_5421,N_4501,N_4696);
and U5422 (N_5422,N_4280,N_4305);
nand U5423 (N_5423,N_4031,N_4599);
or U5424 (N_5424,N_4589,N_4286);
and U5425 (N_5425,N_4806,N_4414);
nand U5426 (N_5426,N_4330,N_4987);
and U5427 (N_5427,N_4442,N_4387);
nor U5428 (N_5428,N_4545,N_4883);
and U5429 (N_5429,N_4042,N_4950);
or U5430 (N_5430,N_4518,N_4880);
xnor U5431 (N_5431,N_4959,N_4441);
xnor U5432 (N_5432,N_4710,N_4080);
nor U5433 (N_5433,N_4887,N_4917);
nand U5434 (N_5434,N_4256,N_4294);
or U5435 (N_5435,N_4482,N_4576);
nor U5436 (N_5436,N_4322,N_4063);
or U5437 (N_5437,N_4475,N_4921);
or U5438 (N_5438,N_4033,N_4437);
xnor U5439 (N_5439,N_4588,N_4461);
and U5440 (N_5440,N_4669,N_4819);
xor U5441 (N_5441,N_4471,N_4781);
and U5442 (N_5442,N_4633,N_4421);
nor U5443 (N_5443,N_4402,N_4925);
xor U5444 (N_5444,N_4053,N_4608);
and U5445 (N_5445,N_4046,N_4721);
xnor U5446 (N_5446,N_4636,N_4162);
xnor U5447 (N_5447,N_4344,N_4605);
xnor U5448 (N_5448,N_4226,N_4434);
nand U5449 (N_5449,N_4171,N_4312);
xor U5450 (N_5450,N_4996,N_4882);
nor U5451 (N_5451,N_4750,N_4551);
and U5452 (N_5452,N_4512,N_4417);
xor U5453 (N_5453,N_4013,N_4032);
xor U5454 (N_5454,N_4362,N_4799);
or U5455 (N_5455,N_4810,N_4906);
nor U5456 (N_5456,N_4444,N_4396);
nor U5457 (N_5457,N_4463,N_4814);
nand U5458 (N_5458,N_4163,N_4916);
nand U5459 (N_5459,N_4761,N_4635);
xor U5460 (N_5460,N_4609,N_4265);
or U5461 (N_5461,N_4548,N_4085);
nor U5462 (N_5462,N_4299,N_4054);
nor U5463 (N_5463,N_4767,N_4544);
or U5464 (N_5464,N_4836,N_4706);
xnor U5465 (N_5465,N_4340,N_4137);
xnor U5466 (N_5466,N_4110,N_4834);
nor U5467 (N_5467,N_4864,N_4049);
or U5468 (N_5468,N_4889,N_4427);
nor U5469 (N_5469,N_4419,N_4552);
or U5470 (N_5470,N_4196,N_4037);
nand U5471 (N_5471,N_4213,N_4251);
nor U5472 (N_5472,N_4069,N_4246);
and U5473 (N_5473,N_4439,N_4267);
xor U5474 (N_5474,N_4188,N_4181);
nor U5475 (N_5475,N_4478,N_4561);
nand U5476 (N_5476,N_4626,N_4628);
nor U5477 (N_5477,N_4817,N_4008);
nor U5478 (N_5478,N_4285,N_4328);
nand U5479 (N_5479,N_4228,N_4369);
or U5480 (N_5480,N_4962,N_4975);
or U5481 (N_5481,N_4874,N_4731);
nor U5482 (N_5482,N_4287,N_4994);
nand U5483 (N_5483,N_4547,N_4440);
or U5484 (N_5484,N_4415,N_4115);
and U5485 (N_5485,N_4831,N_4198);
and U5486 (N_5486,N_4499,N_4102);
nor U5487 (N_5487,N_4899,N_4326);
nand U5488 (N_5488,N_4875,N_4877);
or U5489 (N_5489,N_4898,N_4245);
xor U5490 (N_5490,N_4412,N_4812);
nand U5491 (N_5491,N_4091,N_4853);
nand U5492 (N_5492,N_4025,N_4822);
xor U5493 (N_5493,N_4614,N_4658);
nor U5494 (N_5494,N_4451,N_4502);
nand U5495 (N_5495,N_4537,N_4785);
nand U5496 (N_5496,N_4739,N_4964);
xnor U5497 (N_5497,N_4618,N_4828);
nand U5498 (N_5498,N_4597,N_4900);
nand U5499 (N_5499,N_4838,N_4684);
nor U5500 (N_5500,N_4679,N_4823);
xnor U5501 (N_5501,N_4652,N_4724);
and U5502 (N_5502,N_4007,N_4824);
xnor U5503 (N_5503,N_4029,N_4824);
or U5504 (N_5504,N_4075,N_4458);
nand U5505 (N_5505,N_4035,N_4393);
xor U5506 (N_5506,N_4091,N_4610);
and U5507 (N_5507,N_4465,N_4042);
nand U5508 (N_5508,N_4471,N_4472);
nor U5509 (N_5509,N_4858,N_4994);
nor U5510 (N_5510,N_4290,N_4178);
xor U5511 (N_5511,N_4063,N_4467);
and U5512 (N_5512,N_4406,N_4886);
or U5513 (N_5513,N_4739,N_4668);
nor U5514 (N_5514,N_4137,N_4373);
nand U5515 (N_5515,N_4014,N_4109);
and U5516 (N_5516,N_4681,N_4944);
or U5517 (N_5517,N_4966,N_4518);
or U5518 (N_5518,N_4909,N_4924);
nor U5519 (N_5519,N_4727,N_4454);
or U5520 (N_5520,N_4587,N_4593);
and U5521 (N_5521,N_4344,N_4061);
nand U5522 (N_5522,N_4970,N_4511);
nand U5523 (N_5523,N_4994,N_4971);
nand U5524 (N_5524,N_4461,N_4938);
xor U5525 (N_5525,N_4170,N_4806);
and U5526 (N_5526,N_4711,N_4639);
and U5527 (N_5527,N_4917,N_4076);
and U5528 (N_5528,N_4936,N_4928);
nor U5529 (N_5529,N_4936,N_4784);
nor U5530 (N_5530,N_4538,N_4280);
or U5531 (N_5531,N_4361,N_4027);
nand U5532 (N_5532,N_4390,N_4936);
nand U5533 (N_5533,N_4301,N_4012);
nand U5534 (N_5534,N_4159,N_4113);
xor U5535 (N_5535,N_4978,N_4039);
nor U5536 (N_5536,N_4039,N_4203);
xnor U5537 (N_5537,N_4461,N_4347);
or U5538 (N_5538,N_4529,N_4614);
or U5539 (N_5539,N_4380,N_4663);
xnor U5540 (N_5540,N_4774,N_4516);
nor U5541 (N_5541,N_4836,N_4496);
and U5542 (N_5542,N_4881,N_4285);
or U5543 (N_5543,N_4298,N_4445);
nand U5544 (N_5544,N_4296,N_4989);
or U5545 (N_5545,N_4892,N_4517);
xor U5546 (N_5546,N_4015,N_4683);
or U5547 (N_5547,N_4739,N_4517);
and U5548 (N_5548,N_4065,N_4608);
nand U5549 (N_5549,N_4647,N_4534);
nand U5550 (N_5550,N_4160,N_4469);
nor U5551 (N_5551,N_4725,N_4109);
nor U5552 (N_5552,N_4128,N_4379);
or U5553 (N_5553,N_4922,N_4759);
nand U5554 (N_5554,N_4479,N_4706);
and U5555 (N_5555,N_4800,N_4439);
or U5556 (N_5556,N_4620,N_4478);
or U5557 (N_5557,N_4851,N_4988);
or U5558 (N_5558,N_4916,N_4490);
or U5559 (N_5559,N_4835,N_4458);
nor U5560 (N_5560,N_4088,N_4362);
or U5561 (N_5561,N_4158,N_4178);
nor U5562 (N_5562,N_4240,N_4214);
nand U5563 (N_5563,N_4447,N_4165);
and U5564 (N_5564,N_4559,N_4183);
nor U5565 (N_5565,N_4379,N_4765);
and U5566 (N_5566,N_4965,N_4926);
nand U5567 (N_5567,N_4293,N_4657);
or U5568 (N_5568,N_4156,N_4353);
or U5569 (N_5569,N_4789,N_4209);
xnor U5570 (N_5570,N_4575,N_4610);
nor U5571 (N_5571,N_4584,N_4635);
nor U5572 (N_5572,N_4599,N_4859);
nor U5573 (N_5573,N_4873,N_4862);
nor U5574 (N_5574,N_4574,N_4818);
and U5575 (N_5575,N_4225,N_4453);
or U5576 (N_5576,N_4194,N_4888);
nand U5577 (N_5577,N_4808,N_4406);
nor U5578 (N_5578,N_4900,N_4799);
nor U5579 (N_5579,N_4840,N_4547);
and U5580 (N_5580,N_4160,N_4664);
nor U5581 (N_5581,N_4738,N_4932);
or U5582 (N_5582,N_4414,N_4307);
nor U5583 (N_5583,N_4248,N_4044);
or U5584 (N_5584,N_4508,N_4419);
and U5585 (N_5585,N_4513,N_4905);
nor U5586 (N_5586,N_4427,N_4759);
or U5587 (N_5587,N_4400,N_4328);
or U5588 (N_5588,N_4242,N_4795);
xor U5589 (N_5589,N_4667,N_4621);
xnor U5590 (N_5590,N_4453,N_4572);
xor U5591 (N_5591,N_4811,N_4931);
xor U5592 (N_5592,N_4113,N_4977);
or U5593 (N_5593,N_4910,N_4439);
and U5594 (N_5594,N_4929,N_4455);
and U5595 (N_5595,N_4243,N_4728);
or U5596 (N_5596,N_4745,N_4070);
and U5597 (N_5597,N_4365,N_4686);
xor U5598 (N_5598,N_4161,N_4178);
or U5599 (N_5599,N_4293,N_4125);
xnor U5600 (N_5600,N_4152,N_4517);
xnor U5601 (N_5601,N_4400,N_4412);
nor U5602 (N_5602,N_4919,N_4859);
or U5603 (N_5603,N_4175,N_4202);
xor U5604 (N_5604,N_4290,N_4169);
xor U5605 (N_5605,N_4857,N_4189);
xnor U5606 (N_5606,N_4057,N_4052);
nand U5607 (N_5607,N_4050,N_4189);
nor U5608 (N_5608,N_4472,N_4425);
or U5609 (N_5609,N_4462,N_4940);
or U5610 (N_5610,N_4969,N_4079);
or U5611 (N_5611,N_4230,N_4684);
nor U5612 (N_5612,N_4615,N_4000);
xnor U5613 (N_5613,N_4152,N_4287);
nor U5614 (N_5614,N_4367,N_4282);
and U5615 (N_5615,N_4827,N_4253);
nor U5616 (N_5616,N_4682,N_4827);
nand U5617 (N_5617,N_4648,N_4525);
nor U5618 (N_5618,N_4323,N_4763);
and U5619 (N_5619,N_4327,N_4216);
and U5620 (N_5620,N_4761,N_4580);
and U5621 (N_5621,N_4323,N_4863);
or U5622 (N_5622,N_4805,N_4647);
or U5623 (N_5623,N_4453,N_4632);
nor U5624 (N_5624,N_4809,N_4101);
nand U5625 (N_5625,N_4054,N_4250);
nor U5626 (N_5626,N_4639,N_4214);
xnor U5627 (N_5627,N_4948,N_4712);
nand U5628 (N_5628,N_4453,N_4585);
xor U5629 (N_5629,N_4433,N_4923);
or U5630 (N_5630,N_4341,N_4826);
or U5631 (N_5631,N_4971,N_4624);
or U5632 (N_5632,N_4257,N_4976);
nand U5633 (N_5633,N_4951,N_4579);
xor U5634 (N_5634,N_4943,N_4912);
and U5635 (N_5635,N_4948,N_4768);
and U5636 (N_5636,N_4261,N_4332);
nor U5637 (N_5637,N_4993,N_4571);
nand U5638 (N_5638,N_4966,N_4285);
xor U5639 (N_5639,N_4830,N_4318);
or U5640 (N_5640,N_4494,N_4061);
nand U5641 (N_5641,N_4485,N_4261);
nor U5642 (N_5642,N_4953,N_4304);
or U5643 (N_5643,N_4053,N_4244);
nand U5644 (N_5644,N_4816,N_4658);
xor U5645 (N_5645,N_4706,N_4214);
and U5646 (N_5646,N_4141,N_4136);
and U5647 (N_5647,N_4662,N_4645);
xnor U5648 (N_5648,N_4461,N_4323);
or U5649 (N_5649,N_4068,N_4379);
nor U5650 (N_5650,N_4672,N_4637);
nand U5651 (N_5651,N_4315,N_4679);
and U5652 (N_5652,N_4870,N_4289);
and U5653 (N_5653,N_4919,N_4829);
and U5654 (N_5654,N_4974,N_4650);
nand U5655 (N_5655,N_4641,N_4521);
or U5656 (N_5656,N_4479,N_4910);
and U5657 (N_5657,N_4270,N_4124);
xor U5658 (N_5658,N_4017,N_4676);
nand U5659 (N_5659,N_4862,N_4266);
and U5660 (N_5660,N_4564,N_4126);
and U5661 (N_5661,N_4018,N_4257);
and U5662 (N_5662,N_4868,N_4242);
xor U5663 (N_5663,N_4188,N_4602);
xnor U5664 (N_5664,N_4942,N_4527);
nor U5665 (N_5665,N_4255,N_4488);
and U5666 (N_5666,N_4170,N_4459);
xor U5667 (N_5667,N_4190,N_4447);
nand U5668 (N_5668,N_4468,N_4125);
nor U5669 (N_5669,N_4385,N_4959);
or U5670 (N_5670,N_4262,N_4571);
xor U5671 (N_5671,N_4666,N_4953);
nand U5672 (N_5672,N_4850,N_4817);
xor U5673 (N_5673,N_4292,N_4162);
nand U5674 (N_5674,N_4520,N_4302);
and U5675 (N_5675,N_4728,N_4068);
nor U5676 (N_5676,N_4969,N_4057);
xor U5677 (N_5677,N_4986,N_4140);
and U5678 (N_5678,N_4193,N_4715);
or U5679 (N_5679,N_4915,N_4394);
and U5680 (N_5680,N_4585,N_4796);
xnor U5681 (N_5681,N_4141,N_4030);
or U5682 (N_5682,N_4814,N_4298);
or U5683 (N_5683,N_4757,N_4569);
or U5684 (N_5684,N_4644,N_4802);
and U5685 (N_5685,N_4839,N_4853);
nor U5686 (N_5686,N_4005,N_4250);
nor U5687 (N_5687,N_4685,N_4104);
xnor U5688 (N_5688,N_4946,N_4546);
xor U5689 (N_5689,N_4201,N_4986);
nor U5690 (N_5690,N_4221,N_4175);
xor U5691 (N_5691,N_4307,N_4051);
xnor U5692 (N_5692,N_4110,N_4910);
xor U5693 (N_5693,N_4209,N_4780);
nor U5694 (N_5694,N_4418,N_4310);
nor U5695 (N_5695,N_4477,N_4005);
nand U5696 (N_5696,N_4787,N_4390);
xor U5697 (N_5697,N_4066,N_4294);
nor U5698 (N_5698,N_4527,N_4204);
nand U5699 (N_5699,N_4590,N_4623);
or U5700 (N_5700,N_4909,N_4812);
nand U5701 (N_5701,N_4287,N_4768);
nand U5702 (N_5702,N_4474,N_4130);
xor U5703 (N_5703,N_4905,N_4813);
nor U5704 (N_5704,N_4540,N_4069);
or U5705 (N_5705,N_4073,N_4030);
xnor U5706 (N_5706,N_4713,N_4188);
and U5707 (N_5707,N_4907,N_4203);
and U5708 (N_5708,N_4558,N_4992);
xnor U5709 (N_5709,N_4172,N_4325);
xor U5710 (N_5710,N_4493,N_4942);
and U5711 (N_5711,N_4834,N_4437);
xor U5712 (N_5712,N_4254,N_4732);
nand U5713 (N_5713,N_4509,N_4486);
xnor U5714 (N_5714,N_4537,N_4004);
nor U5715 (N_5715,N_4532,N_4942);
nor U5716 (N_5716,N_4018,N_4850);
and U5717 (N_5717,N_4599,N_4990);
and U5718 (N_5718,N_4560,N_4303);
nor U5719 (N_5719,N_4931,N_4306);
nor U5720 (N_5720,N_4606,N_4672);
and U5721 (N_5721,N_4199,N_4010);
or U5722 (N_5722,N_4759,N_4031);
and U5723 (N_5723,N_4347,N_4725);
nor U5724 (N_5724,N_4157,N_4585);
nor U5725 (N_5725,N_4600,N_4817);
nor U5726 (N_5726,N_4239,N_4961);
nor U5727 (N_5727,N_4304,N_4435);
and U5728 (N_5728,N_4005,N_4403);
and U5729 (N_5729,N_4776,N_4150);
or U5730 (N_5730,N_4488,N_4280);
and U5731 (N_5731,N_4141,N_4010);
nor U5732 (N_5732,N_4320,N_4160);
or U5733 (N_5733,N_4709,N_4882);
nor U5734 (N_5734,N_4681,N_4320);
nor U5735 (N_5735,N_4717,N_4004);
nand U5736 (N_5736,N_4521,N_4354);
nand U5737 (N_5737,N_4971,N_4225);
nand U5738 (N_5738,N_4632,N_4805);
and U5739 (N_5739,N_4393,N_4093);
nand U5740 (N_5740,N_4360,N_4757);
nand U5741 (N_5741,N_4731,N_4017);
and U5742 (N_5742,N_4821,N_4831);
nor U5743 (N_5743,N_4737,N_4005);
nor U5744 (N_5744,N_4132,N_4681);
and U5745 (N_5745,N_4867,N_4566);
and U5746 (N_5746,N_4442,N_4143);
or U5747 (N_5747,N_4408,N_4263);
or U5748 (N_5748,N_4199,N_4710);
nor U5749 (N_5749,N_4458,N_4840);
xor U5750 (N_5750,N_4572,N_4903);
and U5751 (N_5751,N_4596,N_4860);
nand U5752 (N_5752,N_4687,N_4969);
nor U5753 (N_5753,N_4374,N_4324);
or U5754 (N_5754,N_4082,N_4022);
and U5755 (N_5755,N_4273,N_4833);
nand U5756 (N_5756,N_4992,N_4982);
xor U5757 (N_5757,N_4716,N_4929);
or U5758 (N_5758,N_4074,N_4689);
and U5759 (N_5759,N_4681,N_4821);
xor U5760 (N_5760,N_4253,N_4884);
and U5761 (N_5761,N_4708,N_4100);
or U5762 (N_5762,N_4233,N_4812);
or U5763 (N_5763,N_4315,N_4133);
and U5764 (N_5764,N_4149,N_4017);
nand U5765 (N_5765,N_4967,N_4469);
nand U5766 (N_5766,N_4884,N_4349);
nor U5767 (N_5767,N_4120,N_4461);
nand U5768 (N_5768,N_4453,N_4261);
nor U5769 (N_5769,N_4947,N_4836);
and U5770 (N_5770,N_4102,N_4054);
or U5771 (N_5771,N_4231,N_4994);
xnor U5772 (N_5772,N_4636,N_4352);
xnor U5773 (N_5773,N_4556,N_4061);
nor U5774 (N_5774,N_4212,N_4301);
nor U5775 (N_5775,N_4352,N_4668);
xor U5776 (N_5776,N_4478,N_4894);
and U5777 (N_5777,N_4648,N_4428);
or U5778 (N_5778,N_4485,N_4392);
nand U5779 (N_5779,N_4036,N_4561);
nor U5780 (N_5780,N_4300,N_4246);
and U5781 (N_5781,N_4671,N_4117);
or U5782 (N_5782,N_4337,N_4526);
xnor U5783 (N_5783,N_4672,N_4701);
and U5784 (N_5784,N_4842,N_4193);
xor U5785 (N_5785,N_4481,N_4779);
and U5786 (N_5786,N_4900,N_4864);
nor U5787 (N_5787,N_4413,N_4323);
or U5788 (N_5788,N_4842,N_4755);
or U5789 (N_5789,N_4853,N_4124);
nand U5790 (N_5790,N_4715,N_4446);
nand U5791 (N_5791,N_4719,N_4283);
nand U5792 (N_5792,N_4422,N_4859);
and U5793 (N_5793,N_4708,N_4350);
nand U5794 (N_5794,N_4925,N_4989);
xor U5795 (N_5795,N_4002,N_4055);
or U5796 (N_5796,N_4774,N_4395);
nand U5797 (N_5797,N_4575,N_4145);
and U5798 (N_5798,N_4759,N_4152);
nand U5799 (N_5799,N_4162,N_4203);
nand U5800 (N_5800,N_4531,N_4494);
and U5801 (N_5801,N_4668,N_4113);
xnor U5802 (N_5802,N_4769,N_4891);
and U5803 (N_5803,N_4075,N_4778);
or U5804 (N_5804,N_4711,N_4875);
nand U5805 (N_5805,N_4274,N_4898);
nor U5806 (N_5806,N_4895,N_4650);
nor U5807 (N_5807,N_4223,N_4975);
nor U5808 (N_5808,N_4174,N_4596);
nand U5809 (N_5809,N_4083,N_4516);
nor U5810 (N_5810,N_4966,N_4916);
nor U5811 (N_5811,N_4772,N_4604);
and U5812 (N_5812,N_4975,N_4057);
nand U5813 (N_5813,N_4681,N_4485);
or U5814 (N_5814,N_4914,N_4093);
nor U5815 (N_5815,N_4251,N_4921);
xor U5816 (N_5816,N_4040,N_4861);
xor U5817 (N_5817,N_4532,N_4060);
nand U5818 (N_5818,N_4796,N_4415);
or U5819 (N_5819,N_4902,N_4412);
nor U5820 (N_5820,N_4790,N_4561);
and U5821 (N_5821,N_4843,N_4037);
or U5822 (N_5822,N_4866,N_4267);
and U5823 (N_5823,N_4685,N_4553);
xnor U5824 (N_5824,N_4799,N_4877);
and U5825 (N_5825,N_4805,N_4164);
xnor U5826 (N_5826,N_4090,N_4825);
nand U5827 (N_5827,N_4407,N_4527);
nand U5828 (N_5828,N_4001,N_4974);
nor U5829 (N_5829,N_4475,N_4969);
or U5830 (N_5830,N_4506,N_4592);
xor U5831 (N_5831,N_4019,N_4552);
xnor U5832 (N_5832,N_4536,N_4745);
nor U5833 (N_5833,N_4377,N_4538);
and U5834 (N_5834,N_4724,N_4075);
and U5835 (N_5835,N_4010,N_4204);
and U5836 (N_5836,N_4618,N_4002);
or U5837 (N_5837,N_4219,N_4577);
nand U5838 (N_5838,N_4242,N_4435);
xor U5839 (N_5839,N_4672,N_4381);
and U5840 (N_5840,N_4217,N_4892);
nor U5841 (N_5841,N_4780,N_4163);
nand U5842 (N_5842,N_4339,N_4847);
nor U5843 (N_5843,N_4793,N_4521);
or U5844 (N_5844,N_4704,N_4766);
and U5845 (N_5845,N_4695,N_4785);
or U5846 (N_5846,N_4842,N_4108);
nand U5847 (N_5847,N_4049,N_4391);
nor U5848 (N_5848,N_4630,N_4959);
nor U5849 (N_5849,N_4647,N_4531);
nand U5850 (N_5850,N_4074,N_4815);
nand U5851 (N_5851,N_4761,N_4966);
and U5852 (N_5852,N_4656,N_4312);
and U5853 (N_5853,N_4450,N_4624);
nor U5854 (N_5854,N_4025,N_4838);
xor U5855 (N_5855,N_4602,N_4170);
xnor U5856 (N_5856,N_4858,N_4367);
nand U5857 (N_5857,N_4916,N_4792);
nand U5858 (N_5858,N_4734,N_4051);
and U5859 (N_5859,N_4563,N_4334);
nor U5860 (N_5860,N_4066,N_4367);
xnor U5861 (N_5861,N_4140,N_4273);
or U5862 (N_5862,N_4958,N_4915);
and U5863 (N_5863,N_4094,N_4046);
or U5864 (N_5864,N_4606,N_4345);
nand U5865 (N_5865,N_4914,N_4456);
nand U5866 (N_5866,N_4810,N_4292);
nand U5867 (N_5867,N_4782,N_4592);
and U5868 (N_5868,N_4455,N_4720);
nor U5869 (N_5869,N_4308,N_4456);
and U5870 (N_5870,N_4451,N_4701);
or U5871 (N_5871,N_4002,N_4389);
or U5872 (N_5872,N_4960,N_4657);
and U5873 (N_5873,N_4109,N_4106);
or U5874 (N_5874,N_4648,N_4792);
or U5875 (N_5875,N_4364,N_4039);
xnor U5876 (N_5876,N_4922,N_4789);
or U5877 (N_5877,N_4469,N_4846);
and U5878 (N_5878,N_4609,N_4647);
nand U5879 (N_5879,N_4311,N_4340);
nor U5880 (N_5880,N_4877,N_4615);
xnor U5881 (N_5881,N_4052,N_4451);
xor U5882 (N_5882,N_4933,N_4529);
nor U5883 (N_5883,N_4446,N_4855);
nand U5884 (N_5884,N_4833,N_4486);
nand U5885 (N_5885,N_4172,N_4777);
or U5886 (N_5886,N_4257,N_4361);
nor U5887 (N_5887,N_4786,N_4893);
nand U5888 (N_5888,N_4884,N_4192);
nand U5889 (N_5889,N_4437,N_4034);
nor U5890 (N_5890,N_4844,N_4528);
nand U5891 (N_5891,N_4154,N_4647);
or U5892 (N_5892,N_4359,N_4843);
or U5893 (N_5893,N_4152,N_4830);
nor U5894 (N_5894,N_4264,N_4159);
nor U5895 (N_5895,N_4979,N_4267);
or U5896 (N_5896,N_4419,N_4553);
xnor U5897 (N_5897,N_4540,N_4378);
or U5898 (N_5898,N_4750,N_4368);
or U5899 (N_5899,N_4887,N_4607);
nand U5900 (N_5900,N_4769,N_4732);
xnor U5901 (N_5901,N_4418,N_4747);
or U5902 (N_5902,N_4948,N_4154);
or U5903 (N_5903,N_4407,N_4739);
and U5904 (N_5904,N_4001,N_4214);
or U5905 (N_5905,N_4681,N_4882);
or U5906 (N_5906,N_4281,N_4373);
nor U5907 (N_5907,N_4709,N_4858);
xnor U5908 (N_5908,N_4028,N_4319);
or U5909 (N_5909,N_4844,N_4356);
or U5910 (N_5910,N_4710,N_4564);
or U5911 (N_5911,N_4450,N_4741);
and U5912 (N_5912,N_4114,N_4538);
and U5913 (N_5913,N_4239,N_4734);
or U5914 (N_5914,N_4469,N_4524);
or U5915 (N_5915,N_4109,N_4501);
nor U5916 (N_5916,N_4896,N_4883);
xnor U5917 (N_5917,N_4532,N_4150);
and U5918 (N_5918,N_4180,N_4749);
xor U5919 (N_5919,N_4654,N_4764);
or U5920 (N_5920,N_4931,N_4851);
xor U5921 (N_5921,N_4852,N_4433);
and U5922 (N_5922,N_4304,N_4970);
nor U5923 (N_5923,N_4558,N_4744);
or U5924 (N_5924,N_4371,N_4207);
xnor U5925 (N_5925,N_4067,N_4511);
and U5926 (N_5926,N_4650,N_4946);
xor U5927 (N_5927,N_4199,N_4645);
nor U5928 (N_5928,N_4017,N_4750);
nand U5929 (N_5929,N_4525,N_4416);
or U5930 (N_5930,N_4250,N_4771);
xnor U5931 (N_5931,N_4626,N_4246);
xnor U5932 (N_5932,N_4255,N_4230);
nor U5933 (N_5933,N_4946,N_4671);
and U5934 (N_5934,N_4621,N_4751);
xnor U5935 (N_5935,N_4227,N_4848);
nand U5936 (N_5936,N_4135,N_4788);
nor U5937 (N_5937,N_4255,N_4492);
nand U5938 (N_5938,N_4288,N_4183);
and U5939 (N_5939,N_4018,N_4740);
nor U5940 (N_5940,N_4864,N_4870);
nand U5941 (N_5941,N_4557,N_4081);
nor U5942 (N_5942,N_4069,N_4928);
and U5943 (N_5943,N_4855,N_4526);
and U5944 (N_5944,N_4081,N_4436);
or U5945 (N_5945,N_4773,N_4802);
and U5946 (N_5946,N_4511,N_4766);
and U5947 (N_5947,N_4612,N_4962);
and U5948 (N_5948,N_4777,N_4069);
and U5949 (N_5949,N_4918,N_4044);
and U5950 (N_5950,N_4253,N_4395);
nand U5951 (N_5951,N_4252,N_4956);
nand U5952 (N_5952,N_4837,N_4172);
nand U5953 (N_5953,N_4973,N_4962);
and U5954 (N_5954,N_4188,N_4412);
and U5955 (N_5955,N_4677,N_4892);
and U5956 (N_5956,N_4458,N_4476);
xor U5957 (N_5957,N_4764,N_4434);
xor U5958 (N_5958,N_4626,N_4231);
xor U5959 (N_5959,N_4316,N_4534);
nand U5960 (N_5960,N_4367,N_4592);
nand U5961 (N_5961,N_4234,N_4375);
nor U5962 (N_5962,N_4951,N_4708);
nand U5963 (N_5963,N_4696,N_4362);
nand U5964 (N_5964,N_4747,N_4028);
xor U5965 (N_5965,N_4082,N_4518);
or U5966 (N_5966,N_4345,N_4330);
nand U5967 (N_5967,N_4854,N_4499);
xnor U5968 (N_5968,N_4855,N_4381);
and U5969 (N_5969,N_4561,N_4147);
and U5970 (N_5970,N_4856,N_4309);
xnor U5971 (N_5971,N_4362,N_4174);
xnor U5972 (N_5972,N_4443,N_4242);
nor U5973 (N_5973,N_4108,N_4629);
or U5974 (N_5974,N_4079,N_4988);
nor U5975 (N_5975,N_4943,N_4379);
nor U5976 (N_5976,N_4011,N_4776);
and U5977 (N_5977,N_4412,N_4096);
nand U5978 (N_5978,N_4823,N_4654);
xor U5979 (N_5979,N_4784,N_4155);
nor U5980 (N_5980,N_4864,N_4040);
or U5981 (N_5981,N_4004,N_4351);
nor U5982 (N_5982,N_4273,N_4051);
or U5983 (N_5983,N_4399,N_4333);
nor U5984 (N_5984,N_4684,N_4984);
or U5985 (N_5985,N_4578,N_4402);
nor U5986 (N_5986,N_4355,N_4867);
nor U5987 (N_5987,N_4033,N_4475);
or U5988 (N_5988,N_4611,N_4191);
nand U5989 (N_5989,N_4160,N_4256);
nor U5990 (N_5990,N_4356,N_4422);
or U5991 (N_5991,N_4590,N_4954);
xnor U5992 (N_5992,N_4406,N_4056);
xnor U5993 (N_5993,N_4829,N_4047);
or U5994 (N_5994,N_4834,N_4488);
xor U5995 (N_5995,N_4365,N_4201);
or U5996 (N_5996,N_4027,N_4311);
nor U5997 (N_5997,N_4731,N_4250);
nor U5998 (N_5998,N_4035,N_4799);
or U5999 (N_5999,N_4209,N_4856);
and U6000 (N_6000,N_5275,N_5938);
nand U6001 (N_6001,N_5406,N_5887);
nand U6002 (N_6002,N_5774,N_5555);
and U6003 (N_6003,N_5423,N_5797);
nand U6004 (N_6004,N_5223,N_5944);
and U6005 (N_6005,N_5332,N_5409);
nor U6006 (N_6006,N_5230,N_5486);
or U6007 (N_6007,N_5759,N_5351);
nand U6008 (N_6008,N_5478,N_5549);
or U6009 (N_6009,N_5343,N_5510);
xor U6010 (N_6010,N_5123,N_5009);
or U6011 (N_6011,N_5190,N_5043);
nor U6012 (N_6012,N_5619,N_5579);
nor U6013 (N_6013,N_5213,N_5861);
nor U6014 (N_6014,N_5138,N_5808);
nor U6015 (N_6015,N_5833,N_5756);
and U6016 (N_6016,N_5411,N_5207);
or U6017 (N_6017,N_5604,N_5001);
nand U6018 (N_6018,N_5441,N_5254);
nand U6019 (N_6019,N_5057,N_5241);
or U6020 (N_6020,N_5841,N_5975);
nor U6021 (N_6021,N_5313,N_5595);
nor U6022 (N_6022,N_5116,N_5176);
and U6023 (N_6023,N_5139,N_5189);
and U6024 (N_6024,N_5066,N_5939);
and U6025 (N_6025,N_5769,N_5038);
nand U6026 (N_6026,N_5713,N_5762);
xor U6027 (N_6027,N_5840,N_5319);
nand U6028 (N_6028,N_5484,N_5090);
nand U6029 (N_6029,N_5210,N_5581);
and U6030 (N_6030,N_5469,N_5903);
and U6031 (N_6031,N_5105,N_5069);
nand U6032 (N_6032,N_5894,N_5671);
and U6033 (N_6033,N_5747,N_5187);
xnor U6034 (N_6034,N_5659,N_5128);
and U6035 (N_6035,N_5592,N_5528);
nand U6036 (N_6036,N_5442,N_5740);
nand U6037 (N_6037,N_5174,N_5432);
nor U6038 (N_6038,N_5450,N_5687);
nor U6039 (N_6039,N_5382,N_5111);
nor U6040 (N_6040,N_5267,N_5807);
and U6041 (N_6041,N_5929,N_5225);
xnor U6042 (N_6042,N_5074,N_5056);
xor U6043 (N_6043,N_5353,N_5739);
nand U6044 (N_6044,N_5614,N_5996);
or U6045 (N_6045,N_5674,N_5192);
and U6046 (N_6046,N_5723,N_5476);
or U6047 (N_6047,N_5422,N_5133);
or U6048 (N_6048,N_5414,N_5886);
nor U6049 (N_6049,N_5503,N_5053);
xor U6050 (N_6050,N_5271,N_5520);
and U6051 (N_6051,N_5742,N_5599);
or U6052 (N_6052,N_5789,N_5600);
nor U6053 (N_6053,N_5358,N_5475);
xnor U6054 (N_6054,N_5732,N_5295);
nor U6055 (N_6055,N_5185,N_5553);
xnor U6056 (N_6056,N_5735,N_5309);
nor U6057 (N_6057,N_5670,N_5901);
nor U6058 (N_6058,N_5270,N_5218);
nor U6059 (N_6059,N_5052,N_5626);
nor U6060 (N_6060,N_5635,N_5629);
nand U6061 (N_6061,N_5193,N_5183);
nand U6062 (N_6062,N_5997,N_5691);
and U6063 (N_6063,N_5646,N_5080);
nor U6064 (N_6064,N_5155,N_5858);
or U6065 (N_6065,N_5695,N_5203);
or U6066 (N_6066,N_5948,N_5709);
and U6067 (N_6067,N_5387,N_5489);
nor U6068 (N_6068,N_5471,N_5787);
or U6069 (N_6069,N_5796,N_5765);
xor U6070 (N_6070,N_5530,N_5383);
or U6071 (N_6071,N_5424,N_5950);
and U6072 (N_6072,N_5034,N_5263);
or U6073 (N_6073,N_5005,N_5608);
xor U6074 (N_6074,N_5127,N_5630);
nor U6075 (N_6075,N_5633,N_5289);
nand U6076 (N_6076,N_5611,N_5966);
nor U6077 (N_6077,N_5726,N_5542);
nor U6078 (N_6078,N_5303,N_5181);
or U6079 (N_6079,N_5785,N_5577);
nor U6080 (N_6080,N_5438,N_5362);
nor U6081 (N_6081,N_5783,N_5779);
nor U6082 (N_6082,N_5474,N_5638);
xor U6083 (N_6083,N_5851,N_5011);
or U6084 (N_6084,N_5985,N_5433);
and U6085 (N_6085,N_5167,N_5013);
nand U6086 (N_6086,N_5763,N_5410);
xnor U6087 (N_6087,N_5959,N_5045);
nand U6088 (N_6088,N_5463,N_5338);
and U6089 (N_6089,N_5597,N_5136);
nor U6090 (N_6090,N_5810,N_5019);
nor U6091 (N_6091,N_5559,N_5087);
or U6092 (N_6092,N_5465,N_5141);
nor U6093 (N_6093,N_5628,N_5491);
and U6094 (N_6094,N_5046,N_5100);
and U6095 (N_6095,N_5784,N_5169);
nor U6096 (N_6096,N_5692,N_5017);
xnor U6097 (N_6097,N_5305,N_5191);
nor U6098 (N_6098,N_5716,N_5262);
nand U6099 (N_6099,N_5316,N_5989);
xor U6100 (N_6100,N_5277,N_5285);
nor U6101 (N_6101,N_5690,N_5067);
xnor U6102 (N_6102,N_5173,N_5748);
nand U6103 (N_6103,N_5341,N_5664);
xnor U6104 (N_6104,N_5242,N_5964);
or U6105 (N_6105,N_5357,N_5472);
nor U6106 (N_6106,N_5668,N_5879);
and U6107 (N_6107,N_5533,N_5444);
and U6108 (N_6108,N_5591,N_5637);
and U6109 (N_6109,N_5085,N_5578);
xor U6110 (N_6110,N_5803,N_5776);
xor U6111 (N_6111,N_5854,N_5728);
xor U6112 (N_6112,N_5867,N_5391);
nor U6113 (N_6113,N_5522,N_5312);
nor U6114 (N_6114,N_5026,N_5655);
nor U6115 (N_6115,N_5897,N_5296);
nor U6116 (N_6116,N_5331,N_5673);
or U6117 (N_6117,N_5935,N_5392);
nor U6118 (N_6118,N_5027,N_5434);
nor U6119 (N_6119,N_5495,N_5068);
or U6120 (N_6120,N_5758,N_5795);
xor U6121 (N_6121,N_5064,N_5605);
nor U6122 (N_6122,N_5073,N_5171);
xor U6123 (N_6123,N_5425,N_5805);
nand U6124 (N_6124,N_5575,N_5298);
nor U6125 (N_6125,N_5482,N_5968);
nand U6126 (N_6126,N_5365,N_5330);
and U6127 (N_6127,N_5071,N_5681);
xor U6128 (N_6128,N_5396,N_5719);
and U6129 (N_6129,N_5117,N_5221);
and U6130 (N_6130,N_5812,N_5310);
nand U6131 (N_6131,N_5282,N_5957);
nand U6132 (N_6132,N_5609,N_5910);
xor U6133 (N_6133,N_5145,N_5751);
or U6134 (N_6134,N_5946,N_5616);
or U6135 (N_6135,N_5273,N_5895);
nand U6136 (N_6136,N_5443,N_5012);
and U6137 (N_6137,N_5268,N_5024);
and U6138 (N_6138,N_5738,N_5744);
nor U6139 (N_6139,N_5834,N_5882);
nand U6140 (N_6140,N_5694,N_5698);
nand U6141 (N_6141,N_5767,N_5921);
xor U6142 (N_6142,N_5823,N_5844);
xnor U6143 (N_6143,N_5857,N_5827);
nand U6144 (N_6144,N_5016,N_5217);
nand U6145 (N_6145,N_5650,N_5845);
and U6146 (N_6146,N_5048,N_5594);
xnor U6147 (N_6147,N_5927,N_5590);
or U6148 (N_6148,N_5216,N_5567);
xor U6149 (N_6149,N_5194,N_5872);
xnor U6150 (N_6150,N_5371,N_5906);
xnor U6151 (N_6151,N_5545,N_5318);
nand U6152 (N_6152,N_5459,N_5710);
nand U6153 (N_6153,N_5771,N_5822);
nand U6154 (N_6154,N_5551,N_5729);
and U6155 (N_6155,N_5023,N_5222);
and U6156 (N_6156,N_5515,N_5849);
xnor U6157 (N_6157,N_5666,N_5736);
nor U6158 (N_6158,N_5370,N_5924);
nor U6159 (N_6159,N_5306,N_5919);
nor U6160 (N_6160,N_5086,N_5920);
nor U6161 (N_6161,N_5003,N_5202);
xor U6162 (N_6162,N_5519,N_5021);
xor U6163 (N_6163,N_5773,N_5279);
xnor U6164 (N_6164,N_5250,N_5287);
xnor U6165 (N_6165,N_5419,N_5790);
or U6166 (N_6166,N_5407,N_5539);
nand U6167 (N_6167,N_5696,N_5714);
nand U6168 (N_6168,N_5177,N_5570);
or U6169 (N_6169,N_5302,N_5106);
or U6170 (N_6170,N_5199,N_5004);
or U6171 (N_6171,N_5725,N_5516);
nand U6172 (N_6172,N_5248,N_5580);
and U6173 (N_6173,N_5607,N_5794);
or U6174 (N_6174,N_5513,N_5163);
nand U6175 (N_6175,N_5757,N_5084);
or U6176 (N_6176,N_5993,N_5799);
nor U6177 (N_6177,N_5431,N_5317);
nor U6178 (N_6178,N_5109,N_5777);
nand U6179 (N_6179,N_5811,N_5603);
and U6180 (N_6180,N_5446,N_5269);
nor U6181 (N_6181,N_5963,N_5283);
and U6182 (N_6182,N_5126,N_5715);
and U6183 (N_6183,N_5307,N_5627);
or U6184 (N_6184,N_5704,N_5556);
or U6185 (N_6185,N_5639,N_5914);
xor U6186 (N_6186,N_5737,N_5037);
or U6187 (N_6187,N_5240,N_5505);
xnor U6188 (N_6188,N_5149,N_5439);
xnor U6189 (N_6189,N_5654,N_5980);
nand U6190 (N_6190,N_5504,N_5473);
nor U6191 (N_6191,N_5701,N_5036);
xor U6192 (N_6192,N_5855,N_5507);
and U6193 (N_6193,N_5228,N_5909);
and U6194 (N_6194,N_5239,N_5206);
nor U6195 (N_6195,N_5874,N_5417);
nand U6196 (N_6196,N_5684,N_5148);
and U6197 (N_6197,N_5727,N_5569);
and U6198 (N_6198,N_5699,N_5247);
and U6199 (N_6199,N_5294,N_5832);
or U6200 (N_6200,N_5554,N_5214);
and U6201 (N_6201,N_5863,N_5481);
xnor U6202 (N_6202,N_5824,N_5333);
xnor U6203 (N_6203,N_5913,N_5464);
and U6204 (N_6204,N_5081,N_5132);
xor U6205 (N_6205,N_5766,N_5689);
and U6206 (N_6206,N_5429,N_5025);
and U6207 (N_6207,N_5121,N_5791);
or U6208 (N_6208,N_5120,N_5376);
xor U6209 (N_6209,N_5381,N_5224);
xnor U6210 (N_6210,N_5186,N_5538);
or U6211 (N_6211,N_5180,N_5000);
or U6212 (N_6212,N_5678,N_5140);
nand U6213 (N_6213,N_5661,N_5261);
nor U6214 (N_6214,N_5449,N_5028);
or U6215 (N_6215,N_5506,N_5398);
and U6216 (N_6216,N_5793,N_5647);
or U6217 (N_6217,N_5359,N_5992);
and U6218 (N_6218,N_5293,N_5781);
xnor U6219 (N_6219,N_5236,N_5426);
nand U6220 (N_6220,N_5511,N_5488);
nor U6221 (N_6221,N_5831,N_5253);
or U6222 (N_6222,N_5550,N_5995);
xor U6223 (N_6223,N_5030,N_5676);
nor U6224 (N_6224,N_5458,N_5150);
and U6225 (N_6225,N_5462,N_5500);
xnor U6226 (N_6226,N_5092,N_5361);
and U6227 (N_6227,N_5792,N_5020);
or U6228 (N_6228,N_5998,N_5601);
xnor U6229 (N_6229,N_5386,N_5044);
or U6230 (N_6230,N_5420,N_5178);
or U6231 (N_6231,N_5900,N_5645);
nand U6232 (N_6232,N_5705,N_5196);
xnor U6233 (N_6233,N_5750,N_5820);
xor U6234 (N_6234,N_5154,N_5587);
xor U6235 (N_6235,N_5256,N_5683);
or U6236 (N_6236,N_5006,N_5397);
or U6237 (N_6237,N_5299,N_5546);
xor U6238 (N_6238,N_5088,N_5072);
nand U6239 (N_6239,N_5168,N_5898);
nor U6240 (N_6240,N_5007,N_5922);
xor U6241 (N_6241,N_5839,N_5470);
or U6242 (N_6242,N_5369,N_5984);
or U6243 (N_6243,N_5537,N_5165);
nor U6244 (N_6244,N_5987,N_5435);
xor U6245 (N_6245,N_5399,N_5226);
nand U6246 (N_6246,N_5943,N_5238);
xor U6247 (N_6247,N_5098,N_5347);
nand U6248 (N_6248,N_5663,N_5350);
xor U6249 (N_6249,N_5721,N_5846);
and U6250 (N_6250,N_5636,N_5852);
xnor U6251 (N_6251,N_5548,N_5652);
nor U6252 (N_6252,N_5314,N_5368);
or U6253 (N_6253,N_5942,N_5972);
nor U6254 (N_6254,N_5091,N_5304);
xor U6255 (N_6255,N_5348,N_5063);
nand U6256 (N_6256,N_5364,N_5493);
and U6257 (N_6257,N_5170,N_5974);
nand U6258 (N_6258,N_5525,N_5480);
and U6259 (N_6259,N_5926,N_5461);
or U6260 (N_6260,N_5682,N_5835);
nor U6261 (N_6261,N_5014,N_5119);
and U6262 (N_6262,N_5818,N_5868);
or U6263 (N_6263,N_5746,N_5393);
and U6264 (N_6264,N_5385,N_5741);
or U6265 (N_6265,N_5932,N_5990);
and U6266 (N_6266,N_5448,N_5408);
and U6267 (N_6267,N_5363,N_5819);
xnor U6268 (N_6268,N_5643,N_5514);
or U6269 (N_6269,N_5962,N_5770);
xor U6270 (N_6270,N_5552,N_5029);
nand U6271 (N_6271,N_5346,N_5826);
and U6272 (N_6272,N_5568,N_5002);
or U6273 (N_6273,N_5866,N_5981);
nand U6274 (N_6274,N_5617,N_5355);
or U6275 (N_6275,N_5281,N_5908);
nand U6276 (N_6276,N_5143,N_5405);
or U6277 (N_6277,N_5232,N_5437);
and U6278 (N_6278,N_5147,N_5829);
nand U6279 (N_6279,N_5099,N_5184);
xnor U6280 (N_6280,N_5838,N_5097);
nor U6281 (N_6281,N_5669,N_5032);
or U6282 (N_6282,N_5915,N_5907);
nor U6283 (N_6283,N_5227,N_5517);
xnor U6284 (N_6284,N_5323,N_5440);
nand U6285 (N_6285,N_5130,N_5875);
or U6286 (N_6286,N_5334,N_5274);
xnor U6287 (N_6287,N_5830,N_5457);
xor U6288 (N_6288,N_5817,N_5697);
nand U6289 (N_6289,N_5082,N_5156);
xnor U6290 (N_6290,N_5413,N_5060);
nand U6291 (N_6291,N_5717,N_5893);
nor U6292 (N_6292,N_5320,N_5802);
nor U6293 (N_6293,N_5544,N_5576);
xor U6294 (N_6294,N_5675,N_5753);
nor U6295 (N_6295,N_5585,N_5561);
nand U6296 (N_6296,N_5342,N_5152);
nor U6297 (N_6297,N_5394,N_5453);
xnor U6298 (N_6298,N_5535,N_5615);
xor U6299 (N_6299,N_5094,N_5649);
nor U6300 (N_6300,N_5496,N_5912);
nor U6301 (N_6301,N_5752,N_5885);
nor U6302 (N_6302,N_5973,N_5598);
or U6303 (N_6303,N_5102,N_5541);
or U6304 (N_6304,N_5547,N_5315);
and U6305 (N_6305,N_5384,N_5284);
or U6306 (N_6306,N_5718,N_5108);
xor U6307 (N_6307,N_5380,N_5917);
nand U6308 (N_6308,N_5521,N_5436);
xnor U6309 (N_6309,N_5953,N_5878);
nor U6310 (N_6310,N_5814,N_5809);
xor U6311 (N_6311,N_5456,N_5110);
xnor U6312 (N_6312,N_5161,N_5499);
nand U6313 (N_6313,N_5200,N_5883);
nand U6314 (N_6314,N_5237,N_5960);
or U6315 (N_6315,N_5404,N_5050);
nand U6316 (N_6316,N_5234,N_5204);
xor U6317 (N_6317,N_5703,N_5911);
nor U6318 (N_6318,N_5562,N_5452);
xnor U6319 (N_6319,N_5114,N_5502);
xnor U6320 (N_6320,N_5103,N_5772);
and U6321 (N_6321,N_5951,N_5083);
nor U6322 (N_6322,N_5129,N_5859);
and U6323 (N_6323,N_5640,N_5388);
or U6324 (N_6324,N_5850,N_5686);
or U6325 (N_6325,N_5272,N_5212);
and U6326 (N_6326,N_5853,N_5916);
and U6327 (N_6327,N_5712,N_5930);
and U6328 (N_6328,N_5079,N_5815);
xor U6329 (N_6329,N_5527,N_5118);
nor U6330 (N_6330,N_5335,N_5460);
or U6331 (N_6331,N_5033,N_5800);
nor U6332 (N_6332,N_5492,N_5573);
and U6333 (N_6333,N_5049,N_5625);
or U6334 (N_6334,N_5497,N_5925);
and U6335 (N_6335,N_5430,N_5821);
nor U6336 (N_6336,N_5390,N_5326);
nor U6337 (N_6337,N_5612,N_5494);
and U6338 (N_6338,N_5888,N_5172);
nand U6339 (N_6339,N_5624,N_5656);
xor U6340 (N_6340,N_5198,N_5146);
nor U6341 (N_6341,N_5375,N_5095);
nand U6342 (N_6342,N_5941,N_5124);
nand U6343 (N_6343,N_5586,N_5706);
and U6344 (N_6344,N_5078,N_5300);
and U6345 (N_6345,N_5836,N_5377);
nor U6346 (N_6346,N_5509,N_5427);
nor U6347 (N_6347,N_5104,N_5125);
or U6348 (N_6348,N_5367,N_5018);
nor U6349 (N_6349,N_5558,N_5672);
and U6350 (N_6350,N_5899,N_5339);
nand U6351 (N_6351,N_5632,N_5047);
nand U6352 (N_6352,N_5379,N_5374);
nand U6353 (N_6353,N_5142,N_5955);
nor U6354 (N_6354,N_5122,N_5040);
nor U6355 (N_6355,N_5428,N_5041);
and U6356 (N_6356,N_5743,N_5531);
and U6357 (N_6357,N_5644,N_5257);
or U6358 (N_6358,N_5720,N_5991);
nor U6359 (N_6359,N_5035,N_5731);
and U6360 (N_6360,N_5389,N_5584);
and U6361 (N_6361,N_5215,N_5965);
xnor U6362 (N_6362,N_5988,N_5162);
and U6363 (N_6363,N_5837,N_5702);
nor U6364 (N_6364,N_5523,N_5113);
or U6365 (N_6365,N_5373,N_5610);
nand U6366 (N_6366,N_5862,N_5869);
and U6367 (N_6367,N_5015,N_5418);
nor U6368 (N_6368,N_5487,N_5233);
xnor U6369 (N_6369,N_5976,N_5954);
xnor U6370 (N_6370,N_5328,N_5058);
xnor U6371 (N_6371,N_5804,N_5144);
nor U6372 (N_6372,N_5896,N_5498);
nor U6373 (N_6373,N_5970,N_5151);
nand U6374 (N_6374,N_5977,N_5101);
nand U6375 (N_6375,N_5501,N_5708);
or U6376 (N_6376,N_5153,N_5665);
xnor U6377 (N_6377,N_5865,N_5244);
or U6378 (N_6378,N_5873,N_5182);
nand U6379 (N_6379,N_5297,N_5246);
nor U6380 (N_6380,N_5402,N_5884);
and U6381 (N_6381,N_5164,N_5479);
nor U6382 (N_6382,N_5768,N_5813);
nand U6383 (N_6383,N_5602,N_5096);
or U6384 (N_6384,N_5593,N_5971);
nor U6385 (N_6385,N_5280,N_5707);
nor U6386 (N_6386,N_5401,N_5679);
nand U6387 (N_6387,N_5843,N_5540);
or U6388 (N_6388,N_5724,N_5291);
nor U6389 (N_6389,N_5572,N_5571);
nor U6390 (N_6390,N_5642,N_5828);
nand U6391 (N_6391,N_5249,N_5219);
or U6392 (N_6392,N_5158,N_5524);
nor U6393 (N_6393,N_5336,N_5266);
or U6394 (N_6394,N_5220,N_5994);
or U6395 (N_6395,N_5734,N_5089);
and U6396 (N_6396,N_5890,N_5565);
or U6397 (N_6397,N_5065,N_5512);
xor U6398 (N_6398,N_5157,N_5445);
and U6399 (N_6399,N_5325,N_5574);
nand U6400 (N_6400,N_5354,N_5889);
nand U6401 (N_6401,N_5931,N_5983);
or U6402 (N_6402,N_5560,N_5596);
nor U6403 (N_6403,N_5589,N_5211);
nor U6404 (N_6404,N_5508,N_5201);
or U6405 (N_6405,N_5039,N_5945);
xor U6406 (N_6406,N_5543,N_5321);
or U6407 (N_6407,N_5657,N_5412);
nand U6408 (N_6408,N_5563,N_5786);
nand U6409 (N_6409,N_5308,N_5483);
nand U6410 (N_6410,N_5477,N_5135);
or U6411 (N_6411,N_5245,N_5947);
and U6412 (N_6412,N_5641,N_5286);
or U6413 (N_6413,N_5008,N_5967);
or U6414 (N_6414,N_5864,N_5159);
nand U6415 (N_6415,N_5564,N_5311);
xor U6416 (N_6416,N_5243,N_5276);
nor U6417 (N_6417,N_5688,N_5265);
and U6418 (N_6418,N_5952,N_5490);
nor U6419 (N_6419,N_5229,N_5112);
nor U6420 (N_6420,N_5755,N_5749);
nand U6421 (N_6421,N_5902,N_5252);
xor U6422 (N_6422,N_5798,N_5062);
nand U6423 (N_6423,N_5958,N_5179);
xor U6424 (N_6424,N_5621,N_5877);
and U6425 (N_6425,N_5344,N_5761);
and U6426 (N_6426,N_5940,N_5251);
nand U6427 (N_6427,N_5891,N_5415);
nand U6428 (N_6428,N_5054,N_5662);
nand U6429 (N_6429,N_5529,N_5764);
and U6430 (N_6430,N_5107,N_5288);
nor U6431 (N_6431,N_5061,N_5454);
nand U6432 (N_6432,N_5806,N_5447);
and U6433 (N_6433,N_5195,N_5778);
xor U6434 (N_6434,N_5395,N_5631);
nand U6435 (N_6435,N_5292,N_5918);
xor U6436 (N_6436,N_5451,N_5648);
or U6437 (N_6437,N_5131,N_5949);
and U6438 (N_6438,N_5733,N_5816);
and U6439 (N_6439,N_5301,N_5622);
xnor U6440 (N_6440,N_5711,N_5278);
or U6441 (N_6441,N_5936,N_5680);
nor U6442 (N_6442,N_5860,N_5115);
and U6443 (N_6443,N_5618,N_5322);
or U6444 (N_6444,N_5070,N_5485);
nand U6445 (N_6445,N_5209,N_5259);
and U6446 (N_6446,N_5979,N_5623);
nor U6447 (N_6447,N_5583,N_5923);
or U6448 (N_6448,N_5825,N_5197);
nor U6449 (N_6449,N_5175,N_5934);
nor U6450 (N_6450,N_5356,N_5134);
or U6451 (N_6451,N_5059,N_5534);
nor U6452 (N_6452,N_5848,N_5722);
xnor U6453 (N_6453,N_5468,N_5880);
nor U6454 (N_6454,N_5978,N_5076);
nand U6455 (N_6455,N_5260,N_5235);
or U6456 (N_6456,N_5651,N_5536);
or U6457 (N_6457,N_5775,N_5337);
nand U6458 (N_6458,N_5582,N_5290);
or U6459 (N_6459,N_5327,N_5532);
nor U6460 (N_6460,N_5042,N_5366);
nand U6461 (N_6461,N_5403,N_5982);
xnor U6462 (N_6462,N_5137,N_5905);
xnor U6463 (N_6463,N_5372,N_5208);
xnor U6464 (N_6464,N_5986,N_5634);
xnor U6465 (N_6465,N_5700,N_5466);
and U6466 (N_6466,N_5166,N_5653);
or U6467 (N_6467,N_5258,N_5526);
and U6468 (N_6468,N_5400,N_5876);
nor U6469 (N_6469,N_5416,N_5255);
xnor U6470 (N_6470,N_5455,N_5928);
or U6471 (N_6471,N_5856,N_5231);
nor U6472 (N_6472,N_5360,N_5093);
nor U6473 (N_6473,N_5613,N_5693);
nor U6474 (N_6474,N_5847,N_5349);
xnor U6475 (N_6475,N_5588,N_5933);
nor U6476 (N_6476,N_5022,N_5969);
nand U6477 (N_6477,N_5566,N_5467);
xor U6478 (N_6478,N_5557,N_5324);
xnor U6479 (N_6479,N_5205,N_5730);
and U6480 (N_6480,N_5685,N_5892);
nand U6481 (N_6481,N_5904,N_5345);
or U6482 (N_6482,N_5760,N_5780);
nand U6483 (N_6483,N_5378,N_5160);
nand U6484 (N_6484,N_5956,N_5677);
nor U6485 (N_6485,N_5788,N_5660);
nand U6486 (N_6486,N_5842,N_5518);
nor U6487 (N_6487,N_5937,N_5329);
or U6488 (N_6488,N_5881,N_5620);
nor U6489 (N_6489,N_5188,N_5801);
nor U6490 (N_6490,N_5340,N_5870);
nand U6491 (N_6491,N_5075,N_5010);
and U6492 (N_6492,N_5031,N_5754);
nor U6493 (N_6493,N_5055,N_5658);
xnor U6494 (N_6494,N_5051,N_5961);
or U6495 (N_6495,N_5264,N_5667);
nor U6496 (N_6496,N_5745,N_5352);
or U6497 (N_6497,N_5999,N_5871);
nor U6498 (N_6498,N_5782,N_5077);
nor U6499 (N_6499,N_5421,N_5606);
nand U6500 (N_6500,N_5819,N_5887);
or U6501 (N_6501,N_5679,N_5681);
and U6502 (N_6502,N_5709,N_5034);
or U6503 (N_6503,N_5406,N_5987);
and U6504 (N_6504,N_5067,N_5539);
nand U6505 (N_6505,N_5126,N_5531);
or U6506 (N_6506,N_5607,N_5364);
nor U6507 (N_6507,N_5624,N_5117);
and U6508 (N_6508,N_5445,N_5780);
xor U6509 (N_6509,N_5000,N_5830);
and U6510 (N_6510,N_5725,N_5600);
or U6511 (N_6511,N_5071,N_5689);
nand U6512 (N_6512,N_5319,N_5724);
nor U6513 (N_6513,N_5346,N_5875);
or U6514 (N_6514,N_5498,N_5678);
nor U6515 (N_6515,N_5212,N_5341);
nand U6516 (N_6516,N_5265,N_5906);
and U6517 (N_6517,N_5717,N_5171);
and U6518 (N_6518,N_5150,N_5744);
nor U6519 (N_6519,N_5488,N_5064);
xnor U6520 (N_6520,N_5946,N_5277);
nor U6521 (N_6521,N_5554,N_5627);
or U6522 (N_6522,N_5930,N_5190);
nand U6523 (N_6523,N_5413,N_5307);
or U6524 (N_6524,N_5895,N_5588);
nor U6525 (N_6525,N_5047,N_5236);
xor U6526 (N_6526,N_5565,N_5509);
nand U6527 (N_6527,N_5070,N_5510);
and U6528 (N_6528,N_5126,N_5033);
xnor U6529 (N_6529,N_5947,N_5152);
xor U6530 (N_6530,N_5667,N_5685);
xnor U6531 (N_6531,N_5929,N_5774);
nor U6532 (N_6532,N_5197,N_5923);
and U6533 (N_6533,N_5254,N_5051);
and U6534 (N_6534,N_5138,N_5581);
or U6535 (N_6535,N_5719,N_5187);
and U6536 (N_6536,N_5521,N_5485);
nand U6537 (N_6537,N_5588,N_5605);
xnor U6538 (N_6538,N_5738,N_5284);
nor U6539 (N_6539,N_5905,N_5001);
nand U6540 (N_6540,N_5073,N_5977);
nor U6541 (N_6541,N_5481,N_5026);
nand U6542 (N_6542,N_5862,N_5639);
and U6543 (N_6543,N_5601,N_5040);
nor U6544 (N_6544,N_5424,N_5831);
or U6545 (N_6545,N_5044,N_5600);
xnor U6546 (N_6546,N_5399,N_5849);
or U6547 (N_6547,N_5864,N_5106);
nor U6548 (N_6548,N_5258,N_5586);
xnor U6549 (N_6549,N_5376,N_5569);
xor U6550 (N_6550,N_5837,N_5598);
xor U6551 (N_6551,N_5910,N_5649);
and U6552 (N_6552,N_5931,N_5303);
and U6553 (N_6553,N_5833,N_5656);
or U6554 (N_6554,N_5822,N_5574);
nand U6555 (N_6555,N_5134,N_5530);
xor U6556 (N_6556,N_5427,N_5038);
xnor U6557 (N_6557,N_5573,N_5560);
nor U6558 (N_6558,N_5920,N_5882);
and U6559 (N_6559,N_5787,N_5589);
nand U6560 (N_6560,N_5201,N_5392);
nor U6561 (N_6561,N_5096,N_5323);
or U6562 (N_6562,N_5572,N_5128);
nor U6563 (N_6563,N_5342,N_5871);
nor U6564 (N_6564,N_5419,N_5577);
nand U6565 (N_6565,N_5841,N_5954);
nand U6566 (N_6566,N_5087,N_5286);
or U6567 (N_6567,N_5400,N_5399);
or U6568 (N_6568,N_5383,N_5573);
nand U6569 (N_6569,N_5983,N_5591);
nor U6570 (N_6570,N_5757,N_5963);
or U6571 (N_6571,N_5831,N_5399);
nand U6572 (N_6572,N_5870,N_5457);
nor U6573 (N_6573,N_5399,N_5671);
xnor U6574 (N_6574,N_5198,N_5589);
or U6575 (N_6575,N_5921,N_5074);
and U6576 (N_6576,N_5440,N_5905);
nor U6577 (N_6577,N_5199,N_5119);
nor U6578 (N_6578,N_5176,N_5241);
and U6579 (N_6579,N_5133,N_5345);
or U6580 (N_6580,N_5973,N_5094);
nand U6581 (N_6581,N_5064,N_5839);
nor U6582 (N_6582,N_5991,N_5441);
nor U6583 (N_6583,N_5189,N_5710);
nand U6584 (N_6584,N_5807,N_5463);
or U6585 (N_6585,N_5822,N_5021);
xor U6586 (N_6586,N_5099,N_5537);
xnor U6587 (N_6587,N_5540,N_5381);
xor U6588 (N_6588,N_5628,N_5200);
xor U6589 (N_6589,N_5080,N_5559);
xnor U6590 (N_6590,N_5665,N_5248);
nor U6591 (N_6591,N_5231,N_5285);
xnor U6592 (N_6592,N_5128,N_5799);
nand U6593 (N_6593,N_5097,N_5030);
or U6594 (N_6594,N_5613,N_5352);
nand U6595 (N_6595,N_5889,N_5639);
xor U6596 (N_6596,N_5720,N_5055);
and U6597 (N_6597,N_5550,N_5508);
nand U6598 (N_6598,N_5479,N_5597);
xnor U6599 (N_6599,N_5364,N_5718);
and U6600 (N_6600,N_5006,N_5955);
nor U6601 (N_6601,N_5470,N_5962);
nor U6602 (N_6602,N_5198,N_5546);
xor U6603 (N_6603,N_5282,N_5606);
and U6604 (N_6604,N_5029,N_5763);
nor U6605 (N_6605,N_5069,N_5552);
xor U6606 (N_6606,N_5796,N_5623);
nand U6607 (N_6607,N_5137,N_5084);
nor U6608 (N_6608,N_5080,N_5622);
nand U6609 (N_6609,N_5472,N_5556);
or U6610 (N_6610,N_5599,N_5951);
or U6611 (N_6611,N_5549,N_5098);
xnor U6612 (N_6612,N_5293,N_5867);
xnor U6613 (N_6613,N_5898,N_5397);
xor U6614 (N_6614,N_5280,N_5109);
nand U6615 (N_6615,N_5345,N_5694);
or U6616 (N_6616,N_5357,N_5506);
and U6617 (N_6617,N_5396,N_5684);
and U6618 (N_6618,N_5178,N_5170);
nand U6619 (N_6619,N_5600,N_5790);
xor U6620 (N_6620,N_5056,N_5182);
nand U6621 (N_6621,N_5727,N_5173);
nand U6622 (N_6622,N_5298,N_5700);
nand U6623 (N_6623,N_5015,N_5994);
xor U6624 (N_6624,N_5889,N_5254);
or U6625 (N_6625,N_5818,N_5028);
nor U6626 (N_6626,N_5371,N_5068);
nor U6627 (N_6627,N_5516,N_5189);
nor U6628 (N_6628,N_5496,N_5742);
or U6629 (N_6629,N_5185,N_5746);
nand U6630 (N_6630,N_5868,N_5637);
or U6631 (N_6631,N_5367,N_5277);
nor U6632 (N_6632,N_5129,N_5682);
and U6633 (N_6633,N_5296,N_5486);
nor U6634 (N_6634,N_5127,N_5792);
nand U6635 (N_6635,N_5321,N_5579);
nand U6636 (N_6636,N_5845,N_5177);
nand U6637 (N_6637,N_5801,N_5180);
nor U6638 (N_6638,N_5996,N_5367);
and U6639 (N_6639,N_5314,N_5192);
or U6640 (N_6640,N_5148,N_5481);
nand U6641 (N_6641,N_5640,N_5987);
nor U6642 (N_6642,N_5645,N_5828);
and U6643 (N_6643,N_5867,N_5107);
nand U6644 (N_6644,N_5416,N_5940);
xnor U6645 (N_6645,N_5092,N_5754);
and U6646 (N_6646,N_5491,N_5155);
or U6647 (N_6647,N_5313,N_5242);
nor U6648 (N_6648,N_5236,N_5954);
or U6649 (N_6649,N_5383,N_5072);
nand U6650 (N_6650,N_5806,N_5672);
nor U6651 (N_6651,N_5743,N_5267);
or U6652 (N_6652,N_5090,N_5909);
nand U6653 (N_6653,N_5121,N_5359);
and U6654 (N_6654,N_5592,N_5541);
and U6655 (N_6655,N_5934,N_5379);
xnor U6656 (N_6656,N_5533,N_5742);
nand U6657 (N_6657,N_5098,N_5900);
xor U6658 (N_6658,N_5333,N_5806);
or U6659 (N_6659,N_5027,N_5185);
xnor U6660 (N_6660,N_5474,N_5269);
or U6661 (N_6661,N_5513,N_5458);
nor U6662 (N_6662,N_5445,N_5813);
xor U6663 (N_6663,N_5653,N_5113);
or U6664 (N_6664,N_5283,N_5047);
nor U6665 (N_6665,N_5566,N_5984);
xnor U6666 (N_6666,N_5236,N_5766);
nor U6667 (N_6667,N_5675,N_5748);
xor U6668 (N_6668,N_5916,N_5669);
nor U6669 (N_6669,N_5864,N_5462);
nor U6670 (N_6670,N_5209,N_5548);
xor U6671 (N_6671,N_5049,N_5877);
nor U6672 (N_6672,N_5728,N_5426);
and U6673 (N_6673,N_5619,N_5111);
or U6674 (N_6674,N_5660,N_5314);
and U6675 (N_6675,N_5941,N_5010);
nor U6676 (N_6676,N_5857,N_5586);
xnor U6677 (N_6677,N_5696,N_5296);
xnor U6678 (N_6678,N_5749,N_5629);
nor U6679 (N_6679,N_5795,N_5903);
nand U6680 (N_6680,N_5928,N_5689);
and U6681 (N_6681,N_5025,N_5760);
nor U6682 (N_6682,N_5708,N_5883);
nand U6683 (N_6683,N_5423,N_5027);
and U6684 (N_6684,N_5492,N_5789);
and U6685 (N_6685,N_5808,N_5505);
or U6686 (N_6686,N_5333,N_5007);
or U6687 (N_6687,N_5563,N_5686);
xor U6688 (N_6688,N_5079,N_5319);
xnor U6689 (N_6689,N_5790,N_5769);
nor U6690 (N_6690,N_5637,N_5377);
or U6691 (N_6691,N_5895,N_5133);
nand U6692 (N_6692,N_5881,N_5508);
nor U6693 (N_6693,N_5062,N_5997);
xnor U6694 (N_6694,N_5367,N_5150);
xor U6695 (N_6695,N_5579,N_5357);
nand U6696 (N_6696,N_5163,N_5034);
nor U6697 (N_6697,N_5449,N_5344);
nor U6698 (N_6698,N_5787,N_5153);
nor U6699 (N_6699,N_5056,N_5659);
nand U6700 (N_6700,N_5510,N_5430);
nor U6701 (N_6701,N_5552,N_5043);
xnor U6702 (N_6702,N_5597,N_5156);
xor U6703 (N_6703,N_5445,N_5831);
xnor U6704 (N_6704,N_5089,N_5196);
nor U6705 (N_6705,N_5852,N_5645);
or U6706 (N_6706,N_5710,N_5952);
nand U6707 (N_6707,N_5417,N_5768);
xor U6708 (N_6708,N_5379,N_5659);
and U6709 (N_6709,N_5967,N_5307);
or U6710 (N_6710,N_5978,N_5470);
or U6711 (N_6711,N_5242,N_5226);
and U6712 (N_6712,N_5344,N_5125);
nand U6713 (N_6713,N_5439,N_5690);
and U6714 (N_6714,N_5377,N_5245);
and U6715 (N_6715,N_5966,N_5588);
nand U6716 (N_6716,N_5601,N_5613);
and U6717 (N_6717,N_5115,N_5488);
and U6718 (N_6718,N_5589,N_5926);
nand U6719 (N_6719,N_5078,N_5960);
xor U6720 (N_6720,N_5100,N_5773);
and U6721 (N_6721,N_5881,N_5970);
xor U6722 (N_6722,N_5234,N_5833);
nor U6723 (N_6723,N_5588,N_5436);
xnor U6724 (N_6724,N_5054,N_5454);
xnor U6725 (N_6725,N_5965,N_5908);
and U6726 (N_6726,N_5597,N_5069);
or U6727 (N_6727,N_5810,N_5543);
and U6728 (N_6728,N_5626,N_5327);
xnor U6729 (N_6729,N_5732,N_5027);
nand U6730 (N_6730,N_5364,N_5909);
nand U6731 (N_6731,N_5812,N_5032);
xnor U6732 (N_6732,N_5668,N_5827);
nor U6733 (N_6733,N_5985,N_5351);
and U6734 (N_6734,N_5152,N_5762);
nor U6735 (N_6735,N_5770,N_5736);
or U6736 (N_6736,N_5148,N_5759);
nor U6737 (N_6737,N_5669,N_5632);
and U6738 (N_6738,N_5717,N_5205);
or U6739 (N_6739,N_5703,N_5963);
and U6740 (N_6740,N_5950,N_5656);
xor U6741 (N_6741,N_5710,N_5566);
nor U6742 (N_6742,N_5314,N_5064);
nor U6743 (N_6743,N_5169,N_5063);
xnor U6744 (N_6744,N_5673,N_5163);
xor U6745 (N_6745,N_5154,N_5003);
nor U6746 (N_6746,N_5906,N_5995);
nor U6747 (N_6747,N_5832,N_5027);
nand U6748 (N_6748,N_5834,N_5296);
xnor U6749 (N_6749,N_5725,N_5536);
or U6750 (N_6750,N_5439,N_5925);
and U6751 (N_6751,N_5309,N_5623);
nand U6752 (N_6752,N_5705,N_5602);
nor U6753 (N_6753,N_5218,N_5524);
or U6754 (N_6754,N_5585,N_5388);
or U6755 (N_6755,N_5169,N_5682);
and U6756 (N_6756,N_5670,N_5055);
or U6757 (N_6757,N_5511,N_5403);
nand U6758 (N_6758,N_5327,N_5682);
nor U6759 (N_6759,N_5555,N_5270);
and U6760 (N_6760,N_5798,N_5826);
xnor U6761 (N_6761,N_5337,N_5545);
and U6762 (N_6762,N_5767,N_5869);
nor U6763 (N_6763,N_5219,N_5393);
and U6764 (N_6764,N_5487,N_5651);
xnor U6765 (N_6765,N_5750,N_5986);
or U6766 (N_6766,N_5244,N_5060);
or U6767 (N_6767,N_5232,N_5539);
nand U6768 (N_6768,N_5155,N_5707);
nand U6769 (N_6769,N_5835,N_5465);
nor U6770 (N_6770,N_5188,N_5397);
xor U6771 (N_6771,N_5208,N_5601);
and U6772 (N_6772,N_5591,N_5845);
and U6773 (N_6773,N_5087,N_5885);
nand U6774 (N_6774,N_5211,N_5227);
and U6775 (N_6775,N_5012,N_5232);
and U6776 (N_6776,N_5715,N_5574);
and U6777 (N_6777,N_5970,N_5064);
or U6778 (N_6778,N_5196,N_5200);
nand U6779 (N_6779,N_5286,N_5011);
or U6780 (N_6780,N_5157,N_5272);
and U6781 (N_6781,N_5692,N_5124);
nand U6782 (N_6782,N_5839,N_5662);
and U6783 (N_6783,N_5398,N_5454);
or U6784 (N_6784,N_5268,N_5189);
xnor U6785 (N_6785,N_5505,N_5557);
and U6786 (N_6786,N_5383,N_5616);
nand U6787 (N_6787,N_5981,N_5762);
xnor U6788 (N_6788,N_5106,N_5291);
nand U6789 (N_6789,N_5122,N_5838);
nor U6790 (N_6790,N_5829,N_5592);
and U6791 (N_6791,N_5045,N_5363);
and U6792 (N_6792,N_5714,N_5218);
and U6793 (N_6793,N_5308,N_5343);
or U6794 (N_6794,N_5287,N_5838);
nor U6795 (N_6795,N_5873,N_5845);
nor U6796 (N_6796,N_5188,N_5693);
or U6797 (N_6797,N_5181,N_5226);
and U6798 (N_6798,N_5056,N_5108);
xnor U6799 (N_6799,N_5500,N_5106);
nand U6800 (N_6800,N_5470,N_5640);
nand U6801 (N_6801,N_5602,N_5150);
xnor U6802 (N_6802,N_5724,N_5898);
nand U6803 (N_6803,N_5491,N_5493);
nor U6804 (N_6804,N_5059,N_5301);
xnor U6805 (N_6805,N_5887,N_5704);
nor U6806 (N_6806,N_5048,N_5044);
xor U6807 (N_6807,N_5691,N_5806);
nand U6808 (N_6808,N_5632,N_5257);
and U6809 (N_6809,N_5388,N_5596);
or U6810 (N_6810,N_5529,N_5649);
nor U6811 (N_6811,N_5730,N_5406);
and U6812 (N_6812,N_5520,N_5379);
and U6813 (N_6813,N_5679,N_5690);
or U6814 (N_6814,N_5329,N_5201);
or U6815 (N_6815,N_5114,N_5368);
nor U6816 (N_6816,N_5006,N_5957);
and U6817 (N_6817,N_5928,N_5369);
or U6818 (N_6818,N_5415,N_5279);
xor U6819 (N_6819,N_5316,N_5340);
or U6820 (N_6820,N_5992,N_5725);
or U6821 (N_6821,N_5114,N_5311);
nor U6822 (N_6822,N_5647,N_5899);
nor U6823 (N_6823,N_5869,N_5701);
or U6824 (N_6824,N_5757,N_5493);
xor U6825 (N_6825,N_5894,N_5006);
xnor U6826 (N_6826,N_5704,N_5689);
and U6827 (N_6827,N_5713,N_5573);
nand U6828 (N_6828,N_5622,N_5232);
nor U6829 (N_6829,N_5506,N_5219);
and U6830 (N_6830,N_5286,N_5953);
nor U6831 (N_6831,N_5064,N_5702);
or U6832 (N_6832,N_5904,N_5470);
xor U6833 (N_6833,N_5113,N_5252);
or U6834 (N_6834,N_5226,N_5079);
nand U6835 (N_6835,N_5227,N_5139);
or U6836 (N_6836,N_5911,N_5471);
or U6837 (N_6837,N_5800,N_5431);
nor U6838 (N_6838,N_5469,N_5405);
xnor U6839 (N_6839,N_5831,N_5265);
nor U6840 (N_6840,N_5531,N_5368);
and U6841 (N_6841,N_5068,N_5825);
xnor U6842 (N_6842,N_5169,N_5295);
xnor U6843 (N_6843,N_5811,N_5148);
and U6844 (N_6844,N_5878,N_5996);
nand U6845 (N_6845,N_5114,N_5217);
nand U6846 (N_6846,N_5086,N_5772);
nor U6847 (N_6847,N_5878,N_5065);
and U6848 (N_6848,N_5253,N_5535);
nor U6849 (N_6849,N_5382,N_5347);
nor U6850 (N_6850,N_5398,N_5110);
and U6851 (N_6851,N_5181,N_5824);
and U6852 (N_6852,N_5249,N_5640);
and U6853 (N_6853,N_5171,N_5821);
nand U6854 (N_6854,N_5712,N_5496);
nand U6855 (N_6855,N_5769,N_5384);
or U6856 (N_6856,N_5070,N_5396);
and U6857 (N_6857,N_5910,N_5884);
or U6858 (N_6858,N_5939,N_5446);
nor U6859 (N_6859,N_5155,N_5804);
and U6860 (N_6860,N_5610,N_5995);
xor U6861 (N_6861,N_5506,N_5849);
or U6862 (N_6862,N_5918,N_5529);
nand U6863 (N_6863,N_5469,N_5764);
or U6864 (N_6864,N_5234,N_5413);
nor U6865 (N_6865,N_5710,N_5456);
or U6866 (N_6866,N_5190,N_5735);
nor U6867 (N_6867,N_5521,N_5617);
and U6868 (N_6868,N_5446,N_5342);
and U6869 (N_6869,N_5442,N_5696);
xor U6870 (N_6870,N_5910,N_5041);
nand U6871 (N_6871,N_5696,N_5797);
and U6872 (N_6872,N_5961,N_5219);
nand U6873 (N_6873,N_5448,N_5671);
and U6874 (N_6874,N_5469,N_5956);
xnor U6875 (N_6875,N_5146,N_5792);
nand U6876 (N_6876,N_5441,N_5279);
nand U6877 (N_6877,N_5263,N_5312);
nor U6878 (N_6878,N_5263,N_5356);
and U6879 (N_6879,N_5984,N_5162);
nor U6880 (N_6880,N_5234,N_5704);
nand U6881 (N_6881,N_5728,N_5691);
or U6882 (N_6882,N_5299,N_5416);
and U6883 (N_6883,N_5945,N_5485);
nand U6884 (N_6884,N_5714,N_5812);
xor U6885 (N_6885,N_5228,N_5776);
nand U6886 (N_6886,N_5646,N_5384);
nand U6887 (N_6887,N_5530,N_5081);
nand U6888 (N_6888,N_5949,N_5078);
nand U6889 (N_6889,N_5172,N_5156);
or U6890 (N_6890,N_5960,N_5087);
nor U6891 (N_6891,N_5676,N_5503);
and U6892 (N_6892,N_5339,N_5848);
or U6893 (N_6893,N_5480,N_5819);
and U6894 (N_6894,N_5121,N_5970);
nor U6895 (N_6895,N_5784,N_5636);
or U6896 (N_6896,N_5752,N_5941);
nand U6897 (N_6897,N_5813,N_5206);
or U6898 (N_6898,N_5232,N_5138);
xor U6899 (N_6899,N_5015,N_5765);
or U6900 (N_6900,N_5767,N_5471);
and U6901 (N_6901,N_5686,N_5872);
and U6902 (N_6902,N_5400,N_5096);
or U6903 (N_6903,N_5585,N_5402);
and U6904 (N_6904,N_5354,N_5467);
or U6905 (N_6905,N_5693,N_5826);
and U6906 (N_6906,N_5782,N_5150);
or U6907 (N_6907,N_5323,N_5792);
nand U6908 (N_6908,N_5894,N_5970);
nor U6909 (N_6909,N_5278,N_5530);
or U6910 (N_6910,N_5027,N_5404);
and U6911 (N_6911,N_5789,N_5820);
nand U6912 (N_6912,N_5170,N_5364);
and U6913 (N_6913,N_5140,N_5960);
or U6914 (N_6914,N_5034,N_5478);
and U6915 (N_6915,N_5245,N_5853);
nand U6916 (N_6916,N_5222,N_5283);
or U6917 (N_6917,N_5810,N_5452);
or U6918 (N_6918,N_5384,N_5922);
or U6919 (N_6919,N_5174,N_5688);
nor U6920 (N_6920,N_5667,N_5974);
and U6921 (N_6921,N_5293,N_5627);
nor U6922 (N_6922,N_5470,N_5515);
nor U6923 (N_6923,N_5419,N_5132);
and U6924 (N_6924,N_5431,N_5174);
nand U6925 (N_6925,N_5641,N_5655);
nor U6926 (N_6926,N_5160,N_5886);
xnor U6927 (N_6927,N_5819,N_5165);
xor U6928 (N_6928,N_5656,N_5137);
and U6929 (N_6929,N_5932,N_5749);
xor U6930 (N_6930,N_5112,N_5479);
nor U6931 (N_6931,N_5267,N_5043);
nor U6932 (N_6932,N_5864,N_5444);
nand U6933 (N_6933,N_5220,N_5316);
nand U6934 (N_6934,N_5203,N_5973);
xor U6935 (N_6935,N_5364,N_5099);
and U6936 (N_6936,N_5418,N_5866);
and U6937 (N_6937,N_5799,N_5980);
or U6938 (N_6938,N_5116,N_5501);
nand U6939 (N_6939,N_5144,N_5416);
nand U6940 (N_6940,N_5551,N_5723);
and U6941 (N_6941,N_5372,N_5670);
nor U6942 (N_6942,N_5440,N_5370);
and U6943 (N_6943,N_5181,N_5626);
nor U6944 (N_6944,N_5545,N_5406);
and U6945 (N_6945,N_5758,N_5719);
nor U6946 (N_6946,N_5990,N_5573);
nor U6947 (N_6947,N_5528,N_5849);
nor U6948 (N_6948,N_5697,N_5548);
nand U6949 (N_6949,N_5887,N_5620);
nor U6950 (N_6950,N_5771,N_5471);
nor U6951 (N_6951,N_5865,N_5115);
and U6952 (N_6952,N_5350,N_5957);
xor U6953 (N_6953,N_5551,N_5171);
and U6954 (N_6954,N_5796,N_5967);
nor U6955 (N_6955,N_5384,N_5165);
nor U6956 (N_6956,N_5494,N_5912);
nand U6957 (N_6957,N_5806,N_5751);
and U6958 (N_6958,N_5973,N_5190);
xor U6959 (N_6959,N_5102,N_5205);
nor U6960 (N_6960,N_5637,N_5247);
and U6961 (N_6961,N_5736,N_5156);
nand U6962 (N_6962,N_5022,N_5576);
nand U6963 (N_6963,N_5377,N_5401);
and U6964 (N_6964,N_5369,N_5444);
or U6965 (N_6965,N_5708,N_5348);
and U6966 (N_6966,N_5671,N_5010);
nand U6967 (N_6967,N_5765,N_5010);
nand U6968 (N_6968,N_5734,N_5024);
and U6969 (N_6969,N_5257,N_5169);
nand U6970 (N_6970,N_5528,N_5831);
xnor U6971 (N_6971,N_5092,N_5314);
nand U6972 (N_6972,N_5685,N_5917);
nand U6973 (N_6973,N_5213,N_5723);
and U6974 (N_6974,N_5270,N_5550);
nor U6975 (N_6975,N_5569,N_5953);
xnor U6976 (N_6976,N_5150,N_5229);
or U6977 (N_6977,N_5204,N_5132);
and U6978 (N_6978,N_5594,N_5169);
xnor U6979 (N_6979,N_5590,N_5222);
and U6980 (N_6980,N_5981,N_5549);
nor U6981 (N_6981,N_5539,N_5372);
xnor U6982 (N_6982,N_5796,N_5833);
and U6983 (N_6983,N_5258,N_5450);
xor U6984 (N_6984,N_5076,N_5990);
or U6985 (N_6985,N_5915,N_5737);
nor U6986 (N_6986,N_5254,N_5324);
xnor U6987 (N_6987,N_5219,N_5160);
and U6988 (N_6988,N_5984,N_5227);
nor U6989 (N_6989,N_5516,N_5717);
xor U6990 (N_6990,N_5590,N_5297);
nor U6991 (N_6991,N_5744,N_5571);
and U6992 (N_6992,N_5501,N_5635);
xnor U6993 (N_6993,N_5210,N_5349);
or U6994 (N_6994,N_5164,N_5286);
nor U6995 (N_6995,N_5145,N_5437);
and U6996 (N_6996,N_5178,N_5001);
xor U6997 (N_6997,N_5840,N_5628);
or U6998 (N_6998,N_5356,N_5390);
and U6999 (N_6999,N_5408,N_5193);
nor U7000 (N_7000,N_6227,N_6699);
or U7001 (N_7001,N_6274,N_6611);
and U7002 (N_7002,N_6341,N_6400);
or U7003 (N_7003,N_6457,N_6352);
or U7004 (N_7004,N_6226,N_6174);
nand U7005 (N_7005,N_6083,N_6888);
nand U7006 (N_7006,N_6655,N_6740);
and U7007 (N_7007,N_6490,N_6332);
or U7008 (N_7008,N_6092,N_6695);
and U7009 (N_7009,N_6294,N_6283);
xnor U7010 (N_7010,N_6062,N_6266);
nor U7011 (N_7011,N_6839,N_6620);
xor U7012 (N_7012,N_6074,N_6001);
xnor U7013 (N_7013,N_6840,N_6604);
nand U7014 (N_7014,N_6536,N_6656);
xor U7015 (N_7015,N_6265,N_6080);
and U7016 (N_7016,N_6072,N_6220);
and U7017 (N_7017,N_6392,N_6033);
nand U7018 (N_7018,N_6737,N_6638);
or U7019 (N_7019,N_6213,N_6731);
or U7020 (N_7020,N_6712,N_6928);
xor U7021 (N_7021,N_6500,N_6534);
nor U7022 (N_7022,N_6037,N_6187);
xnor U7023 (N_7023,N_6607,N_6152);
nor U7024 (N_7024,N_6235,N_6464);
nor U7025 (N_7025,N_6527,N_6881);
nand U7026 (N_7026,N_6569,N_6866);
nand U7027 (N_7027,N_6264,N_6943);
and U7028 (N_7028,N_6207,N_6519);
or U7029 (N_7029,N_6556,N_6508);
xnor U7030 (N_7030,N_6289,N_6766);
and U7031 (N_7031,N_6125,N_6372);
nor U7032 (N_7032,N_6005,N_6716);
nor U7033 (N_7033,N_6311,N_6538);
xor U7034 (N_7034,N_6568,N_6946);
nand U7035 (N_7035,N_6885,N_6403);
or U7036 (N_7036,N_6804,N_6326);
xor U7037 (N_7037,N_6692,N_6843);
and U7038 (N_7038,N_6271,N_6587);
nor U7039 (N_7039,N_6939,N_6028);
or U7040 (N_7040,N_6432,N_6564);
or U7041 (N_7041,N_6309,N_6325);
or U7042 (N_7042,N_6618,N_6511);
or U7043 (N_7043,N_6348,N_6206);
nand U7044 (N_7044,N_6136,N_6233);
or U7045 (N_7045,N_6886,N_6912);
and U7046 (N_7046,N_6520,N_6635);
xor U7047 (N_7047,N_6544,N_6724);
and U7048 (N_7048,N_6224,N_6720);
nor U7049 (N_7049,N_6871,N_6561);
nand U7050 (N_7050,N_6803,N_6454);
nand U7051 (N_7051,N_6088,N_6095);
and U7052 (N_7052,N_6982,N_6475);
and U7053 (N_7053,N_6239,N_6999);
and U7054 (N_7054,N_6767,N_6217);
nor U7055 (N_7055,N_6507,N_6418);
and U7056 (N_7056,N_6509,N_6112);
nor U7057 (N_7057,N_6698,N_6060);
and U7058 (N_7058,N_6019,N_6176);
nand U7059 (N_7059,N_6191,N_6482);
and U7060 (N_7060,N_6964,N_6055);
xor U7061 (N_7061,N_6503,N_6185);
and U7062 (N_7062,N_6933,N_6230);
and U7063 (N_7063,N_6308,N_6253);
xor U7064 (N_7064,N_6693,N_6257);
nand U7065 (N_7065,N_6063,N_6468);
nand U7066 (N_7066,N_6778,N_6354);
xor U7067 (N_7067,N_6818,N_6355);
or U7068 (N_7068,N_6020,N_6727);
and U7069 (N_7069,N_6387,N_6413);
nor U7070 (N_7070,N_6184,N_6735);
nand U7071 (N_7071,N_6593,N_6109);
xor U7072 (N_7072,N_6915,N_6076);
nor U7073 (N_7073,N_6646,N_6153);
xnor U7074 (N_7074,N_6932,N_6445);
nand U7075 (N_7075,N_6142,N_6874);
or U7076 (N_7076,N_6009,N_6234);
nor U7077 (N_7077,N_6942,N_6087);
nor U7078 (N_7078,N_6730,N_6829);
nor U7079 (N_7079,N_6314,N_6822);
nand U7080 (N_7080,N_6243,N_6399);
xor U7081 (N_7081,N_6713,N_6110);
xnor U7082 (N_7082,N_6524,N_6175);
nor U7083 (N_7083,N_6258,N_6006);
or U7084 (N_7084,N_6754,N_6526);
nand U7085 (N_7085,N_6797,N_6542);
nand U7086 (N_7086,N_6018,N_6002);
nor U7087 (N_7087,N_6390,N_6627);
and U7088 (N_7088,N_6657,N_6976);
xnor U7089 (N_7089,N_6130,N_6780);
nand U7090 (N_7090,N_6472,N_6459);
nand U7091 (N_7091,N_6952,N_6518);
nor U7092 (N_7092,N_6197,N_6192);
or U7093 (N_7093,N_6396,N_6555);
nor U7094 (N_7094,N_6752,N_6451);
or U7095 (N_7095,N_6788,N_6378);
xor U7096 (N_7096,N_6823,N_6267);
nor U7097 (N_7097,N_6800,N_6956);
and U7098 (N_7098,N_6064,N_6375);
nor U7099 (N_7099,N_6733,N_6120);
and U7100 (N_7100,N_6809,N_6113);
xnor U7101 (N_7101,N_6049,N_6669);
nor U7102 (N_7102,N_6750,N_6558);
nand U7103 (N_7103,N_6497,N_6602);
nor U7104 (N_7104,N_6216,N_6521);
and U7105 (N_7105,N_6208,N_6397);
or U7106 (N_7106,N_6414,N_6746);
nor U7107 (N_7107,N_6858,N_6917);
and U7108 (N_7108,N_6862,N_6786);
xor U7109 (N_7109,N_6448,N_6517);
nand U7110 (N_7110,N_6395,N_6742);
and U7111 (N_7111,N_6936,N_6749);
xor U7112 (N_7112,N_6630,N_6697);
and U7113 (N_7113,N_6588,N_6491);
xnor U7114 (N_7114,N_6983,N_6854);
or U7115 (N_7115,N_6545,N_6447);
xor U7116 (N_7116,N_6904,N_6071);
xor U7117 (N_7117,N_6559,N_6957);
nand U7118 (N_7118,N_6950,N_6790);
nor U7119 (N_7119,N_6909,N_6641);
and U7120 (N_7120,N_6209,N_6580);
or U7121 (N_7121,N_6241,N_6969);
nor U7122 (N_7122,N_6248,N_6310);
nand U7123 (N_7123,N_6044,N_6831);
xnor U7124 (N_7124,N_6811,N_6801);
xnor U7125 (N_7125,N_6645,N_6900);
or U7126 (N_7126,N_6812,N_6478);
or U7127 (N_7127,N_6411,N_6628);
nor U7128 (N_7128,N_6144,N_6914);
or U7129 (N_7129,N_6439,N_6993);
nand U7130 (N_7130,N_6863,N_6861);
or U7131 (N_7131,N_6262,N_6869);
and U7132 (N_7132,N_6600,N_6703);
nor U7133 (N_7133,N_6732,N_6003);
or U7134 (N_7134,N_6211,N_6654);
or U7135 (N_7135,N_6436,N_6717);
nand U7136 (N_7136,N_6726,N_6927);
or U7137 (N_7137,N_6642,N_6833);
nand U7138 (N_7138,N_6427,N_6129);
and U7139 (N_7139,N_6896,N_6616);
nand U7140 (N_7140,N_6331,N_6947);
nand U7141 (N_7141,N_6825,N_6919);
xnor U7142 (N_7142,N_6963,N_6237);
xnor U7143 (N_7143,N_6887,N_6596);
xor U7144 (N_7144,N_6968,N_6548);
nand U7145 (N_7145,N_6834,N_6098);
and U7146 (N_7146,N_6270,N_6483);
nand U7147 (N_7147,N_6091,N_6700);
nor U7148 (N_7148,N_6884,N_6941);
and U7149 (N_7149,N_6922,N_6086);
nor U7150 (N_7150,N_6461,N_6054);
or U7151 (N_7151,N_6782,N_6452);
nor U7152 (N_7152,N_6783,N_6614);
nor U7153 (N_7153,N_6127,N_6771);
xnor U7154 (N_7154,N_6386,N_6768);
nand U7155 (N_7155,N_6361,N_6819);
nor U7156 (N_7156,N_6948,N_6402);
or U7157 (N_7157,N_6278,N_6196);
nor U7158 (N_7158,N_6532,N_6624);
nor U7159 (N_7159,N_6004,N_6202);
or U7160 (N_7160,N_6077,N_6991);
nand U7161 (N_7161,N_6017,N_6494);
and U7162 (N_7162,N_6745,N_6841);
nor U7163 (N_7163,N_6813,N_6101);
nand U7164 (N_7164,N_6433,N_6640);
nand U7165 (N_7165,N_6515,N_6553);
nand U7166 (N_7166,N_6140,N_6911);
or U7167 (N_7167,N_6867,N_6444);
nand U7168 (N_7168,N_6530,N_6625);
nor U7169 (N_7169,N_6333,N_6894);
xnor U7170 (N_7170,N_6141,N_6015);
xnor U7171 (N_7171,N_6131,N_6694);
or U7172 (N_7172,N_6706,N_6428);
xnor U7173 (N_7173,N_6617,N_6690);
nand U7174 (N_7174,N_6990,N_6636);
and U7175 (N_7175,N_6225,N_6670);
and U7176 (N_7176,N_6252,N_6193);
or U7177 (N_7177,N_6552,N_6541);
or U7178 (N_7178,N_6073,N_6791);
or U7179 (N_7179,N_6031,N_6830);
or U7180 (N_7180,N_6907,N_6421);
and U7181 (N_7181,N_6998,N_6743);
nand U7182 (N_7182,N_6473,N_6154);
and U7183 (N_7183,N_6393,N_6025);
nand U7184 (N_7184,N_6633,N_6081);
nor U7185 (N_7185,N_6895,N_6210);
or U7186 (N_7186,N_6057,N_6759);
nor U7187 (N_7187,N_6504,N_6644);
or U7188 (N_7188,N_6047,N_6940);
or U7189 (N_7189,N_6238,N_6359);
nor U7190 (N_7190,N_6570,N_6150);
or U7191 (N_7191,N_6868,N_6165);
nand U7192 (N_7192,N_6546,N_6471);
xnor U7193 (N_7193,N_6183,N_6404);
nand U7194 (N_7194,N_6719,N_6371);
nor U7195 (N_7195,N_6835,N_6857);
nand U7196 (N_7196,N_6753,N_6032);
or U7197 (N_7197,N_6997,N_6014);
and U7198 (N_7198,N_6229,N_6499);
xor U7199 (N_7199,N_6067,N_6677);
xor U7200 (N_7200,N_6701,N_6648);
or U7201 (N_7201,N_6551,N_6531);
xor U7202 (N_7202,N_6898,N_6322);
nor U7203 (N_7203,N_6251,N_6851);
nand U7204 (N_7204,N_6498,N_6051);
xnor U7205 (N_7205,N_6079,N_6357);
nor U7206 (N_7206,N_6989,N_6808);
nor U7207 (N_7207,N_6662,N_6302);
or U7208 (N_7208,N_6440,N_6287);
nand U7209 (N_7209,N_6180,N_6889);
or U7210 (N_7210,N_6883,N_6290);
nor U7211 (N_7211,N_6035,N_6902);
xnor U7212 (N_7212,N_6373,N_6685);
and U7213 (N_7213,N_6317,N_6951);
nor U7214 (N_7214,N_6115,N_6805);
or U7215 (N_7215,N_6024,N_6675);
nand U7216 (N_7216,N_6446,N_6415);
or U7217 (N_7217,N_6986,N_6505);
nor U7218 (N_7218,N_6401,N_6050);
and U7219 (N_7219,N_6996,N_6441);
or U7220 (N_7220,N_6242,N_6554);
xnor U7221 (N_7221,N_6784,N_6179);
and U7222 (N_7222,N_6592,N_6897);
and U7223 (N_7223,N_6796,N_6377);
nor U7224 (N_7224,N_6231,N_6350);
nor U7225 (N_7225,N_6299,N_6579);
xor U7226 (N_7226,N_6585,N_6279);
xnor U7227 (N_7227,N_6342,N_6626);
nor U7228 (N_7228,N_6034,N_6222);
or U7229 (N_7229,N_6424,N_6984);
xor U7230 (N_7230,N_6995,N_6022);
xnor U7231 (N_7231,N_6622,N_6108);
nand U7232 (N_7232,N_6802,N_6026);
or U7233 (N_7233,N_6385,N_6219);
xnor U7234 (N_7234,N_6543,N_6351);
nor U7235 (N_7235,N_6970,N_6935);
nor U7236 (N_7236,N_6338,N_6199);
xnor U7237 (N_7237,N_6070,N_6300);
nand U7238 (N_7238,N_6761,N_6277);
nand U7239 (N_7239,N_6945,N_6959);
and U7240 (N_7240,N_6773,N_6434);
or U7241 (N_7241,N_6296,N_6815);
or U7242 (N_7242,N_6806,N_6793);
or U7243 (N_7243,N_6307,N_6059);
xor U7244 (N_7244,N_6085,N_6965);
or U7245 (N_7245,N_6336,N_6876);
or U7246 (N_7246,N_6106,N_6463);
nor U7247 (N_7247,N_6288,N_6123);
and U7248 (N_7248,N_6673,N_6814);
xor U7249 (N_7249,N_6666,N_6540);
or U7250 (N_7250,N_6852,N_6516);
nand U7251 (N_7251,N_6882,N_6488);
nor U7252 (N_7252,N_6056,N_6158);
nor U7253 (N_7253,N_6276,N_6613);
nor U7254 (N_7254,N_6736,N_6107);
or U7255 (N_7255,N_6221,N_6653);
nor U7256 (N_7256,N_6757,N_6537);
nor U7257 (N_7257,N_6715,N_6122);
nor U7258 (N_7258,N_6286,N_6291);
xnor U7259 (N_7259,N_6244,N_6953);
nand U7260 (N_7260,N_6356,N_6755);
and U7261 (N_7261,N_6584,N_6388);
or U7262 (N_7262,N_6103,N_6529);
xnor U7263 (N_7263,N_6744,N_6301);
and U7264 (N_7264,N_6619,N_6937);
nand U7265 (N_7265,N_6621,N_6923);
xnor U7266 (N_7266,N_6828,N_6879);
nor U7267 (N_7267,N_6577,N_6042);
xor U7268 (N_7268,N_6438,N_6925);
xor U7269 (N_7269,N_6921,N_6182);
or U7270 (N_7270,N_6038,N_6789);
xor U7271 (N_7271,N_6161,N_6634);
xor U7272 (N_7272,N_6949,N_6149);
nor U7273 (N_7273,N_6629,N_6875);
and U7274 (N_7274,N_6487,N_6479);
or U7275 (N_7275,N_6610,N_6676);
xnor U7276 (N_7276,N_6683,N_6272);
xnor U7277 (N_7277,N_6606,N_6566);
nand U7278 (N_7278,N_6492,N_6763);
nand U7279 (N_7279,N_6236,N_6118);
xor U7280 (N_7280,N_6495,N_6493);
or U7281 (N_7281,N_6430,N_6668);
nand U7282 (N_7282,N_6159,N_6929);
or U7283 (N_7283,N_6245,N_6533);
nor U7284 (N_7284,N_6799,N_6539);
or U7285 (N_7285,N_6794,N_6985);
nor U7286 (N_7286,N_6160,N_6597);
xor U7287 (N_7287,N_6691,N_6955);
nor U7288 (N_7288,N_6068,N_6714);
or U7289 (N_7289,N_6178,N_6305);
xnor U7290 (N_7290,N_6878,N_6586);
and U7291 (N_7291,N_6156,N_6977);
nor U7292 (N_7292,N_6981,N_6679);
or U7293 (N_7293,N_6816,N_6345);
and U7294 (N_7294,N_6650,N_6194);
or U7295 (N_7295,N_6609,N_6162);
xor U7296 (N_7296,N_6820,N_6329);
nand U7297 (N_7297,N_6320,N_6281);
xnor U7298 (N_7298,N_6481,N_6704);
nor U7299 (N_7299,N_6836,N_6458);
and U7300 (N_7300,N_6261,N_6817);
nor U7301 (N_7301,N_6030,N_6417);
and U7302 (N_7302,N_6164,N_6738);
or U7303 (N_7303,N_6431,N_6708);
nand U7304 (N_7304,N_6637,N_6795);
xor U7305 (N_7305,N_6639,N_6297);
or U7306 (N_7306,N_6844,N_6827);
nor U7307 (N_7307,N_6994,N_6920);
xnor U7308 (N_7308,N_6944,N_6426);
nor U7309 (N_7309,N_6480,N_6383);
and U7310 (N_7310,N_6807,N_6456);
xor U7311 (N_7311,N_6850,N_6573);
nor U7312 (N_7312,N_6254,N_6798);
nand U7313 (N_7313,N_6476,N_6133);
or U7314 (N_7314,N_6340,N_6760);
and U7315 (N_7315,N_6873,N_6785);
xnor U7316 (N_7316,N_6781,N_6126);
xor U7317 (N_7317,N_6412,N_6284);
or U7318 (N_7318,N_6318,N_6398);
or U7319 (N_7319,N_6901,N_6563);
and U7320 (N_7320,N_6962,N_6718);
nand U7321 (N_7321,N_6973,N_6260);
nand U7322 (N_7322,N_6603,N_6409);
xor U7323 (N_7323,N_6339,N_6891);
xor U7324 (N_7324,N_6729,N_6214);
nor U7325 (N_7325,N_6443,N_6293);
and U7326 (N_7326,N_6405,N_6711);
xnor U7327 (N_7327,N_6595,N_6263);
and U7328 (N_7328,N_6615,N_6337);
xnor U7329 (N_7329,N_6723,N_6273);
and U7330 (N_7330,N_6938,N_6572);
nand U7331 (N_7331,N_6751,N_6893);
nand U7332 (N_7332,N_6960,N_6143);
xnor U7333 (N_7333,N_6510,N_6872);
nand U7334 (N_7334,N_6212,N_6041);
nor U7335 (N_7335,N_6145,N_6416);
or U7336 (N_7336,N_6232,N_6096);
xor U7337 (N_7337,N_6249,N_6138);
xnor U7338 (N_7338,N_6292,N_6578);
nand U7339 (N_7339,N_6171,N_6764);
and U7340 (N_7340,N_6847,N_6484);
xor U7341 (N_7341,N_6330,N_6967);
nand U7342 (N_7342,N_6169,N_6389);
nor U7343 (N_7343,N_6899,N_6855);
or U7344 (N_7344,N_6021,N_6364);
nor U7345 (N_7345,N_6215,N_6410);
nor U7346 (N_7346,N_6155,N_6696);
and U7347 (N_7347,N_6363,N_6651);
nand U7348 (N_7348,N_6870,N_6890);
xor U7349 (N_7349,N_6643,N_6369);
or U7350 (N_7350,N_6571,N_6303);
xor U7351 (N_7351,N_6280,N_6173);
nor U7352 (N_7352,N_6687,N_6849);
nand U7353 (N_7353,N_6787,N_6934);
and U7354 (N_7354,N_6407,N_6705);
xor U7355 (N_7355,N_6016,N_6612);
and U7356 (N_7356,N_6528,N_6027);
xnor U7357 (N_7357,N_6078,N_6671);
nor U7358 (N_7358,N_6734,N_6758);
and U7359 (N_7359,N_6157,N_6837);
and U7360 (N_7360,N_6008,N_6605);
xor U7361 (N_7361,N_6775,N_6324);
and U7362 (N_7362,N_6139,N_6061);
xnor U7363 (N_7363,N_6681,N_6343);
nand U7364 (N_7364,N_6574,N_6501);
xnor U7365 (N_7365,N_6470,N_6722);
and U7366 (N_7366,N_6094,N_6474);
xnor U7367 (N_7367,N_6661,N_6465);
nand U7368 (N_7368,N_6043,N_6346);
or U7369 (N_7369,N_6576,N_6710);
nand U7370 (N_7370,N_6181,N_6089);
xnor U7371 (N_7371,N_6664,N_6462);
xor U7372 (N_7372,N_6298,N_6845);
and U7373 (N_7373,N_6581,N_6741);
nor U7374 (N_7374,N_6066,N_6512);
xor U7375 (N_7375,N_6667,N_6678);
nand U7376 (N_7376,N_6368,N_6201);
nor U7377 (N_7377,N_6315,N_6926);
nor U7378 (N_7378,N_6707,N_6082);
or U7379 (N_7379,N_6665,N_6040);
and U7380 (N_7380,N_6104,N_6408);
and U7381 (N_7381,N_6560,N_6362);
and U7382 (N_7382,N_6382,N_6792);
nand U7383 (N_7383,N_6877,N_6598);
xor U7384 (N_7384,N_6374,N_6992);
xnor U7385 (N_7385,N_6370,N_6012);
and U7386 (N_7386,N_6514,N_6918);
xor U7387 (N_7387,N_6334,N_6381);
or U7388 (N_7388,N_6659,N_6198);
nand U7389 (N_7389,N_6429,N_6589);
nor U7390 (N_7390,N_6313,N_6966);
nand U7391 (N_7391,N_6978,N_6376);
and U7392 (N_7392,N_6961,N_6682);
xor U7393 (N_7393,N_6011,N_6958);
and U7394 (N_7394,N_6188,N_6166);
and U7395 (N_7395,N_6367,N_6099);
or U7396 (N_7396,N_6756,N_6349);
and U7397 (N_7397,N_6496,N_6218);
nor U7398 (N_7398,N_6137,N_6748);
or U7399 (N_7399,N_6525,N_6535);
xnor U7400 (N_7400,N_6721,N_6975);
nand U7401 (N_7401,N_6327,N_6590);
and U7402 (N_7402,N_6240,N_6304);
or U7403 (N_7403,N_6916,N_6848);
xnor U7404 (N_7404,N_6972,N_6486);
nand U7405 (N_7405,N_6366,N_6549);
or U7406 (N_7406,N_6846,N_6859);
or U7407 (N_7407,N_6905,N_6599);
nand U7408 (N_7408,N_6203,N_6910);
nand U7409 (N_7409,N_6776,N_6268);
xnor U7410 (N_7410,N_6420,N_6772);
and U7411 (N_7411,N_6777,N_6177);
and U7412 (N_7412,N_6102,N_6762);
and U7413 (N_7413,N_6892,N_6010);
xor U7414 (N_7414,N_6347,N_6663);
and U7415 (N_7415,N_6316,N_6779);
xnor U7416 (N_7416,N_6065,N_6631);
and U7417 (N_7417,N_6608,N_6913);
or U7418 (N_7418,N_6575,N_6450);
nor U7419 (N_7419,N_6660,N_6148);
and U7420 (N_7420,N_6954,N_6048);
nand U7421 (N_7421,N_6709,N_6591);
and U7422 (N_7422,N_6124,N_6146);
or U7423 (N_7423,N_6097,N_6652);
xor U7424 (N_7424,N_6285,N_6105);
nand U7425 (N_7425,N_6513,N_6435);
nor U7426 (N_7426,N_6466,N_6824);
nor U7427 (N_7427,N_6601,N_6980);
and U7428 (N_7428,N_6255,N_6686);
or U7429 (N_7429,N_6151,N_6275);
or U7430 (N_7430,N_6856,N_6128);
nor U7431 (N_7431,N_6582,N_6384);
nand U7432 (N_7432,N_6924,N_6100);
and U7433 (N_7433,N_6931,N_6979);
nand U7434 (N_7434,N_6190,N_6684);
or U7435 (N_7435,N_6728,N_6247);
nand U7436 (N_7436,N_6419,N_6770);
xnor U7437 (N_7437,N_6121,N_6647);
xnor U7438 (N_7438,N_6774,N_6000);
nor U7439 (N_7439,N_6282,N_6455);
nor U7440 (N_7440,N_6172,N_6632);
or U7441 (N_7441,N_6688,N_6036);
nand U7442 (N_7442,N_6195,N_6437);
xor U7443 (N_7443,N_6204,N_6114);
nor U7444 (N_7444,N_6328,N_6246);
or U7445 (N_7445,N_6562,N_6565);
xnor U7446 (N_7446,N_6547,N_6360);
nor U7447 (N_7447,N_6422,N_6117);
or U7448 (N_7448,N_6167,N_6903);
or U7449 (N_7449,N_6013,N_6379);
or U7450 (N_7450,N_6906,N_6550);
xnor U7451 (N_7451,N_6250,N_6987);
or U7452 (N_7452,N_6135,N_6842);
nor U7453 (N_7453,N_6864,N_6406);
nand U7454 (N_7454,N_6522,N_6344);
xnor U7455 (N_7455,N_6594,N_6702);
and U7456 (N_7456,N_6467,N_6200);
xnor U7457 (N_7457,N_6477,N_6658);
xnor U7458 (N_7458,N_6442,N_6306);
nor U7459 (N_7459,N_6323,N_6075);
xor U7460 (N_7460,N_6674,N_6557);
nor U7461 (N_7461,N_6046,N_6423);
and U7462 (N_7462,N_6769,N_6090);
nor U7463 (N_7463,N_6353,N_6052);
xor U7464 (N_7464,N_6039,N_6295);
xor U7465 (N_7465,N_6205,N_6689);
nor U7466 (N_7466,N_6930,N_6132);
or U7467 (N_7467,N_6908,N_6449);
nor U7468 (N_7468,N_6069,N_6739);
xnor U7469 (N_7469,N_6335,N_6319);
nand U7470 (N_7470,N_6007,N_6093);
nand U7471 (N_7471,N_6583,N_6119);
xnor U7472 (N_7472,N_6259,N_6988);
nor U7473 (N_7473,N_6826,N_6058);
xor U7474 (N_7474,N_6453,N_6567);
and U7475 (N_7475,N_6256,N_6269);
xnor U7476 (N_7476,N_6485,N_6725);
xnor U7477 (N_7477,N_6860,N_6672);
xnor U7478 (N_7478,N_6765,N_6228);
nand U7479 (N_7479,N_6321,N_6649);
nor U7480 (N_7480,N_6186,N_6853);
xnor U7481 (N_7481,N_6506,N_6365);
and U7482 (N_7482,N_6111,N_6394);
or U7483 (N_7483,N_6747,N_6189);
or U7484 (N_7484,N_6358,N_6971);
nor U7485 (N_7485,N_6391,N_6023);
and U7486 (N_7486,N_6974,N_6380);
nand U7487 (N_7487,N_6147,N_6832);
xor U7488 (N_7488,N_6163,N_6489);
or U7489 (N_7489,N_6880,N_6460);
or U7490 (N_7490,N_6821,N_6469);
nor U7491 (N_7491,N_6680,N_6045);
or U7492 (N_7492,N_6116,N_6810);
nor U7493 (N_7493,N_6134,N_6502);
nand U7494 (N_7494,N_6223,N_6425);
nand U7495 (N_7495,N_6168,N_6170);
xnor U7496 (N_7496,N_6084,N_6312);
and U7497 (N_7497,N_6865,N_6523);
xnor U7498 (N_7498,N_6838,N_6029);
nand U7499 (N_7499,N_6623,N_6053);
and U7500 (N_7500,N_6619,N_6236);
and U7501 (N_7501,N_6913,N_6955);
nand U7502 (N_7502,N_6867,N_6817);
and U7503 (N_7503,N_6174,N_6286);
and U7504 (N_7504,N_6898,N_6007);
nand U7505 (N_7505,N_6984,N_6992);
xor U7506 (N_7506,N_6178,N_6025);
or U7507 (N_7507,N_6334,N_6692);
nor U7508 (N_7508,N_6344,N_6402);
nor U7509 (N_7509,N_6982,N_6464);
and U7510 (N_7510,N_6146,N_6834);
nor U7511 (N_7511,N_6269,N_6446);
xnor U7512 (N_7512,N_6510,N_6952);
nand U7513 (N_7513,N_6178,N_6050);
nand U7514 (N_7514,N_6093,N_6930);
or U7515 (N_7515,N_6247,N_6803);
and U7516 (N_7516,N_6414,N_6876);
and U7517 (N_7517,N_6125,N_6645);
nor U7518 (N_7518,N_6679,N_6001);
nor U7519 (N_7519,N_6645,N_6746);
nor U7520 (N_7520,N_6137,N_6182);
or U7521 (N_7521,N_6620,N_6770);
or U7522 (N_7522,N_6385,N_6190);
nand U7523 (N_7523,N_6664,N_6415);
and U7524 (N_7524,N_6790,N_6259);
nor U7525 (N_7525,N_6610,N_6426);
nor U7526 (N_7526,N_6708,N_6452);
or U7527 (N_7527,N_6741,N_6175);
xnor U7528 (N_7528,N_6465,N_6329);
and U7529 (N_7529,N_6693,N_6719);
and U7530 (N_7530,N_6243,N_6515);
and U7531 (N_7531,N_6509,N_6919);
nor U7532 (N_7532,N_6577,N_6901);
nand U7533 (N_7533,N_6570,N_6234);
or U7534 (N_7534,N_6808,N_6554);
xnor U7535 (N_7535,N_6555,N_6073);
or U7536 (N_7536,N_6255,N_6488);
or U7537 (N_7537,N_6574,N_6208);
xnor U7538 (N_7538,N_6326,N_6448);
nand U7539 (N_7539,N_6507,N_6302);
xor U7540 (N_7540,N_6972,N_6478);
xnor U7541 (N_7541,N_6643,N_6398);
and U7542 (N_7542,N_6736,N_6416);
nor U7543 (N_7543,N_6497,N_6203);
xnor U7544 (N_7544,N_6231,N_6786);
or U7545 (N_7545,N_6242,N_6115);
xor U7546 (N_7546,N_6019,N_6049);
xnor U7547 (N_7547,N_6254,N_6554);
nand U7548 (N_7548,N_6496,N_6894);
nor U7549 (N_7549,N_6649,N_6778);
xor U7550 (N_7550,N_6710,N_6599);
or U7551 (N_7551,N_6901,N_6122);
nand U7552 (N_7552,N_6465,N_6586);
nor U7553 (N_7553,N_6885,N_6427);
or U7554 (N_7554,N_6420,N_6373);
and U7555 (N_7555,N_6829,N_6815);
and U7556 (N_7556,N_6152,N_6239);
or U7557 (N_7557,N_6253,N_6715);
nor U7558 (N_7558,N_6911,N_6875);
nor U7559 (N_7559,N_6402,N_6478);
nor U7560 (N_7560,N_6794,N_6090);
nand U7561 (N_7561,N_6621,N_6420);
or U7562 (N_7562,N_6263,N_6940);
nand U7563 (N_7563,N_6817,N_6970);
nor U7564 (N_7564,N_6995,N_6234);
nand U7565 (N_7565,N_6453,N_6131);
xor U7566 (N_7566,N_6921,N_6196);
or U7567 (N_7567,N_6234,N_6035);
or U7568 (N_7568,N_6616,N_6191);
nor U7569 (N_7569,N_6523,N_6510);
and U7570 (N_7570,N_6190,N_6437);
and U7571 (N_7571,N_6906,N_6279);
nor U7572 (N_7572,N_6899,N_6064);
nor U7573 (N_7573,N_6032,N_6477);
or U7574 (N_7574,N_6261,N_6546);
nand U7575 (N_7575,N_6826,N_6961);
xor U7576 (N_7576,N_6281,N_6539);
nor U7577 (N_7577,N_6032,N_6333);
nand U7578 (N_7578,N_6585,N_6913);
or U7579 (N_7579,N_6971,N_6199);
nor U7580 (N_7580,N_6351,N_6831);
nand U7581 (N_7581,N_6079,N_6947);
nand U7582 (N_7582,N_6256,N_6947);
nand U7583 (N_7583,N_6789,N_6409);
or U7584 (N_7584,N_6719,N_6321);
xnor U7585 (N_7585,N_6542,N_6199);
nand U7586 (N_7586,N_6954,N_6110);
xor U7587 (N_7587,N_6844,N_6794);
nand U7588 (N_7588,N_6568,N_6553);
xnor U7589 (N_7589,N_6799,N_6588);
nor U7590 (N_7590,N_6674,N_6393);
xnor U7591 (N_7591,N_6008,N_6188);
nand U7592 (N_7592,N_6951,N_6327);
or U7593 (N_7593,N_6439,N_6468);
nor U7594 (N_7594,N_6777,N_6096);
nand U7595 (N_7595,N_6518,N_6730);
nand U7596 (N_7596,N_6244,N_6357);
nor U7597 (N_7597,N_6111,N_6386);
nand U7598 (N_7598,N_6770,N_6187);
and U7599 (N_7599,N_6347,N_6814);
or U7600 (N_7600,N_6664,N_6934);
nor U7601 (N_7601,N_6315,N_6502);
nor U7602 (N_7602,N_6996,N_6262);
and U7603 (N_7603,N_6797,N_6057);
and U7604 (N_7604,N_6762,N_6927);
nor U7605 (N_7605,N_6329,N_6876);
xnor U7606 (N_7606,N_6587,N_6621);
and U7607 (N_7607,N_6831,N_6236);
xor U7608 (N_7608,N_6270,N_6206);
and U7609 (N_7609,N_6353,N_6039);
xor U7610 (N_7610,N_6285,N_6877);
xnor U7611 (N_7611,N_6152,N_6630);
nor U7612 (N_7612,N_6971,N_6889);
nor U7613 (N_7613,N_6876,N_6233);
and U7614 (N_7614,N_6362,N_6424);
nor U7615 (N_7615,N_6974,N_6172);
or U7616 (N_7616,N_6292,N_6515);
xor U7617 (N_7617,N_6158,N_6002);
nor U7618 (N_7618,N_6571,N_6141);
and U7619 (N_7619,N_6135,N_6354);
or U7620 (N_7620,N_6163,N_6106);
xnor U7621 (N_7621,N_6119,N_6068);
nor U7622 (N_7622,N_6944,N_6900);
or U7623 (N_7623,N_6030,N_6560);
or U7624 (N_7624,N_6830,N_6626);
and U7625 (N_7625,N_6556,N_6873);
nand U7626 (N_7626,N_6655,N_6812);
xnor U7627 (N_7627,N_6372,N_6031);
xor U7628 (N_7628,N_6489,N_6838);
nand U7629 (N_7629,N_6379,N_6149);
xnor U7630 (N_7630,N_6415,N_6566);
xnor U7631 (N_7631,N_6134,N_6638);
or U7632 (N_7632,N_6581,N_6273);
or U7633 (N_7633,N_6285,N_6548);
nand U7634 (N_7634,N_6797,N_6101);
nand U7635 (N_7635,N_6185,N_6291);
nor U7636 (N_7636,N_6146,N_6451);
or U7637 (N_7637,N_6621,N_6798);
and U7638 (N_7638,N_6247,N_6322);
or U7639 (N_7639,N_6041,N_6391);
nor U7640 (N_7640,N_6877,N_6768);
xor U7641 (N_7641,N_6245,N_6762);
nand U7642 (N_7642,N_6383,N_6439);
nand U7643 (N_7643,N_6294,N_6789);
or U7644 (N_7644,N_6455,N_6480);
nor U7645 (N_7645,N_6393,N_6787);
or U7646 (N_7646,N_6863,N_6133);
nor U7647 (N_7647,N_6028,N_6369);
nand U7648 (N_7648,N_6746,N_6905);
or U7649 (N_7649,N_6738,N_6980);
and U7650 (N_7650,N_6813,N_6232);
nor U7651 (N_7651,N_6949,N_6064);
and U7652 (N_7652,N_6287,N_6407);
nand U7653 (N_7653,N_6620,N_6166);
xnor U7654 (N_7654,N_6234,N_6832);
and U7655 (N_7655,N_6231,N_6276);
nand U7656 (N_7656,N_6333,N_6471);
and U7657 (N_7657,N_6578,N_6981);
nand U7658 (N_7658,N_6164,N_6370);
nand U7659 (N_7659,N_6549,N_6633);
or U7660 (N_7660,N_6303,N_6977);
or U7661 (N_7661,N_6870,N_6616);
and U7662 (N_7662,N_6034,N_6546);
xnor U7663 (N_7663,N_6761,N_6182);
nor U7664 (N_7664,N_6385,N_6434);
and U7665 (N_7665,N_6799,N_6102);
xor U7666 (N_7666,N_6950,N_6283);
or U7667 (N_7667,N_6059,N_6295);
xor U7668 (N_7668,N_6089,N_6519);
and U7669 (N_7669,N_6861,N_6236);
or U7670 (N_7670,N_6331,N_6763);
or U7671 (N_7671,N_6013,N_6855);
nand U7672 (N_7672,N_6869,N_6189);
nand U7673 (N_7673,N_6841,N_6333);
and U7674 (N_7674,N_6970,N_6217);
and U7675 (N_7675,N_6938,N_6634);
xor U7676 (N_7676,N_6957,N_6716);
xnor U7677 (N_7677,N_6437,N_6358);
and U7678 (N_7678,N_6356,N_6621);
or U7679 (N_7679,N_6952,N_6511);
nor U7680 (N_7680,N_6961,N_6750);
or U7681 (N_7681,N_6258,N_6033);
nor U7682 (N_7682,N_6803,N_6658);
nor U7683 (N_7683,N_6042,N_6795);
and U7684 (N_7684,N_6015,N_6287);
nor U7685 (N_7685,N_6445,N_6828);
and U7686 (N_7686,N_6293,N_6262);
nor U7687 (N_7687,N_6671,N_6978);
xor U7688 (N_7688,N_6683,N_6709);
nor U7689 (N_7689,N_6171,N_6243);
xnor U7690 (N_7690,N_6846,N_6278);
xnor U7691 (N_7691,N_6447,N_6379);
or U7692 (N_7692,N_6449,N_6296);
or U7693 (N_7693,N_6954,N_6557);
nand U7694 (N_7694,N_6946,N_6207);
or U7695 (N_7695,N_6907,N_6395);
xor U7696 (N_7696,N_6801,N_6073);
nand U7697 (N_7697,N_6122,N_6702);
or U7698 (N_7698,N_6235,N_6773);
nor U7699 (N_7699,N_6357,N_6564);
nand U7700 (N_7700,N_6612,N_6972);
and U7701 (N_7701,N_6285,N_6053);
nand U7702 (N_7702,N_6240,N_6696);
xnor U7703 (N_7703,N_6559,N_6282);
and U7704 (N_7704,N_6310,N_6271);
or U7705 (N_7705,N_6240,N_6367);
nor U7706 (N_7706,N_6255,N_6290);
and U7707 (N_7707,N_6873,N_6083);
nand U7708 (N_7708,N_6292,N_6005);
nand U7709 (N_7709,N_6465,N_6026);
or U7710 (N_7710,N_6849,N_6275);
and U7711 (N_7711,N_6947,N_6494);
nor U7712 (N_7712,N_6727,N_6728);
or U7713 (N_7713,N_6686,N_6952);
and U7714 (N_7714,N_6051,N_6907);
and U7715 (N_7715,N_6527,N_6084);
or U7716 (N_7716,N_6273,N_6886);
and U7717 (N_7717,N_6456,N_6190);
and U7718 (N_7718,N_6304,N_6310);
nand U7719 (N_7719,N_6281,N_6974);
and U7720 (N_7720,N_6655,N_6553);
xnor U7721 (N_7721,N_6634,N_6024);
nor U7722 (N_7722,N_6362,N_6677);
nor U7723 (N_7723,N_6302,N_6663);
nand U7724 (N_7724,N_6742,N_6978);
or U7725 (N_7725,N_6707,N_6036);
and U7726 (N_7726,N_6045,N_6322);
nor U7727 (N_7727,N_6270,N_6631);
nor U7728 (N_7728,N_6888,N_6544);
nor U7729 (N_7729,N_6171,N_6319);
nand U7730 (N_7730,N_6885,N_6485);
and U7731 (N_7731,N_6486,N_6969);
or U7732 (N_7732,N_6106,N_6363);
or U7733 (N_7733,N_6990,N_6422);
and U7734 (N_7734,N_6931,N_6213);
nand U7735 (N_7735,N_6661,N_6360);
nor U7736 (N_7736,N_6765,N_6664);
and U7737 (N_7737,N_6250,N_6082);
or U7738 (N_7738,N_6360,N_6354);
or U7739 (N_7739,N_6995,N_6959);
nand U7740 (N_7740,N_6426,N_6300);
xor U7741 (N_7741,N_6435,N_6581);
nor U7742 (N_7742,N_6747,N_6285);
nor U7743 (N_7743,N_6169,N_6861);
and U7744 (N_7744,N_6418,N_6855);
or U7745 (N_7745,N_6472,N_6933);
nor U7746 (N_7746,N_6087,N_6960);
or U7747 (N_7747,N_6404,N_6168);
xor U7748 (N_7748,N_6350,N_6642);
or U7749 (N_7749,N_6425,N_6887);
and U7750 (N_7750,N_6593,N_6641);
and U7751 (N_7751,N_6464,N_6629);
or U7752 (N_7752,N_6830,N_6319);
xor U7753 (N_7753,N_6243,N_6633);
nand U7754 (N_7754,N_6029,N_6646);
and U7755 (N_7755,N_6362,N_6367);
nor U7756 (N_7756,N_6168,N_6099);
nand U7757 (N_7757,N_6819,N_6085);
nor U7758 (N_7758,N_6376,N_6025);
and U7759 (N_7759,N_6881,N_6240);
or U7760 (N_7760,N_6545,N_6407);
and U7761 (N_7761,N_6595,N_6081);
or U7762 (N_7762,N_6940,N_6713);
or U7763 (N_7763,N_6432,N_6337);
nand U7764 (N_7764,N_6039,N_6967);
and U7765 (N_7765,N_6920,N_6489);
xnor U7766 (N_7766,N_6937,N_6905);
nand U7767 (N_7767,N_6380,N_6719);
nand U7768 (N_7768,N_6583,N_6623);
xnor U7769 (N_7769,N_6997,N_6111);
nand U7770 (N_7770,N_6917,N_6414);
nand U7771 (N_7771,N_6639,N_6805);
xnor U7772 (N_7772,N_6056,N_6279);
xnor U7773 (N_7773,N_6798,N_6415);
nor U7774 (N_7774,N_6290,N_6120);
or U7775 (N_7775,N_6653,N_6044);
nor U7776 (N_7776,N_6125,N_6941);
nand U7777 (N_7777,N_6480,N_6754);
or U7778 (N_7778,N_6335,N_6057);
xnor U7779 (N_7779,N_6571,N_6751);
xor U7780 (N_7780,N_6241,N_6938);
nand U7781 (N_7781,N_6840,N_6460);
or U7782 (N_7782,N_6134,N_6747);
nor U7783 (N_7783,N_6556,N_6775);
or U7784 (N_7784,N_6050,N_6846);
xnor U7785 (N_7785,N_6939,N_6077);
and U7786 (N_7786,N_6928,N_6038);
and U7787 (N_7787,N_6169,N_6210);
nor U7788 (N_7788,N_6751,N_6650);
nand U7789 (N_7789,N_6276,N_6565);
or U7790 (N_7790,N_6227,N_6915);
and U7791 (N_7791,N_6239,N_6744);
or U7792 (N_7792,N_6186,N_6272);
or U7793 (N_7793,N_6860,N_6856);
xor U7794 (N_7794,N_6756,N_6551);
or U7795 (N_7795,N_6771,N_6052);
or U7796 (N_7796,N_6401,N_6159);
nor U7797 (N_7797,N_6026,N_6467);
nor U7798 (N_7798,N_6787,N_6469);
and U7799 (N_7799,N_6227,N_6558);
or U7800 (N_7800,N_6987,N_6268);
nand U7801 (N_7801,N_6644,N_6784);
or U7802 (N_7802,N_6054,N_6265);
xor U7803 (N_7803,N_6339,N_6598);
nor U7804 (N_7804,N_6121,N_6813);
nor U7805 (N_7805,N_6218,N_6285);
nor U7806 (N_7806,N_6651,N_6477);
xnor U7807 (N_7807,N_6802,N_6037);
or U7808 (N_7808,N_6068,N_6452);
and U7809 (N_7809,N_6060,N_6825);
or U7810 (N_7810,N_6114,N_6966);
xnor U7811 (N_7811,N_6326,N_6125);
or U7812 (N_7812,N_6605,N_6529);
and U7813 (N_7813,N_6608,N_6864);
nor U7814 (N_7814,N_6301,N_6916);
xor U7815 (N_7815,N_6245,N_6764);
nand U7816 (N_7816,N_6218,N_6396);
xnor U7817 (N_7817,N_6116,N_6722);
or U7818 (N_7818,N_6053,N_6226);
nor U7819 (N_7819,N_6349,N_6232);
and U7820 (N_7820,N_6960,N_6605);
xor U7821 (N_7821,N_6628,N_6723);
nor U7822 (N_7822,N_6419,N_6571);
nor U7823 (N_7823,N_6734,N_6175);
nor U7824 (N_7824,N_6781,N_6592);
or U7825 (N_7825,N_6086,N_6139);
nor U7826 (N_7826,N_6335,N_6272);
nand U7827 (N_7827,N_6726,N_6312);
xnor U7828 (N_7828,N_6542,N_6459);
nand U7829 (N_7829,N_6112,N_6967);
nor U7830 (N_7830,N_6139,N_6290);
nand U7831 (N_7831,N_6390,N_6318);
or U7832 (N_7832,N_6710,N_6069);
or U7833 (N_7833,N_6577,N_6180);
and U7834 (N_7834,N_6358,N_6228);
and U7835 (N_7835,N_6720,N_6318);
xor U7836 (N_7836,N_6064,N_6402);
nor U7837 (N_7837,N_6908,N_6932);
nand U7838 (N_7838,N_6046,N_6405);
nand U7839 (N_7839,N_6844,N_6126);
and U7840 (N_7840,N_6270,N_6752);
nand U7841 (N_7841,N_6728,N_6025);
nor U7842 (N_7842,N_6853,N_6233);
or U7843 (N_7843,N_6165,N_6766);
xor U7844 (N_7844,N_6717,N_6882);
and U7845 (N_7845,N_6645,N_6678);
nor U7846 (N_7846,N_6117,N_6926);
nor U7847 (N_7847,N_6402,N_6391);
or U7848 (N_7848,N_6776,N_6151);
or U7849 (N_7849,N_6918,N_6728);
and U7850 (N_7850,N_6525,N_6157);
xor U7851 (N_7851,N_6976,N_6353);
or U7852 (N_7852,N_6300,N_6840);
and U7853 (N_7853,N_6111,N_6783);
xor U7854 (N_7854,N_6310,N_6004);
or U7855 (N_7855,N_6936,N_6005);
nor U7856 (N_7856,N_6710,N_6825);
and U7857 (N_7857,N_6495,N_6441);
or U7858 (N_7858,N_6126,N_6432);
nand U7859 (N_7859,N_6736,N_6444);
or U7860 (N_7860,N_6543,N_6481);
xnor U7861 (N_7861,N_6579,N_6121);
or U7862 (N_7862,N_6211,N_6680);
or U7863 (N_7863,N_6277,N_6777);
and U7864 (N_7864,N_6733,N_6527);
nor U7865 (N_7865,N_6351,N_6095);
nand U7866 (N_7866,N_6623,N_6317);
nand U7867 (N_7867,N_6823,N_6034);
and U7868 (N_7868,N_6912,N_6840);
and U7869 (N_7869,N_6776,N_6853);
xor U7870 (N_7870,N_6361,N_6877);
or U7871 (N_7871,N_6205,N_6665);
nor U7872 (N_7872,N_6567,N_6756);
and U7873 (N_7873,N_6468,N_6901);
nand U7874 (N_7874,N_6545,N_6340);
or U7875 (N_7875,N_6383,N_6433);
or U7876 (N_7876,N_6408,N_6284);
nand U7877 (N_7877,N_6347,N_6733);
and U7878 (N_7878,N_6005,N_6214);
nor U7879 (N_7879,N_6671,N_6431);
or U7880 (N_7880,N_6402,N_6187);
and U7881 (N_7881,N_6848,N_6016);
nand U7882 (N_7882,N_6080,N_6932);
and U7883 (N_7883,N_6945,N_6283);
xnor U7884 (N_7884,N_6330,N_6894);
nor U7885 (N_7885,N_6861,N_6867);
nor U7886 (N_7886,N_6357,N_6028);
nor U7887 (N_7887,N_6195,N_6946);
and U7888 (N_7888,N_6441,N_6333);
nand U7889 (N_7889,N_6956,N_6159);
and U7890 (N_7890,N_6183,N_6801);
nor U7891 (N_7891,N_6384,N_6167);
nor U7892 (N_7892,N_6155,N_6046);
nor U7893 (N_7893,N_6942,N_6168);
and U7894 (N_7894,N_6300,N_6366);
and U7895 (N_7895,N_6510,N_6719);
nand U7896 (N_7896,N_6634,N_6448);
nand U7897 (N_7897,N_6328,N_6944);
nand U7898 (N_7898,N_6214,N_6417);
or U7899 (N_7899,N_6891,N_6580);
or U7900 (N_7900,N_6873,N_6839);
nand U7901 (N_7901,N_6331,N_6864);
or U7902 (N_7902,N_6926,N_6507);
nor U7903 (N_7903,N_6368,N_6390);
nand U7904 (N_7904,N_6953,N_6106);
or U7905 (N_7905,N_6906,N_6855);
or U7906 (N_7906,N_6178,N_6029);
nor U7907 (N_7907,N_6771,N_6200);
and U7908 (N_7908,N_6233,N_6507);
xor U7909 (N_7909,N_6619,N_6082);
nand U7910 (N_7910,N_6722,N_6806);
nand U7911 (N_7911,N_6844,N_6615);
nor U7912 (N_7912,N_6814,N_6676);
nor U7913 (N_7913,N_6073,N_6477);
nand U7914 (N_7914,N_6450,N_6548);
nand U7915 (N_7915,N_6138,N_6898);
and U7916 (N_7916,N_6927,N_6076);
xor U7917 (N_7917,N_6147,N_6160);
nor U7918 (N_7918,N_6908,N_6000);
nor U7919 (N_7919,N_6425,N_6464);
xor U7920 (N_7920,N_6162,N_6840);
xnor U7921 (N_7921,N_6537,N_6711);
and U7922 (N_7922,N_6068,N_6171);
nor U7923 (N_7923,N_6091,N_6940);
nand U7924 (N_7924,N_6108,N_6914);
or U7925 (N_7925,N_6323,N_6951);
nor U7926 (N_7926,N_6829,N_6132);
nor U7927 (N_7927,N_6122,N_6570);
nand U7928 (N_7928,N_6009,N_6233);
or U7929 (N_7929,N_6170,N_6541);
and U7930 (N_7930,N_6664,N_6609);
and U7931 (N_7931,N_6545,N_6985);
xor U7932 (N_7932,N_6582,N_6600);
nor U7933 (N_7933,N_6338,N_6419);
xnor U7934 (N_7934,N_6587,N_6581);
or U7935 (N_7935,N_6460,N_6612);
nand U7936 (N_7936,N_6535,N_6475);
or U7937 (N_7937,N_6381,N_6894);
nand U7938 (N_7938,N_6068,N_6954);
xnor U7939 (N_7939,N_6936,N_6116);
nand U7940 (N_7940,N_6760,N_6687);
nand U7941 (N_7941,N_6496,N_6551);
xor U7942 (N_7942,N_6687,N_6981);
xor U7943 (N_7943,N_6232,N_6487);
or U7944 (N_7944,N_6915,N_6049);
nand U7945 (N_7945,N_6901,N_6545);
nor U7946 (N_7946,N_6560,N_6631);
nand U7947 (N_7947,N_6949,N_6881);
and U7948 (N_7948,N_6210,N_6794);
xor U7949 (N_7949,N_6488,N_6587);
nor U7950 (N_7950,N_6761,N_6905);
xnor U7951 (N_7951,N_6492,N_6323);
and U7952 (N_7952,N_6002,N_6217);
xnor U7953 (N_7953,N_6321,N_6424);
nor U7954 (N_7954,N_6340,N_6336);
xor U7955 (N_7955,N_6407,N_6246);
xnor U7956 (N_7956,N_6042,N_6084);
xor U7957 (N_7957,N_6286,N_6215);
nand U7958 (N_7958,N_6521,N_6651);
nand U7959 (N_7959,N_6408,N_6330);
nand U7960 (N_7960,N_6867,N_6706);
nand U7961 (N_7961,N_6548,N_6639);
or U7962 (N_7962,N_6876,N_6858);
or U7963 (N_7963,N_6916,N_6582);
xnor U7964 (N_7964,N_6915,N_6398);
or U7965 (N_7965,N_6793,N_6025);
and U7966 (N_7966,N_6972,N_6559);
nand U7967 (N_7967,N_6322,N_6681);
or U7968 (N_7968,N_6811,N_6593);
and U7969 (N_7969,N_6291,N_6594);
or U7970 (N_7970,N_6083,N_6560);
nand U7971 (N_7971,N_6137,N_6965);
or U7972 (N_7972,N_6800,N_6598);
xnor U7973 (N_7973,N_6939,N_6072);
xnor U7974 (N_7974,N_6640,N_6877);
nand U7975 (N_7975,N_6356,N_6013);
xor U7976 (N_7976,N_6515,N_6091);
nor U7977 (N_7977,N_6735,N_6481);
and U7978 (N_7978,N_6745,N_6421);
or U7979 (N_7979,N_6422,N_6430);
xor U7980 (N_7980,N_6870,N_6006);
xor U7981 (N_7981,N_6678,N_6300);
nand U7982 (N_7982,N_6971,N_6765);
or U7983 (N_7983,N_6440,N_6855);
or U7984 (N_7984,N_6049,N_6382);
nor U7985 (N_7985,N_6398,N_6763);
xnor U7986 (N_7986,N_6504,N_6738);
nor U7987 (N_7987,N_6255,N_6679);
and U7988 (N_7988,N_6989,N_6840);
or U7989 (N_7989,N_6542,N_6127);
xnor U7990 (N_7990,N_6803,N_6017);
and U7991 (N_7991,N_6834,N_6599);
nand U7992 (N_7992,N_6988,N_6934);
nand U7993 (N_7993,N_6192,N_6087);
and U7994 (N_7994,N_6990,N_6270);
xnor U7995 (N_7995,N_6591,N_6277);
nand U7996 (N_7996,N_6000,N_6247);
xnor U7997 (N_7997,N_6484,N_6319);
nor U7998 (N_7998,N_6947,N_6109);
nand U7999 (N_7999,N_6854,N_6880);
xor U8000 (N_8000,N_7533,N_7182);
nor U8001 (N_8001,N_7609,N_7655);
and U8002 (N_8002,N_7314,N_7957);
nor U8003 (N_8003,N_7303,N_7376);
xor U8004 (N_8004,N_7174,N_7841);
nor U8005 (N_8005,N_7178,N_7317);
and U8006 (N_8006,N_7733,N_7944);
and U8007 (N_8007,N_7338,N_7346);
xor U8008 (N_8008,N_7834,N_7631);
or U8009 (N_8009,N_7591,N_7861);
and U8010 (N_8010,N_7054,N_7586);
nor U8011 (N_8011,N_7126,N_7752);
xnor U8012 (N_8012,N_7094,N_7941);
and U8013 (N_8013,N_7345,N_7385);
nor U8014 (N_8014,N_7565,N_7230);
and U8015 (N_8015,N_7813,N_7032);
nand U8016 (N_8016,N_7132,N_7811);
nor U8017 (N_8017,N_7500,N_7081);
or U8018 (N_8018,N_7577,N_7173);
and U8019 (N_8019,N_7075,N_7769);
and U8020 (N_8020,N_7724,N_7825);
xor U8021 (N_8021,N_7243,N_7730);
or U8022 (N_8022,N_7531,N_7862);
or U8023 (N_8023,N_7843,N_7904);
nor U8024 (N_8024,N_7845,N_7883);
xor U8025 (N_8025,N_7285,N_7473);
xnor U8026 (N_8026,N_7997,N_7229);
or U8027 (N_8027,N_7302,N_7183);
or U8028 (N_8028,N_7802,N_7538);
xnor U8029 (N_8029,N_7125,N_7495);
nand U8030 (N_8030,N_7606,N_7850);
or U8031 (N_8031,N_7751,N_7480);
nand U8032 (N_8032,N_7910,N_7693);
and U8033 (N_8033,N_7650,N_7152);
and U8034 (N_8034,N_7242,N_7912);
and U8035 (N_8035,N_7455,N_7366);
xor U8036 (N_8036,N_7378,N_7319);
or U8037 (N_8037,N_7857,N_7051);
and U8038 (N_8038,N_7206,N_7477);
nor U8039 (N_8039,N_7421,N_7307);
or U8040 (N_8040,N_7707,N_7170);
nand U8041 (N_8041,N_7049,N_7562);
xnor U8042 (N_8042,N_7914,N_7984);
xnor U8043 (N_8043,N_7444,N_7927);
xnor U8044 (N_8044,N_7062,N_7311);
xor U8045 (N_8045,N_7341,N_7466);
xnor U8046 (N_8046,N_7240,N_7250);
nor U8047 (N_8047,N_7484,N_7248);
and U8048 (N_8048,N_7731,N_7169);
and U8049 (N_8049,N_7375,N_7608);
nor U8050 (N_8050,N_7633,N_7624);
nand U8051 (N_8051,N_7387,N_7635);
nor U8052 (N_8052,N_7476,N_7095);
or U8053 (N_8053,N_7943,N_7982);
nor U8054 (N_8054,N_7419,N_7764);
or U8055 (N_8055,N_7232,N_7791);
nor U8056 (N_8056,N_7519,N_7024);
or U8057 (N_8057,N_7740,N_7467);
and U8058 (N_8058,N_7200,N_7969);
xnor U8059 (N_8059,N_7175,N_7975);
nand U8060 (N_8060,N_7705,N_7348);
nand U8061 (N_8061,N_7884,N_7530);
nor U8062 (N_8062,N_7603,N_7670);
nand U8063 (N_8063,N_7617,N_7691);
or U8064 (N_8064,N_7025,N_7507);
or U8065 (N_8065,N_7863,N_7185);
xnor U8066 (N_8066,N_7050,N_7921);
or U8067 (N_8067,N_7488,N_7765);
or U8068 (N_8068,N_7505,N_7795);
nor U8069 (N_8069,N_7454,N_7753);
or U8070 (N_8070,N_7499,N_7917);
and U8071 (N_8071,N_7715,N_7029);
nand U8072 (N_8072,N_7965,N_7677);
or U8073 (N_8073,N_7590,N_7153);
and U8074 (N_8074,N_7552,N_7047);
xnor U8075 (N_8075,N_7771,N_7865);
nor U8076 (N_8076,N_7363,N_7472);
xnor U8077 (N_8077,N_7461,N_7649);
nor U8078 (N_8078,N_7929,N_7402);
xnor U8079 (N_8079,N_7288,N_7393);
nor U8080 (N_8080,N_7675,N_7362);
and U8081 (N_8081,N_7384,N_7636);
and U8082 (N_8082,N_7607,N_7401);
xnor U8083 (N_8083,N_7414,N_7736);
nor U8084 (N_8084,N_7263,N_7322);
and U8085 (N_8085,N_7137,N_7760);
xnor U8086 (N_8086,N_7284,N_7560);
xnor U8087 (N_8087,N_7517,N_7339);
xor U8088 (N_8088,N_7293,N_7020);
nor U8089 (N_8089,N_7361,N_7864);
or U8090 (N_8090,N_7847,N_7221);
nand U8091 (N_8091,N_7459,N_7882);
xor U8092 (N_8092,N_7231,N_7115);
or U8093 (N_8093,N_7683,N_7329);
and U8094 (N_8094,N_7084,N_7852);
nor U8095 (N_8095,N_7349,N_7256);
nand U8096 (N_8096,N_7096,N_7888);
nand U8097 (N_8097,N_7934,N_7815);
and U8098 (N_8098,N_7604,N_7958);
nor U8099 (N_8099,N_7816,N_7810);
nor U8100 (N_8100,N_7754,N_7687);
and U8101 (N_8101,N_7161,N_7723);
nor U8102 (N_8102,N_7728,N_7732);
nor U8103 (N_8103,N_7891,N_7300);
nor U8104 (N_8104,N_7620,N_7721);
and U8105 (N_8105,N_7867,N_7437);
nor U8106 (N_8106,N_7201,N_7673);
nor U8107 (N_8107,N_7599,N_7144);
and U8108 (N_8108,N_7278,N_7973);
nand U8109 (N_8109,N_7305,N_7452);
nand U8110 (N_8110,N_7219,N_7108);
xor U8111 (N_8111,N_7798,N_7537);
and U8112 (N_8112,N_7199,N_7186);
and U8113 (N_8113,N_7298,N_7700);
and U8114 (N_8114,N_7514,N_7682);
nor U8115 (N_8115,N_7526,N_7093);
xor U8116 (N_8116,N_7669,N_7127);
nor U8117 (N_8117,N_7664,N_7475);
or U8118 (N_8118,N_7851,N_7744);
or U8119 (N_8119,N_7245,N_7748);
xnor U8120 (N_8120,N_7781,N_7897);
nand U8121 (N_8121,N_7309,N_7960);
and U8122 (N_8122,N_7171,N_7701);
and U8123 (N_8123,N_7805,N_7823);
nor U8124 (N_8124,N_7972,N_7438);
nand U8125 (N_8125,N_7907,N_7292);
nor U8126 (N_8126,N_7992,N_7622);
or U8127 (N_8127,N_7991,N_7674);
nor U8128 (N_8128,N_7660,N_7269);
nor U8129 (N_8129,N_7350,N_7112);
nand U8130 (N_8130,N_7895,N_7632);
or U8131 (N_8131,N_7038,N_7168);
nor U8132 (N_8132,N_7788,N_7198);
xor U8133 (N_8133,N_7812,N_7706);
nand U8134 (N_8134,N_7568,N_7540);
nor U8135 (N_8135,N_7177,N_7522);
nand U8136 (N_8136,N_7451,N_7786);
xnor U8137 (N_8137,N_7666,N_7896);
or U8138 (N_8138,N_7006,N_7511);
nand U8139 (N_8139,N_7352,N_7092);
and U8140 (N_8140,N_7592,N_7899);
nor U8141 (N_8141,N_7908,N_7262);
nand U8142 (N_8142,N_7353,N_7237);
xnor U8143 (N_8143,N_7064,N_7978);
nor U8144 (N_8144,N_7091,N_7058);
nand U8145 (N_8145,N_7315,N_7755);
xor U8146 (N_8146,N_7513,N_7116);
or U8147 (N_8147,N_7400,N_7432);
and U8148 (N_8148,N_7197,N_7770);
xor U8149 (N_8149,N_7986,N_7589);
and U8150 (N_8150,N_7931,N_7260);
nor U8151 (N_8151,N_7469,N_7313);
xnor U8152 (N_8152,N_7510,N_7195);
xor U8153 (N_8153,N_7840,N_7021);
nor U8154 (N_8154,N_7924,N_7312);
xor U8155 (N_8155,N_7061,N_7193);
or U8156 (N_8156,N_7903,N_7406);
nor U8157 (N_8157,N_7323,N_7842);
or U8158 (N_8158,N_7060,N_7139);
nor U8159 (N_8159,N_7685,N_7555);
nand U8160 (N_8160,N_7234,N_7779);
xnor U8161 (N_8161,N_7433,N_7690);
and U8162 (N_8162,N_7335,N_7704);
nor U8163 (N_8163,N_7397,N_7699);
xor U8164 (N_8164,N_7196,N_7915);
and U8165 (N_8165,N_7227,N_7324);
nor U8166 (N_8166,N_7386,N_7672);
nand U8167 (N_8167,N_7106,N_7023);
xnor U8168 (N_8168,N_7148,N_7493);
nor U8169 (N_8169,N_7642,N_7963);
and U8170 (N_8170,N_7228,N_7124);
nor U8171 (N_8171,N_7626,N_7483);
and U8172 (N_8172,N_7681,N_7113);
or U8173 (N_8173,N_7547,N_7184);
and U8174 (N_8174,N_7819,N_7207);
or U8175 (N_8175,N_7524,N_7948);
nor U8176 (N_8176,N_7297,N_7080);
or U8177 (N_8177,N_7950,N_7719);
nor U8178 (N_8178,N_7089,N_7370);
and U8179 (N_8179,N_7143,N_7016);
nand U8180 (N_8180,N_7103,N_7470);
nand U8181 (N_8181,N_7520,N_7057);
nand U8182 (N_8182,N_7282,N_7766);
nand U8183 (N_8183,N_7134,N_7775);
and U8184 (N_8184,N_7571,N_7518);
nor U8185 (N_8185,N_7615,N_7255);
nand U8186 (N_8186,N_7365,N_7749);
and U8187 (N_8187,N_7994,N_7588);
nand U8188 (N_8188,N_7928,N_7208);
or U8189 (N_8189,N_7980,N_7226);
nor U8190 (N_8190,N_7835,N_7501);
or U8191 (N_8191,N_7046,N_7878);
nor U8192 (N_8192,N_7176,N_7639);
xnor U8193 (N_8193,N_7031,N_7720);
or U8194 (N_8194,N_7133,N_7553);
or U8195 (N_8195,N_7368,N_7450);
nor U8196 (N_8196,N_7983,N_7120);
nor U8197 (N_8197,N_7964,N_7114);
or U8198 (N_8198,N_7745,N_7281);
nand U8199 (N_8199,N_7204,N_7926);
xor U8200 (N_8200,N_7100,N_7083);
xnor U8201 (N_8201,N_7532,N_7875);
nand U8202 (N_8202,N_7576,N_7778);
and U8203 (N_8203,N_7328,N_7504);
and U8204 (N_8204,N_7979,N_7703);
nor U8205 (N_8205,N_7308,N_7808);
nand U8206 (N_8206,N_7739,N_7034);
nand U8207 (N_8207,N_7102,N_7074);
and U8208 (N_8208,N_7695,N_7164);
nand U8209 (N_8209,N_7082,N_7462);
nand U8210 (N_8210,N_7015,N_7709);
or U8211 (N_8211,N_7162,N_7502);
nor U8212 (N_8212,N_7252,N_7310);
nor U8213 (N_8213,N_7254,N_7981);
and U8214 (N_8214,N_7267,N_7790);
or U8215 (N_8215,N_7383,N_7427);
nand U8216 (N_8216,N_7648,N_7913);
nand U8217 (N_8217,N_7217,N_7828);
xnor U8218 (N_8218,N_7056,N_7712);
and U8219 (N_8219,N_7489,N_7605);
or U8220 (N_8220,N_7342,N_7373);
nor U8221 (N_8221,N_7239,N_7203);
nor U8222 (N_8222,N_7004,N_7409);
nor U8223 (N_8223,N_7296,N_7920);
xnor U8224 (N_8224,N_7244,N_7716);
or U8225 (N_8225,N_7059,N_7990);
and U8226 (N_8226,N_7768,N_7246);
xnor U8227 (N_8227,N_7759,N_7824);
nor U8228 (N_8228,N_7391,N_7336);
xor U8229 (N_8229,N_7069,N_7253);
nand U8230 (N_8230,N_7952,N_7787);
xor U8231 (N_8231,N_7209,N_7377);
and U8232 (N_8232,N_7961,N_7151);
or U8233 (N_8233,N_7431,N_7192);
and U8234 (N_8234,N_7971,N_7128);
and U8235 (N_8235,N_7800,N_7333);
nor U8236 (N_8236,N_7688,N_7412);
and U8237 (N_8237,N_7619,N_7570);
nor U8238 (N_8238,N_7696,N_7838);
xnor U8239 (N_8239,N_7906,N_7018);
or U8240 (N_8240,N_7582,N_7130);
and U8241 (N_8241,N_7774,N_7848);
or U8242 (N_8242,N_7429,N_7596);
nand U8243 (N_8243,N_7694,N_7066);
and U8244 (N_8244,N_7894,N_7157);
or U8245 (N_8245,N_7053,N_7331);
and U8246 (N_8246,N_7548,N_7268);
xnor U8247 (N_8247,N_7601,N_7686);
xor U8248 (N_8248,N_7684,N_7154);
and U8249 (N_8249,N_7909,N_7276);
xor U8250 (N_8250,N_7541,N_7347);
and U8251 (N_8251,N_7970,N_7996);
and U8252 (N_8252,N_7564,N_7418);
and U8253 (N_8253,N_7535,N_7379);
nand U8254 (N_8254,N_7937,N_7354);
nand U8255 (N_8255,N_7408,N_7097);
nand U8256 (N_8256,N_7993,N_7726);
nand U8257 (N_8257,N_7616,N_7492);
xor U8258 (N_8258,N_7776,N_7612);
nor U8259 (N_8259,N_7249,N_7554);
nor U8260 (N_8260,N_7832,N_7792);
and U8261 (N_8261,N_7951,N_7073);
nand U8262 (N_8262,N_7423,N_7523);
nand U8263 (N_8263,N_7750,N_7238);
or U8264 (N_8264,N_7017,N_7529);
nor U8265 (N_8265,N_7039,N_7007);
or U8266 (N_8266,N_7998,N_7647);
nand U8267 (N_8267,N_7357,N_7597);
xor U8268 (N_8268,N_7035,N_7223);
nand U8269 (N_8269,N_7767,N_7141);
nand U8270 (N_8270,N_7509,N_7515);
nor U8271 (N_8271,N_7659,N_7773);
xnor U8272 (N_8272,N_7585,N_7900);
nor U8273 (N_8273,N_7536,N_7539);
xnor U8274 (N_8274,N_7123,N_7022);
nand U8275 (N_8275,N_7563,N_7918);
or U8276 (N_8276,N_7872,N_7135);
and U8277 (N_8277,N_7680,N_7698);
or U8278 (N_8278,N_7661,N_7241);
nand U8279 (N_8279,N_7708,N_7422);
nor U8280 (N_8280,N_7337,N_7945);
or U8281 (N_8281,N_7831,N_7689);
nand U8282 (N_8282,N_7901,N_7463);
nand U8283 (N_8283,N_7627,N_7205);
or U8284 (N_8284,N_7656,N_7777);
nor U8285 (N_8285,N_7321,N_7646);
xnor U8286 (N_8286,N_7413,N_7942);
xor U8287 (N_8287,N_7299,N_7099);
nand U8288 (N_8288,N_7257,N_7887);
nor U8289 (N_8289,N_7465,N_7118);
or U8290 (N_8290,N_7077,N_7938);
nand U8291 (N_8291,N_7692,N_7224);
or U8292 (N_8292,N_7940,N_7119);
and U8293 (N_8293,N_7014,N_7645);
xor U8294 (N_8294,N_7561,N_7420);
xor U8295 (N_8295,N_7294,N_7332);
nor U8296 (N_8296,N_7545,N_7654);
and U8297 (N_8297,N_7042,N_7140);
xnor U8298 (N_8298,N_7330,N_7725);
or U8299 (N_8299,N_7820,N_7155);
nor U8300 (N_8300,N_7559,N_7325);
nand U8301 (N_8301,N_7165,N_7233);
and U8302 (N_8302,N_7761,N_7985);
and U8303 (N_8303,N_7036,N_7210);
or U8304 (N_8304,N_7734,N_7251);
and U8305 (N_8305,N_7180,N_7638);
xor U8306 (N_8306,N_7033,N_7027);
nor U8307 (N_8307,N_7301,N_7999);
and U8308 (N_8308,N_7600,N_7542);
nor U8309 (N_8309,N_7079,N_7212);
nor U8310 (N_8310,N_7388,N_7274);
nand U8311 (N_8311,N_7220,N_7717);
and U8312 (N_8312,N_7403,N_7742);
nand U8313 (N_8313,N_7211,N_7922);
and U8314 (N_8314,N_7844,N_7735);
nor U8315 (N_8315,N_7762,N_7890);
or U8316 (N_8316,N_7512,N_7424);
and U8317 (N_8317,N_7265,N_7087);
or U8318 (N_8318,N_7453,N_7949);
nand U8319 (N_8319,N_7747,N_7052);
nor U8320 (N_8320,N_7111,N_7662);
and U8321 (N_8321,N_7356,N_7236);
or U8322 (N_8322,N_7086,N_7871);
or U8323 (N_8323,N_7959,N_7809);
nor U8324 (N_8324,N_7859,N_7471);
nor U8325 (N_8325,N_7578,N_7587);
or U8326 (N_8326,N_7546,N_7827);
xor U8327 (N_8327,N_7822,N_7486);
nand U8328 (N_8328,N_7078,N_7575);
xnor U8329 (N_8329,N_7923,N_7572);
xnor U8330 (N_8330,N_7187,N_7988);
nand U8331 (N_8331,N_7167,N_7722);
nor U8332 (N_8332,N_7885,N_7490);
nand U8333 (N_8333,N_7491,N_7002);
and U8334 (N_8334,N_7456,N_7028);
nand U8335 (N_8335,N_7458,N_7567);
nor U8336 (N_8336,N_7264,N_7351);
xor U8337 (N_8337,N_7625,N_7030);
and U8338 (N_8338,N_7737,N_7005);
nor U8339 (N_8339,N_7508,N_7574);
xnor U8340 (N_8340,N_7797,N_7291);
xor U8341 (N_8341,N_7886,N_7225);
xnor U8342 (N_8342,N_7644,N_7110);
xnor U8343 (N_8343,N_7068,N_7009);
or U8344 (N_8344,N_7447,N_7785);
nand U8345 (N_8345,N_7758,N_7496);
nor U8346 (N_8346,N_7369,N_7389);
and U8347 (N_8347,N_7594,N_7372);
xor U8348 (N_8348,N_7371,N_7037);
xnor U8349 (N_8349,N_7962,N_7320);
nand U8350 (N_8350,N_7479,N_7355);
xnor U8351 (N_8351,N_7714,N_7464);
nand U8352 (N_8352,N_7869,N_7435);
nand U8353 (N_8353,N_7498,N_7041);
xor U8354 (N_8354,N_7411,N_7191);
xor U8355 (N_8355,N_7602,N_7481);
nor U8356 (N_8356,N_7919,N_7107);
nor U8357 (N_8357,N_7849,N_7782);
and U8358 (N_8358,N_7806,N_7445);
and U8359 (N_8359,N_7287,N_7390);
nand U8360 (N_8360,N_7930,N_7892);
xor U8361 (N_8361,N_7697,N_7277);
xor U8362 (N_8362,N_7550,N_7954);
nor U8363 (N_8363,N_7327,N_7334);
nand U8364 (N_8364,N_7286,N_7131);
nor U8365 (N_8365,N_7449,N_7434);
and U8366 (N_8366,N_7428,N_7441);
nand U8367 (N_8367,N_7395,N_7189);
and U8368 (N_8368,N_7629,N_7836);
nand U8369 (N_8369,N_7266,N_7380);
xnor U8370 (N_8370,N_7573,N_7145);
nor U8371 (N_8371,N_7306,N_7156);
nor U8372 (N_8372,N_7671,N_7976);
xor U8373 (N_8373,N_7966,N_7868);
nor U8374 (N_8374,N_7794,N_7235);
xnor U8375 (N_8375,N_7190,N_7676);
nand U8376 (N_8376,N_7048,N_7663);
or U8377 (N_8377,N_7482,N_7398);
and U8378 (N_8378,N_7359,N_7902);
xor U8379 (N_8379,N_7595,N_7818);
and U8380 (N_8380,N_7989,N_7527);
nand U8381 (N_8381,N_7947,N_7067);
nor U8382 (N_8382,N_7783,N_7440);
nor U8383 (N_8383,N_7045,N_7702);
nand U8384 (N_8384,N_7415,N_7218);
nor U8385 (N_8385,N_7011,N_7874);
or U8386 (N_8386,N_7043,N_7146);
or U8387 (N_8387,N_7487,N_7967);
nand U8388 (N_8388,N_7381,N_7583);
nand U8389 (N_8389,N_7521,N_7630);
xor U8390 (N_8390,N_7544,N_7799);
nand U8391 (N_8391,N_7442,N_7407);
or U8392 (N_8392,N_7516,N_7668);
nand U8393 (N_8393,N_7261,N_7953);
and U8394 (N_8394,N_7443,N_7468);
xor U8395 (N_8395,N_7640,N_7090);
nand U8396 (N_8396,N_7893,N_7634);
xor U8397 (N_8397,N_7678,N_7405);
xor U8398 (N_8398,N_7935,N_7003);
nor U8399 (N_8399,N_7613,N_7713);
nor U8400 (N_8400,N_7977,N_7853);
and U8401 (N_8401,N_7598,N_7880);
or U8402 (N_8402,N_7641,N_7746);
nor U8403 (N_8403,N_7817,N_7122);
or U8404 (N_8404,N_7936,N_7417);
nor U8405 (N_8405,N_7340,N_7457);
nand U8406 (N_8406,N_7946,N_7101);
xnor U8407 (N_8407,N_7877,N_7399);
nand U8408 (N_8408,N_7566,N_7718);
xnor U8409 (N_8409,N_7304,N_7569);
nor U8410 (N_8410,N_7855,N_7525);
and U8411 (N_8411,N_7905,N_7044);
nand U8412 (N_8412,N_7757,N_7839);
nand U8413 (N_8413,N_7741,N_7793);
and U8414 (N_8414,N_7326,N_7055);
or U8415 (N_8415,N_7652,N_7814);
nor U8416 (N_8416,N_7729,N_7367);
or U8417 (N_8417,N_7665,N_7743);
and U8418 (N_8418,N_7803,N_7364);
xnor U8419 (N_8419,N_7129,N_7172);
nor U8420 (N_8420,N_7316,N_7343);
and U8421 (N_8421,N_7117,N_7593);
nand U8422 (N_8422,N_7202,N_7956);
and U8423 (N_8423,N_7436,N_7995);
or U8424 (N_8424,N_7866,N_7136);
or U8425 (N_8425,N_7711,N_7556);
xnor U8426 (N_8426,N_7933,N_7181);
nor U8427 (N_8427,N_7474,N_7846);
and U8428 (N_8428,N_7987,N_7179);
xnor U8429 (N_8429,N_7580,N_7833);
xnor U8430 (N_8430,N_7558,N_7222);
or U8431 (N_8431,N_7772,N_7149);
nor U8432 (N_8432,N_7088,N_7446);
and U8433 (N_8433,N_7109,N_7194);
xnor U8434 (N_8434,N_7679,N_7911);
and U8435 (N_8435,N_7460,N_7829);
or U8436 (N_8436,N_7826,N_7651);
or U8437 (N_8437,N_7040,N_7543);
nand U8438 (N_8438,N_7789,N_7534);
xor U8439 (N_8439,N_7968,N_7158);
and U8440 (N_8440,N_7280,N_7344);
or U8441 (N_8441,N_7780,N_7026);
or U8442 (N_8442,N_7854,N_7008);
xnor U8443 (N_8443,N_7925,N_7318);
nor U8444 (N_8444,N_7653,N_7150);
or U8445 (N_8445,N_7485,N_7098);
nand U8446 (N_8446,N_7410,N_7283);
or U8447 (N_8447,N_7142,N_7939);
nand U8448 (N_8448,N_7621,N_7667);
or U8449 (N_8449,N_7497,N_7738);
or U8450 (N_8450,N_7166,N_7275);
or U8451 (N_8451,N_7494,N_7860);
nor U8452 (N_8452,N_7270,N_7289);
xor U8453 (N_8453,N_7070,N_7549);
or U8454 (N_8454,N_7358,N_7727);
xor U8455 (N_8455,N_7614,N_7528);
xor U8456 (N_8456,N_7643,N_7657);
nor U8457 (N_8457,N_7796,N_7801);
nor U8458 (N_8458,N_7404,N_7756);
nand U8459 (N_8459,N_7856,N_7974);
xnor U8460 (N_8460,N_7439,N_7858);
and U8461 (N_8461,N_7821,N_7076);
and U8462 (N_8462,N_7360,N_7710);
nor U8463 (N_8463,N_7581,N_7396);
or U8464 (N_8464,N_7147,N_7163);
and U8465 (N_8465,N_7898,N_7628);
and U8466 (N_8466,N_7272,N_7271);
xor U8467 (N_8467,N_7105,N_7214);
nor U8468 (N_8468,N_7273,N_7121);
or U8469 (N_8469,N_7215,N_7012);
xor U8470 (N_8470,N_7584,N_7426);
and U8471 (N_8471,N_7104,N_7279);
nand U8472 (N_8472,N_7506,N_7295);
xnor U8473 (N_8473,N_7579,N_7448);
or U8474 (N_8474,N_7955,N_7932);
and U8475 (N_8475,N_7430,N_7159);
and U8476 (N_8476,N_7478,N_7138);
or U8477 (N_8477,N_7394,N_7830);
nand U8478 (N_8478,N_7010,N_7072);
or U8479 (N_8479,N_7870,N_7259);
xor U8480 (N_8480,N_7085,N_7557);
nand U8481 (N_8481,N_7889,N_7065);
or U8482 (N_8482,N_7916,N_7216);
xnor U8483 (N_8483,N_7382,N_7551);
or U8484 (N_8484,N_7019,N_7881);
xor U8485 (N_8485,N_7610,N_7000);
and U8486 (N_8486,N_7416,N_7618);
nand U8487 (N_8487,N_7188,N_7213);
and U8488 (N_8488,N_7611,N_7876);
nand U8489 (N_8489,N_7013,N_7392);
or U8490 (N_8490,N_7160,N_7873);
nand U8491 (N_8491,N_7763,N_7784);
or U8492 (N_8492,N_7658,N_7637);
nand U8493 (N_8493,N_7837,N_7063);
nor U8494 (N_8494,N_7503,N_7374);
or U8495 (N_8495,N_7247,N_7807);
nand U8496 (N_8496,N_7425,N_7290);
or U8497 (N_8497,N_7804,N_7001);
xor U8498 (N_8498,N_7071,N_7623);
or U8499 (N_8499,N_7258,N_7879);
nand U8500 (N_8500,N_7804,N_7770);
nor U8501 (N_8501,N_7807,N_7616);
nand U8502 (N_8502,N_7649,N_7782);
xor U8503 (N_8503,N_7603,N_7780);
or U8504 (N_8504,N_7707,N_7234);
nand U8505 (N_8505,N_7905,N_7967);
xnor U8506 (N_8506,N_7302,N_7287);
and U8507 (N_8507,N_7302,N_7687);
or U8508 (N_8508,N_7055,N_7284);
xor U8509 (N_8509,N_7156,N_7034);
and U8510 (N_8510,N_7697,N_7984);
xnor U8511 (N_8511,N_7257,N_7756);
or U8512 (N_8512,N_7249,N_7584);
nand U8513 (N_8513,N_7214,N_7498);
nor U8514 (N_8514,N_7533,N_7440);
nor U8515 (N_8515,N_7669,N_7136);
xor U8516 (N_8516,N_7946,N_7179);
nor U8517 (N_8517,N_7060,N_7610);
nand U8518 (N_8518,N_7042,N_7604);
and U8519 (N_8519,N_7396,N_7390);
or U8520 (N_8520,N_7155,N_7942);
nor U8521 (N_8521,N_7427,N_7818);
xnor U8522 (N_8522,N_7195,N_7386);
nand U8523 (N_8523,N_7951,N_7800);
nor U8524 (N_8524,N_7653,N_7180);
nor U8525 (N_8525,N_7453,N_7976);
xnor U8526 (N_8526,N_7277,N_7766);
nor U8527 (N_8527,N_7690,N_7460);
nor U8528 (N_8528,N_7110,N_7585);
and U8529 (N_8529,N_7187,N_7404);
xor U8530 (N_8530,N_7393,N_7153);
nand U8531 (N_8531,N_7106,N_7779);
or U8532 (N_8532,N_7251,N_7375);
nand U8533 (N_8533,N_7537,N_7020);
xor U8534 (N_8534,N_7484,N_7319);
nor U8535 (N_8535,N_7496,N_7307);
or U8536 (N_8536,N_7620,N_7169);
nor U8537 (N_8537,N_7627,N_7197);
xnor U8538 (N_8538,N_7016,N_7588);
and U8539 (N_8539,N_7212,N_7272);
xnor U8540 (N_8540,N_7265,N_7142);
xor U8541 (N_8541,N_7071,N_7966);
or U8542 (N_8542,N_7297,N_7393);
nand U8543 (N_8543,N_7440,N_7564);
or U8544 (N_8544,N_7776,N_7788);
xor U8545 (N_8545,N_7751,N_7162);
and U8546 (N_8546,N_7769,N_7292);
nor U8547 (N_8547,N_7803,N_7734);
or U8548 (N_8548,N_7610,N_7638);
xor U8549 (N_8549,N_7643,N_7455);
nand U8550 (N_8550,N_7344,N_7218);
nand U8551 (N_8551,N_7097,N_7101);
nand U8552 (N_8552,N_7881,N_7830);
nor U8553 (N_8553,N_7549,N_7100);
xor U8554 (N_8554,N_7522,N_7471);
and U8555 (N_8555,N_7649,N_7114);
nand U8556 (N_8556,N_7310,N_7492);
or U8557 (N_8557,N_7567,N_7160);
nand U8558 (N_8558,N_7319,N_7045);
nand U8559 (N_8559,N_7939,N_7765);
and U8560 (N_8560,N_7934,N_7440);
nand U8561 (N_8561,N_7097,N_7644);
nor U8562 (N_8562,N_7392,N_7320);
nor U8563 (N_8563,N_7799,N_7229);
or U8564 (N_8564,N_7680,N_7096);
nand U8565 (N_8565,N_7620,N_7474);
nand U8566 (N_8566,N_7404,N_7794);
nor U8567 (N_8567,N_7328,N_7013);
nand U8568 (N_8568,N_7044,N_7059);
xor U8569 (N_8569,N_7361,N_7330);
xor U8570 (N_8570,N_7795,N_7808);
nand U8571 (N_8571,N_7412,N_7916);
or U8572 (N_8572,N_7310,N_7266);
nor U8573 (N_8573,N_7624,N_7294);
xnor U8574 (N_8574,N_7154,N_7772);
or U8575 (N_8575,N_7098,N_7174);
and U8576 (N_8576,N_7369,N_7319);
nor U8577 (N_8577,N_7379,N_7397);
and U8578 (N_8578,N_7763,N_7431);
xnor U8579 (N_8579,N_7578,N_7803);
xor U8580 (N_8580,N_7394,N_7727);
or U8581 (N_8581,N_7795,N_7877);
xor U8582 (N_8582,N_7661,N_7006);
and U8583 (N_8583,N_7713,N_7628);
or U8584 (N_8584,N_7180,N_7807);
nor U8585 (N_8585,N_7019,N_7275);
nor U8586 (N_8586,N_7399,N_7884);
nor U8587 (N_8587,N_7991,N_7364);
nor U8588 (N_8588,N_7980,N_7816);
xor U8589 (N_8589,N_7056,N_7511);
and U8590 (N_8590,N_7837,N_7106);
and U8591 (N_8591,N_7112,N_7421);
or U8592 (N_8592,N_7334,N_7929);
xnor U8593 (N_8593,N_7748,N_7970);
nand U8594 (N_8594,N_7960,N_7816);
nand U8595 (N_8595,N_7338,N_7994);
or U8596 (N_8596,N_7757,N_7360);
or U8597 (N_8597,N_7386,N_7458);
and U8598 (N_8598,N_7453,N_7914);
xnor U8599 (N_8599,N_7305,N_7097);
xnor U8600 (N_8600,N_7716,N_7972);
nor U8601 (N_8601,N_7975,N_7346);
and U8602 (N_8602,N_7972,N_7435);
xor U8603 (N_8603,N_7436,N_7210);
xor U8604 (N_8604,N_7129,N_7358);
xnor U8605 (N_8605,N_7945,N_7305);
nor U8606 (N_8606,N_7130,N_7008);
nand U8607 (N_8607,N_7682,N_7124);
and U8608 (N_8608,N_7534,N_7054);
and U8609 (N_8609,N_7341,N_7936);
or U8610 (N_8610,N_7409,N_7282);
and U8611 (N_8611,N_7986,N_7408);
and U8612 (N_8612,N_7391,N_7101);
nor U8613 (N_8613,N_7498,N_7459);
and U8614 (N_8614,N_7666,N_7977);
xor U8615 (N_8615,N_7661,N_7239);
nand U8616 (N_8616,N_7514,N_7987);
and U8617 (N_8617,N_7128,N_7589);
and U8618 (N_8618,N_7296,N_7017);
nor U8619 (N_8619,N_7552,N_7907);
nor U8620 (N_8620,N_7536,N_7789);
nand U8621 (N_8621,N_7043,N_7932);
xor U8622 (N_8622,N_7343,N_7624);
xor U8623 (N_8623,N_7294,N_7143);
nand U8624 (N_8624,N_7782,N_7133);
and U8625 (N_8625,N_7371,N_7680);
nand U8626 (N_8626,N_7147,N_7463);
nand U8627 (N_8627,N_7844,N_7826);
and U8628 (N_8628,N_7994,N_7436);
xor U8629 (N_8629,N_7707,N_7214);
nor U8630 (N_8630,N_7557,N_7871);
and U8631 (N_8631,N_7603,N_7050);
nand U8632 (N_8632,N_7598,N_7112);
nand U8633 (N_8633,N_7914,N_7810);
or U8634 (N_8634,N_7538,N_7449);
nand U8635 (N_8635,N_7585,N_7998);
nor U8636 (N_8636,N_7083,N_7327);
xnor U8637 (N_8637,N_7704,N_7023);
or U8638 (N_8638,N_7142,N_7761);
xnor U8639 (N_8639,N_7160,N_7022);
nor U8640 (N_8640,N_7732,N_7069);
nor U8641 (N_8641,N_7181,N_7371);
nor U8642 (N_8642,N_7633,N_7278);
nand U8643 (N_8643,N_7907,N_7306);
nand U8644 (N_8644,N_7522,N_7771);
nand U8645 (N_8645,N_7189,N_7975);
and U8646 (N_8646,N_7157,N_7282);
nand U8647 (N_8647,N_7843,N_7498);
nor U8648 (N_8648,N_7335,N_7065);
nor U8649 (N_8649,N_7807,N_7289);
or U8650 (N_8650,N_7042,N_7116);
xnor U8651 (N_8651,N_7259,N_7385);
xor U8652 (N_8652,N_7003,N_7608);
or U8653 (N_8653,N_7469,N_7515);
and U8654 (N_8654,N_7384,N_7895);
xor U8655 (N_8655,N_7803,N_7728);
and U8656 (N_8656,N_7000,N_7520);
or U8657 (N_8657,N_7909,N_7555);
and U8658 (N_8658,N_7159,N_7942);
nor U8659 (N_8659,N_7994,N_7437);
and U8660 (N_8660,N_7843,N_7491);
or U8661 (N_8661,N_7074,N_7793);
xnor U8662 (N_8662,N_7644,N_7256);
and U8663 (N_8663,N_7140,N_7775);
and U8664 (N_8664,N_7127,N_7988);
nand U8665 (N_8665,N_7166,N_7997);
or U8666 (N_8666,N_7087,N_7052);
or U8667 (N_8667,N_7330,N_7193);
and U8668 (N_8668,N_7893,N_7112);
xor U8669 (N_8669,N_7573,N_7014);
or U8670 (N_8670,N_7308,N_7257);
and U8671 (N_8671,N_7647,N_7192);
xor U8672 (N_8672,N_7179,N_7022);
and U8673 (N_8673,N_7151,N_7470);
or U8674 (N_8674,N_7832,N_7685);
nand U8675 (N_8675,N_7258,N_7764);
nand U8676 (N_8676,N_7829,N_7935);
xor U8677 (N_8677,N_7408,N_7295);
nand U8678 (N_8678,N_7510,N_7769);
xnor U8679 (N_8679,N_7838,N_7665);
or U8680 (N_8680,N_7237,N_7647);
or U8681 (N_8681,N_7276,N_7304);
xnor U8682 (N_8682,N_7429,N_7639);
nand U8683 (N_8683,N_7924,N_7024);
nand U8684 (N_8684,N_7696,N_7625);
nor U8685 (N_8685,N_7926,N_7861);
xnor U8686 (N_8686,N_7124,N_7245);
xor U8687 (N_8687,N_7457,N_7145);
or U8688 (N_8688,N_7895,N_7820);
nor U8689 (N_8689,N_7490,N_7655);
or U8690 (N_8690,N_7445,N_7353);
and U8691 (N_8691,N_7568,N_7865);
and U8692 (N_8692,N_7308,N_7683);
and U8693 (N_8693,N_7238,N_7333);
or U8694 (N_8694,N_7856,N_7307);
nor U8695 (N_8695,N_7532,N_7297);
nor U8696 (N_8696,N_7153,N_7336);
and U8697 (N_8697,N_7151,N_7327);
nor U8698 (N_8698,N_7595,N_7772);
xor U8699 (N_8699,N_7385,N_7226);
xor U8700 (N_8700,N_7364,N_7432);
nor U8701 (N_8701,N_7025,N_7418);
or U8702 (N_8702,N_7563,N_7265);
xnor U8703 (N_8703,N_7489,N_7801);
nand U8704 (N_8704,N_7758,N_7557);
nand U8705 (N_8705,N_7924,N_7447);
nor U8706 (N_8706,N_7461,N_7351);
xnor U8707 (N_8707,N_7167,N_7677);
and U8708 (N_8708,N_7847,N_7541);
xnor U8709 (N_8709,N_7536,N_7481);
and U8710 (N_8710,N_7821,N_7813);
or U8711 (N_8711,N_7887,N_7057);
nor U8712 (N_8712,N_7488,N_7517);
or U8713 (N_8713,N_7180,N_7272);
xor U8714 (N_8714,N_7051,N_7984);
nor U8715 (N_8715,N_7446,N_7396);
nor U8716 (N_8716,N_7467,N_7553);
or U8717 (N_8717,N_7814,N_7276);
or U8718 (N_8718,N_7988,N_7133);
and U8719 (N_8719,N_7532,N_7918);
nand U8720 (N_8720,N_7596,N_7314);
and U8721 (N_8721,N_7549,N_7931);
nand U8722 (N_8722,N_7633,N_7982);
nand U8723 (N_8723,N_7004,N_7571);
xor U8724 (N_8724,N_7972,N_7336);
or U8725 (N_8725,N_7216,N_7464);
xor U8726 (N_8726,N_7424,N_7592);
xnor U8727 (N_8727,N_7935,N_7738);
or U8728 (N_8728,N_7013,N_7974);
xnor U8729 (N_8729,N_7541,N_7207);
nand U8730 (N_8730,N_7732,N_7150);
or U8731 (N_8731,N_7597,N_7193);
nand U8732 (N_8732,N_7000,N_7938);
nand U8733 (N_8733,N_7824,N_7365);
xnor U8734 (N_8734,N_7288,N_7781);
xnor U8735 (N_8735,N_7850,N_7073);
or U8736 (N_8736,N_7160,N_7689);
or U8737 (N_8737,N_7207,N_7060);
nand U8738 (N_8738,N_7980,N_7896);
xnor U8739 (N_8739,N_7805,N_7428);
nand U8740 (N_8740,N_7891,N_7842);
and U8741 (N_8741,N_7163,N_7351);
nand U8742 (N_8742,N_7510,N_7461);
nand U8743 (N_8743,N_7835,N_7701);
nand U8744 (N_8744,N_7817,N_7822);
nand U8745 (N_8745,N_7682,N_7732);
or U8746 (N_8746,N_7287,N_7237);
or U8747 (N_8747,N_7876,N_7379);
or U8748 (N_8748,N_7148,N_7826);
nor U8749 (N_8749,N_7504,N_7487);
xnor U8750 (N_8750,N_7403,N_7697);
xor U8751 (N_8751,N_7327,N_7026);
nand U8752 (N_8752,N_7066,N_7561);
nor U8753 (N_8753,N_7024,N_7865);
and U8754 (N_8754,N_7915,N_7688);
nand U8755 (N_8755,N_7634,N_7194);
or U8756 (N_8756,N_7907,N_7641);
and U8757 (N_8757,N_7970,N_7184);
nor U8758 (N_8758,N_7647,N_7365);
xnor U8759 (N_8759,N_7501,N_7807);
nor U8760 (N_8760,N_7428,N_7740);
nor U8761 (N_8761,N_7578,N_7201);
or U8762 (N_8762,N_7382,N_7599);
or U8763 (N_8763,N_7456,N_7406);
and U8764 (N_8764,N_7172,N_7038);
or U8765 (N_8765,N_7456,N_7818);
or U8766 (N_8766,N_7168,N_7196);
nor U8767 (N_8767,N_7282,N_7303);
nor U8768 (N_8768,N_7648,N_7252);
or U8769 (N_8769,N_7364,N_7602);
nor U8770 (N_8770,N_7842,N_7732);
and U8771 (N_8771,N_7242,N_7925);
xor U8772 (N_8772,N_7625,N_7334);
or U8773 (N_8773,N_7822,N_7628);
xnor U8774 (N_8774,N_7582,N_7685);
xor U8775 (N_8775,N_7219,N_7658);
xnor U8776 (N_8776,N_7007,N_7013);
nand U8777 (N_8777,N_7488,N_7542);
nand U8778 (N_8778,N_7193,N_7164);
xnor U8779 (N_8779,N_7016,N_7380);
or U8780 (N_8780,N_7939,N_7864);
nor U8781 (N_8781,N_7436,N_7252);
xor U8782 (N_8782,N_7232,N_7940);
xnor U8783 (N_8783,N_7137,N_7966);
nor U8784 (N_8784,N_7479,N_7865);
or U8785 (N_8785,N_7677,N_7139);
or U8786 (N_8786,N_7577,N_7738);
xor U8787 (N_8787,N_7413,N_7304);
nor U8788 (N_8788,N_7724,N_7650);
nor U8789 (N_8789,N_7998,N_7299);
nor U8790 (N_8790,N_7427,N_7691);
nand U8791 (N_8791,N_7571,N_7457);
and U8792 (N_8792,N_7290,N_7770);
nand U8793 (N_8793,N_7829,N_7017);
or U8794 (N_8794,N_7489,N_7776);
or U8795 (N_8795,N_7503,N_7020);
nand U8796 (N_8796,N_7227,N_7946);
xnor U8797 (N_8797,N_7586,N_7085);
nor U8798 (N_8798,N_7488,N_7957);
nand U8799 (N_8799,N_7018,N_7572);
nor U8800 (N_8800,N_7121,N_7438);
or U8801 (N_8801,N_7961,N_7551);
nand U8802 (N_8802,N_7404,N_7488);
nand U8803 (N_8803,N_7937,N_7646);
nor U8804 (N_8804,N_7001,N_7496);
and U8805 (N_8805,N_7066,N_7640);
nor U8806 (N_8806,N_7003,N_7271);
nand U8807 (N_8807,N_7605,N_7911);
or U8808 (N_8808,N_7878,N_7250);
nor U8809 (N_8809,N_7491,N_7715);
or U8810 (N_8810,N_7399,N_7827);
and U8811 (N_8811,N_7980,N_7681);
xnor U8812 (N_8812,N_7584,N_7463);
xnor U8813 (N_8813,N_7905,N_7396);
and U8814 (N_8814,N_7998,N_7924);
nor U8815 (N_8815,N_7724,N_7940);
or U8816 (N_8816,N_7205,N_7043);
or U8817 (N_8817,N_7328,N_7252);
or U8818 (N_8818,N_7925,N_7913);
or U8819 (N_8819,N_7438,N_7627);
nand U8820 (N_8820,N_7702,N_7803);
xor U8821 (N_8821,N_7957,N_7541);
nor U8822 (N_8822,N_7920,N_7793);
or U8823 (N_8823,N_7330,N_7881);
nor U8824 (N_8824,N_7507,N_7707);
or U8825 (N_8825,N_7551,N_7581);
or U8826 (N_8826,N_7892,N_7924);
or U8827 (N_8827,N_7471,N_7112);
xor U8828 (N_8828,N_7967,N_7499);
and U8829 (N_8829,N_7311,N_7820);
xor U8830 (N_8830,N_7320,N_7620);
nor U8831 (N_8831,N_7515,N_7354);
xor U8832 (N_8832,N_7061,N_7746);
nor U8833 (N_8833,N_7470,N_7057);
nand U8834 (N_8834,N_7487,N_7932);
or U8835 (N_8835,N_7112,N_7763);
xor U8836 (N_8836,N_7205,N_7744);
xor U8837 (N_8837,N_7578,N_7821);
and U8838 (N_8838,N_7811,N_7228);
nand U8839 (N_8839,N_7093,N_7360);
and U8840 (N_8840,N_7121,N_7848);
and U8841 (N_8841,N_7467,N_7145);
xor U8842 (N_8842,N_7271,N_7291);
nor U8843 (N_8843,N_7908,N_7207);
nor U8844 (N_8844,N_7311,N_7665);
nand U8845 (N_8845,N_7690,N_7288);
and U8846 (N_8846,N_7624,N_7162);
nand U8847 (N_8847,N_7251,N_7491);
xor U8848 (N_8848,N_7386,N_7125);
nand U8849 (N_8849,N_7616,N_7020);
nor U8850 (N_8850,N_7806,N_7128);
nand U8851 (N_8851,N_7206,N_7413);
and U8852 (N_8852,N_7962,N_7484);
nand U8853 (N_8853,N_7308,N_7164);
nand U8854 (N_8854,N_7786,N_7519);
xor U8855 (N_8855,N_7475,N_7738);
and U8856 (N_8856,N_7605,N_7318);
nor U8857 (N_8857,N_7273,N_7239);
xnor U8858 (N_8858,N_7995,N_7377);
or U8859 (N_8859,N_7116,N_7668);
nor U8860 (N_8860,N_7423,N_7756);
and U8861 (N_8861,N_7360,N_7156);
nor U8862 (N_8862,N_7387,N_7605);
nand U8863 (N_8863,N_7189,N_7248);
or U8864 (N_8864,N_7877,N_7764);
xor U8865 (N_8865,N_7359,N_7922);
nor U8866 (N_8866,N_7976,N_7009);
nor U8867 (N_8867,N_7274,N_7598);
nand U8868 (N_8868,N_7082,N_7524);
or U8869 (N_8869,N_7242,N_7013);
and U8870 (N_8870,N_7334,N_7651);
xor U8871 (N_8871,N_7360,N_7915);
or U8872 (N_8872,N_7818,N_7875);
and U8873 (N_8873,N_7473,N_7712);
xor U8874 (N_8874,N_7496,N_7334);
and U8875 (N_8875,N_7029,N_7707);
and U8876 (N_8876,N_7592,N_7105);
and U8877 (N_8877,N_7253,N_7304);
nand U8878 (N_8878,N_7816,N_7569);
xor U8879 (N_8879,N_7548,N_7955);
or U8880 (N_8880,N_7561,N_7244);
or U8881 (N_8881,N_7846,N_7273);
nand U8882 (N_8882,N_7579,N_7738);
nand U8883 (N_8883,N_7634,N_7881);
xor U8884 (N_8884,N_7123,N_7603);
or U8885 (N_8885,N_7902,N_7635);
nand U8886 (N_8886,N_7357,N_7748);
nor U8887 (N_8887,N_7635,N_7063);
xor U8888 (N_8888,N_7129,N_7953);
and U8889 (N_8889,N_7789,N_7371);
xor U8890 (N_8890,N_7354,N_7400);
nand U8891 (N_8891,N_7952,N_7028);
nor U8892 (N_8892,N_7176,N_7183);
xor U8893 (N_8893,N_7999,N_7415);
xnor U8894 (N_8894,N_7942,N_7621);
nor U8895 (N_8895,N_7605,N_7359);
xor U8896 (N_8896,N_7660,N_7206);
or U8897 (N_8897,N_7606,N_7540);
nor U8898 (N_8898,N_7604,N_7974);
nor U8899 (N_8899,N_7371,N_7354);
or U8900 (N_8900,N_7772,N_7491);
xnor U8901 (N_8901,N_7384,N_7673);
nand U8902 (N_8902,N_7138,N_7811);
nand U8903 (N_8903,N_7786,N_7189);
xor U8904 (N_8904,N_7671,N_7703);
or U8905 (N_8905,N_7651,N_7540);
and U8906 (N_8906,N_7408,N_7855);
and U8907 (N_8907,N_7661,N_7875);
and U8908 (N_8908,N_7185,N_7683);
and U8909 (N_8909,N_7292,N_7075);
or U8910 (N_8910,N_7620,N_7513);
nand U8911 (N_8911,N_7870,N_7409);
xnor U8912 (N_8912,N_7584,N_7011);
and U8913 (N_8913,N_7691,N_7842);
nand U8914 (N_8914,N_7601,N_7102);
xor U8915 (N_8915,N_7533,N_7169);
nor U8916 (N_8916,N_7544,N_7374);
xor U8917 (N_8917,N_7145,N_7504);
or U8918 (N_8918,N_7829,N_7760);
nor U8919 (N_8919,N_7377,N_7607);
xnor U8920 (N_8920,N_7946,N_7113);
and U8921 (N_8921,N_7805,N_7766);
nor U8922 (N_8922,N_7357,N_7581);
and U8923 (N_8923,N_7373,N_7638);
nand U8924 (N_8924,N_7581,N_7042);
xor U8925 (N_8925,N_7346,N_7610);
nor U8926 (N_8926,N_7694,N_7683);
nor U8927 (N_8927,N_7784,N_7372);
nand U8928 (N_8928,N_7712,N_7581);
or U8929 (N_8929,N_7837,N_7385);
or U8930 (N_8930,N_7902,N_7000);
or U8931 (N_8931,N_7793,N_7642);
or U8932 (N_8932,N_7315,N_7061);
xnor U8933 (N_8933,N_7195,N_7930);
and U8934 (N_8934,N_7679,N_7984);
nor U8935 (N_8935,N_7848,N_7174);
nand U8936 (N_8936,N_7259,N_7862);
xnor U8937 (N_8937,N_7283,N_7585);
nor U8938 (N_8938,N_7005,N_7400);
nor U8939 (N_8939,N_7572,N_7187);
or U8940 (N_8940,N_7365,N_7192);
nor U8941 (N_8941,N_7927,N_7960);
or U8942 (N_8942,N_7007,N_7392);
and U8943 (N_8943,N_7848,N_7002);
and U8944 (N_8944,N_7510,N_7885);
xnor U8945 (N_8945,N_7749,N_7541);
nor U8946 (N_8946,N_7314,N_7578);
and U8947 (N_8947,N_7462,N_7796);
nor U8948 (N_8948,N_7206,N_7929);
xor U8949 (N_8949,N_7747,N_7849);
nor U8950 (N_8950,N_7613,N_7943);
xnor U8951 (N_8951,N_7417,N_7797);
nor U8952 (N_8952,N_7314,N_7127);
and U8953 (N_8953,N_7428,N_7290);
nand U8954 (N_8954,N_7838,N_7100);
nor U8955 (N_8955,N_7684,N_7211);
or U8956 (N_8956,N_7602,N_7012);
nor U8957 (N_8957,N_7969,N_7265);
or U8958 (N_8958,N_7137,N_7355);
nor U8959 (N_8959,N_7044,N_7495);
nand U8960 (N_8960,N_7948,N_7889);
nor U8961 (N_8961,N_7544,N_7481);
or U8962 (N_8962,N_7646,N_7171);
nand U8963 (N_8963,N_7516,N_7714);
xor U8964 (N_8964,N_7267,N_7563);
xnor U8965 (N_8965,N_7085,N_7529);
and U8966 (N_8966,N_7088,N_7368);
and U8967 (N_8967,N_7739,N_7297);
and U8968 (N_8968,N_7096,N_7422);
nor U8969 (N_8969,N_7343,N_7553);
xnor U8970 (N_8970,N_7134,N_7672);
nor U8971 (N_8971,N_7665,N_7022);
and U8972 (N_8972,N_7711,N_7000);
and U8973 (N_8973,N_7957,N_7696);
nor U8974 (N_8974,N_7768,N_7618);
nand U8975 (N_8975,N_7089,N_7481);
or U8976 (N_8976,N_7865,N_7415);
nor U8977 (N_8977,N_7946,N_7713);
nor U8978 (N_8978,N_7293,N_7390);
xor U8979 (N_8979,N_7902,N_7083);
nor U8980 (N_8980,N_7767,N_7699);
or U8981 (N_8981,N_7456,N_7982);
nor U8982 (N_8982,N_7171,N_7652);
or U8983 (N_8983,N_7655,N_7007);
nand U8984 (N_8984,N_7521,N_7024);
and U8985 (N_8985,N_7763,N_7752);
nor U8986 (N_8986,N_7056,N_7546);
or U8987 (N_8987,N_7938,N_7260);
and U8988 (N_8988,N_7283,N_7581);
and U8989 (N_8989,N_7577,N_7584);
or U8990 (N_8990,N_7194,N_7374);
xnor U8991 (N_8991,N_7455,N_7998);
and U8992 (N_8992,N_7431,N_7766);
or U8993 (N_8993,N_7434,N_7534);
xor U8994 (N_8994,N_7140,N_7157);
xnor U8995 (N_8995,N_7988,N_7619);
nand U8996 (N_8996,N_7474,N_7549);
xnor U8997 (N_8997,N_7600,N_7284);
or U8998 (N_8998,N_7947,N_7074);
and U8999 (N_8999,N_7320,N_7132);
and U9000 (N_9000,N_8007,N_8712);
and U9001 (N_9001,N_8137,N_8512);
nand U9002 (N_9002,N_8290,N_8126);
nand U9003 (N_9003,N_8501,N_8513);
and U9004 (N_9004,N_8106,N_8220);
and U9005 (N_9005,N_8689,N_8688);
or U9006 (N_9006,N_8066,N_8603);
and U9007 (N_9007,N_8541,N_8910);
xor U9008 (N_9008,N_8895,N_8870);
or U9009 (N_9009,N_8468,N_8619);
nand U9010 (N_9010,N_8620,N_8476);
nand U9011 (N_9011,N_8558,N_8314);
xor U9012 (N_9012,N_8877,N_8426);
xor U9013 (N_9013,N_8643,N_8112);
nor U9014 (N_9014,N_8103,N_8294);
nand U9015 (N_9015,N_8746,N_8592);
or U9016 (N_9016,N_8141,N_8665);
and U9017 (N_9017,N_8334,N_8146);
or U9018 (N_9018,N_8824,N_8660);
or U9019 (N_9019,N_8659,N_8523);
nand U9020 (N_9020,N_8219,N_8439);
nand U9021 (N_9021,N_8390,N_8804);
nor U9022 (N_9022,N_8424,N_8559);
and U9023 (N_9023,N_8863,N_8122);
xor U9024 (N_9024,N_8465,N_8196);
and U9025 (N_9025,N_8125,N_8860);
xnor U9026 (N_9026,N_8456,N_8254);
nor U9027 (N_9027,N_8675,N_8599);
and U9028 (N_9028,N_8186,N_8736);
or U9029 (N_9029,N_8449,N_8943);
and U9030 (N_9030,N_8886,N_8401);
nor U9031 (N_9031,N_8145,N_8790);
and U9032 (N_9032,N_8434,N_8792);
nand U9033 (N_9033,N_8964,N_8984);
and U9034 (N_9034,N_8742,N_8772);
nand U9035 (N_9035,N_8621,N_8887);
and U9036 (N_9036,N_8636,N_8349);
nor U9037 (N_9037,N_8844,N_8306);
or U9038 (N_9038,N_8394,N_8857);
and U9039 (N_9039,N_8816,N_8990);
or U9040 (N_9040,N_8545,N_8717);
and U9041 (N_9041,N_8515,N_8041);
or U9042 (N_9042,N_8276,N_8068);
xnor U9043 (N_9043,N_8738,N_8817);
and U9044 (N_9044,N_8261,N_8960);
and U9045 (N_9045,N_8775,N_8312);
nor U9046 (N_9046,N_8319,N_8562);
and U9047 (N_9047,N_8819,N_8947);
and U9048 (N_9048,N_8427,N_8575);
nand U9049 (N_9049,N_8134,N_8307);
or U9050 (N_9050,N_8783,N_8295);
or U9051 (N_9051,N_8030,N_8168);
nor U9052 (N_9052,N_8358,N_8693);
nor U9053 (N_9053,N_8798,N_8357);
nand U9054 (N_9054,N_8705,N_8935);
or U9055 (N_9055,N_8520,N_8001);
and U9056 (N_9056,N_8104,N_8799);
nor U9057 (N_9057,N_8078,N_8518);
and U9058 (N_9058,N_8878,N_8566);
xnor U9059 (N_9059,N_8521,N_8360);
xnor U9060 (N_9060,N_8152,N_8876);
nand U9061 (N_9061,N_8371,N_8789);
or U9062 (N_9062,N_8653,N_8179);
or U9063 (N_9063,N_8377,N_8040);
and U9064 (N_9064,N_8242,N_8215);
and U9065 (N_9065,N_8634,N_8206);
nor U9066 (N_9066,N_8011,N_8998);
xnor U9067 (N_9067,N_8904,N_8210);
nand U9068 (N_9068,N_8542,N_8346);
and U9069 (N_9069,N_8847,N_8241);
xnor U9070 (N_9070,N_8576,N_8669);
xnor U9071 (N_9071,N_8353,N_8631);
nor U9072 (N_9072,N_8662,N_8075);
xnor U9073 (N_9073,N_8709,N_8683);
xnor U9074 (N_9074,N_8671,N_8996);
nor U9075 (N_9075,N_8667,N_8815);
nor U9076 (N_9076,N_8065,N_8114);
xor U9077 (N_9077,N_8766,N_8590);
nand U9078 (N_9078,N_8869,N_8664);
nand U9079 (N_9079,N_8282,N_8980);
and U9080 (N_9080,N_8005,N_8999);
and U9081 (N_9081,N_8981,N_8063);
nor U9082 (N_9082,N_8135,N_8684);
or U9083 (N_9083,N_8555,N_8781);
or U9084 (N_9084,N_8837,N_8931);
or U9085 (N_9085,N_8718,N_8691);
and U9086 (N_9086,N_8916,N_8605);
or U9087 (N_9087,N_8893,N_8187);
and U9088 (N_9088,N_8280,N_8822);
nor U9089 (N_9089,N_8796,N_8383);
nand U9090 (N_9090,N_8949,N_8052);
and U9091 (N_9091,N_8406,N_8903);
nand U9092 (N_9092,N_8909,N_8800);
or U9093 (N_9093,N_8900,N_8354);
nand U9094 (N_9094,N_8431,N_8169);
nor U9095 (N_9095,N_8247,N_8164);
and U9096 (N_9096,N_8938,N_8258);
nor U9097 (N_9097,N_8674,N_8047);
and U9098 (N_9098,N_8534,N_8986);
and U9099 (N_9099,N_8514,N_8531);
xnor U9100 (N_9100,N_8832,N_8277);
and U9101 (N_9101,N_8079,N_8739);
or U9102 (N_9102,N_8069,N_8271);
xnor U9103 (N_9103,N_8754,N_8230);
or U9104 (N_9104,N_8029,N_8611);
nor U9105 (N_9105,N_8922,N_8447);
nand U9106 (N_9106,N_8330,N_8544);
and U9107 (N_9107,N_8151,N_8706);
and U9108 (N_9108,N_8711,N_8504);
and U9109 (N_9109,N_8823,N_8630);
nand U9110 (N_9110,N_8036,N_8726);
xnor U9111 (N_9111,N_8156,N_8745);
and U9112 (N_9112,N_8661,N_8749);
xnor U9113 (N_9113,N_8255,N_8451);
nor U9114 (N_9114,N_8090,N_8213);
xor U9115 (N_9115,N_8563,N_8171);
and U9116 (N_9116,N_8509,N_8647);
or U9117 (N_9117,N_8948,N_8853);
nor U9118 (N_9118,N_8296,N_8919);
or U9119 (N_9119,N_8490,N_8583);
nand U9120 (N_9120,N_8205,N_8627);
and U9121 (N_9121,N_8245,N_8238);
and U9122 (N_9122,N_8233,N_8160);
xnor U9123 (N_9123,N_8912,N_8644);
or U9124 (N_9124,N_8037,N_8459);
nor U9125 (N_9125,N_8725,N_8564);
nor U9126 (N_9126,N_8951,N_8226);
nor U9127 (N_9127,N_8686,N_8430);
nor U9128 (N_9128,N_8232,N_8682);
nor U9129 (N_9129,N_8941,N_8764);
nor U9130 (N_9130,N_8281,N_8510);
and U9131 (N_9131,N_8157,N_8165);
and U9132 (N_9132,N_8535,N_8582);
or U9133 (N_9133,N_8622,N_8017);
nand U9134 (N_9134,N_8496,N_8687);
or U9135 (N_9135,N_8851,N_8864);
xnor U9136 (N_9136,N_8410,N_8082);
nor U9137 (N_9137,N_8801,N_8194);
or U9138 (N_9138,N_8928,N_8148);
nor U9139 (N_9139,N_8379,N_8552);
or U9140 (N_9140,N_8142,N_8761);
xor U9141 (N_9141,N_8498,N_8652);
nor U9142 (N_9142,N_8568,N_8989);
and U9143 (N_9143,N_8607,N_8975);
nor U9144 (N_9144,N_8797,N_8362);
xor U9145 (N_9145,N_8757,N_8888);
xor U9146 (N_9146,N_8364,N_8820);
xnor U9147 (N_9147,N_8778,N_8250);
xnor U9148 (N_9148,N_8884,N_8366);
and U9149 (N_9149,N_8270,N_8855);
xor U9150 (N_9150,N_8750,N_8656);
nor U9151 (N_9151,N_8429,N_8010);
or U9152 (N_9152,N_8972,N_8291);
xnor U9153 (N_9153,N_8163,N_8715);
xor U9154 (N_9154,N_8861,N_8225);
nor U9155 (N_9155,N_8043,N_8388);
or U9156 (N_9156,N_8483,N_8901);
nand U9157 (N_9157,N_8987,N_8601);
xnor U9158 (N_9158,N_8409,N_8615);
and U9159 (N_9159,N_8180,N_8032);
or U9160 (N_9160,N_8214,N_8486);
or U9161 (N_9161,N_8256,N_8785);
nor U9162 (N_9162,N_8111,N_8119);
xnor U9163 (N_9163,N_8042,N_8985);
or U9164 (N_9164,N_8272,N_8842);
nor U9165 (N_9165,N_8421,N_8262);
nor U9166 (N_9166,N_8774,N_8556);
nand U9167 (N_9167,N_8899,N_8529);
nand U9168 (N_9168,N_8392,N_8204);
nand U9169 (N_9169,N_8020,N_8056);
nor U9170 (N_9170,N_8500,N_8086);
and U9171 (N_9171,N_8051,N_8301);
and U9172 (N_9172,N_8059,N_8672);
nand U9173 (N_9173,N_8110,N_8978);
nand U9174 (N_9174,N_8062,N_8268);
or U9175 (N_9175,N_8532,N_8329);
and U9176 (N_9176,N_8932,N_8172);
nand U9177 (N_9177,N_8002,N_8965);
nor U9178 (N_9178,N_8993,N_8199);
and U9179 (N_9179,N_8829,N_8979);
nor U9180 (N_9180,N_8216,N_8067);
nor U9181 (N_9181,N_8095,N_8517);
xor U9182 (N_9182,N_8298,N_8218);
and U9183 (N_9183,N_8278,N_8389);
xor U9184 (N_9184,N_8403,N_8419);
or U9185 (N_9185,N_8707,N_8162);
nor U9186 (N_9186,N_8791,N_8629);
xor U9187 (N_9187,N_8963,N_8311);
or U9188 (N_9188,N_8848,N_8257);
xnor U9189 (N_9189,N_8641,N_8317);
nor U9190 (N_9190,N_8628,N_8028);
nor U9191 (N_9191,N_8463,N_8417);
nand U9192 (N_9192,N_8759,N_8839);
xor U9193 (N_9193,N_8516,N_8253);
or U9194 (N_9194,N_8954,N_8604);
nor U9195 (N_9195,N_8109,N_8957);
nor U9196 (N_9196,N_8795,N_8956);
xnor U9197 (N_9197,N_8868,N_8655);
nand U9198 (N_9198,N_8344,N_8033);
or U9199 (N_9199,N_8006,N_8885);
or U9200 (N_9200,N_8663,N_8339);
xnor U9201 (N_9201,N_8175,N_8201);
and U9202 (N_9202,N_8805,N_8098);
xnor U9203 (N_9203,N_8335,N_8915);
xor U9204 (N_9204,N_8769,N_8983);
xnor U9205 (N_9205,N_8991,N_8573);
xnor U9206 (N_9206,N_8438,N_8473);
nor U9207 (N_9207,N_8115,N_8747);
nor U9208 (N_9208,N_8753,N_8658);
nor U9209 (N_9209,N_8748,N_8012);
xor U9210 (N_9210,N_8588,N_8359);
and U9211 (N_9211,N_8154,N_8091);
nor U9212 (N_9212,N_8235,N_8026);
or U9213 (N_9213,N_8391,N_8913);
nor U9214 (N_9214,N_8945,N_8466);
and U9215 (N_9215,N_8279,N_8879);
and U9216 (N_9216,N_8287,N_8246);
or U9217 (N_9217,N_8616,N_8679);
or U9218 (N_9218,N_8549,N_8461);
or U9219 (N_9219,N_8714,N_8713);
nor U9220 (N_9220,N_8762,N_8321);
or U9221 (N_9221,N_8740,N_8132);
or U9222 (N_9222,N_8347,N_8153);
and U9223 (N_9223,N_8898,N_8374);
nand U9224 (N_9224,N_8807,N_8252);
and U9225 (N_9225,N_8297,N_8835);
xor U9226 (N_9226,N_8070,N_8474);
xor U9227 (N_9227,N_8144,N_8120);
nand U9228 (N_9228,N_8440,N_8399);
and U9229 (N_9229,N_8131,N_8015);
xnor U9230 (N_9230,N_8966,N_8458);
or U9231 (N_9231,N_8578,N_8177);
or U9232 (N_9232,N_8944,N_8891);
and U9233 (N_9233,N_8589,N_8591);
and U9234 (N_9234,N_8397,N_8836);
xnor U9235 (N_9235,N_8872,N_8393);
and U9236 (N_9236,N_8786,N_8969);
and U9237 (N_9237,N_8982,N_8955);
and U9238 (N_9238,N_8727,N_8721);
xnor U9239 (N_9239,N_8690,N_8997);
nand U9240 (N_9240,N_8814,N_8914);
and U9241 (N_9241,N_8923,N_8022);
nor U9242 (N_9242,N_8019,N_8387);
xor U9243 (N_9243,N_8097,N_8973);
or U9244 (N_9244,N_8405,N_8570);
xnor U9245 (N_9245,N_8696,N_8341);
nor U9246 (N_9246,N_8723,N_8074);
and U9247 (N_9247,N_8318,N_8170);
and U9248 (N_9248,N_8720,N_8854);
or U9249 (N_9249,N_8402,N_8755);
nand U9250 (N_9250,N_8849,N_8994);
and U9251 (N_9251,N_8093,N_8380);
nor U9252 (N_9252,N_8569,N_8737);
nor U9253 (N_9253,N_8767,N_8927);
xnor U9254 (N_9254,N_8480,N_8046);
xor U9255 (N_9255,N_8827,N_8055);
nand U9256 (N_9256,N_8875,N_8333);
nand U9257 (N_9257,N_8852,N_8009);
and U9258 (N_9258,N_8049,N_8073);
and U9259 (N_9259,N_8124,N_8651);
xor U9260 (N_9260,N_8072,N_8600);
and U9261 (N_9261,N_8522,N_8018);
xnor U9262 (N_9262,N_8765,N_8231);
nand U9263 (N_9263,N_8100,N_8004);
or U9264 (N_9264,N_8053,N_8299);
nor U9265 (N_9265,N_8203,N_8221);
nor U9266 (N_9266,N_8929,N_8760);
and U9267 (N_9267,N_8489,N_8937);
or U9268 (N_9268,N_8084,N_8469);
nand U9269 (N_9269,N_8833,N_8952);
nand U9270 (N_9270,N_8743,N_8236);
and U9271 (N_9271,N_8442,N_8127);
xnor U9272 (N_9272,N_8361,N_8701);
nor U9273 (N_9273,N_8788,N_8382);
nand U9274 (N_9274,N_8161,N_8096);
or U9275 (N_9275,N_8525,N_8441);
or U9276 (N_9276,N_8475,N_8167);
xnor U9277 (N_9277,N_8071,N_8326);
nor U9278 (N_9278,N_8099,N_8492);
nand U9279 (N_9279,N_8654,N_8471);
nor U9280 (N_9280,N_8495,N_8905);
nor U9281 (N_9281,N_8728,N_8585);
nor U9282 (N_9282,N_8593,N_8327);
nand U9283 (N_9283,N_8284,N_8064);
nand U9284 (N_9284,N_8034,N_8770);
or U9285 (N_9285,N_8497,N_8692);
and U9286 (N_9286,N_8646,N_8894);
or U9287 (N_9287,N_8060,N_8414);
nor U9288 (N_9288,N_8025,N_8195);
nor U9289 (N_9289,N_8453,N_8618);
nand U9290 (N_9290,N_8435,N_8208);
or U9291 (N_9291,N_8251,N_8130);
xor U9292 (N_9292,N_8702,N_8027);
or U9293 (N_9293,N_8560,N_8303);
nand U9294 (N_9294,N_8638,N_8117);
xor U9295 (N_9295,N_8524,N_8176);
and U9296 (N_9296,N_8088,N_8315);
xnor U9297 (N_9297,N_8462,N_8094);
or U9298 (N_9298,N_8264,N_8337);
or U9299 (N_9299,N_8035,N_8023);
nor U9300 (N_9300,N_8472,N_8386);
or U9301 (N_9301,N_8266,N_8433);
nor U9302 (N_9302,N_8880,N_8376);
nor U9303 (N_9303,N_8087,N_8484);
xnor U9304 (N_9304,N_8645,N_8336);
xor U9305 (N_9305,N_8408,N_8331);
nor U9306 (N_9306,N_8540,N_8609);
and U9307 (N_9307,N_8602,N_8198);
or U9308 (N_9308,N_8967,N_8794);
nor U9309 (N_9309,N_8340,N_8508);
and U9310 (N_9310,N_8356,N_8313);
nand U9311 (N_9311,N_8077,N_8862);
and U9312 (N_9312,N_8464,N_8921);
nand U9313 (N_9313,N_8649,N_8384);
or U9314 (N_9314,N_8874,N_8274);
xor U9315 (N_9315,N_8507,N_8482);
nor U9316 (N_9316,N_8812,N_8673);
nand U9317 (N_9317,N_8116,N_8437);
nand U9318 (N_9318,N_8809,N_8565);
or U9319 (N_9319,N_8428,N_8906);
or U9320 (N_9320,N_8273,N_8918);
or U9321 (N_9321,N_8808,N_8352);
or U9322 (N_9322,N_8606,N_8302);
nor U9323 (N_9323,N_8048,N_8806);
or U9324 (N_9324,N_8722,N_8460);
xnor U9325 (N_9325,N_8971,N_8443);
nor U9326 (N_9326,N_8933,N_8803);
nor U9327 (N_9327,N_8625,N_8581);
or U9328 (N_9328,N_8958,N_8639);
and U9329 (N_9329,N_8128,N_8320);
nand U9330 (N_9330,N_8724,N_8940);
xor U9331 (N_9331,N_8348,N_8719);
nand U9332 (N_9332,N_8793,N_8821);
xor U9333 (N_9333,N_8092,N_8838);
xor U9334 (N_9334,N_8123,N_8396);
xor U9335 (N_9335,N_8085,N_8873);
or U9336 (N_9336,N_8452,N_8189);
nor U9337 (N_9337,N_8557,N_8289);
xor U9338 (N_9338,N_8548,N_8446);
nand U9339 (N_9339,N_8102,N_8666);
nand U9340 (N_9340,N_8547,N_8735);
and U9341 (N_9341,N_8398,N_8533);
nand U9342 (N_9342,N_8248,N_8732);
xnor U9343 (N_9343,N_8478,N_8670);
or U9344 (N_9344,N_8866,N_8269);
and U9345 (N_9345,N_8704,N_8676);
nand U9346 (N_9346,N_8351,N_8946);
or U9347 (N_9347,N_8200,N_8411);
nor U9348 (N_9348,N_8695,N_8328);
nor U9349 (N_9349,N_8703,N_8920);
and U9350 (N_9350,N_8181,N_8892);
or U9351 (N_9351,N_8917,N_8197);
nand U9352 (N_9352,N_8239,N_8595);
and U9353 (N_9353,N_8538,N_8355);
or U9354 (N_9354,N_8418,N_8243);
nand U9355 (N_9355,N_8890,N_8897);
nor U9356 (N_9356,N_8924,N_8716);
and U9357 (N_9357,N_8050,N_8267);
or U9358 (N_9358,N_8155,N_8343);
or U9359 (N_9359,N_8528,N_8694);
nand U9360 (N_9360,N_8404,N_8292);
nand U9361 (N_9361,N_8322,N_8561);
and U9362 (N_9362,N_8567,N_8378);
and U9363 (N_9363,N_8422,N_8977);
nand U9364 (N_9364,N_8623,N_8211);
xnor U9365 (N_9365,N_8741,N_8734);
or U9366 (N_9366,N_8249,N_8229);
nand U9367 (N_9367,N_8626,N_8385);
and U9368 (N_9368,N_8288,N_8038);
or U9369 (N_9369,N_8485,N_8223);
or U9370 (N_9370,N_8502,N_8519);
nand U9371 (N_9371,N_8310,N_8150);
xor U9372 (N_9372,N_8685,N_8858);
and U9373 (N_9373,N_8598,N_8217);
or U9374 (N_9374,N_8584,N_8436);
nand U9375 (N_9375,N_8416,N_8420);
xnor U9376 (N_9376,N_8014,N_8147);
or U9377 (N_9377,N_8058,N_8698);
xnor U9378 (N_9378,N_8237,N_8637);
xnor U9379 (N_9379,N_8970,N_8448);
and U9380 (N_9380,N_8285,N_8190);
and U9381 (N_9381,N_8024,N_8974);
nand U9382 (N_9382,N_8577,N_8697);
and U9383 (N_9383,N_8286,N_8871);
nand U9384 (N_9384,N_8784,N_8499);
or U9385 (N_9385,N_8733,N_8304);
nor U9386 (N_9386,N_8744,N_8503);
and U9387 (N_9387,N_8608,N_8939);
nand U9388 (N_9388,N_8061,N_8587);
nor U9389 (N_9389,N_8551,N_8423);
xor U9390 (N_9390,N_8612,N_8959);
nand U9391 (N_9391,N_8222,N_8536);
and U9392 (N_9392,N_8368,N_8305);
xor U9393 (N_9393,N_8107,N_8710);
xor U9394 (N_9394,N_8491,N_8202);
nand U9395 (N_9395,N_8140,N_8526);
nand U9396 (N_9396,N_8412,N_8158);
and U9397 (N_9397,N_8826,N_8907);
or U9398 (N_9398,N_8166,N_8045);
and U9399 (N_9399,N_8457,N_8081);
nor U9400 (N_9400,N_8228,N_8080);
nand U9401 (N_9401,N_8992,N_8934);
nor U9402 (N_9402,N_8013,N_8425);
nand U9403 (N_9403,N_8730,N_8136);
xor U9404 (N_9404,N_8293,N_8381);
nor U9405 (N_9405,N_8811,N_8942);
and U9406 (N_9406,N_8108,N_8481);
and U9407 (N_9407,N_8976,N_8260);
nand U9408 (N_9408,N_8192,N_8830);
nand U9409 (N_9409,N_8700,N_8968);
xor U9410 (N_9410,N_8375,N_8756);
nand U9411 (N_9411,N_8632,N_8908);
nand U9412 (N_9412,N_8118,N_8139);
xnor U9413 (N_9413,N_8083,N_8834);
xnor U9414 (N_9414,N_8859,N_8207);
nor U9415 (N_9415,N_8773,N_8610);
nor U9416 (N_9416,N_8624,N_8574);
nand U9417 (N_9417,N_8454,N_8962);
and U9418 (N_9418,N_8044,N_8370);
nor U9419 (N_9419,N_8530,N_8263);
nor U9420 (N_9420,N_8003,N_8546);
and U9421 (N_9421,N_8184,N_8596);
nand U9422 (N_9422,N_8613,N_8185);
nand U9423 (N_9423,N_8089,N_8537);
xnor U9424 (N_9424,N_8283,N_8057);
or U9425 (N_9425,N_8494,N_8432);
or U9426 (N_9426,N_8450,N_8648);
or U9427 (N_9427,N_8902,N_8810);
nor U9428 (N_9428,N_8149,N_8961);
or U9429 (N_9429,N_8527,N_8455);
nor U9430 (N_9430,N_8758,N_8777);
xnor U9431 (N_9431,N_8493,N_8677);
or U9432 (N_9432,N_8586,N_8309);
nor U9433 (N_9433,N_8244,N_8678);
xor U9434 (N_9434,N_8597,N_8543);
nand U9435 (N_9435,N_8768,N_8445);
nor U9436 (N_9436,N_8182,N_8867);
xnor U9437 (N_9437,N_8550,N_8444);
nor U9438 (N_9438,N_8642,N_8259);
xnor U9439 (N_9439,N_8325,N_8787);
and U9440 (N_9440,N_8174,N_8731);
and U9441 (N_9441,N_8988,N_8300);
or U9442 (N_9442,N_8553,N_8771);
and U9443 (N_9443,N_8668,N_8400);
nor U9444 (N_9444,N_8138,N_8227);
nand U9445 (N_9445,N_8479,N_8209);
xor U9446 (N_9446,N_8372,N_8413);
nand U9447 (N_9447,N_8039,N_8580);
or U9448 (N_9448,N_8752,N_8212);
nor U9449 (N_9449,N_8021,N_8594);
nor U9450 (N_9450,N_8571,N_8159);
nor U9451 (N_9451,N_8845,N_8308);
nand U9452 (N_9452,N_8173,N_8825);
and U9453 (N_9453,N_8617,N_8572);
nor U9454 (N_9454,N_8316,N_8345);
xnor U9455 (N_9455,N_8143,N_8802);
and U9456 (N_9456,N_8846,N_8188);
xor U9457 (N_9457,N_8640,N_8657);
or U9458 (N_9458,N_8925,N_8883);
or U9459 (N_9459,N_8763,N_8323);
nand U9460 (N_9460,N_8031,N_8129);
nor U9461 (N_9461,N_8133,N_8539);
xor U9462 (N_9462,N_8470,N_8505);
xor U9463 (N_9463,N_8275,N_8776);
xor U9464 (N_9464,N_8234,N_8729);
and U9465 (N_9465,N_8350,N_8782);
nor U9466 (N_9466,N_8000,N_8882);
and U9467 (N_9467,N_8016,N_8407);
nand U9468 (N_9468,N_8554,N_8614);
and U9469 (N_9469,N_8680,N_8841);
nor U9470 (N_9470,N_8193,N_8183);
nand U9471 (N_9471,N_8511,N_8105);
and U9472 (N_9472,N_8831,N_8113);
or U9473 (N_9473,N_8840,N_8342);
xnor U9474 (N_9474,N_8477,N_8265);
xnor U9475 (N_9475,N_8324,N_8751);
nand U9476 (N_9476,N_8936,N_8889);
or U9477 (N_9477,N_8365,N_8488);
xor U9478 (N_9478,N_8681,N_8467);
nand U9479 (N_9479,N_8076,N_8635);
and U9480 (N_9480,N_8101,N_8843);
and U9481 (N_9481,N_8850,N_8856);
nor U9482 (N_9482,N_8369,N_8911);
and U9483 (N_9483,N_8373,N_8332);
nand U9484 (N_9484,N_8708,N_8224);
or U9485 (N_9485,N_8865,N_8953);
xnor U9486 (N_9486,N_8633,N_8487);
or U9487 (N_9487,N_8818,N_8828);
or U9488 (N_9488,N_8896,N_8779);
nand U9489 (N_9489,N_8506,N_8338);
nor U9490 (N_9490,N_8950,N_8650);
and U9491 (N_9491,N_8178,N_8881);
xnor U9492 (N_9492,N_8054,N_8191);
nor U9493 (N_9493,N_8363,N_8813);
or U9494 (N_9494,N_8995,N_8699);
xnor U9495 (N_9495,N_8780,N_8121);
or U9496 (N_9496,N_8395,N_8579);
or U9497 (N_9497,N_8240,N_8930);
xnor U9498 (N_9498,N_8926,N_8415);
or U9499 (N_9499,N_8367,N_8008);
nor U9500 (N_9500,N_8556,N_8695);
xnor U9501 (N_9501,N_8157,N_8972);
nand U9502 (N_9502,N_8663,N_8592);
nor U9503 (N_9503,N_8254,N_8205);
nor U9504 (N_9504,N_8998,N_8784);
xor U9505 (N_9505,N_8707,N_8239);
nand U9506 (N_9506,N_8999,N_8643);
nor U9507 (N_9507,N_8886,N_8019);
nor U9508 (N_9508,N_8642,N_8154);
and U9509 (N_9509,N_8962,N_8211);
and U9510 (N_9510,N_8263,N_8645);
or U9511 (N_9511,N_8401,N_8028);
and U9512 (N_9512,N_8901,N_8588);
xnor U9513 (N_9513,N_8556,N_8871);
xor U9514 (N_9514,N_8911,N_8916);
and U9515 (N_9515,N_8238,N_8533);
and U9516 (N_9516,N_8967,N_8443);
and U9517 (N_9517,N_8293,N_8107);
nand U9518 (N_9518,N_8875,N_8012);
xnor U9519 (N_9519,N_8446,N_8306);
and U9520 (N_9520,N_8787,N_8375);
nand U9521 (N_9521,N_8788,N_8252);
nand U9522 (N_9522,N_8405,N_8432);
nor U9523 (N_9523,N_8962,N_8124);
nand U9524 (N_9524,N_8652,N_8061);
nand U9525 (N_9525,N_8802,N_8268);
nor U9526 (N_9526,N_8772,N_8839);
nand U9527 (N_9527,N_8138,N_8027);
xnor U9528 (N_9528,N_8037,N_8993);
and U9529 (N_9529,N_8145,N_8014);
nand U9530 (N_9530,N_8702,N_8555);
xor U9531 (N_9531,N_8065,N_8216);
and U9532 (N_9532,N_8392,N_8824);
xor U9533 (N_9533,N_8339,N_8639);
or U9534 (N_9534,N_8468,N_8678);
nor U9535 (N_9535,N_8104,N_8010);
nand U9536 (N_9536,N_8599,N_8212);
nand U9537 (N_9537,N_8321,N_8474);
nor U9538 (N_9538,N_8330,N_8530);
nor U9539 (N_9539,N_8982,N_8729);
nand U9540 (N_9540,N_8934,N_8235);
xor U9541 (N_9541,N_8383,N_8384);
xnor U9542 (N_9542,N_8005,N_8271);
or U9543 (N_9543,N_8843,N_8249);
nor U9544 (N_9544,N_8708,N_8987);
and U9545 (N_9545,N_8672,N_8333);
nor U9546 (N_9546,N_8862,N_8263);
and U9547 (N_9547,N_8186,N_8116);
and U9548 (N_9548,N_8115,N_8776);
nor U9549 (N_9549,N_8519,N_8701);
nor U9550 (N_9550,N_8411,N_8804);
nand U9551 (N_9551,N_8116,N_8969);
nor U9552 (N_9552,N_8883,N_8723);
xor U9553 (N_9553,N_8184,N_8996);
and U9554 (N_9554,N_8384,N_8272);
or U9555 (N_9555,N_8561,N_8661);
nand U9556 (N_9556,N_8713,N_8842);
nor U9557 (N_9557,N_8096,N_8247);
or U9558 (N_9558,N_8263,N_8825);
nand U9559 (N_9559,N_8554,N_8574);
nor U9560 (N_9560,N_8369,N_8922);
xor U9561 (N_9561,N_8057,N_8187);
nand U9562 (N_9562,N_8371,N_8876);
and U9563 (N_9563,N_8485,N_8271);
xnor U9564 (N_9564,N_8654,N_8310);
nor U9565 (N_9565,N_8443,N_8871);
or U9566 (N_9566,N_8410,N_8156);
or U9567 (N_9567,N_8713,N_8674);
nand U9568 (N_9568,N_8639,N_8651);
xnor U9569 (N_9569,N_8194,N_8276);
or U9570 (N_9570,N_8682,N_8582);
nand U9571 (N_9571,N_8241,N_8841);
nor U9572 (N_9572,N_8767,N_8391);
xor U9573 (N_9573,N_8168,N_8471);
or U9574 (N_9574,N_8135,N_8510);
and U9575 (N_9575,N_8133,N_8792);
nand U9576 (N_9576,N_8525,N_8437);
nor U9577 (N_9577,N_8946,N_8601);
and U9578 (N_9578,N_8886,N_8942);
nor U9579 (N_9579,N_8551,N_8888);
or U9580 (N_9580,N_8528,N_8158);
xnor U9581 (N_9581,N_8358,N_8956);
or U9582 (N_9582,N_8578,N_8261);
nor U9583 (N_9583,N_8923,N_8428);
nand U9584 (N_9584,N_8475,N_8552);
nand U9585 (N_9585,N_8641,N_8203);
and U9586 (N_9586,N_8947,N_8527);
nand U9587 (N_9587,N_8438,N_8202);
nor U9588 (N_9588,N_8830,N_8254);
nand U9589 (N_9589,N_8353,N_8441);
nor U9590 (N_9590,N_8078,N_8565);
and U9591 (N_9591,N_8548,N_8773);
xor U9592 (N_9592,N_8100,N_8516);
xor U9593 (N_9593,N_8890,N_8610);
xor U9594 (N_9594,N_8728,N_8939);
or U9595 (N_9595,N_8955,N_8306);
nand U9596 (N_9596,N_8495,N_8171);
xor U9597 (N_9597,N_8593,N_8015);
or U9598 (N_9598,N_8244,N_8783);
and U9599 (N_9599,N_8856,N_8263);
and U9600 (N_9600,N_8434,N_8225);
nor U9601 (N_9601,N_8053,N_8468);
or U9602 (N_9602,N_8069,N_8613);
and U9603 (N_9603,N_8862,N_8032);
and U9604 (N_9604,N_8911,N_8174);
or U9605 (N_9605,N_8024,N_8386);
nand U9606 (N_9606,N_8997,N_8890);
nor U9607 (N_9607,N_8898,N_8852);
and U9608 (N_9608,N_8202,N_8322);
xor U9609 (N_9609,N_8772,N_8237);
nor U9610 (N_9610,N_8220,N_8645);
or U9611 (N_9611,N_8065,N_8274);
nor U9612 (N_9612,N_8336,N_8388);
nor U9613 (N_9613,N_8566,N_8661);
nand U9614 (N_9614,N_8805,N_8964);
xnor U9615 (N_9615,N_8259,N_8415);
xor U9616 (N_9616,N_8068,N_8776);
or U9617 (N_9617,N_8112,N_8762);
nor U9618 (N_9618,N_8365,N_8678);
xnor U9619 (N_9619,N_8962,N_8786);
or U9620 (N_9620,N_8197,N_8810);
nor U9621 (N_9621,N_8552,N_8748);
nor U9622 (N_9622,N_8023,N_8348);
nand U9623 (N_9623,N_8800,N_8769);
and U9624 (N_9624,N_8591,N_8608);
or U9625 (N_9625,N_8221,N_8421);
and U9626 (N_9626,N_8668,N_8785);
nor U9627 (N_9627,N_8371,N_8121);
nor U9628 (N_9628,N_8528,N_8733);
and U9629 (N_9629,N_8873,N_8198);
xor U9630 (N_9630,N_8792,N_8079);
and U9631 (N_9631,N_8078,N_8531);
or U9632 (N_9632,N_8244,N_8363);
xor U9633 (N_9633,N_8510,N_8145);
and U9634 (N_9634,N_8674,N_8976);
nand U9635 (N_9635,N_8278,N_8957);
nand U9636 (N_9636,N_8253,N_8568);
nor U9637 (N_9637,N_8781,N_8791);
nor U9638 (N_9638,N_8036,N_8140);
nand U9639 (N_9639,N_8913,N_8053);
nand U9640 (N_9640,N_8884,N_8293);
nand U9641 (N_9641,N_8732,N_8788);
nand U9642 (N_9642,N_8780,N_8697);
xor U9643 (N_9643,N_8588,N_8103);
xnor U9644 (N_9644,N_8464,N_8365);
or U9645 (N_9645,N_8211,N_8849);
nor U9646 (N_9646,N_8541,N_8512);
or U9647 (N_9647,N_8833,N_8335);
nand U9648 (N_9648,N_8519,N_8779);
and U9649 (N_9649,N_8717,N_8468);
xor U9650 (N_9650,N_8297,N_8617);
and U9651 (N_9651,N_8438,N_8644);
nor U9652 (N_9652,N_8828,N_8366);
nor U9653 (N_9653,N_8843,N_8788);
nand U9654 (N_9654,N_8497,N_8437);
or U9655 (N_9655,N_8118,N_8755);
nand U9656 (N_9656,N_8387,N_8164);
or U9657 (N_9657,N_8675,N_8124);
and U9658 (N_9658,N_8280,N_8723);
xor U9659 (N_9659,N_8156,N_8531);
xor U9660 (N_9660,N_8186,N_8004);
xnor U9661 (N_9661,N_8663,N_8666);
nand U9662 (N_9662,N_8043,N_8108);
nor U9663 (N_9663,N_8285,N_8160);
xor U9664 (N_9664,N_8441,N_8121);
and U9665 (N_9665,N_8965,N_8019);
nor U9666 (N_9666,N_8548,N_8704);
xor U9667 (N_9667,N_8266,N_8981);
xor U9668 (N_9668,N_8372,N_8416);
nand U9669 (N_9669,N_8546,N_8370);
or U9670 (N_9670,N_8714,N_8246);
xnor U9671 (N_9671,N_8778,N_8641);
and U9672 (N_9672,N_8900,N_8040);
nor U9673 (N_9673,N_8892,N_8399);
or U9674 (N_9674,N_8990,N_8653);
nand U9675 (N_9675,N_8324,N_8986);
and U9676 (N_9676,N_8418,N_8638);
or U9677 (N_9677,N_8112,N_8149);
xor U9678 (N_9678,N_8880,N_8257);
xnor U9679 (N_9679,N_8567,N_8911);
nand U9680 (N_9680,N_8969,N_8469);
nand U9681 (N_9681,N_8896,N_8233);
nor U9682 (N_9682,N_8741,N_8841);
nand U9683 (N_9683,N_8928,N_8415);
or U9684 (N_9684,N_8136,N_8041);
and U9685 (N_9685,N_8749,N_8981);
and U9686 (N_9686,N_8373,N_8211);
nor U9687 (N_9687,N_8422,N_8647);
xnor U9688 (N_9688,N_8286,N_8736);
and U9689 (N_9689,N_8659,N_8121);
nand U9690 (N_9690,N_8873,N_8863);
or U9691 (N_9691,N_8915,N_8963);
nand U9692 (N_9692,N_8369,N_8846);
or U9693 (N_9693,N_8470,N_8382);
nand U9694 (N_9694,N_8633,N_8238);
xnor U9695 (N_9695,N_8236,N_8856);
xor U9696 (N_9696,N_8611,N_8905);
or U9697 (N_9697,N_8108,N_8009);
nand U9698 (N_9698,N_8117,N_8458);
nor U9699 (N_9699,N_8341,N_8892);
nand U9700 (N_9700,N_8683,N_8688);
and U9701 (N_9701,N_8003,N_8461);
or U9702 (N_9702,N_8397,N_8619);
nand U9703 (N_9703,N_8275,N_8685);
xnor U9704 (N_9704,N_8615,N_8082);
or U9705 (N_9705,N_8571,N_8613);
and U9706 (N_9706,N_8567,N_8021);
or U9707 (N_9707,N_8932,N_8746);
xor U9708 (N_9708,N_8516,N_8271);
and U9709 (N_9709,N_8321,N_8195);
nand U9710 (N_9710,N_8924,N_8312);
nand U9711 (N_9711,N_8335,N_8371);
or U9712 (N_9712,N_8972,N_8469);
xor U9713 (N_9713,N_8087,N_8388);
xor U9714 (N_9714,N_8609,N_8874);
and U9715 (N_9715,N_8992,N_8322);
and U9716 (N_9716,N_8595,N_8039);
nand U9717 (N_9717,N_8798,N_8434);
xnor U9718 (N_9718,N_8555,N_8109);
or U9719 (N_9719,N_8422,N_8355);
and U9720 (N_9720,N_8715,N_8055);
xor U9721 (N_9721,N_8834,N_8012);
or U9722 (N_9722,N_8804,N_8270);
nor U9723 (N_9723,N_8072,N_8531);
nand U9724 (N_9724,N_8033,N_8796);
and U9725 (N_9725,N_8533,N_8865);
nand U9726 (N_9726,N_8574,N_8886);
xor U9727 (N_9727,N_8744,N_8045);
nor U9728 (N_9728,N_8785,N_8861);
xnor U9729 (N_9729,N_8773,N_8462);
or U9730 (N_9730,N_8574,N_8060);
or U9731 (N_9731,N_8096,N_8419);
xor U9732 (N_9732,N_8224,N_8817);
and U9733 (N_9733,N_8527,N_8575);
nor U9734 (N_9734,N_8875,N_8533);
nor U9735 (N_9735,N_8159,N_8521);
xnor U9736 (N_9736,N_8964,N_8051);
xnor U9737 (N_9737,N_8666,N_8977);
nor U9738 (N_9738,N_8822,N_8857);
nor U9739 (N_9739,N_8917,N_8550);
and U9740 (N_9740,N_8782,N_8813);
nor U9741 (N_9741,N_8939,N_8589);
nor U9742 (N_9742,N_8211,N_8311);
xor U9743 (N_9743,N_8691,N_8381);
nor U9744 (N_9744,N_8350,N_8806);
and U9745 (N_9745,N_8035,N_8879);
and U9746 (N_9746,N_8684,N_8157);
nor U9747 (N_9747,N_8169,N_8604);
nand U9748 (N_9748,N_8778,N_8402);
nand U9749 (N_9749,N_8885,N_8403);
xnor U9750 (N_9750,N_8034,N_8272);
or U9751 (N_9751,N_8443,N_8055);
xor U9752 (N_9752,N_8974,N_8142);
nand U9753 (N_9753,N_8113,N_8036);
and U9754 (N_9754,N_8377,N_8461);
nand U9755 (N_9755,N_8966,N_8035);
xnor U9756 (N_9756,N_8476,N_8981);
nor U9757 (N_9757,N_8383,N_8873);
or U9758 (N_9758,N_8375,N_8965);
nand U9759 (N_9759,N_8060,N_8627);
and U9760 (N_9760,N_8626,N_8677);
nor U9761 (N_9761,N_8572,N_8197);
and U9762 (N_9762,N_8616,N_8671);
or U9763 (N_9763,N_8462,N_8089);
xor U9764 (N_9764,N_8983,N_8275);
nor U9765 (N_9765,N_8056,N_8264);
or U9766 (N_9766,N_8949,N_8408);
xor U9767 (N_9767,N_8505,N_8358);
nand U9768 (N_9768,N_8874,N_8930);
or U9769 (N_9769,N_8145,N_8736);
or U9770 (N_9770,N_8144,N_8783);
nand U9771 (N_9771,N_8922,N_8955);
xnor U9772 (N_9772,N_8705,N_8838);
or U9773 (N_9773,N_8597,N_8920);
nand U9774 (N_9774,N_8047,N_8927);
nand U9775 (N_9775,N_8857,N_8350);
or U9776 (N_9776,N_8201,N_8584);
or U9777 (N_9777,N_8442,N_8465);
nor U9778 (N_9778,N_8209,N_8808);
nand U9779 (N_9779,N_8387,N_8724);
or U9780 (N_9780,N_8229,N_8407);
or U9781 (N_9781,N_8997,N_8081);
nor U9782 (N_9782,N_8865,N_8315);
xor U9783 (N_9783,N_8037,N_8345);
or U9784 (N_9784,N_8909,N_8274);
xnor U9785 (N_9785,N_8848,N_8288);
nor U9786 (N_9786,N_8893,N_8644);
or U9787 (N_9787,N_8596,N_8925);
and U9788 (N_9788,N_8979,N_8387);
nand U9789 (N_9789,N_8503,N_8131);
and U9790 (N_9790,N_8281,N_8776);
xnor U9791 (N_9791,N_8839,N_8500);
nand U9792 (N_9792,N_8130,N_8053);
nor U9793 (N_9793,N_8431,N_8600);
nand U9794 (N_9794,N_8622,N_8101);
or U9795 (N_9795,N_8928,N_8745);
xnor U9796 (N_9796,N_8348,N_8193);
xor U9797 (N_9797,N_8515,N_8282);
nand U9798 (N_9798,N_8066,N_8332);
and U9799 (N_9799,N_8129,N_8188);
nor U9800 (N_9800,N_8109,N_8343);
or U9801 (N_9801,N_8006,N_8480);
xnor U9802 (N_9802,N_8803,N_8414);
and U9803 (N_9803,N_8600,N_8280);
or U9804 (N_9804,N_8109,N_8564);
nor U9805 (N_9805,N_8870,N_8434);
xor U9806 (N_9806,N_8556,N_8171);
xnor U9807 (N_9807,N_8591,N_8681);
and U9808 (N_9808,N_8818,N_8665);
and U9809 (N_9809,N_8008,N_8003);
nand U9810 (N_9810,N_8996,N_8646);
and U9811 (N_9811,N_8563,N_8876);
or U9812 (N_9812,N_8843,N_8183);
nand U9813 (N_9813,N_8160,N_8451);
and U9814 (N_9814,N_8966,N_8159);
nor U9815 (N_9815,N_8617,N_8386);
nor U9816 (N_9816,N_8916,N_8500);
nor U9817 (N_9817,N_8865,N_8329);
xor U9818 (N_9818,N_8209,N_8745);
xnor U9819 (N_9819,N_8828,N_8934);
xor U9820 (N_9820,N_8374,N_8404);
or U9821 (N_9821,N_8816,N_8770);
and U9822 (N_9822,N_8327,N_8747);
nand U9823 (N_9823,N_8551,N_8384);
nor U9824 (N_9824,N_8290,N_8589);
nor U9825 (N_9825,N_8760,N_8567);
and U9826 (N_9826,N_8855,N_8073);
and U9827 (N_9827,N_8162,N_8577);
xor U9828 (N_9828,N_8732,N_8066);
nand U9829 (N_9829,N_8715,N_8437);
and U9830 (N_9830,N_8849,N_8606);
or U9831 (N_9831,N_8667,N_8316);
xor U9832 (N_9832,N_8385,N_8397);
nand U9833 (N_9833,N_8029,N_8001);
nand U9834 (N_9834,N_8963,N_8551);
or U9835 (N_9835,N_8503,N_8940);
nor U9836 (N_9836,N_8186,N_8299);
nand U9837 (N_9837,N_8735,N_8425);
nand U9838 (N_9838,N_8363,N_8400);
nand U9839 (N_9839,N_8062,N_8800);
nand U9840 (N_9840,N_8849,N_8825);
nor U9841 (N_9841,N_8374,N_8264);
nand U9842 (N_9842,N_8721,N_8709);
or U9843 (N_9843,N_8178,N_8535);
or U9844 (N_9844,N_8300,N_8970);
or U9845 (N_9845,N_8011,N_8765);
nand U9846 (N_9846,N_8056,N_8702);
or U9847 (N_9847,N_8815,N_8607);
or U9848 (N_9848,N_8713,N_8575);
xor U9849 (N_9849,N_8606,N_8198);
nand U9850 (N_9850,N_8201,N_8447);
xnor U9851 (N_9851,N_8779,N_8495);
or U9852 (N_9852,N_8889,N_8691);
nor U9853 (N_9853,N_8251,N_8892);
and U9854 (N_9854,N_8493,N_8233);
nor U9855 (N_9855,N_8843,N_8140);
and U9856 (N_9856,N_8459,N_8308);
and U9857 (N_9857,N_8204,N_8583);
or U9858 (N_9858,N_8508,N_8012);
nor U9859 (N_9859,N_8252,N_8699);
nand U9860 (N_9860,N_8034,N_8343);
xnor U9861 (N_9861,N_8303,N_8931);
or U9862 (N_9862,N_8403,N_8143);
xor U9863 (N_9863,N_8388,N_8813);
and U9864 (N_9864,N_8318,N_8296);
nor U9865 (N_9865,N_8244,N_8419);
nand U9866 (N_9866,N_8240,N_8029);
xor U9867 (N_9867,N_8306,N_8533);
nand U9868 (N_9868,N_8921,N_8845);
nor U9869 (N_9869,N_8316,N_8514);
and U9870 (N_9870,N_8489,N_8518);
or U9871 (N_9871,N_8601,N_8966);
nand U9872 (N_9872,N_8065,N_8113);
and U9873 (N_9873,N_8687,N_8778);
nand U9874 (N_9874,N_8313,N_8104);
nand U9875 (N_9875,N_8040,N_8713);
or U9876 (N_9876,N_8367,N_8723);
and U9877 (N_9877,N_8822,N_8425);
or U9878 (N_9878,N_8914,N_8699);
nor U9879 (N_9879,N_8589,N_8542);
nor U9880 (N_9880,N_8301,N_8971);
xnor U9881 (N_9881,N_8075,N_8412);
and U9882 (N_9882,N_8714,N_8996);
nand U9883 (N_9883,N_8907,N_8280);
xnor U9884 (N_9884,N_8638,N_8897);
or U9885 (N_9885,N_8169,N_8683);
nor U9886 (N_9886,N_8793,N_8351);
nand U9887 (N_9887,N_8322,N_8043);
xor U9888 (N_9888,N_8257,N_8137);
xor U9889 (N_9889,N_8419,N_8781);
or U9890 (N_9890,N_8421,N_8272);
or U9891 (N_9891,N_8589,N_8239);
nand U9892 (N_9892,N_8783,N_8836);
or U9893 (N_9893,N_8979,N_8441);
nand U9894 (N_9894,N_8139,N_8448);
nor U9895 (N_9895,N_8912,N_8472);
or U9896 (N_9896,N_8886,N_8868);
or U9897 (N_9897,N_8161,N_8534);
xor U9898 (N_9898,N_8359,N_8412);
and U9899 (N_9899,N_8649,N_8700);
nor U9900 (N_9900,N_8840,N_8274);
or U9901 (N_9901,N_8496,N_8696);
nor U9902 (N_9902,N_8767,N_8984);
xnor U9903 (N_9903,N_8426,N_8594);
and U9904 (N_9904,N_8966,N_8407);
or U9905 (N_9905,N_8970,N_8064);
and U9906 (N_9906,N_8487,N_8994);
nor U9907 (N_9907,N_8583,N_8019);
and U9908 (N_9908,N_8137,N_8743);
xnor U9909 (N_9909,N_8686,N_8882);
xor U9910 (N_9910,N_8951,N_8181);
nor U9911 (N_9911,N_8242,N_8733);
xnor U9912 (N_9912,N_8220,N_8573);
or U9913 (N_9913,N_8649,N_8851);
nand U9914 (N_9914,N_8057,N_8539);
nor U9915 (N_9915,N_8552,N_8152);
and U9916 (N_9916,N_8463,N_8605);
or U9917 (N_9917,N_8831,N_8324);
xnor U9918 (N_9918,N_8390,N_8019);
or U9919 (N_9919,N_8168,N_8426);
or U9920 (N_9920,N_8611,N_8578);
xnor U9921 (N_9921,N_8831,N_8001);
and U9922 (N_9922,N_8992,N_8799);
nor U9923 (N_9923,N_8571,N_8631);
or U9924 (N_9924,N_8252,N_8394);
xor U9925 (N_9925,N_8822,N_8995);
nand U9926 (N_9926,N_8734,N_8607);
xor U9927 (N_9927,N_8243,N_8913);
and U9928 (N_9928,N_8620,N_8426);
xor U9929 (N_9929,N_8674,N_8186);
nand U9930 (N_9930,N_8887,N_8153);
nand U9931 (N_9931,N_8596,N_8440);
and U9932 (N_9932,N_8129,N_8041);
and U9933 (N_9933,N_8783,N_8389);
nand U9934 (N_9934,N_8661,N_8559);
nor U9935 (N_9935,N_8734,N_8083);
nand U9936 (N_9936,N_8897,N_8634);
or U9937 (N_9937,N_8199,N_8578);
nor U9938 (N_9938,N_8453,N_8174);
nand U9939 (N_9939,N_8278,N_8981);
or U9940 (N_9940,N_8421,N_8597);
or U9941 (N_9941,N_8509,N_8102);
or U9942 (N_9942,N_8820,N_8150);
or U9943 (N_9943,N_8639,N_8904);
or U9944 (N_9944,N_8748,N_8379);
nand U9945 (N_9945,N_8774,N_8609);
nand U9946 (N_9946,N_8004,N_8312);
nand U9947 (N_9947,N_8141,N_8650);
nor U9948 (N_9948,N_8095,N_8119);
or U9949 (N_9949,N_8757,N_8354);
and U9950 (N_9950,N_8519,N_8974);
nand U9951 (N_9951,N_8494,N_8287);
xnor U9952 (N_9952,N_8349,N_8205);
nor U9953 (N_9953,N_8912,N_8902);
or U9954 (N_9954,N_8983,N_8850);
and U9955 (N_9955,N_8079,N_8673);
xnor U9956 (N_9956,N_8603,N_8304);
nand U9957 (N_9957,N_8681,N_8555);
xor U9958 (N_9958,N_8319,N_8004);
xnor U9959 (N_9959,N_8442,N_8344);
or U9960 (N_9960,N_8347,N_8433);
or U9961 (N_9961,N_8129,N_8568);
or U9962 (N_9962,N_8838,N_8440);
or U9963 (N_9963,N_8050,N_8053);
or U9964 (N_9964,N_8979,N_8783);
nand U9965 (N_9965,N_8117,N_8057);
or U9966 (N_9966,N_8381,N_8920);
xor U9967 (N_9967,N_8133,N_8114);
nor U9968 (N_9968,N_8664,N_8263);
and U9969 (N_9969,N_8030,N_8789);
xnor U9970 (N_9970,N_8755,N_8190);
nor U9971 (N_9971,N_8955,N_8001);
nand U9972 (N_9972,N_8490,N_8916);
or U9973 (N_9973,N_8859,N_8054);
and U9974 (N_9974,N_8851,N_8156);
nor U9975 (N_9975,N_8494,N_8082);
and U9976 (N_9976,N_8337,N_8944);
nand U9977 (N_9977,N_8150,N_8315);
xnor U9978 (N_9978,N_8456,N_8885);
and U9979 (N_9979,N_8868,N_8676);
nor U9980 (N_9980,N_8548,N_8577);
and U9981 (N_9981,N_8272,N_8371);
and U9982 (N_9982,N_8143,N_8123);
or U9983 (N_9983,N_8930,N_8808);
and U9984 (N_9984,N_8776,N_8416);
xor U9985 (N_9985,N_8789,N_8738);
nor U9986 (N_9986,N_8921,N_8898);
nand U9987 (N_9987,N_8301,N_8484);
or U9988 (N_9988,N_8763,N_8125);
and U9989 (N_9989,N_8924,N_8966);
xor U9990 (N_9990,N_8854,N_8210);
nand U9991 (N_9991,N_8801,N_8568);
and U9992 (N_9992,N_8550,N_8210);
nor U9993 (N_9993,N_8708,N_8246);
xor U9994 (N_9994,N_8237,N_8490);
and U9995 (N_9995,N_8520,N_8172);
and U9996 (N_9996,N_8171,N_8304);
nand U9997 (N_9997,N_8557,N_8669);
nor U9998 (N_9998,N_8323,N_8210);
nor U9999 (N_9999,N_8996,N_8143);
nor U10000 (N_10000,N_9826,N_9607);
and U10001 (N_10001,N_9158,N_9401);
and U10002 (N_10002,N_9244,N_9575);
or U10003 (N_10003,N_9009,N_9679);
xor U10004 (N_10004,N_9530,N_9506);
or U10005 (N_10005,N_9662,N_9921);
and U10006 (N_10006,N_9043,N_9296);
or U10007 (N_10007,N_9061,N_9204);
and U10008 (N_10008,N_9238,N_9508);
nand U10009 (N_10009,N_9068,N_9150);
nand U10010 (N_10010,N_9383,N_9710);
nor U10011 (N_10011,N_9487,N_9300);
xnor U10012 (N_10012,N_9420,N_9926);
and U10013 (N_10013,N_9769,N_9876);
or U10014 (N_10014,N_9527,N_9391);
nand U10015 (N_10015,N_9587,N_9106);
nor U10016 (N_10016,N_9291,N_9614);
nand U10017 (N_10017,N_9877,N_9036);
nand U10018 (N_10018,N_9138,N_9865);
or U10019 (N_10019,N_9202,N_9483);
or U10020 (N_10020,N_9501,N_9638);
and U10021 (N_10021,N_9741,N_9059);
and U10022 (N_10022,N_9367,N_9313);
and U10023 (N_10023,N_9133,N_9813);
and U10024 (N_10024,N_9262,N_9547);
xor U10025 (N_10025,N_9311,N_9035);
xnor U10026 (N_10026,N_9408,N_9688);
xor U10027 (N_10027,N_9753,N_9943);
or U10028 (N_10028,N_9867,N_9681);
xor U10029 (N_10029,N_9003,N_9720);
nand U10030 (N_10030,N_9208,N_9087);
nor U10031 (N_10031,N_9413,N_9891);
xnor U10032 (N_10032,N_9493,N_9498);
nor U10033 (N_10033,N_9694,N_9132);
nand U10034 (N_10034,N_9522,N_9334);
or U10035 (N_10035,N_9496,N_9653);
and U10036 (N_10036,N_9934,N_9800);
or U10037 (N_10037,N_9794,N_9310);
and U10038 (N_10038,N_9905,N_9161);
nand U10039 (N_10039,N_9916,N_9576);
xnor U10040 (N_10040,N_9193,N_9386);
or U10041 (N_10041,N_9349,N_9376);
or U10042 (N_10042,N_9528,N_9181);
nand U10043 (N_10043,N_9615,N_9260);
nor U10044 (N_10044,N_9987,N_9006);
xor U10045 (N_10045,N_9786,N_9140);
nor U10046 (N_10046,N_9257,N_9904);
xnor U10047 (N_10047,N_9821,N_9321);
and U10048 (N_10048,N_9422,N_9971);
nand U10049 (N_10049,N_9596,N_9569);
nor U10050 (N_10050,N_9728,N_9689);
and U10051 (N_10051,N_9466,N_9154);
nand U10052 (N_10052,N_9079,N_9130);
nand U10053 (N_10053,N_9517,N_9234);
or U10054 (N_10054,N_9960,N_9935);
nand U10055 (N_10055,N_9211,N_9892);
and U10056 (N_10056,N_9481,N_9388);
nand U10057 (N_10057,N_9286,N_9840);
nand U10058 (N_10058,N_9024,N_9718);
and U10059 (N_10059,N_9463,N_9669);
xor U10060 (N_10060,N_9210,N_9472);
and U10061 (N_10061,N_9439,N_9478);
xor U10062 (N_10062,N_9649,N_9324);
nand U10063 (N_10063,N_9788,N_9924);
nor U10064 (N_10064,N_9185,N_9082);
and U10065 (N_10065,N_9727,N_9419);
xnor U10066 (N_10066,N_9127,N_9872);
or U10067 (N_10067,N_9529,N_9806);
or U10068 (N_10068,N_9621,N_9965);
or U10069 (N_10069,N_9426,N_9574);
or U10070 (N_10070,N_9243,N_9881);
or U10071 (N_10071,N_9812,N_9016);
nor U10072 (N_10072,N_9803,N_9091);
nand U10073 (N_10073,N_9565,N_9578);
nor U10074 (N_10074,N_9562,N_9038);
xor U10075 (N_10075,N_9863,N_9785);
nor U10076 (N_10076,N_9392,N_9414);
and U10077 (N_10077,N_9768,N_9586);
xor U10078 (N_10078,N_9982,N_9437);
and U10079 (N_10079,N_9882,N_9817);
or U10080 (N_10080,N_9983,N_9331);
xor U10081 (N_10081,N_9326,N_9719);
xor U10082 (N_10082,N_9250,N_9609);
and U10083 (N_10083,N_9017,N_9278);
or U10084 (N_10084,N_9111,N_9510);
or U10085 (N_10085,N_9630,N_9455);
nand U10086 (N_10086,N_9054,N_9946);
and U10087 (N_10087,N_9680,N_9378);
and U10088 (N_10088,N_9101,N_9595);
nand U10089 (N_10089,N_9169,N_9667);
nand U10090 (N_10090,N_9665,N_9717);
and U10091 (N_10091,N_9359,N_9362);
nor U10092 (N_10092,N_9115,N_9103);
and U10093 (N_10093,N_9668,N_9382);
nand U10094 (N_10094,N_9824,N_9002);
xor U10095 (N_10095,N_9648,N_9950);
or U10096 (N_10096,N_9105,N_9637);
nor U10097 (N_10097,N_9956,N_9818);
xor U10098 (N_10098,N_9886,N_9352);
xnor U10099 (N_10099,N_9789,N_9754);
nand U10100 (N_10100,N_9799,N_9771);
and U10101 (N_10101,N_9592,N_9116);
and U10102 (N_10102,N_9053,N_9209);
or U10103 (N_10103,N_9471,N_9235);
and U10104 (N_10104,N_9676,N_9585);
xor U10105 (N_10105,N_9333,N_9879);
xnor U10106 (N_10106,N_9692,N_9602);
nand U10107 (N_10107,N_9525,N_9029);
xor U10108 (N_10108,N_9344,N_9294);
nand U10109 (N_10109,N_9486,N_9268);
nand U10110 (N_10110,N_9857,N_9889);
and U10111 (N_10111,N_9675,N_9329);
or U10112 (N_10112,N_9948,N_9086);
and U10113 (N_10113,N_9521,N_9046);
nand U10114 (N_10114,N_9171,N_9492);
xnor U10115 (N_10115,N_9514,N_9224);
nor U10116 (N_10116,N_9792,N_9148);
nand U10117 (N_10117,N_9758,N_9027);
nand U10118 (N_10118,N_9804,N_9540);
nor U10119 (N_10119,N_9639,N_9139);
and U10120 (N_10120,N_9128,N_9125);
and U10121 (N_10121,N_9845,N_9536);
nand U10122 (N_10122,N_9307,N_9220);
or U10123 (N_10123,N_9656,N_9096);
xnor U10124 (N_10124,N_9743,N_9914);
nor U10125 (N_10125,N_9584,N_9494);
nand U10126 (N_10126,N_9146,N_9573);
nor U10127 (N_10127,N_9511,N_9825);
and U10128 (N_10128,N_9020,N_9760);
and U10129 (N_10129,N_9631,N_9069);
or U10130 (N_10130,N_9572,N_9791);
xor U10131 (N_10131,N_9843,N_9099);
nor U10132 (N_10132,N_9242,N_9301);
or U10133 (N_10133,N_9773,N_9348);
and U10134 (N_10134,N_9178,N_9438);
or U10135 (N_10135,N_9165,N_9962);
and U10136 (N_10136,N_9449,N_9998);
xor U10137 (N_10137,N_9339,N_9822);
xnor U10138 (N_10138,N_9714,N_9842);
or U10139 (N_10139,N_9942,N_9315);
xnor U10140 (N_10140,N_9075,N_9205);
nand U10141 (N_10141,N_9733,N_9920);
nor U10142 (N_10142,N_9289,N_9980);
nor U10143 (N_10143,N_9734,N_9861);
nor U10144 (N_10144,N_9070,N_9040);
nand U10145 (N_10145,N_9659,N_9698);
nand U10146 (N_10146,N_9505,N_9940);
and U10147 (N_10147,N_9526,N_9440);
or U10148 (N_10148,N_9259,N_9599);
or U10149 (N_10149,N_9938,N_9080);
xor U10150 (N_10150,N_9322,N_9306);
nor U10151 (N_10151,N_9447,N_9513);
nor U10152 (N_10152,N_9197,N_9135);
nor U10153 (N_10153,N_9869,N_9913);
nor U10154 (N_10154,N_9093,N_9851);
nand U10155 (N_10155,N_9502,N_9958);
nand U10156 (N_10156,N_9194,N_9251);
and U10157 (N_10157,N_9738,N_9853);
or U10158 (N_10158,N_9121,N_9593);
xnor U10159 (N_10159,N_9247,N_9222);
nor U10160 (N_10160,N_9370,N_9763);
nor U10161 (N_10161,N_9484,N_9335);
or U10162 (N_10162,N_9088,N_9073);
and U10163 (N_10163,N_9775,N_9037);
or U10164 (N_10164,N_9828,N_9542);
xnor U10165 (N_10165,N_9774,N_9605);
xor U10166 (N_10166,N_9767,N_9873);
nor U10167 (N_10167,N_9240,N_9462);
nor U10168 (N_10168,N_9395,N_9500);
nand U10169 (N_10169,N_9149,N_9212);
nor U10170 (N_10170,N_9100,N_9163);
nor U10171 (N_10171,N_9868,N_9044);
nor U10172 (N_10172,N_9827,N_9600);
nand U10173 (N_10173,N_9880,N_9625);
and U10174 (N_10174,N_9480,N_9063);
or U10175 (N_10175,N_9730,N_9279);
xnor U10176 (N_10176,N_9001,N_9495);
nand U10177 (N_10177,N_9545,N_9424);
nand U10178 (N_10178,N_9673,N_9102);
nor U10179 (N_10179,N_9287,N_9923);
xnor U10180 (N_10180,N_9459,N_9475);
nor U10181 (N_10181,N_9107,N_9622);
or U10182 (N_10182,N_9026,N_9328);
and U10183 (N_10183,N_9752,N_9110);
and U10184 (N_10184,N_9490,N_9559);
and U10185 (N_10185,N_9065,N_9470);
or U10186 (N_10186,N_9353,N_9729);
nor U10187 (N_10187,N_9742,N_9355);
and U10188 (N_10188,N_9795,N_9532);
nand U10189 (N_10189,N_9085,N_9317);
xnor U10190 (N_10190,N_9270,N_9885);
or U10191 (N_10191,N_9167,N_9953);
nand U10192 (N_10192,N_9837,N_9174);
and U10193 (N_10193,N_9901,N_9398);
and U10194 (N_10194,N_9314,N_9014);
nor U10195 (N_10195,N_9340,N_9011);
nand U10196 (N_10196,N_9485,N_9531);
xor U10197 (N_10197,N_9083,N_9271);
or U10198 (N_10198,N_9354,N_9590);
or U10199 (N_10199,N_9189,N_9008);
xor U10200 (N_10200,N_9482,N_9779);
xnor U10201 (N_10201,N_9970,N_9476);
or U10202 (N_10202,N_9062,N_9261);
and U10203 (N_10203,N_9968,N_9830);
xnor U10204 (N_10204,N_9316,N_9410);
and U10205 (N_10205,N_9090,N_9556);
and U10206 (N_10206,N_9553,N_9337);
nand U10207 (N_10207,N_9223,N_9706);
nand U10208 (N_10208,N_9267,N_9726);
xnor U10209 (N_10209,N_9831,N_9524);
or U10210 (N_10210,N_9922,N_9216);
and U10211 (N_10211,N_9276,N_9474);
or U10212 (N_10212,N_9191,N_9379);
nor U10213 (N_10213,N_9429,N_9421);
and U10214 (N_10214,N_9497,N_9409);
or U10215 (N_10215,N_9433,N_9134);
and U10216 (N_10216,N_9263,N_9911);
xnor U10217 (N_10217,N_9693,N_9985);
xor U10218 (N_10218,N_9722,N_9887);
or U10219 (N_10219,N_9218,N_9076);
and U10220 (N_10220,N_9539,N_9520);
nand U10221 (N_10221,N_9180,N_9533);
nor U10222 (N_10222,N_9973,N_9254);
nor U10223 (N_10223,N_9118,N_9384);
and U10224 (N_10224,N_9012,N_9320);
xnor U10225 (N_10225,N_9336,N_9452);
nand U10226 (N_10226,N_9032,N_9173);
or U10227 (N_10227,N_9974,N_9347);
xor U10228 (N_10228,N_9708,N_9890);
nand U10229 (N_10229,N_9430,N_9229);
xor U10230 (N_10230,N_9835,N_9757);
or U10231 (N_10231,N_9509,N_9207);
or U10232 (N_10232,N_9780,N_9518);
xor U10233 (N_10233,N_9350,N_9156);
xor U10234 (N_10234,N_9512,N_9147);
and U10235 (N_10235,N_9385,N_9947);
nor U10236 (N_10236,N_9666,N_9214);
and U10237 (N_10237,N_9927,N_9168);
nand U10238 (N_10238,N_9071,N_9796);
or U10239 (N_10239,N_9141,N_9390);
nand U10240 (N_10240,N_9227,N_9696);
xor U10241 (N_10241,N_9523,N_9707);
and U10242 (N_10242,N_9626,N_9435);
nor U10243 (N_10243,N_9119,N_9641);
and U10244 (N_10244,N_9781,N_9416);
xor U10245 (N_10245,N_9755,N_9374);
and U10246 (N_10246,N_9451,N_9023);
nor U10247 (N_10247,N_9672,N_9381);
xnor U10248 (N_10248,N_9721,N_9588);
xnor U10249 (N_10249,N_9396,N_9635);
nand U10250 (N_10250,N_9613,N_9897);
xnor U10251 (N_10251,N_9961,N_9256);
nand U10252 (N_10252,N_9245,N_9343);
nand U10253 (N_10253,N_9810,N_9015);
nand U10254 (N_10254,N_9954,N_9175);
and U10255 (N_10255,N_9503,N_9671);
nand U10256 (N_10256,N_9856,N_9691);
and U10257 (N_10257,N_9361,N_9554);
or U10258 (N_10258,N_9823,N_9820);
or U10259 (N_10259,N_9561,N_9488);
and U10260 (N_10260,N_9018,N_9941);
or U10261 (N_10261,N_9461,N_9878);
and U10262 (N_10262,N_9364,N_9644);
and U10263 (N_10263,N_9284,N_9855);
nor U10264 (N_10264,N_9273,N_9577);
and U10265 (N_10265,N_9725,N_9418);
nor U10266 (N_10266,N_9790,N_9995);
and U10267 (N_10267,N_9177,N_9237);
and U10268 (N_10268,N_9969,N_9479);
xnor U10269 (N_10269,N_9893,N_9051);
nor U10270 (N_10270,N_9366,N_9351);
or U10271 (N_10271,N_9039,N_9744);
xnor U10272 (N_10272,N_9811,N_9809);
nor U10273 (N_10273,N_9685,N_9318);
nand U10274 (N_10274,N_9467,N_9807);
or U10275 (N_10275,N_9010,N_9682);
and U10276 (N_10276,N_9930,N_9750);
nor U10277 (N_10277,N_9406,N_9658);
nand U10278 (N_10278,N_9967,N_9829);
nor U10279 (N_10279,N_9761,N_9661);
or U10280 (N_10280,N_9589,N_9996);
and U10281 (N_10281,N_9655,N_9183);
and U10282 (N_10282,N_9702,N_9136);
nor U10283 (N_10283,N_9028,N_9898);
or U10284 (N_10284,N_9866,N_9852);
or U10285 (N_10285,N_9888,N_9737);
or U10286 (N_10286,N_9489,N_9144);
or U10287 (N_10287,N_9269,N_9356);
xor U10288 (N_10288,N_9756,N_9157);
and U10289 (N_10289,N_9432,N_9371);
nand U10290 (N_10290,N_9917,N_9951);
nand U10291 (N_10291,N_9603,N_9298);
and U10292 (N_10292,N_9928,N_9735);
and U10293 (N_10293,N_9551,N_9399);
or U10294 (N_10294,N_9153,N_9411);
xor U10295 (N_10295,N_9113,N_9616);
xnor U10296 (N_10296,N_9957,N_9124);
xnor U10297 (N_10297,N_9544,N_9883);
nor U10298 (N_10298,N_9777,N_9670);
or U10299 (N_10299,N_9910,N_9404);
and U10300 (N_10300,N_9798,N_9277);
xnor U10301 (N_10301,N_9412,N_9977);
xnor U10302 (N_10302,N_9206,N_9034);
xnor U10303 (N_10303,N_9465,N_9221);
nor U10304 (N_10304,N_9999,N_9199);
and U10305 (N_10305,N_9709,N_9048);
nand U10306 (N_10306,N_9050,N_9057);
nor U10307 (N_10307,N_9764,N_9152);
or U10308 (N_10308,N_9550,N_9937);
and U10309 (N_10309,N_9089,N_9389);
or U10310 (N_10310,N_9142,N_9417);
nor U10311 (N_10311,N_9198,N_9581);
and U10312 (N_10312,N_9902,N_9187);
xnor U10313 (N_10313,N_9072,N_9989);
xnor U10314 (N_10314,N_9802,N_9699);
nor U10315 (N_10315,N_9074,N_9580);
xor U10316 (N_10316,N_9537,N_9594);
nor U10317 (N_10317,N_9959,N_9716);
xnor U10318 (N_10318,N_9179,N_9870);
xnor U10319 (N_10319,N_9081,N_9192);
and U10320 (N_10320,N_9458,N_9058);
or U10321 (N_10321,N_9731,N_9285);
xor U10322 (N_10322,N_9442,N_9566);
xor U10323 (N_10323,N_9686,N_9543);
nor U10324 (N_10324,N_9647,N_9363);
nor U10325 (N_10325,N_9516,N_9253);
xnor U10326 (N_10326,N_9988,N_9991);
and U10327 (N_10327,N_9703,N_9078);
nor U10328 (N_10328,N_9723,N_9295);
and U10329 (N_10329,N_9117,N_9299);
and U10330 (N_10330,N_9736,N_9929);
or U10331 (N_10331,N_9583,N_9143);
or U10332 (N_10332,N_9782,N_9713);
xnor U10333 (N_10333,N_9712,N_9617);
xor U10334 (N_10334,N_9456,N_9745);
nor U10335 (N_10335,N_9770,N_9357);
and U10336 (N_10336,N_9978,N_9558);
xor U10337 (N_10337,N_9041,N_9415);
nand U10338 (N_10338,N_9232,N_9330);
nand U10339 (N_10339,N_9684,N_9847);
and U10340 (N_10340,N_9473,N_9975);
nand U10341 (N_10341,N_9979,N_9808);
nand U10342 (N_10342,N_9900,N_9939);
or U10343 (N_10343,N_9815,N_9265);
xor U10344 (N_10344,N_9226,N_9077);
xor U10345 (N_10345,N_9604,N_9955);
or U10346 (N_10346,N_9700,N_9084);
and U10347 (N_10347,N_9444,N_9407);
and U10348 (N_10348,N_9325,N_9453);
nand U10349 (N_10349,N_9292,N_9519);
or U10350 (N_10350,N_9994,N_9787);
and U10351 (N_10351,N_9591,N_9990);
nor U10352 (N_10352,N_9908,N_9114);
and U10353 (N_10353,N_9402,N_9838);
nand U10354 (N_10354,N_9912,N_9097);
nor U10355 (N_10355,N_9186,N_9184);
nor U10356 (N_10356,N_9674,N_9264);
nor U10357 (N_10357,N_9844,N_9190);
or U10358 (N_10358,N_9515,N_9427);
xor U10359 (N_10359,N_9358,N_9992);
and U10360 (N_10360,N_9534,N_9369);
nor U10361 (N_10361,N_9652,N_9695);
or U10362 (N_10362,N_9448,N_9195);
nand U10363 (N_10363,N_9309,N_9664);
xnor U10364 (N_10364,N_9098,N_9567);
or U10365 (N_10365,N_9176,N_9007);
nand U10366 (N_10366,N_9464,N_9772);
nand U10367 (N_10367,N_9746,N_9281);
or U10368 (N_10368,N_9606,N_9196);
nand U10369 (N_10369,N_9332,N_9846);
xor U10370 (N_10370,N_9360,N_9170);
nor U10371 (N_10371,N_9836,N_9643);
nor U10372 (N_10372,N_9833,N_9619);
and U10373 (N_10373,N_9640,N_9431);
nor U10374 (N_10374,N_9832,N_9850);
or U10375 (N_10375,N_9632,N_9443);
or U10376 (N_10376,N_9571,N_9302);
nor U10377 (N_10377,N_9095,N_9568);
or U10378 (N_10378,N_9159,N_9859);
nor U10379 (N_10379,N_9748,N_9793);
xnor U10380 (N_10380,N_9236,N_9239);
xor U10381 (N_10381,N_9896,N_9932);
or U10382 (N_10382,N_9283,N_9188);
nor U10383 (N_10383,N_9499,N_9747);
xnor U10384 (N_10384,N_9327,N_9555);
nor U10385 (N_10385,N_9687,N_9200);
and U10386 (N_10386,N_9172,N_9249);
nor U10387 (N_10387,N_9004,N_9884);
or U10388 (N_10388,N_9005,N_9303);
nand U10389 (N_10389,N_9397,N_9894);
nor U10390 (N_10390,N_9766,N_9031);
and U10391 (N_10391,N_9919,N_9255);
or U10392 (N_10392,N_9657,N_9628);
nor U10393 (N_10393,N_9778,N_9160);
and U10394 (N_10394,N_9019,N_9634);
or U10395 (N_10395,N_9582,N_9246);
or U10396 (N_10396,N_9981,N_9290);
nand U10397 (N_10397,N_9491,N_9964);
nand U10398 (N_10398,N_9552,N_9557);
nand U10399 (N_10399,N_9875,N_9131);
xnor U10400 (N_10400,N_9848,N_9541);
or U10401 (N_10401,N_9784,N_9066);
nand U10402 (N_10402,N_9740,N_9776);
and U10403 (N_10403,N_9436,N_9400);
or U10404 (N_10404,N_9112,N_9660);
or U10405 (N_10405,N_9819,N_9274);
nand U10406 (N_10406,N_9936,N_9393);
or U10407 (N_10407,N_9839,N_9762);
nor U10408 (N_10408,N_9445,N_9368);
xor U10409 (N_10409,N_9457,N_9230);
xnor U10410 (N_10410,N_9899,N_9627);
xnor U10411 (N_10411,N_9252,N_9013);
and U10412 (N_10412,N_9697,N_9504);
or U10413 (N_10413,N_9346,N_9394);
nor U10414 (N_10414,N_9166,N_9874);
xnor U10415 (N_10415,N_9963,N_9732);
nand U10416 (N_10416,N_9570,N_9341);
nand U10417 (N_10417,N_9538,N_9871);
or U10418 (N_10418,N_9104,N_9123);
nor U10419 (N_10419,N_9145,N_9535);
nor U10420 (N_10420,N_9201,N_9642);
and U10421 (N_10421,N_9129,N_9620);
and U10422 (N_10422,N_9765,N_9654);
or U10423 (N_10423,N_9909,N_9507);
or U10424 (N_10424,N_9816,N_9446);
or U10425 (N_10425,N_9288,N_9560);
or U10426 (N_10426,N_9715,N_9441);
nor U10427 (N_10427,N_9425,N_9258);
nand U10428 (N_10428,N_9164,N_9225);
or U10429 (N_10429,N_9906,N_9618);
xor U10430 (N_10430,N_9579,N_9109);
nor U10431 (N_10431,N_9651,N_9387);
xor U10432 (N_10432,N_9986,N_9049);
xor U10433 (N_10433,N_9862,N_9460);
and U10434 (N_10434,N_9549,N_9000);
nor U10435 (N_10435,N_9933,N_9182);
and U10436 (N_10436,N_9155,N_9949);
or U10437 (N_10437,N_9380,N_9372);
xor U10438 (N_10438,N_9203,N_9984);
and U10439 (N_10439,N_9375,N_9052);
and U10440 (N_10440,N_9952,N_9612);
nor U10441 (N_10441,N_9993,N_9849);
nand U10442 (N_10442,N_9711,N_9945);
xor U10443 (N_10443,N_9297,N_9704);
or U10444 (N_10444,N_9597,N_9151);
xor U10445 (N_10445,N_9428,N_9636);
nor U10446 (N_10446,N_9304,N_9564);
xnor U10447 (N_10447,N_9841,N_9423);
or U10448 (N_10448,N_9308,N_9997);
xor U10449 (N_10449,N_9546,N_9217);
and U10450 (N_10450,N_9976,N_9864);
xnor U10451 (N_10451,N_9280,N_9373);
and U10452 (N_10452,N_9025,N_9690);
or U10453 (N_10453,N_9282,N_9055);
nand U10454 (N_10454,N_9275,N_9042);
xnor U10455 (N_10455,N_9266,N_9601);
or U10456 (N_10456,N_9323,N_9895);
nor U10457 (N_10457,N_9092,N_9548);
and U10458 (N_10458,N_9108,N_9563);
nor U10459 (N_10459,N_9293,N_9434);
xor U10460 (N_10460,N_9468,N_9623);
nand U10461 (N_10461,N_9215,N_9272);
nand U10462 (N_10462,N_9783,N_9759);
nor U10463 (N_10463,N_9701,N_9598);
xor U10464 (N_10464,N_9047,N_9751);
nand U10465 (N_10465,N_9228,N_9645);
nor U10466 (N_10466,N_9972,N_9858);
nor U10467 (N_10467,N_9122,N_9724);
or U10468 (N_10468,N_9477,N_9749);
xor U10469 (N_10469,N_9405,N_9338);
and U10470 (N_10470,N_9705,N_9126);
or U10471 (N_10471,N_9739,N_9925);
nor U10472 (N_10472,N_9021,N_9342);
xnor U10473 (N_10473,N_9064,N_9162);
or U10474 (N_10474,N_9045,N_9931);
and U10475 (N_10475,N_9305,N_9377);
nand U10476 (N_10476,N_9611,N_9022);
and U10477 (N_10477,N_9137,N_9629);
or U10478 (N_10478,N_9403,N_9454);
or U10479 (N_10479,N_9450,N_9345);
nand U10480 (N_10480,N_9834,N_9797);
nand U10481 (N_10481,N_9120,N_9663);
and U10482 (N_10482,N_9067,N_9319);
nand U10483 (N_10483,N_9918,N_9094);
and U10484 (N_10484,N_9610,N_9241);
and U10485 (N_10485,N_9860,N_9801);
or U10486 (N_10486,N_9213,N_9633);
and U10487 (N_10487,N_9608,N_9365);
nor U10488 (N_10488,N_9312,N_9650);
and U10489 (N_10489,N_9805,N_9469);
nor U10490 (N_10490,N_9678,N_9966);
or U10491 (N_10491,N_9944,N_9915);
and U10492 (N_10492,N_9233,N_9854);
nor U10493 (N_10493,N_9677,N_9248);
nor U10494 (N_10494,N_9033,N_9030);
or U10495 (N_10495,N_9056,N_9231);
or U10496 (N_10496,N_9624,N_9683);
nor U10497 (N_10497,N_9814,N_9907);
and U10498 (N_10498,N_9219,N_9903);
xnor U10499 (N_10499,N_9060,N_9646);
nand U10500 (N_10500,N_9154,N_9540);
or U10501 (N_10501,N_9040,N_9098);
or U10502 (N_10502,N_9438,N_9038);
nand U10503 (N_10503,N_9485,N_9045);
and U10504 (N_10504,N_9639,N_9651);
and U10505 (N_10505,N_9522,N_9600);
or U10506 (N_10506,N_9017,N_9687);
nand U10507 (N_10507,N_9918,N_9106);
or U10508 (N_10508,N_9587,N_9431);
xor U10509 (N_10509,N_9071,N_9966);
xnor U10510 (N_10510,N_9556,N_9493);
xor U10511 (N_10511,N_9333,N_9462);
nand U10512 (N_10512,N_9153,N_9475);
nand U10513 (N_10513,N_9329,N_9917);
nand U10514 (N_10514,N_9340,N_9159);
and U10515 (N_10515,N_9993,N_9458);
nand U10516 (N_10516,N_9870,N_9468);
or U10517 (N_10517,N_9157,N_9115);
nand U10518 (N_10518,N_9092,N_9002);
nor U10519 (N_10519,N_9400,N_9991);
or U10520 (N_10520,N_9066,N_9341);
and U10521 (N_10521,N_9616,N_9365);
nand U10522 (N_10522,N_9771,N_9440);
xor U10523 (N_10523,N_9830,N_9368);
or U10524 (N_10524,N_9745,N_9987);
or U10525 (N_10525,N_9561,N_9265);
or U10526 (N_10526,N_9717,N_9826);
xor U10527 (N_10527,N_9576,N_9332);
nand U10528 (N_10528,N_9874,N_9555);
and U10529 (N_10529,N_9731,N_9269);
nor U10530 (N_10530,N_9574,N_9745);
nand U10531 (N_10531,N_9689,N_9321);
nor U10532 (N_10532,N_9877,N_9508);
nor U10533 (N_10533,N_9975,N_9775);
or U10534 (N_10534,N_9691,N_9002);
nand U10535 (N_10535,N_9561,N_9199);
and U10536 (N_10536,N_9886,N_9759);
nor U10537 (N_10537,N_9059,N_9529);
and U10538 (N_10538,N_9365,N_9923);
nor U10539 (N_10539,N_9463,N_9676);
nor U10540 (N_10540,N_9373,N_9346);
xnor U10541 (N_10541,N_9625,N_9718);
or U10542 (N_10542,N_9961,N_9822);
and U10543 (N_10543,N_9187,N_9161);
nor U10544 (N_10544,N_9162,N_9034);
and U10545 (N_10545,N_9415,N_9034);
nand U10546 (N_10546,N_9512,N_9178);
and U10547 (N_10547,N_9855,N_9803);
nand U10548 (N_10548,N_9525,N_9787);
or U10549 (N_10549,N_9751,N_9829);
nand U10550 (N_10550,N_9844,N_9984);
nand U10551 (N_10551,N_9003,N_9610);
nor U10552 (N_10552,N_9565,N_9771);
and U10553 (N_10553,N_9614,N_9075);
xor U10554 (N_10554,N_9888,N_9552);
nor U10555 (N_10555,N_9927,N_9398);
xor U10556 (N_10556,N_9438,N_9276);
nor U10557 (N_10557,N_9146,N_9171);
nor U10558 (N_10558,N_9447,N_9975);
or U10559 (N_10559,N_9790,N_9944);
nand U10560 (N_10560,N_9717,N_9362);
or U10561 (N_10561,N_9027,N_9255);
nor U10562 (N_10562,N_9622,N_9367);
xor U10563 (N_10563,N_9478,N_9768);
and U10564 (N_10564,N_9421,N_9466);
and U10565 (N_10565,N_9449,N_9597);
nand U10566 (N_10566,N_9034,N_9148);
nand U10567 (N_10567,N_9672,N_9503);
and U10568 (N_10568,N_9792,N_9152);
nand U10569 (N_10569,N_9664,N_9310);
nand U10570 (N_10570,N_9993,N_9056);
or U10571 (N_10571,N_9619,N_9708);
and U10572 (N_10572,N_9112,N_9669);
and U10573 (N_10573,N_9317,N_9800);
and U10574 (N_10574,N_9834,N_9603);
nand U10575 (N_10575,N_9323,N_9333);
xnor U10576 (N_10576,N_9205,N_9671);
nand U10577 (N_10577,N_9998,N_9597);
and U10578 (N_10578,N_9575,N_9267);
or U10579 (N_10579,N_9815,N_9714);
and U10580 (N_10580,N_9372,N_9401);
nor U10581 (N_10581,N_9706,N_9850);
nand U10582 (N_10582,N_9281,N_9708);
nand U10583 (N_10583,N_9999,N_9383);
nand U10584 (N_10584,N_9045,N_9249);
nor U10585 (N_10585,N_9469,N_9097);
xnor U10586 (N_10586,N_9042,N_9383);
nand U10587 (N_10587,N_9921,N_9756);
and U10588 (N_10588,N_9387,N_9172);
xor U10589 (N_10589,N_9213,N_9510);
or U10590 (N_10590,N_9876,N_9167);
xor U10591 (N_10591,N_9456,N_9628);
and U10592 (N_10592,N_9462,N_9890);
and U10593 (N_10593,N_9187,N_9534);
and U10594 (N_10594,N_9225,N_9092);
xor U10595 (N_10595,N_9742,N_9896);
and U10596 (N_10596,N_9276,N_9787);
nor U10597 (N_10597,N_9890,N_9217);
and U10598 (N_10598,N_9061,N_9437);
nand U10599 (N_10599,N_9439,N_9862);
nand U10600 (N_10600,N_9484,N_9094);
nor U10601 (N_10601,N_9379,N_9201);
or U10602 (N_10602,N_9774,N_9513);
nand U10603 (N_10603,N_9016,N_9027);
or U10604 (N_10604,N_9250,N_9886);
nand U10605 (N_10605,N_9907,N_9054);
xor U10606 (N_10606,N_9915,N_9374);
or U10607 (N_10607,N_9395,N_9725);
xor U10608 (N_10608,N_9249,N_9369);
and U10609 (N_10609,N_9758,N_9502);
xor U10610 (N_10610,N_9617,N_9682);
and U10611 (N_10611,N_9849,N_9900);
nor U10612 (N_10612,N_9845,N_9822);
or U10613 (N_10613,N_9079,N_9640);
or U10614 (N_10614,N_9797,N_9513);
or U10615 (N_10615,N_9702,N_9623);
or U10616 (N_10616,N_9112,N_9860);
or U10617 (N_10617,N_9089,N_9337);
xnor U10618 (N_10618,N_9686,N_9237);
and U10619 (N_10619,N_9731,N_9000);
and U10620 (N_10620,N_9185,N_9748);
xnor U10621 (N_10621,N_9827,N_9552);
nand U10622 (N_10622,N_9982,N_9583);
or U10623 (N_10623,N_9213,N_9419);
nor U10624 (N_10624,N_9259,N_9543);
nor U10625 (N_10625,N_9848,N_9654);
xor U10626 (N_10626,N_9143,N_9008);
nor U10627 (N_10627,N_9136,N_9510);
and U10628 (N_10628,N_9719,N_9253);
nand U10629 (N_10629,N_9772,N_9617);
and U10630 (N_10630,N_9632,N_9308);
nand U10631 (N_10631,N_9672,N_9325);
and U10632 (N_10632,N_9707,N_9824);
nand U10633 (N_10633,N_9061,N_9193);
nand U10634 (N_10634,N_9703,N_9718);
nand U10635 (N_10635,N_9863,N_9092);
nand U10636 (N_10636,N_9470,N_9678);
nand U10637 (N_10637,N_9879,N_9934);
nor U10638 (N_10638,N_9382,N_9915);
xor U10639 (N_10639,N_9652,N_9666);
xnor U10640 (N_10640,N_9257,N_9953);
nand U10641 (N_10641,N_9093,N_9868);
nor U10642 (N_10642,N_9217,N_9876);
nand U10643 (N_10643,N_9791,N_9883);
nor U10644 (N_10644,N_9988,N_9631);
nand U10645 (N_10645,N_9451,N_9463);
xnor U10646 (N_10646,N_9063,N_9709);
and U10647 (N_10647,N_9122,N_9074);
nor U10648 (N_10648,N_9975,N_9860);
nand U10649 (N_10649,N_9751,N_9561);
xnor U10650 (N_10650,N_9781,N_9577);
nand U10651 (N_10651,N_9747,N_9107);
or U10652 (N_10652,N_9852,N_9449);
xor U10653 (N_10653,N_9770,N_9294);
nand U10654 (N_10654,N_9930,N_9573);
nor U10655 (N_10655,N_9560,N_9407);
nand U10656 (N_10656,N_9159,N_9735);
nand U10657 (N_10657,N_9029,N_9422);
and U10658 (N_10658,N_9972,N_9829);
and U10659 (N_10659,N_9048,N_9304);
or U10660 (N_10660,N_9048,N_9188);
and U10661 (N_10661,N_9734,N_9001);
or U10662 (N_10662,N_9350,N_9619);
nor U10663 (N_10663,N_9441,N_9362);
xor U10664 (N_10664,N_9341,N_9258);
and U10665 (N_10665,N_9924,N_9709);
xor U10666 (N_10666,N_9696,N_9935);
or U10667 (N_10667,N_9810,N_9750);
and U10668 (N_10668,N_9728,N_9971);
nor U10669 (N_10669,N_9520,N_9467);
nand U10670 (N_10670,N_9004,N_9965);
nor U10671 (N_10671,N_9089,N_9429);
or U10672 (N_10672,N_9832,N_9559);
nand U10673 (N_10673,N_9711,N_9538);
and U10674 (N_10674,N_9476,N_9634);
nor U10675 (N_10675,N_9180,N_9492);
nand U10676 (N_10676,N_9527,N_9051);
or U10677 (N_10677,N_9687,N_9432);
or U10678 (N_10678,N_9321,N_9441);
or U10679 (N_10679,N_9498,N_9107);
xnor U10680 (N_10680,N_9110,N_9585);
nand U10681 (N_10681,N_9055,N_9555);
nor U10682 (N_10682,N_9882,N_9742);
and U10683 (N_10683,N_9376,N_9733);
xor U10684 (N_10684,N_9857,N_9738);
and U10685 (N_10685,N_9894,N_9364);
or U10686 (N_10686,N_9299,N_9815);
nand U10687 (N_10687,N_9229,N_9107);
nand U10688 (N_10688,N_9579,N_9554);
nand U10689 (N_10689,N_9365,N_9397);
or U10690 (N_10690,N_9416,N_9855);
nand U10691 (N_10691,N_9219,N_9168);
or U10692 (N_10692,N_9835,N_9412);
nor U10693 (N_10693,N_9458,N_9861);
nor U10694 (N_10694,N_9669,N_9261);
and U10695 (N_10695,N_9088,N_9297);
or U10696 (N_10696,N_9150,N_9412);
or U10697 (N_10697,N_9692,N_9353);
nor U10698 (N_10698,N_9965,N_9072);
xnor U10699 (N_10699,N_9568,N_9251);
nor U10700 (N_10700,N_9971,N_9537);
or U10701 (N_10701,N_9992,N_9133);
and U10702 (N_10702,N_9406,N_9758);
or U10703 (N_10703,N_9789,N_9864);
nand U10704 (N_10704,N_9060,N_9491);
nor U10705 (N_10705,N_9194,N_9581);
xnor U10706 (N_10706,N_9573,N_9078);
or U10707 (N_10707,N_9901,N_9159);
xnor U10708 (N_10708,N_9219,N_9115);
xor U10709 (N_10709,N_9310,N_9770);
xor U10710 (N_10710,N_9681,N_9233);
and U10711 (N_10711,N_9674,N_9628);
and U10712 (N_10712,N_9952,N_9778);
xnor U10713 (N_10713,N_9050,N_9526);
nand U10714 (N_10714,N_9577,N_9023);
and U10715 (N_10715,N_9179,N_9078);
nor U10716 (N_10716,N_9838,N_9202);
nor U10717 (N_10717,N_9297,N_9882);
and U10718 (N_10718,N_9117,N_9730);
nand U10719 (N_10719,N_9360,N_9632);
or U10720 (N_10720,N_9213,N_9581);
nor U10721 (N_10721,N_9668,N_9633);
or U10722 (N_10722,N_9972,N_9228);
nand U10723 (N_10723,N_9242,N_9899);
nor U10724 (N_10724,N_9154,N_9334);
or U10725 (N_10725,N_9925,N_9193);
nand U10726 (N_10726,N_9607,N_9431);
nand U10727 (N_10727,N_9567,N_9857);
and U10728 (N_10728,N_9286,N_9516);
nor U10729 (N_10729,N_9956,N_9423);
or U10730 (N_10730,N_9802,N_9066);
and U10731 (N_10731,N_9103,N_9601);
xor U10732 (N_10732,N_9771,N_9296);
xor U10733 (N_10733,N_9070,N_9263);
and U10734 (N_10734,N_9128,N_9512);
or U10735 (N_10735,N_9965,N_9784);
xnor U10736 (N_10736,N_9815,N_9442);
nand U10737 (N_10737,N_9788,N_9670);
nor U10738 (N_10738,N_9315,N_9264);
nand U10739 (N_10739,N_9489,N_9573);
xnor U10740 (N_10740,N_9495,N_9084);
nand U10741 (N_10741,N_9683,N_9464);
xnor U10742 (N_10742,N_9931,N_9057);
and U10743 (N_10743,N_9547,N_9052);
or U10744 (N_10744,N_9747,N_9529);
or U10745 (N_10745,N_9913,N_9473);
nor U10746 (N_10746,N_9924,N_9329);
nand U10747 (N_10747,N_9124,N_9437);
nand U10748 (N_10748,N_9695,N_9125);
and U10749 (N_10749,N_9956,N_9643);
or U10750 (N_10750,N_9218,N_9744);
or U10751 (N_10751,N_9411,N_9230);
and U10752 (N_10752,N_9366,N_9462);
xor U10753 (N_10753,N_9311,N_9537);
or U10754 (N_10754,N_9103,N_9812);
nand U10755 (N_10755,N_9380,N_9214);
xor U10756 (N_10756,N_9899,N_9549);
or U10757 (N_10757,N_9915,N_9421);
or U10758 (N_10758,N_9885,N_9573);
xor U10759 (N_10759,N_9247,N_9978);
and U10760 (N_10760,N_9808,N_9727);
and U10761 (N_10761,N_9093,N_9707);
nor U10762 (N_10762,N_9959,N_9674);
nand U10763 (N_10763,N_9885,N_9997);
or U10764 (N_10764,N_9404,N_9893);
xor U10765 (N_10765,N_9618,N_9550);
or U10766 (N_10766,N_9898,N_9526);
and U10767 (N_10767,N_9754,N_9019);
nor U10768 (N_10768,N_9359,N_9139);
or U10769 (N_10769,N_9509,N_9581);
nor U10770 (N_10770,N_9143,N_9704);
or U10771 (N_10771,N_9949,N_9153);
nor U10772 (N_10772,N_9074,N_9314);
xor U10773 (N_10773,N_9527,N_9927);
nor U10774 (N_10774,N_9664,N_9995);
nor U10775 (N_10775,N_9080,N_9615);
and U10776 (N_10776,N_9543,N_9168);
or U10777 (N_10777,N_9827,N_9176);
nor U10778 (N_10778,N_9013,N_9496);
xnor U10779 (N_10779,N_9295,N_9115);
nor U10780 (N_10780,N_9495,N_9203);
and U10781 (N_10781,N_9862,N_9744);
xnor U10782 (N_10782,N_9202,N_9622);
or U10783 (N_10783,N_9260,N_9978);
and U10784 (N_10784,N_9714,N_9154);
or U10785 (N_10785,N_9969,N_9652);
or U10786 (N_10786,N_9583,N_9970);
and U10787 (N_10787,N_9445,N_9809);
xor U10788 (N_10788,N_9165,N_9960);
xnor U10789 (N_10789,N_9251,N_9081);
nand U10790 (N_10790,N_9956,N_9866);
nand U10791 (N_10791,N_9755,N_9922);
or U10792 (N_10792,N_9540,N_9549);
or U10793 (N_10793,N_9795,N_9200);
nor U10794 (N_10794,N_9478,N_9385);
or U10795 (N_10795,N_9010,N_9400);
nand U10796 (N_10796,N_9046,N_9370);
nor U10797 (N_10797,N_9628,N_9328);
and U10798 (N_10798,N_9210,N_9013);
nand U10799 (N_10799,N_9812,N_9891);
xor U10800 (N_10800,N_9482,N_9565);
or U10801 (N_10801,N_9940,N_9356);
xnor U10802 (N_10802,N_9504,N_9579);
nor U10803 (N_10803,N_9442,N_9736);
nor U10804 (N_10804,N_9396,N_9129);
xor U10805 (N_10805,N_9180,N_9317);
or U10806 (N_10806,N_9095,N_9164);
or U10807 (N_10807,N_9836,N_9005);
or U10808 (N_10808,N_9880,N_9310);
and U10809 (N_10809,N_9373,N_9334);
nand U10810 (N_10810,N_9078,N_9995);
nor U10811 (N_10811,N_9377,N_9046);
nor U10812 (N_10812,N_9602,N_9656);
nor U10813 (N_10813,N_9956,N_9605);
xor U10814 (N_10814,N_9776,N_9712);
xnor U10815 (N_10815,N_9890,N_9554);
xor U10816 (N_10816,N_9001,N_9648);
or U10817 (N_10817,N_9953,N_9205);
nand U10818 (N_10818,N_9434,N_9457);
nand U10819 (N_10819,N_9843,N_9916);
or U10820 (N_10820,N_9374,N_9159);
or U10821 (N_10821,N_9147,N_9821);
xnor U10822 (N_10822,N_9201,N_9008);
nand U10823 (N_10823,N_9105,N_9125);
nand U10824 (N_10824,N_9927,N_9561);
nand U10825 (N_10825,N_9749,N_9109);
and U10826 (N_10826,N_9093,N_9558);
and U10827 (N_10827,N_9235,N_9319);
or U10828 (N_10828,N_9410,N_9291);
or U10829 (N_10829,N_9069,N_9004);
and U10830 (N_10830,N_9667,N_9180);
and U10831 (N_10831,N_9335,N_9063);
nand U10832 (N_10832,N_9809,N_9335);
nor U10833 (N_10833,N_9102,N_9976);
nor U10834 (N_10834,N_9086,N_9259);
nand U10835 (N_10835,N_9838,N_9299);
nor U10836 (N_10836,N_9218,N_9809);
nand U10837 (N_10837,N_9084,N_9244);
nand U10838 (N_10838,N_9624,N_9474);
xnor U10839 (N_10839,N_9407,N_9464);
nand U10840 (N_10840,N_9701,N_9563);
nand U10841 (N_10841,N_9715,N_9403);
or U10842 (N_10842,N_9342,N_9636);
nand U10843 (N_10843,N_9481,N_9636);
nand U10844 (N_10844,N_9303,N_9249);
and U10845 (N_10845,N_9528,N_9479);
and U10846 (N_10846,N_9795,N_9620);
nand U10847 (N_10847,N_9676,N_9014);
or U10848 (N_10848,N_9098,N_9700);
nand U10849 (N_10849,N_9307,N_9522);
xor U10850 (N_10850,N_9500,N_9869);
nand U10851 (N_10851,N_9954,N_9284);
nor U10852 (N_10852,N_9902,N_9354);
nor U10853 (N_10853,N_9729,N_9526);
xnor U10854 (N_10854,N_9528,N_9881);
or U10855 (N_10855,N_9218,N_9758);
or U10856 (N_10856,N_9669,N_9088);
and U10857 (N_10857,N_9592,N_9149);
and U10858 (N_10858,N_9634,N_9517);
nand U10859 (N_10859,N_9634,N_9516);
or U10860 (N_10860,N_9994,N_9814);
nor U10861 (N_10861,N_9818,N_9231);
xnor U10862 (N_10862,N_9845,N_9328);
or U10863 (N_10863,N_9841,N_9406);
or U10864 (N_10864,N_9136,N_9452);
xnor U10865 (N_10865,N_9910,N_9986);
nand U10866 (N_10866,N_9349,N_9435);
xor U10867 (N_10867,N_9161,N_9930);
xor U10868 (N_10868,N_9813,N_9438);
xnor U10869 (N_10869,N_9625,N_9386);
nand U10870 (N_10870,N_9007,N_9342);
or U10871 (N_10871,N_9414,N_9832);
nor U10872 (N_10872,N_9589,N_9655);
nor U10873 (N_10873,N_9162,N_9905);
or U10874 (N_10874,N_9653,N_9324);
nor U10875 (N_10875,N_9270,N_9578);
xnor U10876 (N_10876,N_9048,N_9164);
nor U10877 (N_10877,N_9902,N_9739);
nand U10878 (N_10878,N_9893,N_9273);
or U10879 (N_10879,N_9524,N_9617);
xor U10880 (N_10880,N_9258,N_9547);
nand U10881 (N_10881,N_9212,N_9899);
and U10882 (N_10882,N_9803,N_9760);
or U10883 (N_10883,N_9383,N_9882);
nor U10884 (N_10884,N_9729,N_9033);
nor U10885 (N_10885,N_9281,N_9484);
nand U10886 (N_10886,N_9153,N_9518);
nor U10887 (N_10887,N_9366,N_9775);
xor U10888 (N_10888,N_9865,N_9178);
nor U10889 (N_10889,N_9231,N_9000);
nand U10890 (N_10890,N_9624,N_9478);
and U10891 (N_10891,N_9698,N_9919);
nand U10892 (N_10892,N_9654,N_9450);
xor U10893 (N_10893,N_9592,N_9563);
xnor U10894 (N_10894,N_9231,N_9280);
nand U10895 (N_10895,N_9881,N_9998);
nor U10896 (N_10896,N_9580,N_9924);
xor U10897 (N_10897,N_9485,N_9209);
nor U10898 (N_10898,N_9022,N_9625);
nor U10899 (N_10899,N_9858,N_9086);
xor U10900 (N_10900,N_9874,N_9346);
xnor U10901 (N_10901,N_9766,N_9870);
or U10902 (N_10902,N_9374,N_9353);
xor U10903 (N_10903,N_9144,N_9609);
nor U10904 (N_10904,N_9015,N_9957);
xnor U10905 (N_10905,N_9882,N_9092);
xor U10906 (N_10906,N_9000,N_9728);
nand U10907 (N_10907,N_9251,N_9740);
nand U10908 (N_10908,N_9650,N_9277);
nand U10909 (N_10909,N_9611,N_9054);
nor U10910 (N_10910,N_9254,N_9672);
xor U10911 (N_10911,N_9950,N_9082);
nor U10912 (N_10912,N_9838,N_9886);
and U10913 (N_10913,N_9612,N_9426);
nand U10914 (N_10914,N_9778,N_9488);
nor U10915 (N_10915,N_9107,N_9068);
nand U10916 (N_10916,N_9351,N_9474);
or U10917 (N_10917,N_9546,N_9901);
or U10918 (N_10918,N_9105,N_9611);
and U10919 (N_10919,N_9100,N_9560);
or U10920 (N_10920,N_9719,N_9790);
and U10921 (N_10921,N_9500,N_9112);
and U10922 (N_10922,N_9828,N_9245);
nand U10923 (N_10923,N_9276,N_9465);
xnor U10924 (N_10924,N_9964,N_9139);
nand U10925 (N_10925,N_9108,N_9811);
or U10926 (N_10926,N_9148,N_9881);
nor U10927 (N_10927,N_9690,N_9428);
or U10928 (N_10928,N_9631,N_9425);
xnor U10929 (N_10929,N_9548,N_9897);
and U10930 (N_10930,N_9009,N_9337);
and U10931 (N_10931,N_9312,N_9674);
or U10932 (N_10932,N_9070,N_9949);
xor U10933 (N_10933,N_9620,N_9656);
or U10934 (N_10934,N_9048,N_9265);
and U10935 (N_10935,N_9382,N_9379);
or U10936 (N_10936,N_9689,N_9135);
xnor U10937 (N_10937,N_9349,N_9114);
and U10938 (N_10938,N_9571,N_9882);
nand U10939 (N_10939,N_9005,N_9589);
and U10940 (N_10940,N_9656,N_9553);
and U10941 (N_10941,N_9141,N_9308);
and U10942 (N_10942,N_9456,N_9545);
xor U10943 (N_10943,N_9713,N_9566);
or U10944 (N_10944,N_9734,N_9492);
xor U10945 (N_10945,N_9214,N_9821);
nor U10946 (N_10946,N_9424,N_9263);
and U10947 (N_10947,N_9191,N_9563);
nor U10948 (N_10948,N_9560,N_9772);
nand U10949 (N_10949,N_9034,N_9543);
nand U10950 (N_10950,N_9867,N_9199);
nor U10951 (N_10951,N_9433,N_9720);
nand U10952 (N_10952,N_9579,N_9555);
nand U10953 (N_10953,N_9553,N_9088);
nand U10954 (N_10954,N_9873,N_9166);
nor U10955 (N_10955,N_9913,N_9716);
nand U10956 (N_10956,N_9966,N_9381);
or U10957 (N_10957,N_9005,N_9823);
nor U10958 (N_10958,N_9906,N_9162);
xnor U10959 (N_10959,N_9572,N_9286);
xor U10960 (N_10960,N_9743,N_9552);
xnor U10961 (N_10961,N_9365,N_9367);
xor U10962 (N_10962,N_9475,N_9008);
nor U10963 (N_10963,N_9190,N_9037);
xor U10964 (N_10964,N_9144,N_9968);
nor U10965 (N_10965,N_9578,N_9255);
and U10966 (N_10966,N_9525,N_9821);
xnor U10967 (N_10967,N_9042,N_9839);
xnor U10968 (N_10968,N_9389,N_9245);
xor U10969 (N_10969,N_9389,N_9206);
nand U10970 (N_10970,N_9923,N_9902);
nor U10971 (N_10971,N_9411,N_9623);
and U10972 (N_10972,N_9895,N_9230);
nand U10973 (N_10973,N_9247,N_9906);
or U10974 (N_10974,N_9141,N_9154);
nor U10975 (N_10975,N_9227,N_9569);
and U10976 (N_10976,N_9564,N_9370);
and U10977 (N_10977,N_9582,N_9860);
xor U10978 (N_10978,N_9555,N_9240);
or U10979 (N_10979,N_9304,N_9166);
nor U10980 (N_10980,N_9546,N_9393);
or U10981 (N_10981,N_9402,N_9126);
or U10982 (N_10982,N_9142,N_9637);
xor U10983 (N_10983,N_9963,N_9176);
xor U10984 (N_10984,N_9684,N_9682);
nor U10985 (N_10985,N_9980,N_9049);
nor U10986 (N_10986,N_9800,N_9703);
or U10987 (N_10987,N_9024,N_9239);
or U10988 (N_10988,N_9888,N_9212);
and U10989 (N_10989,N_9107,N_9297);
or U10990 (N_10990,N_9143,N_9762);
xnor U10991 (N_10991,N_9113,N_9457);
nand U10992 (N_10992,N_9896,N_9604);
nor U10993 (N_10993,N_9171,N_9060);
or U10994 (N_10994,N_9223,N_9161);
nor U10995 (N_10995,N_9409,N_9519);
nor U10996 (N_10996,N_9265,N_9267);
and U10997 (N_10997,N_9458,N_9503);
or U10998 (N_10998,N_9910,N_9274);
and U10999 (N_10999,N_9273,N_9452);
xnor U11000 (N_11000,N_10705,N_10404);
nand U11001 (N_11001,N_10952,N_10296);
nand U11002 (N_11002,N_10895,N_10996);
or U11003 (N_11003,N_10077,N_10676);
nand U11004 (N_11004,N_10392,N_10401);
or U11005 (N_11005,N_10968,N_10416);
nor U11006 (N_11006,N_10728,N_10292);
or U11007 (N_11007,N_10935,N_10500);
nor U11008 (N_11008,N_10125,N_10736);
xor U11009 (N_11009,N_10320,N_10408);
and U11010 (N_11010,N_10235,N_10467);
or U11011 (N_11011,N_10661,N_10974);
xnor U11012 (N_11012,N_10941,N_10424);
nor U11013 (N_11013,N_10759,N_10236);
nor U11014 (N_11014,N_10315,N_10792);
or U11015 (N_11015,N_10999,N_10619);
nand U11016 (N_11016,N_10490,N_10695);
xnor U11017 (N_11017,N_10382,N_10609);
or U11018 (N_11018,N_10568,N_10923);
xnor U11019 (N_11019,N_10215,N_10354);
or U11020 (N_11020,N_10272,N_10722);
xnor U11021 (N_11021,N_10946,N_10209);
or U11022 (N_11022,N_10868,N_10945);
nor U11023 (N_11023,N_10993,N_10270);
and U11024 (N_11024,N_10387,N_10169);
nor U11025 (N_11025,N_10233,N_10506);
or U11026 (N_11026,N_10052,N_10116);
xor U11027 (N_11027,N_10561,N_10028);
xnor U11028 (N_11028,N_10822,N_10029);
nand U11029 (N_11029,N_10217,N_10083);
nor U11030 (N_11030,N_10297,N_10636);
xnor U11031 (N_11031,N_10326,N_10281);
and U11032 (N_11032,N_10943,N_10111);
nand U11033 (N_11033,N_10495,N_10585);
nand U11034 (N_11034,N_10237,N_10606);
xnor U11035 (N_11035,N_10892,N_10815);
and U11036 (N_11036,N_10406,N_10551);
or U11037 (N_11037,N_10790,N_10214);
and U11038 (N_11038,N_10545,N_10699);
xor U11039 (N_11039,N_10266,N_10223);
or U11040 (N_11040,N_10452,N_10095);
nor U11041 (N_11041,N_10801,N_10906);
and U11042 (N_11042,N_10578,N_10374);
nor U11043 (N_11043,N_10924,N_10574);
nand U11044 (N_11044,N_10159,N_10626);
nor U11045 (N_11045,N_10625,N_10091);
xnor U11046 (N_11046,N_10510,N_10087);
nand U11047 (N_11047,N_10536,N_10316);
xnor U11048 (N_11048,N_10793,N_10967);
xor U11049 (N_11049,N_10668,N_10024);
xor U11050 (N_11050,N_10836,N_10934);
or U11051 (N_11051,N_10030,N_10082);
nand U11052 (N_11052,N_10644,N_10937);
nand U11053 (N_11053,N_10716,N_10352);
or U11054 (N_11054,N_10157,N_10365);
nand U11055 (N_11055,N_10958,N_10818);
nor U11056 (N_11056,N_10837,N_10718);
or U11057 (N_11057,N_10012,N_10537);
or U11058 (N_11058,N_10673,N_10770);
or U11059 (N_11059,N_10980,N_10757);
or U11060 (N_11060,N_10805,N_10620);
and U11061 (N_11061,N_10966,N_10624);
xor U11062 (N_11062,N_10927,N_10114);
xor U11063 (N_11063,N_10437,N_10804);
or U11064 (N_11064,N_10991,N_10998);
nor U11065 (N_11065,N_10230,N_10848);
and U11066 (N_11066,N_10959,N_10711);
or U11067 (N_11067,N_10696,N_10194);
nor U11068 (N_11068,N_10954,N_10747);
nor U11069 (N_11069,N_10575,N_10552);
xnor U11070 (N_11070,N_10810,N_10202);
and U11071 (N_11071,N_10242,N_10861);
or U11072 (N_11072,N_10745,N_10459);
or U11073 (N_11073,N_10838,N_10762);
nand U11074 (N_11074,N_10364,N_10827);
xnor U11075 (N_11075,N_10834,N_10454);
and U11076 (N_11076,N_10148,N_10262);
nor U11077 (N_11077,N_10803,N_10504);
and U11078 (N_11078,N_10328,N_10294);
and U11079 (N_11079,N_10957,N_10948);
or U11080 (N_11080,N_10807,N_10756);
xnor U11081 (N_11081,N_10713,N_10174);
and U11082 (N_11082,N_10698,N_10345);
xnor U11083 (N_11083,N_10391,N_10766);
or U11084 (N_11084,N_10285,N_10896);
and U11085 (N_11085,N_10278,N_10851);
nand U11086 (N_11086,N_10309,N_10332);
nand U11087 (N_11087,N_10652,N_10257);
and U11088 (N_11088,N_10965,N_10357);
nand U11089 (N_11089,N_10630,N_10327);
nor U11090 (N_11090,N_10254,N_10465);
nand U11091 (N_11091,N_10127,N_10780);
nor U11092 (N_11092,N_10498,N_10334);
or U11093 (N_11093,N_10146,N_10022);
xnor U11094 (N_11094,N_10553,N_10201);
and U11095 (N_11095,N_10592,N_10156);
xor U11096 (N_11096,N_10068,N_10462);
xor U11097 (N_11097,N_10386,N_10884);
and U11098 (N_11098,N_10246,N_10640);
and U11099 (N_11099,N_10003,N_10261);
or U11100 (N_11100,N_10450,N_10092);
or U11101 (N_11101,N_10155,N_10020);
and U11102 (N_11102,N_10341,N_10191);
nor U11103 (N_11103,N_10724,N_10050);
xnor U11104 (N_11104,N_10653,N_10494);
xor U11105 (N_11105,N_10066,N_10213);
nand U11106 (N_11106,N_10632,N_10007);
nand U11107 (N_11107,N_10337,N_10989);
nor U11108 (N_11108,N_10306,N_10950);
or U11109 (N_11109,N_10182,N_10754);
nand U11110 (N_11110,N_10026,N_10623);
nand U11111 (N_11111,N_10346,N_10583);
and U11112 (N_11112,N_10514,N_10388);
nand U11113 (N_11113,N_10929,N_10389);
nor U11114 (N_11114,N_10918,N_10046);
or U11115 (N_11115,N_10889,N_10817);
xor U11116 (N_11116,N_10516,N_10013);
xnor U11117 (N_11117,N_10176,N_10683);
or U11118 (N_11118,N_10515,N_10751);
nor U11119 (N_11119,N_10276,N_10723);
nand U11120 (N_11120,N_10897,N_10582);
xnor U11121 (N_11121,N_10249,N_10166);
xnor U11122 (N_11122,N_10032,N_10813);
or U11123 (N_11123,N_10163,N_10308);
nand U11124 (N_11124,N_10329,N_10882);
nand U11125 (N_11125,N_10840,N_10369);
and U11126 (N_11126,N_10288,N_10375);
nor U11127 (N_11127,N_10821,N_10547);
or U11128 (N_11128,N_10005,N_10115);
nand U11129 (N_11129,N_10360,N_10611);
or U11130 (N_11130,N_10137,N_10691);
xnor U11131 (N_11131,N_10660,N_10422);
nand U11132 (N_11132,N_10844,N_10232);
nor U11133 (N_11133,N_10160,N_10887);
nand U11134 (N_11134,N_10634,N_10291);
nor U11135 (N_11135,N_10353,N_10709);
or U11136 (N_11136,N_10904,N_10643);
xnor U11137 (N_11137,N_10311,N_10587);
xor U11138 (N_11138,N_10662,N_10199);
and U11139 (N_11139,N_10496,N_10684);
nand U11140 (N_11140,N_10167,N_10638);
xor U11141 (N_11141,N_10631,N_10655);
nor U11142 (N_11142,N_10796,N_10343);
xnor U11143 (N_11143,N_10118,N_10136);
nand U11144 (N_11144,N_10128,N_10930);
and U11145 (N_11145,N_10405,N_10384);
nand U11146 (N_11146,N_10976,N_10446);
xor U11147 (N_11147,N_10732,N_10295);
and U11148 (N_11148,N_10689,N_10750);
nand U11149 (N_11149,N_10403,N_10314);
nand U11150 (N_11150,N_10277,N_10608);
xnor U11151 (N_11151,N_10062,N_10555);
xnor U11152 (N_11152,N_10324,N_10340);
nand U11153 (N_11153,N_10441,N_10371);
or U11154 (N_11154,N_10594,N_10216);
nor U11155 (N_11155,N_10431,N_10258);
and U11156 (N_11156,N_10806,N_10627);
and U11157 (N_11157,N_10415,N_10075);
xor U11158 (N_11158,N_10491,N_10679);
xnor U11159 (N_11159,N_10764,N_10729);
nor U11160 (N_11160,N_10121,N_10414);
nand U11161 (N_11161,N_10603,N_10646);
nor U11162 (N_11162,N_10043,N_10741);
nand U11163 (N_11163,N_10106,N_10483);
or U11164 (N_11164,N_10411,N_10748);
nand U11165 (N_11165,N_10955,N_10862);
and U11166 (N_11166,N_10178,N_10669);
nor U11167 (N_11167,N_10244,N_10180);
xnor U11168 (N_11168,N_10196,N_10443);
nand U11169 (N_11169,N_10616,N_10702);
nor U11170 (N_11170,N_10263,N_10936);
or U11171 (N_11171,N_10218,N_10298);
xor U11172 (N_11172,N_10678,N_10580);
nand U11173 (N_11173,N_10845,N_10189);
xor U11174 (N_11174,N_10381,N_10737);
and U11175 (N_11175,N_10081,N_10610);
nand U11176 (N_11176,N_10428,N_10657);
and U11177 (N_11177,N_10949,N_10572);
nor U11178 (N_11178,N_10356,N_10132);
nor U11179 (N_11179,N_10883,N_10531);
nand U11180 (N_11180,N_10534,N_10025);
or U11181 (N_11181,N_10396,N_10060);
and U11182 (N_11182,N_10186,N_10107);
xor U11183 (N_11183,N_10874,N_10567);
nor U11184 (N_11184,N_10322,N_10184);
or U11185 (N_11185,N_10198,N_10675);
nor U11186 (N_11186,N_10753,N_10820);
and U11187 (N_11187,N_10170,N_10870);
nor U11188 (N_11188,N_10970,N_10379);
or U11189 (N_11189,N_10681,N_10018);
nor U11190 (N_11190,N_10588,N_10865);
or U11191 (N_11191,N_10987,N_10212);
nand U11192 (N_11192,N_10973,N_10727);
nor U11193 (N_11193,N_10692,N_10385);
nor U11194 (N_11194,N_10775,N_10240);
xor U11195 (N_11195,N_10794,N_10816);
nor U11196 (N_11196,N_10548,N_10476);
and U11197 (N_11197,N_10589,N_10541);
nand U11198 (N_11198,N_10501,N_10597);
nor U11199 (N_11199,N_10687,N_10562);
xor U11200 (N_11200,N_10744,N_10720);
nand U11201 (N_11201,N_10635,N_10477);
or U11202 (N_11202,N_10535,N_10427);
nand U11203 (N_11203,N_10021,N_10546);
or U11204 (N_11204,N_10071,N_10873);
nor U11205 (N_11205,N_10429,N_10253);
or U11206 (N_11206,N_10529,N_10089);
xnor U11207 (N_11207,N_10256,N_10911);
nand U11208 (N_11208,N_10857,N_10774);
nor U11209 (N_11209,N_10785,N_10351);
or U11210 (N_11210,N_10394,N_10872);
nand U11211 (N_11211,N_10090,N_10522);
nand U11212 (N_11212,N_10761,N_10234);
xnor U11213 (N_11213,N_10972,N_10448);
or U11214 (N_11214,N_10584,N_10074);
or U11215 (N_11215,N_10119,N_10318);
and U11216 (N_11216,N_10440,N_10953);
and U11217 (N_11217,N_10304,N_10888);
nand U11218 (N_11218,N_10282,N_10893);
or U11219 (N_11219,N_10344,N_10786);
nor U11220 (N_11220,N_10172,N_10983);
or U11221 (N_11221,N_10502,N_10085);
nor U11222 (N_11222,N_10487,N_10512);
xnor U11223 (N_11223,N_10366,N_10361);
xor U11224 (N_11224,N_10791,N_10839);
nor U11225 (N_11225,N_10975,N_10962);
nand U11226 (N_11226,N_10864,N_10185);
or U11227 (N_11227,N_10015,N_10947);
and U11228 (N_11228,N_10768,N_10393);
nor U11229 (N_11229,N_10795,N_10434);
xor U11230 (N_11230,N_10425,N_10614);
nor U11231 (N_11231,N_10449,N_10842);
nand U11232 (N_11232,N_10700,N_10777);
nor U11233 (N_11233,N_10543,N_10685);
and U11234 (N_11234,N_10310,N_10878);
or U11235 (N_11235,N_10139,N_10508);
nor U11236 (N_11236,N_10355,N_10843);
nand U11237 (N_11237,N_10171,N_10942);
xnor U11238 (N_11238,N_10037,N_10641);
xor U11239 (N_11239,N_10130,N_10468);
and U11240 (N_11240,N_10463,N_10034);
nand U11241 (N_11241,N_10505,N_10289);
nand U11242 (N_11242,N_10313,N_10981);
xor U11243 (N_11243,N_10565,N_10057);
or U11244 (N_11244,N_10161,N_10633);
nor U11245 (N_11245,N_10688,N_10549);
nor U11246 (N_11246,N_10150,N_10841);
xor U11247 (N_11247,N_10855,N_10607);
xor U11248 (N_11248,N_10370,N_10397);
and U11249 (N_11249,N_10469,N_10472);
nor U11250 (N_11250,N_10204,N_10112);
and U11251 (N_11251,N_10177,N_10471);
xor U11252 (N_11252,N_10758,N_10173);
xnor U11253 (N_11253,N_10359,N_10339);
nand U11254 (N_11254,N_10251,N_10084);
or U11255 (N_11255,N_10303,N_10482);
nand U11256 (N_11256,N_10649,N_10760);
or U11257 (N_11257,N_10238,N_10479);
and U11258 (N_11258,N_10210,N_10601);
xnor U11259 (N_11259,N_10152,N_10544);
xnor U11260 (N_11260,N_10988,N_10302);
and U11261 (N_11261,N_10599,N_10336);
nand U11262 (N_11262,N_10717,N_10533);
or U11263 (N_11263,N_10847,N_10763);
and U11264 (N_11264,N_10558,N_10402);
and U11265 (N_11265,N_10853,N_10069);
or U11266 (N_11266,N_10600,N_10708);
nor U11267 (N_11267,N_10099,N_10714);
nor U11268 (N_11268,N_10693,N_10746);
xnor U11269 (N_11269,N_10880,N_10255);
and U11270 (N_11270,N_10628,N_10466);
and U11271 (N_11271,N_10879,N_10367);
nand U11272 (N_11272,N_10735,N_10731);
or U11273 (N_11273,N_10765,N_10348);
and U11274 (N_11274,N_10590,N_10239);
nor U11275 (N_11275,N_10478,N_10444);
nor U11276 (N_11276,N_10530,N_10755);
or U11277 (N_11277,N_10113,N_10009);
and U11278 (N_11278,N_10995,N_10123);
nor U11279 (N_11279,N_10824,N_10586);
nand U11280 (N_11280,N_10409,N_10784);
nand U11281 (N_11281,N_10104,N_10321);
xnor U11282 (N_11282,N_10473,N_10856);
nand U11283 (N_11283,N_10985,N_10053);
xor U11284 (N_11284,N_10442,N_10330);
or U11285 (N_11285,N_10509,N_10951);
or U11286 (N_11286,N_10200,N_10867);
xor U11287 (N_11287,N_10475,N_10800);
or U11288 (N_11288,N_10000,N_10267);
nand U11289 (N_11289,N_10241,N_10165);
and U11290 (N_11290,N_10650,N_10849);
and U11291 (N_11291,N_10789,N_10871);
and U11292 (N_11292,N_10109,N_10776);
xor U11293 (N_11293,N_10602,N_10526);
and U11294 (N_11294,N_10563,N_10268);
and U11295 (N_11295,N_10153,N_10835);
nor U11296 (N_11296,N_10591,N_10902);
and U11297 (N_11297,N_10300,N_10252);
and U11298 (N_11298,N_10538,N_10604);
nand U11299 (N_11299,N_10484,N_10260);
nand U11300 (N_11300,N_10063,N_10788);
nor U11301 (N_11301,N_10206,N_10248);
nor U11302 (N_11302,N_10006,N_10208);
xnor U11303 (N_11303,N_10154,N_10108);
nand U11304 (N_11304,N_10061,N_10307);
nand U11305 (N_11305,N_10539,N_10832);
nor U11306 (N_11306,N_10220,N_10890);
nand U11307 (N_11307,N_10299,N_10305);
nor U11308 (N_11308,N_10418,N_10637);
nor U11309 (N_11309,N_10489,N_10520);
nand U11310 (N_11310,N_10400,N_10560);
and U11311 (N_11311,N_10464,N_10876);
xor U11312 (N_11312,N_10067,N_10101);
nor U11313 (N_11313,N_10219,N_10457);
nor U11314 (N_11314,N_10909,N_10460);
or U11315 (N_11315,N_10138,N_10192);
or U11316 (N_11316,N_10492,N_10131);
nor U11317 (N_11317,N_10044,N_10122);
xnor U11318 (N_11318,N_10197,N_10666);
xnor U11319 (N_11319,N_10742,N_10680);
xor U11320 (N_11320,N_10140,N_10903);
and U11321 (N_11321,N_10542,N_10885);
nand U11322 (N_11322,N_10671,N_10380);
nor U11323 (N_11323,N_10149,N_10629);
or U11324 (N_11324,N_10245,N_10706);
or U11325 (N_11325,N_10928,N_10038);
nor U11326 (N_11326,N_10850,N_10098);
nor U11327 (N_11327,N_10550,N_10485);
nand U11328 (N_11328,N_10617,N_10179);
and U11329 (N_11329,N_10771,N_10135);
or U11330 (N_11330,N_10497,N_10672);
or U11331 (N_11331,N_10554,N_10481);
nand U11332 (N_11332,N_10439,N_10126);
or U11333 (N_11333,N_10417,N_10187);
nand U11334 (N_11334,N_10333,N_10054);
nor U11335 (N_11335,N_10259,N_10914);
xnor U11336 (N_11336,N_10721,N_10690);
and U11337 (N_11337,N_10019,N_10188);
xor U11338 (N_11338,N_10016,N_10004);
and U11339 (N_11339,N_10808,N_10779);
nor U11340 (N_11340,N_10726,N_10183);
nand U11341 (N_11341,N_10323,N_10499);
and U11342 (N_11342,N_10056,N_10042);
xnor U11343 (N_11343,N_10919,N_10944);
xor U11344 (N_11344,N_10273,N_10994);
and U11345 (N_11345,N_10931,N_10227);
or U11346 (N_11346,N_10642,N_10373);
or U11347 (N_11347,N_10990,N_10694);
xor U11348 (N_11348,N_10105,N_10017);
and U11349 (N_11349,N_10474,N_10458);
and U11350 (N_11350,N_10697,N_10781);
and U11351 (N_11351,N_10719,N_10193);
and U11352 (N_11352,N_10243,N_10102);
nand U11353 (N_11353,N_10809,N_10814);
xnor U11354 (N_11354,N_10971,N_10907);
xor U11355 (N_11355,N_10826,N_10701);
or U11356 (N_11356,N_10577,N_10621);
nor U11357 (N_11357,N_10556,N_10349);
or U11358 (N_11358,N_10639,N_10581);
xor U11359 (N_11359,N_10040,N_10390);
nand U11360 (N_11360,N_10513,N_10961);
and U11361 (N_11361,N_10982,N_10134);
xor U11362 (N_11362,N_10264,N_10286);
and U11363 (N_11363,N_10686,N_10969);
or U11364 (N_11364,N_10312,N_10410);
and U11365 (N_11365,N_10271,N_10269);
nor U11366 (N_11366,N_10058,N_10596);
nand U11367 (N_11367,N_10203,N_10939);
nor U11368 (N_11368,N_10051,N_10358);
xnor U11369 (N_11369,N_10540,N_10147);
nor U11370 (N_11370,N_10986,N_10593);
and U11371 (N_11371,N_10877,N_10579);
and U11372 (N_11372,N_10124,N_10912);
nand U11373 (N_11373,N_10738,N_10730);
nor U11374 (N_11374,N_10925,N_10035);
or U11375 (N_11375,N_10080,N_10103);
nor U11376 (N_11376,N_10226,N_10899);
xor U11377 (N_11377,N_10413,N_10287);
xnor U11378 (N_11378,N_10651,N_10451);
and U11379 (N_11379,N_10350,N_10031);
nor U11380 (N_11380,N_10455,N_10778);
or U11381 (N_11381,N_10715,N_10325);
or U11382 (N_11382,N_10674,N_10819);
xor U11383 (N_11383,N_10979,N_10423);
nand U11384 (N_11384,N_10221,N_10963);
nor U11385 (N_11385,N_10461,N_10383);
xor U11386 (N_11386,N_10093,N_10096);
and U11387 (N_11387,N_10921,N_10846);
or U11388 (N_11388,N_10622,N_10618);
nor U11389 (N_11389,N_10036,N_10211);
or U11390 (N_11390,N_10279,N_10065);
and U11391 (N_11391,N_10070,N_10347);
or U11392 (N_11392,N_10648,N_10910);
xor U11393 (N_11393,N_10677,N_10377);
nor U11394 (N_11394,N_10863,N_10117);
xnor U11395 (N_11395,N_10158,N_10802);
nand U11396 (N_11396,N_10783,N_10866);
or U11397 (N_11397,N_10734,N_10229);
nand U11398 (N_11398,N_10576,N_10707);
xor U11399 (N_11399,N_10280,N_10725);
nand U11400 (N_11400,N_10368,N_10421);
xnor U11401 (N_11401,N_10860,N_10225);
xor U11402 (N_11402,N_10704,N_10894);
or U11403 (N_11403,N_10564,N_10488);
nand U11404 (N_11404,N_10797,N_10480);
and U11405 (N_11405,N_10228,N_10335);
and U11406 (N_11406,N_10517,N_10086);
and U11407 (N_11407,N_10833,N_10045);
nand U11408 (N_11408,N_10932,N_10059);
xor U11409 (N_11409,N_10453,N_10828);
and U11410 (N_11410,N_10523,N_10926);
xnor U11411 (N_11411,N_10331,N_10231);
nand U11412 (N_11412,N_10670,N_10023);
or U11413 (N_11413,N_10749,N_10205);
or U11414 (N_11414,N_10100,N_10598);
and U11415 (N_11415,N_10917,N_10033);
and U11416 (N_11416,N_10898,N_10011);
and U11417 (N_11417,N_10047,N_10740);
nor U11418 (N_11418,N_10830,N_10647);
nand U11419 (N_11419,N_10145,N_10164);
xor U11420 (N_11420,N_10787,N_10859);
nand U11421 (N_11421,N_10445,N_10293);
xor U11422 (N_11422,N_10407,N_10120);
nor U11423 (N_11423,N_10048,N_10773);
nor U11424 (N_11424,N_10072,N_10664);
nor U11425 (N_11425,N_10014,N_10559);
xor U11426 (N_11426,N_10055,N_10436);
xor U11427 (N_11427,N_10521,N_10984);
nor U11428 (N_11428,N_10767,N_10524);
nand U11429 (N_11429,N_10605,N_10869);
and U11430 (N_11430,N_10891,N_10831);
nor U11431 (N_11431,N_10275,N_10190);
nand U11432 (N_11432,N_10265,N_10078);
nor U11433 (N_11433,N_10195,N_10992);
or U11434 (N_11434,N_10079,N_10772);
or U11435 (N_11435,N_10110,N_10378);
and U11436 (N_11436,N_10739,N_10854);
or U11437 (N_11437,N_10752,N_10825);
nor U11438 (N_11438,N_10881,N_10852);
xor U11439 (N_11439,N_10920,N_10141);
nor U11440 (N_11440,N_10142,N_10570);
nand U11441 (N_11441,N_10319,N_10181);
or U11442 (N_11442,N_10486,N_10659);
nor U11443 (N_11443,N_10525,N_10435);
xnor U11444 (N_11444,N_10076,N_10615);
and U11445 (N_11445,N_10144,N_10571);
nand U11446 (N_11446,N_10710,N_10733);
or U11447 (N_11447,N_10399,N_10342);
nor U11448 (N_11448,N_10977,N_10456);
xor U11449 (N_11449,N_10799,N_10913);
xnor U11450 (N_11450,N_10284,N_10247);
and U11451 (N_11451,N_10811,N_10039);
xnor U11452 (N_11452,N_10372,N_10224);
nor U11453 (N_11453,N_10557,N_10470);
nand U11454 (N_11454,N_10097,N_10656);
and U11455 (N_11455,N_10823,N_10875);
or U11456 (N_11456,N_10094,N_10419);
or U11457 (N_11457,N_10916,N_10613);
or U11458 (N_11458,N_10412,N_10207);
and U11459 (N_11459,N_10027,N_10438);
xnor U11460 (N_11460,N_10940,N_10507);
nor U11461 (N_11461,N_10447,N_10682);
xor U11462 (N_11462,N_10168,N_10064);
and U11463 (N_11463,N_10129,N_10964);
nor U11464 (N_11464,N_10712,N_10908);
or U11465 (N_11465,N_10363,N_10008);
nand U11466 (N_11466,N_10049,N_10301);
nand U11467 (N_11467,N_10769,N_10915);
xor U11468 (N_11468,N_10151,N_10665);
nand U11469 (N_11469,N_10362,N_10978);
xnor U11470 (N_11470,N_10663,N_10283);
or U11471 (N_11471,N_10519,N_10518);
nand U11472 (N_11472,N_10088,N_10782);
or U11473 (N_11473,N_10503,N_10338);
nor U11474 (N_11474,N_10426,N_10133);
nor U11475 (N_11475,N_10010,N_10143);
or U11476 (N_11476,N_10395,N_10658);
or U11477 (N_11477,N_10743,N_10703);
nor U11478 (N_11478,N_10162,N_10667);
nand U11479 (N_11479,N_10933,N_10595);
and U11480 (N_11480,N_10493,N_10001);
xor U11481 (N_11481,N_10645,N_10956);
nand U11482 (N_11482,N_10398,N_10905);
and U11483 (N_11483,N_10829,N_10886);
and U11484 (N_11484,N_10654,N_10430);
or U11485 (N_11485,N_10433,N_10527);
and U11486 (N_11486,N_10175,N_10002);
or U11487 (N_11487,N_10222,N_10528);
nand U11488 (N_11488,N_10573,N_10511);
nor U11489 (N_11489,N_10566,N_10812);
xor U11490 (N_11490,N_10420,N_10938);
and U11491 (N_11491,N_10290,N_10612);
nor U11492 (N_11492,N_10569,N_10900);
or U11493 (N_11493,N_10376,N_10250);
nand U11494 (N_11494,N_10041,N_10432);
and U11495 (N_11495,N_10997,N_10858);
and U11496 (N_11496,N_10532,N_10901);
nand U11497 (N_11497,N_10960,N_10798);
and U11498 (N_11498,N_10274,N_10922);
nand U11499 (N_11499,N_10317,N_10073);
or U11500 (N_11500,N_10752,N_10485);
and U11501 (N_11501,N_10416,N_10814);
nand U11502 (N_11502,N_10783,N_10862);
xnor U11503 (N_11503,N_10094,N_10775);
xor U11504 (N_11504,N_10067,N_10990);
nor U11505 (N_11505,N_10955,N_10046);
or U11506 (N_11506,N_10848,N_10789);
and U11507 (N_11507,N_10402,N_10076);
xnor U11508 (N_11508,N_10631,N_10296);
nor U11509 (N_11509,N_10671,N_10352);
or U11510 (N_11510,N_10730,N_10468);
nor U11511 (N_11511,N_10377,N_10913);
nand U11512 (N_11512,N_10986,N_10867);
nand U11513 (N_11513,N_10024,N_10036);
nand U11514 (N_11514,N_10695,N_10581);
and U11515 (N_11515,N_10918,N_10741);
or U11516 (N_11516,N_10621,N_10021);
or U11517 (N_11517,N_10166,N_10231);
nand U11518 (N_11518,N_10729,N_10963);
and U11519 (N_11519,N_10363,N_10072);
xnor U11520 (N_11520,N_10257,N_10856);
or U11521 (N_11521,N_10021,N_10562);
or U11522 (N_11522,N_10153,N_10543);
and U11523 (N_11523,N_10372,N_10958);
nand U11524 (N_11524,N_10186,N_10612);
nor U11525 (N_11525,N_10008,N_10150);
and U11526 (N_11526,N_10742,N_10265);
or U11527 (N_11527,N_10517,N_10944);
nand U11528 (N_11528,N_10521,N_10952);
xnor U11529 (N_11529,N_10043,N_10160);
or U11530 (N_11530,N_10549,N_10230);
nor U11531 (N_11531,N_10337,N_10854);
or U11532 (N_11532,N_10583,N_10993);
or U11533 (N_11533,N_10158,N_10834);
nand U11534 (N_11534,N_10815,N_10009);
and U11535 (N_11535,N_10965,N_10784);
or U11536 (N_11536,N_10943,N_10208);
xnor U11537 (N_11537,N_10870,N_10458);
xnor U11538 (N_11538,N_10029,N_10163);
nor U11539 (N_11539,N_10427,N_10875);
nand U11540 (N_11540,N_10229,N_10721);
and U11541 (N_11541,N_10654,N_10167);
nand U11542 (N_11542,N_10074,N_10357);
and U11543 (N_11543,N_10524,N_10124);
nand U11544 (N_11544,N_10192,N_10804);
xor U11545 (N_11545,N_10620,N_10003);
and U11546 (N_11546,N_10650,N_10792);
or U11547 (N_11547,N_10918,N_10414);
nand U11548 (N_11548,N_10911,N_10604);
nand U11549 (N_11549,N_10061,N_10496);
or U11550 (N_11550,N_10977,N_10179);
and U11551 (N_11551,N_10386,N_10298);
and U11552 (N_11552,N_10288,N_10136);
or U11553 (N_11553,N_10449,N_10964);
and U11554 (N_11554,N_10220,N_10521);
nand U11555 (N_11555,N_10085,N_10949);
nor U11556 (N_11556,N_10805,N_10420);
nor U11557 (N_11557,N_10399,N_10953);
nor U11558 (N_11558,N_10318,N_10047);
xor U11559 (N_11559,N_10589,N_10742);
xnor U11560 (N_11560,N_10067,N_10898);
nand U11561 (N_11561,N_10230,N_10167);
or U11562 (N_11562,N_10758,N_10076);
nor U11563 (N_11563,N_10033,N_10790);
or U11564 (N_11564,N_10920,N_10973);
nor U11565 (N_11565,N_10310,N_10236);
or U11566 (N_11566,N_10216,N_10551);
or U11567 (N_11567,N_10773,N_10731);
xor U11568 (N_11568,N_10577,N_10287);
nor U11569 (N_11569,N_10794,N_10365);
and U11570 (N_11570,N_10010,N_10135);
and U11571 (N_11571,N_10699,N_10311);
nand U11572 (N_11572,N_10608,N_10749);
or U11573 (N_11573,N_10837,N_10146);
and U11574 (N_11574,N_10399,N_10922);
nand U11575 (N_11575,N_10578,N_10585);
nand U11576 (N_11576,N_10745,N_10947);
or U11577 (N_11577,N_10877,N_10554);
nand U11578 (N_11578,N_10929,N_10570);
xor U11579 (N_11579,N_10157,N_10234);
xnor U11580 (N_11580,N_10390,N_10148);
or U11581 (N_11581,N_10478,N_10090);
nand U11582 (N_11582,N_10545,N_10764);
and U11583 (N_11583,N_10274,N_10372);
nand U11584 (N_11584,N_10730,N_10479);
nand U11585 (N_11585,N_10359,N_10304);
nand U11586 (N_11586,N_10410,N_10192);
and U11587 (N_11587,N_10197,N_10192);
xnor U11588 (N_11588,N_10755,N_10260);
and U11589 (N_11589,N_10855,N_10938);
or U11590 (N_11590,N_10433,N_10652);
xnor U11591 (N_11591,N_10516,N_10619);
or U11592 (N_11592,N_10661,N_10524);
xor U11593 (N_11593,N_10192,N_10464);
xor U11594 (N_11594,N_10580,N_10152);
nand U11595 (N_11595,N_10014,N_10752);
xnor U11596 (N_11596,N_10713,N_10965);
xor U11597 (N_11597,N_10228,N_10286);
nor U11598 (N_11598,N_10118,N_10423);
and U11599 (N_11599,N_10707,N_10639);
or U11600 (N_11600,N_10378,N_10516);
nand U11601 (N_11601,N_10006,N_10858);
nor U11602 (N_11602,N_10250,N_10156);
and U11603 (N_11603,N_10334,N_10557);
nand U11604 (N_11604,N_10828,N_10700);
nand U11605 (N_11605,N_10126,N_10521);
nor U11606 (N_11606,N_10570,N_10835);
and U11607 (N_11607,N_10053,N_10391);
nand U11608 (N_11608,N_10738,N_10352);
or U11609 (N_11609,N_10874,N_10018);
nor U11610 (N_11610,N_10517,N_10315);
nand U11611 (N_11611,N_10346,N_10169);
xnor U11612 (N_11612,N_10380,N_10458);
and U11613 (N_11613,N_10407,N_10459);
xor U11614 (N_11614,N_10901,N_10132);
and U11615 (N_11615,N_10856,N_10977);
and U11616 (N_11616,N_10254,N_10795);
nor U11617 (N_11617,N_10949,N_10316);
xnor U11618 (N_11618,N_10980,N_10439);
xor U11619 (N_11619,N_10646,N_10889);
xor U11620 (N_11620,N_10763,N_10406);
nand U11621 (N_11621,N_10413,N_10082);
nor U11622 (N_11622,N_10549,N_10786);
xor U11623 (N_11623,N_10933,N_10322);
xnor U11624 (N_11624,N_10669,N_10150);
or U11625 (N_11625,N_10128,N_10145);
and U11626 (N_11626,N_10534,N_10594);
xor U11627 (N_11627,N_10519,N_10343);
nand U11628 (N_11628,N_10492,N_10776);
nor U11629 (N_11629,N_10156,N_10545);
nand U11630 (N_11630,N_10913,N_10409);
xnor U11631 (N_11631,N_10330,N_10046);
xor U11632 (N_11632,N_10927,N_10300);
and U11633 (N_11633,N_10404,N_10973);
xor U11634 (N_11634,N_10023,N_10283);
and U11635 (N_11635,N_10646,N_10521);
xnor U11636 (N_11636,N_10723,N_10893);
nor U11637 (N_11637,N_10905,N_10782);
nor U11638 (N_11638,N_10485,N_10016);
nand U11639 (N_11639,N_10155,N_10515);
or U11640 (N_11640,N_10070,N_10172);
or U11641 (N_11641,N_10812,N_10859);
nor U11642 (N_11642,N_10816,N_10075);
xor U11643 (N_11643,N_10360,N_10091);
or U11644 (N_11644,N_10324,N_10980);
nor U11645 (N_11645,N_10311,N_10515);
or U11646 (N_11646,N_10300,N_10143);
and U11647 (N_11647,N_10796,N_10631);
nor U11648 (N_11648,N_10853,N_10100);
or U11649 (N_11649,N_10759,N_10140);
or U11650 (N_11650,N_10509,N_10658);
xor U11651 (N_11651,N_10993,N_10983);
and U11652 (N_11652,N_10485,N_10930);
xnor U11653 (N_11653,N_10424,N_10592);
nand U11654 (N_11654,N_10355,N_10992);
nand U11655 (N_11655,N_10046,N_10005);
nand U11656 (N_11656,N_10052,N_10013);
and U11657 (N_11657,N_10968,N_10260);
nand U11658 (N_11658,N_10993,N_10487);
and U11659 (N_11659,N_10122,N_10843);
and U11660 (N_11660,N_10795,N_10998);
nand U11661 (N_11661,N_10861,N_10243);
nor U11662 (N_11662,N_10640,N_10288);
xor U11663 (N_11663,N_10416,N_10689);
nand U11664 (N_11664,N_10838,N_10406);
or U11665 (N_11665,N_10363,N_10168);
nand U11666 (N_11666,N_10022,N_10722);
and U11667 (N_11667,N_10439,N_10451);
nor U11668 (N_11668,N_10212,N_10911);
and U11669 (N_11669,N_10586,N_10344);
or U11670 (N_11670,N_10830,N_10270);
or U11671 (N_11671,N_10759,N_10305);
xor U11672 (N_11672,N_10289,N_10793);
nand U11673 (N_11673,N_10693,N_10402);
and U11674 (N_11674,N_10026,N_10022);
or U11675 (N_11675,N_10964,N_10655);
xor U11676 (N_11676,N_10079,N_10081);
nand U11677 (N_11677,N_10480,N_10485);
nor U11678 (N_11678,N_10880,N_10450);
or U11679 (N_11679,N_10587,N_10146);
nor U11680 (N_11680,N_10081,N_10618);
nor U11681 (N_11681,N_10157,N_10865);
nor U11682 (N_11682,N_10492,N_10496);
and U11683 (N_11683,N_10222,N_10751);
nand U11684 (N_11684,N_10342,N_10073);
nor U11685 (N_11685,N_10516,N_10033);
or U11686 (N_11686,N_10994,N_10648);
nand U11687 (N_11687,N_10138,N_10240);
or U11688 (N_11688,N_10496,N_10780);
and U11689 (N_11689,N_10212,N_10139);
nand U11690 (N_11690,N_10875,N_10463);
nand U11691 (N_11691,N_10109,N_10388);
nand U11692 (N_11692,N_10382,N_10136);
xor U11693 (N_11693,N_10361,N_10391);
and U11694 (N_11694,N_10274,N_10496);
and U11695 (N_11695,N_10174,N_10518);
nand U11696 (N_11696,N_10492,N_10886);
and U11697 (N_11697,N_10346,N_10210);
nand U11698 (N_11698,N_10556,N_10531);
or U11699 (N_11699,N_10723,N_10128);
nand U11700 (N_11700,N_10188,N_10299);
and U11701 (N_11701,N_10519,N_10185);
or U11702 (N_11702,N_10690,N_10850);
nor U11703 (N_11703,N_10021,N_10436);
and U11704 (N_11704,N_10952,N_10492);
and U11705 (N_11705,N_10650,N_10451);
xnor U11706 (N_11706,N_10728,N_10199);
xnor U11707 (N_11707,N_10557,N_10343);
or U11708 (N_11708,N_10672,N_10988);
or U11709 (N_11709,N_10380,N_10513);
and U11710 (N_11710,N_10348,N_10309);
nand U11711 (N_11711,N_10210,N_10563);
xor U11712 (N_11712,N_10218,N_10695);
and U11713 (N_11713,N_10846,N_10694);
xor U11714 (N_11714,N_10473,N_10961);
nand U11715 (N_11715,N_10454,N_10591);
or U11716 (N_11716,N_10582,N_10111);
nand U11717 (N_11717,N_10197,N_10342);
xor U11718 (N_11718,N_10567,N_10066);
nand U11719 (N_11719,N_10211,N_10464);
xnor U11720 (N_11720,N_10209,N_10186);
xnor U11721 (N_11721,N_10512,N_10828);
or U11722 (N_11722,N_10056,N_10886);
nand U11723 (N_11723,N_10787,N_10252);
or U11724 (N_11724,N_10036,N_10146);
xnor U11725 (N_11725,N_10138,N_10353);
or U11726 (N_11726,N_10603,N_10983);
and U11727 (N_11727,N_10917,N_10982);
and U11728 (N_11728,N_10534,N_10954);
nand U11729 (N_11729,N_10446,N_10497);
xor U11730 (N_11730,N_10607,N_10799);
or U11731 (N_11731,N_10242,N_10114);
nor U11732 (N_11732,N_10678,N_10141);
nand U11733 (N_11733,N_10416,N_10382);
xor U11734 (N_11734,N_10101,N_10103);
and U11735 (N_11735,N_10578,N_10149);
and U11736 (N_11736,N_10195,N_10166);
xnor U11737 (N_11737,N_10792,N_10003);
xnor U11738 (N_11738,N_10537,N_10560);
or U11739 (N_11739,N_10364,N_10331);
and U11740 (N_11740,N_10952,N_10804);
or U11741 (N_11741,N_10230,N_10363);
and U11742 (N_11742,N_10948,N_10098);
nand U11743 (N_11743,N_10889,N_10450);
or U11744 (N_11744,N_10986,N_10983);
or U11745 (N_11745,N_10941,N_10207);
nand U11746 (N_11746,N_10624,N_10408);
nand U11747 (N_11747,N_10252,N_10211);
nor U11748 (N_11748,N_10424,N_10738);
or U11749 (N_11749,N_10015,N_10833);
and U11750 (N_11750,N_10124,N_10778);
nor U11751 (N_11751,N_10175,N_10852);
nand U11752 (N_11752,N_10091,N_10571);
or U11753 (N_11753,N_10044,N_10527);
nor U11754 (N_11754,N_10019,N_10250);
nand U11755 (N_11755,N_10705,N_10857);
nor U11756 (N_11756,N_10810,N_10560);
and U11757 (N_11757,N_10546,N_10925);
nand U11758 (N_11758,N_10459,N_10340);
nand U11759 (N_11759,N_10888,N_10916);
and U11760 (N_11760,N_10834,N_10961);
xor U11761 (N_11761,N_10872,N_10287);
xor U11762 (N_11762,N_10521,N_10830);
and U11763 (N_11763,N_10996,N_10298);
xor U11764 (N_11764,N_10810,N_10903);
xor U11765 (N_11765,N_10836,N_10060);
xor U11766 (N_11766,N_10581,N_10680);
and U11767 (N_11767,N_10709,N_10403);
nor U11768 (N_11768,N_10473,N_10725);
nor U11769 (N_11769,N_10086,N_10766);
nand U11770 (N_11770,N_10127,N_10902);
xor U11771 (N_11771,N_10315,N_10138);
nor U11772 (N_11772,N_10119,N_10251);
and U11773 (N_11773,N_10949,N_10725);
nor U11774 (N_11774,N_10984,N_10554);
and U11775 (N_11775,N_10204,N_10284);
and U11776 (N_11776,N_10270,N_10343);
xor U11777 (N_11777,N_10725,N_10288);
or U11778 (N_11778,N_10070,N_10321);
or U11779 (N_11779,N_10890,N_10111);
and U11780 (N_11780,N_10090,N_10441);
nor U11781 (N_11781,N_10302,N_10719);
nor U11782 (N_11782,N_10665,N_10380);
or U11783 (N_11783,N_10035,N_10881);
and U11784 (N_11784,N_10056,N_10870);
xor U11785 (N_11785,N_10857,N_10081);
xor U11786 (N_11786,N_10290,N_10336);
xnor U11787 (N_11787,N_10795,N_10516);
xor U11788 (N_11788,N_10290,N_10042);
nand U11789 (N_11789,N_10824,N_10872);
xnor U11790 (N_11790,N_10499,N_10431);
nor U11791 (N_11791,N_10695,N_10897);
nand U11792 (N_11792,N_10950,N_10722);
nor U11793 (N_11793,N_10421,N_10931);
nand U11794 (N_11794,N_10995,N_10632);
nand U11795 (N_11795,N_10182,N_10331);
nand U11796 (N_11796,N_10903,N_10044);
xor U11797 (N_11797,N_10048,N_10497);
nand U11798 (N_11798,N_10855,N_10650);
nor U11799 (N_11799,N_10726,N_10262);
nor U11800 (N_11800,N_10330,N_10048);
xor U11801 (N_11801,N_10725,N_10412);
or U11802 (N_11802,N_10588,N_10260);
xnor U11803 (N_11803,N_10227,N_10349);
nor U11804 (N_11804,N_10092,N_10309);
nor U11805 (N_11805,N_10048,N_10401);
and U11806 (N_11806,N_10936,N_10626);
nand U11807 (N_11807,N_10858,N_10927);
xnor U11808 (N_11808,N_10362,N_10248);
and U11809 (N_11809,N_10865,N_10333);
nor U11810 (N_11810,N_10508,N_10894);
or U11811 (N_11811,N_10959,N_10936);
nand U11812 (N_11812,N_10643,N_10592);
nand U11813 (N_11813,N_10060,N_10922);
nor U11814 (N_11814,N_10184,N_10042);
and U11815 (N_11815,N_10466,N_10658);
or U11816 (N_11816,N_10233,N_10687);
and U11817 (N_11817,N_10643,N_10465);
nor U11818 (N_11818,N_10911,N_10602);
nand U11819 (N_11819,N_10917,N_10469);
and U11820 (N_11820,N_10443,N_10428);
nand U11821 (N_11821,N_10625,N_10187);
and U11822 (N_11822,N_10633,N_10764);
nand U11823 (N_11823,N_10736,N_10456);
nor U11824 (N_11824,N_10399,N_10388);
and U11825 (N_11825,N_10436,N_10758);
nand U11826 (N_11826,N_10968,N_10216);
or U11827 (N_11827,N_10798,N_10929);
nand U11828 (N_11828,N_10501,N_10912);
or U11829 (N_11829,N_10025,N_10133);
nor U11830 (N_11830,N_10980,N_10959);
xnor U11831 (N_11831,N_10626,N_10928);
nand U11832 (N_11832,N_10881,N_10651);
nand U11833 (N_11833,N_10975,N_10515);
xnor U11834 (N_11834,N_10465,N_10949);
nand U11835 (N_11835,N_10971,N_10161);
or U11836 (N_11836,N_10614,N_10077);
and U11837 (N_11837,N_10383,N_10869);
xnor U11838 (N_11838,N_10957,N_10062);
and U11839 (N_11839,N_10398,N_10729);
xnor U11840 (N_11840,N_10962,N_10404);
nor U11841 (N_11841,N_10784,N_10561);
xor U11842 (N_11842,N_10605,N_10079);
nand U11843 (N_11843,N_10927,N_10424);
nand U11844 (N_11844,N_10552,N_10353);
or U11845 (N_11845,N_10664,N_10085);
xor U11846 (N_11846,N_10223,N_10195);
xor U11847 (N_11847,N_10522,N_10385);
or U11848 (N_11848,N_10923,N_10306);
xor U11849 (N_11849,N_10095,N_10275);
xor U11850 (N_11850,N_10796,N_10339);
and U11851 (N_11851,N_10212,N_10082);
xnor U11852 (N_11852,N_10583,N_10457);
nand U11853 (N_11853,N_10461,N_10722);
nor U11854 (N_11854,N_10208,N_10385);
or U11855 (N_11855,N_10910,N_10215);
nand U11856 (N_11856,N_10384,N_10507);
or U11857 (N_11857,N_10484,N_10154);
or U11858 (N_11858,N_10450,N_10133);
nand U11859 (N_11859,N_10811,N_10873);
or U11860 (N_11860,N_10930,N_10655);
nor U11861 (N_11861,N_10772,N_10340);
and U11862 (N_11862,N_10464,N_10454);
xor U11863 (N_11863,N_10422,N_10492);
nand U11864 (N_11864,N_10971,N_10369);
and U11865 (N_11865,N_10373,N_10412);
xor U11866 (N_11866,N_10503,N_10441);
xor U11867 (N_11867,N_10811,N_10520);
and U11868 (N_11868,N_10981,N_10161);
nor U11869 (N_11869,N_10203,N_10114);
or U11870 (N_11870,N_10072,N_10701);
or U11871 (N_11871,N_10181,N_10231);
and U11872 (N_11872,N_10589,N_10637);
xor U11873 (N_11873,N_10910,N_10567);
nor U11874 (N_11874,N_10616,N_10555);
or U11875 (N_11875,N_10796,N_10731);
nand U11876 (N_11876,N_10263,N_10075);
xor U11877 (N_11877,N_10199,N_10097);
and U11878 (N_11878,N_10990,N_10921);
or U11879 (N_11879,N_10273,N_10415);
or U11880 (N_11880,N_10840,N_10797);
xnor U11881 (N_11881,N_10187,N_10238);
nor U11882 (N_11882,N_10886,N_10664);
nand U11883 (N_11883,N_10585,N_10995);
xnor U11884 (N_11884,N_10770,N_10847);
xor U11885 (N_11885,N_10399,N_10719);
xor U11886 (N_11886,N_10718,N_10472);
and U11887 (N_11887,N_10254,N_10834);
and U11888 (N_11888,N_10154,N_10477);
nor U11889 (N_11889,N_10400,N_10102);
or U11890 (N_11890,N_10051,N_10538);
and U11891 (N_11891,N_10047,N_10905);
nor U11892 (N_11892,N_10151,N_10993);
nand U11893 (N_11893,N_10777,N_10024);
nand U11894 (N_11894,N_10827,N_10993);
nand U11895 (N_11895,N_10892,N_10328);
nand U11896 (N_11896,N_10011,N_10194);
and U11897 (N_11897,N_10702,N_10293);
or U11898 (N_11898,N_10880,N_10252);
nor U11899 (N_11899,N_10059,N_10915);
or U11900 (N_11900,N_10140,N_10975);
and U11901 (N_11901,N_10543,N_10529);
xnor U11902 (N_11902,N_10015,N_10376);
xnor U11903 (N_11903,N_10692,N_10334);
nor U11904 (N_11904,N_10538,N_10400);
xnor U11905 (N_11905,N_10383,N_10036);
xnor U11906 (N_11906,N_10911,N_10580);
and U11907 (N_11907,N_10294,N_10455);
xnor U11908 (N_11908,N_10334,N_10165);
and U11909 (N_11909,N_10980,N_10706);
and U11910 (N_11910,N_10569,N_10407);
or U11911 (N_11911,N_10226,N_10123);
nor U11912 (N_11912,N_10679,N_10931);
and U11913 (N_11913,N_10256,N_10999);
or U11914 (N_11914,N_10990,N_10855);
nand U11915 (N_11915,N_10250,N_10514);
and U11916 (N_11916,N_10199,N_10391);
xor U11917 (N_11917,N_10284,N_10184);
and U11918 (N_11918,N_10669,N_10208);
or U11919 (N_11919,N_10968,N_10263);
or U11920 (N_11920,N_10627,N_10247);
nor U11921 (N_11921,N_10674,N_10882);
nor U11922 (N_11922,N_10421,N_10831);
and U11923 (N_11923,N_10729,N_10296);
xnor U11924 (N_11924,N_10721,N_10265);
xnor U11925 (N_11925,N_10472,N_10633);
and U11926 (N_11926,N_10996,N_10331);
xor U11927 (N_11927,N_10956,N_10757);
or U11928 (N_11928,N_10603,N_10204);
xnor U11929 (N_11929,N_10814,N_10211);
nor U11930 (N_11930,N_10618,N_10315);
and U11931 (N_11931,N_10903,N_10461);
and U11932 (N_11932,N_10375,N_10033);
or U11933 (N_11933,N_10247,N_10116);
nor U11934 (N_11934,N_10141,N_10336);
and U11935 (N_11935,N_10063,N_10950);
xnor U11936 (N_11936,N_10138,N_10556);
nor U11937 (N_11937,N_10622,N_10578);
or U11938 (N_11938,N_10491,N_10889);
or U11939 (N_11939,N_10049,N_10137);
nand U11940 (N_11940,N_10795,N_10984);
and U11941 (N_11941,N_10677,N_10536);
and U11942 (N_11942,N_10836,N_10092);
xor U11943 (N_11943,N_10771,N_10685);
nor U11944 (N_11944,N_10317,N_10417);
and U11945 (N_11945,N_10174,N_10998);
xor U11946 (N_11946,N_10495,N_10028);
or U11947 (N_11947,N_10071,N_10914);
xor U11948 (N_11948,N_10252,N_10640);
and U11949 (N_11949,N_10922,N_10357);
nor U11950 (N_11950,N_10612,N_10868);
and U11951 (N_11951,N_10170,N_10399);
nand U11952 (N_11952,N_10621,N_10136);
and U11953 (N_11953,N_10932,N_10227);
and U11954 (N_11954,N_10926,N_10991);
nand U11955 (N_11955,N_10698,N_10278);
or U11956 (N_11956,N_10232,N_10535);
or U11957 (N_11957,N_10499,N_10163);
xnor U11958 (N_11958,N_10793,N_10656);
and U11959 (N_11959,N_10020,N_10346);
xor U11960 (N_11960,N_10900,N_10744);
or U11961 (N_11961,N_10979,N_10066);
or U11962 (N_11962,N_10487,N_10502);
or U11963 (N_11963,N_10473,N_10847);
xor U11964 (N_11964,N_10896,N_10413);
and U11965 (N_11965,N_10136,N_10534);
or U11966 (N_11966,N_10471,N_10373);
nor U11967 (N_11967,N_10441,N_10027);
or U11968 (N_11968,N_10192,N_10630);
xnor U11969 (N_11969,N_10453,N_10417);
nor U11970 (N_11970,N_10826,N_10188);
nor U11971 (N_11971,N_10663,N_10253);
and U11972 (N_11972,N_10197,N_10624);
nand U11973 (N_11973,N_10950,N_10125);
nor U11974 (N_11974,N_10826,N_10544);
nor U11975 (N_11975,N_10474,N_10136);
or U11976 (N_11976,N_10437,N_10297);
and U11977 (N_11977,N_10844,N_10022);
nor U11978 (N_11978,N_10728,N_10850);
or U11979 (N_11979,N_10733,N_10764);
nand U11980 (N_11980,N_10674,N_10454);
nor U11981 (N_11981,N_10565,N_10413);
xor U11982 (N_11982,N_10660,N_10167);
nand U11983 (N_11983,N_10991,N_10422);
or U11984 (N_11984,N_10154,N_10400);
nor U11985 (N_11985,N_10893,N_10201);
nor U11986 (N_11986,N_10329,N_10845);
and U11987 (N_11987,N_10773,N_10148);
nor U11988 (N_11988,N_10970,N_10364);
xnor U11989 (N_11989,N_10109,N_10076);
and U11990 (N_11990,N_10523,N_10356);
and U11991 (N_11991,N_10480,N_10667);
xor U11992 (N_11992,N_10593,N_10911);
nor U11993 (N_11993,N_10697,N_10593);
nand U11994 (N_11994,N_10205,N_10049);
nand U11995 (N_11995,N_10388,N_10041);
nand U11996 (N_11996,N_10500,N_10340);
xnor U11997 (N_11997,N_10786,N_10740);
and U11998 (N_11998,N_10691,N_10483);
and U11999 (N_11999,N_10964,N_10123);
nand U12000 (N_12000,N_11604,N_11884);
or U12001 (N_12001,N_11331,N_11127);
nand U12002 (N_12002,N_11566,N_11206);
nand U12003 (N_12003,N_11301,N_11834);
or U12004 (N_12004,N_11845,N_11435);
xor U12005 (N_12005,N_11973,N_11449);
and U12006 (N_12006,N_11412,N_11151);
nor U12007 (N_12007,N_11810,N_11040);
or U12008 (N_12008,N_11643,N_11669);
nor U12009 (N_12009,N_11912,N_11098);
or U12010 (N_12010,N_11764,N_11808);
and U12011 (N_12011,N_11546,N_11740);
or U12012 (N_12012,N_11996,N_11051);
xnor U12013 (N_12013,N_11796,N_11277);
xnor U12014 (N_12014,N_11362,N_11134);
or U12015 (N_12015,N_11373,N_11261);
or U12016 (N_12016,N_11711,N_11610);
nand U12017 (N_12017,N_11258,N_11313);
nand U12018 (N_12018,N_11188,N_11940);
or U12019 (N_12019,N_11284,N_11763);
nor U12020 (N_12020,N_11914,N_11426);
nand U12021 (N_12021,N_11527,N_11640);
or U12022 (N_12022,N_11798,N_11081);
and U12023 (N_12023,N_11992,N_11090);
or U12024 (N_12024,N_11406,N_11096);
xnor U12025 (N_12025,N_11153,N_11780);
xor U12026 (N_12026,N_11960,N_11541);
nor U12027 (N_12027,N_11178,N_11728);
nor U12028 (N_12028,N_11447,N_11901);
or U12029 (N_12029,N_11201,N_11918);
or U12030 (N_12030,N_11242,N_11887);
nand U12031 (N_12031,N_11743,N_11502);
nor U12032 (N_12032,N_11715,N_11524);
and U12033 (N_12033,N_11485,N_11142);
nor U12034 (N_12034,N_11194,N_11755);
and U12035 (N_12035,N_11461,N_11110);
or U12036 (N_12036,N_11994,N_11182);
nand U12037 (N_12037,N_11737,N_11727);
nand U12038 (N_12038,N_11686,N_11470);
nor U12039 (N_12039,N_11529,N_11172);
nand U12040 (N_12040,N_11868,N_11703);
and U12041 (N_12041,N_11947,N_11050);
or U12042 (N_12042,N_11220,N_11788);
xnor U12043 (N_12043,N_11468,N_11100);
nand U12044 (N_12044,N_11067,N_11121);
and U12045 (N_12045,N_11583,N_11942);
nor U12046 (N_12046,N_11817,N_11801);
xnor U12047 (N_12047,N_11783,N_11186);
and U12048 (N_12048,N_11518,N_11465);
nand U12049 (N_12049,N_11049,N_11870);
nand U12050 (N_12050,N_11593,N_11516);
xnor U12051 (N_12051,N_11733,N_11166);
xnor U12052 (N_12052,N_11818,N_11722);
nor U12053 (N_12053,N_11253,N_11423);
nor U12054 (N_12054,N_11981,N_11893);
xor U12055 (N_12055,N_11978,N_11421);
xnor U12056 (N_12056,N_11070,N_11894);
nor U12057 (N_12057,N_11547,N_11779);
xor U12058 (N_12058,N_11000,N_11397);
and U12059 (N_12059,N_11299,N_11858);
and U12060 (N_12060,N_11735,N_11768);
or U12061 (N_12061,N_11929,N_11891);
and U12062 (N_12062,N_11410,N_11056);
and U12063 (N_12063,N_11348,N_11137);
nor U12064 (N_12064,N_11745,N_11377);
nand U12065 (N_12065,N_11479,N_11445);
xor U12066 (N_12066,N_11118,N_11897);
xnor U12067 (N_12067,N_11544,N_11133);
nand U12068 (N_12068,N_11382,N_11545);
or U12069 (N_12069,N_11751,N_11682);
and U12070 (N_12070,N_11148,N_11179);
or U12071 (N_12071,N_11951,N_11287);
xnor U12072 (N_12072,N_11577,N_11268);
nand U12073 (N_12073,N_11343,N_11217);
nand U12074 (N_12074,N_11875,N_11175);
and U12075 (N_12075,N_11334,N_11214);
nor U12076 (N_12076,N_11102,N_11538);
nand U12077 (N_12077,N_11212,N_11814);
xor U12078 (N_12078,N_11670,N_11020);
nand U12079 (N_12079,N_11629,N_11741);
or U12080 (N_12080,N_11630,N_11184);
nand U12081 (N_12081,N_11187,N_11970);
and U12082 (N_12082,N_11847,N_11687);
nand U12083 (N_12083,N_11128,N_11480);
and U12084 (N_12084,N_11422,N_11309);
or U12085 (N_12085,N_11109,N_11841);
or U12086 (N_12086,N_11369,N_11559);
or U12087 (N_12087,N_11854,N_11155);
or U12088 (N_12088,N_11197,N_11667);
nor U12089 (N_12089,N_11896,N_11636);
and U12090 (N_12090,N_11407,N_11451);
nor U12091 (N_12091,N_11260,N_11785);
and U12092 (N_12092,N_11856,N_11596);
or U12093 (N_12093,N_11744,N_11395);
and U12094 (N_12094,N_11556,N_11558);
nand U12095 (N_12095,N_11292,N_11831);
or U12096 (N_12096,N_11936,N_11709);
nor U12097 (N_12097,N_11708,N_11235);
nand U12098 (N_12098,N_11554,N_11075);
or U12099 (N_12099,N_11999,N_11086);
nand U12100 (N_12100,N_11939,N_11651);
nor U12101 (N_12101,N_11296,N_11729);
nor U12102 (N_12102,N_11052,N_11104);
and U12103 (N_12103,N_11710,N_11601);
or U12104 (N_12104,N_11846,N_11227);
or U12105 (N_12105,N_11762,N_11922);
nor U12106 (N_12106,N_11913,N_11565);
nand U12107 (N_12107,N_11365,N_11748);
nand U12108 (N_12108,N_11338,N_11530);
nand U12109 (N_12109,N_11631,N_11467);
nor U12110 (N_12110,N_11816,N_11433);
nand U12111 (N_12111,N_11514,N_11493);
or U12112 (N_12112,N_11652,N_11648);
xor U12113 (N_12113,N_11797,N_11821);
nor U12114 (N_12114,N_11460,N_11419);
and U12115 (N_12115,N_11649,N_11482);
and U12116 (N_12116,N_11938,N_11865);
xnor U12117 (N_12117,N_11903,N_11676);
xnor U12118 (N_12118,N_11626,N_11813);
xnor U12119 (N_12119,N_11581,N_11697);
and U12120 (N_12120,N_11095,N_11146);
nand U12121 (N_12121,N_11700,N_11196);
nand U12122 (N_12122,N_11368,N_11572);
nor U12123 (N_12123,N_11222,N_11523);
xor U12124 (N_12124,N_11666,N_11615);
and U12125 (N_12125,N_11325,N_11066);
and U12126 (N_12126,N_11843,N_11671);
or U12127 (N_12127,N_11754,N_11414);
xor U12128 (N_12128,N_11563,N_11082);
or U12129 (N_12129,N_11275,N_11290);
nand U12130 (N_12130,N_11114,N_11394);
and U12131 (N_12131,N_11018,N_11276);
nand U12132 (N_12132,N_11580,N_11043);
and U12133 (N_12133,N_11927,N_11135);
or U12134 (N_12134,N_11370,N_11835);
and U12135 (N_12135,N_11691,N_11655);
xor U12136 (N_12136,N_11683,N_11163);
nor U12137 (N_12137,N_11047,N_11508);
nor U12138 (N_12138,N_11739,N_11665);
nand U12139 (N_12139,N_11526,N_11320);
xnor U12140 (N_12140,N_11209,N_11006);
nand U12141 (N_12141,N_11769,N_11004);
and U12142 (N_12142,N_11717,N_11827);
and U12143 (N_12143,N_11982,N_11925);
or U12144 (N_12144,N_11859,N_11656);
nor U12145 (N_12145,N_11282,N_11809);
xnor U12146 (N_12146,N_11264,N_11991);
nand U12147 (N_12147,N_11357,N_11415);
nor U12148 (N_12148,N_11466,N_11063);
nand U12149 (N_12149,N_11899,N_11356);
nor U12150 (N_12150,N_11490,N_11622);
and U12151 (N_12151,N_11753,N_11107);
xnor U12152 (N_12152,N_11007,N_11408);
nor U12153 (N_12153,N_11943,N_11010);
and U12154 (N_12154,N_11725,N_11304);
xnor U12155 (N_12155,N_11723,N_11418);
nand U12156 (N_12156,N_11624,N_11826);
or U12157 (N_12157,N_11795,N_11329);
nand U12158 (N_12158,N_11457,N_11602);
or U12159 (N_12159,N_11849,N_11488);
or U12160 (N_12160,N_11385,N_11337);
nor U12161 (N_12161,N_11034,N_11424);
xnor U12162 (N_12162,N_11861,N_11730);
or U12163 (N_12163,N_11009,N_11106);
nand U12164 (N_12164,N_11800,N_11611);
nand U12165 (N_12165,N_11384,N_11911);
nand U12166 (N_12166,N_11316,N_11409);
nor U12167 (N_12167,N_11200,N_11330);
nor U12168 (N_12168,N_11437,N_11807);
nand U12169 (N_12169,N_11044,N_11087);
xnor U12170 (N_12170,N_11573,N_11789);
and U12171 (N_12171,N_11949,N_11477);
and U12172 (N_12172,N_11885,N_11061);
or U12173 (N_12173,N_11674,N_11761);
or U12174 (N_12174,N_11877,N_11623);
and U12175 (N_12175,N_11513,N_11905);
xor U12176 (N_12176,N_11165,N_11672);
xnor U12177 (N_12177,N_11312,N_11126);
nand U12178 (N_12178,N_11873,N_11192);
nor U12179 (N_12179,N_11012,N_11819);
nand U12180 (N_12180,N_11968,N_11463);
xnor U12181 (N_12181,N_11644,N_11986);
or U12182 (N_12182,N_11079,N_11219);
or U12183 (N_12183,N_11802,N_11690);
and U12184 (N_12184,N_11678,N_11294);
or U12185 (N_12185,N_11995,N_11976);
nand U12186 (N_12186,N_11306,N_11123);
and U12187 (N_12187,N_11937,N_11120);
nand U12188 (N_12188,N_11113,N_11396);
and U12189 (N_12189,N_11767,N_11575);
nand U12190 (N_12190,N_11045,N_11383);
and U12191 (N_12191,N_11077,N_11675);
nand U12192 (N_12192,N_11928,N_11237);
xnor U12193 (N_12193,N_11042,N_11352);
or U12194 (N_12194,N_11204,N_11857);
or U12195 (N_12195,N_11791,N_11129);
xor U12196 (N_12196,N_11980,N_11517);
xnor U12197 (N_12197,N_11833,N_11907);
or U12198 (N_12198,N_11141,N_11578);
xnor U12199 (N_12199,N_11039,N_11944);
or U12200 (N_12200,N_11786,N_11895);
or U12201 (N_12201,N_11244,N_11747);
nor U12202 (N_12202,N_11698,N_11487);
nor U12203 (N_12203,N_11074,N_11612);
xnor U12204 (N_12204,N_11144,N_11974);
nand U12205 (N_12205,N_11257,N_11256);
and U12206 (N_12206,N_11898,N_11030);
xnor U12207 (N_12207,N_11302,N_11021);
nor U12208 (N_12208,N_11758,N_11668);
nand U12209 (N_12209,N_11681,N_11600);
nor U12210 (N_12210,N_11228,N_11363);
nand U12211 (N_12211,N_11387,N_11332);
xnor U12212 (N_12212,N_11948,N_11933);
or U12213 (N_12213,N_11505,N_11378);
xor U12214 (N_12214,N_11398,N_11029);
nor U12215 (N_12215,N_11945,N_11811);
nand U12216 (N_12216,N_11111,N_11489);
or U12217 (N_12217,N_11354,N_11225);
or U12218 (N_12218,N_11579,N_11055);
nand U12219 (N_12219,N_11374,N_11660);
xor U12220 (N_12220,N_11026,N_11654);
xor U12221 (N_12221,N_11318,N_11072);
nand U12222 (N_12222,N_11438,N_11536);
nand U12223 (N_12223,N_11176,N_11829);
nor U12224 (N_12224,N_11230,N_11375);
xnor U12225 (N_12225,N_11125,N_11707);
nand U12226 (N_12226,N_11956,N_11367);
nand U12227 (N_12227,N_11250,N_11420);
xor U12228 (N_12228,N_11574,N_11695);
or U12229 (N_12229,N_11543,N_11932);
nor U12230 (N_12230,N_11427,N_11019);
nand U12231 (N_12231,N_11286,N_11255);
and U12232 (N_12232,N_11634,N_11108);
or U12233 (N_12233,N_11335,N_11202);
and U12234 (N_12234,N_11360,N_11871);
or U12235 (N_12235,N_11564,N_11342);
or U12236 (N_12236,N_11168,N_11499);
xnor U12237 (N_12237,N_11492,N_11381);
nor U12238 (N_12238,N_11115,N_11850);
and U12239 (N_12239,N_11955,N_11389);
or U12240 (N_12240,N_11706,N_11853);
and U12241 (N_12241,N_11851,N_11150);
nand U12242 (N_12242,N_11439,N_11252);
xor U12243 (N_12243,N_11005,N_11453);
xnor U12244 (N_12244,N_11376,N_11411);
xnor U12245 (N_12245,N_11097,N_11825);
and U12246 (N_12246,N_11372,N_11160);
xor U12247 (N_12247,N_11716,N_11509);
nand U12248 (N_12248,N_11229,N_11249);
or U12249 (N_12249,N_11952,N_11475);
nand U12250 (N_12250,N_11860,N_11347);
nor U12251 (N_12251,N_11832,N_11481);
xnor U12252 (N_12252,N_11300,N_11507);
nand U12253 (N_12253,N_11720,N_11283);
nand U12254 (N_12254,N_11993,N_11112);
and U12255 (N_12255,N_11458,N_11156);
nor U12256 (N_12256,N_11173,N_11990);
nand U12257 (N_12257,N_11548,N_11193);
nand U12258 (N_12258,N_11588,N_11772);
nand U12259 (N_12259,N_11532,N_11361);
nor U12260 (N_12260,N_11662,N_11586);
and U12261 (N_12261,N_11533,N_11787);
xnor U12262 (N_12262,N_11595,N_11093);
xnor U12263 (N_12263,N_11659,N_11673);
nor U12264 (N_12264,N_11842,N_11921);
nor U12265 (N_12265,N_11984,N_11966);
or U12266 (N_12266,N_11303,N_11963);
and U12267 (N_12267,N_11340,N_11650);
xor U12268 (N_12268,N_11658,N_11958);
or U12269 (N_12269,N_11280,N_11476);
or U12270 (N_12270,N_11169,N_11664);
or U12271 (N_12271,N_11692,N_11719);
nor U12272 (N_12272,N_11770,N_11635);
and U12273 (N_12273,N_11326,N_11621);
nor U12274 (N_12274,N_11497,N_11035);
nor U12275 (N_12275,N_11031,N_11254);
nand U12276 (N_12276,N_11919,N_11027);
xnor U12277 (N_12277,N_11511,N_11679);
nand U12278 (N_12278,N_11525,N_11677);
nor U12279 (N_12279,N_11391,N_11613);
nor U12280 (N_12280,N_11778,N_11033);
nand U12281 (N_12281,N_11207,N_11568);
and U12282 (N_12282,N_11701,N_11210);
nor U12283 (N_12283,N_11218,N_11353);
xor U12284 (N_12284,N_11119,N_11147);
xor U12285 (N_12285,N_11443,N_11799);
and U12286 (N_12286,N_11239,N_11321);
nor U12287 (N_12287,N_11472,N_11486);
nand U12288 (N_12288,N_11346,N_11632);
nand U12289 (N_12289,N_11305,N_11646);
nor U12290 (N_12290,N_11550,N_11852);
nand U12291 (N_12291,N_11866,N_11567);
nand U12292 (N_12292,N_11089,N_11224);
or U12293 (N_12293,N_11902,N_11270);
and U12294 (N_12294,N_11024,N_11088);
nor U12295 (N_12295,N_11638,N_11483);
or U12296 (N_12296,N_11965,N_11162);
xnor U12297 (N_12297,N_11724,N_11822);
and U12298 (N_12298,N_11117,N_11085);
nor U12299 (N_12299,N_11234,N_11869);
nor U12300 (N_12300,N_11614,N_11776);
nand U12301 (N_12301,N_11388,N_11103);
xor U12302 (N_12302,N_11618,N_11551);
nor U12303 (N_12303,N_11587,N_11713);
or U12304 (N_12304,N_11130,N_11450);
nand U12305 (N_12305,N_11402,N_11404);
and U12306 (N_12306,N_11251,N_11699);
or U12307 (N_12307,N_11878,N_11247);
xnor U12308 (N_12308,N_11584,N_11881);
or U12309 (N_12309,N_11883,N_11961);
and U12310 (N_12310,N_11812,N_11528);
and U12311 (N_12311,N_11071,N_11805);
nor U12312 (N_12312,N_11653,N_11452);
nand U12313 (N_12313,N_11132,N_11607);
nor U12314 (N_12314,N_11281,N_11904);
xnor U12315 (N_12315,N_11641,N_11645);
nand U12316 (N_12316,N_11569,N_11998);
and U12317 (N_12317,N_11185,N_11983);
xnor U12318 (N_12318,N_11366,N_11782);
and U12319 (N_12319,N_11215,N_11073);
xnor U12320 (N_12320,N_11617,N_11359);
nor U12321 (N_12321,N_11985,N_11562);
nor U12322 (N_12322,N_11590,N_11417);
nor U12323 (N_12323,N_11444,N_11003);
xnor U12324 (N_12324,N_11862,N_11962);
nand U12325 (N_12325,N_11358,N_11585);
or U12326 (N_12326,N_11140,N_11693);
xor U12327 (N_12327,N_11867,N_11879);
xnor U12328 (N_12328,N_11279,N_11882);
or U12329 (N_12329,N_11262,N_11293);
nor U12330 (N_12330,N_11803,N_11272);
or U12331 (N_12331,N_11597,N_11022);
xnor U12332 (N_12332,N_11464,N_11498);
or U12333 (N_12333,N_11941,N_11839);
nor U12334 (N_12334,N_11017,N_11931);
xor U12335 (N_12335,N_11759,N_11092);
nand U12336 (N_12336,N_11392,N_11267);
and U12337 (N_12337,N_11243,N_11344);
nand U12338 (N_12338,N_11001,N_11355);
nor U12339 (N_12339,N_11263,N_11471);
nor U12340 (N_12340,N_11149,N_11350);
nor U12341 (N_12341,N_11539,N_11917);
nor U12342 (N_12342,N_11386,N_11760);
nand U12343 (N_12343,N_11553,N_11161);
nor U12344 (N_12344,N_11273,N_11552);
or U12345 (N_12345,N_11122,N_11934);
and U12346 (N_12346,N_11164,N_11425);
xnor U12347 (N_12347,N_11637,N_11351);
and U12348 (N_12348,N_11484,N_11519);
and U12349 (N_12349,N_11589,N_11742);
xnor U12350 (N_12350,N_11837,N_11848);
and U12351 (N_12351,N_11434,N_11057);
and U12352 (N_12352,N_11815,N_11393);
and U12353 (N_12353,N_11278,N_11496);
or U12354 (N_12354,N_11307,N_11766);
and U12355 (N_12355,N_11333,N_11619);
nor U12356 (N_12356,N_11756,N_11910);
xnor U12357 (N_12357,N_11512,N_11864);
and U12358 (N_12358,N_11555,N_11793);
nor U12359 (N_12359,N_11231,N_11696);
nand U12360 (N_12360,N_11198,N_11876);
and U12361 (N_12361,N_11221,N_11731);
nand U12362 (N_12362,N_11591,N_11721);
xor U12363 (N_12363,N_11345,N_11459);
nand U12364 (N_12364,N_11311,N_11454);
nand U12365 (N_12365,N_11926,N_11310);
xnor U12366 (N_12366,N_11399,N_11116);
and U12367 (N_12367,N_11967,N_11099);
nand U12368 (N_12368,N_11013,N_11792);
or U12369 (N_12369,N_11083,N_11226);
nor U12370 (N_12370,N_11874,N_11872);
or U12371 (N_12371,N_11062,N_11171);
nor U12372 (N_12372,N_11180,N_11380);
nand U12373 (N_12373,N_11238,N_11510);
nor U12374 (N_12374,N_11540,N_11094);
nand U12375 (N_12375,N_11236,N_11271);
nor U12376 (N_12376,N_11462,N_11064);
nor U12377 (N_12377,N_11964,N_11806);
nor U12378 (N_12378,N_11908,N_11339);
or U12379 (N_12379,N_11364,N_11322);
nor U12380 (N_12380,N_11515,N_11836);
and U12381 (N_12381,N_11076,N_11987);
nor U12382 (N_12382,N_11469,N_11946);
and U12383 (N_12383,N_11771,N_11432);
or U12384 (N_12384,N_11923,N_11223);
nand U12385 (N_12385,N_11011,N_11138);
or U12386 (N_12386,N_11400,N_11537);
xnor U12387 (N_12387,N_11131,N_11712);
or U12388 (N_12388,N_11975,N_11157);
and U12389 (N_12389,N_11065,N_11265);
and U12390 (N_12390,N_11718,N_11642);
and U12391 (N_12391,N_11319,N_11431);
xnor U12392 (N_12392,N_11101,N_11205);
and U12393 (N_12393,N_11336,N_11749);
nand U12394 (N_12394,N_11890,N_11246);
xor U12395 (N_12395,N_11416,N_11016);
nor U12396 (N_12396,N_11048,N_11892);
and U12397 (N_12397,N_11734,N_11576);
and U12398 (N_12398,N_11054,N_11213);
and U12399 (N_12399,N_11023,N_11765);
and U12400 (N_12400,N_11297,N_11259);
nand U12401 (N_12401,N_11080,N_11143);
nand U12402 (N_12402,N_11139,N_11920);
nand U12403 (N_12403,N_11534,N_11323);
nand U12404 (N_12404,N_11957,N_11053);
xnor U12405 (N_12405,N_11379,N_11328);
xor U12406 (N_12406,N_11840,N_11954);
xor U12407 (N_12407,N_11774,N_11609);
xor U12408 (N_12408,N_11495,N_11429);
xor U12409 (N_12409,N_11446,N_11289);
nand U12410 (N_12410,N_11561,N_11136);
and U12411 (N_12411,N_11661,N_11032);
and U12412 (N_12412,N_11582,N_11308);
nand U12413 (N_12413,N_11969,N_11189);
and U12414 (N_12414,N_11170,N_11473);
and U12415 (N_12415,N_11784,N_11828);
nor U12416 (N_12416,N_11038,N_11405);
nor U12417 (N_12417,N_11327,N_11124);
nor U12418 (N_12418,N_11503,N_11159);
xor U12419 (N_12419,N_11041,N_11091);
or U12420 (N_12420,N_11248,N_11324);
nor U12421 (N_12421,N_11199,N_11240);
nand U12422 (N_12422,N_11531,N_11491);
or U12423 (N_12423,N_11455,N_11314);
nand U12424 (N_12424,N_11522,N_11245);
and U12425 (N_12425,N_11752,N_11736);
xor U12426 (N_12426,N_11935,N_11820);
xor U12427 (N_12427,N_11838,N_11570);
xor U12428 (N_12428,N_11605,N_11977);
or U12429 (N_12429,N_11971,N_11274);
nor U12430 (N_12430,N_11233,N_11060);
nor U12431 (N_12431,N_11633,N_11500);
nand U12432 (N_12432,N_11900,N_11506);
and U12433 (N_12433,N_11906,N_11191);
xnor U12434 (N_12434,N_11542,N_11608);
xnor U12435 (N_12435,N_11824,N_11298);
xor U12436 (N_12436,N_11068,N_11183);
xnor U12437 (N_12437,N_11688,N_11989);
and U12438 (N_12438,N_11880,N_11804);
and U12439 (N_12439,N_11950,N_11037);
nand U12440 (N_12440,N_11441,N_11657);
and U12441 (N_12441,N_11501,N_11195);
xor U12442 (N_12442,N_11078,N_11105);
nor U12443 (N_12443,N_11823,N_11403);
nor U12444 (N_12444,N_11285,N_11015);
or U12445 (N_12445,N_11775,N_11606);
xor U12446 (N_12446,N_11241,N_11909);
nand U12447 (N_12447,N_11520,N_11599);
and U12448 (N_12448,N_11371,N_11535);
or U12449 (N_12449,N_11889,N_11997);
xnor U12450 (N_12450,N_11430,N_11401);
and U12451 (N_12451,N_11436,N_11478);
xor U12452 (N_12452,N_11959,N_11058);
nor U12453 (N_12453,N_11794,N_11028);
nand U12454 (N_12454,N_11266,N_11440);
nand U12455 (N_12455,N_11726,N_11177);
nand U12456 (N_12456,N_11521,N_11494);
and U12457 (N_12457,N_11689,N_11924);
and U12458 (N_12458,N_11341,N_11639);
xnor U12459 (N_12459,N_11694,N_11773);
xor U12460 (N_12460,N_11930,N_11625);
xnor U12461 (N_12461,N_11916,N_11428);
and U12462 (N_12462,N_11211,N_11154);
xor U12463 (N_12463,N_11456,N_11069);
xor U12464 (N_12464,N_11680,N_11746);
nand U12465 (N_12465,N_11855,N_11190);
nand U12466 (N_12466,N_11777,N_11504);
or U12467 (N_12467,N_11474,N_11972);
and U12468 (N_12468,N_11152,N_11413);
or U12469 (N_12469,N_11830,N_11603);
nor U12470 (N_12470,N_11232,N_11036);
nor U12471 (N_12471,N_11560,N_11216);
nand U12472 (N_12472,N_11750,N_11685);
nand U12473 (N_12473,N_11014,N_11208);
nor U12474 (N_12474,N_11557,N_11442);
nand U12475 (N_12475,N_11663,N_11627);
or U12476 (N_12476,N_11349,N_11620);
nor U12477 (N_12477,N_11781,N_11145);
and U12478 (N_12478,N_11571,N_11288);
nand U12479 (N_12479,N_11174,N_11647);
or U12480 (N_12480,N_11979,N_11628);
nand U12481 (N_12481,N_11702,N_11592);
xnor U12482 (N_12482,N_11705,N_11158);
nor U12483 (N_12483,N_11084,N_11616);
nand U12484 (N_12484,N_11714,N_11317);
and U12485 (N_12485,N_11448,N_11886);
or U12486 (N_12486,N_11988,N_11684);
nor U12487 (N_12487,N_11390,N_11594);
xor U12488 (N_12488,N_11025,N_11844);
xor U12489 (N_12489,N_11291,N_11738);
nor U12490 (N_12490,N_11167,N_11863);
or U12491 (N_12491,N_11046,N_11704);
nor U12492 (N_12492,N_11953,N_11203);
xor U12493 (N_12493,N_11757,N_11732);
xnor U12494 (N_12494,N_11790,N_11059);
xor U12495 (N_12495,N_11002,N_11269);
nand U12496 (N_12496,N_11181,N_11915);
nor U12497 (N_12497,N_11549,N_11295);
xor U12498 (N_12498,N_11598,N_11008);
nor U12499 (N_12499,N_11315,N_11888);
nor U12500 (N_12500,N_11104,N_11396);
and U12501 (N_12501,N_11846,N_11603);
xnor U12502 (N_12502,N_11966,N_11121);
or U12503 (N_12503,N_11792,N_11782);
nand U12504 (N_12504,N_11961,N_11721);
xor U12505 (N_12505,N_11443,N_11421);
xnor U12506 (N_12506,N_11325,N_11218);
nor U12507 (N_12507,N_11060,N_11201);
xnor U12508 (N_12508,N_11584,N_11541);
or U12509 (N_12509,N_11156,N_11896);
xnor U12510 (N_12510,N_11250,N_11097);
xor U12511 (N_12511,N_11113,N_11109);
or U12512 (N_12512,N_11413,N_11815);
nand U12513 (N_12513,N_11085,N_11423);
xor U12514 (N_12514,N_11238,N_11152);
xor U12515 (N_12515,N_11397,N_11918);
xnor U12516 (N_12516,N_11523,N_11459);
nand U12517 (N_12517,N_11070,N_11443);
xnor U12518 (N_12518,N_11431,N_11213);
nor U12519 (N_12519,N_11984,N_11280);
nor U12520 (N_12520,N_11783,N_11010);
xnor U12521 (N_12521,N_11351,N_11119);
or U12522 (N_12522,N_11676,N_11640);
nor U12523 (N_12523,N_11225,N_11378);
or U12524 (N_12524,N_11812,N_11738);
and U12525 (N_12525,N_11095,N_11956);
or U12526 (N_12526,N_11318,N_11113);
nand U12527 (N_12527,N_11190,N_11196);
nor U12528 (N_12528,N_11315,N_11430);
nand U12529 (N_12529,N_11394,N_11984);
or U12530 (N_12530,N_11984,N_11001);
nand U12531 (N_12531,N_11592,N_11618);
or U12532 (N_12532,N_11676,N_11107);
xnor U12533 (N_12533,N_11681,N_11736);
xnor U12534 (N_12534,N_11507,N_11164);
and U12535 (N_12535,N_11417,N_11288);
and U12536 (N_12536,N_11694,N_11247);
or U12537 (N_12537,N_11815,N_11375);
or U12538 (N_12538,N_11088,N_11670);
nand U12539 (N_12539,N_11508,N_11255);
xnor U12540 (N_12540,N_11681,N_11547);
or U12541 (N_12541,N_11605,N_11780);
xor U12542 (N_12542,N_11015,N_11271);
nand U12543 (N_12543,N_11142,N_11000);
and U12544 (N_12544,N_11946,N_11776);
nand U12545 (N_12545,N_11391,N_11612);
and U12546 (N_12546,N_11354,N_11485);
nand U12547 (N_12547,N_11505,N_11272);
nand U12548 (N_12548,N_11608,N_11939);
nand U12549 (N_12549,N_11252,N_11095);
or U12550 (N_12550,N_11304,N_11564);
or U12551 (N_12551,N_11601,N_11867);
nand U12552 (N_12552,N_11552,N_11400);
and U12553 (N_12553,N_11969,N_11228);
nor U12554 (N_12554,N_11289,N_11829);
or U12555 (N_12555,N_11397,N_11296);
and U12556 (N_12556,N_11638,N_11130);
or U12557 (N_12557,N_11118,N_11274);
nand U12558 (N_12558,N_11450,N_11309);
nand U12559 (N_12559,N_11728,N_11057);
nor U12560 (N_12560,N_11039,N_11826);
and U12561 (N_12561,N_11524,N_11063);
nor U12562 (N_12562,N_11166,N_11358);
xor U12563 (N_12563,N_11280,N_11495);
nand U12564 (N_12564,N_11551,N_11495);
nand U12565 (N_12565,N_11460,N_11629);
nand U12566 (N_12566,N_11034,N_11967);
or U12567 (N_12567,N_11845,N_11268);
nor U12568 (N_12568,N_11990,N_11261);
or U12569 (N_12569,N_11550,N_11375);
or U12570 (N_12570,N_11852,N_11952);
nor U12571 (N_12571,N_11102,N_11824);
and U12572 (N_12572,N_11082,N_11422);
nor U12573 (N_12573,N_11530,N_11664);
xnor U12574 (N_12574,N_11692,N_11600);
nor U12575 (N_12575,N_11544,N_11324);
nor U12576 (N_12576,N_11878,N_11490);
and U12577 (N_12577,N_11799,N_11576);
nand U12578 (N_12578,N_11267,N_11262);
nor U12579 (N_12579,N_11227,N_11156);
xnor U12580 (N_12580,N_11715,N_11069);
and U12581 (N_12581,N_11390,N_11389);
and U12582 (N_12582,N_11776,N_11750);
or U12583 (N_12583,N_11453,N_11908);
nand U12584 (N_12584,N_11387,N_11937);
nand U12585 (N_12585,N_11558,N_11800);
and U12586 (N_12586,N_11110,N_11843);
nor U12587 (N_12587,N_11843,N_11541);
nor U12588 (N_12588,N_11758,N_11542);
or U12589 (N_12589,N_11749,N_11476);
or U12590 (N_12590,N_11172,N_11906);
or U12591 (N_12591,N_11731,N_11638);
xnor U12592 (N_12592,N_11829,N_11269);
or U12593 (N_12593,N_11301,N_11750);
and U12594 (N_12594,N_11782,N_11029);
and U12595 (N_12595,N_11968,N_11496);
xnor U12596 (N_12596,N_11434,N_11550);
nand U12597 (N_12597,N_11648,N_11378);
and U12598 (N_12598,N_11740,N_11210);
or U12599 (N_12599,N_11162,N_11072);
and U12600 (N_12600,N_11083,N_11275);
and U12601 (N_12601,N_11066,N_11879);
and U12602 (N_12602,N_11056,N_11871);
xor U12603 (N_12603,N_11247,N_11858);
and U12604 (N_12604,N_11208,N_11356);
xnor U12605 (N_12605,N_11444,N_11263);
or U12606 (N_12606,N_11512,N_11226);
nand U12607 (N_12607,N_11078,N_11448);
nor U12608 (N_12608,N_11830,N_11320);
and U12609 (N_12609,N_11539,N_11963);
nor U12610 (N_12610,N_11708,N_11274);
nor U12611 (N_12611,N_11910,N_11473);
nor U12612 (N_12612,N_11947,N_11409);
and U12613 (N_12613,N_11203,N_11506);
and U12614 (N_12614,N_11202,N_11733);
xor U12615 (N_12615,N_11437,N_11725);
xnor U12616 (N_12616,N_11446,N_11444);
xnor U12617 (N_12617,N_11974,N_11957);
xor U12618 (N_12618,N_11942,N_11350);
and U12619 (N_12619,N_11483,N_11133);
and U12620 (N_12620,N_11887,N_11345);
nand U12621 (N_12621,N_11457,N_11750);
nor U12622 (N_12622,N_11609,N_11702);
nand U12623 (N_12623,N_11158,N_11259);
nor U12624 (N_12624,N_11172,N_11982);
or U12625 (N_12625,N_11504,N_11691);
and U12626 (N_12626,N_11257,N_11761);
and U12627 (N_12627,N_11817,N_11406);
nor U12628 (N_12628,N_11296,N_11352);
and U12629 (N_12629,N_11040,N_11562);
nor U12630 (N_12630,N_11888,N_11601);
nand U12631 (N_12631,N_11523,N_11906);
nand U12632 (N_12632,N_11492,N_11237);
nand U12633 (N_12633,N_11944,N_11005);
nor U12634 (N_12634,N_11658,N_11440);
or U12635 (N_12635,N_11837,N_11366);
and U12636 (N_12636,N_11088,N_11659);
nor U12637 (N_12637,N_11936,N_11839);
and U12638 (N_12638,N_11279,N_11240);
and U12639 (N_12639,N_11653,N_11613);
nor U12640 (N_12640,N_11338,N_11453);
and U12641 (N_12641,N_11393,N_11262);
or U12642 (N_12642,N_11179,N_11019);
or U12643 (N_12643,N_11513,N_11188);
nand U12644 (N_12644,N_11606,N_11414);
or U12645 (N_12645,N_11083,N_11852);
or U12646 (N_12646,N_11383,N_11323);
or U12647 (N_12647,N_11196,N_11826);
and U12648 (N_12648,N_11365,N_11782);
xnor U12649 (N_12649,N_11868,N_11610);
xnor U12650 (N_12650,N_11660,N_11651);
nor U12651 (N_12651,N_11523,N_11961);
nand U12652 (N_12652,N_11675,N_11082);
nor U12653 (N_12653,N_11936,N_11235);
and U12654 (N_12654,N_11269,N_11615);
nor U12655 (N_12655,N_11874,N_11788);
nand U12656 (N_12656,N_11798,N_11732);
or U12657 (N_12657,N_11066,N_11634);
nand U12658 (N_12658,N_11258,N_11846);
and U12659 (N_12659,N_11440,N_11136);
or U12660 (N_12660,N_11507,N_11312);
xnor U12661 (N_12661,N_11202,N_11975);
nor U12662 (N_12662,N_11338,N_11936);
and U12663 (N_12663,N_11550,N_11948);
nand U12664 (N_12664,N_11348,N_11282);
nand U12665 (N_12665,N_11964,N_11459);
nor U12666 (N_12666,N_11978,N_11308);
nor U12667 (N_12667,N_11479,N_11383);
nand U12668 (N_12668,N_11201,N_11486);
nand U12669 (N_12669,N_11099,N_11247);
nand U12670 (N_12670,N_11539,N_11347);
and U12671 (N_12671,N_11991,N_11043);
nand U12672 (N_12672,N_11365,N_11262);
nand U12673 (N_12673,N_11773,N_11136);
nor U12674 (N_12674,N_11795,N_11115);
nand U12675 (N_12675,N_11771,N_11249);
xnor U12676 (N_12676,N_11608,N_11629);
and U12677 (N_12677,N_11367,N_11282);
and U12678 (N_12678,N_11224,N_11011);
and U12679 (N_12679,N_11657,N_11423);
and U12680 (N_12680,N_11636,N_11080);
xnor U12681 (N_12681,N_11619,N_11267);
and U12682 (N_12682,N_11465,N_11737);
xor U12683 (N_12683,N_11771,N_11728);
or U12684 (N_12684,N_11896,N_11136);
nand U12685 (N_12685,N_11238,N_11527);
and U12686 (N_12686,N_11006,N_11062);
xnor U12687 (N_12687,N_11926,N_11197);
xor U12688 (N_12688,N_11621,N_11384);
nor U12689 (N_12689,N_11537,N_11386);
and U12690 (N_12690,N_11670,N_11496);
nand U12691 (N_12691,N_11654,N_11139);
and U12692 (N_12692,N_11516,N_11726);
or U12693 (N_12693,N_11764,N_11451);
nor U12694 (N_12694,N_11812,N_11823);
or U12695 (N_12695,N_11109,N_11803);
nor U12696 (N_12696,N_11898,N_11310);
nand U12697 (N_12697,N_11311,N_11702);
nand U12698 (N_12698,N_11958,N_11094);
or U12699 (N_12699,N_11557,N_11494);
xor U12700 (N_12700,N_11348,N_11389);
nand U12701 (N_12701,N_11735,N_11027);
and U12702 (N_12702,N_11032,N_11890);
xor U12703 (N_12703,N_11009,N_11368);
nand U12704 (N_12704,N_11905,N_11771);
and U12705 (N_12705,N_11769,N_11635);
xnor U12706 (N_12706,N_11837,N_11259);
nand U12707 (N_12707,N_11083,N_11399);
xor U12708 (N_12708,N_11719,N_11979);
or U12709 (N_12709,N_11149,N_11146);
or U12710 (N_12710,N_11098,N_11782);
and U12711 (N_12711,N_11934,N_11632);
and U12712 (N_12712,N_11747,N_11570);
nand U12713 (N_12713,N_11388,N_11747);
xor U12714 (N_12714,N_11805,N_11052);
nand U12715 (N_12715,N_11035,N_11146);
xor U12716 (N_12716,N_11354,N_11620);
and U12717 (N_12717,N_11818,N_11857);
nand U12718 (N_12718,N_11001,N_11334);
nor U12719 (N_12719,N_11371,N_11313);
nor U12720 (N_12720,N_11560,N_11380);
nor U12721 (N_12721,N_11856,N_11343);
nand U12722 (N_12722,N_11393,N_11903);
xnor U12723 (N_12723,N_11654,N_11595);
and U12724 (N_12724,N_11725,N_11669);
and U12725 (N_12725,N_11727,N_11203);
xor U12726 (N_12726,N_11342,N_11954);
xnor U12727 (N_12727,N_11725,N_11072);
nand U12728 (N_12728,N_11916,N_11733);
nor U12729 (N_12729,N_11668,N_11832);
nor U12730 (N_12730,N_11718,N_11188);
or U12731 (N_12731,N_11142,N_11589);
nor U12732 (N_12732,N_11026,N_11892);
xor U12733 (N_12733,N_11921,N_11073);
or U12734 (N_12734,N_11250,N_11125);
or U12735 (N_12735,N_11689,N_11828);
or U12736 (N_12736,N_11433,N_11321);
or U12737 (N_12737,N_11572,N_11197);
xnor U12738 (N_12738,N_11063,N_11224);
nor U12739 (N_12739,N_11679,N_11248);
nor U12740 (N_12740,N_11208,N_11089);
or U12741 (N_12741,N_11685,N_11510);
xor U12742 (N_12742,N_11173,N_11150);
or U12743 (N_12743,N_11995,N_11564);
xor U12744 (N_12744,N_11035,N_11469);
and U12745 (N_12745,N_11358,N_11904);
nand U12746 (N_12746,N_11401,N_11104);
nor U12747 (N_12747,N_11056,N_11798);
nand U12748 (N_12748,N_11768,N_11333);
and U12749 (N_12749,N_11504,N_11291);
xnor U12750 (N_12750,N_11259,N_11159);
nand U12751 (N_12751,N_11963,N_11872);
xnor U12752 (N_12752,N_11297,N_11599);
nand U12753 (N_12753,N_11789,N_11635);
nand U12754 (N_12754,N_11845,N_11640);
xnor U12755 (N_12755,N_11701,N_11652);
nand U12756 (N_12756,N_11562,N_11839);
nor U12757 (N_12757,N_11723,N_11714);
and U12758 (N_12758,N_11643,N_11636);
nand U12759 (N_12759,N_11000,N_11096);
and U12760 (N_12760,N_11698,N_11989);
or U12761 (N_12761,N_11795,N_11288);
xnor U12762 (N_12762,N_11532,N_11189);
nand U12763 (N_12763,N_11960,N_11565);
nor U12764 (N_12764,N_11545,N_11132);
and U12765 (N_12765,N_11564,N_11045);
and U12766 (N_12766,N_11531,N_11391);
xnor U12767 (N_12767,N_11422,N_11144);
and U12768 (N_12768,N_11743,N_11789);
nor U12769 (N_12769,N_11392,N_11165);
nor U12770 (N_12770,N_11177,N_11840);
nor U12771 (N_12771,N_11172,N_11799);
nor U12772 (N_12772,N_11552,N_11524);
nor U12773 (N_12773,N_11473,N_11478);
or U12774 (N_12774,N_11075,N_11520);
and U12775 (N_12775,N_11523,N_11124);
or U12776 (N_12776,N_11269,N_11475);
xor U12777 (N_12777,N_11612,N_11881);
and U12778 (N_12778,N_11514,N_11574);
or U12779 (N_12779,N_11090,N_11641);
nor U12780 (N_12780,N_11107,N_11645);
nand U12781 (N_12781,N_11421,N_11658);
or U12782 (N_12782,N_11380,N_11255);
and U12783 (N_12783,N_11437,N_11155);
and U12784 (N_12784,N_11757,N_11559);
and U12785 (N_12785,N_11837,N_11126);
and U12786 (N_12786,N_11446,N_11939);
nand U12787 (N_12787,N_11505,N_11247);
nor U12788 (N_12788,N_11412,N_11843);
nor U12789 (N_12789,N_11347,N_11510);
and U12790 (N_12790,N_11609,N_11858);
nand U12791 (N_12791,N_11730,N_11252);
and U12792 (N_12792,N_11204,N_11568);
and U12793 (N_12793,N_11731,N_11649);
and U12794 (N_12794,N_11497,N_11086);
nand U12795 (N_12795,N_11821,N_11297);
nand U12796 (N_12796,N_11477,N_11969);
and U12797 (N_12797,N_11888,N_11132);
nor U12798 (N_12798,N_11246,N_11488);
and U12799 (N_12799,N_11545,N_11654);
and U12800 (N_12800,N_11781,N_11129);
and U12801 (N_12801,N_11942,N_11919);
nor U12802 (N_12802,N_11817,N_11396);
nor U12803 (N_12803,N_11835,N_11785);
xnor U12804 (N_12804,N_11940,N_11457);
or U12805 (N_12805,N_11959,N_11501);
and U12806 (N_12806,N_11820,N_11342);
and U12807 (N_12807,N_11572,N_11496);
nor U12808 (N_12808,N_11291,N_11957);
and U12809 (N_12809,N_11574,N_11217);
xnor U12810 (N_12810,N_11791,N_11517);
xnor U12811 (N_12811,N_11069,N_11301);
and U12812 (N_12812,N_11572,N_11708);
and U12813 (N_12813,N_11365,N_11667);
and U12814 (N_12814,N_11772,N_11617);
and U12815 (N_12815,N_11900,N_11964);
nand U12816 (N_12816,N_11402,N_11601);
xor U12817 (N_12817,N_11213,N_11773);
nor U12818 (N_12818,N_11624,N_11614);
and U12819 (N_12819,N_11818,N_11098);
nor U12820 (N_12820,N_11324,N_11677);
and U12821 (N_12821,N_11646,N_11997);
nor U12822 (N_12822,N_11126,N_11591);
nand U12823 (N_12823,N_11595,N_11524);
nor U12824 (N_12824,N_11787,N_11888);
and U12825 (N_12825,N_11530,N_11232);
and U12826 (N_12826,N_11569,N_11991);
xor U12827 (N_12827,N_11947,N_11168);
nand U12828 (N_12828,N_11730,N_11278);
or U12829 (N_12829,N_11219,N_11382);
or U12830 (N_12830,N_11326,N_11536);
or U12831 (N_12831,N_11156,N_11897);
xor U12832 (N_12832,N_11980,N_11973);
or U12833 (N_12833,N_11025,N_11366);
nor U12834 (N_12834,N_11375,N_11482);
and U12835 (N_12835,N_11884,N_11994);
or U12836 (N_12836,N_11088,N_11691);
and U12837 (N_12837,N_11525,N_11550);
and U12838 (N_12838,N_11945,N_11956);
nand U12839 (N_12839,N_11769,N_11573);
and U12840 (N_12840,N_11890,N_11708);
and U12841 (N_12841,N_11568,N_11174);
nor U12842 (N_12842,N_11671,N_11431);
nand U12843 (N_12843,N_11068,N_11071);
and U12844 (N_12844,N_11080,N_11529);
and U12845 (N_12845,N_11073,N_11717);
nand U12846 (N_12846,N_11284,N_11963);
or U12847 (N_12847,N_11834,N_11092);
and U12848 (N_12848,N_11540,N_11784);
nor U12849 (N_12849,N_11190,N_11248);
xnor U12850 (N_12850,N_11306,N_11556);
or U12851 (N_12851,N_11185,N_11816);
xnor U12852 (N_12852,N_11889,N_11780);
and U12853 (N_12853,N_11073,N_11220);
and U12854 (N_12854,N_11481,N_11065);
and U12855 (N_12855,N_11210,N_11555);
xor U12856 (N_12856,N_11510,N_11521);
or U12857 (N_12857,N_11537,N_11224);
xnor U12858 (N_12858,N_11430,N_11361);
or U12859 (N_12859,N_11717,N_11307);
nor U12860 (N_12860,N_11914,N_11223);
and U12861 (N_12861,N_11039,N_11417);
nand U12862 (N_12862,N_11554,N_11633);
or U12863 (N_12863,N_11109,N_11065);
nand U12864 (N_12864,N_11934,N_11610);
nand U12865 (N_12865,N_11497,N_11247);
and U12866 (N_12866,N_11744,N_11683);
and U12867 (N_12867,N_11993,N_11664);
nor U12868 (N_12868,N_11755,N_11914);
nor U12869 (N_12869,N_11135,N_11039);
xnor U12870 (N_12870,N_11450,N_11593);
nor U12871 (N_12871,N_11989,N_11890);
or U12872 (N_12872,N_11889,N_11744);
and U12873 (N_12873,N_11837,N_11106);
or U12874 (N_12874,N_11800,N_11142);
xor U12875 (N_12875,N_11947,N_11197);
nor U12876 (N_12876,N_11331,N_11698);
or U12877 (N_12877,N_11080,N_11972);
or U12878 (N_12878,N_11075,N_11747);
xnor U12879 (N_12879,N_11684,N_11263);
or U12880 (N_12880,N_11233,N_11518);
nor U12881 (N_12881,N_11989,N_11935);
nor U12882 (N_12882,N_11579,N_11521);
xor U12883 (N_12883,N_11946,N_11530);
and U12884 (N_12884,N_11496,N_11609);
and U12885 (N_12885,N_11849,N_11787);
nor U12886 (N_12886,N_11020,N_11140);
or U12887 (N_12887,N_11701,N_11260);
and U12888 (N_12888,N_11205,N_11806);
or U12889 (N_12889,N_11329,N_11566);
nand U12890 (N_12890,N_11245,N_11035);
and U12891 (N_12891,N_11024,N_11014);
or U12892 (N_12892,N_11315,N_11476);
nor U12893 (N_12893,N_11604,N_11404);
xor U12894 (N_12894,N_11245,N_11811);
nand U12895 (N_12895,N_11299,N_11257);
and U12896 (N_12896,N_11711,N_11365);
xor U12897 (N_12897,N_11943,N_11535);
or U12898 (N_12898,N_11371,N_11548);
nand U12899 (N_12899,N_11186,N_11278);
xor U12900 (N_12900,N_11402,N_11279);
nand U12901 (N_12901,N_11713,N_11767);
and U12902 (N_12902,N_11729,N_11924);
and U12903 (N_12903,N_11030,N_11396);
and U12904 (N_12904,N_11204,N_11257);
nor U12905 (N_12905,N_11206,N_11728);
and U12906 (N_12906,N_11140,N_11421);
xnor U12907 (N_12907,N_11253,N_11045);
and U12908 (N_12908,N_11194,N_11691);
xor U12909 (N_12909,N_11751,N_11785);
xor U12910 (N_12910,N_11060,N_11755);
and U12911 (N_12911,N_11013,N_11551);
and U12912 (N_12912,N_11797,N_11246);
nor U12913 (N_12913,N_11923,N_11559);
nor U12914 (N_12914,N_11322,N_11627);
and U12915 (N_12915,N_11762,N_11287);
nor U12916 (N_12916,N_11392,N_11136);
xor U12917 (N_12917,N_11974,N_11539);
nor U12918 (N_12918,N_11042,N_11414);
nor U12919 (N_12919,N_11351,N_11806);
nand U12920 (N_12920,N_11369,N_11806);
and U12921 (N_12921,N_11062,N_11310);
nor U12922 (N_12922,N_11808,N_11584);
or U12923 (N_12923,N_11279,N_11884);
and U12924 (N_12924,N_11945,N_11364);
or U12925 (N_12925,N_11976,N_11312);
and U12926 (N_12926,N_11334,N_11013);
or U12927 (N_12927,N_11048,N_11973);
nand U12928 (N_12928,N_11211,N_11834);
or U12929 (N_12929,N_11379,N_11963);
or U12930 (N_12930,N_11112,N_11807);
nor U12931 (N_12931,N_11229,N_11324);
nor U12932 (N_12932,N_11485,N_11069);
nand U12933 (N_12933,N_11761,N_11660);
nand U12934 (N_12934,N_11829,N_11642);
and U12935 (N_12935,N_11720,N_11075);
nor U12936 (N_12936,N_11285,N_11085);
and U12937 (N_12937,N_11259,N_11116);
nand U12938 (N_12938,N_11347,N_11995);
xnor U12939 (N_12939,N_11062,N_11678);
nor U12940 (N_12940,N_11450,N_11109);
nand U12941 (N_12941,N_11919,N_11177);
xor U12942 (N_12942,N_11441,N_11621);
or U12943 (N_12943,N_11285,N_11602);
xnor U12944 (N_12944,N_11249,N_11402);
and U12945 (N_12945,N_11831,N_11329);
xnor U12946 (N_12946,N_11281,N_11516);
xnor U12947 (N_12947,N_11556,N_11113);
or U12948 (N_12948,N_11200,N_11767);
and U12949 (N_12949,N_11593,N_11533);
and U12950 (N_12950,N_11973,N_11518);
and U12951 (N_12951,N_11688,N_11502);
nand U12952 (N_12952,N_11821,N_11606);
xor U12953 (N_12953,N_11782,N_11341);
nor U12954 (N_12954,N_11429,N_11559);
or U12955 (N_12955,N_11339,N_11294);
xor U12956 (N_12956,N_11298,N_11389);
xnor U12957 (N_12957,N_11643,N_11126);
and U12958 (N_12958,N_11764,N_11053);
and U12959 (N_12959,N_11301,N_11376);
and U12960 (N_12960,N_11463,N_11769);
or U12961 (N_12961,N_11461,N_11712);
nor U12962 (N_12962,N_11154,N_11791);
nor U12963 (N_12963,N_11903,N_11495);
nor U12964 (N_12964,N_11848,N_11956);
or U12965 (N_12965,N_11091,N_11485);
xor U12966 (N_12966,N_11381,N_11534);
or U12967 (N_12967,N_11800,N_11845);
nor U12968 (N_12968,N_11368,N_11907);
nand U12969 (N_12969,N_11708,N_11636);
or U12970 (N_12970,N_11890,N_11617);
nor U12971 (N_12971,N_11417,N_11447);
and U12972 (N_12972,N_11534,N_11879);
or U12973 (N_12973,N_11956,N_11169);
or U12974 (N_12974,N_11389,N_11443);
nor U12975 (N_12975,N_11770,N_11052);
xnor U12976 (N_12976,N_11814,N_11392);
nor U12977 (N_12977,N_11778,N_11194);
nand U12978 (N_12978,N_11147,N_11586);
or U12979 (N_12979,N_11614,N_11036);
xnor U12980 (N_12980,N_11666,N_11895);
nand U12981 (N_12981,N_11503,N_11672);
nand U12982 (N_12982,N_11912,N_11151);
nor U12983 (N_12983,N_11332,N_11702);
nand U12984 (N_12984,N_11425,N_11290);
xnor U12985 (N_12985,N_11734,N_11315);
or U12986 (N_12986,N_11745,N_11540);
and U12987 (N_12987,N_11629,N_11817);
nand U12988 (N_12988,N_11603,N_11741);
and U12989 (N_12989,N_11826,N_11953);
nor U12990 (N_12990,N_11004,N_11180);
xnor U12991 (N_12991,N_11430,N_11312);
nand U12992 (N_12992,N_11947,N_11968);
nor U12993 (N_12993,N_11836,N_11291);
or U12994 (N_12994,N_11004,N_11999);
nand U12995 (N_12995,N_11987,N_11460);
nand U12996 (N_12996,N_11457,N_11433);
nand U12997 (N_12997,N_11685,N_11718);
and U12998 (N_12998,N_11452,N_11358);
xnor U12999 (N_12999,N_11661,N_11263);
nand U13000 (N_13000,N_12273,N_12262);
nor U13001 (N_13001,N_12597,N_12233);
nor U13002 (N_13002,N_12850,N_12056);
or U13003 (N_13003,N_12250,N_12317);
nor U13004 (N_13004,N_12138,N_12826);
and U13005 (N_13005,N_12249,N_12482);
xnor U13006 (N_13006,N_12432,N_12076);
nand U13007 (N_13007,N_12321,N_12707);
nor U13008 (N_13008,N_12187,N_12116);
nor U13009 (N_13009,N_12906,N_12928);
and U13010 (N_13010,N_12100,N_12157);
xor U13011 (N_13011,N_12823,N_12182);
and U13012 (N_13012,N_12111,N_12419);
nand U13013 (N_13013,N_12325,N_12203);
nand U13014 (N_13014,N_12260,N_12082);
xnor U13015 (N_13015,N_12980,N_12350);
xnor U13016 (N_13016,N_12814,N_12745);
and U13017 (N_13017,N_12037,N_12238);
nor U13018 (N_13018,N_12429,N_12957);
nor U13019 (N_13019,N_12228,N_12589);
and U13020 (N_13020,N_12889,N_12099);
nand U13021 (N_13021,N_12715,N_12806);
nand U13022 (N_13022,N_12398,N_12127);
xor U13023 (N_13023,N_12593,N_12668);
and U13024 (N_13024,N_12684,N_12710);
or U13025 (N_13025,N_12909,N_12275);
nor U13026 (N_13026,N_12034,N_12102);
and U13027 (N_13027,N_12208,N_12641);
nand U13028 (N_13028,N_12501,N_12782);
nor U13029 (N_13029,N_12759,N_12800);
nor U13030 (N_13030,N_12451,N_12898);
or U13031 (N_13031,N_12513,N_12504);
or U13032 (N_13032,N_12661,N_12708);
xor U13033 (N_13033,N_12590,N_12302);
and U13034 (N_13034,N_12573,N_12952);
nor U13035 (N_13035,N_12109,N_12761);
nor U13036 (N_13036,N_12825,N_12071);
xor U13037 (N_13037,N_12447,N_12380);
and U13038 (N_13038,N_12498,N_12882);
and U13039 (N_13039,N_12490,N_12990);
nor U13040 (N_13040,N_12748,N_12562);
xor U13041 (N_13041,N_12306,N_12159);
nand U13042 (N_13042,N_12692,N_12899);
nor U13043 (N_13043,N_12625,N_12023);
and U13044 (N_13044,N_12881,N_12717);
or U13045 (N_13045,N_12489,N_12267);
nor U13046 (N_13046,N_12971,N_12731);
xnor U13047 (N_13047,N_12105,N_12272);
nand U13048 (N_13048,N_12393,N_12564);
or U13049 (N_13049,N_12751,N_12179);
nor U13050 (N_13050,N_12902,N_12506);
nor U13051 (N_13051,N_12862,N_12367);
nand U13052 (N_13052,N_12728,N_12336);
and U13053 (N_13053,N_12505,N_12770);
nand U13054 (N_13054,N_12199,N_12397);
nor U13055 (N_13055,N_12491,N_12665);
nor U13056 (N_13056,N_12757,N_12720);
xnor U13057 (N_13057,N_12470,N_12112);
or U13058 (N_13058,N_12932,N_12176);
nor U13059 (N_13059,N_12209,N_12561);
or U13060 (N_13060,N_12531,N_12270);
and U13061 (N_13061,N_12614,N_12469);
or U13062 (N_13062,N_12872,N_12602);
and U13063 (N_13063,N_12320,N_12162);
xor U13064 (N_13064,N_12258,N_12125);
or U13065 (N_13065,N_12153,N_12274);
nand U13066 (N_13066,N_12938,N_12297);
nand U13067 (N_13067,N_12309,N_12402);
nor U13068 (N_13068,N_12815,N_12205);
and U13069 (N_13069,N_12345,N_12920);
xnor U13070 (N_13070,N_12647,N_12401);
nor U13071 (N_13071,N_12636,N_12310);
nor U13072 (N_13072,N_12655,N_12113);
nor U13073 (N_13073,N_12416,N_12523);
and U13074 (N_13074,N_12128,N_12992);
xor U13075 (N_13075,N_12388,N_12542);
nand U13076 (N_13076,N_12132,N_12328);
nand U13077 (N_13077,N_12516,N_12444);
or U13078 (N_13078,N_12958,N_12443);
nand U13079 (N_13079,N_12421,N_12148);
nor U13080 (N_13080,N_12340,N_12555);
nor U13081 (N_13081,N_12772,N_12338);
nand U13082 (N_13082,N_12846,N_12394);
xor U13083 (N_13083,N_12925,N_12033);
and U13084 (N_13084,N_12893,N_12546);
nor U13085 (N_13085,N_12241,N_12239);
or U13086 (N_13086,N_12824,N_12658);
or U13087 (N_13087,N_12609,N_12522);
xor U13088 (N_13088,N_12372,N_12299);
xnor U13089 (N_13089,N_12006,N_12487);
and U13090 (N_13090,N_12790,N_12866);
or U13091 (N_13091,N_12064,N_12956);
nor U13092 (N_13092,N_12103,N_12045);
nor U13093 (N_13093,N_12901,N_12106);
xnor U13094 (N_13094,N_12383,N_12156);
xor U13095 (N_13095,N_12089,N_12833);
nand U13096 (N_13096,N_12428,N_12507);
nor U13097 (N_13097,N_12934,N_12718);
nor U13098 (N_13098,N_12566,N_12189);
xnor U13099 (N_13099,N_12648,N_12769);
nor U13100 (N_13100,N_12596,N_12828);
or U13101 (N_13101,N_12514,N_12892);
xnor U13102 (N_13102,N_12931,N_12459);
and U13103 (N_13103,N_12049,N_12544);
and U13104 (N_13104,N_12400,N_12600);
nand U13105 (N_13105,N_12849,N_12797);
nor U13106 (N_13106,N_12948,N_12486);
and U13107 (N_13107,N_12694,N_12038);
xor U13108 (N_13108,N_12098,N_12151);
nand U13109 (N_13109,N_12509,N_12768);
or U13110 (N_13110,N_12879,N_12508);
or U13111 (N_13111,N_12622,N_12784);
or U13112 (N_13112,N_12677,N_12221);
nor U13113 (N_13113,N_12188,N_12155);
nand U13114 (N_13114,N_12888,N_12294);
nor U13115 (N_13115,N_12282,N_12935);
or U13116 (N_13116,N_12052,N_12407);
xor U13117 (N_13117,N_12540,N_12682);
and U13118 (N_13118,N_12142,N_12364);
and U13119 (N_13119,N_12235,N_12860);
or U13120 (N_13120,N_12805,N_12289);
or U13121 (N_13121,N_12462,N_12377);
nand U13122 (N_13122,N_12167,N_12081);
and U13123 (N_13123,N_12563,N_12281);
xnor U13124 (N_13124,N_12737,N_12870);
xor U13125 (N_13125,N_12859,N_12438);
xor U13126 (N_13126,N_12858,N_12979);
nor U13127 (N_13127,N_12568,N_12588);
or U13128 (N_13128,N_12532,N_12615);
and U13129 (N_13129,N_12816,N_12541);
nor U13130 (N_13130,N_12845,N_12936);
nand U13131 (N_13131,N_12864,N_12991);
xnor U13132 (N_13132,N_12131,N_12493);
and U13133 (N_13133,N_12732,N_12070);
and U13134 (N_13134,N_12043,N_12699);
nor U13135 (N_13135,N_12821,N_12019);
nor U13136 (N_13136,N_12868,N_12512);
nor U13137 (N_13137,N_12365,N_12631);
and U13138 (N_13138,N_12666,N_12766);
or U13139 (N_13139,N_12527,N_12242);
xnor U13140 (N_13140,N_12629,N_12255);
or U13141 (N_13141,N_12587,N_12009);
xnor U13142 (N_13142,N_12431,N_12724);
xor U13143 (N_13143,N_12164,N_12358);
xnor U13144 (N_13144,N_12765,N_12133);
nor U13145 (N_13145,N_12607,N_12366);
xnor U13146 (N_13146,N_12403,N_12729);
xnor U13147 (N_13147,N_12223,N_12706);
or U13148 (N_13148,N_12477,N_12954);
or U13149 (N_13149,N_12974,N_12497);
xnor U13150 (N_13150,N_12475,N_12329);
xnor U13151 (N_13151,N_12061,N_12580);
nand U13152 (N_13152,N_12093,N_12252);
nand U13153 (N_13153,N_12332,N_12022);
nand U13154 (N_13154,N_12547,N_12669);
nor U13155 (N_13155,N_12251,N_12474);
nand U13156 (N_13156,N_12080,N_12248);
nand U13157 (N_13157,N_12016,N_12741);
or U13158 (N_13158,N_12068,N_12192);
and U13159 (N_13159,N_12690,N_12680);
or U13160 (N_13160,N_12010,N_12337);
nand U13161 (N_13161,N_12617,N_12307);
nand U13162 (N_13162,N_12915,N_12288);
nor U13163 (N_13163,N_12437,N_12863);
xor U13164 (N_13164,N_12305,N_12619);
nor U13165 (N_13165,N_12108,N_12518);
nor U13166 (N_13166,N_12856,N_12054);
nor U13167 (N_13167,N_12807,N_12565);
or U13168 (N_13168,N_12802,N_12295);
nand U13169 (N_13169,N_12911,N_12704);
and U13170 (N_13170,N_12218,N_12002);
nand U13171 (N_13171,N_12472,N_12785);
xnor U13172 (N_13172,N_12018,N_12917);
and U13173 (N_13173,N_12375,N_12293);
or U13174 (N_13174,N_12650,N_12656);
and U13175 (N_13175,N_12308,N_12413);
nor U13176 (N_13176,N_12572,N_12749);
or U13177 (N_13177,N_12586,N_12492);
and U13178 (N_13178,N_12280,N_12986);
or U13179 (N_13179,N_12183,N_12149);
nor U13180 (N_13180,N_12534,N_12007);
xnor U13181 (N_13181,N_12129,N_12545);
or U13182 (N_13182,N_12869,N_12456);
nor U13183 (N_13183,N_12135,N_12659);
xor U13184 (N_13184,N_12319,N_12126);
nand U13185 (N_13185,N_12254,N_12977);
or U13186 (N_13186,N_12422,N_12570);
and U13187 (N_13187,N_12798,N_12657);
nor U13188 (N_13188,N_12754,N_12940);
xnor U13189 (N_13189,N_12137,N_12789);
nor U13190 (N_13190,N_12165,N_12743);
xnor U13191 (N_13191,N_12663,N_12044);
and U13192 (N_13192,N_12907,N_12341);
xor U13193 (N_13193,N_12993,N_12084);
nor U13194 (N_13194,N_12434,N_12670);
xnor U13195 (N_13195,N_12496,N_12796);
or U13196 (N_13196,N_12683,N_12623);
nand U13197 (N_13197,N_12723,N_12467);
and U13198 (N_13198,N_12458,N_12236);
and U13199 (N_13199,N_12463,N_12794);
or U13200 (N_13200,N_12894,N_12230);
and U13201 (N_13201,N_12628,N_12050);
or U13202 (N_13202,N_12713,N_12412);
and U13203 (N_13203,N_12689,N_12644);
xor U13204 (N_13204,N_12471,N_12696);
or U13205 (N_13205,N_12996,N_12829);
nor U13206 (N_13206,N_12842,N_12788);
xnor U13207 (N_13207,N_12021,N_12175);
nor U13208 (N_13208,N_12120,N_12261);
nand U13209 (N_13209,N_12312,N_12152);
xnor U13210 (N_13210,N_12466,N_12982);
nor U13211 (N_13211,N_12995,N_12722);
xor U13212 (N_13212,N_12853,N_12679);
xor U13213 (N_13213,N_12637,N_12180);
or U13214 (N_13214,N_12985,N_12781);
xnor U13215 (N_13215,N_12595,N_12897);
and U13216 (N_13216,N_12304,N_12296);
xnor U13217 (N_13217,N_12285,N_12537);
xnor U13218 (N_13218,N_12001,N_12483);
and U13219 (N_13219,N_12278,N_12613);
nor U13220 (N_13220,N_12652,N_12210);
or U13221 (N_13221,N_12989,N_12730);
or U13222 (N_13222,N_12225,N_12604);
xnor U13223 (N_13223,N_12951,N_12104);
nor U13224 (N_13224,N_12173,N_12725);
xor U13225 (N_13225,N_12583,N_12926);
xnor U13226 (N_13226,N_12791,N_12543);
nand U13227 (N_13227,N_12075,N_12237);
or U13228 (N_13228,N_12214,N_12793);
or U13229 (N_13229,N_12240,N_12479);
nor U13230 (N_13230,N_12921,N_12417);
nor U13231 (N_13231,N_12517,N_12929);
or U13232 (N_13232,N_12712,N_12257);
nor U13233 (N_13233,N_12141,N_12777);
nor U13234 (N_13234,N_12811,N_12392);
or U13235 (N_13235,N_12215,N_12753);
and U13236 (N_13236,N_12645,N_12716);
and U13237 (N_13237,N_12433,N_12124);
nor U13238 (N_13238,N_12763,N_12778);
nand U13239 (N_13239,N_12426,N_12334);
and U13240 (N_13240,N_12143,N_12758);
nand U13241 (N_13241,N_12220,N_12854);
and U13242 (N_13242,N_12158,N_12286);
and U13243 (N_13243,N_12762,N_12485);
nor U13244 (N_13244,N_12356,N_12502);
and U13245 (N_13245,N_12026,N_12499);
xor U13246 (N_13246,N_12174,N_12896);
and U13247 (N_13247,N_12119,N_12351);
or U13248 (N_13248,N_12681,N_12114);
or U13249 (N_13249,N_12391,N_12359);
nand U13250 (N_13250,N_12488,N_12072);
and U13251 (N_13251,N_12343,N_12736);
xor U13252 (N_13252,N_12714,N_12300);
nand U13253 (N_13253,N_12804,N_12840);
or U13254 (N_13254,N_12357,N_12454);
xor U13255 (N_13255,N_12315,N_12955);
nand U13256 (N_13256,N_12408,N_12646);
nor U13257 (N_13257,N_12943,N_12764);
nor U13258 (N_13258,N_12750,N_12515);
and U13259 (N_13259,N_12455,N_12322);
nand U13260 (N_13260,N_12352,N_12396);
nor U13261 (N_13261,N_12755,N_12626);
nand U13262 (N_13262,N_12145,N_12031);
xor U13263 (N_13263,N_12535,N_12301);
nor U13264 (N_13264,N_12953,N_12767);
xor U13265 (N_13265,N_12330,N_12548);
nand U13266 (N_13266,N_12110,N_12029);
nand U13267 (N_13267,N_12721,N_12354);
and U13268 (N_13268,N_12835,N_12115);
nor U13269 (N_13269,N_12344,N_12571);
nand U13270 (N_13270,N_12975,N_12405);
or U13271 (N_13271,N_12530,N_12083);
xnor U13272 (N_13272,N_12476,N_12290);
xor U13273 (N_13273,N_12937,N_12910);
nor U13274 (N_13274,N_12965,N_12933);
nand U13275 (N_13275,N_12253,N_12409);
nand U13276 (N_13276,N_12269,N_12808);
or U13277 (N_13277,N_12335,N_12945);
and U13278 (N_13278,N_12903,N_12386);
nand U13279 (N_13279,N_12101,N_12703);
nor U13280 (N_13280,N_12839,N_12967);
nor U13281 (N_13281,N_12424,N_12678);
nor U13282 (N_13282,N_12923,N_12976);
and U13283 (N_13283,N_12942,N_12983);
nor U13284 (N_13284,N_12649,N_12886);
or U13285 (N_13285,N_12349,N_12526);
or U13286 (N_13286,N_12449,N_12040);
xor U13287 (N_13287,N_12560,N_12078);
nor U13288 (N_13288,N_12012,N_12464);
nand U13289 (N_13289,N_12247,N_12074);
or U13290 (N_13290,N_12598,N_12177);
or U13291 (N_13291,N_12460,N_12771);
or U13292 (N_13292,N_12154,N_12196);
or U13293 (N_13293,N_12461,N_12369);
nand U13294 (N_13294,N_12733,N_12524);
nand U13295 (N_13295,N_12107,N_12674);
and U13296 (N_13296,N_12311,N_12918);
or U13297 (N_13297,N_12324,N_12867);
nand U13298 (N_13298,N_12066,N_12318);
or U13299 (N_13299,N_12117,N_12635);
xor U13300 (N_13300,N_12908,N_12355);
and U13301 (N_13301,N_12373,N_12582);
nor U13302 (N_13302,N_12191,N_12053);
nor U13303 (N_13303,N_12370,N_12848);
and U13304 (N_13304,N_12711,N_12667);
nor U13305 (N_13305,N_12146,N_12865);
nand U13306 (N_13306,N_12121,N_12139);
xnor U13307 (N_13307,N_12841,N_12944);
and U13308 (N_13308,N_12746,N_12618);
xor U13309 (N_13309,N_12640,N_12495);
or U13310 (N_13310,N_12973,N_12510);
xnor U13311 (N_13311,N_12435,N_12591);
and U13312 (N_13312,N_12144,N_12077);
or U13313 (N_13313,N_12246,N_12122);
nor U13314 (N_13314,N_12701,N_12441);
or U13315 (N_13315,N_12533,N_12567);
nand U13316 (N_13316,N_12291,N_12259);
and U13317 (N_13317,N_12283,N_12700);
xor U13318 (N_13318,N_12970,N_12327);
xnor U13319 (N_13319,N_12787,N_12818);
xnor U13320 (N_13320,N_12234,N_12981);
or U13321 (N_13321,N_12984,N_12653);
or U13322 (N_13322,N_12550,N_12091);
nor U13323 (N_13323,N_12672,N_12887);
nor U13324 (N_13324,N_12671,N_12776);
nand U13325 (N_13325,N_12691,N_12760);
nand U13326 (N_13326,N_12207,N_12381);
xnor U13327 (N_13327,N_12611,N_12685);
xor U13328 (N_13328,N_12738,N_12172);
xor U13329 (N_13329,N_12442,N_12195);
xor U13330 (N_13330,N_12994,N_12642);
and U13331 (N_13331,N_12592,N_12809);
or U13332 (N_13332,N_12536,N_12453);
xor U13333 (N_13333,N_12004,N_12844);
and U13334 (N_13334,N_12118,N_12065);
and U13335 (N_13335,N_12895,N_12185);
xor U13336 (N_13336,N_12206,N_12003);
nand U13337 (N_13337,N_12450,N_12316);
nor U13338 (N_13338,N_12877,N_12200);
nor U13339 (N_13339,N_12972,N_12035);
nand U13340 (N_13340,N_12968,N_12446);
nor U13341 (N_13341,N_12389,N_12384);
or U13342 (N_13342,N_12348,N_12688);
or U13343 (N_13343,N_12404,N_12079);
nand U13344 (N_13344,N_12998,N_12930);
xnor U13345 (N_13345,N_12222,N_12059);
xor U13346 (N_13346,N_12201,N_12660);
xnor U13347 (N_13347,N_12585,N_12439);
nand U13348 (N_13348,N_12014,N_12406);
nor U13349 (N_13349,N_12232,N_12773);
xor U13350 (N_13350,N_12134,N_12047);
xor U13351 (N_13351,N_12216,N_12181);
nor U13352 (N_13352,N_12525,N_12584);
xor U13353 (N_13353,N_12032,N_12468);
and U13354 (N_13354,N_12927,N_12742);
nand U13355 (N_13355,N_12639,N_12919);
nand U13356 (N_13356,N_12675,N_12436);
or U13357 (N_13357,N_12579,N_12997);
and U13358 (N_13358,N_12634,N_12687);
or U13359 (N_13359,N_12939,N_12184);
xor U13360 (N_13360,N_12612,N_12651);
or U13361 (N_13361,N_12632,N_12085);
xnor U13362 (N_13362,N_12339,N_12912);
and U13363 (N_13363,N_12385,N_12719);
nand U13364 (N_13364,N_12969,N_12415);
and U13365 (N_13365,N_12264,N_12539);
nor U13366 (N_13366,N_12136,N_12069);
and U13367 (N_13367,N_12204,N_12353);
or U13368 (N_13368,N_12734,N_12171);
and U13369 (N_13369,N_12884,N_12430);
xor U13370 (N_13370,N_12166,N_12051);
and U13371 (N_13371,N_12213,N_12374);
nor U13372 (N_13372,N_12905,N_12874);
or U13373 (N_13373,N_12511,N_12727);
or U13374 (N_13374,N_12654,N_12371);
nor U13375 (N_13375,N_12528,N_12662);
xnor U13376 (N_13376,N_12265,N_12000);
nand U13377 (N_13377,N_12620,N_12219);
and U13378 (N_13378,N_12160,N_12020);
or U13379 (N_13379,N_12123,N_12150);
nor U13380 (N_13380,N_12039,N_12017);
nand U13381 (N_13381,N_12287,N_12559);
nand U13382 (N_13382,N_12780,N_12838);
and U13383 (N_13383,N_12529,N_12057);
nand U13384 (N_13384,N_12941,N_12904);
and U13385 (N_13385,N_12852,N_12606);
nand U13386 (N_13386,N_12445,N_12411);
and U13387 (N_13387,N_12279,N_12885);
nor U13388 (N_13388,N_12871,N_12963);
nor U13389 (N_13389,N_12387,N_12817);
or U13390 (N_13390,N_12876,N_12420);
nor U13391 (N_13391,N_12030,N_12726);
or U13392 (N_13392,N_12538,N_12558);
nand U13393 (N_13393,N_12092,N_12055);
xnor U13394 (N_13394,N_12610,N_12088);
xor U13395 (N_13395,N_12601,N_12478);
nand U13396 (N_13396,N_12624,N_12575);
nor U13397 (N_13397,N_12520,N_12812);
nor U13398 (N_13398,N_12425,N_12028);
nand U13399 (N_13399,N_12735,N_12494);
nor U13400 (N_13400,N_12594,N_12630);
or U13401 (N_13401,N_12830,N_12914);
and U13402 (N_13402,N_12519,N_12783);
nand U13403 (N_13403,N_12827,N_12382);
or U13404 (N_13404,N_12966,N_12041);
xnor U13405 (N_13405,N_12695,N_12633);
or U13406 (N_13406,N_12803,N_12861);
and U13407 (N_13407,N_12553,N_12423);
or U13408 (N_13408,N_12605,N_12457);
nand U13409 (N_13409,N_12313,N_12087);
nor U13410 (N_13410,N_12978,N_12194);
xnor U13411 (N_13411,N_12913,N_12178);
nor U13412 (N_13412,N_12792,N_12857);
nor U13413 (N_13413,N_12097,N_12616);
or U13414 (N_13414,N_12950,N_12752);
nand U13415 (N_13415,N_12831,N_12130);
nor U13416 (N_13416,N_12303,N_12946);
or U13417 (N_13417,N_12747,N_12015);
or U13418 (N_13418,N_12961,N_12900);
nor U13419 (N_13419,N_12608,N_12024);
nand U13420 (N_13420,N_12922,N_12603);
or U13421 (N_13421,N_12227,N_12245);
nor U13422 (N_13422,N_12005,N_12569);
xnor U13423 (N_13423,N_12578,N_12576);
xor U13424 (N_13424,N_12577,N_12193);
xnor U13425 (N_13425,N_12465,N_12368);
nand U13426 (N_13426,N_12025,N_12036);
nand U13427 (N_13427,N_12820,N_12673);
nand U13428 (N_13428,N_12500,N_12964);
nand U13429 (N_13429,N_12774,N_12362);
nor U13430 (N_13430,N_12292,N_12410);
and U13431 (N_13431,N_12924,N_12027);
and U13432 (N_13432,N_12399,N_12073);
and U13433 (N_13433,N_12395,N_12202);
and U13434 (N_13434,N_12740,N_12836);
nand U13435 (N_13435,N_12008,N_12390);
nor U13436 (N_13436,N_12378,N_12484);
or U13437 (N_13437,N_12062,N_12481);
nand U13438 (N_13438,N_12161,N_12843);
or U13439 (N_13439,N_12891,N_12581);
nor U13440 (N_13440,N_12810,N_12452);
xnor U13441 (N_13441,N_12756,N_12949);
xnor U13442 (N_13442,N_12556,N_12880);
xnor U13443 (N_13443,N_12211,N_12284);
and U13444 (N_13444,N_12427,N_12873);
or U13445 (N_13445,N_12847,N_12224);
xor U13446 (N_13446,N_12627,N_12890);
nor U13447 (N_13447,N_12331,N_12060);
xor U13448 (N_13448,N_12298,N_12834);
nor U13449 (N_13449,N_12063,N_12960);
or U13450 (N_13450,N_12163,N_12086);
nor U13451 (N_13451,N_12226,N_12702);
and U13452 (N_13452,N_12801,N_12414);
nand U13453 (N_13453,N_12875,N_12878);
xnor U13454 (N_13454,N_12779,N_12169);
or U13455 (N_13455,N_12376,N_12947);
nand U13456 (N_13456,N_12744,N_12266);
xnor U13457 (N_13457,N_12686,N_12883);
nand U13458 (N_13458,N_12090,N_12314);
nand U13459 (N_13459,N_12698,N_12799);
or U13460 (N_13460,N_12094,N_12705);
nand U13461 (N_13461,N_12379,N_12557);
and U13462 (N_13462,N_12346,N_12418);
nor U13463 (N_13463,N_12697,N_12168);
and U13464 (N_13464,N_12231,N_12186);
nor U13465 (N_13465,N_12095,N_12813);
and U13466 (N_13466,N_12503,N_12048);
xor U13467 (N_13467,N_12277,N_12011);
nor U13468 (N_13468,N_12271,N_12837);
xor U13469 (N_13469,N_12551,N_12987);
nor U13470 (N_13470,N_12256,N_12521);
xor U13471 (N_13471,N_12323,N_12058);
and U13472 (N_13472,N_12212,N_12999);
and U13473 (N_13473,N_12147,N_12243);
or U13474 (N_13474,N_12440,N_12229);
xnor U13475 (N_13475,N_12347,N_12676);
or U13476 (N_13476,N_12709,N_12448);
or U13477 (N_13477,N_12197,N_12851);
xnor U13478 (N_13478,N_12096,N_12959);
nor U13479 (N_13479,N_12333,N_12962);
xnor U13480 (N_13480,N_12263,N_12822);
nand U13481 (N_13481,N_12276,N_12342);
nor U13482 (N_13482,N_12693,N_12190);
xnor U13483 (N_13483,N_12042,N_12046);
nand U13484 (N_13484,N_12574,N_12170);
or U13485 (N_13485,N_12916,N_12217);
nor U13486 (N_13486,N_12786,N_12361);
and U13487 (N_13487,N_12795,N_12664);
nand U13488 (N_13488,N_12198,N_12988);
xor U13489 (N_13489,N_12855,N_12326);
and U13490 (N_13490,N_12244,N_12599);
and U13491 (N_13491,N_12067,N_12621);
or U13492 (N_13492,N_12268,N_12013);
xnor U13493 (N_13493,N_12554,N_12480);
nor U13494 (N_13494,N_12360,N_12363);
nor U13495 (N_13495,N_12638,N_12140);
nand U13496 (N_13496,N_12552,N_12473);
or U13497 (N_13497,N_12739,N_12775);
nor U13498 (N_13498,N_12819,N_12832);
xnor U13499 (N_13499,N_12643,N_12549);
or U13500 (N_13500,N_12142,N_12289);
or U13501 (N_13501,N_12563,N_12067);
nand U13502 (N_13502,N_12352,N_12736);
nand U13503 (N_13503,N_12472,N_12743);
nor U13504 (N_13504,N_12621,N_12405);
or U13505 (N_13505,N_12314,N_12412);
nor U13506 (N_13506,N_12613,N_12538);
or U13507 (N_13507,N_12693,N_12579);
nor U13508 (N_13508,N_12522,N_12829);
xnor U13509 (N_13509,N_12286,N_12796);
nor U13510 (N_13510,N_12327,N_12493);
xor U13511 (N_13511,N_12257,N_12152);
xor U13512 (N_13512,N_12606,N_12775);
xor U13513 (N_13513,N_12007,N_12547);
or U13514 (N_13514,N_12380,N_12037);
xor U13515 (N_13515,N_12146,N_12724);
xor U13516 (N_13516,N_12644,N_12185);
nor U13517 (N_13517,N_12145,N_12641);
xor U13518 (N_13518,N_12964,N_12650);
xor U13519 (N_13519,N_12193,N_12619);
nor U13520 (N_13520,N_12507,N_12418);
or U13521 (N_13521,N_12093,N_12923);
or U13522 (N_13522,N_12069,N_12229);
and U13523 (N_13523,N_12930,N_12110);
or U13524 (N_13524,N_12576,N_12735);
and U13525 (N_13525,N_12036,N_12510);
nand U13526 (N_13526,N_12601,N_12144);
nor U13527 (N_13527,N_12894,N_12274);
nor U13528 (N_13528,N_12558,N_12070);
nand U13529 (N_13529,N_12330,N_12589);
or U13530 (N_13530,N_12315,N_12157);
and U13531 (N_13531,N_12271,N_12366);
xor U13532 (N_13532,N_12780,N_12473);
xnor U13533 (N_13533,N_12974,N_12610);
nor U13534 (N_13534,N_12105,N_12037);
nor U13535 (N_13535,N_12812,N_12636);
nor U13536 (N_13536,N_12222,N_12314);
xnor U13537 (N_13537,N_12401,N_12479);
nor U13538 (N_13538,N_12897,N_12901);
xnor U13539 (N_13539,N_12498,N_12586);
nor U13540 (N_13540,N_12354,N_12993);
nand U13541 (N_13541,N_12503,N_12919);
or U13542 (N_13542,N_12146,N_12760);
nor U13543 (N_13543,N_12618,N_12027);
nor U13544 (N_13544,N_12294,N_12788);
nand U13545 (N_13545,N_12977,N_12443);
nor U13546 (N_13546,N_12129,N_12696);
nor U13547 (N_13547,N_12040,N_12192);
nand U13548 (N_13548,N_12130,N_12083);
or U13549 (N_13549,N_12329,N_12993);
nand U13550 (N_13550,N_12720,N_12312);
and U13551 (N_13551,N_12274,N_12373);
xor U13552 (N_13552,N_12082,N_12662);
nand U13553 (N_13553,N_12405,N_12182);
xor U13554 (N_13554,N_12875,N_12782);
or U13555 (N_13555,N_12830,N_12863);
nand U13556 (N_13556,N_12168,N_12523);
xnor U13557 (N_13557,N_12567,N_12391);
and U13558 (N_13558,N_12760,N_12907);
nor U13559 (N_13559,N_12000,N_12103);
and U13560 (N_13560,N_12321,N_12195);
nor U13561 (N_13561,N_12572,N_12435);
nor U13562 (N_13562,N_12505,N_12020);
nor U13563 (N_13563,N_12673,N_12889);
xor U13564 (N_13564,N_12371,N_12087);
and U13565 (N_13565,N_12472,N_12473);
nor U13566 (N_13566,N_12845,N_12876);
nand U13567 (N_13567,N_12260,N_12802);
xnor U13568 (N_13568,N_12244,N_12999);
nor U13569 (N_13569,N_12102,N_12785);
nor U13570 (N_13570,N_12879,N_12828);
xnor U13571 (N_13571,N_12096,N_12860);
xor U13572 (N_13572,N_12842,N_12797);
nor U13573 (N_13573,N_12610,N_12592);
nor U13574 (N_13574,N_12455,N_12641);
or U13575 (N_13575,N_12832,N_12871);
nor U13576 (N_13576,N_12853,N_12115);
nor U13577 (N_13577,N_12102,N_12463);
nor U13578 (N_13578,N_12852,N_12676);
and U13579 (N_13579,N_12446,N_12895);
nand U13580 (N_13580,N_12408,N_12613);
nor U13581 (N_13581,N_12239,N_12880);
nor U13582 (N_13582,N_12543,N_12041);
xor U13583 (N_13583,N_12393,N_12659);
or U13584 (N_13584,N_12839,N_12798);
and U13585 (N_13585,N_12723,N_12554);
nor U13586 (N_13586,N_12494,N_12884);
or U13587 (N_13587,N_12087,N_12578);
or U13588 (N_13588,N_12629,N_12444);
or U13589 (N_13589,N_12273,N_12658);
xnor U13590 (N_13590,N_12203,N_12693);
and U13591 (N_13591,N_12091,N_12997);
nand U13592 (N_13592,N_12773,N_12328);
nand U13593 (N_13593,N_12026,N_12731);
and U13594 (N_13594,N_12179,N_12404);
xnor U13595 (N_13595,N_12488,N_12776);
nand U13596 (N_13596,N_12165,N_12094);
nor U13597 (N_13597,N_12064,N_12351);
and U13598 (N_13598,N_12725,N_12108);
xor U13599 (N_13599,N_12325,N_12125);
and U13600 (N_13600,N_12784,N_12372);
or U13601 (N_13601,N_12676,N_12130);
or U13602 (N_13602,N_12627,N_12882);
xnor U13603 (N_13603,N_12055,N_12564);
nand U13604 (N_13604,N_12096,N_12275);
xnor U13605 (N_13605,N_12074,N_12300);
xor U13606 (N_13606,N_12588,N_12333);
or U13607 (N_13607,N_12423,N_12451);
or U13608 (N_13608,N_12318,N_12975);
nand U13609 (N_13609,N_12657,N_12522);
or U13610 (N_13610,N_12413,N_12090);
and U13611 (N_13611,N_12667,N_12063);
and U13612 (N_13612,N_12203,N_12602);
nor U13613 (N_13613,N_12543,N_12144);
nand U13614 (N_13614,N_12426,N_12240);
or U13615 (N_13615,N_12551,N_12568);
nand U13616 (N_13616,N_12731,N_12734);
xnor U13617 (N_13617,N_12902,N_12006);
nand U13618 (N_13618,N_12140,N_12290);
and U13619 (N_13619,N_12625,N_12316);
nand U13620 (N_13620,N_12817,N_12135);
and U13621 (N_13621,N_12157,N_12140);
or U13622 (N_13622,N_12847,N_12684);
or U13623 (N_13623,N_12320,N_12530);
or U13624 (N_13624,N_12169,N_12857);
and U13625 (N_13625,N_12346,N_12161);
nor U13626 (N_13626,N_12896,N_12687);
and U13627 (N_13627,N_12874,N_12004);
nor U13628 (N_13628,N_12073,N_12380);
nand U13629 (N_13629,N_12858,N_12990);
xnor U13630 (N_13630,N_12776,N_12516);
nand U13631 (N_13631,N_12337,N_12067);
nor U13632 (N_13632,N_12766,N_12028);
nand U13633 (N_13633,N_12233,N_12057);
and U13634 (N_13634,N_12576,N_12510);
nor U13635 (N_13635,N_12197,N_12187);
nor U13636 (N_13636,N_12477,N_12614);
nand U13637 (N_13637,N_12143,N_12624);
nor U13638 (N_13638,N_12988,N_12366);
and U13639 (N_13639,N_12295,N_12019);
nand U13640 (N_13640,N_12139,N_12851);
nor U13641 (N_13641,N_12533,N_12094);
nand U13642 (N_13642,N_12706,N_12076);
and U13643 (N_13643,N_12549,N_12446);
and U13644 (N_13644,N_12276,N_12852);
nor U13645 (N_13645,N_12835,N_12545);
nor U13646 (N_13646,N_12362,N_12903);
nand U13647 (N_13647,N_12967,N_12906);
nor U13648 (N_13648,N_12692,N_12068);
xnor U13649 (N_13649,N_12994,N_12900);
nor U13650 (N_13650,N_12374,N_12369);
nor U13651 (N_13651,N_12696,N_12027);
and U13652 (N_13652,N_12464,N_12832);
nor U13653 (N_13653,N_12730,N_12922);
nand U13654 (N_13654,N_12019,N_12626);
xor U13655 (N_13655,N_12846,N_12774);
and U13656 (N_13656,N_12743,N_12871);
and U13657 (N_13657,N_12411,N_12738);
and U13658 (N_13658,N_12334,N_12997);
and U13659 (N_13659,N_12124,N_12689);
or U13660 (N_13660,N_12320,N_12621);
nor U13661 (N_13661,N_12599,N_12414);
nor U13662 (N_13662,N_12327,N_12787);
nor U13663 (N_13663,N_12355,N_12190);
nand U13664 (N_13664,N_12438,N_12834);
or U13665 (N_13665,N_12401,N_12630);
xor U13666 (N_13666,N_12645,N_12443);
nand U13667 (N_13667,N_12331,N_12479);
or U13668 (N_13668,N_12657,N_12541);
xor U13669 (N_13669,N_12168,N_12833);
and U13670 (N_13670,N_12445,N_12121);
nor U13671 (N_13671,N_12017,N_12621);
xor U13672 (N_13672,N_12302,N_12300);
or U13673 (N_13673,N_12136,N_12862);
and U13674 (N_13674,N_12360,N_12257);
nand U13675 (N_13675,N_12703,N_12760);
xor U13676 (N_13676,N_12467,N_12241);
or U13677 (N_13677,N_12178,N_12213);
nand U13678 (N_13678,N_12426,N_12816);
or U13679 (N_13679,N_12676,N_12762);
or U13680 (N_13680,N_12508,N_12106);
nand U13681 (N_13681,N_12582,N_12256);
xor U13682 (N_13682,N_12005,N_12586);
nor U13683 (N_13683,N_12979,N_12648);
xnor U13684 (N_13684,N_12358,N_12157);
xor U13685 (N_13685,N_12739,N_12508);
xor U13686 (N_13686,N_12777,N_12573);
or U13687 (N_13687,N_12850,N_12520);
or U13688 (N_13688,N_12162,N_12866);
and U13689 (N_13689,N_12468,N_12381);
and U13690 (N_13690,N_12757,N_12911);
nor U13691 (N_13691,N_12870,N_12559);
or U13692 (N_13692,N_12648,N_12530);
xnor U13693 (N_13693,N_12380,N_12422);
and U13694 (N_13694,N_12425,N_12758);
nor U13695 (N_13695,N_12109,N_12131);
and U13696 (N_13696,N_12578,N_12016);
and U13697 (N_13697,N_12702,N_12830);
or U13698 (N_13698,N_12129,N_12534);
or U13699 (N_13699,N_12223,N_12452);
nor U13700 (N_13700,N_12334,N_12284);
nor U13701 (N_13701,N_12812,N_12062);
xnor U13702 (N_13702,N_12509,N_12026);
nand U13703 (N_13703,N_12795,N_12717);
nand U13704 (N_13704,N_12834,N_12133);
xor U13705 (N_13705,N_12689,N_12096);
nand U13706 (N_13706,N_12943,N_12311);
xnor U13707 (N_13707,N_12568,N_12023);
nor U13708 (N_13708,N_12026,N_12558);
or U13709 (N_13709,N_12281,N_12826);
or U13710 (N_13710,N_12085,N_12666);
and U13711 (N_13711,N_12200,N_12653);
nand U13712 (N_13712,N_12624,N_12025);
nand U13713 (N_13713,N_12194,N_12499);
nand U13714 (N_13714,N_12937,N_12807);
xnor U13715 (N_13715,N_12725,N_12652);
or U13716 (N_13716,N_12746,N_12666);
or U13717 (N_13717,N_12726,N_12290);
or U13718 (N_13718,N_12393,N_12163);
xnor U13719 (N_13719,N_12079,N_12939);
xor U13720 (N_13720,N_12797,N_12159);
xor U13721 (N_13721,N_12648,N_12379);
xnor U13722 (N_13722,N_12402,N_12577);
or U13723 (N_13723,N_12876,N_12145);
xor U13724 (N_13724,N_12752,N_12723);
nor U13725 (N_13725,N_12858,N_12399);
or U13726 (N_13726,N_12734,N_12305);
nand U13727 (N_13727,N_12757,N_12172);
and U13728 (N_13728,N_12679,N_12955);
and U13729 (N_13729,N_12813,N_12264);
or U13730 (N_13730,N_12431,N_12539);
nand U13731 (N_13731,N_12821,N_12222);
or U13732 (N_13732,N_12885,N_12018);
or U13733 (N_13733,N_12825,N_12550);
or U13734 (N_13734,N_12959,N_12395);
xnor U13735 (N_13735,N_12250,N_12229);
and U13736 (N_13736,N_12541,N_12609);
nand U13737 (N_13737,N_12405,N_12314);
and U13738 (N_13738,N_12930,N_12188);
xnor U13739 (N_13739,N_12223,N_12726);
xnor U13740 (N_13740,N_12616,N_12153);
and U13741 (N_13741,N_12273,N_12833);
nand U13742 (N_13742,N_12900,N_12576);
or U13743 (N_13743,N_12275,N_12810);
xor U13744 (N_13744,N_12757,N_12046);
nor U13745 (N_13745,N_12143,N_12958);
xor U13746 (N_13746,N_12478,N_12711);
xor U13747 (N_13747,N_12671,N_12632);
and U13748 (N_13748,N_12633,N_12966);
and U13749 (N_13749,N_12658,N_12530);
nor U13750 (N_13750,N_12897,N_12878);
nor U13751 (N_13751,N_12624,N_12645);
and U13752 (N_13752,N_12081,N_12971);
nand U13753 (N_13753,N_12329,N_12802);
xnor U13754 (N_13754,N_12795,N_12827);
or U13755 (N_13755,N_12790,N_12912);
or U13756 (N_13756,N_12612,N_12665);
nand U13757 (N_13757,N_12626,N_12642);
xor U13758 (N_13758,N_12086,N_12921);
and U13759 (N_13759,N_12070,N_12815);
and U13760 (N_13760,N_12882,N_12568);
and U13761 (N_13761,N_12438,N_12051);
or U13762 (N_13762,N_12385,N_12847);
xnor U13763 (N_13763,N_12026,N_12822);
and U13764 (N_13764,N_12500,N_12229);
nor U13765 (N_13765,N_12891,N_12417);
xnor U13766 (N_13766,N_12671,N_12388);
xnor U13767 (N_13767,N_12878,N_12019);
and U13768 (N_13768,N_12043,N_12169);
nor U13769 (N_13769,N_12023,N_12258);
or U13770 (N_13770,N_12875,N_12162);
nor U13771 (N_13771,N_12085,N_12275);
xnor U13772 (N_13772,N_12656,N_12832);
and U13773 (N_13773,N_12932,N_12671);
and U13774 (N_13774,N_12521,N_12974);
nand U13775 (N_13775,N_12179,N_12422);
nor U13776 (N_13776,N_12630,N_12496);
nand U13777 (N_13777,N_12682,N_12410);
and U13778 (N_13778,N_12451,N_12736);
nand U13779 (N_13779,N_12425,N_12299);
or U13780 (N_13780,N_12131,N_12425);
nor U13781 (N_13781,N_12585,N_12995);
xor U13782 (N_13782,N_12382,N_12060);
or U13783 (N_13783,N_12435,N_12381);
xor U13784 (N_13784,N_12710,N_12060);
nand U13785 (N_13785,N_12608,N_12207);
nor U13786 (N_13786,N_12125,N_12625);
nor U13787 (N_13787,N_12956,N_12631);
nor U13788 (N_13788,N_12381,N_12168);
nand U13789 (N_13789,N_12197,N_12276);
or U13790 (N_13790,N_12759,N_12156);
and U13791 (N_13791,N_12089,N_12483);
nand U13792 (N_13792,N_12356,N_12898);
and U13793 (N_13793,N_12285,N_12290);
nor U13794 (N_13794,N_12827,N_12069);
nor U13795 (N_13795,N_12440,N_12694);
xor U13796 (N_13796,N_12217,N_12215);
nor U13797 (N_13797,N_12875,N_12920);
or U13798 (N_13798,N_12550,N_12212);
nor U13799 (N_13799,N_12631,N_12529);
or U13800 (N_13800,N_12038,N_12523);
nand U13801 (N_13801,N_12477,N_12032);
nor U13802 (N_13802,N_12308,N_12613);
or U13803 (N_13803,N_12269,N_12689);
and U13804 (N_13804,N_12567,N_12316);
nor U13805 (N_13805,N_12800,N_12691);
nand U13806 (N_13806,N_12948,N_12227);
xnor U13807 (N_13807,N_12250,N_12829);
or U13808 (N_13808,N_12100,N_12269);
xor U13809 (N_13809,N_12139,N_12953);
nor U13810 (N_13810,N_12349,N_12957);
xnor U13811 (N_13811,N_12970,N_12406);
nand U13812 (N_13812,N_12653,N_12609);
and U13813 (N_13813,N_12399,N_12595);
nand U13814 (N_13814,N_12762,N_12304);
and U13815 (N_13815,N_12230,N_12984);
and U13816 (N_13816,N_12778,N_12083);
nand U13817 (N_13817,N_12273,N_12035);
xor U13818 (N_13818,N_12506,N_12895);
nor U13819 (N_13819,N_12245,N_12065);
xor U13820 (N_13820,N_12374,N_12519);
or U13821 (N_13821,N_12905,N_12371);
xor U13822 (N_13822,N_12066,N_12250);
nor U13823 (N_13823,N_12480,N_12187);
or U13824 (N_13824,N_12673,N_12402);
nand U13825 (N_13825,N_12786,N_12189);
nor U13826 (N_13826,N_12132,N_12568);
or U13827 (N_13827,N_12825,N_12271);
xnor U13828 (N_13828,N_12636,N_12230);
nor U13829 (N_13829,N_12504,N_12793);
nand U13830 (N_13830,N_12671,N_12039);
nor U13831 (N_13831,N_12551,N_12268);
xor U13832 (N_13832,N_12429,N_12702);
nor U13833 (N_13833,N_12620,N_12845);
or U13834 (N_13834,N_12897,N_12377);
and U13835 (N_13835,N_12124,N_12174);
nor U13836 (N_13836,N_12163,N_12597);
and U13837 (N_13837,N_12122,N_12881);
nand U13838 (N_13838,N_12186,N_12442);
nand U13839 (N_13839,N_12189,N_12515);
xnor U13840 (N_13840,N_12430,N_12348);
and U13841 (N_13841,N_12591,N_12576);
and U13842 (N_13842,N_12952,N_12091);
xor U13843 (N_13843,N_12052,N_12648);
or U13844 (N_13844,N_12983,N_12246);
or U13845 (N_13845,N_12924,N_12384);
or U13846 (N_13846,N_12375,N_12266);
or U13847 (N_13847,N_12803,N_12889);
xnor U13848 (N_13848,N_12487,N_12877);
nand U13849 (N_13849,N_12602,N_12776);
nor U13850 (N_13850,N_12099,N_12787);
nor U13851 (N_13851,N_12941,N_12630);
or U13852 (N_13852,N_12573,N_12634);
xnor U13853 (N_13853,N_12932,N_12043);
xnor U13854 (N_13854,N_12225,N_12383);
and U13855 (N_13855,N_12320,N_12797);
nor U13856 (N_13856,N_12967,N_12679);
or U13857 (N_13857,N_12461,N_12959);
nand U13858 (N_13858,N_12089,N_12824);
xnor U13859 (N_13859,N_12736,N_12095);
nand U13860 (N_13860,N_12196,N_12640);
nor U13861 (N_13861,N_12591,N_12731);
or U13862 (N_13862,N_12618,N_12601);
nor U13863 (N_13863,N_12309,N_12888);
xor U13864 (N_13864,N_12283,N_12361);
nor U13865 (N_13865,N_12344,N_12231);
nor U13866 (N_13866,N_12320,N_12930);
and U13867 (N_13867,N_12310,N_12566);
nor U13868 (N_13868,N_12948,N_12212);
and U13869 (N_13869,N_12506,N_12037);
nand U13870 (N_13870,N_12052,N_12612);
nand U13871 (N_13871,N_12741,N_12231);
nand U13872 (N_13872,N_12355,N_12314);
or U13873 (N_13873,N_12002,N_12085);
nand U13874 (N_13874,N_12260,N_12071);
xor U13875 (N_13875,N_12938,N_12148);
or U13876 (N_13876,N_12015,N_12362);
xnor U13877 (N_13877,N_12586,N_12591);
nor U13878 (N_13878,N_12410,N_12261);
nand U13879 (N_13879,N_12182,N_12852);
or U13880 (N_13880,N_12799,N_12096);
nand U13881 (N_13881,N_12899,N_12902);
xor U13882 (N_13882,N_12829,N_12817);
xnor U13883 (N_13883,N_12676,N_12164);
and U13884 (N_13884,N_12117,N_12068);
or U13885 (N_13885,N_12182,N_12320);
nor U13886 (N_13886,N_12505,N_12498);
xnor U13887 (N_13887,N_12792,N_12500);
or U13888 (N_13888,N_12788,N_12013);
nor U13889 (N_13889,N_12137,N_12280);
nand U13890 (N_13890,N_12582,N_12818);
and U13891 (N_13891,N_12161,N_12252);
nor U13892 (N_13892,N_12511,N_12400);
nor U13893 (N_13893,N_12101,N_12631);
nor U13894 (N_13894,N_12982,N_12674);
nor U13895 (N_13895,N_12961,N_12140);
nor U13896 (N_13896,N_12135,N_12476);
xnor U13897 (N_13897,N_12434,N_12374);
nor U13898 (N_13898,N_12092,N_12504);
nand U13899 (N_13899,N_12631,N_12711);
xor U13900 (N_13900,N_12010,N_12091);
nor U13901 (N_13901,N_12090,N_12599);
or U13902 (N_13902,N_12921,N_12864);
and U13903 (N_13903,N_12663,N_12118);
or U13904 (N_13904,N_12808,N_12991);
or U13905 (N_13905,N_12055,N_12316);
xor U13906 (N_13906,N_12905,N_12472);
nor U13907 (N_13907,N_12857,N_12717);
nor U13908 (N_13908,N_12211,N_12405);
xnor U13909 (N_13909,N_12121,N_12296);
and U13910 (N_13910,N_12152,N_12445);
and U13911 (N_13911,N_12671,N_12436);
nor U13912 (N_13912,N_12119,N_12696);
nand U13913 (N_13913,N_12844,N_12363);
xnor U13914 (N_13914,N_12887,N_12581);
or U13915 (N_13915,N_12953,N_12271);
nand U13916 (N_13916,N_12711,N_12175);
and U13917 (N_13917,N_12348,N_12262);
nor U13918 (N_13918,N_12190,N_12146);
nand U13919 (N_13919,N_12061,N_12906);
nor U13920 (N_13920,N_12016,N_12417);
xnor U13921 (N_13921,N_12718,N_12304);
nor U13922 (N_13922,N_12428,N_12697);
and U13923 (N_13923,N_12228,N_12645);
or U13924 (N_13924,N_12991,N_12010);
xnor U13925 (N_13925,N_12851,N_12039);
or U13926 (N_13926,N_12705,N_12303);
or U13927 (N_13927,N_12857,N_12146);
and U13928 (N_13928,N_12568,N_12843);
or U13929 (N_13929,N_12505,N_12074);
or U13930 (N_13930,N_12610,N_12380);
or U13931 (N_13931,N_12410,N_12783);
nor U13932 (N_13932,N_12061,N_12131);
nor U13933 (N_13933,N_12741,N_12008);
and U13934 (N_13934,N_12784,N_12366);
nand U13935 (N_13935,N_12307,N_12762);
xor U13936 (N_13936,N_12327,N_12208);
or U13937 (N_13937,N_12554,N_12853);
xnor U13938 (N_13938,N_12327,N_12369);
nor U13939 (N_13939,N_12321,N_12329);
xor U13940 (N_13940,N_12206,N_12311);
or U13941 (N_13941,N_12660,N_12802);
nor U13942 (N_13942,N_12978,N_12101);
nand U13943 (N_13943,N_12777,N_12584);
or U13944 (N_13944,N_12648,N_12936);
nand U13945 (N_13945,N_12165,N_12846);
and U13946 (N_13946,N_12804,N_12737);
nand U13947 (N_13947,N_12293,N_12699);
nor U13948 (N_13948,N_12884,N_12163);
or U13949 (N_13949,N_12533,N_12910);
nor U13950 (N_13950,N_12692,N_12561);
nor U13951 (N_13951,N_12061,N_12290);
and U13952 (N_13952,N_12652,N_12320);
or U13953 (N_13953,N_12645,N_12225);
and U13954 (N_13954,N_12188,N_12604);
nand U13955 (N_13955,N_12283,N_12312);
nor U13956 (N_13956,N_12878,N_12519);
nor U13957 (N_13957,N_12346,N_12654);
and U13958 (N_13958,N_12331,N_12581);
nand U13959 (N_13959,N_12458,N_12664);
nor U13960 (N_13960,N_12739,N_12053);
or U13961 (N_13961,N_12140,N_12169);
xor U13962 (N_13962,N_12343,N_12876);
nand U13963 (N_13963,N_12473,N_12664);
xnor U13964 (N_13964,N_12351,N_12245);
xor U13965 (N_13965,N_12945,N_12332);
nor U13966 (N_13966,N_12886,N_12244);
xor U13967 (N_13967,N_12263,N_12345);
and U13968 (N_13968,N_12631,N_12745);
nand U13969 (N_13969,N_12298,N_12036);
xnor U13970 (N_13970,N_12018,N_12101);
and U13971 (N_13971,N_12319,N_12661);
and U13972 (N_13972,N_12872,N_12050);
and U13973 (N_13973,N_12975,N_12420);
nand U13974 (N_13974,N_12633,N_12338);
and U13975 (N_13975,N_12389,N_12960);
or U13976 (N_13976,N_12157,N_12390);
and U13977 (N_13977,N_12562,N_12933);
xnor U13978 (N_13978,N_12372,N_12243);
nand U13979 (N_13979,N_12375,N_12129);
nor U13980 (N_13980,N_12809,N_12176);
xor U13981 (N_13981,N_12623,N_12111);
xor U13982 (N_13982,N_12239,N_12108);
nor U13983 (N_13983,N_12587,N_12439);
xnor U13984 (N_13984,N_12363,N_12184);
and U13985 (N_13985,N_12290,N_12659);
or U13986 (N_13986,N_12309,N_12214);
and U13987 (N_13987,N_12174,N_12554);
xnor U13988 (N_13988,N_12419,N_12897);
and U13989 (N_13989,N_12926,N_12174);
or U13990 (N_13990,N_12705,N_12958);
and U13991 (N_13991,N_12570,N_12460);
nand U13992 (N_13992,N_12320,N_12158);
or U13993 (N_13993,N_12507,N_12083);
or U13994 (N_13994,N_12136,N_12045);
xnor U13995 (N_13995,N_12941,N_12690);
and U13996 (N_13996,N_12292,N_12817);
and U13997 (N_13997,N_12422,N_12396);
and U13998 (N_13998,N_12010,N_12463);
nand U13999 (N_13999,N_12490,N_12550);
xor U14000 (N_14000,N_13935,N_13765);
and U14001 (N_14001,N_13952,N_13597);
nor U14002 (N_14002,N_13556,N_13640);
nor U14003 (N_14003,N_13668,N_13087);
xnor U14004 (N_14004,N_13543,N_13938);
nand U14005 (N_14005,N_13633,N_13139);
nand U14006 (N_14006,N_13726,N_13253);
xnor U14007 (N_14007,N_13538,N_13666);
nor U14008 (N_14008,N_13697,N_13770);
or U14009 (N_14009,N_13573,N_13165);
nor U14010 (N_14010,N_13810,N_13424);
or U14011 (N_14011,N_13958,N_13558);
nor U14012 (N_14012,N_13653,N_13654);
nor U14013 (N_14013,N_13117,N_13960);
nor U14014 (N_14014,N_13414,N_13379);
or U14015 (N_14015,N_13874,N_13814);
nand U14016 (N_14016,N_13360,N_13883);
nor U14017 (N_14017,N_13127,N_13063);
nor U14018 (N_14018,N_13079,N_13122);
nand U14019 (N_14019,N_13428,N_13769);
or U14020 (N_14020,N_13111,N_13094);
or U14021 (N_14021,N_13818,N_13483);
or U14022 (N_14022,N_13959,N_13083);
nand U14023 (N_14023,N_13477,N_13189);
nand U14024 (N_14024,N_13491,N_13452);
nor U14025 (N_14025,N_13157,N_13010);
nor U14026 (N_14026,N_13036,N_13455);
xnor U14027 (N_14027,N_13182,N_13578);
or U14028 (N_14028,N_13449,N_13739);
or U14029 (N_14029,N_13511,N_13313);
nand U14030 (N_14030,N_13329,N_13848);
xnor U14031 (N_14031,N_13762,N_13011);
or U14032 (N_14032,N_13126,N_13112);
xnor U14033 (N_14033,N_13922,N_13432);
and U14034 (N_14034,N_13445,N_13199);
nand U14035 (N_14035,N_13598,N_13893);
or U14036 (N_14036,N_13289,N_13949);
nor U14037 (N_14037,N_13916,N_13977);
or U14038 (N_14038,N_13942,N_13048);
xor U14039 (N_14039,N_13995,N_13150);
and U14040 (N_14040,N_13110,N_13172);
nand U14041 (N_14041,N_13179,N_13557);
nand U14042 (N_14042,N_13567,N_13847);
nand U14043 (N_14043,N_13105,N_13368);
xor U14044 (N_14044,N_13377,N_13203);
or U14045 (N_14045,N_13616,N_13669);
and U14046 (N_14046,N_13019,N_13525);
and U14047 (N_14047,N_13894,N_13453);
nor U14048 (N_14048,N_13131,N_13324);
or U14049 (N_14049,N_13887,N_13056);
nand U14050 (N_14050,N_13718,N_13576);
and U14051 (N_14051,N_13146,N_13061);
and U14052 (N_14052,N_13185,N_13068);
nand U14053 (N_14053,N_13343,N_13008);
nor U14054 (N_14054,N_13706,N_13863);
or U14055 (N_14055,N_13420,N_13430);
or U14056 (N_14056,N_13659,N_13918);
or U14057 (N_14057,N_13541,N_13690);
nand U14058 (N_14058,N_13717,N_13701);
nand U14059 (N_14059,N_13806,N_13415);
nand U14060 (N_14060,N_13362,N_13018);
nand U14061 (N_14061,N_13702,N_13378);
and U14062 (N_14062,N_13221,N_13943);
and U14063 (N_14063,N_13171,N_13373);
nand U14064 (N_14064,N_13064,N_13475);
or U14065 (N_14065,N_13840,N_13315);
xnor U14066 (N_14066,N_13191,N_13035);
and U14067 (N_14067,N_13907,N_13745);
nor U14068 (N_14068,N_13497,N_13988);
and U14069 (N_14069,N_13211,N_13071);
or U14070 (N_14070,N_13369,N_13707);
or U14071 (N_14071,N_13159,N_13239);
nor U14072 (N_14072,N_13996,N_13429);
or U14073 (N_14073,N_13046,N_13851);
or U14074 (N_14074,N_13344,N_13820);
nand U14075 (N_14075,N_13651,N_13976);
and U14076 (N_14076,N_13534,N_13506);
or U14077 (N_14077,N_13784,N_13248);
xor U14078 (N_14078,N_13961,N_13200);
and U14079 (N_14079,N_13622,N_13412);
or U14080 (N_14080,N_13735,N_13861);
nor U14081 (N_14081,N_13882,N_13438);
and U14082 (N_14082,N_13299,N_13778);
or U14083 (N_14083,N_13895,N_13613);
nand U14084 (N_14084,N_13004,N_13711);
xnor U14085 (N_14085,N_13007,N_13852);
xnor U14086 (N_14086,N_13338,N_13950);
and U14087 (N_14087,N_13891,N_13107);
nand U14088 (N_14088,N_13715,N_13471);
nor U14089 (N_14089,N_13496,N_13650);
xor U14090 (N_14090,N_13716,N_13294);
and U14091 (N_14091,N_13772,N_13410);
or U14092 (N_14092,N_13161,N_13969);
nand U14093 (N_14093,N_13017,N_13662);
nor U14094 (N_14094,N_13067,N_13908);
xor U14095 (N_14095,N_13621,N_13151);
nand U14096 (N_14096,N_13584,N_13099);
or U14097 (N_14097,N_13560,N_13407);
nor U14098 (N_14098,N_13825,N_13572);
nand U14099 (N_14099,N_13508,N_13130);
or U14100 (N_14100,N_13740,N_13624);
nor U14101 (N_14101,N_13078,N_13678);
nor U14102 (N_14102,N_13437,N_13886);
or U14103 (N_14103,N_13404,N_13986);
and U14104 (N_14104,N_13054,N_13266);
or U14105 (N_14105,N_13476,N_13354);
nand U14106 (N_14106,N_13877,N_13837);
nor U14107 (N_14107,N_13785,N_13252);
or U14108 (N_14108,N_13489,N_13775);
and U14109 (N_14109,N_13897,N_13192);
nand U14110 (N_14110,N_13644,N_13569);
nand U14111 (N_14111,N_13355,N_13325);
xor U14112 (N_14112,N_13839,N_13804);
nand U14113 (N_14113,N_13792,N_13413);
nand U14114 (N_14114,N_13904,N_13311);
and U14115 (N_14115,N_13675,N_13815);
and U14116 (N_14116,N_13272,N_13521);
and U14117 (N_14117,N_13781,N_13963);
and U14118 (N_14118,N_13967,N_13198);
xor U14119 (N_14119,N_13532,N_13244);
xor U14120 (N_14120,N_13230,N_13892);
xnor U14121 (N_14121,N_13218,N_13256);
or U14122 (N_14122,N_13583,N_13389);
and U14123 (N_14123,N_13579,N_13507);
and U14124 (N_14124,N_13733,N_13615);
nand U14125 (N_14125,N_13206,N_13856);
nand U14126 (N_14126,N_13411,N_13260);
or U14127 (N_14127,N_13780,N_13732);
or U14128 (N_14128,N_13392,N_13997);
or U14129 (N_14129,N_13454,N_13059);
or U14130 (N_14130,N_13630,N_13381);
xor U14131 (N_14131,N_13065,N_13441);
nor U14132 (N_14132,N_13636,N_13764);
and U14133 (N_14133,N_13610,N_13082);
nor U14134 (N_14134,N_13481,N_13990);
nand U14135 (N_14135,N_13470,N_13393);
nor U14136 (N_14136,N_13293,N_13186);
or U14137 (N_14137,N_13822,N_13366);
and U14138 (N_14138,N_13915,N_13562);
nor U14139 (N_14139,N_13872,N_13013);
and U14140 (N_14140,N_13912,N_13955);
nand U14141 (N_14141,N_13208,N_13401);
and U14142 (N_14142,N_13603,N_13727);
or U14143 (N_14143,N_13468,N_13279);
or U14144 (N_14144,N_13217,N_13081);
nand U14145 (N_14145,N_13479,N_13375);
and U14146 (N_14146,N_13276,N_13667);
nand U14147 (N_14147,N_13403,N_13228);
nand U14148 (N_14148,N_13526,N_13298);
nand U14149 (N_14149,N_13318,N_13542);
and U14150 (N_14150,N_13994,N_13210);
nor U14151 (N_14151,N_13509,N_13209);
or U14152 (N_14152,N_13529,N_13442);
nand U14153 (N_14153,N_13634,N_13869);
nand U14154 (N_14154,N_13234,N_13531);
nand U14155 (N_14155,N_13728,N_13871);
nand U14156 (N_14156,N_13484,N_13750);
xnor U14157 (N_14157,N_13451,N_13749);
or U14158 (N_14158,N_13805,N_13027);
nand U14159 (N_14159,N_13844,N_13359);
nor U14160 (N_14160,N_13271,N_13015);
and U14161 (N_14161,N_13282,N_13353);
and U14162 (N_14162,N_13328,N_13547);
xor U14163 (N_14163,N_13190,N_13098);
and U14164 (N_14164,N_13889,N_13487);
or U14165 (N_14165,N_13400,N_13671);
or U14166 (N_14166,N_13817,N_13632);
nand U14167 (N_14167,N_13236,N_13371);
nor U14168 (N_14168,N_13333,N_13841);
nand U14169 (N_14169,N_13828,N_13267);
xnor U14170 (N_14170,N_13979,N_13149);
and U14171 (N_14171,N_13884,N_13187);
nand U14172 (N_14172,N_13292,N_13406);
nand U14173 (N_14173,N_13050,N_13347);
nand U14174 (N_14174,N_13195,N_13283);
and U14175 (N_14175,N_13763,N_13639);
or U14176 (N_14176,N_13647,N_13215);
nand U14177 (N_14177,N_13029,N_13743);
or U14178 (N_14178,N_13188,N_13327);
and U14179 (N_14179,N_13040,N_13049);
or U14180 (N_14180,N_13306,N_13431);
nor U14181 (N_14181,N_13937,N_13168);
nor U14182 (N_14182,N_13748,N_13480);
or U14183 (N_14183,N_13034,N_13114);
xor U14184 (N_14184,N_13356,N_13962);
nor U14185 (N_14185,N_13258,N_13080);
nand U14186 (N_14186,N_13791,N_13753);
or U14187 (N_14187,N_13223,N_13024);
xnor U14188 (N_14188,N_13596,N_13277);
and U14189 (N_14189,N_13364,N_13593);
nand U14190 (N_14190,N_13794,N_13383);
and U14191 (N_14191,N_13801,N_13559);
or U14192 (N_14192,N_13473,N_13308);
nand U14193 (N_14193,N_13535,N_13694);
and U14194 (N_14194,N_13077,N_13025);
or U14195 (N_14195,N_13953,N_13231);
and U14196 (N_14196,N_13340,N_13896);
xnor U14197 (N_14197,N_13570,N_13954);
nand U14198 (N_14198,N_13900,N_13873);
xnor U14199 (N_14199,N_13586,N_13095);
nand U14200 (N_14200,N_13088,N_13365);
and U14201 (N_14201,N_13688,N_13561);
nand U14202 (N_14202,N_13838,N_13734);
xnor U14203 (N_14203,N_13700,N_13133);
nand U14204 (N_14204,N_13564,N_13867);
or U14205 (N_14205,N_13673,N_13462);
nor U14206 (N_14206,N_13574,N_13929);
nand U14207 (N_14207,N_13776,N_13044);
and U14208 (N_14208,N_13227,N_13280);
xor U14209 (N_14209,N_13156,N_13175);
or U14210 (N_14210,N_13917,N_13782);
nand U14211 (N_14211,N_13670,N_13555);
nor U14212 (N_14212,N_13720,N_13257);
nand U14213 (N_14213,N_13488,N_13695);
nor U14214 (N_14214,N_13522,N_13229);
or U14215 (N_14215,N_13605,N_13545);
nor U14216 (N_14216,N_13513,N_13809);
and U14217 (N_14217,N_13826,N_13472);
nand U14218 (N_14218,N_13971,N_13419);
xor U14219 (N_14219,N_13663,N_13899);
or U14220 (N_14220,N_13719,N_13337);
and U14221 (N_14221,N_13273,N_13802);
nor U14222 (N_14222,N_13222,N_13070);
nand U14223 (N_14223,N_13982,N_13577);
nand U14224 (N_14224,N_13879,N_13803);
xor U14225 (N_14225,N_13320,N_13296);
or U14226 (N_14226,N_13425,N_13224);
and U14227 (N_14227,N_13020,N_13197);
or U14228 (N_14228,N_13787,N_13363);
or U14229 (N_14229,N_13274,N_13387);
xnor U14230 (N_14230,N_13269,N_13384);
and U14231 (N_14231,N_13498,N_13262);
nand U14232 (N_14232,N_13124,N_13587);
nand U14233 (N_14233,N_13641,N_13786);
and U14234 (N_14234,N_13652,N_13264);
nor U14235 (N_14235,N_13858,N_13875);
and U14236 (N_14236,N_13037,N_13946);
or U14237 (N_14237,N_13842,N_13499);
nand U14238 (N_14238,N_13242,N_13618);
nand U14239 (N_14239,N_13495,N_13225);
or U14240 (N_14240,N_13309,N_13478);
xor U14241 (N_14241,N_13713,N_13297);
and U14242 (N_14242,N_13811,N_13000);
nor U14243 (N_14243,N_13003,N_13617);
and U14244 (N_14244,N_13287,N_13450);
xor U14245 (N_14245,N_13902,N_13709);
and U14246 (N_14246,N_13370,N_13703);
nand U14247 (N_14247,N_13170,N_13736);
xnor U14248 (N_14248,N_13395,N_13866);
nand U14249 (N_14249,N_13464,N_13947);
nor U14250 (N_14250,N_13723,N_13014);
xnor U14251 (N_14251,N_13235,N_13604);
nand U14252 (N_14252,N_13756,N_13196);
nor U14253 (N_14253,N_13909,N_13850);
xor U14254 (N_14254,N_13456,N_13101);
nand U14255 (N_14255,N_13458,N_13626);
and U14256 (N_14256,N_13463,N_13397);
and U14257 (N_14257,N_13600,N_13086);
and U14258 (N_14258,N_13933,N_13345);
xor U14259 (N_14259,N_13581,N_13357);
nor U14260 (N_14260,N_13968,N_13092);
nand U14261 (N_14261,N_13349,N_13254);
and U14262 (N_14262,N_13518,N_13849);
nor U14263 (N_14263,N_13699,N_13819);
or U14264 (N_14264,N_13629,N_13993);
or U14265 (N_14265,N_13989,N_13399);
and U14266 (N_14266,N_13342,N_13539);
xnor U14267 (N_14267,N_13864,N_13268);
or U14268 (N_14268,N_13402,N_13358);
nor U14269 (N_14269,N_13291,N_13853);
and U14270 (N_14270,N_13436,N_13164);
or U14271 (N_14271,N_13985,N_13301);
and U14272 (N_14272,N_13813,N_13623);
xor U14273 (N_14273,N_13683,N_13351);
and U14274 (N_14274,N_13664,N_13661);
or U14275 (N_14275,N_13777,N_13625);
and U14276 (N_14276,N_13552,N_13265);
or U14277 (N_14277,N_13691,N_13631);
or U14278 (N_14278,N_13136,N_13113);
xnor U14279 (N_14279,N_13612,N_13466);
or U14280 (N_14280,N_13143,N_13154);
nor U14281 (N_14281,N_13550,N_13372);
or U14282 (N_14282,N_13398,N_13119);
or U14283 (N_14283,N_13072,N_13174);
nor U14284 (N_14284,N_13243,N_13544);
xnor U14285 (N_14285,N_13057,N_13898);
xor U14286 (N_14286,N_13658,N_13021);
xor U14287 (N_14287,N_13376,N_13972);
nor U14288 (N_14288,N_13417,N_13674);
and U14289 (N_14289,N_13001,N_13862);
xor U14290 (N_14290,N_13028,N_13038);
or U14291 (N_14291,N_13091,N_13295);
nor U14292 (N_14292,N_13833,N_13469);
and U14293 (N_14293,N_13194,N_13676);
nor U14294 (N_14294,N_13519,N_13055);
xnor U14295 (N_14295,N_13606,N_13931);
nand U14296 (N_14296,N_13767,N_13832);
nand U14297 (N_14297,N_13053,N_13115);
xor U14298 (N_14298,N_13876,N_13284);
nor U14299 (N_14299,N_13913,N_13388);
nand U14300 (N_14300,N_13836,N_13374);
nand U14301 (N_14301,N_13435,N_13033);
or U14302 (N_14302,N_13684,N_13835);
xor U14303 (N_14303,N_13457,N_13237);
and U14304 (N_14304,N_13485,N_13738);
and U14305 (N_14305,N_13032,N_13155);
and U14306 (N_14306,N_13288,N_13797);
and U14307 (N_14307,N_13125,N_13533);
xor U14308 (N_14308,N_13744,N_13824);
and U14309 (N_14309,N_13692,N_13108);
nand U14310 (N_14310,N_13408,N_13073);
or U14311 (N_14311,N_13178,N_13689);
xnor U14312 (N_14312,N_13255,N_13181);
nor U14313 (N_14313,N_13494,N_13798);
or U14314 (N_14314,N_13731,N_13890);
nor U14315 (N_14315,N_13220,N_13321);
nand U14316 (N_14316,N_13440,N_13045);
and U14317 (N_14317,N_13643,N_13537);
and U14318 (N_14318,N_13725,N_13981);
or U14319 (N_14319,N_13162,N_13870);
nor U14320 (N_14320,N_13052,N_13924);
or U14321 (N_14321,N_13426,N_13760);
and U14322 (N_14322,N_13729,N_13314);
nor U14323 (N_14323,N_13281,N_13698);
or U14324 (N_14324,N_13493,N_13649);
nand U14325 (N_14325,N_13704,N_13951);
or U14326 (N_14326,N_13588,N_13416);
or U14327 (N_14327,N_13207,N_13134);
and U14328 (N_14328,N_13076,N_13147);
nor U14329 (N_14329,N_13554,N_13386);
or U14330 (N_14330,N_13304,N_13568);
and U14331 (N_14331,N_13026,N_13226);
nor U14332 (N_14332,N_13066,N_13602);
nand U14333 (N_14333,N_13779,N_13607);
xnor U14334 (N_14334,N_13352,N_13807);
and U14335 (N_14335,N_13030,N_13970);
and U14336 (N_14336,N_13465,N_13580);
nand U14337 (N_14337,N_13752,N_13714);
nand U14338 (N_14338,N_13409,N_13655);
nand U14339 (N_14339,N_13530,N_13682);
or U14340 (N_14340,N_13141,N_13788);
nor U14341 (N_14341,N_13240,N_13705);
and U14342 (N_14342,N_13184,N_13755);
xor U14343 (N_14343,N_13421,N_13627);
or U14344 (N_14344,N_13620,N_13920);
nor U14345 (N_14345,N_13514,N_13058);
xnor U14346 (N_14346,N_13905,N_13773);
nor U14347 (N_14347,N_13808,N_13911);
xnor U14348 (N_14348,N_13548,N_13628);
nand U14349 (N_14349,N_13249,N_13965);
nor U14350 (N_14350,N_13216,N_13444);
nor U14351 (N_14351,N_13214,N_13660);
nor U14352 (N_14352,N_13339,N_13829);
or U14353 (N_14353,N_13524,N_13885);
nand U14354 (N_14354,N_13648,N_13051);
nor U14355 (N_14355,N_13250,N_13241);
nor U14356 (N_14356,N_13551,N_13656);
xor U14357 (N_14357,N_13270,N_13062);
nor U14358 (N_14358,N_13085,N_13768);
nand U14359 (N_14359,N_13118,N_13232);
and U14360 (N_14360,N_13747,N_13043);
and U14361 (N_14361,N_13834,N_13305);
xor U14362 (N_14362,N_13590,N_13757);
nand U14363 (N_14363,N_13546,N_13391);
or U14364 (N_14364,N_13914,N_13759);
nand U14365 (N_14365,N_13219,N_13923);
xor U14366 (N_14366,N_13880,N_13183);
nor U14367 (N_14367,N_13932,N_13312);
nand U14368 (N_14368,N_13992,N_13322);
and U14369 (N_14369,N_13336,N_13303);
xor U14370 (N_14370,N_13926,N_13816);
xnor U14371 (N_14371,N_13857,N_13300);
and U14372 (N_14372,N_13361,N_13341);
nor U14373 (N_14373,N_13859,N_13978);
and U14374 (N_14374,N_13158,N_13998);
nor U14375 (N_14375,N_13202,N_13930);
or U14376 (N_14376,N_13427,N_13637);
nand U14377 (N_14377,N_13956,N_13665);
and U14378 (N_14378,N_13945,N_13830);
xnor U14379 (N_14379,N_13941,N_13503);
xnor U14380 (N_14380,N_13823,N_13614);
nand U14381 (N_14381,N_13482,N_13921);
xor U14382 (N_14382,N_13638,N_13275);
and U14383 (N_14383,N_13317,N_13504);
and U14384 (N_14384,N_13939,N_13039);
nor U14385 (N_14385,N_13973,N_13233);
nand U14386 (N_14386,N_13582,N_13104);
or U14387 (N_14387,N_13766,N_13611);
and U14388 (N_14388,N_13129,N_13135);
nand U14389 (N_14389,N_13901,N_13925);
nand U14390 (N_14390,N_13443,N_13681);
xnor U14391 (N_14391,N_13642,N_13679);
xnor U14392 (N_14392,N_13944,N_13367);
or U14393 (N_14393,N_13331,N_13585);
nor U14394 (N_14394,N_13510,N_13138);
xnor U14395 (N_14395,N_13193,N_13999);
xnor U14396 (N_14396,N_13023,N_13201);
xor U14397 (N_14397,N_13263,N_13761);
nand U14398 (N_14398,N_13084,N_13173);
and U14399 (N_14399,N_13335,N_13446);
and U14400 (N_14400,N_13536,N_13153);
xor U14401 (N_14401,N_13865,N_13672);
xor U14402 (N_14402,N_13163,N_13474);
xor U14403 (N_14403,N_13601,N_13492);
or U14404 (N_14404,N_13589,N_13940);
nand U14405 (N_14405,N_13459,N_13075);
and U14406 (N_14406,N_13319,N_13074);
or U14407 (N_14407,N_13594,N_13460);
nand U14408 (N_14408,N_13527,N_13903);
or U14409 (N_14409,N_13486,N_13680);
xnor U14410 (N_14410,N_13860,N_13845);
and U14411 (N_14411,N_13204,N_13285);
nand U14412 (N_14412,N_13754,N_13396);
or U14413 (N_14413,N_13323,N_13783);
nand U14414 (N_14414,N_13854,N_13974);
or U14415 (N_14415,N_13646,N_13927);
nor U14416 (N_14416,N_13948,N_13793);
or U14417 (N_14417,N_13516,N_13247);
nand U14418 (N_14418,N_13106,N_13751);
nand U14419 (N_14419,N_13505,N_13330);
nand U14420 (N_14420,N_13563,N_13710);
nand U14421 (N_14421,N_13418,N_13109);
or U14422 (N_14422,N_13987,N_13100);
nor U14423 (N_14423,N_13685,N_13348);
nor U14424 (N_14424,N_13167,N_13878);
nand U14425 (N_14425,N_13160,N_13176);
xor U14426 (N_14426,N_13919,N_13575);
and U14427 (N_14427,N_13910,N_13102);
or U14428 (N_14428,N_13332,N_13888);
xnor U14429 (N_14429,N_13461,N_13380);
and U14430 (N_14430,N_13261,N_13737);
nand U14431 (N_14431,N_13047,N_13500);
or U14432 (N_14432,N_13385,N_13595);
nand U14433 (N_14433,N_13645,N_13796);
and U14434 (N_14434,N_13212,N_13934);
nor U14435 (N_14435,N_13553,N_13148);
xor U14436 (N_14436,N_13591,N_13696);
nor U14437 (N_14437,N_13121,N_13041);
nand U14438 (N_14438,N_13278,N_13346);
nor U14439 (N_14439,N_13936,N_13448);
nand U14440 (N_14440,N_13540,N_13120);
and U14441 (N_14441,N_13307,N_13843);
nor U14442 (N_14442,N_13290,N_13693);
nand U14443 (N_14443,N_13687,N_13549);
and U14444 (N_14444,N_13022,N_13928);
nand U14445 (N_14445,N_13423,N_13005);
xnor U14446 (N_14446,N_13246,N_13145);
nor U14447 (N_14447,N_13501,N_13984);
nor U14448 (N_14448,N_13742,N_13090);
or U14449 (N_14449,N_13140,N_13964);
nand U14450 (N_14450,N_13881,N_13592);
xor U14451 (N_14451,N_13245,N_13093);
nor U14452 (N_14452,N_13042,N_13599);
nor U14453 (N_14453,N_13350,N_13657);
nand U14454 (N_14454,N_13741,N_13434);
xnor U14455 (N_14455,N_13609,N_13238);
nor U14456 (N_14456,N_13002,N_13137);
nand U14457 (N_14457,N_13251,N_13439);
nor U14458 (N_14458,N_13069,N_13991);
or U14459 (N_14459,N_13334,N_13758);
and U14460 (N_14460,N_13966,N_13800);
or U14461 (N_14461,N_13957,N_13980);
and U14462 (N_14462,N_13405,N_13467);
xnor U14463 (N_14463,N_13123,N_13790);
xnor U14464 (N_14464,N_13259,N_13490);
or U14465 (N_14465,N_13712,N_13447);
or U14466 (N_14466,N_13310,N_13103);
xnor U14467 (N_14467,N_13302,N_13515);
or U14468 (N_14468,N_13132,N_13774);
xnor U14469 (N_14469,N_13635,N_13096);
nor U14470 (N_14470,N_13528,N_13619);
nand U14471 (N_14471,N_13502,N_13089);
or U14472 (N_14472,N_13382,N_13746);
xnor U14473 (N_14473,N_13708,N_13394);
xor U14474 (N_14474,N_13846,N_13169);
nand U14475 (N_14475,N_13983,N_13144);
nand U14476 (N_14476,N_13520,N_13205);
nor U14477 (N_14477,N_13722,N_13812);
xnor U14478 (N_14478,N_13686,N_13166);
or U14479 (N_14479,N_13326,N_13097);
or U14480 (N_14480,N_13142,N_13975);
nand U14481 (N_14481,N_13512,N_13721);
or U14482 (N_14482,N_13827,N_13868);
nor U14483 (N_14483,N_13517,N_13390);
xor U14484 (N_14484,N_13006,N_13116);
xor U14485 (N_14485,N_13795,N_13771);
nor U14486 (N_14486,N_13060,N_13906);
xor U14487 (N_14487,N_13422,N_13152);
or U14488 (N_14488,N_13789,N_13316);
nand U14489 (N_14489,N_13855,N_13677);
or U14490 (N_14490,N_13016,N_13433);
and U14491 (N_14491,N_13571,N_13831);
and U14492 (N_14492,N_13177,N_13009);
nor U14493 (N_14493,N_13523,N_13608);
nor U14494 (N_14494,N_13799,N_13821);
xor U14495 (N_14495,N_13286,N_13730);
nand U14496 (N_14496,N_13180,N_13012);
nor U14497 (N_14497,N_13031,N_13724);
and U14498 (N_14498,N_13128,N_13565);
nor U14499 (N_14499,N_13213,N_13566);
xnor U14500 (N_14500,N_13210,N_13587);
nor U14501 (N_14501,N_13143,N_13584);
or U14502 (N_14502,N_13615,N_13001);
or U14503 (N_14503,N_13212,N_13801);
nor U14504 (N_14504,N_13450,N_13138);
nor U14505 (N_14505,N_13928,N_13809);
or U14506 (N_14506,N_13697,N_13839);
xnor U14507 (N_14507,N_13176,N_13302);
and U14508 (N_14508,N_13833,N_13658);
nor U14509 (N_14509,N_13014,N_13162);
or U14510 (N_14510,N_13866,N_13881);
and U14511 (N_14511,N_13534,N_13851);
and U14512 (N_14512,N_13054,N_13591);
and U14513 (N_14513,N_13905,N_13619);
and U14514 (N_14514,N_13483,N_13740);
nor U14515 (N_14515,N_13832,N_13837);
and U14516 (N_14516,N_13569,N_13936);
nand U14517 (N_14517,N_13353,N_13511);
or U14518 (N_14518,N_13829,N_13508);
xnor U14519 (N_14519,N_13264,N_13593);
nor U14520 (N_14520,N_13464,N_13619);
xor U14521 (N_14521,N_13884,N_13407);
xnor U14522 (N_14522,N_13571,N_13201);
nand U14523 (N_14523,N_13286,N_13937);
nand U14524 (N_14524,N_13791,N_13956);
xnor U14525 (N_14525,N_13234,N_13168);
nand U14526 (N_14526,N_13042,N_13683);
and U14527 (N_14527,N_13001,N_13906);
or U14528 (N_14528,N_13109,N_13181);
or U14529 (N_14529,N_13259,N_13730);
or U14530 (N_14530,N_13417,N_13977);
or U14531 (N_14531,N_13949,N_13804);
nor U14532 (N_14532,N_13448,N_13595);
nor U14533 (N_14533,N_13809,N_13443);
xnor U14534 (N_14534,N_13404,N_13317);
xnor U14535 (N_14535,N_13318,N_13664);
and U14536 (N_14536,N_13121,N_13748);
nand U14537 (N_14537,N_13963,N_13818);
or U14538 (N_14538,N_13970,N_13266);
nand U14539 (N_14539,N_13319,N_13131);
or U14540 (N_14540,N_13736,N_13335);
or U14541 (N_14541,N_13589,N_13984);
and U14542 (N_14542,N_13570,N_13206);
nand U14543 (N_14543,N_13966,N_13523);
nand U14544 (N_14544,N_13796,N_13976);
and U14545 (N_14545,N_13103,N_13427);
and U14546 (N_14546,N_13478,N_13220);
and U14547 (N_14547,N_13659,N_13706);
or U14548 (N_14548,N_13881,N_13725);
nor U14549 (N_14549,N_13705,N_13313);
xnor U14550 (N_14550,N_13781,N_13251);
or U14551 (N_14551,N_13646,N_13763);
nand U14552 (N_14552,N_13160,N_13568);
nor U14553 (N_14553,N_13501,N_13915);
nor U14554 (N_14554,N_13231,N_13319);
nand U14555 (N_14555,N_13493,N_13325);
and U14556 (N_14556,N_13673,N_13132);
nor U14557 (N_14557,N_13708,N_13741);
or U14558 (N_14558,N_13828,N_13480);
and U14559 (N_14559,N_13509,N_13665);
and U14560 (N_14560,N_13658,N_13432);
nor U14561 (N_14561,N_13372,N_13195);
and U14562 (N_14562,N_13598,N_13618);
nand U14563 (N_14563,N_13744,N_13300);
nor U14564 (N_14564,N_13923,N_13519);
or U14565 (N_14565,N_13549,N_13211);
or U14566 (N_14566,N_13711,N_13556);
or U14567 (N_14567,N_13129,N_13808);
nor U14568 (N_14568,N_13249,N_13552);
xor U14569 (N_14569,N_13709,N_13604);
and U14570 (N_14570,N_13809,N_13017);
nor U14571 (N_14571,N_13288,N_13737);
or U14572 (N_14572,N_13505,N_13828);
nor U14573 (N_14573,N_13145,N_13684);
nand U14574 (N_14574,N_13205,N_13046);
or U14575 (N_14575,N_13752,N_13539);
or U14576 (N_14576,N_13433,N_13712);
xnor U14577 (N_14577,N_13022,N_13258);
nor U14578 (N_14578,N_13174,N_13782);
and U14579 (N_14579,N_13739,N_13217);
nor U14580 (N_14580,N_13006,N_13688);
and U14581 (N_14581,N_13386,N_13129);
nor U14582 (N_14582,N_13661,N_13663);
or U14583 (N_14583,N_13049,N_13094);
nand U14584 (N_14584,N_13015,N_13407);
nor U14585 (N_14585,N_13577,N_13591);
nor U14586 (N_14586,N_13256,N_13754);
xnor U14587 (N_14587,N_13951,N_13799);
xor U14588 (N_14588,N_13476,N_13821);
and U14589 (N_14589,N_13920,N_13388);
or U14590 (N_14590,N_13995,N_13790);
nand U14591 (N_14591,N_13376,N_13887);
and U14592 (N_14592,N_13690,N_13052);
or U14593 (N_14593,N_13695,N_13043);
or U14594 (N_14594,N_13116,N_13210);
and U14595 (N_14595,N_13216,N_13155);
nand U14596 (N_14596,N_13498,N_13960);
and U14597 (N_14597,N_13376,N_13322);
nor U14598 (N_14598,N_13065,N_13327);
xnor U14599 (N_14599,N_13330,N_13222);
nor U14600 (N_14600,N_13929,N_13180);
and U14601 (N_14601,N_13692,N_13258);
and U14602 (N_14602,N_13642,N_13064);
nor U14603 (N_14603,N_13800,N_13349);
xnor U14604 (N_14604,N_13476,N_13175);
nor U14605 (N_14605,N_13144,N_13539);
and U14606 (N_14606,N_13450,N_13502);
or U14607 (N_14607,N_13990,N_13374);
and U14608 (N_14608,N_13388,N_13153);
or U14609 (N_14609,N_13175,N_13796);
or U14610 (N_14610,N_13063,N_13565);
nand U14611 (N_14611,N_13252,N_13640);
nand U14612 (N_14612,N_13975,N_13787);
xor U14613 (N_14613,N_13260,N_13832);
or U14614 (N_14614,N_13221,N_13791);
nand U14615 (N_14615,N_13772,N_13090);
and U14616 (N_14616,N_13243,N_13817);
or U14617 (N_14617,N_13956,N_13763);
and U14618 (N_14618,N_13042,N_13523);
nand U14619 (N_14619,N_13192,N_13365);
and U14620 (N_14620,N_13899,N_13137);
and U14621 (N_14621,N_13933,N_13704);
nor U14622 (N_14622,N_13050,N_13913);
xnor U14623 (N_14623,N_13295,N_13522);
or U14624 (N_14624,N_13056,N_13768);
nor U14625 (N_14625,N_13499,N_13264);
nor U14626 (N_14626,N_13502,N_13299);
and U14627 (N_14627,N_13919,N_13783);
nor U14628 (N_14628,N_13646,N_13849);
xor U14629 (N_14629,N_13446,N_13876);
or U14630 (N_14630,N_13583,N_13398);
nand U14631 (N_14631,N_13896,N_13337);
xnor U14632 (N_14632,N_13505,N_13531);
and U14633 (N_14633,N_13743,N_13260);
or U14634 (N_14634,N_13819,N_13785);
nor U14635 (N_14635,N_13218,N_13289);
nor U14636 (N_14636,N_13783,N_13612);
and U14637 (N_14637,N_13146,N_13999);
nor U14638 (N_14638,N_13109,N_13883);
nor U14639 (N_14639,N_13127,N_13276);
and U14640 (N_14640,N_13844,N_13910);
and U14641 (N_14641,N_13756,N_13111);
nand U14642 (N_14642,N_13556,N_13008);
xor U14643 (N_14643,N_13790,N_13994);
and U14644 (N_14644,N_13044,N_13273);
xor U14645 (N_14645,N_13155,N_13059);
nand U14646 (N_14646,N_13519,N_13728);
nor U14647 (N_14647,N_13159,N_13224);
nand U14648 (N_14648,N_13549,N_13755);
xor U14649 (N_14649,N_13517,N_13535);
and U14650 (N_14650,N_13602,N_13379);
nor U14651 (N_14651,N_13103,N_13659);
or U14652 (N_14652,N_13499,N_13722);
nor U14653 (N_14653,N_13059,N_13870);
and U14654 (N_14654,N_13295,N_13818);
xnor U14655 (N_14655,N_13145,N_13006);
and U14656 (N_14656,N_13235,N_13534);
nand U14657 (N_14657,N_13677,N_13464);
nor U14658 (N_14658,N_13628,N_13618);
or U14659 (N_14659,N_13072,N_13269);
or U14660 (N_14660,N_13166,N_13192);
xor U14661 (N_14661,N_13449,N_13391);
nor U14662 (N_14662,N_13635,N_13046);
or U14663 (N_14663,N_13837,N_13548);
nor U14664 (N_14664,N_13251,N_13018);
xnor U14665 (N_14665,N_13839,N_13444);
nand U14666 (N_14666,N_13274,N_13647);
xor U14667 (N_14667,N_13479,N_13828);
xor U14668 (N_14668,N_13091,N_13744);
nand U14669 (N_14669,N_13869,N_13676);
nand U14670 (N_14670,N_13734,N_13072);
nand U14671 (N_14671,N_13424,N_13114);
nor U14672 (N_14672,N_13243,N_13283);
nor U14673 (N_14673,N_13363,N_13188);
nor U14674 (N_14674,N_13955,N_13277);
nor U14675 (N_14675,N_13887,N_13097);
or U14676 (N_14676,N_13350,N_13115);
and U14677 (N_14677,N_13304,N_13142);
xor U14678 (N_14678,N_13148,N_13933);
or U14679 (N_14679,N_13234,N_13072);
xor U14680 (N_14680,N_13934,N_13585);
and U14681 (N_14681,N_13042,N_13675);
nand U14682 (N_14682,N_13223,N_13884);
and U14683 (N_14683,N_13296,N_13884);
nand U14684 (N_14684,N_13933,N_13339);
or U14685 (N_14685,N_13435,N_13394);
and U14686 (N_14686,N_13276,N_13404);
nor U14687 (N_14687,N_13119,N_13278);
nand U14688 (N_14688,N_13546,N_13506);
or U14689 (N_14689,N_13460,N_13150);
xor U14690 (N_14690,N_13032,N_13197);
and U14691 (N_14691,N_13365,N_13206);
and U14692 (N_14692,N_13855,N_13745);
nand U14693 (N_14693,N_13682,N_13957);
and U14694 (N_14694,N_13040,N_13020);
nand U14695 (N_14695,N_13928,N_13882);
and U14696 (N_14696,N_13382,N_13176);
nor U14697 (N_14697,N_13899,N_13609);
nor U14698 (N_14698,N_13496,N_13203);
or U14699 (N_14699,N_13320,N_13142);
nor U14700 (N_14700,N_13953,N_13898);
or U14701 (N_14701,N_13927,N_13737);
xnor U14702 (N_14702,N_13537,N_13812);
xnor U14703 (N_14703,N_13888,N_13650);
nor U14704 (N_14704,N_13195,N_13432);
nand U14705 (N_14705,N_13109,N_13411);
or U14706 (N_14706,N_13287,N_13403);
or U14707 (N_14707,N_13641,N_13398);
or U14708 (N_14708,N_13134,N_13531);
or U14709 (N_14709,N_13896,N_13272);
nand U14710 (N_14710,N_13065,N_13338);
nor U14711 (N_14711,N_13801,N_13886);
and U14712 (N_14712,N_13896,N_13712);
or U14713 (N_14713,N_13201,N_13448);
nand U14714 (N_14714,N_13980,N_13017);
xnor U14715 (N_14715,N_13362,N_13375);
nor U14716 (N_14716,N_13979,N_13759);
and U14717 (N_14717,N_13239,N_13333);
nand U14718 (N_14718,N_13159,N_13145);
nor U14719 (N_14719,N_13317,N_13343);
or U14720 (N_14720,N_13889,N_13805);
xnor U14721 (N_14721,N_13369,N_13980);
nand U14722 (N_14722,N_13194,N_13814);
or U14723 (N_14723,N_13933,N_13844);
or U14724 (N_14724,N_13550,N_13599);
nand U14725 (N_14725,N_13786,N_13569);
and U14726 (N_14726,N_13749,N_13731);
and U14727 (N_14727,N_13369,N_13828);
xor U14728 (N_14728,N_13341,N_13733);
nand U14729 (N_14729,N_13140,N_13218);
nor U14730 (N_14730,N_13362,N_13405);
and U14731 (N_14731,N_13560,N_13238);
nand U14732 (N_14732,N_13405,N_13227);
nor U14733 (N_14733,N_13242,N_13354);
and U14734 (N_14734,N_13880,N_13457);
nor U14735 (N_14735,N_13272,N_13855);
and U14736 (N_14736,N_13852,N_13458);
xor U14737 (N_14737,N_13350,N_13517);
xor U14738 (N_14738,N_13896,N_13091);
and U14739 (N_14739,N_13547,N_13255);
xor U14740 (N_14740,N_13582,N_13608);
nand U14741 (N_14741,N_13810,N_13233);
nor U14742 (N_14742,N_13881,N_13929);
or U14743 (N_14743,N_13109,N_13845);
nand U14744 (N_14744,N_13865,N_13816);
and U14745 (N_14745,N_13816,N_13917);
xor U14746 (N_14746,N_13730,N_13296);
nand U14747 (N_14747,N_13608,N_13220);
nand U14748 (N_14748,N_13844,N_13313);
nor U14749 (N_14749,N_13595,N_13013);
or U14750 (N_14750,N_13758,N_13484);
nand U14751 (N_14751,N_13078,N_13207);
xnor U14752 (N_14752,N_13916,N_13319);
nand U14753 (N_14753,N_13149,N_13311);
xnor U14754 (N_14754,N_13856,N_13402);
nor U14755 (N_14755,N_13096,N_13658);
nor U14756 (N_14756,N_13146,N_13645);
or U14757 (N_14757,N_13787,N_13558);
or U14758 (N_14758,N_13678,N_13379);
nor U14759 (N_14759,N_13818,N_13008);
and U14760 (N_14760,N_13715,N_13661);
or U14761 (N_14761,N_13461,N_13357);
and U14762 (N_14762,N_13217,N_13977);
nor U14763 (N_14763,N_13606,N_13452);
or U14764 (N_14764,N_13131,N_13953);
nor U14765 (N_14765,N_13110,N_13759);
or U14766 (N_14766,N_13655,N_13643);
nor U14767 (N_14767,N_13697,N_13634);
nor U14768 (N_14768,N_13063,N_13725);
nor U14769 (N_14769,N_13397,N_13047);
nor U14770 (N_14770,N_13217,N_13691);
or U14771 (N_14771,N_13020,N_13192);
and U14772 (N_14772,N_13364,N_13392);
nor U14773 (N_14773,N_13179,N_13830);
nand U14774 (N_14774,N_13116,N_13559);
nand U14775 (N_14775,N_13498,N_13653);
nand U14776 (N_14776,N_13269,N_13762);
nor U14777 (N_14777,N_13994,N_13327);
xnor U14778 (N_14778,N_13092,N_13646);
and U14779 (N_14779,N_13209,N_13734);
nor U14780 (N_14780,N_13964,N_13979);
and U14781 (N_14781,N_13236,N_13359);
xnor U14782 (N_14782,N_13355,N_13003);
xnor U14783 (N_14783,N_13166,N_13285);
nor U14784 (N_14784,N_13664,N_13055);
xor U14785 (N_14785,N_13407,N_13762);
nor U14786 (N_14786,N_13713,N_13179);
nand U14787 (N_14787,N_13364,N_13090);
nand U14788 (N_14788,N_13594,N_13849);
xnor U14789 (N_14789,N_13669,N_13369);
nor U14790 (N_14790,N_13016,N_13902);
xor U14791 (N_14791,N_13593,N_13341);
nand U14792 (N_14792,N_13694,N_13124);
and U14793 (N_14793,N_13234,N_13116);
nor U14794 (N_14794,N_13367,N_13633);
or U14795 (N_14795,N_13643,N_13150);
xnor U14796 (N_14796,N_13146,N_13027);
and U14797 (N_14797,N_13753,N_13712);
xor U14798 (N_14798,N_13803,N_13043);
xnor U14799 (N_14799,N_13792,N_13234);
and U14800 (N_14800,N_13209,N_13856);
or U14801 (N_14801,N_13963,N_13168);
and U14802 (N_14802,N_13133,N_13763);
nor U14803 (N_14803,N_13405,N_13485);
or U14804 (N_14804,N_13454,N_13147);
xnor U14805 (N_14805,N_13543,N_13698);
or U14806 (N_14806,N_13165,N_13714);
nor U14807 (N_14807,N_13574,N_13300);
xor U14808 (N_14808,N_13325,N_13709);
and U14809 (N_14809,N_13360,N_13124);
or U14810 (N_14810,N_13259,N_13729);
or U14811 (N_14811,N_13276,N_13723);
or U14812 (N_14812,N_13539,N_13646);
xnor U14813 (N_14813,N_13898,N_13741);
and U14814 (N_14814,N_13275,N_13296);
nand U14815 (N_14815,N_13634,N_13709);
and U14816 (N_14816,N_13356,N_13155);
and U14817 (N_14817,N_13717,N_13626);
xnor U14818 (N_14818,N_13732,N_13454);
or U14819 (N_14819,N_13265,N_13986);
xor U14820 (N_14820,N_13983,N_13777);
and U14821 (N_14821,N_13192,N_13924);
nor U14822 (N_14822,N_13283,N_13223);
xnor U14823 (N_14823,N_13378,N_13797);
nor U14824 (N_14824,N_13561,N_13508);
nor U14825 (N_14825,N_13218,N_13870);
or U14826 (N_14826,N_13140,N_13702);
nand U14827 (N_14827,N_13420,N_13653);
or U14828 (N_14828,N_13309,N_13756);
or U14829 (N_14829,N_13366,N_13342);
nor U14830 (N_14830,N_13852,N_13157);
xor U14831 (N_14831,N_13627,N_13207);
nand U14832 (N_14832,N_13963,N_13972);
and U14833 (N_14833,N_13079,N_13260);
or U14834 (N_14834,N_13690,N_13125);
or U14835 (N_14835,N_13414,N_13172);
or U14836 (N_14836,N_13927,N_13437);
nand U14837 (N_14837,N_13101,N_13439);
or U14838 (N_14838,N_13733,N_13560);
nor U14839 (N_14839,N_13622,N_13093);
and U14840 (N_14840,N_13173,N_13579);
xor U14841 (N_14841,N_13791,N_13200);
and U14842 (N_14842,N_13299,N_13129);
nor U14843 (N_14843,N_13553,N_13857);
nor U14844 (N_14844,N_13757,N_13638);
xnor U14845 (N_14845,N_13689,N_13855);
and U14846 (N_14846,N_13172,N_13533);
nor U14847 (N_14847,N_13808,N_13252);
nor U14848 (N_14848,N_13349,N_13693);
and U14849 (N_14849,N_13193,N_13057);
nor U14850 (N_14850,N_13473,N_13283);
and U14851 (N_14851,N_13735,N_13264);
and U14852 (N_14852,N_13978,N_13597);
and U14853 (N_14853,N_13714,N_13605);
or U14854 (N_14854,N_13666,N_13103);
nand U14855 (N_14855,N_13679,N_13286);
and U14856 (N_14856,N_13196,N_13260);
nand U14857 (N_14857,N_13771,N_13877);
nand U14858 (N_14858,N_13396,N_13043);
or U14859 (N_14859,N_13591,N_13551);
or U14860 (N_14860,N_13185,N_13516);
and U14861 (N_14861,N_13982,N_13747);
nor U14862 (N_14862,N_13008,N_13104);
nand U14863 (N_14863,N_13235,N_13142);
xnor U14864 (N_14864,N_13497,N_13463);
nand U14865 (N_14865,N_13199,N_13538);
or U14866 (N_14866,N_13579,N_13687);
and U14867 (N_14867,N_13644,N_13952);
xor U14868 (N_14868,N_13852,N_13165);
or U14869 (N_14869,N_13024,N_13801);
and U14870 (N_14870,N_13380,N_13559);
and U14871 (N_14871,N_13186,N_13228);
xnor U14872 (N_14872,N_13296,N_13038);
and U14873 (N_14873,N_13600,N_13096);
nand U14874 (N_14874,N_13538,N_13346);
and U14875 (N_14875,N_13684,N_13390);
and U14876 (N_14876,N_13331,N_13621);
and U14877 (N_14877,N_13637,N_13697);
nor U14878 (N_14878,N_13886,N_13538);
nor U14879 (N_14879,N_13716,N_13961);
xnor U14880 (N_14880,N_13197,N_13039);
xnor U14881 (N_14881,N_13955,N_13364);
xnor U14882 (N_14882,N_13055,N_13396);
and U14883 (N_14883,N_13303,N_13278);
xor U14884 (N_14884,N_13047,N_13771);
nor U14885 (N_14885,N_13651,N_13176);
or U14886 (N_14886,N_13161,N_13253);
xor U14887 (N_14887,N_13852,N_13396);
or U14888 (N_14888,N_13435,N_13661);
xnor U14889 (N_14889,N_13035,N_13246);
nor U14890 (N_14890,N_13756,N_13767);
nor U14891 (N_14891,N_13761,N_13087);
nand U14892 (N_14892,N_13843,N_13892);
and U14893 (N_14893,N_13972,N_13609);
and U14894 (N_14894,N_13021,N_13003);
nand U14895 (N_14895,N_13659,N_13364);
or U14896 (N_14896,N_13842,N_13403);
or U14897 (N_14897,N_13760,N_13438);
or U14898 (N_14898,N_13063,N_13678);
or U14899 (N_14899,N_13994,N_13365);
xor U14900 (N_14900,N_13402,N_13548);
and U14901 (N_14901,N_13633,N_13328);
nand U14902 (N_14902,N_13240,N_13653);
nor U14903 (N_14903,N_13065,N_13776);
or U14904 (N_14904,N_13918,N_13934);
xor U14905 (N_14905,N_13034,N_13765);
and U14906 (N_14906,N_13946,N_13795);
nand U14907 (N_14907,N_13426,N_13732);
and U14908 (N_14908,N_13557,N_13674);
and U14909 (N_14909,N_13493,N_13357);
xor U14910 (N_14910,N_13174,N_13298);
or U14911 (N_14911,N_13002,N_13806);
nor U14912 (N_14912,N_13756,N_13419);
and U14913 (N_14913,N_13613,N_13176);
nand U14914 (N_14914,N_13446,N_13085);
nor U14915 (N_14915,N_13514,N_13858);
and U14916 (N_14916,N_13406,N_13975);
nand U14917 (N_14917,N_13285,N_13207);
xnor U14918 (N_14918,N_13575,N_13440);
or U14919 (N_14919,N_13870,N_13785);
or U14920 (N_14920,N_13970,N_13207);
nor U14921 (N_14921,N_13054,N_13864);
or U14922 (N_14922,N_13066,N_13750);
and U14923 (N_14923,N_13577,N_13698);
or U14924 (N_14924,N_13912,N_13110);
or U14925 (N_14925,N_13588,N_13239);
or U14926 (N_14926,N_13873,N_13332);
xor U14927 (N_14927,N_13437,N_13401);
nor U14928 (N_14928,N_13386,N_13808);
nor U14929 (N_14929,N_13964,N_13352);
xnor U14930 (N_14930,N_13210,N_13554);
nand U14931 (N_14931,N_13205,N_13732);
or U14932 (N_14932,N_13128,N_13095);
or U14933 (N_14933,N_13979,N_13035);
and U14934 (N_14934,N_13740,N_13283);
and U14935 (N_14935,N_13810,N_13175);
and U14936 (N_14936,N_13736,N_13207);
xnor U14937 (N_14937,N_13401,N_13990);
xnor U14938 (N_14938,N_13128,N_13004);
nand U14939 (N_14939,N_13188,N_13799);
xnor U14940 (N_14940,N_13430,N_13719);
xor U14941 (N_14941,N_13939,N_13044);
and U14942 (N_14942,N_13823,N_13964);
xor U14943 (N_14943,N_13678,N_13825);
and U14944 (N_14944,N_13321,N_13745);
nor U14945 (N_14945,N_13276,N_13601);
or U14946 (N_14946,N_13603,N_13976);
xor U14947 (N_14947,N_13355,N_13587);
nor U14948 (N_14948,N_13561,N_13637);
or U14949 (N_14949,N_13397,N_13974);
or U14950 (N_14950,N_13533,N_13105);
or U14951 (N_14951,N_13217,N_13047);
or U14952 (N_14952,N_13513,N_13345);
and U14953 (N_14953,N_13644,N_13714);
nor U14954 (N_14954,N_13021,N_13535);
nand U14955 (N_14955,N_13948,N_13768);
nand U14956 (N_14956,N_13910,N_13928);
nor U14957 (N_14957,N_13191,N_13733);
nor U14958 (N_14958,N_13175,N_13615);
or U14959 (N_14959,N_13676,N_13825);
and U14960 (N_14960,N_13369,N_13189);
and U14961 (N_14961,N_13467,N_13626);
and U14962 (N_14962,N_13095,N_13436);
nand U14963 (N_14963,N_13861,N_13481);
or U14964 (N_14964,N_13431,N_13331);
nor U14965 (N_14965,N_13552,N_13980);
xnor U14966 (N_14966,N_13809,N_13405);
nand U14967 (N_14967,N_13064,N_13313);
or U14968 (N_14968,N_13214,N_13851);
or U14969 (N_14969,N_13827,N_13649);
nor U14970 (N_14970,N_13749,N_13409);
and U14971 (N_14971,N_13350,N_13774);
and U14972 (N_14972,N_13214,N_13566);
nand U14973 (N_14973,N_13979,N_13286);
or U14974 (N_14974,N_13466,N_13374);
and U14975 (N_14975,N_13110,N_13253);
nand U14976 (N_14976,N_13296,N_13017);
nor U14977 (N_14977,N_13536,N_13812);
or U14978 (N_14978,N_13830,N_13486);
nor U14979 (N_14979,N_13283,N_13230);
xor U14980 (N_14980,N_13634,N_13116);
xnor U14981 (N_14981,N_13023,N_13254);
xnor U14982 (N_14982,N_13184,N_13156);
nand U14983 (N_14983,N_13424,N_13316);
nor U14984 (N_14984,N_13064,N_13880);
and U14985 (N_14985,N_13581,N_13324);
or U14986 (N_14986,N_13769,N_13571);
nor U14987 (N_14987,N_13460,N_13383);
xnor U14988 (N_14988,N_13125,N_13554);
xnor U14989 (N_14989,N_13618,N_13307);
nor U14990 (N_14990,N_13114,N_13594);
nor U14991 (N_14991,N_13868,N_13289);
and U14992 (N_14992,N_13838,N_13530);
nor U14993 (N_14993,N_13126,N_13601);
xor U14994 (N_14994,N_13175,N_13998);
xnor U14995 (N_14995,N_13501,N_13431);
xnor U14996 (N_14996,N_13203,N_13259);
and U14997 (N_14997,N_13421,N_13526);
nor U14998 (N_14998,N_13973,N_13498);
or U14999 (N_14999,N_13580,N_13723);
nand U15000 (N_15000,N_14917,N_14305);
or U15001 (N_15001,N_14892,N_14093);
xnor U15002 (N_15002,N_14272,N_14865);
nand U15003 (N_15003,N_14783,N_14938);
or U15004 (N_15004,N_14220,N_14110);
or U15005 (N_15005,N_14544,N_14844);
or U15006 (N_15006,N_14129,N_14121);
nand U15007 (N_15007,N_14323,N_14540);
nor U15008 (N_15008,N_14712,N_14051);
nand U15009 (N_15009,N_14022,N_14391);
and U15010 (N_15010,N_14192,N_14805);
or U15011 (N_15011,N_14592,N_14874);
nand U15012 (N_15012,N_14378,N_14873);
xor U15013 (N_15013,N_14909,N_14743);
xor U15014 (N_15014,N_14269,N_14566);
and U15015 (N_15015,N_14530,N_14700);
xnor U15016 (N_15016,N_14039,N_14058);
xor U15017 (N_15017,N_14036,N_14406);
and U15018 (N_15018,N_14173,N_14932);
xnor U15019 (N_15019,N_14726,N_14381);
nand U15020 (N_15020,N_14621,N_14005);
xor U15021 (N_15021,N_14738,N_14496);
xor U15022 (N_15022,N_14382,N_14214);
and U15023 (N_15023,N_14798,N_14950);
nor U15024 (N_15024,N_14218,N_14000);
nand U15025 (N_15025,N_14067,N_14984);
and U15026 (N_15026,N_14646,N_14167);
nand U15027 (N_15027,N_14597,N_14209);
xor U15028 (N_15028,N_14778,N_14763);
nand U15029 (N_15029,N_14516,N_14190);
xor U15030 (N_15030,N_14359,N_14452);
nand U15031 (N_15031,N_14575,N_14432);
xor U15032 (N_15032,N_14979,N_14273);
or U15033 (N_15033,N_14425,N_14593);
nand U15034 (N_15034,N_14056,N_14640);
and U15035 (N_15035,N_14910,N_14714);
xor U15036 (N_15036,N_14741,N_14681);
and U15037 (N_15037,N_14752,N_14825);
nor U15038 (N_15038,N_14729,N_14390);
nor U15039 (N_15039,N_14493,N_14508);
nand U15040 (N_15040,N_14528,N_14655);
nor U15041 (N_15041,N_14806,N_14164);
and U15042 (N_15042,N_14716,N_14614);
and U15043 (N_15043,N_14298,N_14311);
nor U15044 (N_15044,N_14072,N_14629);
or U15045 (N_15045,N_14466,N_14510);
and U15046 (N_15046,N_14046,N_14203);
nor U15047 (N_15047,N_14157,N_14135);
or U15048 (N_15048,N_14771,N_14394);
xor U15049 (N_15049,N_14478,N_14561);
nand U15050 (N_15050,N_14703,N_14413);
xnor U15051 (N_15051,N_14310,N_14520);
nor U15052 (N_15052,N_14849,N_14212);
nand U15053 (N_15053,N_14125,N_14319);
or U15054 (N_15054,N_14078,N_14997);
xor U15055 (N_15055,N_14579,N_14563);
nor U15056 (N_15056,N_14309,N_14816);
or U15057 (N_15057,N_14337,N_14833);
xor U15058 (N_15058,N_14952,N_14471);
nor U15059 (N_15059,N_14601,N_14670);
or U15060 (N_15060,N_14815,N_14596);
and U15061 (N_15061,N_14534,N_14559);
and U15062 (N_15062,N_14308,N_14789);
and U15063 (N_15063,N_14573,N_14436);
and U15064 (N_15064,N_14202,N_14299);
and U15065 (N_15065,N_14194,N_14188);
nor U15066 (N_15066,N_14928,N_14731);
or U15067 (N_15067,N_14554,N_14047);
nand U15068 (N_15068,N_14132,N_14043);
or U15069 (N_15069,N_14669,N_14662);
or U15070 (N_15070,N_14724,N_14506);
xnor U15071 (N_15071,N_14024,N_14230);
and U15072 (N_15072,N_14503,N_14542);
or U15073 (N_15073,N_14238,N_14946);
and U15074 (N_15074,N_14571,N_14913);
and U15075 (N_15075,N_14907,N_14021);
nand U15076 (N_15076,N_14992,N_14007);
or U15077 (N_15077,N_14967,N_14820);
nor U15078 (N_15078,N_14585,N_14514);
nor U15079 (N_15079,N_14822,N_14410);
and U15080 (N_15080,N_14229,N_14297);
and U15081 (N_15081,N_14006,N_14600);
or U15082 (N_15082,N_14341,N_14695);
nor U15083 (N_15083,N_14965,N_14330);
nor U15084 (N_15084,N_14282,N_14186);
or U15085 (N_15085,N_14964,N_14504);
nor U15086 (N_15086,N_14901,N_14953);
xnor U15087 (N_15087,N_14792,N_14444);
or U15088 (N_15088,N_14624,N_14620);
or U15089 (N_15089,N_14161,N_14197);
or U15090 (N_15090,N_14656,N_14259);
nor U15091 (N_15091,N_14782,N_14615);
and U15092 (N_15092,N_14607,N_14667);
or U15093 (N_15093,N_14940,N_14483);
nor U15094 (N_15094,N_14160,N_14603);
xor U15095 (N_15095,N_14112,N_14799);
nand U15096 (N_15096,N_14012,N_14899);
or U15097 (N_15097,N_14252,N_14883);
nor U15098 (N_15098,N_14458,N_14787);
nor U15099 (N_15099,N_14963,N_14491);
and U15100 (N_15100,N_14035,N_14602);
or U15101 (N_15101,N_14584,N_14316);
nor U15102 (N_15102,N_14463,N_14288);
or U15103 (N_15103,N_14296,N_14709);
or U15104 (N_15104,N_14393,N_14059);
xor U15105 (N_15105,N_14980,N_14420);
nor U15106 (N_15106,N_14985,N_14786);
and U15107 (N_15107,N_14268,N_14589);
nor U15108 (N_15108,N_14598,N_14223);
or U15109 (N_15109,N_14742,N_14176);
nor U15110 (N_15110,N_14399,N_14156);
nand U15111 (N_15111,N_14912,N_14405);
and U15112 (N_15112,N_14877,N_14306);
nor U15113 (N_15113,N_14948,N_14148);
nand U15114 (N_15114,N_14389,N_14092);
nand U15115 (N_15115,N_14210,N_14746);
and U15116 (N_15116,N_14501,N_14085);
xnor U15117 (N_15117,N_14758,N_14224);
nand U15118 (N_15118,N_14802,N_14438);
and U15119 (N_15119,N_14234,N_14766);
and U15120 (N_15120,N_14395,N_14529);
or U15121 (N_15121,N_14527,N_14141);
nand U15122 (N_15122,N_14809,N_14146);
nor U15123 (N_15123,N_14240,N_14077);
and U15124 (N_15124,N_14130,N_14179);
nand U15125 (N_15125,N_14287,N_14026);
nand U15126 (N_15126,N_14930,N_14631);
nor U15127 (N_15127,N_14718,N_14834);
xnor U15128 (N_15128,N_14537,N_14352);
nor U15129 (N_15129,N_14237,N_14578);
nand U15130 (N_15130,N_14266,N_14847);
nor U15131 (N_15131,N_14497,N_14418);
and U15132 (N_15132,N_14217,N_14808);
nor U15133 (N_15133,N_14574,N_14842);
and U15134 (N_15134,N_14256,N_14293);
nand U15135 (N_15135,N_14680,N_14991);
and U15136 (N_15136,N_14064,N_14430);
xor U15137 (N_15137,N_14871,N_14660);
or U15138 (N_15138,N_14856,N_14857);
xor U15139 (N_15139,N_14696,N_14375);
xnor U15140 (N_15140,N_14138,N_14705);
xnor U15141 (N_15141,N_14253,N_14890);
and U15142 (N_15142,N_14443,N_14276);
xnor U15143 (N_15143,N_14748,N_14502);
nor U15144 (N_15144,N_14469,N_14710);
and U15145 (N_15145,N_14962,N_14102);
and U15146 (N_15146,N_14292,N_14960);
or U15147 (N_15147,N_14550,N_14313);
and U15148 (N_15148,N_14082,N_14042);
or U15149 (N_15149,N_14264,N_14285);
nor U15150 (N_15150,N_14100,N_14115);
nor U15151 (N_15151,N_14307,N_14289);
nor U15152 (N_15152,N_14546,N_14380);
xor U15153 (N_15153,N_14027,N_14236);
and U15154 (N_15154,N_14470,N_14442);
xor U15155 (N_15155,N_14701,N_14541);
or U15156 (N_15156,N_14075,N_14242);
or U15157 (N_15157,N_14248,N_14807);
xnor U15158 (N_15158,N_14676,N_14780);
or U15159 (N_15159,N_14525,N_14531);
and U15160 (N_15160,N_14122,N_14685);
nand U15161 (N_15161,N_14126,N_14467);
or U15162 (N_15162,N_14657,N_14623);
and U15163 (N_15163,N_14207,N_14038);
nand U15164 (N_15164,N_14446,N_14290);
xnor U15165 (N_15165,N_14383,N_14166);
nor U15166 (N_15166,N_14903,N_14532);
nor U15167 (N_15167,N_14972,N_14066);
nor U15168 (N_15168,N_14011,N_14127);
nand U15169 (N_15169,N_14793,N_14835);
nor U15170 (N_15170,N_14401,N_14206);
and U15171 (N_15171,N_14136,N_14008);
xnor U15172 (N_15172,N_14734,N_14565);
nand U15173 (N_15173,N_14016,N_14211);
xnor U15174 (N_15174,N_14906,N_14109);
or U15175 (N_15175,N_14029,N_14587);
and U15176 (N_15176,N_14402,N_14949);
nand U15177 (N_15177,N_14325,N_14751);
nor U15178 (N_15178,N_14978,N_14174);
nor U15179 (N_15179,N_14454,N_14317);
and U15180 (N_15180,N_14117,N_14908);
nor U15181 (N_15181,N_14988,N_14694);
and U15182 (N_15182,N_14435,N_14411);
or U15183 (N_15183,N_14990,N_14720);
nor U15184 (N_15184,N_14241,N_14335);
nor U15185 (N_15185,N_14878,N_14526);
nor U15186 (N_15186,N_14827,N_14208);
nand U15187 (N_15187,N_14699,N_14374);
nand U15188 (N_15188,N_14279,N_14398);
nand U15189 (N_15189,N_14576,N_14353);
or U15190 (N_15190,N_14215,N_14538);
nor U15191 (N_15191,N_14774,N_14314);
nand U15192 (N_15192,N_14545,N_14989);
and U15193 (N_15193,N_14665,N_14858);
nor U15194 (N_15194,N_14781,N_14582);
nand U15195 (N_15195,N_14180,N_14688);
nor U15196 (N_15196,N_14547,N_14143);
and U15197 (N_15197,N_14139,N_14057);
nor U15198 (N_15198,N_14934,N_14977);
xnor U15199 (N_15199,N_14070,N_14089);
and U15200 (N_15200,N_14837,N_14653);
or U15201 (N_15201,N_14227,N_14684);
and U15202 (N_15202,N_14733,N_14864);
xnor U15203 (N_15203,N_14823,N_14678);
nor U15204 (N_15204,N_14618,N_14111);
xnor U15205 (N_15205,N_14348,N_14982);
nor U15206 (N_15206,N_14044,N_14113);
nor U15207 (N_15207,N_14756,N_14155);
xor U15208 (N_15208,N_14866,N_14668);
nand U15209 (N_15209,N_14409,N_14826);
xnor U15210 (N_15210,N_14365,N_14959);
nor U15211 (N_15211,N_14830,N_14052);
xnor U15212 (N_15212,N_14097,N_14628);
and U15213 (N_15213,N_14862,N_14069);
and U15214 (N_15214,N_14191,N_14717);
xor U15215 (N_15215,N_14358,N_14889);
nand U15216 (N_15216,N_14009,N_14679);
and U15217 (N_15217,N_14996,N_14107);
xor U15218 (N_15218,N_14686,N_14448);
nand U15219 (N_15219,N_14961,N_14507);
nor U15220 (N_15220,N_14854,N_14450);
nand U15221 (N_15221,N_14187,N_14321);
and U15222 (N_15222,N_14821,N_14281);
nand U15223 (N_15223,N_14388,N_14020);
or U15224 (N_15224,N_14079,N_14274);
nand U15225 (N_15225,N_14441,N_14755);
nor U15226 (N_15226,N_14622,N_14697);
or U15227 (N_15227,N_14706,N_14745);
nand U15228 (N_15228,N_14536,N_14294);
nand U15229 (N_15229,N_14225,N_14567);
or U15230 (N_15230,N_14926,N_14345);
nand U15231 (N_15231,N_14836,N_14555);
or U15232 (N_15232,N_14715,N_14776);
nand U15233 (N_15233,N_14951,N_14730);
nor U15234 (N_15234,N_14108,N_14796);
xnor U15235 (N_15235,N_14219,N_14429);
and U15236 (N_15236,N_14087,N_14464);
nand U15237 (N_15237,N_14178,N_14922);
xor U15238 (N_15238,N_14015,N_14719);
xor U15239 (N_15239,N_14832,N_14881);
xnor U15240 (N_15240,N_14152,N_14053);
or U15241 (N_15241,N_14683,N_14553);
and U15242 (N_15242,N_14765,N_14642);
and U15243 (N_15243,N_14385,N_14558);
or U15244 (N_15244,N_14548,N_14270);
and U15245 (N_15245,N_14200,N_14872);
nor U15246 (N_15246,N_14480,N_14371);
nor U15247 (N_15247,N_14791,N_14260);
nand U15248 (N_15248,N_14017,N_14437);
and U15249 (N_15249,N_14168,N_14476);
or U15250 (N_15250,N_14407,N_14772);
or U15251 (N_15251,N_14853,N_14898);
nor U15252 (N_15252,N_14386,N_14328);
and U15253 (N_15253,N_14736,N_14687);
or U15254 (N_15254,N_14754,N_14761);
and U15255 (N_15255,N_14784,N_14482);
nor U15256 (N_15256,N_14654,N_14300);
nor U15257 (N_15257,N_14904,N_14326);
nor U15258 (N_15258,N_14134,N_14415);
xor U15259 (N_15259,N_14580,N_14451);
nor U15260 (N_15260,N_14495,N_14283);
and U15261 (N_15261,N_14340,N_14769);
nand U15262 (N_15262,N_14900,N_14088);
and U15263 (N_15263,N_14408,N_14427);
and U15264 (N_15264,N_14885,N_14098);
or U15265 (N_15265,N_14804,N_14499);
or U15266 (N_15266,N_14037,N_14551);
or U15267 (N_15267,N_14076,N_14817);
nand U15268 (N_15268,N_14249,N_14879);
nor U15269 (N_15269,N_14239,N_14184);
or U15270 (N_15270,N_14397,N_14172);
nor U15271 (N_15271,N_14061,N_14128);
or U15272 (N_15272,N_14515,N_14032);
or U15273 (N_15273,N_14018,N_14324);
xnor U15274 (N_15274,N_14050,N_14315);
nor U15275 (N_15275,N_14728,N_14970);
and U15276 (N_15276,N_14301,N_14658);
nand U15277 (N_15277,N_14942,N_14644);
xor U15278 (N_15278,N_14993,N_14773);
nand U15279 (N_15279,N_14490,N_14263);
nand U15280 (N_15280,N_14447,N_14303);
or U15281 (N_15281,N_14468,N_14376);
nand U15282 (N_15282,N_14205,N_14201);
nand U15283 (N_15283,N_14366,N_14759);
nand U15284 (N_15284,N_14351,N_14974);
xor U15285 (N_15285,N_14481,N_14255);
or U15286 (N_15286,N_14981,N_14868);
xor U15287 (N_15287,N_14513,N_14533);
nand U15288 (N_15288,N_14711,N_14419);
or U15289 (N_15289,N_14170,N_14257);
nand U15290 (N_15290,N_14251,N_14159);
nand U15291 (N_15291,N_14944,N_14936);
or U15292 (N_15292,N_14360,N_14633);
nor U15293 (N_15293,N_14231,N_14610);
xnor U15294 (N_15294,N_14671,N_14054);
xor U15295 (N_15295,N_14275,N_14845);
and U15296 (N_15296,N_14570,N_14333);
nand U15297 (N_15297,N_14947,N_14151);
or U15298 (N_15298,N_14803,N_14673);
and U15299 (N_15299,N_14594,N_14431);
or U15300 (N_15300,N_14829,N_14235);
and U15301 (N_15301,N_14639,N_14691);
or U15302 (N_15302,N_14638,N_14071);
and U15303 (N_15303,N_14019,N_14065);
nor U15304 (N_15304,N_14492,N_14414);
nand U15305 (N_15305,N_14440,N_14147);
and U15306 (N_15306,N_14265,N_14969);
and U15307 (N_15307,N_14318,N_14902);
nand U15308 (N_15308,N_14295,N_14955);
nor U15309 (N_15309,N_14943,N_14937);
nand U15310 (N_15310,N_14261,N_14939);
nand U15311 (N_15311,N_14216,N_14739);
and U15312 (N_15312,N_14403,N_14521);
xor U15313 (N_15313,N_14707,N_14617);
and U15314 (N_15314,N_14312,N_14882);
and U15315 (N_15315,N_14355,N_14221);
xnor U15316 (N_15316,N_14732,N_14713);
xnor U15317 (N_15317,N_14023,N_14114);
xor U15318 (N_15318,N_14094,N_14228);
nand U15319 (N_15319,N_14971,N_14609);
nor U15320 (N_15320,N_14831,N_14770);
and U15321 (N_15321,N_14370,N_14457);
nand U15322 (N_15322,N_14271,N_14762);
xor U15323 (N_15323,N_14119,N_14606);
xnor U15324 (N_15324,N_14124,N_14935);
or U15325 (N_15325,N_14474,N_14643);
or U15326 (N_15326,N_14332,N_14404);
xnor U15327 (N_15327,N_14625,N_14999);
and U15328 (N_15328,N_14557,N_14095);
nand U15329 (N_15329,N_14811,N_14552);
nand U15330 (N_15330,N_14976,N_14986);
nand U15331 (N_15331,N_14177,N_14494);
xor U15332 (N_15332,N_14084,N_14635);
nor U15333 (N_15333,N_14189,N_14041);
nor U15334 (N_15334,N_14925,N_14387);
and U15335 (N_15335,N_14475,N_14560);
and U15336 (N_15336,N_14338,N_14428);
nor U15337 (N_15337,N_14749,N_14118);
nand U15338 (N_15338,N_14747,N_14768);
nor U15339 (N_15339,N_14244,N_14373);
or U15340 (N_15340,N_14672,N_14462);
xor U15341 (N_15341,N_14392,N_14727);
or U15342 (N_15342,N_14488,N_14895);
or U15343 (N_15343,N_14891,N_14975);
xnor U15344 (N_15344,N_14183,N_14336);
or U15345 (N_15345,N_14896,N_14813);
nor U15346 (N_15346,N_14002,N_14245);
xnor U15347 (N_15347,N_14568,N_14083);
xnor U15348 (N_15348,N_14846,N_14461);
or U15349 (N_15349,N_14556,N_14855);
and U15350 (N_15350,N_14740,N_14233);
or U15351 (N_15351,N_14851,N_14923);
xor U15352 (N_15352,N_14445,N_14887);
or U15353 (N_15353,N_14344,N_14543);
and U15354 (N_15354,N_14222,N_14204);
and U15355 (N_15355,N_14449,N_14357);
nor U15356 (N_15356,N_14915,N_14852);
nor U15357 (N_15357,N_14572,N_14025);
nand U15358 (N_15358,N_14422,N_14801);
nor U15359 (N_15359,N_14708,N_14302);
nor U15360 (N_15360,N_14841,N_14611);
and U15361 (N_15361,N_14648,N_14818);
xnor U15362 (N_15362,N_14870,N_14247);
or U15363 (N_15363,N_14931,N_14421);
xor U15364 (N_15364,N_14367,N_14800);
xor U15365 (N_15365,N_14439,N_14327);
and U15366 (N_15366,N_14797,N_14987);
nand U15367 (N_15367,N_14175,N_14090);
nand U15368 (N_15368,N_14919,N_14356);
or U15369 (N_15369,N_14651,N_14663);
nand U15370 (N_15370,N_14396,N_14914);
nor U15371 (N_15371,N_14933,N_14116);
nor U15372 (N_15372,N_14060,N_14106);
xnor U15373 (N_15373,N_14911,N_14775);
nor U15374 (N_15374,N_14814,N_14661);
or U15375 (N_15375,N_14767,N_14860);
xor U15376 (N_15376,N_14171,N_14182);
nand U15377 (N_15377,N_14875,N_14423);
and U15378 (N_15378,N_14929,N_14604);
xor U15379 (N_15379,N_14158,N_14484);
nand U15380 (N_15380,N_14839,N_14918);
nand U15381 (N_15381,N_14810,N_14957);
nand U15382 (N_15382,N_14905,N_14369);
nor U15383 (N_15383,N_14674,N_14562);
nand U15384 (N_15384,N_14838,N_14472);
nor U15385 (N_15385,N_14627,N_14916);
xnor U15386 (N_15386,N_14322,N_14522);
nor U15387 (N_15387,N_14048,N_14198);
or U15388 (N_15388,N_14487,N_14062);
nand U15389 (N_15389,N_14757,N_14489);
nand U15390 (N_15390,N_14068,N_14049);
or U15391 (N_15391,N_14894,N_14725);
xor U15392 (N_15392,N_14101,N_14819);
nor U15393 (N_15393,N_14460,N_14859);
nor U15394 (N_15394,N_14346,N_14744);
and U15395 (N_15395,N_14014,N_14523);
xnor U15396 (N_15396,N_14412,N_14790);
and U15397 (N_15397,N_14954,N_14500);
nand U15398 (N_15398,N_14692,N_14081);
xnor U15399 (N_15399,N_14840,N_14320);
or U15400 (N_15400,N_14723,N_14595);
nor U15401 (N_15401,N_14196,N_14581);
nand U15402 (N_15402,N_14511,N_14379);
nor U15403 (N_15403,N_14013,N_14998);
xnor U15404 (N_15404,N_14433,N_14181);
nor U15405 (N_15405,N_14400,N_14664);
nor U15406 (N_15406,N_14945,N_14650);
nand U15407 (N_15407,N_14347,N_14368);
nand U15408 (N_15408,N_14030,N_14505);
or U15409 (N_15409,N_14063,N_14258);
or U15410 (N_15410,N_14142,N_14613);
xnor U15411 (N_15411,N_14956,N_14331);
and U15412 (N_15412,N_14794,N_14193);
or U15413 (N_15413,N_14619,N_14304);
xnor U15414 (N_15414,N_14973,N_14632);
nor U15415 (N_15415,N_14213,N_14384);
xnor U15416 (N_15416,N_14569,N_14073);
nand U15417 (N_15417,N_14086,N_14893);
nor U15418 (N_15418,N_14055,N_14848);
nand U15419 (N_15419,N_14983,N_14417);
and U15420 (N_15420,N_14091,N_14267);
or U15421 (N_15421,N_14941,N_14535);
nor U15422 (N_15422,N_14284,N_14120);
and U15423 (N_15423,N_14162,N_14693);
nor U15424 (N_15424,N_14140,N_14666);
nand U15425 (N_15425,N_14608,N_14634);
xnor U15426 (N_15426,N_14698,N_14163);
xnor U15427 (N_15427,N_14583,N_14485);
nor U15428 (N_15428,N_14144,N_14812);
or U15429 (N_15429,N_14010,N_14329);
nand U15430 (N_15430,N_14372,N_14103);
nor U15431 (N_15431,N_14477,N_14034);
and U15432 (N_15432,N_14777,N_14785);
or U15433 (N_15433,N_14185,N_14519);
xor U15434 (N_15434,N_14465,N_14517);
and U15435 (N_15435,N_14123,N_14364);
nand U15436 (N_15436,N_14867,N_14137);
nand U15437 (N_15437,N_14040,N_14001);
xor U15438 (N_15438,N_14764,N_14652);
xnor U15439 (N_15439,N_14869,N_14647);
and U15440 (N_15440,N_14649,N_14645);
nand U15441 (N_15441,N_14291,N_14512);
nor U15442 (N_15442,N_14850,N_14362);
xor U15443 (N_15443,N_14659,N_14145);
xor U15444 (N_15444,N_14455,N_14690);
or U15445 (N_15445,N_14524,N_14722);
nand U15446 (N_15446,N_14721,N_14966);
nand U15447 (N_15447,N_14486,N_14350);
xnor U15448 (N_15448,N_14795,N_14277);
nor U15449 (N_15449,N_14884,N_14897);
nor U15450 (N_15450,N_14080,N_14843);
xnor U15451 (N_15451,N_14586,N_14753);
nand U15452 (N_15452,N_14434,N_14150);
xnor U15453 (N_15453,N_14920,N_14689);
nand U15454 (N_15454,N_14612,N_14637);
xnor U15455 (N_15455,N_14149,N_14031);
xor U15456 (N_15456,N_14424,N_14195);
xnor U15457 (N_15457,N_14677,N_14096);
nand U15458 (N_15458,N_14828,N_14682);
and U15459 (N_15459,N_14286,N_14074);
xnor U15460 (N_15460,N_14927,N_14921);
nor U15461 (N_15461,N_14339,N_14824);
or U15462 (N_15462,N_14426,N_14165);
nor U15463 (N_15463,N_14243,N_14342);
or U15464 (N_15464,N_14099,N_14377);
nor U15465 (N_15465,N_14641,N_14958);
and U15466 (N_15466,N_14924,N_14363);
and U15467 (N_15467,N_14456,N_14453);
xnor U15468 (N_15468,N_14254,N_14549);
xor U15469 (N_15469,N_14232,N_14735);
nand U15470 (N_15470,N_14226,N_14599);
xnor U15471 (N_15471,N_14737,N_14564);
and U15472 (N_15472,N_14888,N_14995);
xnor U15473 (N_15473,N_14133,N_14169);
and U15474 (N_15474,N_14250,N_14105);
and U15475 (N_15475,N_14262,N_14591);
nand U15476 (N_15476,N_14033,N_14886);
nor U15477 (N_15477,N_14577,N_14630);
or U15478 (N_15478,N_14863,N_14479);
and U15479 (N_15479,N_14760,N_14518);
nor U15480 (N_15480,N_14880,N_14509);
xor U15481 (N_15481,N_14876,N_14459);
xnor U15482 (N_15482,N_14003,N_14153);
xor U15483 (N_15483,N_14704,N_14539);
and U15484 (N_15484,N_14280,N_14675);
nand U15485 (N_15485,N_14199,N_14045);
xnor U15486 (N_15486,N_14590,N_14131);
xor U15487 (N_15487,N_14246,N_14104);
nor U15488 (N_15488,N_14354,N_14343);
nor U15489 (N_15489,N_14278,N_14004);
nor U15490 (N_15490,N_14788,N_14626);
or U15491 (N_15491,N_14750,N_14605);
nor U15492 (N_15492,N_14636,N_14361);
nor U15493 (N_15493,N_14154,N_14968);
nand U15494 (N_15494,N_14416,N_14498);
nor U15495 (N_15495,N_14779,N_14588);
xnor U15496 (N_15496,N_14028,N_14334);
nor U15497 (N_15497,N_14702,N_14616);
nand U15498 (N_15498,N_14994,N_14473);
xor U15499 (N_15499,N_14349,N_14861);
nor U15500 (N_15500,N_14716,N_14892);
or U15501 (N_15501,N_14695,N_14211);
or U15502 (N_15502,N_14669,N_14161);
or U15503 (N_15503,N_14044,N_14952);
nand U15504 (N_15504,N_14042,N_14283);
and U15505 (N_15505,N_14009,N_14361);
and U15506 (N_15506,N_14751,N_14900);
nand U15507 (N_15507,N_14891,N_14309);
xor U15508 (N_15508,N_14034,N_14150);
nor U15509 (N_15509,N_14365,N_14728);
xnor U15510 (N_15510,N_14131,N_14408);
and U15511 (N_15511,N_14870,N_14522);
or U15512 (N_15512,N_14588,N_14098);
nand U15513 (N_15513,N_14026,N_14464);
or U15514 (N_15514,N_14684,N_14908);
and U15515 (N_15515,N_14681,N_14651);
nor U15516 (N_15516,N_14345,N_14453);
and U15517 (N_15517,N_14278,N_14417);
or U15518 (N_15518,N_14929,N_14534);
and U15519 (N_15519,N_14184,N_14483);
and U15520 (N_15520,N_14275,N_14151);
nand U15521 (N_15521,N_14501,N_14316);
and U15522 (N_15522,N_14430,N_14346);
nor U15523 (N_15523,N_14887,N_14690);
nor U15524 (N_15524,N_14352,N_14303);
nor U15525 (N_15525,N_14194,N_14486);
and U15526 (N_15526,N_14691,N_14230);
nor U15527 (N_15527,N_14579,N_14392);
xor U15528 (N_15528,N_14033,N_14640);
nand U15529 (N_15529,N_14334,N_14359);
nor U15530 (N_15530,N_14786,N_14769);
nand U15531 (N_15531,N_14389,N_14767);
nor U15532 (N_15532,N_14462,N_14282);
and U15533 (N_15533,N_14597,N_14946);
or U15534 (N_15534,N_14820,N_14005);
or U15535 (N_15535,N_14976,N_14837);
nand U15536 (N_15536,N_14448,N_14723);
or U15537 (N_15537,N_14671,N_14124);
xnor U15538 (N_15538,N_14476,N_14154);
nor U15539 (N_15539,N_14466,N_14473);
or U15540 (N_15540,N_14629,N_14774);
nand U15541 (N_15541,N_14810,N_14762);
xor U15542 (N_15542,N_14773,N_14265);
nor U15543 (N_15543,N_14158,N_14016);
nor U15544 (N_15544,N_14689,N_14401);
nand U15545 (N_15545,N_14149,N_14289);
and U15546 (N_15546,N_14420,N_14113);
xor U15547 (N_15547,N_14284,N_14538);
xor U15548 (N_15548,N_14812,N_14637);
nor U15549 (N_15549,N_14082,N_14338);
or U15550 (N_15550,N_14844,N_14941);
nor U15551 (N_15551,N_14236,N_14957);
and U15552 (N_15552,N_14992,N_14866);
nor U15553 (N_15553,N_14929,N_14971);
xor U15554 (N_15554,N_14624,N_14886);
nor U15555 (N_15555,N_14590,N_14342);
nand U15556 (N_15556,N_14514,N_14232);
and U15557 (N_15557,N_14646,N_14287);
nand U15558 (N_15558,N_14130,N_14509);
and U15559 (N_15559,N_14061,N_14325);
xor U15560 (N_15560,N_14799,N_14506);
nor U15561 (N_15561,N_14375,N_14246);
nand U15562 (N_15562,N_14198,N_14505);
or U15563 (N_15563,N_14723,N_14933);
xor U15564 (N_15564,N_14655,N_14363);
and U15565 (N_15565,N_14984,N_14846);
nand U15566 (N_15566,N_14206,N_14568);
xnor U15567 (N_15567,N_14416,N_14624);
nand U15568 (N_15568,N_14640,N_14324);
nand U15569 (N_15569,N_14363,N_14898);
or U15570 (N_15570,N_14328,N_14223);
xnor U15571 (N_15571,N_14471,N_14970);
xor U15572 (N_15572,N_14120,N_14267);
xor U15573 (N_15573,N_14295,N_14713);
nor U15574 (N_15574,N_14184,N_14265);
or U15575 (N_15575,N_14759,N_14117);
or U15576 (N_15576,N_14880,N_14341);
and U15577 (N_15577,N_14777,N_14801);
nand U15578 (N_15578,N_14759,N_14420);
nand U15579 (N_15579,N_14724,N_14764);
and U15580 (N_15580,N_14328,N_14339);
nor U15581 (N_15581,N_14653,N_14727);
xnor U15582 (N_15582,N_14224,N_14324);
nand U15583 (N_15583,N_14486,N_14278);
or U15584 (N_15584,N_14021,N_14116);
xor U15585 (N_15585,N_14245,N_14465);
nand U15586 (N_15586,N_14299,N_14217);
nor U15587 (N_15587,N_14099,N_14957);
and U15588 (N_15588,N_14815,N_14001);
or U15589 (N_15589,N_14387,N_14468);
and U15590 (N_15590,N_14465,N_14280);
or U15591 (N_15591,N_14984,N_14206);
nand U15592 (N_15592,N_14169,N_14058);
nand U15593 (N_15593,N_14907,N_14268);
nor U15594 (N_15594,N_14336,N_14956);
and U15595 (N_15595,N_14756,N_14917);
xnor U15596 (N_15596,N_14742,N_14621);
or U15597 (N_15597,N_14595,N_14337);
nand U15598 (N_15598,N_14275,N_14066);
xnor U15599 (N_15599,N_14908,N_14576);
or U15600 (N_15600,N_14992,N_14186);
xnor U15601 (N_15601,N_14015,N_14640);
nand U15602 (N_15602,N_14252,N_14608);
xnor U15603 (N_15603,N_14600,N_14371);
nor U15604 (N_15604,N_14778,N_14000);
xnor U15605 (N_15605,N_14139,N_14491);
and U15606 (N_15606,N_14778,N_14733);
xnor U15607 (N_15607,N_14960,N_14666);
xor U15608 (N_15608,N_14710,N_14538);
nor U15609 (N_15609,N_14772,N_14192);
or U15610 (N_15610,N_14738,N_14722);
or U15611 (N_15611,N_14503,N_14552);
and U15612 (N_15612,N_14166,N_14847);
xor U15613 (N_15613,N_14557,N_14647);
or U15614 (N_15614,N_14009,N_14298);
nor U15615 (N_15615,N_14346,N_14206);
nor U15616 (N_15616,N_14951,N_14760);
xnor U15617 (N_15617,N_14636,N_14473);
xor U15618 (N_15618,N_14460,N_14998);
nor U15619 (N_15619,N_14702,N_14436);
xnor U15620 (N_15620,N_14012,N_14412);
xnor U15621 (N_15621,N_14634,N_14850);
nand U15622 (N_15622,N_14243,N_14677);
nor U15623 (N_15623,N_14862,N_14568);
and U15624 (N_15624,N_14237,N_14228);
or U15625 (N_15625,N_14695,N_14137);
xnor U15626 (N_15626,N_14205,N_14694);
or U15627 (N_15627,N_14829,N_14450);
or U15628 (N_15628,N_14137,N_14755);
xnor U15629 (N_15629,N_14693,N_14802);
nor U15630 (N_15630,N_14193,N_14905);
and U15631 (N_15631,N_14372,N_14788);
or U15632 (N_15632,N_14037,N_14309);
or U15633 (N_15633,N_14717,N_14146);
nor U15634 (N_15634,N_14819,N_14261);
nand U15635 (N_15635,N_14710,N_14849);
and U15636 (N_15636,N_14427,N_14288);
nor U15637 (N_15637,N_14708,N_14467);
or U15638 (N_15638,N_14291,N_14905);
or U15639 (N_15639,N_14471,N_14801);
nor U15640 (N_15640,N_14481,N_14731);
or U15641 (N_15641,N_14631,N_14456);
and U15642 (N_15642,N_14180,N_14333);
and U15643 (N_15643,N_14246,N_14684);
or U15644 (N_15644,N_14341,N_14429);
or U15645 (N_15645,N_14408,N_14366);
nand U15646 (N_15646,N_14953,N_14769);
nand U15647 (N_15647,N_14561,N_14751);
nor U15648 (N_15648,N_14848,N_14743);
xor U15649 (N_15649,N_14553,N_14294);
nor U15650 (N_15650,N_14885,N_14533);
xor U15651 (N_15651,N_14163,N_14007);
or U15652 (N_15652,N_14885,N_14399);
xor U15653 (N_15653,N_14863,N_14491);
and U15654 (N_15654,N_14038,N_14268);
or U15655 (N_15655,N_14598,N_14325);
nand U15656 (N_15656,N_14825,N_14945);
nand U15657 (N_15657,N_14586,N_14082);
nor U15658 (N_15658,N_14212,N_14729);
xor U15659 (N_15659,N_14172,N_14232);
xnor U15660 (N_15660,N_14058,N_14945);
xor U15661 (N_15661,N_14479,N_14907);
nand U15662 (N_15662,N_14567,N_14413);
or U15663 (N_15663,N_14084,N_14657);
nand U15664 (N_15664,N_14365,N_14586);
and U15665 (N_15665,N_14931,N_14479);
or U15666 (N_15666,N_14883,N_14245);
xnor U15667 (N_15667,N_14963,N_14494);
nand U15668 (N_15668,N_14257,N_14453);
nor U15669 (N_15669,N_14388,N_14769);
xor U15670 (N_15670,N_14555,N_14974);
and U15671 (N_15671,N_14994,N_14980);
nand U15672 (N_15672,N_14836,N_14693);
nand U15673 (N_15673,N_14452,N_14468);
nand U15674 (N_15674,N_14284,N_14508);
nor U15675 (N_15675,N_14850,N_14983);
xor U15676 (N_15676,N_14476,N_14246);
nand U15677 (N_15677,N_14495,N_14196);
nand U15678 (N_15678,N_14527,N_14456);
and U15679 (N_15679,N_14141,N_14904);
nor U15680 (N_15680,N_14383,N_14006);
or U15681 (N_15681,N_14661,N_14955);
or U15682 (N_15682,N_14724,N_14523);
xnor U15683 (N_15683,N_14980,N_14354);
and U15684 (N_15684,N_14803,N_14170);
nand U15685 (N_15685,N_14871,N_14499);
nor U15686 (N_15686,N_14385,N_14830);
nor U15687 (N_15687,N_14624,N_14117);
nand U15688 (N_15688,N_14530,N_14120);
or U15689 (N_15689,N_14230,N_14086);
or U15690 (N_15690,N_14309,N_14018);
or U15691 (N_15691,N_14980,N_14158);
nand U15692 (N_15692,N_14543,N_14580);
nand U15693 (N_15693,N_14483,N_14820);
xnor U15694 (N_15694,N_14890,N_14148);
and U15695 (N_15695,N_14576,N_14939);
and U15696 (N_15696,N_14979,N_14928);
and U15697 (N_15697,N_14025,N_14005);
or U15698 (N_15698,N_14452,N_14802);
nor U15699 (N_15699,N_14041,N_14001);
nand U15700 (N_15700,N_14575,N_14565);
or U15701 (N_15701,N_14271,N_14300);
or U15702 (N_15702,N_14548,N_14924);
nor U15703 (N_15703,N_14035,N_14461);
and U15704 (N_15704,N_14372,N_14573);
xor U15705 (N_15705,N_14250,N_14338);
or U15706 (N_15706,N_14761,N_14021);
or U15707 (N_15707,N_14417,N_14987);
and U15708 (N_15708,N_14144,N_14919);
and U15709 (N_15709,N_14389,N_14966);
nor U15710 (N_15710,N_14366,N_14487);
and U15711 (N_15711,N_14938,N_14244);
and U15712 (N_15712,N_14271,N_14725);
or U15713 (N_15713,N_14126,N_14021);
xor U15714 (N_15714,N_14455,N_14861);
nor U15715 (N_15715,N_14865,N_14371);
nor U15716 (N_15716,N_14896,N_14739);
or U15717 (N_15717,N_14116,N_14518);
or U15718 (N_15718,N_14284,N_14025);
or U15719 (N_15719,N_14695,N_14079);
nor U15720 (N_15720,N_14992,N_14924);
nand U15721 (N_15721,N_14069,N_14729);
or U15722 (N_15722,N_14934,N_14020);
or U15723 (N_15723,N_14342,N_14281);
nand U15724 (N_15724,N_14570,N_14703);
nand U15725 (N_15725,N_14280,N_14211);
nand U15726 (N_15726,N_14883,N_14651);
or U15727 (N_15727,N_14083,N_14414);
and U15728 (N_15728,N_14489,N_14136);
nand U15729 (N_15729,N_14894,N_14927);
and U15730 (N_15730,N_14168,N_14097);
xor U15731 (N_15731,N_14972,N_14883);
xnor U15732 (N_15732,N_14816,N_14286);
xnor U15733 (N_15733,N_14319,N_14183);
and U15734 (N_15734,N_14331,N_14881);
xnor U15735 (N_15735,N_14628,N_14258);
nand U15736 (N_15736,N_14554,N_14967);
nor U15737 (N_15737,N_14354,N_14804);
nand U15738 (N_15738,N_14519,N_14852);
xnor U15739 (N_15739,N_14719,N_14670);
nor U15740 (N_15740,N_14863,N_14563);
nand U15741 (N_15741,N_14724,N_14085);
xnor U15742 (N_15742,N_14033,N_14873);
nor U15743 (N_15743,N_14131,N_14223);
nor U15744 (N_15744,N_14915,N_14958);
xnor U15745 (N_15745,N_14194,N_14870);
nand U15746 (N_15746,N_14832,N_14819);
or U15747 (N_15747,N_14559,N_14495);
nor U15748 (N_15748,N_14726,N_14502);
or U15749 (N_15749,N_14908,N_14122);
nor U15750 (N_15750,N_14362,N_14521);
nand U15751 (N_15751,N_14106,N_14337);
or U15752 (N_15752,N_14982,N_14700);
and U15753 (N_15753,N_14060,N_14412);
nor U15754 (N_15754,N_14340,N_14107);
nor U15755 (N_15755,N_14882,N_14611);
nor U15756 (N_15756,N_14940,N_14528);
nand U15757 (N_15757,N_14543,N_14260);
and U15758 (N_15758,N_14742,N_14461);
nand U15759 (N_15759,N_14165,N_14956);
nand U15760 (N_15760,N_14057,N_14976);
nor U15761 (N_15761,N_14006,N_14998);
nor U15762 (N_15762,N_14749,N_14115);
or U15763 (N_15763,N_14093,N_14052);
nand U15764 (N_15764,N_14016,N_14305);
xnor U15765 (N_15765,N_14643,N_14211);
nor U15766 (N_15766,N_14417,N_14622);
and U15767 (N_15767,N_14979,N_14429);
and U15768 (N_15768,N_14372,N_14269);
xnor U15769 (N_15769,N_14989,N_14550);
nand U15770 (N_15770,N_14076,N_14243);
xnor U15771 (N_15771,N_14463,N_14350);
xnor U15772 (N_15772,N_14279,N_14053);
and U15773 (N_15773,N_14019,N_14128);
or U15774 (N_15774,N_14375,N_14180);
and U15775 (N_15775,N_14030,N_14734);
xor U15776 (N_15776,N_14336,N_14495);
or U15777 (N_15777,N_14028,N_14188);
xor U15778 (N_15778,N_14097,N_14496);
and U15779 (N_15779,N_14716,N_14765);
nor U15780 (N_15780,N_14545,N_14596);
nor U15781 (N_15781,N_14297,N_14590);
nand U15782 (N_15782,N_14599,N_14310);
or U15783 (N_15783,N_14750,N_14670);
and U15784 (N_15784,N_14949,N_14142);
nor U15785 (N_15785,N_14953,N_14709);
xor U15786 (N_15786,N_14258,N_14294);
and U15787 (N_15787,N_14573,N_14867);
and U15788 (N_15788,N_14100,N_14239);
xnor U15789 (N_15789,N_14536,N_14621);
nor U15790 (N_15790,N_14647,N_14914);
nand U15791 (N_15791,N_14413,N_14227);
and U15792 (N_15792,N_14704,N_14420);
or U15793 (N_15793,N_14957,N_14921);
nand U15794 (N_15794,N_14574,N_14216);
nand U15795 (N_15795,N_14298,N_14164);
nand U15796 (N_15796,N_14298,N_14092);
xnor U15797 (N_15797,N_14480,N_14736);
or U15798 (N_15798,N_14667,N_14628);
xnor U15799 (N_15799,N_14299,N_14598);
or U15800 (N_15800,N_14768,N_14777);
nand U15801 (N_15801,N_14933,N_14587);
xor U15802 (N_15802,N_14663,N_14198);
nand U15803 (N_15803,N_14364,N_14444);
nor U15804 (N_15804,N_14687,N_14392);
nor U15805 (N_15805,N_14625,N_14721);
xor U15806 (N_15806,N_14505,N_14124);
xnor U15807 (N_15807,N_14494,N_14308);
nor U15808 (N_15808,N_14489,N_14264);
and U15809 (N_15809,N_14063,N_14182);
and U15810 (N_15810,N_14580,N_14491);
nand U15811 (N_15811,N_14017,N_14927);
xnor U15812 (N_15812,N_14293,N_14250);
nor U15813 (N_15813,N_14576,N_14366);
xor U15814 (N_15814,N_14000,N_14228);
xor U15815 (N_15815,N_14068,N_14562);
xor U15816 (N_15816,N_14964,N_14743);
or U15817 (N_15817,N_14226,N_14058);
nor U15818 (N_15818,N_14424,N_14937);
and U15819 (N_15819,N_14550,N_14238);
or U15820 (N_15820,N_14714,N_14652);
nand U15821 (N_15821,N_14543,N_14035);
nor U15822 (N_15822,N_14331,N_14435);
xor U15823 (N_15823,N_14231,N_14426);
or U15824 (N_15824,N_14430,N_14917);
xnor U15825 (N_15825,N_14300,N_14525);
nand U15826 (N_15826,N_14139,N_14869);
and U15827 (N_15827,N_14028,N_14415);
xnor U15828 (N_15828,N_14994,N_14858);
xnor U15829 (N_15829,N_14797,N_14383);
nor U15830 (N_15830,N_14425,N_14900);
xor U15831 (N_15831,N_14708,N_14489);
nand U15832 (N_15832,N_14157,N_14295);
and U15833 (N_15833,N_14573,N_14106);
xnor U15834 (N_15834,N_14747,N_14112);
and U15835 (N_15835,N_14665,N_14549);
xnor U15836 (N_15836,N_14038,N_14853);
xnor U15837 (N_15837,N_14666,N_14529);
xnor U15838 (N_15838,N_14428,N_14384);
or U15839 (N_15839,N_14153,N_14853);
or U15840 (N_15840,N_14528,N_14384);
nor U15841 (N_15841,N_14541,N_14477);
and U15842 (N_15842,N_14094,N_14449);
nor U15843 (N_15843,N_14815,N_14620);
nor U15844 (N_15844,N_14673,N_14826);
xor U15845 (N_15845,N_14755,N_14185);
nor U15846 (N_15846,N_14585,N_14761);
or U15847 (N_15847,N_14299,N_14187);
or U15848 (N_15848,N_14219,N_14596);
and U15849 (N_15849,N_14757,N_14761);
nand U15850 (N_15850,N_14783,N_14205);
nand U15851 (N_15851,N_14946,N_14458);
nor U15852 (N_15852,N_14172,N_14175);
nand U15853 (N_15853,N_14839,N_14149);
and U15854 (N_15854,N_14403,N_14428);
xnor U15855 (N_15855,N_14602,N_14244);
xnor U15856 (N_15856,N_14744,N_14650);
and U15857 (N_15857,N_14148,N_14411);
xor U15858 (N_15858,N_14972,N_14811);
and U15859 (N_15859,N_14584,N_14848);
or U15860 (N_15860,N_14546,N_14097);
and U15861 (N_15861,N_14544,N_14596);
xnor U15862 (N_15862,N_14334,N_14433);
xor U15863 (N_15863,N_14435,N_14880);
and U15864 (N_15864,N_14208,N_14632);
or U15865 (N_15865,N_14088,N_14764);
nor U15866 (N_15866,N_14573,N_14127);
nor U15867 (N_15867,N_14354,N_14003);
or U15868 (N_15868,N_14061,N_14056);
nand U15869 (N_15869,N_14543,N_14275);
xnor U15870 (N_15870,N_14666,N_14803);
nor U15871 (N_15871,N_14650,N_14915);
nor U15872 (N_15872,N_14387,N_14449);
or U15873 (N_15873,N_14983,N_14048);
xnor U15874 (N_15874,N_14948,N_14393);
nand U15875 (N_15875,N_14855,N_14630);
nand U15876 (N_15876,N_14525,N_14121);
or U15877 (N_15877,N_14265,N_14336);
nor U15878 (N_15878,N_14686,N_14544);
or U15879 (N_15879,N_14597,N_14900);
xor U15880 (N_15880,N_14568,N_14062);
or U15881 (N_15881,N_14562,N_14310);
and U15882 (N_15882,N_14673,N_14716);
nand U15883 (N_15883,N_14441,N_14346);
and U15884 (N_15884,N_14348,N_14152);
nand U15885 (N_15885,N_14274,N_14231);
nand U15886 (N_15886,N_14939,N_14191);
and U15887 (N_15887,N_14018,N_14420);
nor U15888 (N_15888,N_14043,N_14676);
xor U15889 (N_15889,N_14258,N_14113);
and U15890 (N_15890,N_14529,N_14707);
and U15891 (N_15891,N_14439,N_14740);
nand U15892 (N_15892,N_14898,N_14931);
or U15893 (N_15893,N_14879,N_14668);
xor U15894 (N_15894,N_14428,N_14520);
nand U15895 (N_15895,N_14897,N_14621);
or U15896 (N_15896,N_14602,N_14484);
nand U15897 (N_15897,N_14445,N_14671);
nor U15898 (N_15898,N_14722,N_14170);
xnor U15899 (N_15899,N_14909,N_14983);
xnor U15900 (N_15900,N_14026,N_14730);
and U15901 (N_15901,N_14061,N_14941);
nor U15902 (N_15902,N_14153,N_14591);
nand U15903 (N_15903,N_14436,N_14551);
nor U15904 (N_15904,N_14140,N_14221);
nor U15905 (N_15905,N_14473,N_14491);
nor U15906 (N_15906,N_14027,N_14880);
xnor U15907 (N_15907,N_14371,N_14030);
nor U15908 (N_15908,N_14467,N_14490);
or U15909 (N_15909,N_14379,N_14407);
and U15910 (N_15910,N_14713,N_14448);
xor U15911 (N_15911,N_14442,N_14313);
and U15912 (N_15912,N_14172,N_14849);
xor U15913 (N_15913,N_14516,N_14662);
nor U15914 (N_15914,N_14347,N_14195);
nand U15915 (N_15915,N_14078,N_14941);
nor U15916 (N_15916,N_14485,N_14275);
nand U15917 (N_15917,N_14647,N_14231);
nand U15918 (N_15918,N_14347,N_14385);
or U15919 (N_15919,N_14771,N_14370);
nor U15920 (N_15920,N_14073,N_14717);
nand U15921 (N_15921,N_14801,N_14268);
and U15922 (N_15922,N_14034,N_14162);
nand U15923 (N_15923,N_14322,N_14923);
nand U15924 (N_15924,N_14965,N_14249);
xnor U15925 (N_15925,N_14855,N_14875);
or U15926 (N_15926,N_14202,N_14257);
xnor U15927 (N_15927,N_14334,N_14613);
nor U15928 (N_15928,N_14341,N_14791);
or U15929 (N_15929,N_14816,N_14224);
nand U15930 (N_15930,N_14068,N_14491);
nor U15931 (N_15931,N_14765,N_14634);
nor U15932 (N_15932,N_14448,N_14297);
and U15933 (N_15933,N_14543,N_14794);
or U15934 (N_15934,N_14615,N_14778);
xor U15935 (N_15935,N_14881,N_14019);
and U15936 (N_15936,N_14725,N_14872);
or U15937 (N_15937,N_14445,N_14177);
xor U15938 (N_15938,N_14937,N_14414);
nand U15939 (N_15939,N_14884,N_14080);
and U15940 (N_15940,N_14549,N_14205);
nand U15941 (N_15941,N_14539,N_14077);
nand U15942 (N_15942,N_14747,N_14159);
xor U15943 (N_15943,N_14086,N_14078);
xnor U15944 (N_15944,N_14863,N_14456);
nand U15945 (N_15945,N_14823,N_14668);
nand U15946 (N_15946,N_14018,N_14963);
and U15947 (N_15947,N_14064,N_14110);
or U15948 (N_15948,N_14268,N_14681);
nor U15949 (N_15949,N_14463,N_14941);
nand U15950 (N_15950,N_14450,N_14245);
or U15951 (N_15951,N_14487,N_14194);
and U15952 (N_15952,N_14921,N_14339);
xor U15953 (N_15953,N_14471,N_14078);
or U15954 (N_15954,N_14453,N_14530);
or U15955 (N_15955,N_14014,N_14321);
and U15956 (N_15956,N_14260,N_14493);
nand U15957 (N_15957,N_14602,N_14745);
xor U15958 (N_15958,N_14509,N_14665);
nand U15959 (N_15959,N_14264,N_14200);
nor U15960 (N_15960,N_14236,N_14059);
nor U15961 (N_15961,N_14398,N_14720);
xnor U15962 (N_15962,N_14934,N_14945);
or U15963 (N_15963,N_14151,N_14553);
nor U15964 (N_15964,N_14596,N_14800);
nor U15965 (N_15965,N_14842,N_14883);
or U15966 (N_15966,N_14106,N_14223);
nor U15967 (N_15967,N_14239,N_14218);
nor U15968 (N_15968,N_14575,N_14628);
nor U15969 (N_15969,N_14635,N_14232);
nand U15970 (N_15970,N_14495,N_14322);
nor U15971 (N_15971,N_14840,N_14381);
xor U15972 (N_15972,N_14512,N_14219);
nor U15973 (N_15973,N_14891,N_14398);
nor U15974 (N_15974,N_14537,N_14901);
or U15975 (N_15975,N_14313,N_14819);
or U15976 (N_15976,N_14179,N_14030);
nand U15977 (N_15977,N_14996,N_14239);
nor U15978 (N_15978,N_14708,N_14904);
nand U15979 (N_15979,N_14592,N_14837);
and U15980 (N_15980,N_14070,N_14460);
nor U15981 (N_15981,N_14422,N_14344);
and U15982 (N_15982,N_14547,N_14294);
nand U15983 (N_15983,N_14489,N_14226);
and U15984 (N_15984,N_14276,N_14115);
nand U15985 (N_15985,N_14745,N_14950);
nor U15986 (N_15986,N_14035,N_14531);
xor U15987 (N_15987,N_14371,N_14586);
or U15988 (N_15988,N_14504,N_14126);
or U15989 (N_15989,N_14959,N_14559);
and U15990 (N_15990,N_14236,N_14364);
or U15991 (N_15991,N_14335,N_14266);
or U15992 (N_15992,N_14139,N_14430);
and U15993 (N_15993,N_14781,N_14025);
nand U15994 (N_15994,N_14473,N_14920);
nor U15995 (N_15995,N_14920,N_14324);
and U15996 (N_15996,N_14997,N_14934);
nand U15997 (N_15997,N_14721,N_14251);
xnor U15998 (N_15998,N_14989,N_14781);
or U15999 (N_15999,N_14402,N_14461);
xor U16000 (N_16000,N_15173,N_15437);
and U16001 (N_16001,N_15561,N_15078);
and U16002 (N_16002,N_15762,N_15274);
xor U16003 (N_16003,N_15519,N_15029);
xnor U16004 (N_16004,N_15421,N_15791);
nand U16005 (N_16005,N_15592,N_15833);
nand U16006 (N_16006,N_15272,N_15027);
or U16007 (N_16007,N_15244,N_15972);
nor U16008 (N_16008,N_15706,N_15373);
nor U16009 (N_16009,N_15821,N_15179);
and U16010 (N_16010,N_15966,N_15683);
nand U16011 (N_16011,N_15948,N_15451);
nand U16012 (N_16012,N_15379,N_15709);
or U16013 (N_16013,N_15154,N_15792);
xnor U16014 (N_16014,N_15215,N_15284);
xor U16015 (N_16015,N_15168,N_15465);
nand U16016 (N_16016,N_15603,N_15739);
nand U16017 (N_16017,N_15780,N_15692);
and U16018 (N_16018,N_15193,N_15130);
or U16019 (N_16019,N_15288,N_15461);
or U16020 (N_16020,N_15090,N_15488);
xor U16021 (N_16021,N_15329,N_15482);
or U16022 (N_16022,N_15336,N_15365);
nand U16023 (N_16023,N_15197,N_15449);
and U16024 (N_16024,N_15162,N_15563);
nand U16025 (N_16025,N_15270,N_15467);
or U16026 (N_16026,N_15656,N_15546);
nor U16027 (N_16027,N_15832,N_15909);
and U16028 (N_16028,N_15504,N_15915);
and U16029 (N_16029,N_15797,N_15899);
nor U16030 (N_16030,N_15898,N_15030);
and U16031 (N_16031,N_15978,N_15590);
or U16032 (N_16032,N_15399,N_15132);
nor U16033 (N_16033,N_15069,N_15572);
and U16034 (N_16034,N_15655,N_15989);
and U16035 (N_16035,N_15033,N_15633);
and U16036 (N_16036,N_15190,N_15887);
xor U16037 (N_16037,N_15153,N_15850);
and U16038 (N_16038,N_15549,N_15089);
or U16039 (N_16039,N_15388,N_15851);
nand U16040 (N_16040,N_15494,N_15386);
nor U16041 (N_16041,N_15072,N_15144);
or U16042 (N_16042,N_15218,N_15836);
and U16043 (N_16043,N_15847,N_15216);
nand U16044 (N_16044,N_15729,N_15790);
and U16045 (N_16045,N_15105,N_15106);
or U16046 (N_16046,N_15439,N_15026);
nor U16047 (N_16047,N_15375,N_15536);
nor U16048 (N_16048,N_15834,N_15827);
nand U16049 (N_16049,N_15621,N_15707);
and U16050 (N_16050,N_15844,N_15586);
and U16051 (N_16051,N_15010,N_15472);
nor U16052 (N_16052,N_15974,N_15508);
or U16053 (N_16053,N_15092,N_15685);
xor U16054 (N_16054,N_15309,N_15903);
or U16055 (N_16055,N_15073,N_15347);
and U16056 (N_16056,N_15487,N_15798);
nand U16057 (N_16057,N_15538,N_15318);
and U16058 (N_16058,N_15061,N_15083);
and U16059 (N_16059,N_15265,N_15865);
nor U16060 (N_16060,N_15734,N_15659);
xor U16061 (N_16061,N_15870,N_15484);
nor U16062 (N_16062,N_15743,N_15455);
nand U16063 (N_16063,N_15943,N_15940);
and U16064 (N_16064,N_15250,N_15941);
nor U16065 (N_16065,N_15404,N_15977);
and U16066 (N_16066,N_15378,N_15102);
xnor U16067 (N_16067,N_15766,N_15861);
or U16068 (N_16068,N_15917,N_15161);
xnor U16069 (N_16069,N_15891,N_15335);
and U16070 (N_16070,N_15169,N_15890);
xor U16071 (N_16071,N_15624,N_15242);
xor U16072 (N_16072,N_15142,N_15885);
nor U16073 (N_16073,N_15584,N_15376);
and U16074 (N_16074,N_15846,N_15098);
and U16075 (N_16075,N_15372,N_15160);
or U16076 (N_16076,N_15393,N_15704);
nor U16077 (N_16077,N_15327,N_15413);
and U16078 (N_16078,N_15280,N_15279);
nor U16079 (N_16079,N_15454,N_15658);
xor U16080 (N_16080,N_15104,N_15814);
nor U16081 (N_16081,N_15911,N_15959);
and U16082 (N_16082,N_15431,N_15875);
and U16083 (N_16083,N_15062,N_15390);
nand U16084 (N_16084,N_15093,N_15843);
nand U16085 (N_16085,N_15637,N_15053);
nand U16086 (N_16086,N_15323,N_15298);
xnor U16087 (N_16087,N_15096,N_15261);
or U16088 (N_16088,N_15294,N_15511);
nor U16089 (N_16089,N_15634,N_15680);
nor U16090 (N_16090,N_15320,N_15363);
xnor U16091 (N_16091,N_15855,N_15411);
and U16092 (N_16092,N_15246,N_15292);
or U16093 (N_16093,N_15016,N_15183);
and U16094 (N_16094,N_15001,N_15587);
xor U16095 (N_16095,N_15570,N_15579);
and U16096 (N_16096,N_15693,N_15551);
or U16097 (N_16097,N_15207,N_15585);
and U16098 (N_16098,N_15632,N_15651);
xor U16099 (N_16099,N_15969,N_15631);
and U16100 (N_16100,N_15604,N_15992);
or U16101 (N_16101,N_15512,N_15949);
nand U16102 (N_16102,N_15297,N_15815);
or U16103 (N_16103,N_15853,N_15353);
or U16104 (N_16104,N_15740,N_15781);
xor U16105 (N_16105,N_15123,N_15236);
nor U16106 (N_16106,N_15965,N_15448);
and U16107 (N_16107,N_15471,N_15937);
nor U16108 (N_16108,N_15406,N_15492);
nand U16109 (N_16109,N_15023,N_15559);
and U16110 (N_16110,N_15436,N_15548);
nor U16111 (N_16111,N_15533,N_15984);
nand U16112 (N_16112,N_15702,N_15573);
xnor U16113 (N_16113,N_15237,N_15477);
xnor U16114 (N_16114,N_15800,N_15896);
and U16115 (N_16115,N_15313,N_15607);
and U16116 (N_16116,N_15883,N_15809);
and U16117 (N_16117,N_15211,N_15761);
nand U16118 (N_16118,N_15126,N_15922);
xor U16119 (N_16119,N_15750,N_15565);
or U16120 (N_16120,N_15295,N_15979);
xnor U16121 (N_16121,N_15269,N_15352);
and U16122 (N_16122,N_15470,N_15544);
nor U16123 (N_16123,N_15934,N_15332);
nand U16124 (N_16124,N_15418,N_15227);
xnor U16125 (N_16125,N_15907,N_15071);
or U16126 (N_16126,N_15498,N_15485);
and U16127 (N_16127,N_15793,N_15860);
xor U16128 (N_16128,N_15524,N_15755);
nor U16129 (N_16129,N_15645,N_15121);
nor U16130 (N_16130,N_15003,N_15848);
and U16131 (N_16131,N_15321,N_15080);
xor U16132 (N_16132,N_15505,N_15688);
xnor U16133 (N_16133,N_15159,N_15194);
and U16134 (N_16134,N_15474,N_15869);
nor U16135 (N_16135,N_15356,N_15196);
nor U16136 (N_16136,N_15660,N_15530);
xor U16137 (N_16137,N_15571,N_15610);
nand U16138 (N_16138,N_15562,N_15859);
and U16139 (N_16139,N_15479,N_15784);
or U16140 (N_16140,N_15231,N_15960);
xnor U16141 (N_16141,N_15598,N_15745);
nor U16142 (N_16142,N_15264,N_15201);
nor U16143 (N_16143,N_15368,N_15031);
nand U16144 (N_16144,N_15513,N_15346);
and U16145 (N_16145,N_15999,N_15803);
and U16146 (N_16146,N_15450,N_15878);
nor U16147 (N_16147,N_15462,N_15839);
or U16148 (N_16148,N_15650,N_15810);
xnor U16149 (N_16149,N_15599,N_15695);
xor U16150 (N_16150,N_15808,N_15021);
or U16151 (N_16151,N_15925,N_15856);
or U16152 (N_16152,N_15124,N_15697);
or U16153 (N_16153,N_15752,N_15625);
and U16154 (N_16154,N_15234,N_15322);
or U16155 (N_16155,N_15243,N_15727);
or U16156 (N_16156,N_15456,N_15344);
and U16157 (N_16157,N_15954,N_15464);
xnor U16158 (N_16158,N_15155,N_15145);
or U16159 (N_16159,N_15996,N_15048);
or U16160 (N_16160,N_15066,N_15543);
xnor U16161 (N_16161,N_15849,N_15483);
xor U16162 (N_16162,N_15217,N_15140);
nand U16163 (N_16163,N_15701,N_15720);
xor U16164 (N_16164,N_15486,N_15493);
xnor U16165 (N_16165,N_15109,N_15050);
nand U16166 (N_16166,N_15018,N_15595);
xnor U16167 (N_16167,N_15764,N_15622);
or U16168 (N_16168,N_15646,N_15933);
nor U16169 (N_16169,N_15382,N_15741);
or U16170 (N_16170,N_15514,N_15820);
nor U16171 (N_16171,N_15558,N_15259);
and U16172 (N_16172,N_15111,N_15845);
or U16173 (N_16173,N_15747,N_15768);
xor U16174 (N_16174,N_15141,N_15936);
nand U16175 (N_16175,N_15601,N_15401);
and U16176 (N_16176,N_15986,N_15691);
and U16177 (N_16177,N_15678,N_15895);
nor U16178 (N_16178,N_15175,N_15824);
or U16179 (N_16179,N_15331,N_15249);
or U16180 (N_16180,N_15838,N_15221);
xnor U16181 (N_16181,N_15229,N_15723);
and U16182 (N_16182,N_15556,N_15235);
xnor U16183 (N_16183,N_15084,N_15415);
nand U16184 (N_16184,N_15433,N_15428);
and U16185 (N_16185,N_15064,N_15367);
xnor U16186 (N_16186,N_15760,N_15863);
nand U16187 (N_16187,N_15611,N_15636);
xnor U16188 (N_16188,N_15478,N_15308);
nand U16189 (N_16189,N_15164,N_15725);
nand U16190 (N_16190,N_15112,N_15613);
or U16191 (N_16191,N_15226,N_15362);
nor U16192 (N_16192,N_15531,N_15757);
and U16193 (N_16193,N_15276,N_15682);
or U16194 (N_16194,N_15606,N_15623);
or U16195 (N_16195,N_15831,N_15334);
xor U16196 (N_16196,N_15137,N_15758);
or U16197 (N_16197,N_15058,N_15928);
nor U16198 (N_16198,N_15967,N_15041);
and U16199 (N_16199,N_15147,N_15176);
nor U16200 (N_16200,N_15174,N_15342);
nand U16201 (N_16201,N_15247,N_15547);
and U16202 (N_16202,N_15358,N_15047);
nand U16203 (N_16203,N_15995,N_15879);
nand U16204 (N_16204,N_15662,N_15253);
or U16205 (N_16205,N_15343,N_15326);
and U16206 (N_16206,N_15872,N_15854);
or U16207 (N_16207,N_15736,N_15912);
or U16208 (N_16208,N_15717,N_15350);
xor U16209 (N_16209,N_15686,N_15654);
nand U16210 (N_16210,N_15886,N_15608);
xor U16211 (N_16211,N_15997,N_15732);
nand U16212 (N_16212,N_15157,N_15000);
nand U16213 (N_16213,N_15212,N_15639);
and U16214 (N_16214,N_15567,N_15749);
or U16215 (N_16215,N_15374,N_15705);
nand U16216 (N_16216,N_15038,N_15040);
xnor U16217 (N_16217,N_15640,N_15541);
and U16218 (N_16218,N_15357,N_15316);
nor U16219 (N_16219,N_15830,N_15735);
or U16220 (N_16220,N_15476,N_15165);
xnor U16221 (N_16221,N_15529,N_15299);
or U16222 (N_16222,N_15629,N_15238);
and U16223 (N_16223,N_15054,N_15674);
or U16224 (N_16224,N_15262,N_15866);
xnor U16225 (N_16225,N_15290,N_15576);
or U16226 (N_16226,N_15713,N_15395);
xnor U16227 (N_16227,N_15306,N_15588);
xor U16228 (N_16228,N_15285,N_15075);
and U16229 (N_16229,N_15289,N_15976);
nand U16230 (N_16230,N_15774,N_15022);
nor U16231 (N_16231,N_15942,N_15841);
nand U16232 (N_16232,N_15273,N_15523);
and U16233 (N_16233,N_15554,N_15746);
nor U16234 (N_16234,N_15818,N_15769);
nor U16235 (N_16235,N_15118,N_15935);
or U16236 (N_16236,N_15015,N_15826);
or U16237 (N_16237,N_15366,N_15794);
nor U16238 (N_16238,N_15699,N_15076);
or U16239 (N_16239,N_15947,N_15927);
nor U16240 (N_16240,N_15728,N_15108);
nand U16241 (N_16241,N_15409,N_15962);
and U16242 (N_16242,N_15268,N_15871);
and U16243 (N_16243,N_15981,N_15122);
xnor U16244 (N_16244,N_15407,N_15189);
xnor U16245 (N_16245,N_15921,N_15125);
or U16246 (N_16246,N_15210,N_15490);
nand U16247 (N_16247,N_15241,N_15239);
nor U16248 (N_16248,N_15481,N_15025);
nor U16249 (N_16249,N_15172,N_15497);
xor U16250 (N_16250,N_15897,N_15443);
and U16251 (N_16251,N_15718,N_15900);
or U16252 (N_16252,N_15055,N_15534);
and U16253 (N_16253,N_15518,N_15819);
nor U16254 (N_16254,N_15609,N_15812);
and U16255 (N_16255,N_15881,N_15591);
and U16256 (N_16256,N_15296,N_15767);
or U16257 (N_16257,N_15240,N_15004);
and U16258 (N_16258,N_15385,N_15620);
and U16259 (N_16259,N_15923,N_15913);
and U16260 (N_16260,N_15703,N_15167);
or U16261 (N_16261,N_15391,N_15068);
and U16262 (N_16262,N_15920,N_15039);
nand U16263 (N_16263,N_15648,N_15177);
or U16264 (N_16264,N_15158,N_15230);
or U16265 (N_16265,N_15527,N_15582);
nor U16266 (N_16266,N_15840,N_15684);
nor U16267 (N_16267,N_15150,N_15463);
or U16268 (N_16268,N_15113,N_15187);
nor U16269 (N_16269,N_15384,N_15056);
or U16270 (N_16270,N_15007,N_15744);
xor U16271 (N_16271,N_15447,N_15924);
or U16272 (N_16272,N_15894,N_15387);
nand U16273 (N_16273,N_15596,N_15771);
or U16274 (N_16274,N_15630,N_15858);
or U16275 (N_16275,N_15129,N_15852);
xor U16276 (N_16276,N_15807,N_15698);
or U16277 (N_16277,N_15722,N_15203);
and U16278 (N_16278,N_15635,N_15013);
and U16279 (N_16279,N_15453,N_15835);
nand U16280 (N_16280,N_15670,N_15577);
xnor U16281 (N_16281,N_15438,N_15181);
and U16282 (N_16282,N_15065,N_15339);
and U16283 (N_16283,N_15991,N_15904);
and U16284 (N_16284,N_15687,N_15501);
xnor U16285 (N_16285,N_15419,N_15202);
or U16286 (N_16286,N_15184,N_15772);
xnor U16287 (N_16287,N_15786,N_15627);
xor U16288 (N_16288,N_15120,N_15560);
and U16289 (N_16289,N_15506,N_15348);
or U16290 (N_16290,N_15889,N_15307);
xor U16291 (N_16291,N_15097,N_15661);
xnor U16292 (N_16292,N_15874,N_15063);
xnor U16293 (N_16293,N_15710,N_15602);
nor U16294 (N_16294,N_15918,N_15252);
nor U16295 (N_16295,N_15916,N_15349);
nand U16296 (N_16296,N_15028,N_15914);
or U16297 (N_16297,N_15163,N_15857);
xnor U16298 (N_16298,N_15127,N_15982);
nor U16299 (N_16299,N_15074,N_15128);
xor U16300 (N_16300,N_15788,N_15371);
xnor U16301 (N_16301,N_15816,N_15260);
and U16302 (N_16302,N_15219,N_15796);
and U16303 (N_16303,N_15146,N_15873);
or U16304 (N_16304,N_15876,N_15983);
nor U16305 (N_16305,N_15223,N_15271);
or U16306 (N_16306,N_15908,N_15254);
nor U16307 (N_16307,N_15499,N_15328);
or U16308 (N_16308,N_15005,N_15430);
nor U16309 (N_16309,N_15994,N_15138);
nor U16310 (N_16310,N_15059,N_15380);
xor U16311 (N_16311,N_15555,N_15930);
xnor U16312 (N_16312,N_15738,N_15696);
or U16313 (N_16313,N_15643,N_15293);
and U16314 (N_16314,N_15458,N_15776);
nor U16315 (N_16315,N_15716,N_15107);
xnor U16316 (N_16316,N_15460,N_15867);
and U16317 (N_16317,N_15011,N_15191);
or U16318 (N_16318,N_15364,N_15708);
xor U16319 (N_16319,N_15939,N_15532);
nand U16320 (N_16320,N_15232,N_15975);
or U16321 (N_16321,N_15502,N_15491);
xnor U16322 (N_16322,N_15341,N_15429);
nor U16323 (N_16323,N_15892,N_15469);
and U16324 (N_16324,N_15952,N_15480);
xnor U16325 (N_16325,N_15990,N_15423);
nand U16326 (N_16326,N_15303,N_15103);
and U16327 (N_16327,N_15711,N_15139);
or U16328 (N_16328,N_15644,N_15081);
nand U16329 (N_16329,N_15446,N_15282);
or U16330 (N_16330,N_15310,N_15426);
and U16331 (N_16331,N_15405,N_15457);
xor U16332 (N_16332,N_15652,N_15700);
xnor U16333 (N_16333,N_15770,N_15580);
xor U16334 (N_16334,N_15756,N_15077);
nor U16335 (N_16335,N_15192,N_15314);
nor U16336 (N_16336,N_15616,N_15525);
nor U16337 (N_16337,N_15811,N_15445);
xor U16338 (N_16338,N_15961,N_15020);
and U16339 (N_16339,N_15805,N_15006);
or U16340 (N_16340,N_15963,N_15473);
nor U16341 (N_16341,N_15719,N_15665);
nor U16342 (N_16342,N_15578,N_15325);
and U16343 (N_16343,N_15862,N_15638);
and U16344 (N_16344,N_15452,N_15557);
and U16345 (N_16345,N_15724,N_15496);
nor U16346 (N_16346,N_15731,N_15500);
or U16347 (N_16347,N_15837,N_15581);
and U16348 (N_16348,N_15402,N_15266);
and U16349 (N_16349,N_15220,N_15251);
nor U16350 (N_16350,N_15152,N_15115);
or U16351 (N_16351,N_15829,N_15550);
xnor U16352 (N_16352,N_15642,N_15663);
xnor U16353 (N_16353,N_15919,N_15045);
or U16354 (N_16354,N_15574,N_15060);
and U16355 (N_16355,N_15675,N_15256);
nor U16356 (N_16356,N_15381,N_15209);
nand U16357 (N_16357,N_15195,N_15789);
or U16358 (N_16358,N_15971,N_15225);
or U16359 (N_16359,N_15052,N_15079);
nor U16360 (N_16360,N_15087,N_15910);
nor U16361 (N_16361,N_15689,N_15422);
xnor U16362 (N_16362,N_15337,N_15114);
nand U16363 (N_16363,N_15206,N_15082);
xor U16364 (N_16364,N_15459,N_15324);
or U16365 (N_16365,N_15715,N_15275);
and U16366 (N_16366,N_15714,N_15057);
or U16367 (N_16367,N_15302,N_15410);
or U16368 (N_16368,N_15667,N_15657);
nand U16369 (N_16369,N_15046,N_15278);
nor U16370 (N_16370,N_15392,N_15753);
or U16371 (N_16371,N_15291,N_15136);
nor U16372 (N_16372,N_15002,N_15777);
or U16373 (N_16373,N_15605,N_15135);
or U16374 (N_16374,N_15806,N_15931);
xor U16375 (N_16375,N_15009,N_15782);
or U16376 (N_16376,N_15035,N_15377);
nand U16377 (N_16377,N_15509,N_15775);
and U16378 (N_16378,N_15117,N_15394);
nand U16379 (N_16379,N_15042,N_15679);
nor U16380 (N_16380,N_15412,N_15044);
xor U16381 (N_16381,N_15510,N_15403);
and U16382 (N_16382,N_15263,N_15442);
nor U16383 (N_16383,N_15905,N_15198);
and U16384 (N_16384,N_15049,N_15178);
or U16385 (N_16385,N_15317,N_15441);
or U16386 (N_16386,N_15964,N_15754);
nor U16387 (N_16387,N_15526,N_15932);
nand U16388 (N_16388,N_15864,N_15690);
or U16389 (N_16389,N_15528,N_15795);
nor U16390 (N_16390,N_15950,N_15095);
or U16391 (N_16391,N_15726,N_15614);
nand U16392 (N_16392,N_15495,N_15641);
nand U16393 (N_16393,N_15233,N_15134);
nand U16394 (N_16394,N_15205,N_15338);
nand U16395 (N_16395,N_15998,N_15304);
nand U16396 (N_16396,N_15204,N_15424);
or U16397 (N_16397,N_15319,N_15503);
nand U16398 (N_16398,N_15956,N_15267);
or U16399 (N_16399,N_15171,N_15185);
nor U16400 (N_16400,N_15801,N_15618);
nand U16401 (N_16401,N_15186,N_15987);
and U16402 (N_16402,N_15765,N_15417);
nor U16403 (N_16403,N_15149,N_15012);
nand U16404 (N_16404,N_15545,N_15369);
nand U16405 (N_16405,N_15330,N_15973);
xor U16406 (N_16406,N_15520,N_15257);
nand U16407 (N_16407,N_15957,N_15258);
xnor U16408 (N_16408,N_15893,N_15408);
xor U16409 (N_16409,N_15116,N_15199);
and U16410 (N_16410,N_15583,N_15564);
xor U16411 (N_16411,N_15355,N_15721);
or U16412 (N_16412,N_15817,N_15799);
nand U16413 (N_16413,N_15813,N_15619);
or U16414 (N_16414,N_15383,N_15748);
nor U16415 (N_16415,N_15993,N_15101);
xor U16416 (N_16416,N_15649,N_15664);
nand U16417 (N_16417,N_15489,N_15414);
xor U16418 (N_16418,N_15759,N_15156);
xor U16419 (N_16419,N_15435,N_15589);
nand U16420 (N_16420,N_15612,N_15085);
xnor U16421 (N_16421,N_15345,N_15311);
nand U16422 (N_16422,N_15397,N_15946);
nand U16423 (N_16423,N_15842,N_15389);
nor U16424 (N_16424,N_15737,N_15213);
nor U16425 (N_16425,N_15593,N_15968);
nand U16426 (N_16426,N_15988,N_15515);
xor U16427 (N_16427,N_15420,N_15507);
or U16428 (N_16428,N_15301,N_15131);
and U16429 (N_16429,N_15245,N_15475);
xor U16430 (N_16430,N_15901,N_15416);
xnor U16431 (N_16431,N_15425,N_15133);
or U16432 (N_16432,N_15773,N_15051);
nand U16433 (N_16433,N_15575,N_15110);
or U16434 (N_16434,N_15091,N_15440);
xor U16435 (N_16435,N_15166,N_15359);
and U16436 (N_16436,N_15312,N_15017);
xor U16437 (N_16437,N_15730,N_15617);
or U16438 (N_16438,N_15672,N_15539);
xnor U16439 (N_16439,N_15938,N_15751);
nor U16440 (N_16440,N_15929,N_15008);
and U16441 (N_16441,N_15677,N_15712);
and U16442 (N_16442,N_15255,N_15427);
or U16443 (N_16443,N_15868,N_15783);
nor U16444 (N_16444,N_15822,N_15398);
nor U16445 (N_16445,N_15985,N_15787);
or U16446 (N_16446,N_15200,N_15669);
nor U16447 (N_16447,N_15902,N_15676);
xnor U16448 (N_16448,N_15880,N_15944);
xor U16449 (N_16449,N_15779,N_15351);
nand U16450 (N_16450,N_15516,N_15569);
or U16451 (N_16451,N_15955,N_15067);
and U16452 (N_16452,N_15884,N_15980);
and U16453 (N_16453,N_15354,N_15535);
or U16454 (N_16454,N_15287,N_15600);
and U16455 (N_16455,N_15228,N_15626);
and U16456 (N_16456,N_15432,N_15553);
xor U16457 (N_16457,N_15628,N_15537);
nand U16458 (N_16458,N_15951,N_15305);
nand U16459 (N_16459,N_15953,N_15647);
or U16460 (N_16460,N_15170,N_15094);
nand U16461 (N_16461,N_15014,N_15521);
xor U16462 (N_16462,N_15182,N_15277);
nand U16463 (N_16463,N_15906,N_15088);
and U16464 (N_16464,N_15882,N_15597);
nand U16465 (N_16465,N_15032,N_15733);
nand U16466 (N_16466,N_15333,N_15360);
nor U16467 (N_16467,N_15281,N_15099);
nor U16468 (N_16468,N_15742,N_15542);
nand U16469 (N_16469,N_15673,N_15804);
nor U16470 (N_16470,N_15802,N_15361);
or U16471 (N_16471,N_15888,N_15444);
xnor U16472 (N_16472,N_15522,N_15037);
xor U16473 (N_16473,N_15466,N_15143);
and U16474 (N_16474,N_15828,N_15552);
nand U16475 (N_16475,N_15148,N_15036);
and U16476 (N_16476,N_15119,N_15400);
or U16477 (N_16477,N_15945,N_15566);
nor U16478 (N_16478,N_15763,N_15300);
and U16479 (N_16479,N_15434,N_15100);
xnor U16480 (N_16480,N_15653,N_15222);
nand U16481 (N_16481,N_15370,N_15034);
and U16482 (N_16482,N_15180,N_15188);
or U16483 (N_16483,N_15019,N_15214);
nand U16484 (N_16484,N_15594,N_15681);
nand U16485 (N_16485,N_15070,N_15086);
nand U16486 (N_16486,N_15877,N_15286);
xnor U16487 (N_16487,N_15825,N_15043);
xnor U16488 (N_16488,N_15151,N_15615);
nand U16489 (N_16489,N_15208,N_15823);
xnor U16490 (N_16490,N_15517,N_15468);
or U16491 (N_16491,N_15671,N_15668);
xnor U16492 (N_16492,N_15024,N_15958);
nand U16493 (N_16493,N_15248,N_15540);
and U16494 (N_16494,N_15340,N_15785);
or U16495 (N_16495,N_15694,N_15778);
xor U16496 (N_16496,N_15283,N_15568);
xor U16497 (N_16497,N_15224,N_15396);
or U16498 (N_16498,N_15666,N_15315);
nand U16499 (N_16499,N_15926,N_15970);
xnor U16500 (N_16500,N_15289,N_15636);
nor U16501 (N_16501,N_15256,N_15994);
or U16502 (N_16502,N_15115,N_15819);
xnor U16503 (N_16503,N_15580,N_15758);
and U16504 (N_16504,N_15616,N_15230);
nand U16505 (N_16505,N_15689,N_15611);
and U16506 (N_16506,N_15739,N_15119);
nor U16507 (N_16507,N_15719,N_15165);
or U16508 (N_16508,N_15104,N_15572);
and U16509 (N_16509,N_15737,N_15366);
xor U16510 (N_16510,N_15473,N_15911);
or U16511 (N_16511,N_15292,N_15877);
nor U16512 (N_16512,N_15720,N_15145);
nand U16513 (N_16513,N_15304,N_15254);
nand U16514 (N_16514,N_15097,N_15418);
or U16515 (N_16515,N_15595,N_15069);
nor U16516 (N_16516,N_15405,N_15795);
nand U16517 (N_16517,N_15121,N_15775);
and U16518 (N_16518,N_15221,N_15495);
xor U16519 (N_16519,N_15362,N_15737);
xor U16520 (N_16520,N_15154,N_15864);
xor U16521 (N_16521,N_15643,N_15867);
nand U16522 (N_16522,N_15491,N_15339);
nor U16523 (N_16523,N_15224,N_15014);
or U16524 (N_16524,N_15741,N_15679);
and U16525 (N_16525,N_15226,N_15939);
nand U16526 (N_16526,N_15352,N_15123);
xor U16527 (N_16527,N_15374,N_15894);
nand U16528 (N_16528,N_15567,N_15193);
xor U16529 (N_16529,N_15337,N_15119);
nor U16530 (N_16530,N_15623,N_15716);
or U16531 (N_16531,N_15088,N_15078);
nand U16532 (N_16532,N_15091,N_15823);
nor U16533 (N_16533,N_15738,N_15190);
and U16534 (N_16534,N_15984,N_15798);
or U16535 (N_16535,N_15204,N_15802);
nor U16536 (N_16536,N_15889,N_15765);
nand U16537 (N_16537,N_15878,N_15371);
xor U16538 (N_16538,N_15709,N_15409);
or U16539 (N_16539,N_15368,N_15213);
nand U16540 (N_16540,N_15262,N_15466);
xnor U16541 (N_16541,N_15533,N_15025);
nand U16542 (N_16542,N_15281,N_15793);
xnor U16543 (N_16543,N_15399,N_15124);
xnor U16544 (N_16544,N_15913,N_15717);
nor U16545 (N_16545,N_15303,N_15199);
and U16546 (N_16546,N_15097,N_15076);
xor U16547 (N_16547,N_15140,N_15224);
xor U16548 (N_16548,N_15664,N_15129);
xnor U16549 (N_16549,N_15528,N_15289);
xor U16550 (N_16550,N_15137,N_15423);
and U16551 (N_16551,N_15629,N_15368);
and U16552 (N_16552,N_15406,N_15918);
and U16553 (N_16553,N_15828,N_15256);
and U16554 (N_16554,N_15058,N_15106);
or U16555 (N_16555,N_15641,N_15132);
xor U16556 (N_16556,N_15576,N_15337);
xnor U16557 (N_16557,N_15302,N_15900);
xor U16558 (N_16558,N_15309,N_15315);
and U16559 (N_16559,N_15743,N_15648);
and U16560 (N_16560,N_15188,N_15080);
nor U16561 (N_16561,N_15254,N_15335);
xnor U16562 (N_16562,N_15039,N_15007);
xor U16563 (N_16563,N_15608,N_15195);
nand U16564 (N_16564,N_15924,N_15282);
and U16565 (N_16565,N_15745,N_15092);
nand U16566 (N_16566,N_15442,N_15210);
and U16567 (N_16567,N_15208,N_15476);
nor U16568 (N_16568,N_15602,N_15554);
nand U16569 (N_16569,N_15578,N_15134);
xnor U16570 (N_16570,N_15005,N_15626);
nor U16571 (N_16571,N_15343,N_15652);
and U16572 (N_16572,N_15298,N_15555);
or U16573 (N_16573,N_15831,N_15657);
and U16574 (N_16574,N_15100,N_15071);
xor U16575 (N_16575,N_15845,N_15694);
or U16576 (N_16576,N_15662,N_15302);
nor U16577 (N_16577,N_15670,N_15932);
and U16578 (N_16578,N_15982,N_15081);
nand U16579 (N_16579,N_15192,N_15823);
nand U16580 (N_16580,N_15503,N_15255);
xnor U16581 (N_16581,N_15495,N_15413);
nand U16582 (N_16582,N_15752,N_15426);
xor U16583 (N_16583,N_15838,N_15554);
nor U16584 (N_16584,N_15572,N_15573);
and U16585 (N_16585,N_15037,N_15683);
xor U16586 (N_16586,N_15507,N_15446);
xnor U16587 (N_16587,N_15059,N_15817);
xnor U16588 (N_16588,N_15124,N_15283);
and U16589 (N_16589,N_15266,N_15112);
nand U16590 (N_16590,N_15420,N_15352);
or U16591 (N_16591,N_15113,N_15938);
xor U16592 (N_16592,N_15600,N_15299);
or U16593 (N_16593,N_15993,N_15111);
and U16594 (N_16594,N_15685,N_15945);
nor U16595 (N_16595,N_15492,N_15182);
and U16596 (N_16596,N_15689,N_15164);
nand U16597 (N_16597,N_15295,N_15891);
nand U16598 (N_16598,N_15660,N_15531);
nor U16599 (N_16599,N_15296,N_15338);
xnor U16600 (N_16600,N_15252,N_15059);
nor U16601 (N_16601,N_15967,N_15656);
nand U16602 (N_16602,N_15899,N_15763);
nor U16603 (N_16603,N_15512,N_15925);
nand U16604 (N_16604,N_15575,N_15358);
xor U16605 (N_16605,N_15472,N_15245);
and U16606 (N_16606,N_15868,N_15250);
nand U16607 (N_16607,N_15961,N_15728);
nand U16608 (N_16608,N_15539,N_15852);
and U16609 (N_16609,N_15486,N_15057);
and U16610 (N_16610,N_15578,N_15938);
and U16611 (N_16611,N_15545,N_15872);
and U16612 (N_16612,N_15822,N_15505);
xor U16613 (N_16613,N_15299,N_15152);
xor U16614 (N_16614,N_15302,N_15934);
or U16615 (N_16615,N_15545,N_15172);
and U16616 (N_16616,N_15258,N_15265);
nand U16617 (N_16617,N_15913,N_15303);
nor U16618 (N_16618,N_15526,N_15211);
nand U16619 (N_16619,N_15826,N_15356);
xnor U16620 (N_16620,N_15352,N_15029);
nand U16621 (N_16621,N_15037,N_15543);
xnor U16622 (N_16622,N_15123,N_15781);
or U16623 (N_16623,N_15147,N_15891);
or U16624 (N_16624,N_15219,N_15308);
nand U16625 (N_16625,N_15100,N_15153);
nor U16626 (N_16626,N_15763,N_15600);
nand U16627 (N_16627,N_15052,N_15589);
xor U16628 (N_16628,N_15060,N_15975);
or U16629 (N_16629,N_15015,N_15836);
nand U16630 (N_16630,N_15369,N_15497);
xnor U16631 (N_16631,N_15057,N_15501);
or U16632 (N_16632,N_15470,N_15504);
or U16633 (N_16633,N_15364,N_15694);
nor U16634 (N_16634,N_15389,N_15450);
or U16635 (N_16635,N_15884,N_15454);
xor U16636 (N_16636,N_15137,N_15060);
nor U16637 (N_16637,N_15728,N_15012);
or U16638 (N_16638,N_15084,N_15595);
and U16639 (N_16639,N_15695,N_15351);
nor U16640 (N_16640,N_15757,N_15798);
xor U16641 (N_16641,N_15067,N_15099);
and U16642 (N_16642,N_15357,N_15656);
and U16643 (N_16643,N_15004,N_15712);
and U16644 (N_16644,N_15210,N_15237);
xnor U16645 (N_16645,N_15004,N_15530);
and U16646 (N_16646,N_15591,N_15304);
and U16647 (N_16647,N_15341,N_15872);
nor U16648 (N_16648,N_15904,N_15054);
or U16649 (N_16649,N_15381,N_15506);
or U16650 (N_16650,N_15200,N_15402);
nand U16651 (N_16651,N_15859,N_15238);
or U16652 (N_16652,N_15548,N_15512);
nor U16653 (N_16653,N_15793,N_15290);
and U16654 (N_16654,N_15268,N_15334);
nand U16655 (N_16655,N_15028,N_15054);
and U16656 (N_16656,N_15444,N_15484);
or U16657 (N_16657,N_15823,N_15570);
xor U16658 (N_16658,N_15413,N_15461);
or U16659 (N_16659,N_15700,N_15745);
xnor U16660 (N_16660,N_15174,N_15284);
xnor U16661 (N_16661,N_15668,N_15502);
and U16662 (N_16662,N_15248,N_15228);
nor U16663 (N_16663,N_15836,N_15394);
nor U16664 (N_16664,N_15331,N_15469);
xnor U16665 (N_16665,N_15939,N_15264);
or U16666 (N_16666,N_15198,N_15598);
or U16667 (N_16667,N_15995,N_15785);
xnor U16668 (N_16668,N_15319,N_15594);
or U16669 (N_16669,N_15478,N_15873);
and U16670 (N_16670,N_15503,N_15655);
nor U16671 (N_16671,N_15454,N_15096);
and U16672 (N_16672,N_15832,N_15516);
and U16673 (N_16673,N_15660,N_15824);
or U16674 (N_16674,N_15255,N_15668);
nand U16675 (N_16675,N_15587,N_15632);
xor U16676 (N_16676,N_15426,N_15537);
or U16677 (N_16677,N_15230,N_15697);
or U16678 (N_16678,N_15853,N_15965);
xor U16679 (N_16679,N_15215,N_15466);
or U16680 (N_16680,N_15546,N_15992);
xor U16681 (N_16681,N_15358,N_15014);
nor U16682 (N_16682,N_15729,N_15206);
and U16683 (N_16683,N_15696,N_15586);
or U16684 (N_16684,N_15978,N_15586);
nand U16685 (N_16685,N_15175,N_15608);
xnor U16686 (N_16686,N_15222,N_15941);
and U16687 (N_16687,N_15257,N_15022);
nor U16688 (N_16688,N_15299,N_15619);
xor U16689 (N_16689,N_15033,N_15160);
nor U16690 (N_16690,N_15262,N_15875);
xnor U16691 (N_16691,N_15148,N_15205);
and U16692 (N_16692,N_15069,N_15682);
xnor U16693 (N_16693,N_15494,N_15331);
nor U16694 (N_16694,N_15258,N_15741);
nor U16695 (N_16695,N_15669,N_15169);
or U16696 (N_16696,N_15302,N_15260);
nor U16697 (N_16697,N_15281,N_15823);
or U16698 (N_16698,N_15806,N_15900);
or U16699 (N_16699,N_15550,N_15156);
xnor U16700 (N_16700,N_15685,N_15303);
nand U16701 (N_16701,N_15557,N_15514);
and U16702 (N_16702,N_15075,N_15977);
nor U16703 (N_16703,N_15939,N_15447);
or U16704 (N_16704,N_15994,N_15167);
or U16705 (N_16705,N_15908,N_15172);
xor U16706 (N_16706,N_15752,N_15605);
nor U16707 (N_16707,N_15173,N_15027);
nor U16708 (N_16708,N_15785,N_15065);
or U16709 (N_16709,N_15760,N_15268);
xor U16710 (N_16710,N_15990,N_15142);
nand U16711 (N_16711,N_15769,N_15980);
or U16712 (N_16712,N_15854,N_15946);
and U16713 (N_16713,N_15262,N_15126);
nand U16714 (N_16714,N_15943,N_15577);
xor U16715 (N_16715,N_15749,N_15714);
or U16716 (N_16716,N_15603,N_15121);
nand U16717 (N_16717,N_15067,N_15865);
nor U16718 (N_16718,N_15122,N_15998);
xor U16719 (N_16719,N_15848,N_15613);
or U16720 (N_16720,N_15356,N_15044);
nor U16721 (N_16721,N_15519,N_15076);
and U16722 (N_16722,N_15034,N_15301);
or U16723 (N_16723,N_15507,N_15916);
xor U16724 (N_16724,N_15122,N_15113);
xnor U16725 (N_16725,N_15658,N_15335);
or U16726 (N_16726,N_15810,N_15121);
nand U16727 (N_16727,N_15572,N_15232);
and U16728 (N_16728,N_15975,N_15377);
nand U16729 (N_16729,N_15999,N_15598);
or U16730 (N_16730,N_15000,N_15544);
nand U16731 (N_16731,N_15578,N_15135);
xnor U16732 (N_16732,N_15145,N_15689);
nor U16733 (N_16733,N_15617,N_15248);
nand U16734 (N_16734,N_15451,N_15329);
xnor U16735 (N_16735,N_15421,N_15574);
and U16736 (N_16736,N_15268,N_15165);
nand U16737 (N_16737,N_15546,N_15425);
nand U16738 (N_16738,N_15700,N_15124);
or U16739 (N_16739,N_15690,N_15596);
nand U16740 (N_16740,N_15212,N_15652);
xor U16741 (N_16741,N_15191,N_15422);
or U16742 (N_16742,N_15070,N_15001);
xor U16743 (N_16743,N_15043,N_15360);
and U16744 (N_16744,N_15826,N_15325);
and U16745 (N_16745,N_15999,N_15562);
xnor U16746 (N_16746,N_15145,N_15940);
nor U16747 (N_16747,N_15788,N_15434);
or U16748 (N_16748,N_15818,N_15923);
nand U16749 (N_16749,N_15525,N_15550);
or U16750 (N_16750,N_15577,N_15499);
and U16751 (N_16751,N_15400,N_15964);
xor U16752 (N_16752,N_15320,N_15355);
or U16753 (N_16753,N_15078,N_15387);
nor U16754 (N_16754,N_15385,N_15440);
and U16755 (N_16755,N_15697,N_15745);
and U16756 (N_16756,N_15605,N_15532);
xor U16757 (N_16757,N_15423,N_15533);
xor U16758 (N_16758,N_15734,N_15666);
xnor U16759 (N_16759,N_15498,N_15916);
nor U16760 (N_16760,N_15444,N_15241);
and U16761 (N_16761,N_15441,N_15268);
nor U16762 (N_16762,N_15989,N_15947);
nand U16763 (N_16763,N_15498,N_15331);
nand U16764 (N_16764,N_15764,N_15540);
xor U16765 (N_16765,N_15620,N_15009);
nor U16766 (N_16766,N_15301,N_15695);
xnor U16767 (N_16767,N_15732,N_15559);
or U16768 (N_16768,N_15592,N_15323);
and U16769 (N_16769,N_15960,N_15557);
nor U16770 (N_16770,N_15508,N_15614);
xnor U16771 (N_16771,N_15894,N_15819);
xnor U16772 (N_16772,N_15828,N_15182);
and U16773 (N_16773,N_15714,N_15593);
nor U16774 (N_16774,N_15556,N_15616);
or U16775 (N_16775,N_15704,N_15686);
xnor U16776 (N_16776,N_15489,N_15109);
nor U16777 (N_16777,N_15076,N_15274);
nand U16778 (N_16778,N_15134,N_15739);
xor U16779 (N_16779,N_15112,N_15101);
nand U16780 (N_16780,N_15228,N_15743);
nor U16781 (N_16781,N_15146,N_15867);
xnor U16782 (N_16782,N_15485,N_15859);
or U16783 (N_16783,N_15115,N_15918);
nor U16784 (N_16784,N_15484,N_15917);
nand U16785 (N_16785,N_15519,N_15520);
or U16786 (N_16786,N_15257,N_15353);
xnor U16787 (N_16787,N_15597,N_15083);
xor U16788 (N_16788,N_15555,N_15083);
nor U16789 (N_16789,N_15647,N_15628);
nor U16790 (N_16790,N_15230,N_15831);
nor U16791 (N_16791,N_15778,N_15356);
and U16792 (N_16792,N_15447,N_15581);
nand U16793 (N_16793,N_15323,N_15047);
and U16794 (N_16794,N_15675,N_15896);
xor U16795 (N_16795,N_15908,N_15209);
and U16796 (N_16796,N_15401,N_15330);
or U16797 (N_16797,N_15786,N_15018);
xor U16798 (N_16798,N_15829,N_15227);
nand U16799 (N_16799,N_15373,N_15957);
and U16800 (N_16800,N_15315,N_15823);
xnor U16801 (N_16801,N_15031,N_15678);
and U16802 (N_16802,N_15721,N_15915);
nor U16803 (N_16803,N_15442,N_15294);
nand U16804 (N_16804,N_15552,N_15669);
nor U16805 (N_16805,N_15956,N_15943);
nor U16806 (N_16806,N_15520,N_15754);
xnor U16807 (N_16807,N_15329,N_15952);
and U16808 (N_16808,N_15585,N_15842);
and U16809 (N_16809,N_15747,N_15788);
or U16810 (N_16810,N_15290,N_15582);
nand U16811 (N_16811,N_15245,N_15485);
xnor U16812 (N_16812,N_15284,N_15712);
or U16813 (N_16813,N_15907,N_15459);
nand U16814 (N_16814,N_15323,N_15720);
or U16815 (N_16815,N_15675,N_15510);
xor U16816 (N_16816,N_15227,N_15031);
xnor U16817 (N_16817,N_15008,N_15751);
nand U16818 (N_16818,N_15566,N_15840);
nand U16819 (N_16819,N_15159,N_15997);
xnor U16820 (N_16820,N_15923,N_15236);
xor U16821 (N_16821,N_15049,N_15976);
nor U16822 (N_16822,N_15508,N_15875);
and U16823 (N_16823,N_15992,N_15065);
xor U16824 (N_16824,N_15177,N_15160);
and U16825 (N_16825,N_15614,N_15917);
xnor U16826 (N_16826,N_15720,N_15127);
nand U16827 (N_16827,N_15979,N_15009);
xor U16828 (N_16828,N_15779,N_15111);
nand U16829 (N_16829,N_15374,N_15779);
and U16830 (N_16830,N_15211,N_15446);
and U16831 (N_16831,N_15532,N_15880);
nand U16832 (N_16832,N_15010,N_15165);
nor U16833 (N_16833,N_15476,N_15825);
xnor U16834 (N_16834,N_15409,N_15745);
and U16835 (N_16835,N_15665,N_15046);
nand U16836 (N_16836,N_15219,N_15612);
or U16837 (N_16837,N_15298,N_15830);
or U16838 (N_16838,N_15421,N_15018);
and U16839 (N_16839,N_15215,N_15277);
and U16840 (N_16840,N_15142,N_15469);
and U16841 (N_16841,N_15590,N_15835);
xnor U16842 (N_16842,N_15098,N_15141);
xor U16843 (N_16843,N_15476,N_15562);
nor U16844 (N_16844,N_15419,N_15784);
nand U16845 (N_16845,N_15673,N_15668);
nor U16846 (N_16846,N_15941,N_15691);
and U16847 (N_16847,N_15027,N_15905);
nor U16848 (N_16848,N_15008,N_15523);
nand U16849 (N_16849,N_15751,N_15604);
nor U16850 (N_16850,N_15157,N_15221);
and U16851 (N_16851,N_15189,N_15650);
nor U16852 (N_16852,N_15779,N_15743);
nand U16853 (N_16853,N_15171,N_15385);
nand U16854 (N_16854,N_15917,N_15171);
or U16855 (N_16855,N_15523,N_15268);
or U16856 (N_16856,N_15049,N_15833);
xnor U16857 (N_16857,N_15040,N_15562);
xor U16858 (N_16858,N_15991,N_15881);
or U16859 (N_16859,N_15036,N_15494);
and U16860 (N_16860,N_15386,N_15292);
or U16861 (N_16861,N_15838,N_15270);
xor U16862 (N_16862,N_15298,N_15645);
xnor U16863 (N_16863,N_15822,N_15277);
nor U16864 (N_16864,N_15472,N_15276);
xnor U16865 (N_16865,N_15633,N_15889);
nand U16866 (N_16866,N_15343,N_15575);
xor U16867 (N_16867,N_15860,N_15009);
and U16868 (N_16868,N_15519,N_15364);
xnor U16869 (N_16869,N_15984,N_15114);
or U16870 (N_16870,N_15320,N_15917);
nor U16871 (N_16871,N_15841,N_15432);
or U16872 (N_16872,N_15306,N_15877);
and U16873 (N_16873,N_15773,N_15311);
nand U16874 (N_16874,N_15958,N_15774);
nand U16875 (N_16875,N_15632,N_15477);
nor U16876 (N_16876,N_15809,N_15944);
nor U16877 (N_16877,N_15107,N_15502);
nor U16878 (N_16878,N_15269,N_15791);
and U16879 (N_16879,N_15965,N_15704);
or U16880 (N_16880,N_15274,N_15503);
nor U16881 (N_16881,N_15659,N_15864);
and U16882 (N_16882,N_15647,N_15303);
or U16883 (N_16883,N_15904,N_15640);
nor U16884 (N_16884,N_15505,N_15789);
nor U16885 (N_16885,N_15827,N_15460);
xor U16886 (N_16886,N_15946,N_15812);
xnor U16887 (N_16887,N_15095,N_15966);
nand U16888 (N_16888,N_15981,N_15898);
nand U16889 (N_16889,N_15088,N_15972);
nand U16890 (N_16890,N_15112,N_15778);
nor U16891 (N_16891,N_15737,N_15893);
nand U16892 (N_16892,N_15844,N_15921);
nand U16893 (N_16893,N_15382,N_15974);
nor U16894 (N_16894,N_15324,N_15466);
and U16895 (N_16895,N_15245,N_15952);
nor U16896 (N_16896,N_15775,N_15442);
nor U16897 (N_16897,N_15789,N_15724);
xor U16898 (N_16898,N_15413,N_15622);
nor U16899 (N_16899,N_15065,N_15918);
nor U16900 (N_16900,N_15275,N_15617);
or U16901 (N_16901,N_15713,N_15180);
and U16902 (N_16902,N_15221,N_15874);
and U16903 (N_16903,N_15821,N_15852);
xnor U16904 (N_16904,N_15785,N_15339);
xnor U16905 (N_16905,N_15538,N_15133);
nand U16906 (N_16906,N_15460,N_15767);
or U16907 (N_16907,N_15359,N_15817);
and U16908 (N_16908,N_15280,N_15066);
xor U16909 (N_16909,N_15273,N_15935);
nor U16910 (N_16910,N_15219,N_15753);
nand U16911 (N_16911,N_15746,N_15582);
and U16912 (N_16912,N_15531,N_15801);
xor U16913 (N_16913,N_15489,N_15987);
or U16914 (N_16914,N_15875,N_15323);
and U16915 (N_16915,N_15323,N_15320);
nor U16916 (N_16916,N_15972,N_15065);
nand U16917 (N_16917,N_15134,N_15840);
and U16918 (N_16918,N_15614,N_15967);
nand U16919 (N_16919,N_15540,N_15733);
and U16920 (N_16920,N_15071,N_15596);
and U16921 (N_16921,N_15184,N_15892);
or U16922 (N_16922,N_15024,N_15163);
or U16923 (N_16923,N_15346,N_15750);
or U16924 (N_16924,N_15972,N_15659);
or U16925 (N_16925,N_15097,N_15277);
nor U16926 (N_16926,N_15631,N_15353);
and U16927 (N_16927,N_15023,N_15469);
nand U16928 (N_16928,N_15905,N_15165);
or U16929 (N_16929,N_15427,N_15934);
nor U16930 (N_16930,N_15730,N_15573);
and U16931 (N_16931,N_15927,N_15315);
nor U16932 (N_16932,N_15314,N_15858);
nor U16933 (N_16933,N_15999,N_15547);
and U16934 (N_16934,N_15285,N_15218);
nor U16935 (N_16935,N_15803,N_15080);
nor U16936 (N_16936,N_15408,N_15768);
nor U16937 (N_16937,N_15693,N_15878);
nor U16938 (N_16938,N_15643,N_15287);
xnor U16939 (N_16939,N_15089,N_15113);
and U16940 (N_16940,N_15321,N_15624);
or U16941 (N_16941,N_15569,N_15123);
and U16942 (N_16942,N_15700,N_15976);
nor U16943 (N_16943,N_15196,N_15941);
xor U16944 (N_16944,N_15931,N_15507);
xnor U16945 (N_16945,N_15282,N_15765);
and U16946 (N_16946,N_15664,N_15209);
xor U16947 (N_16947,N_15016,N_15318);
and U16948 (N_16948,N_15012,N_15086);
xor U16949 (N_16949,N_15969,N_15693);
or U16950 (N_16950,N_15304,N_15735);
or U16951 (N_16951,N_15202,N_15279);
nand U16952 (N_16952,N_15332,N_15995);
xor U16953 (N_16953,N_15318,N_15989);
and U16954 (N_16954,N_15747,N_15056);
nor U16955 (N_16955,N_15595,N_15144);
xnor U16956 (N_16956,N_15774,N_15303);
xor U16957 (N_16957,N_15607,N_15375);
nor U16958 (N_16958,N_15674,N_15042);
nor U16959 (N_16959,N_15699,N_15526);
nor U16960 (N_16960,N_15438,N_15909);
and U16961 (N_16961,N_15276,N_15783);
or U16962 (N_16962,N_15228,N_15318);
or U16963 (N_16963,N_15904,N_15050);
or U16964 (N_16964,N_15432,N_15726);
xnor U16965 (N_16965,N_15956,N_15902);
nand U16966 (N_16966,N_15790,N_15920);
nand U16967 (N_16967,N_15194,N_15665);
or U16968 (N_16968,N_15079,N_15936);
nand U16969 (N_16969,N_15883,N_15506);
xnor U16970 (N_16970,N_15274,N_15580);
nand U16971 (N_16971,N_15056,N_15624);
nand U16972 (N_16972,N_15682,N_15135);
xor U16973 (N_16973,N_15862,N_15219);
and U16974 (N_16974,N_15405,N_15428);
or U16975 (N_16975,N_15802,N_15635);
and U16976 (N_16976,N_15265,N_15168);
nor U16977 (N_16977,N_15610,N_15783);
and U16978 (N_16978,N_15303,N_15690);
or U16979 (N_16979,N_15205,N_15395);
xor U16980 (N_16980,N_15161,N_15413);
nor U16981 (N_16981,N_15555,N_15549);
nand U16982 (N_16982,N_15963,N_15598);
and U16983 (N_16983,N_15383,N_15935);
nor U16984 (N_16984,N_15919,N_15114);
nor U16985 (N_16985,N_15576,N_15486);
or U16986 (N_16986,N_15998,N_15372);
nand U16987 (N_16987,N_15258,N_15445);
nand U16988 (N_16988,N_15796,N_15706);
nor U16989 (N_16989,N_15094,N_15912);
and U16990 (N_16990,N_15989,N_15058);
and U16991 (N_16991,N_15067,N_15780);
nor U16992 (N_16992,N_15799,N_15053);
and U16993 (N_16993,N_15781,N_15725);
nor U16994 (N_16994,N_15258,N_15876);
or U16995 (N_16995,N_15550,N_15914);
nor U16996 (N_16996,N_15086,N_15722);
and U16997 (N_16997,N_15466,N_15970);
xnor U16998 (N_16998,N_15676,N_15316);
or U16999 (N_16999,N_15741,N_15172);
nand U17000 (N_17000,N_16951,N_16938);
nand U17001 (N_17001,N_16833,N_16140);
or U17002 (N_17002,N_16040,N_16479);
nor U17003 (N_17003,N_16043,N_16076);
nor U17004 (N_17004,N_16394,N_16760);
nand U17005 (N_17005,N_16415,N_16834);
nand U17006 (N_17006,N_16175,N_16227);
nor U17007 (N_17007,N_16462,N_16574);
xor U17008 (N_17008,N_16799,N_16783);
nor U17009 (N_17009,N_16813,N_16994);
and U17010 (N_17010,N_16587,N_16680);
nand U17011 (N_17011,N_16048,N_16715);
or U17012 (N_17012,N_16422,N_16859);
nand U17013 (N_17013,N_16558,N_16351);
nor U17014 (N_17014,N_16643,N_16662);
xnor U17015 (N_17015,N_16114,N_16473);
nand U17016 (N_17016,N_16821,N_16283);
nand U17017 (N_17017,N_16614,N_16285);
or U17018 (N_17018,N_16107,N_16890);
nor U17019 (N_17019,N_16915,N_16252);
or U17020 (N_17020,N_16204,N_16009);
and U17021 (N_17021,N_16554,N_16383);
and U17022 (N_17022,N_16709,N_16518);
and U17023 (N_17023,N_16499,N_16545);
nand U17024 (N_17024,N_16676,N_16253);
and U17025 (N_17025,N_16646,N_16376);
or U17026 (N_17026,N_16630,N_16322);
or U17027 (N_17027,N_16379,N_16069);
and U17028 (N_17028,N_16404,N_16240);
xnor U17029 (N_17029,N_16004,N_16976);
nor U17030 (N_17030,N_16918,N_16644);
xor U17031 (N_17031,N_16192,N_16441);
nor U17032 (N_17032,N_16496,N_16812);
or U17033 (N_17033,N_16233,N_16455);
or U17034 (N_17034,N_16300,N_16008);
or U17035 (N_17035,N_16958,N_16274);
or U17036 (N_17036,N_16012,N_16461);
nor U17037 (N_17037,N_16276,N_16758);
xor U17038 (N_17038,N_16442,N_16722);
and U17039 (N_17039,N_16143,N_16905);
xnor U17040 (N_17040,N_16210,N_16961);
nor U17041 (N_17041,N_16216,N_16016);
nor U17042 (N_17042,N_16932,N_16158);
nor U17043 (N_17043,N_16585,N_16549);
and U17044 (N_17044,N_16542,N_16962);
or U17045 (N_17045,N_16317,N_16567);
nor U17046 (N_17046,N_16242,N_16960);
xor U17047 (N_17047,N_16561,N_16718);
nor U17048 (N_17048,N_16658,N_16551);
and U17049 (N_17049,N_16267,N_16953);
xor U17050 (N_17050,N_16922,N_16031);
and U17051 (N_17051,N_16625,N_16544);
xor U17052 (N_17052,N_16772,N_16740);
and U17053 (N_17053,N_16973,N_16743);
and U17054 (N_17054,N_16309,N_16271);
xor U17055 (N_17055,N_16099,N_16801);
and U17056 (N_17056,N_16478,N_16495);
nand U17057 (N_17057,N_16494,N_16678);
xor U17058 (N_17058,N_16717,N_16051);
xnor U17059 (N_17059,N_16893,N_16897);
nor U17060 (N_17060,N_16703,N_16657);
and U17061 (N_17061,N_16557,N_16301);
and U17062 (N_17062,N_16452,N_16001);
nand U17063 (N_17063,N_16581,N_16806);
nand U17064 (N_17064,N_16590,N_16110);
nand U17065 (N_17065,N_16515,N_16367);
nand U17066 (N_17066,N_16524,N_16273);
xnor U17067 (N_17067,N_16900,N_16692);
xnor U17068 (N_17068,N_16446,N_16816);
and U17069 (N_17069,N_16521,N_16481);
nand U17070 (N_17070,N_16778,N_16347);
and U17071 (N_17071,N_16096,N_16117);
or U17072 (N_17072,N_16492,N_16670);
xnor U17073 (N_17073,N_16789,N_16203);
xor U17074 (N_17074,N_16675,N_16637);
nand U17075 (N_17075,N_16133,N_16293);
nand U17076 (N_17076,N_16519,N_16393);
xnor U17077 (N_17077,N_16366,N_16484);
nor U17078 (N_17078,N_16304,N_16170);
nand U17079 (N_17079,N_16250,N_16700);
nand U17080 (N_17080,N_16901,N_16705);
xor U17081 (N_17081,N_16123,N_16400);
xnor U17082 (N_17082,N_16919,N_16934);
nand U17083 (N_17083,N_16259,N_16555);
xnor U17084 (N_17084,N_16520,N_16889);
xnor U17085 (N_17085,N_16762,N_16371);
or U17086 (N_17086,N_16674,N_16916);
nand U17087 (N_17087,N_16505,N_16995);
nor U17088 (N_17088,N_16305,N_16981);
xor U17089 (N_17089,N_16723,N_16629);
and U17090 (N_17090,N_16620,N_16380);
and U17091 (N_17091,N_16530,N_16825);
nand U17092 (N_17092,N_16493,N_16539);
nand U17093 (N_17093,N_16337,N_16513);
nor U17094 (N_17094,N_16753,N_16419);
and U17095 (N_17095,N_16475,N_16179);
or U17096 (N_17096,N_16598,N_16594);
and U17097 (N_17097,N_16262,N_16209);
and U17098 (N_17098,N_16592,N_16792);
xor U17099 (N_17099,N_16306,N_16328);
nand U17100 (N_17100,N_16669,N_16164);
or U17101 (N_17101,N_16313,N_16220);
and U17102 (N_17102,N_16850,N_16200);
nor U17103 (N_17103,N_16318,N_16467);
nand U17104 (N_17104,N_16272,N_16876);
nand U17105 (N_17105,N_16432,N_16745);
and U17106 (N_17106,N_16390,N_16042);
nor U17107 (N_17107,N_16489,N_16485);
or U17108 (N_17108,N_16696,N_16898);
nor U17109 (N_17109,N_16018,N_16565);
or U17110 (N_17110,N_16427,N_16977);
nor U17111 (N_17111,N_16027,N_16580);
and U17112 (N_17112,N_16111,N_16136);
and U17113 (N_17113,N_16755,N_16023);
and U17114 (N_17114,N_16765,N_16997);
or U17115 (N_17115,N_16634,N_16720);
nor U17116 (N_17116,N_16661,N_16509);
nor U17117 (N_17117,N_16236,N_16451);
xnor U17118 (N_17118,N_16217,N_16221);
xnor U17119 (N_17119,N_16194,N_16529);
nor U17120 (N_17120,N_16168,N_16677);
nor U17121 (N_17121,N_16085,N_16497);
nor U17122 (N_17122,N_16845,N_16296);
nand U17123 (N_17123,N_16928,N_16548);
xnor U17124 (N_17124,N_16603,N_16989);
or U17125 (N_17125,N_16754,N_16647);
and U17126 (N_17126,N_16576,N_16345);
xnor U17127 (N_17127,N_16161,N_16418);
nand U17128 (N_17128,N_16104,N_16829);
nor U17129 (N_17129,N_16207,N_16819);
xnor U17130 (N_17130,N_16483,N_16095);
nor U17131 (N_17131,N_16358,N_16132);
nand U17132 (N_17132,N_16279,N_16109);
or U17133 (N_17133,N_16502,N_16206);
or U17134 (N_17134,N_16399,N_16959);
nand U17135 (N_17135,N_16269,N_16438);
and U17136 (N_17136,N_16795,N_16189);
xnor U17137 (N_17137,N_16965,N_16730);
nand U17138 (N_17138,N_16550,N_16857);
xor U17139 (N_17139,N_16425,N_16270);
nor U17140 (N_17140,N_16124,N_16612);
nand U17141 (N_17141,N_16011,N_16865);
and U17142 (N_17142,N_16844,N_16190);
or U17143 (N_17143,N_16057,N_16556);
and U17144 (N_17144,N_16824,N_16421);
or U17145 (N_17145,N_16453,N_16688);
or U17146 (N_17146,N_16909,N_16992);
or U17147 (N_17147,N_16343,N_16039);
and U17148 (N_17148,N_16943,N_16516);
or U17149 (N_17149,N_16106,N_16346);
nand U17150 (N_17150,N_16781,N_16780);
or U17151 (N_17151,N_16022,N_16239);
nand U17152 (N_17152,N_16407,N_16002);
or U17153 (N_17153,N_16146,N_16249);
and U17154 (N_17154,N_16144,N_16998);
xor U17155 (N_17155,N_16195,N_16906);
nor U17156 (N_17156,N_16609,N_16284);
and U17157 (N_17157,N_16639,N_16289);
and U17158 (N_17158,N_16796,N_16385);
nand U17159 (N_17159,N_16822,N_16986);
xnor U17160 (N_17160,N_16948,N_16842);
or U17161 (N_17161,N_16817,N_16097);
nand U17162 (N_17162,N_16130,N_16735);
xnor U17163 (N_17163,N_16560,N_16682);
xor U17164 (N_17164,N_16840,N_16779);
or U17165 (N_17165,N_16984,N_16597);
nand U17166 (N_17166,N_16666,N_16826);
nand U17167 (N_17167,N_16389,N_16626);
nor U17168 (N_17168,N_16913,N_16884);
xnor U17169 (N_17169,N_16155,N_16980);
or U17170 (N_17170,N_16299,N_16342);
or U17171 (N_17171,N_16782,N_16751);
and U17172 (N_17172,N_16532,N_16761);
nor U17173 (N_17173,N_16686,N_16064);
nor U17174 (N_17174,N_16511,N_16664);
and U17175 (N_17175,N_16727,N_16465);
nor U17176 (N_17176,N_16635,N_16794);
or U17177 (N_17177,N_16444,N_16098);
nand U17178 (N_17178,N_16904,N_16330);
or U17179 (N_17179,N_16184,N_16134);
xor U17180 (N_17180,N_16266,N_16858);
nor U17181 (N_17181,N_16923,N_16186);
or U17182 (N_17182,N_16288,N_16355);
xor U17183 (N_17183,N_16215,N_16294);
and U17184 (N_17184,N_16159,N_16254);
and U17185 (N_17185,N_16768,N_16747);
and U17186 (N_17186,N_16382,N_16596);
and U17187 (N_17187,N_16238,N_16401);
and U17188 (N_17188,N_16264,N_16854);
nand U17189 (N_17189,N_16275,N_16936);
nor U17190 (N_17190,N_16641,N_16245);
nor U17191 (N_17191,N_16457,N_16145);
and U17192 (N_17192,N_16650,N_16756);
and U17193 (N_17193,N_16610,N_16954);
xor U17194 (N_17194,N_16410,N_16374);
or U17195 (N_17195,N_16331,N_16402);
and U17196 (N_17196,N_16939,N_16258);
or U17197 (N_17197,N_16899,N_16608);
xor U17198 (N_17198,N_16291,N_16131);
nor U17199 (N_17199,N_16873,N_16029);
and U17200 (N_17200,N_16292,N_16055);
and U17201 (N_17201,N_16032,N_16437);
and U17202 (N_17202,N_16510,N_16126);
nor U17203 (N_17203,N_16800,N_16871);
or U17204 (N_17204,N_16020,N_16870);
nand U17205 (N_17205,N_16482,N_16037);
and U17206 (N_17206,N_16454,N_16571);
or U17207 (N_17207,N_16538,N_16531);
nand U17208 (N_17208,N_16263,N_16471);
xnor U17209 (N_17209,N_16070,N_16714);
xor U17210 (N_17210,N_16514,N_16562);
nor U17211 (N_17211,N_16791,N_16083);
or U17212 (N_17212,N_16757,N_16185);
xnor U17213 (N_17213,N_16147,N_16044);
xnor U17214 (N_17214,N_16137,N_16708);
xnor U17215 (N_17215,N_16302,N_16972);
nor U17216 (N_17216,N_16656,N_16623);
and U17217 (N_17217,N_16108,N_16935);
xnor U17218 (N_17218,N_16681,N_16573);
nor U17219 (N_17219,N_16828,N_16719);
xnor U17220 (N_17220,N_16447,N_16695);
or U17221 (N_17221,N_16710,N_16088);
nand U17222 (N_17222,N_16112,N_16320);
nor U17223 (N_17223,N_16063,N_16926);
nor U17224 (N_17224,N_16885,N_16163);
and U17225 (N_17225,N_16030,N_16196);
and U17226 (N_17226,N_16578,N_16640);
and U17227 (N_17227,N_16802,N_16982);
xor U17228 (N_17228,N_16075,N_16701);
nand U17229 (N_17229,N_16600,N_16153);
nand U17230 (N_17230,N_16653,N_16769);
nor U17231 (N_17231,N_16171,N_16183);
or U17232 (N_17232,N_16663,N_16373);
or U17233 (N_17233,N_16894,N_16752);
or U17234 (N_17234,N_16809,N_16181);
nand U17235 (N_17235,N_16101,N_16784);
xor U17236 (N_17236,N_16428,N_16135);
nand U17237 (N_17237,N_16082,N_16440);
or U17238 (N_17238,N_16248,N_16771);
or U17239 (N_17239,N_16308,N_16119);
and U17240 (N_17240,N_16583,N_16775);
or U17241 (N_17241,N_16472,N_16235);
xnor U17242 (N_17242,N_16952,N_16021);
nand U17243 (N_17243,N_16742,N_16823);
xor U17244 (N_17244,N_16464,N_16856);
nor U17245 (N_17245,N_16968,N_16247);
nor U17246 (N_17246,N_16738,N_16193);
xnor U17247 (N_17247,N_16282,N_16668);
and U17248 (N_17248,N_16324,N_16024);
or U17249 (N_17249,N_16586,N_16156);
nand U17250 (N_17250,N_16672,N_16173);
and U17251 (N_17251,N_16177,N_16855);
xnor U17252 (N_17252,N_16746,N_16166);
xnor U17253 (N_17253,N_16933,N_16729);
and U17254 (N_17254,N_16141,N_16007);
and U17255 (N_17255,N_16636,N_16671);
and U17256 (N_17256,N_16724,N_16359);
nor U17257 (N_17257,N_16244,N_16543);
nand U17258 (N_17258,N_16537,N_16246);
nor U17259 (N_17259,N_16602,N_16038);
or U17260 (N_17260,N_16748,N_16569);
and U17261 (N_17261,N_16526,N_16278);
nand U17262 (N_17262,N_16231,N_16632);
and U17263 (N_17263,N_16361,N_16956);
xor U17264 (N_17264,N_16501,N_16365);
nand U17265 (N_17265,N_16536,N_16619);
and U17266 (N_17266,N_16323,N_16793);
nor U17267 (N_17267,N_16103,N_16086);
xor U17268 (N_17268,N_16290,N_16102);
xnor U17269 (N_17269,N_16387,N_16559);
nand U17270 (N_17270,N_16469,N_16584);
nand U17271 (N_17271,N_16065,N_16955);
xnor U17272 (N_17272,N_16148,N_16862);
nand U17273 (N_17273,N_16903,N_16120);
or U17274 (N_17274,N_16533,N_16169);
nor U17275 (N_17275,N_16967,N_16439);
nand U17276 (N_17276,N_16176,N_16191);
nor U17277 (N_17277,N_16396,N_16835);
and U17278 (N_17278,N_16202,N_16251);
and U17279 (N_17279,N_16116,N_16491);
nand U17280 (N_17280,N_16080,N_16160);
and U17281 (N_17281,N_16412,N_16409);
or U17282 (N_17282,N_16414,N_16832);
and U17283 (N_17283,N_16566,N_16090);
xnor U17284 (N_17284,N_16458,N_16113);
nor U17285 (N_17285,N_16649,N_16622);
or U17286 (N_17286,N_16572,N_16797);
nand U17287 (N_17287,N_16974,N_16920);
nor U17288 (N_17288,N_16237,N_16424);
nor U17289 (N_17289,N_16297,N_16356);
xnor U17290 (N_17290,N_16613,N_16776);
xor U17291 (N_17291,N_16687,N_16887);
nor U17292 (N_17292,N_16333,N_16895);
xnor U17293 (N_17293,N_16525,N_16917);
xnor U17294 (N_17294,N_16459,N_16445);
and U17295 (N_17295,N_16852,N_16487);
nand U17296 (N_17296,N_16314,N_16049);
and U17297 (N_17297,N_16434,N_16931);
xnor U17298 (N_17298,N_16332,N_16881);
nor U17299 (N_17299,N_16225,N_16691);
and U17300 (N_17300,N_16831,N_16077);
and U17301 (N_17301,N_16413,N_16642);
nor U17302 (N_17302,N_16503,N_16712);
nand U17303 (N_17303,N_16803,N_16528);
xor U17304 (N_17304,N_16256,N_16138);
or U17305 (N_17305,N_16770,N_16734);
or U17306 (N_17306,N_16838,N_16019);
nand U17307 (N_17307,N_16033,N_16908);
nand U17308 (N_17308,N_16129,N_16564);
nand U17309 (N_17309,N_16633,N_16941);
nor U17310 (N_17310,N_16281,N_16942);
nor U17311 (N_17311,N_16218,N_16336);
nor U17312 (N_17312,N_16739,N_16589);
xnor U17313 (N_17313,N_16100,N_16224);
or U17314 (N_17314,N_16888,N_16398);
nor U17315 (N_17315,N_16352,N_16645);
xnor U17316 (N_17316,N_16326,N_16523);
nor U17317 (N_17317,N_16325,N_16966);
or U17318 (N_17318,N_16988,N_16693);
nor U17319 (N_17319,N_16456,N_16648);
and U17320 (N_17320,N_16257,N_16839);
nor U17321 (N_17321,N_16744,N_16041);
nor U17322 (N_17322,N_16068,N_16595);
and U17323 (N_17323,N_16848,N_16072);
nand U17324 (N_17324,N_16286,N_16035);
nand U17325 (N_17325,N_16201,N_16534);
nand U17326 (N_17326,N_16504,N_16577);
xor U17327 (N_17327,N_16711,N_16830);
or U17328 (N_17328,N_16690,N_16255);
and U17329 (N_17329,N_16728,N_16624);
nand U17330 (N_17330,N_16420,N_16386);
and U17331 (N_17331,N_16384,N_16867);
or U17332 (N_17332,N_16721,N_16945);
or U17333 (N_17333,N_16071,N_16853);
nor U17334 (N_17334,N_16378,N_16725);
xor U17335 (N_17335,N_16488,N_16214);
nor U17336 (N_17336,N_16621,N_16912);
nand U17337 (N_17337,N_16851,N_16774);
xor U17338 (N_17338,N_16868,N_16073);
xnor U17339 (N_17339,N_16448,N_16094);
xnor U17340 (N_17340,N_16869,N_16498);
or U17341 (N_17341,N_16655,N_16172);
nand U17342 (N_17342,N_16260,N_16363);
or U17343 (N_17343,N_16969,N_16814);
xor U17344 (N_17344,N_16733,N_16205);
or U17345 (N_17345,N_16990,N_16078);
nor U17346 (N_17346,N_16050,N_16927);
nand U17347 (N_17347,N_16341,N_16512);
nor U17348 (N_17348,N_16949,N_16836);
nand U17349 (N_17349,N_16843,N_16684);
xnor U17350 (N_17350,N_16327,N_16431);
nand U17351 (N_17351,N_16535,N_16615);
nor U17352 (N_17352,N_16391,N_16180);
nor U17353 (N_17353,N_16056,N_16470);
nor U17354 (N_17354,N_16174,N_16015);
nor U17355 (N_17355,N_16892,N_16921);
or U17356 (N_17356,N_16369,N_16010);
xnor U17357 (N_17357,N_16993,N_16226);
nor U17358 (N_17358,N_16058,N_16066);
and U17359 (N_17359,N_16879,N_16139);
xnor U17360 (N_17360,N_16785,N_16883);
nand U17361 (N_17361,N_16477,N_16570);
nor U17362 (N_17362,N_16875,N_16243);
nor U17363 (N_17363,N_16092,N_16679);
and U17364 (N_17364,N_16527,N_16790);
xor U17365 (N_17365,N_16430,N_16372);
xnor U17366 (N_17366,N_16187,N_16874);
nor U17367 (N_17367,N_16880,N_16810);
nor U17368 (N_17368,N_16408,N_16067);
xor U17369 (N_17369,N_16303,N_16907);
nor U17370 (N_17370,N_16999,N_16084);
or U17371 (N_17371,N_16277,N_16811);
nor U17372 (N_17372,N_16547,N_16368);
nand U17373 (N_17373,N_16486,N_16311);
or U17374 (N_17374,N_16540,N_16228);
and U17375 (N_17375,N_16213,N_16872);
or U17376 (N_17376,N_16338,N_16767);
nand U17377 (N_17377,N_16105,N_16506);
nand U17378 (N_17378,N_16081,N_16996);
or U17379 (N_17379,N_16659,N_16607);
nor U17380 (N_17380,N_16435,N_16468);
nor U17381 (N_17381,N_16449,N_16773);
nand U17382 (N_17382,N_16344,N_16759);
nor U17383 (N_17383,N_16517,N_16005);
xor U17384 (N_17384,N_16241,N_16052);
or U17385 (N_17385,N_16741,N_16925);
or U17386 (N_17386,N_16463,N_16706);
nand U17387 (N_17387,N_16827,N_16766);
or U17388 (N_17388,N_16298,N_16698);
nor U17389 (N_17389,N_16460,N_16093);
or U17390 (N_17390,N_16364,N_16047);
xnor U17391 (N_17391,N_16417,N_16651);
nor U17392 (N_17392,N_16152,N_16230);
or U17393 (N_17393,N_16697,N_16268);
nor U17394 (N_17394,N_16787,N_16307);
and U17395 (N_17395,N_16786,N_16059);
or U17396 (N_17396,N_16265,N_16234);
and U17397 (N_17397,N_16349,N_16036);
nand U17398 (N_17398,N_16028,N_16128);
xnor U17399 (N_17399,N_16060,N_16849);
xor U17400 (N_17400,N_16937,N_16074);
nand U17401 (N_17401,N_16388,N_16397);
nor U17402 (N_17402,N_16319,N_16947);
nor U17403 (N_17403,N_16929,N_16357);
or U17404 (N_17404,N_16553,N_16568);
nor U17405 (N_17405,N_16329,N_16142);
nor U17406 (N_17406,N_16611,N_16591);
and U17407 (N_17407,N_16654,N_16579);
nand U17408 (N_17408,N_16006,N_16987);
nand U17409 (N_17409,N_16749,N_16150);
nor U17410 (N_17410,N_16392,N_16353);
nor U17411 (N_17411,N_16370,N_16466);
and U17412 (N_17412,N_16866,N_16087);
and U17413 (N_17413,N_16025,N_16013);
xor U17414 (N_17414,N_16552,N_16606);
or U17415 (N_17415,N_16375,N_16593);
and U17416 (N_17416,N_16575,N_16985);
and U17417 (N_17417,N_16212,N_16122);
xnor U17418 (N_17418,N_16713,N_16726);
nand U17419 (N_17419,N_16798,N_16541);
and U17420 (N_17420,N_16704,N_16702);
or U17421 (N_17421,N_16991,N_16321);
or U17422 (N_17422,N_16436,N_16983);
xnor U17423 (N_17423,N_16588,N_16652);
or U17424 (N_17424,N_16683,N_16405);
nor U17425 (N_17425,N_16115,N_16522);
and U17426 (N_17426,N_16546,N_16053);
and U17427 (N_17427,N_16211,N_16699);
nand U17428 (N_17428,N_16685,N_16165);
nor U17429 (N_17429,N_16846,N_16911);
nand U17430 (N_17430,N_16601,N_16443);
or U17431 (N_17431,N_16638,N_16627);
nand U17432 (N_17432,N_16350,N_16154);
xnor U17433 (N_17433,N_16763,N_16805);
and U17434 (N_17434,N_16280,N_16978);
xnor U17435 (N_17435,N_16416,N_16157);
or U17436 (N_17436,N_16162,N_16360);
or U17437 (N_17437,N_16089,N_16979);
or U17438 (N_17438,N_16863,N_16310);
and U17439 (N_17439,N_16315,N_16062);
or U17440 (N_17440,N_16118,N_16667);
xnor U17441 (N_17441,N_16732,N_16970);
and U17442 (N_17442,N_16891,N_16957);
nor U17443 (N_17443,N_16930,N_16411);
nand U17444 (N_17444,N_16716,N_16563);
nand U17445 (N_17445,N_16000,N_16046);
or U17446 (N_17446,N_16689,N_16815);
nor U17447 (N_17447,N_16837,N_16731);
nand U17448 (N_17448,N_16229,N_16964);
or U17449 (N_17449,N_16232,N_16199);
nand U17450 (N_17450,N_16223,N_16339);
nor U17451 (N_17451,N_16673,N_16381);
nand U17452 (N_17452,N_16423,N_16335);
or U17453 (N_17453,N_16222,N_16508);
nand U17454 (N_17454,N_16354,N_16944);
nor U17455 (N_17455,N_16197,N_16014);
xnor U17456 (N_17456,N_16219,N_16582);
or U17457 (N_17457,N_16034,N_16334);
xor U17458 (N_17458,N_16707,N_16054);
or U17459 (N_17459,N_16861,N_16261);
nand U17460 (N_17460,N_16946,N_16188);
and U17461 (N_17461,N_16618,N_16198);
xor U17462 (N_17462,N_16631,N_16924);
xor U17463 (N_17463,N_16476,N_16149);
or U17464 (N_17464,N_16963,N_16295);
nor U17465 (N_17465,N_16807,N_16121);
nand U17466 (N_17466,N_16507,N_16788);
nand U17467 (N_17467,N_16061,N_16003);
xnor U17468 (N_17468,N_16841,N_16045);
nand U17469 (N_17469,N_16340,N_16617);
nand U17470 (N_17470,N_16808,N_16971);
or U17471 (N_17471,N_16450,N_16737);
xor U17472 (N_17472,N_16864,N_16480);
nand U17473 (N_17473,N_16820,N_16777);
and U17474 (N_17474,N_16599,N_16628);
xor U17475 (N_17475,N_16017,N_16605);
xor U17476 (N_17476,N_16125,N_16026);
xnor U17477 (N_17477,N_16604,N_16818);
xor U17478 (N_17478,N_16474,N_16665);
xnor U17479 (N_17479,N_16914,N_16886);
nand U17480 (N_17480,N_16616,N_16847);
or U17481 (N_17481,N_16287,N_16860);
xnor U17482 (N_17482,N_16377,N_16490);
nor U17483 (N_17483,N_16896,N_16312);
xor U17484 (N_17484,N_16975,N_16182);
nand U17485 (N_17485,N_16950,N_16736);
or U17486 (N_17486,N_16878,N_16750);
and U17487 (N_17487,N_16178,N_16433);
and U17488 (N_17488,N_16208,N_16902);
or U17489 (N_17489,N_16348,N_16316);
nand U17490 (N_17490,N_16764,N_16877);
or U17491 (N_17491,N_16500,N_16362);
nor U17492 (N_17492,N_16395,N_16940);
xnor U17493 (N_17493,N_16403,N_16079);
nand U17494 (N_17494,N_16167,N_16804);
nor U17495 (N_17495,N_16091,N_16406);
and U17496 (N_17496,N_16694,N_16127);
or U17497 (N_17497,N_16882,N_16910);
nand U17498 (N_17498,N_16151,N_16660);
xor U17499 (N_17499,N_16429,N_16426);
and U17500 (N_17500,N_16650,N_16368);
nand U17501 (N_17501,N_16169,N_16442);
xnor U17502 (N_17502,N_16550,N_16886);
xor U17503 (N_17503,N_16864,N_16991);
xnor U17504 (N_17504,N_16935,N_16711);
and U17505 (N_17505,N_16465,N_16777);
nor U17506 (N_17506,N_16864,N_16968);
and U17507 (N_17507,N_16006,N_16642);
xnor U17508 (N_17508,N_16592,N_16247);
xnor U17509 (N_17509,N_16074,N_16512);
nor U17510 (N_17510,N_16737,N_16165);
nand U17511 (N_17511,N_16061,N_16929);
nand U17512 (N_17512,N_16469,N_16409);
nand U17513 (N_17513,N_16616,N_16022);
and U17514 (N_17514,N_16953,N_16962);
xnor U17515 (N_17515,N_16141,N_16956);
xnor U17516 (N_17516,N_16259,N_16159);
nor U17517 (N_17517,N_16207,N_16858);
xnor U17518 (N_17518,N_16859,N_16136);
nand U17519 (N_17519,N_16501,N_16737);
and U17520 (N_17520,N_16652,N_16967);
xor U17521 (N_17521,N_16647,N_16477);
xnor U17522 (N_17522,N_16571,N_16669);
nor U17523 (N_17523,N_16123,N_16641);
nand U17524 (N_17524,N_16874,N_16827);
xnor U17525 (N_17525,N_16779,N_16269);
and U17526 (N_17526,N_16590,N_16156);
and U17527 (N_17527,N_16540,N_16282);
nand U17528 (N_17528,N_16732,N_16401);
nand U17529 (N_17529,N_16181,N_16396);
xor U17530 (N_17530,N_16172,N_16700);
nor U17531 (N_17531,N_16699,N_16334);
and U17532 (N_17532,N_16717,N_16917);
nor U17533 (N_17533,N_16076,N_16107);
nand U17534 (N_17534,N_16555,N_16813);
nand U17535 (N_17535,N_16786,N_16921);
nor U17536 (N_17536,N_16295,N_16516);
and U17537 (N_17537,N_16416,N_16516);
or U17538 (N_17538,N_16633,N_16145);
or U17539 (N_17539,N_16763,N_16992);
or U17540 (N_17540,N_16093,N_16233);
xnor U17541 (N_17541,N_16567,N_16445);
nand U17542 (N_17542,N_16268,N_16073);
or U17543 (N_17543,N_16125,N_16690);
and U17544 (N_17544,N_16558,N_16952);
nor U17545 (N_17545,N_16132,N_16618);
xor U17546 (N_17546,N_16661,N_16902);
or U17547 (N_17547,N_16848,N_16912);
or U17548 (N_17548,N_16611,N_16194);
or U17549 (N_17549,N_16846,N_16661);
or U17550 (N_17550,N_16856,N_16473);
and U17551 (N_17551,N_16806,N_16249);
nor U17552 (N_17552,N_16309,N_16318);
nand U17553 (N_17553,N_16071,N_16351);
nand U17554 (N_17554,N_16515,N_16373);
and U17555 (N_17555,N_16302,N_16737);
nand U17556 (N_17556,N_16214,N_16234);
xnor U17557 (N_17557,N_16888,N_16571);
xnor U17558 (N_17558,N_16240,N_16486);
nand U17559 (N_17559,N_16689,N_16733);
and U17560 (N_17560,N_16277,N_16712);
and U17561 (N_17561,N_16023,N_16787);
nor U17562 (N_17562,N_16572,N_16215);
and U17563 (N_17563,N_16752,N_16286);
xor U17564 (N_17564,N_16653,N_16915);
and U17565 (N_17565,N_16407,N_16553);
nor U17566 (N_17566,N_16955,N_16175);
xor U17567 (N_17567,N_16906,N_16248);
or U17568 (N_17568,N_16509,N_16229);
xor U17569 (N_17569,N_16142,N_16537);
or U17570 (N_17570,N_16678,N_16055);
nor U17571 (N_17571,N_16664,N_16869);
or U17572 (N_17572,N_16048,N_16244);
and U17573 (N_17573,N_16443,N_16242);
and U17574 (N_17574,N_16290,N_16391);
or U17575 (N_17575,N_16819,N_16958);
xor U17576 (N_17576,N_16336,N_16253);
nand U17577 (N_17577,N_16327,N_16430);
nor U17578 (N_17578,N_16957,N_16823);
and U17579 (N_17579,N_16180,N_16772);
xnor U17580 (N_17580,N_16489,N_16193);
and U17581 (N_17581,N_16020,N_16340);
xor U17582 (N_17582,N_16745,N_16254);
xnor U17583 (N_17583,N_16389,N_16711);
or U17584 (N_17584,N_16297,N_16358);
or U17585 (N_17585,N_16135,N_16367);
xnor U17586 (N_17586,N_16761,N_16555);
nor U17587 (N_17587,N_16327,N_16301);
nor U17588 (N_17588,N_16880,N_16245);
nor U17589 (N_17589,N_16376,N_16976);
or U17590 (N_17590,N_16584,N_16373);
or U17591 (N_17591,N_16397,N_16443);
and U17592 (N_17592,N_16953,N_16143);
and U17593 (N_17593,N_16304,N_16830);
xor U17594 (N_17594,N_16960,N_16821);
nand U17595 (N_17595,N_16988,N_16964);
or U17596 (N_17596,N_16260,N_16162);
nor U17597 (N_17597,N_16781,N_16291);
or U17598 (N_17598,N_16510,N_16133);
nand U17599 (N_17599,N_16060,N_16789);
nand U17600 (N_17600,N_16445,N_16128);
nand U17601 (N_17601,N_16820,N_16234);
and U17602 (N_17602,N_16964,N_16627);
nand U17603 (N_17603,N_16018,N_16803);
nor U17604 (N_17604,N_16886,N_16132);
or U17605 (N_17605,N_16829,N_16551);
nand U17606 (N_17606,N_16433,N_16977);
nor U17607 (N_17607,N_16861,N_16766);
nand U17608 (N_17608,N_16118,N_16797);
and U17609 (N_17609,N_16633,N_16264);
nor U17610 (N_17610,N_16073,N_16949);
nand U17611 (N_17611,N_16372,N_16402);
and U17612 (N_17612,N_16570,N_16785);
xnor U17613 (N_17613,N_16419,N_16991);
nand U17614 (N_17614,N_16371,N_16177);
and U17615 (N_17615,N_16025,N_16864);
nand U17616 (N_17616,N_16017,N_16157);
or U17617 (N_17617,N_16819,N_16470);
nand U17618 (N_17618,N_16777,N_16069);
nor U17619 (N_17619,N_16090,N_16856);
xnor U17620 (N_17620,N_16187,N_16425);
nor U17621 (N_17621,N_16594,N_16081);
or U17622 (N_17622,N_16872,N_16858);
and U17623 (N_17623,N_16540,N_16923);
or U17624 (N_17624,N_16359,N_16209);
nand U17625 (N_17625,N_16510,N_16614);
or U17626 (N_17626,N_16028,N_16862);
or U17627 (N_17627,N_16285,N_16083);
nand U17628 (N_17628,N_16680,N_16703);
and U17629 (N_17629,N_16904,N_16259);
nand U17630 (N_17630,N_16734,N_16148);
xor U17631 (N_17631,N_16631,N_16011);
nor U17632 (N_17632,N_16021,N_16745);
nor U17633 (N_17633,N_16265,N_16863);
nand U17634 (N_17634,N_16334,N_16083);
xnor U17635 (N_17635,N_16209,N_16596);
or U17636 (N_17636,N_16245,N_16813);
nor U17637 (N_17637,N_16151,N_16162);
nand U17638 (N_17638,N_16411,N_16312);
and U17639 (N_17639,N_16576,N_16256);
nand U17640 (N_17640,N_16302,N_16958);
nor U17641 (N_17641,N_16358,N_16305);
nand U17642 (N_17642,N_16362,N_16169);
nand U17643 (N_17643,N_16422,N_16644);
and U17644 (N_17644,N_16486,N_16828);
and U17645 (N_17645,N_16917,N_16972);
nand U17646 (N_17646,N_16950,N_16561);
nor U17647 (N_17647,N_16784,N_16064);
and U17648 (N_17648,N_16643,N_16913);
nor U17649 (N_17649,N_16405,N_16953);
and U17650 (N_17650,N_16846,N_16697);
xnor U17651 (N_17651,N_16910,N_16468);
nand U17652 (N_17652,N_16235,N_16272);
or U17653 (N_17653,N_16852,N_16397);
nand U17654 (N_17654,N_16427,N_16570);
nor U17655 (N_17655,N_16732,N_16132);
or U17656 (N_17656,N_16400,N_16517);
or U17657 (N_17657,N_16261,N_16626);
nand U17658 (N_17658,N_16789,N_16537);
or U17659 (N_17659,N_16537,N_16261);
or U17660 (N_17660,N_16869,N_16469);
nor U17661 (N_17661,N_16669,N_16883);
nand U17662 (N_17662,N_16007,N_16158);
and U17663 (N_17663,N_16804,N_16346);
nor U17664 (N_17664,N_16748,N_16867);
nand U17665 (N_17665,N_16031,N_16593);
nor U17666 (N_17666,N_16487,N_16171);
xor U17667 (N_17667,N_16758,N_16334);
nand U17668 (N_17668,N_16205,N_16562);
xnor U17669 (N_17669,N_16397,N_16653);
nor U17670 (N_17670,N_16264,N_16638);
nor U17671 (N_17671,N_16144,N_16041);
nor U17672 (N_17672,N_16287,N_16377);
nor U17673 (N_17673,N_16853,N_16469);
nor U17674 (N_17674,N_16886,N_16921);
xor U17675 (N_17675,N_16228,N_16311);
and U17676 (N_17676,N_16131,N_16611);
or U17677 (N_17677,N_16991,N_16805);
xor U17678 (N_17678,N_16401,N_16639);
xnor U17679 (N_17679,N_16450,N_16464);
or U17680 (N_17680,N_16107,N_16453);
xor U17681 (N_17681,N_16140,N_16776);
or U17682 (N_17682,N_16027,N_16045);
or U17683 (N_17683,N_16029,N_16556);
or U17684 (N_17684,N_16412,N_16869);
and U17685 (N_17685,N_16421,N_16278);
and U17686 (N_17686,N_16532,N_16374);
nand U17687 (N_17687,N_16710,N_16802);
xnor U17688 (N_17688,N_16352,N_16721);
nand U17689 (N_17689,N_16834,N_16570);
or U17690 (N_17690,N_16512,N_16871);
or U17691 (N_17691,N_16315,N_16303);
nand U17692 (N_17692,N_16034,N_16112);
and U17693 (N_17693,N_16531,N_16884);
xor U17694 (N_17694,N_16283,N_16254);
nand U17695 (N_17695,N_16131,N_16957);
and U17696 (N_17696,N_16907,N_16198);
nor U17697 (N_17697,N_16408,N_16587);
or U17698 (N_17698,N_16096,N_16194);
xnor U17699 (N_17699,N_16250,N_16364);
xnor U17700 (N_17700,N_16528,N_16715);
nor U17701 (N_17701,N_16883,N_16116);
xnor U17702 (N_17702,N_16731,N_16603);
or U17703 (N_17703,N_16243,N_16649);
and U17704 (N_17704,N_16163,N_16060);
or U17705 (N_17705,N_16274,N_16820);
or U17706 (N_17706,N_16662,N_16434);
nor U17707 (N_17707,N_16447,N_16974);
or U17708 (N_17708,N_16597,N_16100);
and U17709 (N_17709,N_16409,N_16300);
and U17710 (N_17710,N_16088,N_16308);
xor U17711 (N_17711,N_16858,N_16953);
and U17712 (N_17712,N_16305,N_16463);
or U17713 (N_17713,N_16674,N_16262);
nand U17714 (N_17714,N_16535,N_16477);
or U17715 (N_17715,N_16495,N_16439);
or U17716 (N_17716,N_16321,N_16566);
nor U17717 (N_17717,N_16863,N_16546);
nor U17718 (N_17718,N_16002,N_16039);
or U17719 (N_17719,N_16622,N_16716);
or U17720 (N_17720,N_16392,N_16896);
or U17721 (N_17721,N_16872,N_16890);
or U17722 (N_17722,N_16993,N_16141);
and U17723 (N_17723,N_16284,N_16734);
nor U17724 (N_17724,N_16625,N_16757);
nand U17725 (N_17725,N_16157,N_16585);
or U17726 (N_17726,N_16865,N_16607);
xnor U17727 (N_17727,N_16248,N_16025);
or U17728 (N_17728,N_16916,N_16814);
or U17729 (N_17729,N_16303,N_16406);
or U17730 (N_17730,N_16023,N_16799);
nor U17731 (N_17731,N_16744,N_16371);
nand U17732 (N_17732,N_16866,N_16713);
and U17733 (N_17733,N_16878,N_16234);
nor U17734 (N_17734,N_16427,N_16478);
nand U17735 (N_17735,N_16413,N_16357);
nor U17736 (N_17736,N_16790,N_16705);
xnor U17737 (N_17737,N_16846,N_16024);
xor U17738 (N_17738,N_16150,N_16538);
and U17739 (N_17739,N_16629,N_16303);
or U17740 (N_17740,N_16213,N_16603);
nor U17741 (N_17741,N_16114,N_16853);
nor U17742 (N_17742,N_16685,N_16285);
nand U17743 (N_17743,N_16311,N_16508);
nand U17744 (N_17744,N_16623,N_16005);
nand U17745 (N_17745,N_16078,N_16697);
xor U17746 (N_17746,N_16801,N_16005);
xor U17747 (N_17747,N_16289,N_16103);
or U17748 (N_17748,N_16047,N_16244);
xnor U17749 (N_17749,N_16498,N_16645);
or U17750 (N_17750,N_16876,N_16799);
nor U17751 (N_17751,N_16958,N_16459);
or U17752 (N_17752,N_16899,N_16801);
nand U17753 (N_17753,N_16307,N_16707);
xor U17754 (N_17754,N_16525,N_16390);
or U17755 (N_17755,N_16522,N_16948);
xor U17756 (N_17756,N_16448,N_16394);
or U17757 (N_17757,N_16759,N_16631);
nor U17758 (N_17758,N_16770,N_16991);
xnor U17759 (N_17759,N_16804,N_16364);
nand U17760 (N_17760,N_16768,N_16047);
nor U17761 (N_17761,N_16511,N_16073);
and U17762 (N_17762,N_16132,N_16104);
nor U17763 (N_17763,N_16984,N_16401);
nand U17764 (N_17764,N_16423,N_16017);
nor U17765 (N_17765,N_16581,N_16394);
xnor U17766 (N_17766,N_16277,N_16315);
xor U17767 (N_17767,N_16221,N_16860);
or U17768 (N_17768,N_16798,N_16521);
xnor U17769 (N_17769,N_16422,N_16238);
and U17770 (N_17770,N_16177,N_16158);
nand U17771 (N_17771,N_16867,N_16299);
nor U17772 (N_17772,N_16801,N_16558);
or U17773 (N_17773,N_16586,N_16972);
or U17774 (N_17774,N_16771,N_16039);
xnor U17775 (N_17775,N_16825,N_16302);
nor U17776 (N_17776,N_16309,N_16870);
or U17777 (N_17777,N_16875,N_16161);
or U17778 (N_17778,N_16708,N_16913);
and U17779 (N_17779,N_16998,N_16685);
nor U17780 (N_17780,N_16841,N_16693);
nand U17781 (N_17781,N_16127,N_16253);
xnor U17782 (N_17782,N_16882,N_16947);
and U17783 (N_17783,N_16858,N_16662);
xnor U17784 (N_17784,N_16816,N_16203);
xnor U17785 (N_17785,N_16391,N_16958);
xor U17786 (N_17786,N_16749,N_16263);
and U17787 (N_17787,N_16161,N_16296);
nor U17788 (N_17788,N_16370,N_16903);
and U17789 (N_17789,N_16727,N_16651);
and U17790 (N_17790,N_16097,N_16908);
xnor U17791 (N_17791,N_16404,N_16938);
xnor U17792 (N_17792,N_16215,N_16317);
xor U17793 (N_17793,N_16641,N_16025);
and U17794 (N_17794,N_16819,N_16180);
xnor U17795 (N_17795,N_16999,N_16221);
or U17796 (N_17796,N_16487,N_16482);
nand U17797 (N_17797,N_16662,N_16488);
and U17798 (N_17798,N_16732,N_16878);
nor U17799 (N_17799,N_16683,N_16072);
xnor U17800 (N_17800,N_16953,N_16939);
nor U17801 (N_17801,N_16599,N_16966);
xnor U17802 (N_17802,N_16155,N_16373);
and U17803 (N_17803,N_16655,N_16139);
and U17804 (N_17804,N_16779,N_16944);
nand U17805 (N_17805,N_16520,N_16426);
nor U17806 (N_17806,N_16333,N_16382);
xnor U17807 (N_17807,N_16210,N_16817);
xor U17808 (N_17808,N_16169,N_16022);
nor U17809 (N_17809,N_16268,N_16050);
or U17810 (N_17810,N_16370,N_16100);
xnor U17811 (N_17811,N_16098,N_16532);
nor U17812 (N_17812,N_16497,N_16415);
and U17813 (N_17813,N_16186,N_16819);
nand U17814 (N_17814,N_16690,N_16119);
xor U17815 (N_17815,N_16059,N_16870);
nand U17816 (N_17816,N_16437,N_16296);
nor U17817 (N_17817,N_16050,N_16619);
nand U17818 (N_17818,N_16282,N_16374);
nand U17819 (N_17819,N_16487,N_16714);
nor U17820 (N_17820,N_16692,N_16000);
and U17821 (N_17821,N_16126,N_16061);
nor U17822 (N_17822,N_16255,N_16254);
xnor U17823 (N_17823,N_16198,N_16288);
nor U17824 (N_17824,N_16732,N_16386);
or U17825 (N_17825,N_16412,N_16638);
and U17826 (N_17826,N_16466,N_16840);
nor U17827 (N_17827,N_16199,N_16485);
nand U17828 (N_17828,N_16674,N_16124);
or U17829 (N_17829,N_16993,N_16598);
and U17830 (N_17830,N_16399,N_16542);
nor U17831 (N_17831,N_16968,N_16822);
and U17832 (N_17832,N_16651,N_16098);
nor U17833 (N_17833,N_16932,N_16003);
or U17834 (N_17834,N_16891,N_16424);
and U17835 (N_17835,N_16250,N_16632);
or U17836 (N_17836,N_16286,N_16973);
xnor U17837 (N_17837,N_16538,N_16454);
xor U17838 (N_17838,N_16203,N_16349);
nor U17839 (N_17839,N_16607,N_16586);
or U17840 (N_17840,N_16816,N_16416);
nor U17841 (N_17841,N_16839,N_16123);
nor U17842 (N_17842,N_16186,N_16489);
or U17843 (N_17843,N_16642,N_16724);
nand U17844 (N_17844,N_16740,N_16130);
xnor U17845 (N_17845,N_16707,N_16390);
and U17846 (N_17846,N_16165,N_16935);
or U17847 (N_17847,N_16962,N_16591);
and U17848 (N_17848,N_16277,N_16736);
xor U17849 (N_17849,N_16398,N_16144);
and U17850 (N_17850,N_16961,N_16790);
and U17851 (N_17851,N_16031,N_16899);
nor U17852 (N_17852,N_16292,N_16137);
and U17853 (N_17853,N_16737,N_16073);
or U17854 (N_17854,N_16015,N_16949);
nand U17855 (N_17855,N_16543,N_16252);
nand U17856 (N_17856,N_16634,N_16633);
nor U17857 (N_17857,N_16989,N_16515);
nand U17858 (N_17858,N_16617,N_16170);
and U17859 (N_17859,N_16352,N_16365);
xnor U17860 (N_17860,N_16861,N_16155);
xnor U17861 (N_17861,N_16190,N_16249);
and U17862 (N_17862,N_16341,N_16950);
and U17863 (N_17863,N_16876,N_16760);
xnor U17864 (N_17864,N_16477,N_16882);
nor U17865 (N_17865,N_16431,N_16539);
nand U17866 (N_17866,N_16108,N_16252);
or U17867 (N_17867,N_16645,N_16043);
or U17868 (N_17868,N_16068,N_16904);
and U17869 (N_17869,N_16295,N_16977);
xor U17870 (N_17870,N_16674,N_16512);
or U17871 (N_17871,N_16530,N_16140);
nor U17872 (N_17872,N_16764,N_16269);
or U17873 (N_17873,N_16685,N_16971);
nor U17874 (N_17874,N_16330,N_16687);
xor U17875 (N_17875,N_16751,N_16034);
nand U17876 (N_17876,N_16500,N_16069);
nand U17877 (N_17877,N_16750,N_16796);
nor U17878 (N_17878,N_16964,N_16266);
nand U17879 (N_17879,N_16272,N_16803);
or U17880 (N_17880,N_16827,N_16978);
xnor U17881 (N_17881,N_16489,N_16347);
or U17882 (N_17882,N_16152,N_16213);
nand U17883 (N_17883,N_16029,N_16680);
xor U17884 (N_17884,N_16063,N_16804);
nand U17885 (N_17885,N_16340,N_16525);
or U17886 (N_17886,N_16697,N_16685);
or U17887 (N_17887,N_16785,N_16954);
or U17888 (N_17888,N_16632,N_16448);
or U17889 (N_17889,N_16783,N_16178);
and U17890 (N_17890,N_16976,N_16392);
or U17891 (N_17891,N_16320,N_16875);
nand U17892 (N_17892,N_16106,N_16017);
or U17893 (N_17893,N_16419,N_16768);
xor U17894 (N_17894,N_16834,N_16897);
nand U17895 (N_17895,N_16751,N_16667);
and U17896 (N_17896,N_16060,N_16188);
nor U17897 (N_17897,N_16696,N_16559);
or U17898 (N_17898,N_16174,N_16117);
nand U17899 (N_17899,N_16485,N_16848);
nor U17900 (N_17900,N_16895,N_16973);
or U17901 (N_17901,N_16649,N_16502);
nand U17902 (N_17902,N_16986,N_16466);
or U17903 (N_17903,N_16047,N_16392);
or U17904 (N_17904,N_16299,N_16856);
nor U17905 (N_17905,N_16238,N_16079);
nor U17906 (N_17906,N_16059,N_16846);
nand U17907 (N_17907,N_16267,N_16133);
xnor U17908 (N_17908,N_16540,N_16685);
xnor U17909 (N_17909,N_16344,N_16332);
nor U17910 (N_17910,N_16332,N_16769);
and U17911 (N_17911,N_16978,N_16023);
or U17912 (N_17912,N_16614,N_16778);
nand U17913 (N_17913,N_16144,N_16251);
xnor U17914 (N_17914,N_16223,N_16361);
nor U17915 (N_17915,N_16019,N_16172);
and U17916 (N_17916,N_16457,N_16152);
nand U17917 (N_17917,N_16003,N_16439);
nand U17918 (N_17918,N_16658,N_16362);
xnor U17919 (N_17919,N_16444,N_16421);
nor U17920 (N_17920,N_16616,N_16179);
xnor U17921 (N_17921,N_16104,N_16451);
and U17922 (N_17922,N_16029,N_16875);
nand U17923 (N_17923,N_16441,N_16497);
nand U17924 (N_17924,N_16167,N_16318);
and U17925 (N_17925,N_16982,N_16409);
and U17926 (N_17926,N_16812,N_16351);
nand U17927 (N_17927,N_16217,N_16937);
xor U17928 (N_17928,N_16783,N_16766);
and U17929 (N_17929,N_16262,N_16848);
or U17930 (N_17930,N_16917,N_16695);
xnor U17931 (N_17931,N_16765,N_16577);
nor U17932 (N_17932,N_16015,N_16763);
xnor U17933 (N_17933,N_16880,N_16346);
and U17934 (N_17934,N_16174,N_16277);
and U17935 (N_17935,N_16798,N_16461);
nand U17936 (N_17936,N_16254,N_16269);
xnor U17937 (N_17937,N_16900,N_16983);
nor U17938 (N_17938,N_16433,N_16096);
nand U17939 (N_17939,N_16646,N_16874);
nand U17940 (N_17940,N_16471,N_16916);
or U17941 (N_17941,N_16356,N_16388);
and U17942 (N_17942,N_16504,N_16578);
and U17943 (N_17943,N_16072,N_16488);
and U17944 (N_17944,N_16769,N_16920);
and U17945 (N_17945,N_16548,N_16072);
and U17946 (N_17946,N_16709,N_16931);
and U17947 (N_17947,N_16935,N_16508);
nor U17948 (N_17948,N_16100,N_16089);
and U17949 (N_17949,N_16126,N_16440);
xnor U17950 (N_17950,N_16762,N_16572);
and U17951 (N_17951,N_16263,N_16103);
and U17952 (N_17952,N_16300,N_16188);
nor U17953 (N_17953,N_16476,N_16469);
xnor U17954 (N_17954,N_16901,N_16027);
nand U17955 (N_17955,N_16452,N_16006);
or U17956 (N_17956,N_16807,N_16558);
or U17957 (N_17957,N_16135,N_16199);
and U17958 (N_17958,N_16241,N_16875);
or U17959 (N_17959,N_16545,N_16419);
nand U17960 (N_17960,N_16093,N_16341);
xnor U17961 (N_17961,N_16874,N_16982);
nand U17962 (N_17962,N_16577,N_16338);
nand U17963 (N_17963,N_16359,N_16331);
and U17964 (N_17964,N_16170,N_16159);
and U17965 (N_17965,N_16792,N_16746);
and U17966 (N_17966,N_16971,N_16655);
xor U17967 (N_17967,N_16750,N_16887);
nor U17968 (N_17968,N_16277,N_16100);
nor U17969 (N_17969,N_16126,N_16288);
or U17970 (N_17970,N_16156,N_16044);
xnor U17971 (N_17971,N_16800,N_16257);
xor U17972 (N_17972,N_16605,N_16930);
nand U17973 (N_17973,N_16705,N_16673);
and U17974 (N_17974,N_16723,N_16025);
nand U17975 (N_17975,N_16050,N_16664);
and U17976 (N_17976,N_16480,N_16705);
xnor U17977 (N_17977,N_16197,N_16104);
and U17978 (N_17978,N_16966,N_16214);
or U17979 (N_17979,N_16138,N_16571);
and U17980 (N_17980,N_16345,N_16313);
nor U17981 (N_17981,N_16850,N_16752);
and U17982 (N_17982,N_16800,N_16685);
and U17983 (N_17983,N_16616,N_16114);
nor U17984 (N_17984,N_16934,N_16285);
nand U17985 (N_17985,N_16529,N_16306);
nor U17986 (N_17986,N_16710,N_16415);
xor U17987 (N_17987,N_16947,N_16084);
nand U17988 (N_17988,N_16892,N_16010);
nor U17989 (N_17989,N_16868,N_16682);
xnor U17990 (N_17990,N_16357,N_16458);
xnor U17991 (N_17991,N_16199,N_16974);
or U17992 (N_17992,N_16266,N_16907);
or U17993 (N_17993,N_16168,N_16637);
nor U17994 (N_17994,N_16908,N_16437);
and U17995 (N_17995,N_16949,N_16848);
or U17996 (N_17996,N_16574,N_16454);
xnor U17997 (N_17997,N_16195,N_16127);
or U17998 (N_17998,N_16761,N_16627);
and U17999 (N_17999,N_16742,N_16829);
nand U18000 (N_18000,N_17759,N_17947);
nor U18001 (N_18001,N_17832,N_17580);
xnor U18002 (N_18002,N_17754,N_17084);
or U18003 (N_18003,N_17596,N_17955);
or U18004 (N_18004,N_17593,N_17862);
xnor U18005 (N_18005,N_17121,N_17150);
xnor U18006 (N_18006,N_17119,N_17191);
and U18007 (N_18007,N_17679,N_17309);
nand U18008 (N_18008,N_17196,N_17108);
nand U18009 (N_18009,N_17723,N_17939);
xnor U18010 (N_18010,N_17384,N_17612);
nand U18011 (N_18011,N_17331,N_17681);
nand U18012 (N_18012,N_17987,N_17020);
nand U18013 (N_18013,N_17653,N_17619);
or U18014 (N_18014,N_17787,N_17005);
and U18015 (N_18015,N_17297,N_17184);
xnor U18016 (N_18016,N_17595,N_17290);
xor U18017 (N_18017,N_17490,N_17823);
or U18018 (N_18018,N_17994,N_17684);
xnor U18019 (N_18019,N_17537,N_17019);
and U18020 (N_18020,N_17457,N_17228);
and U18021 (N_18021,N_17935,N_17948);
nor U18022 (N_18022,N_17086,N_17934);
xor U18023 (N_18023,N_17039,N_17986);
or U18024 (N_18024,N_17971,N_17784);
or U18025 (N_18025,N_17185,N_17911);
or U18026 (N_18026,N_17786,N_17954);
nand U18027 (N_18027,N_17928,N_17422);
nand U18028 (N_18028,N_17300,N_17138);
or U18029 (N_18029,N_17673,N_17703);
or U18030 (N_18030,N_17852,N_17391);
nand U18031 (N_18031,N_17842,N_17743);
nand U18032 (N_18032,N_17072,N_17804);
and U18033 (N_18033,N_17508,N_17449);
nor U18034 (N_18034,N_17085,N_17912);
or U18035 (N_18035,N_17492,N_17690);
or U18036 (N_18036,N_17937,N_17231);
or U18037 (N_18037,N_17791,N_17818);
or U18038 (N_18038,N_17843,N_17240);
nand U18039 (N_18039,N_17658,N_17340);
nor U18040 (N_18040,N_17571,N_17888);
nand U18041 (N_18041,N_17182,N_17963);
xnor U18042 (N_18042,N_17124,N_17661);
nand U18043 (N_18043,N_17411,N_17962);
nand U18044 (N_18044,N_17193,N_17311);
nor U18045 (N_18045,N_17866,N_17822);
nor U18046 (N_18046,N_17825,N_17079);
nand U18047 (N_18047,N_17172,N_17988);
xnor U18048 (N_18048,N_17530,N_17914);
xor U18049 (N_18049,N_17610,N_17874);
xor U18050 (N_18050,N_17414,N_17499);
nor U18051 (N_18051,N_17348,N_17943);
nand U18052 (N_18052,N_17400,N_17873);
xor U18053 (N_18053,N_17143,N_17261);
or U18054 (N_18054,N_17260,N_17718);
nand U18055 (N_18055,N_17753,N_17775);
xnor U18056 (N_18056,N_17513,N_17237);
xor U18057 (N_18057,N_17051,N_17274);
and U18058 (N_18058,N_17905,N_17915);
and U18059 (N_18059,N_17324,N_17033);
xor U18060 (N_18060,N_17319,N_17314);
and U18061 (N_18061,N_17996,N_17900);
xor U18062 (N_18062,N_17253,N_17587);
xnor U18063 (N_18063,N_17533,N_17696);
nor U18064 (N_18064,N_17840,N_17399);
xor U18065 (N_18065,N_17747,N_17047);
nand U18066 (N_18066,N_17878,N_17369);
nor U18067 (N_18067,N_17337,N_17173);
nand U18068 (N_18068,N_17484,N_17567);
and U18069 (N_18069,N_17927,N_17975);
nand U18070 (N_18070,N_17305,N_17437);
nand U18071 (N_18071,N_17083,N_17286);
nand U18072 (N_18072,N_17435,N_17313);
xor U18073 (N_18073,N_17930,N_17220);
xnor U18074 (N_18074,N_17575,N_17224);
and U18075 (N_18075,N_17027,N_17054);
or U18076 (N_18076,N_17758,N_17712);
or U18077 (N_18077,N_17504,N_17371);
nor U18078 (N_18078,N_17110,N_17133);
xor U18079 (N_18079,N_17769,N_17557);
or U18080 (N_18080,N_17764,N_17739);
or U18081 (N_18081,N_17746,N_17024);
xor U18082 (N_18082,N_17957,N_17232);
nor U18083 (N_18083,N_17989,N_17613);
nor U18084 (N_18084,N_17132,N_17330);
and U18085 (N_18085,N_17523,N_17071);
and U18086 (N_18086,N_17856,N_17001);
and U18087 (N_18087,N_17181,N_17545);
or U18088 (N_18088,N_17548,N_17230);
xor U18089 (N_18089,N_17158,N_17826);
nor U18090 (N_18090,N_17385,N_17099);
nand U18091 (N_18091,N_17360,N_17502);
and U18092 (N_18092,N_17810,N_17461);
nor U18093 (N_18093,N_17570,N_17303);
or U18094 (N_18094,N_17168,N_17659);
and U18095 (N_18095,N_17773,N_17456);
xnor U18096 (N_18096,N_17316,N_17419);
nor U18097 (N_18097,N_17816,N_17332);
and U18098 (N_18098,N_17387,N_17388);
and U18099 (N_18099,N_17701,N_17302);
and U18100 (N_18100,N_17800,N_17632);
or U18101 (N_18101,N_17736,N_17973);
or U18102 (N_18102,N_17691,N_17091);
nor U18103 (N_18103,N_17453,N_17445);
nor U18104 (N_18104,N_17689,N_17926);
xnor U18105 (N_18105,N_17827,N_17134);
nand U18106 (N_18106,N_17563,N_17644);
xor U18107 (N_18107,N_17640,N_17722);
and U18108 (N_18108,N_17846,N_17105);
nor U18109 (N_18109,N_17361,N_17217);
nand U18110 (N_18110,N_17126,N_17117);
xor U18111 (N_18111,N_17817,N_17294);
nor U18112 (N_18112,N_17030,N_17569);
xnor U18113 (N_18113,N_17062,N_17656);
or U18114 (N_18114,N_17732,N_17997);
nand U18115 (N_18115,N_17426,N_17917);
xor U18116 (N_18116,N_17269,N_17544);
nor U18117 (N_18117,N_17886,N_17284);
nor U18118 (N_18118,N_17541,N_17931);
or U18119 (N_18119,N_17093,N_17296);
or U18120 (N_18120,N_17946,N_17783);
nand U18121 (N_18121,N_17667,N_17519);
and U18122 (N_18122,N_17098,N_17861);
nand U18123 (N_18123,N_17795,N_17710);
nand U18124 (N_18124,N_17851,N_17467);
or U18125 (N_18125,N_17552,N_17892);
or U18126 (N_18126,N_17351,N_17500);
xnor U18127 (N_18127,N_17985,N_17708);
and U18128 (N_18128,N_17762,N_17607);
or U18129 (N_18129,N_17245,N_17442);
or U18130 (N_18130,N_17497,N_17950);
nand U18131 (N_18131,N_17568,N_17899);
nor U18132 (N_18132,N_17199,N_17068);
nand U18133 (N_18133,N_17958,N_17518);
nor U18134 (N_18134,N_17944,N_17287);
nand U18135 (N_18135,N_17668,N_17207);
nor U18136 (N_18136,N_17216,N_17932);
xor U18137 (N_18137,N_17893,N_17829);
and U18138 (N_18138,N_17647,N_17967);
nor U18139 (N_18139,N_17774,N_17789);
nand U18140 (N_18140,N_17195,N_17562);
and U18141 (N_18141,N_17772,N_17582);
xnor U18142 (N_18142,N_17321,N_17771);
xnor U18143 (N_18143,N_17646,N_17009);
nand U18144 (N_18144,N_17410,N_17729);
and U18145 (N_18145,N_17142,N_17394);
or U18146 (N_18146,N_17853,N_17601);
and U18147 (N_18147,N_17560,N_17599);
xnor U18148 (N_18148,N_17909,N_17821);
and U18149 (N_18149,N_17365,N_17163);
nand U18150 (N_18150,N_17836,N_17877);
nand U18151 (N_18151,N_17976,N_17700);
nand U18152 (N_18152,N_17278,N_17586);
and U18153 (N_18153,N_17424,N_17811);
nor U18154 (N_18154,N_17263,N_17841);
or U18155 (N_18155,N_17855,N_17782);
nand U18156 (N_18156,N_17995,N_17210);
or U18157 (N_18157,N_17686,N_17551);
or U18158 (N_18158,N_17285,N_17355);
and U18159 (N_18159,N_17487,N_17397);
nand U18160 (N_18160,N_17112,N_17434);
nor U18161 (N_18161,N_17517,N_17413);
nor U18162 (N_18162,N_17022,N_17336);
xor U18163 (N_18163,N_17326,N_17250);
xor U18164 (N_18164,N_17585,N_17222);
nor U18165 (N_18165,N_17695,N_17243);
or U18166 (N_18166,N_17777,N_17289);
and U18167 (N_18167,N_17699,N_17167);
nor U18168 (N_18168,N_17312,N_17378);
or U18169 (N_18169,N_17583,N_17357);
nand U18170 (N_18170,N_17735,N_17096);
and U18171 (N_18171,N_17961,N_17629);
or U18172 (N_18172,N_17706,N_17871);
nor U18173 (N_18173,N_17055,N_17614);
or U18174 (N_18174,N_17042,N_17409);
nand U18175 (N_18175,N_17574,N_17145);
xor U18176 (N_18176,N_17443,N_17641);
xnor U18177 (N_18177,N_17002,N_17180);
xnor U18178 (N_18178,N_17881,N_17494);
nand U18179 (N_18179,N_17952,N_17916);
and U18180 (N_18180,N_17671,N_17526);
xnor U18181 (N_18181,N_17919,N_17910);
nand U18182 (N_18182,N_17465,N_17209);
xor U18183 (N_18183,N_17863,N_17577);
or U18184 (N_18184,N_17999,N_17187);
nor U18185 (N_18185,N_17432,N_17064);
nand U18186 (N_18186,N_17488,N_17704);
or U18187 (N_18187,N_17707,N_17186);
xor U18188 (N_18188,N_17462,N_17156);
xor U18189 (N_18189,N_17146,N_17651);
or U18190 (N_18190,N_17713,N_17724);
nor U18191 (N_18191,N_17923,N_17628);
or U18192 (N_18192,N_17404,N_17719);
xnor U18193 (N_18193,N_17320,N_17493);
nor U18194 (N_18194,N_17130,N_17776);
and U18195 (N_18195,N_17244,N_17978);
and U18196 (N_18196,N_17377,N_17048);
nor U18197 (N_18197,N_17779,N_17547);
nand U18198 (N_18198,N_17844,N_17660);
and U18199 (N_18199,N_17430,N_17839);
nand U18200 (N_18200,N_17714,N_17023);
nor U18201 (N_18201,N_17676,N_17534);
xor U18202 (N_18202,N_17597,N_17740);
and U18203 (N_18203,N_17591,N_17342);
xor U18204 (N_18204,N_17137,N_17299);
and U18205 (N_18205,N_17383,N_17848);
and U18206 (N_18206,N_17011,N_17218);
or U18207 (N_18207,N_17466,N_17233);
nor U18208 (N_18208,N_17389,N_17643);
xnor U18209 (N_18209,N_17868,N_17352);
nor U18210 (N_18210,N_17529,N_17440);
nor U18211 (N_18211,N_17760,N_17205);
or U18212 (N_18212,N_17428,N_17041);
and U18213 (N_18213,N_17749,N_17705);
xnor U18214 (N_18214,N_17206,N_17398);
nand U18215 (N_18215,N_17179,N_17883);
nor U18216 (N_18216,N_17857,N_17665);
xor U18217 (N_18217,N_17716,N_17157);
and U18218 (N_18218,N_17590,N_17675);
and U18219 (N_18219,N_17604,N_17390);
xor U18220 (N_18220,N_17439,N_17095);
and U18221 (N_18221,N_17505,N_17252);
or U18222 (N_18222,N_17584,N_17869);
nor U18223 (N_18223,N_17188,N_17970);
xor U18224 (N_18224,N_17446,N_17213);
nor U18225 (N_18225,N_17837,N_17247);
and U18226 (N_18226,N_17160,N_17630);
and U18227 (N_18227,N_17097,N_17315);
xor U18228 (N_18228,N_17026,N_17964);
and U18229 (N_18229,N_17801,N_17329);
and U18230 (N_18230,N_17876,N_17059);
and U18231 (N_18231,N_17201,N_17692);
and U18232 (N_18232,N_17304,N_17662);
nand U18233 (N_18233,N_17983,N_17203);
and U18234 (N_18234,N_17219,N_17564);
or U18235 (N_18235,N_17008,N_17347);
xor U18236 (N_18236,N_17645,N_17012);
xor U18237 (N_18237,N_17128,N_17685);
nand U18238 (N_18238,N_17364,N_17589);
and U18239 (N_18239,N_17058,N_17566);
xor U18240 (N_18240,N_17004,N_17460);
nor U18241 (N_18241,N_17122,N_17765);
xor U18242 (N_18242,N_17929,N_17473);
nor U18243 (N_18243,N_17170,N_17264);
and U18244 (N_18244,N_17458,N_17674);
or U18245 (N_18245,N_17366,N_17524);
nand U18246 (N_18246,N_17509,N_17745);
or U18247 (N_18247,N_17021,N_17949);
or U18248 (N_18248,N_17522,N_17100);
nand U18249 (N_18249,N_17034,N_17794);
or U18250 (N_18250,N_17543,N_17682);
nor U18251 (N_18251,N_17808,N_17993);
nor U18252 (N_18252,N_17406,N_17858);
nor U18253 (N_18253,N_17813,N_17924);
xnor U18254 (N_18254,N_17942,N_17281);
and U18255 (N_18255,N_17438,N_17270);
xor U18256 (N_18256,N_17968,N_17491);
nor U18257 (N_18257,N_17666,N_17379);
nor U18258 (N_18258,N_17756,N_17239);
nor U18259 (N_18259,N_17652,N_17087);
and U18260 (N_18260,N_17781,N_17073);
nor U18261 (N_18261,N_17074,N_17835);
and U18262 (N_18262,N_17080,N_17057);
or U18263 (N_18263,N_17828,N_17452);
and U18264 (N_18264,N_17344,N_17697);
nand U18265 (N_18265,N_17238,N_17531);
xnor U18266 (N_18266,N_17907,N_17190);
and U18267 (N_18267,N_17370,N_17757);
or U18268 (N_18268,N_17895,N_17367);
or U18269 (N_18269,N_17657,N_17918);
nand U18270 (N_18270,N_17265,N_17798);
or U18271 (N_18271,N_17556,N_17401);
nand U18272 (N_18272,N_17755,N_17214);
nor U18273 (N_18273,N_17965,N_17104);
and U18274 (N_18274,N_17600,N_17903);
xnor U18275 (N_18275,N_17511,N_17474);
xnor U18276 (N_18276,N_17625,N_17793);
or U18277 (N_18277,N_17885,N_17386);
nand U18278 (N_18278,N_17788,N_17578);
nor U18279 (N_18279,N_17730,N_17468);
xor U18280 (N_18280,N_17197,N_17129);
nor U18281 (N_18281,N_17200,N_17737);
xor U18282 (N_18282,N_17972,N_17242);
and U18283 (N_18283,N_17075,N_17166);
and U18284 (N_18284,N_17249,N_17815);
and U18285 (N_18285,N_17992,N_17901);
and U18286 (N_18286,N_17154,N_17115);
and U18287 (N_18287,N_17392,N_17444);
xor U18288 (N_18288,N_17183,N_17687);
or U18289 (N_18289,N_17018,N_17295);
nand U18290 (N_18290,N_17481,N_17017);
xnor U18291 (N_18291,N_17626,N_17381);
xor U18292 (N_18292,N_17717,N_17000);
or U18293 (N_18293,N_17272,N_17951);
nor U18294 (N_18294,N_17709,N_17898);
or U18295 (N_18295,N_17880,N_17506);
nand U18296 (N_18296,N_17616,N_17617);
and U18297 (N_18297,N_17078,N_17663);
nand U18298 (N_18298,N_17540,N_17807);
xnor U18299 (N_18299,N_17982,N_17149);
and U18300 (N_18300,N_17454,N_17007);
nor U18301 (N_18301,N_17711,N_17094);
nor U18302 (N_18302,N_17338,N_17169);
or U18303 (N_18303,N_17472,N_17120);
nand U18304 (N_18304,N_17559,N_17380);
and U18305 (N_18305,N_17480,N_17485);
or U18306 (N_18306,N_17376,N_17118);
xor U18307 (N_18307,N_17744,N_17748);
xnor U18308 (N_18308,N_17867,N_17192);
or U18309 (N_18309,N_17553,N_17627);
and U18310 (N_18310,N_17353,N_17897);
nand U18311 (N_18311,N_17198,N_17050);
nand U18312 (N_18312,N_17956,N_17592);
nor U18313 (N_18313,N_17266,N_17208);
nor U18314 (N_18314,N_17922,N_17114);
nand U18315 (N_18315,N_17849,N_17279);
xnor U18316 (N_18316,N_17036,N_17891);
nor U18317 (N_18317,N_17417,N_17546);
or U18318 (N_18318,N_17693,N_17780);
or U18319 (N_18319,N_17479,N_17980);
xor U18320 (N_18320,N_17865,N_17148);
or U18321 (N_18321,N_17362,N_17741);
nor U18322 (N_18322,N_17268,N_17101);
nor U18323 (N_18323,N_17043,N_17555);
nand U18324 (N_18324,N_17423,N_17532);
nor U18325 (N_18325,N_17766,N_17953);
and U18326 (N_18326,N_17257,N_17291);
and U18327 (N_18327,N_17408,N_17678);
or U18328 (N_18328,N_17715,N_17175);
or U18329 (N_18329,N_17609,N_17637);
nor U18330 (N_18330,N_17921,N_17421);
nand U18331 (N_18331,N_17763,N_17561);
xor U18332 (N_18332,N_17292,N_17622);
and U18333 (N_18333,N_17516,N_17139);
nand U18334 (N_18334,N_17611,N_17650);
xor U18335 (N_18335,N_17450,N_17368);
nand U18336 (N_18336,N_17136,N_17038);
and U18337 (N_18337,N_17259,N_17416);
nand U18338 (N_18338,N_17677,N_17824);
xor U18339 (N_18339,N_17334,N_17029);
and U18340 (N_18340,N_17447,N_17694);
or U18341 (N_18341,N_17945,N_17061);
and U18342 (N_18342,N_17670,N_17752);
and U18343 (N_18343,N_17306,N_17418);
or U18344 (N_18344,N_17615,N_17672);
nor U18345 (N_18345,N_17464,N_17135);
nand U18346 (N_18346,N_17335,N_17698);
xnor U18347 (N_18347,N_17803,N_17106);
nor U18348 (N_18348,N_17525,N_17477);
or U18349 (N_18349,N_17991,N_17407);
nand U18350 (N_18350,N_17236,N_17860);
or U18351 (N_18351,N_17037,N_17496);
nand U18352 (N_18352,N_17427,N_17204);
or U18353 (N_18353,N_17702,N_17006);
nand U18354 (N_18354,N_17116,N_17960);
nand U18355 (N_18355,N_17280,N_17805);
or U18356 (N_18356,N_17634,N_17177);
and U18357 (N_18357,N_17016,N_17429);
nand U18358 (N_18358,N_17638,N_17489);
or U18359 (N_18359,N_17354,N_17107);
or U18360 (N_18360,N_17171,N_17202);
nor U18361 (N_18361,N_17345,N_17738);
nor U18362 (N_18362,N_17872,N_17273);
nand U18363 (N_18363,N_17014,N_17904);
and U18364 (N_18364,N_17212,N_17831);
nor U18365 (N_18365,N_17322,N_17598);
nand U18366 (N_18366,N_17293,N_17141);
or U18367 (N_18367,N_17520,N_17325);
nand U18368 (N_18368,N_17984,N_17402);
nor U18369 (N_18369,N_17113,N_17875);
or U18370 (N_18370,N_17870,N_17307);
nor U18371 (N_18371,N_17475,N_17375);
nor U18372 (N_18372,N_17642,N_17503);
xor U18373 (N_18373,N_17979,N_17809);
xnor U18374 (N_18374,N_17153,N_17028);
or U18375 (N_18375,N_17536,N_17636);
nand U18376 (N_18376,N_17317,N_17550);
xor U18377 (N_18377,N_17221,N_17301);
nand U18378 (N_18378,N_17393,N_17833);
xnor U18379 (N_18379,N_17654,N_17558);
nand U18380 (N_18380,N_17147,N_17065);
nor U18381 (N_18381,N_17358,N_17267);
and U18382 (N_18382,N_17013,N_17069);
or U18383 (N_18383,N_17602,N_17298);
or U18384 (N_18384,N_17814,N_17076);
nor U18385 (N_18385,N_17581,N_17731);
nand U18386 (N_18386,N_17189,N_17415);
nor U18387 (N_18387,N_17246,N_17123);
nor U18388 (N_18388,N_17925,N_17178);
xnor U18389 (N_18389,N_17031,N_17648);
nor U18390 (N_18390,N_17639,N_17834);
nand U18391 (N_18391,N_17799,N_17056);
and U18392 (N_18392,N_17433,N_17588);
nor U18393 (N_18393,N_17633,N_17721);
and U18394 (N_18394,N_17174,N_17151);
nand U18395 (N_18395,N_17277,N_17276);
nor U18396 (N_18396,N_17092,N_17425);
and U18397 (N_18397,N_17283,N_17431);
and U18398 (N_18398,N_17346,N_17288);
and U18399 (N_18399,N_17920,N_17887);
xor U18400 (N_18400,N_17327,N_17412);
xnor U18401 (N_18401,N_17908,N_17229);
xor U18402 (N_18402,N_17608,N_17081);
nand U18403 (N_18403,N_17211,N_17469);
or U18404 (N_18404,N_17161,N_17049);
nand U18405 (N_18405,N_17063,N_17554);
or U18406 (N_18406,N_17720,N_17850);
and U18407 (N_18407,N_17045,N_17785);
nor U18408 (N_18408,N_17688,N_17089);
or U18409 (N_18409,N_17339,N_17549);
nor U18410 (N_18410,N_17356,N_17941);
or U18411 (N_18411,N_17215,N_17535);
or U18412 (N_18412,N_17164,N_17683);
nor U18413 (N_18413,N_17734,N_17470);
nand U18414 (N_18414,N_17066,N_17176);
nand U18415 (N_18415,N_17802,N_17070);
and U18416 (N_18416,N_17728,N_17884);
or U18417 (N_18417,N_17420,N_17792);
nand U18418 (N_18418,N_17889,N_17990);
xnor U18419 (N_18419,N_17859,N_17981);
xor U18420 (N_18420,N_17864,N_17271);
nand U18421 (N_18421,N_17998,N_17374);
nor U18422 (N_18422,N_17538,N_17977);
and U18423 (N_18423,N_17631,N_17894);
or U18424 (N_18424,N_17082,N_17372);
and U18425 (N_18425,N_17605,N_17936);
nor U18426 (N_18426,N_17512,N_17155);
nor U18427 (N_18427,N_17680,N_17282);
xnor U18428 (N_18428,N_17090,N_17539);
or U18429 (N_18429,N_17498,N_17254);
xnor U18430 (N_18430,N_17733,N_17655);
xor U18431 (N_18431,N_17767,N_17256);
and U18432 (N_18432,N_17225,N_17618);
nand U18433 (N_18433,N_17275,N_17241);
nand U18434 (N_18434,N_17103,N_17742);
nor U18435 (N_18435,N_17726,N_17528);
xnor U18436 (N_18436,N_17255,N_17165);
or U18437 (N_18437,N_17323,N_17025);
nor U18438 (N_18438,N_17162,N_17603);
nor U18439 (N_18439,N_17521,N_17879);
nand U18440 (N_18440,N_17797,N_17770);
and U18441 (N_18441,N_17594,N_17507);
xor U18442 (N_18442,N_17373,N_17812);
xor U18443 (N_18443,N_17969,N_17258);
or U18444 (N_18444,N_17318,N_17436);
or U18445 (N_18445,N_17902,N_17664);
and U18446 (N_18446,N_17478,N_17396);
or U18447 (N_18447,N_17966,N_17542);
xor U18448 (N_18448,N_17035,N_17565);
nand U18449 (N_18449,N_17959,N_17194);
and U18450 (N_18450,N_17913,N_17350);
or U18451 (N_18451,N_17854,N_17111);
xor U18452 (N_18452,N_17819,N_17234);
nor U18453 (N_18453,N_17761,N_17649);
nand U18454 (N_18454,N_17144,N_17363);
or U18455 (N_18455,N_17838,N_17003);
and U18456 (N_18456,N_17044,N_17806);
and U18457 (N_18457,N_17455,N_17040);
nor U18458 (N_18458,N_17890,N_17974);
nor U18459 (N_18459,N_17403,N_17778);
or U18460 (N_18460,N_17343,N_17750);
nor U18461 (N_18461,N_17606,N_17441);
or U18462 (N_18462,N_17052,N_17088);
nor U18463 (N_18463,N_17906,N_17152);
nor U18464 (N_18464,N_17333,N_17576);
nor U18465 (N_18465,N_17127,N_17067);
and U18466 (N_18466,N_17405,N_17463);
or U18467 (N_18467,N_17046,N_17933);
or U18468 (N_18468,N_17235,N_17109);
xnor U18469 (N_18469,N_17882,N_17010);
nor U18470 (N_18470,N_17725,N_17077);
nor U18471 (N_18471,N_17125,N_17451);
nor U18472 (N_18472,N_17471,N_17845);
xnor U18473 (N_18473,N_17573,N_17032);
and U18474 (N_18474,N_17341,N_17830);
nor U18475 (N_18475,N_17248,N_17620);
xor U18476 (N_18476,N_17820,N_17768);
nor U18477 (N_18477,N_17940,N_17053);
or U18478 (N_18478,N_17482,N_17159);
or U18479 (N_18479,N_17495,N_17140);
or U18480 (N_18480,N_17476,N_17310);
and U18481 (N_18481,N_17251,N_17448);
and U18482 (N_18482,N_17359,N_17015);
nor U18483 (N_18483,N_17486,N_17727);
xor U18484 (N_18484,N_17382,N_17102);
and U18485 (N_18485,N_17514,N_17262);
and U18486 (N_18486,N_17227,N_17510);
nand U18487 (N_18487,N_17060,N_17226);
nor U18488 (N_18488,N_17624,N_17223);
xnor U18489 (N_18489,N_17796,N_17790);
and U18490 (N_18490,N_17395,N_17131);
or U18491 (N_18491,N_17459,N_17847);
and U18492 (N_18492,N_17328,N_17579);
nand U18493 (N_18493,N_17623,N_17527);
xnor U18494 (N_18494,N_17669,N_17751);
and U18495 (N_18495,N_17308,N_17896);
or U18496 (N_18496,N_17635,N_17572);
or U18497 (N_18497,N_17621,N_17501);
xor U18498 (N_18498,N_17938,N_17349);
nor U18499 (N_18499,N_17483,N_17515);
or U18500 (N_18500,N_17406,N_17898);
and U18501 (N_18501,N_17582,N_17403);
xnor U18502 (N_18502,N_17980,N_17138);
xnor U18503 (N_18503,N_17504,N_17672);
and U18504 (N_18504,N_17283,N_17433);
or U18505 (N_18505,N_17787,N_17080);
and U18506 (N_18506,N_17988,N_17672);
nand U18507 (N_18507,N_17526,N_17414);
and U18508 (N_18508,N_17714,N_17540);
nor U18509 (N_18509,N_17958,N_17349);
nor U18510 (N_18510,N_17109,N_17123);
nor U18511 (N_18511,N_17567,N_17066);
and U18512 (N_18512,N_17157,N_17267);
nor U18513 (N_18513,N_17349,N_17916);
xor U18514 (N_18514,N_17662,N_17102);
xnor U18515 (N_18515,N_17365,N_17529);
nand U18516 (N_18516,N_17691,N_17303);
nor U18517 (N_18517,N_17437,N_17082);
or U18518 (N_18518,N_17848,N_17720);
and U18519 (N_18519,N_17686,N_17210);
and U18520 (N_18520,N_17465,N_17599);
or U18521 (N_18521,N_17702,N_17376);
xnor U18522 (N_18522,N_17003,N_17429);
nand U18523 (N_18523,N_17459,N_17283);
and U18524 (N_18524,N_17601,N_17339);
and U18525 (N_18525,N_17387,N_17653);
or U18526 (N_18526,N_17043,N_17209);
nand U18527 (N_18527,N_17213,N_17566);
xnor U18528 (N_18528,N_17925,N_17864);
nor U18529 (N_18529,N_17906,N_17493);
and U18530 (N_18530,N_17619,N_17811);
nor U18531 (N_18531,N_17877,N_17807);
nor U18532 (N_18532,N_17539,N_17295);
and U18533 (N_18533,N_17312,N_17600);
nand U18534 (N_18534,N_17968,N_17674);
nor U18535 (N_18535,N_17060,N_17244);
xor U18536 (N_18536,N_17059,N_17074);
xor U18537 (N_18537,N_17383,N_17161);
nor U18538 (N_18538,N_17157,N_17840);
xor U18539 (N_18539,N_17672,N_17517);
and U18540 (N_18540,N_17246,N_17075);
nand U18541 (N_18541,N_17941,N_17072);
nand U18542 (N_18542,N_17375,N_17403);
or U18543 (N_18543,N_17032,N_17483);
nand U18544 (N_18544,N_17426,N_17418);
or U18545 (N_18545,N_17901,N_17530);
xnor U18546 (N_18546,N_17157,N_17855);
or U18547 (N_18547,N_17667,N_17067);
or U18548 (N_18548,N_17050,N_17029);
xor U18549 (N_18549,N_17766,N_17666);
nand U18550 (N_18550,N_17145,N_17390);
xor U18551 (N_18551,N_17592,N_17836);
nor U18552 (N_18552,N_17352,N_17805);
or U18553 (N_18553,N_17432,N_17633);
nor U18554 (N_18554,N_17714,N_17001);
or U18555 (N_18555,N_17955,N_17820);
nor U18556 (N_18556,N_17351,N_17522);
xor U18557 (N_18557,N_17530,N_17698);
nand U18558 (N_18558,N_17361,N_17387);
nor U18559 (N_18559,N_17165,N_17884);
nand U18560 (N_18560,N_17732,N_17993);
xor U18561 (N_18561,N_17626,N_17375);
and U18562 (N_18562,N_17467,N_17204);
xnor U18563 (N_18563,N_17410,N_17221);
nor U18564 (N_18564,N_17818,N_17527);
or U18565 (N_18565,N_17944,N_17079);
nor U18566 (N_18566,N_17224,N_17062);
xor U18567 (N_18567,N_17880,N_17252);
and U18568 (N_18568,N_17811,N_17599);
xor U18569 (N_18569,N_17352,N_17882);
xor U18570 (N_18570,N_17855,N_17404);
or U18571 (N_18571,N_17093,N_17777);
and U18572 (N_18572,N_17380,N_17556);
nor U18573 (N_18573,N_17902,N_17146);
xor U18574 (N_18574,N_17108,N_17554);
xor U18575 (N_18575,N_17080,N_17306);
nor U18576 (N_18576,N_17986,N_17707);
nand U18577 (N_18577,N_17417,N_17049);
nor U18578 (N_18578,N_17781,N_17667);
nor U18579 (N_18579,N_17938,N_17540);
and U18580 (N_18580,N_17212,N_17816);
nor U18581 (N_18581,N_17220,N_17067);
xnor U18582 (N_18582,N_17896,N_17911);
and U18583 (N_18583,N_17357,N_17350);
xnor U18584 (N_18584,N_17430,N_17491);
nand U18585 (N_18585,N_17475,N_17574);
or U18586 (N_18586,N_17837,N_17349);
nor U18587 (N_18587,N_17009,N_17200);
nor U18588 (N_18588,N_17336,N_17153);
nor U18589 (N_18589,N_17152,N_17570);
or U18590 (N_18590,N_17421,N_17003);
and U18591 (N_18591,N_17811,N_17550);
and U18592 (N_18592,N_17176,N_17746);
nor U18593 (N_18593,N_17137,N_17714);
and U18594 (N_18594,N_17288,N_17472);
or U18595 (N_18595,N_17410,N_17642);
nand U18596 (N_18596,N_17183,N_17821);
nor U18597 (N_18597,N_17915,N_17117);
nor U18598 (N_18598,N_17653,N_17203);
and U18599 (N_18599,N_17413,N_17830);
or U18600 (N_18600,N_17415,N_17370);
or U18601 (N_18601,N_17590,N_17281);
xnor U18602 (N_18602,N_17907,N_17433);
nand U18603 (N_18603,N_17680,N_17362);
nand U18604 (N_18604,N_17699,N_17636);
xnor U18605 (N_18605,N_17541,N_17255);
nand U18606 (N_18606,N_17655,N_17340);
and U18607 (N_18607,N_17209,N_17369);
nor U18608 (N_18608,N_17800,N_17578);
nor U18609 (N_18609,N_17742,N_17752);
and U18610 (N_18610,N_17696,N_17145);
or U18611 (N_18611,N_17575,N_17346);
xnor U18612 (N_18612,N_17420,N_17796);
and U18613 (N_18613,N_17228,N_17379);
nand U18614 (N_18614,N_17803,N_17303);
xnor U18615 (N_18615,N_17672,N_17336);
xor U18616 (N_18616,N_17707,N_17047);
xor U18617 (N_18617,N_17319,N_17439);
nand U18618 (N_18618,N_17375,N_17145);
nand U18619 (N_18619,N_17987,N_17249);
and U18620 (N_18620,N_17496,N_17655);
or U18621 (N_18621,N_17032,N_17637);
and U18622 (N_18622,N_17712,N_17678);
and U18623 (N_18623,N_17245,N_17183);
xor U18624 (N_18624,N_17403,N_17007);
and U18625 (N_18625,N_17513,N_17827);
nor U18626 (N_18626,N_17963,N_17473);
nand U18627 (N_18627,N_17579,N_17548);
or U18628 (N_18628,N_17062,N_17342);
xor U18629 (N_18629,N_17857,N_17822);
or U18630 (N_18630,N_17059,N_17922);
xnor U18631 (N_18631,N_17567,N_17322);
or U18632 (N_18632,N_17326,N_17107);
or U18633 (N_18633,N_17819,N_17927);
xnor U18634 (N_18634,N_17274,N_17884);
xnor U18635 (N_18635,N_17671,N_17643);
xnor U18636 (N_18636,N_17451,N_17706);
nor U18637 (N_18637,N_17410,N_17929);
and U18638 (N_18638,N_17859,N_17547);
nand U18639 (N_18639,N_17697,N_17200);
xor U18640 (N_18640,N_17809,N_17159);
nand U18641 (N_18641,N_17178,N_17900);
nand U18642 (N_18642,N_17789,N_17238);
xnor U18643 (N_18643,N_17371,N_17830);
or U18644 (N_18644,N_17343,N_17058);
or U18645 (N_18645,N_17013,N_17959);
and U18646 (N_18646,N_17486,N_17818);
and U18647 (N_18647,N_17507,N_17096);
and U18648 (N_18648,N_17870,N_17422);
or U18649 (N_18649,N_17898,N_17691);
nand U18650 (N_18650,N_17473,N_17200);
nand U18651 (N_18651,N_17100,N_17736);
xor U18652 (N_18652,N_17773,N_17967);
or U18653 (N_18653,N_17186,N_17247);
xor U18654 (N_18654,N_17768,N_17003);
or U18655 (N_18655,N_17965,N_17493);
nand U18656 (N_18656,N_17173,N_17360);
nand U18657 (N_18657,N_17988,N_17678);
xor U18658 (N_18658,N_17836,N_17317);
nor U18659 (N_18659,N_17552,N_17066);
nor U18660 (N_18660,N_17645,N_17098);
xor U18661 (N_18661,N_17949,N_17693);
and U18662 (N_18662,N_17097,N_17086);
xor U18663 (N_18663,N_17809,N_17787);
nor U18664 (N_18664,N_17867,N_17863);
nor U18665 (N_18665,N_17566,N_17512);
and U18666 (N_18666,N_17612,N_17599);
nor U18667 (N_18667,N_17582,N_17885);
and U18668 (N_18668,N_17634,N_17407);
nand U18669 (N_18669,N_17245,N_17001);
nor U18670 (N_18670,N_17791,N_17198);
nand U18671 (N_18671,N_17566,N_17507);
nand U18672 (N_18672,N_17115,N_17870);
or U18673 (N_18673,N_17861,N_17965);
nand U18674 (N_18674,N_17935,N_17112);
or U18675 (N_18675,N_17006,N_17803);
or U18676 (N_18676,N_17996,N_17136);
and U18677 (N_18677,N_17606,N_17400);
xnor U18678 (N_18678,N_17460,N_17782);
nand U18679 (N_18679,N_17202,N_17696);
xnor U18680 (N_18680,N_17618,N_17975);
nor U18681 (N_18681,N_17498,N_17349);
or U18682 (N_18682,N_17984,N_17008);
nor U18683 (N_18683,N_17758,N_17665);
or U18684 (N_18684,N_17652,N_17081);
nor U18685 (N_18685,N_17143,N_17938);
nor U18686 (N_18686,N_17047,N_17494);
and U18687 (N_18687,N_17839,N_17094);
and U18688 (N_18688,N_17696,N_17836);
nand U18689 (N_18689,N_17756,N_17114);
or U18690 (N_18690,N_17709,N_17079);
nand U18691 (N_18691,N_17601,N_17624);
and U18692 (N_18692,N_17060,N_17231);
or U18693 (N_18693,N_17833,N_17794);
xor U18694 (N_18694,N_17250,N_17886);
xor U18695 (N_18695,N_17528,N_17211);
nand U18696 (N_18696,N_17508,N_17960);
and U18697 (N_18697,N_17216,N_17895);
nand U18698 (N_18698,N_17802,N_17476);
and U18699 (N_18699,N_17671,N_17240);
and U18700 (N_18700,N_17951,N_17977);
nor U18701 (N_18701,N_17073,N_17188);
nand U18702 (N_18702,N_17744,N_17705);
xor U18703 (N_18703,N_17453,N_17568);
nand U18704 (N_18704,N_17280,N_17935);
nor U18705 (N_18705,N_17705,N_17417);
xor U18706 (N_18706,N_17066,N_17614);
and U18707 (N_18707,N_17038,N_17640);
and U18708 (N_18708,N_17500,N_17405);
and U18709 (N_18709,N_17216,N_17989);
xnor U18710 (N_18710,N_17588,N_17608);
or U18711 (N_18711,N_17064,N_17213);
or U18712 (N_18712,N_17097,N_17337);
or U18713 (N_18713,N_17226,N_17084);
and U18714 (N_18714,N_17040,N_17120);
nand U18715 (N_18715,N_17691,N_17191);
nand U18716 (N_18716,N_17935,N_17912);
and U18717 (N_18717,N_17604,N_17879);
or U18718 (N_18718,N_17992,N_17476);
xor U18719 (N_18719,N_17260,N_17612);
or U18720 (N_18720,N_17907,N_17537);
and U18721 (N_18721,N_17576,N_17023);
nor U18722 (N_18722,N_17186,N_17777);
or U18723 (N_18723,N_17138,N_17575);
xor U18724 (N_18724,N_17877,N_17432);
or U18725 (N_18725,N_17204,N_17470);
and U18726 (N_18726,N_17664,N_17998);
nor U18727 (N_18727,N_17166,N_17899);
or U18728 (N_18728,N_17676,N_17941);
and U18729 (N_18729,N_17498,N_17129);
xor U18730 (N_18730,N_17842,N_17205);
xnor U18731 (N_18731,N_17967,N_17091);
and U18732 (N_18732,N_17293,N_17858);
xnor U18733 (N_18733,N_17760,N_17222);
and U18734 (N_18734,N_17932,N_17388);
nand U18735 (N_18735,N_17978,N_17430);
xnor U18736 (N_18736,N_17145,N_17251);
and U18737 (N_18737,N_17786,N_17514);
xor U18738 (N_18738,N_17145,N_17447);
or U18739 (N_18739,N_17514,N_17054);
nor U18740 (N_18740,N_17629,N_17262);
nand U18741 (N_18741,N_17851,N_17681);
and U18742 (N_18742,N_17495,N_17871);
nand U18743 (N_18743,N_17615,N_17933);
and U18744 (N_18744,N_17680,N_17499);
nand U18745 (N_18745,N_17858,N_17504);
nor U18746 (N_18746,N_17148,N_17650);
nor U18747 (N_18747,N_17995,N_17479);
and U18748 (N_18748,N_17717,N_17792);
or U18749 (N_18749,N_17198,N_17456);
nand U18750 (N_18750,N_17888,N_17091);
and U18751 (N_18751,N_17441,N_17024);
nand U18752 (N_18752,N_17286,N_17792);
nand U18753 (N_18753,N_17615,N_17110);
nand U18754 (N_18754,N_17182,N_17727);
nand U18755 (N_18755,N_17871,N_17470);
nand U18756 (N_18756,N_17391,N_17412);
nor U18757 (N_18757,N_17215,N_17329);
nand U18758 (N_18758,N_17511,N_17616);
nor U18759 (N_18759,N_17802,N_17816);
or U18760 (N_18760,N_17585,N_17214);
and U18761 (N_18761,N_17655,N_17475);
nor U18762 (N_18762,N_17376,N_17007);
and U18763 (N_18763,N_17481,N_17307);
nor U18764 (N_18764,N_17114,N_17412);
xnor U18765 (N_18765,N_17904,N_17470);
or U18766 (N_18766,N_17492,N_17183);
nor U18767 (N_18767,N_17981,N_17523);
and U18768 (N_18768,N_17358,N_17223);
or U18769 (N_18769,N_17388,N_17063);
nor U18770 (N_18770,N_17229,N_17906);
nand U18771 (N_18771,N_17583,N_17645);
or U18772 (N_18772,N_17502,N_17304);
nor U18773 (N_18773,N_17067,N_17452);
xor U18774 (N_18774,N_17912,N_17813);
nand U18775 (N_18775,N_17805,N_17986);
nor U18776 (N_18776,N_17838,N_17878);
or U18777 (N_18777,N_17268,N_17803);
nor U18778 (N_18778,N_17277,N_17156);
and U18779 (N_18779,N_17641,N_17626);
xnor U18780 (N_18780,N_17778,N_17716);
nand U18781 (N_18781,N_17658,N_17263);
nor U18782 (N_18782,N_17329,N_17680);
xor U18783 (N_18783,N_17647,N_17907);
xor U18784 (N_18784,N_17824,N_17530);
xor U18785 (N_18785,N_17062,N_17866);
nor U18786 (N_18786,N_17246,N_17751);
and U18787 (N_18787,N_17910,N_17975);
nand U18788 (N_18788,N_17074,N_17105);
and U18789 (N_18789,N_17425,N_17062);
nand U18790 (N_18790,N_17340,N_17527);
or U18791 (N_18791,N_17414,N_17577);
nor U18792 (N_18792,N_17564,N_17960);
nor U18793 (N_18793,N_17791,N_17013);
and U18794 (N_18794,N_17379,N_17186);
xnor U18795 (N_18795,N_17875,N_17451);
or U18796 (N_18796,N_17222,N_17566);
nor U18797 (N_18797,N_17303,N_17992);
nand U18798 (N_18798,N_17654,N_17839);
or U18799 (N_18799,N_17499,N_17390);
nor U18800 (N_18800,N_17456,N_17339);
nor U18801 (N_18801,N_17095,N_17512);
or U18802 (N_18802,N_17923,N_17544);
nand U18803 (N_18803,N_17688,N_17454);
and U18804 (N_18804,N_17814,N_17995);
and U18805 (N_18805,N_17038,N_17246);
or U18806 (N_18806,N_17222,N_17214);
nor U18807 (N_18807,N_17331,N_17132);
xnor U18808 (N_18808,N_17601,N_17701);
or U18809 (N_18809,N_17643,N_17905);
nand U18810 (N_18810,N_17353,N_17805);
or U18811 (N_18811,N_17244,N_17376);
or U18812 (N_18812,N_17682,N_17652);
or U18813 (N_18813,N_17672,N_17174);
and U18814 (N_18814,N_17324,N_17481);
or U18815 (N_18815,N_17863,N_17659);
or U18816 (N_18816,N_17070,N_17435);
xnor U18817 (N_18817,N_17135,N_17213);
nor U18818 (N_18818,N_17422,N_17998);
nor U18819 (N_18819,N_17984,N_17726);
or U18820 (N_18820,N_17408,N_17062);
xor U18821 (N_18821,N_17440,N_17055);
nand U18822 (N_18822,N_17572,N_17288);
or U18823 (N_18823,N_17649,N_17686);
nor U18824 (N_18824,N_17258,N_17183);
nand U18825 (N_18825,N_17176,N_17029);
or U18826 (N_18826,N_17083,N_17300);
or U18827 (N_18827,N_17739,N_17272);
nor U18828 (N_18828,N_17309,N_17770);
nand U18829 (N_18829,N_17361,N_17616);
and U18830 (N_18830,N_17269,N_17585);
and U18831 (N_18831,N_17501,N_17265);
nand U18832 (N_18832,N_17551,N_17912);
and U18833 (N_18833,N_17981,N_17348);
or U18834 (N_18834,N_17162,N_17231);
nand U18835 (N_18835,N_17101,N_17510);
and U18836 (N_18836,N_17731,N_17998);
or U18837 (N_18837,N_17576,N_17938);
and U18838 (N_18838,N_17822,N_17806);
or U18839 (N_18839,N_17859,N_17731);
or U18840 (N_18840,N_17805,N_17062);
nand U18841 (N_18841,N_17566,N_17335);
nand U18842 (N_18842,N_17918,N_17922);
or U18843 (N_18843,N_17440,N_17094);
or U18844 (N_18844,N_17930,N_17536);
xnor U18845 (N_18845,N_17773,N_17597);
or U18846 (N_18846,N_17760,N_17752);
or U18847 (N_18847,N_17544,N_17587);
or U18848 (N_18848,N_17659,N_17083);
and U18849 (N_18849,N_17839,N_17437);
xor U18850 (N_18850,N_17989,N_17345);
xor U18851 (N_18851,N_17984,N_17167);
xnor U18852 (N_18852,N_17956,N_17249);
xor U18853 (N_18853,N_17262,N_17993);
xnor U18854 (N_18854,N_17806,N_17938);
or U18855 (N_18855,N_17611,N_17416);
or U18856 (N_18856,N_17012,N_17437);
xor U18857 (N_18857,N_17218,N_17507);
or U18858 (N_18858,N_17186,N_17609);
xnor U18859 (N_18859,N_17729,N_17533);
nand U18860 (N_18860,N_17156,N_17887);
nor U18861 (N_18861,N_17565,N_17998);
xor U18862 (N_18862,N_17780,N_17696);
and U18863 (N_18863,N_17156,N_17933);
or U18864 (N_18864,N_17677,N_17112);
or U18865 (N_18865,N_17099,N_17561);
xor U18866 (N_18866,N_17023,N_17050);
nand U18867 (N_18867,N_17410,N_17524);
xnor U18868 (N_18868,N_17371,N_17472);
or U18869 (N_18869,N_17502,N_17813);
nor U18870 (N_18870,N_17400,N_17069);
and U18871 (N_18871,N_17714,N_17326);
or U18872 (N_18872,N_17837,N_17697);
xnor U18873 (N_18873,N_17982,N_17385);
nand U18874 (N_18874,N_17904,N_17870);
nor U18875 (N_18875,N_17313,N_17931);
xor U18876 (N_18876,N_17539,N_17155);
or U18877 (N_18877,N_17414,N_17228);
nor U18878 (N_18878,N_17232,N_17595);
or U18879 (N_18879,N_17925,N_17343);
nand U18880 (N_18880,N_17536,N_17415);
xnor U18881 (N_18881,N_17509,N_17911);
nand U18882 (N_18882,N_17071,N_17229);
xor U18883 (N_18883,N_17243,N_17267);
nor U18884 (N_18884,N_17412,N_17431);
xor U18885 (N_18885,N_17946,N_17520);
nor U18886 (N_18886,N_17636,N_17852);
nor U18887 (N_18887,N_17718,N_17607);
nand U18888 (N_18888,N_17175,N_17937);
or U18889 (N_18889,N_17647,N_17319);
nor U18890 (N_18890,N_17484,N_17901);
nor U18891 (N_18891,N_17965,N_17257);
and U18892 (N_18892,N_17855,N_17471);
xnor U18893 (N_18893,N_17589,N_17875);
nand U18894 (N_18894,N_17150,N_17250);
or U18895 (N_18895,N_17311,N_17504);
or U18896 (N_18896,N_17978,N_17846);
or U18897 (N_18897,N_17384,N_17527);
xnor U18898 (N_18898,N_17144,N_17757);
nor U18899 (N_18899,N_17031,N_17746);
and U18900 (N_18900,N_17116,N_17383);
or U18901 (N_18901,N_17428,N_17932);
nor U18902 (N_18902,N_17400,N_17407);
and U18903 (N_18903,N_17096,N_17465);
nor U18904 (N_18904,N_17197,N_17977);
xnor U18905 (N_18905,N_17913,N_17053);
nand U18906 (N_18906,N_17654,N_17092);
nor U18907 (N_18907,N_17391,N_17379);
nand U18908 (N_18908,N_17594,N_17946);
or U18909 (N_18909,N_17980,N_17070);
nor U18910 (N_18910,N_17386,N_17874);
xor U18911 (N_18911,N_17455,N_17539);
xnor U18912 (N_18912,N_17365,N_17071);
and U18913 (N_18913,N_17063,N_17704);
and U18914 (N_18914,N_17476,N_17506);
nand U18915 (N_18915,N_17959,N_17335);
nand U18916 (N_18916,N_17007,N_17742);
and U18917 (N_18917,N_17588,N_17180);
xor U18918 (N_18918,N_17652,N_17797);
or U18919 (N_18919,N_17264,N_17445);
and U18920 (N_18920,N_17666,N_17661);
and U18921 (N_18921,N_17071,N_17454);
and U18922 (N_18922,N_17558,N_17195);
nand U18923 (N_18923,N_17541,N_17543);
nand U18924 (N_18924,N_17694,N_17718);
nand U18925 (N_18925,N_17523,N_17440);
nand U18926 (N_18926,N_17524,N_17430);
nand U18927 (N_18927,N_17048,N_17128);
nand U18928 (N_18928,N_17612,N_17115);
or U18929 (N_18929,N_17014,N_17416);
xor U18930 (N_18930,N_17925,N_17736);
nand U18931 (N_18931,N_17413,N_17402);
nor U18932 (N_18932,N_17849,N_17161);
nor U18933 (N_18933,N_17706,N_17201);
nand U18934 (N_18934,N_17280,N_17978);
xnor U18935 (N_18935,N_17224,N_17894);
or U18936 (N_18936,N_17004,N_17798);
xnor U18937 (N_18937,N_17288,N_17505);
or U18938 (N_18938,N_17231,N_17490);
or U18939 (N_18939,N_17789,N_17957);
nand U18940 (N_18940,N_17275,N_17293);
nand U18941 (N_18941,N_17342,N_17740);
or U18942 (N_18942,N_17915,N_17061);
or U18943 (N_18943,N_17476,N_17882);
and U18944 (N_18944,N_17475,N_17862);
xor U18945 (N_18945,N_17132,N_17546);
nor U18946 (N_18946,N_17625,N_17004);
xnor U18947 (N_18947,N_17717,N_17261);
xor U18948 (N_18948,N_17662,N_17956);
xnor U18949 (N_18949,N_17505,N_17346);
nand U18950 (N_18950,N_17286,N_17018);
or U18951 (N_18951,N_17316,N_17483);
nor U18952 (N_18952,N_17624,N_17028);
nand U18953 (N_18953,N_17563,N_17088);
nor U18954 (N_18954,N_17187,N_17424);
or U18955 (N_18955,N_17218,N_17968);
nand U18956 (N_18956,N_17486,N_17719);
nor U18957 (N_18957,N_17631,N_17166);
nor U18958 (N_18958,N_17750,N_17520);
nor U18959 (N_18959,N_17401,N_17405);
nand U18960 (N_18960,N_17236,N_17889);
and U18961 (N_18961,N_17159,N_17513);
or U18962 (N_18962,N_17887,N_17220);
or U18963 (N_18963,N_17871,N_17103);
xnor U18964 (N_18964,N_17939,N_17501);
xnor U18965 (N_18965,N_17765,N_17007);
or U18966 (N_18966,N_17783,N_17387);
or U18967 (N_18967,N_17498,N_17608);
nand U18968 (N_18968,N_17299,N_17616);
and U18969 (N_18969,N_17714,N_17595);
and U18970 (N_18970,N_17773,N_17218);
or U18971 (N_18971,N_17558,N_17089);
xnor U18972 (N_18972,N_17667,N_17884);
xnor U18973 (N_18973,N_17511,N_17223);
nand U18974 (N_18974,N_17935,N_17410);
nor U18975 (N_18975,N_17122,N_17449);
xor U18976 (N_18976,N_17329,N_17088);
or U18977 (N_18977,N_17743,N_17321);
and U18978 (N_18978,N_17661,N_17873);
nor U18979 (N_18979,N_17810,N_17212);
and U18980 (N_18980,N_17407,N_17726);
xor U18981 (N_18981,N_17367,N_17836);
nor U18982 (N_18982,N_17187,N_17396);
or U18983 (N_18983,N_17586,N_17355);
xor U18984 (N_18984,N_17161,N_17535);
or U18985 (N_18985,N_17811,N_17754);
or U18986 (N_18986,N_17909,N_17787);
nand U18987 (N_18987,N_17452,N_17999);
or U18988 (N_18988,N_17048,N_17878);
nand U18989 (N_18989,N_17810,N_17186);
and U18990 (N_18990,N_17782,N_17528);
nor U18991 (N_18991,N_17655,N_17380);
nand U18992 (N_18992,N_17523,N_17127);
and U18993 (N_18993,N_17894,N_17210);
xor U18994 (N_18994,N_17028,N_17452);
or U18995 (N_18995,N_17824,N_17243);
and U18996 (N_18996,N_17299,N_17271);
xor U18997 (N_18997,N_17089,N_17680);
nor U18998 (N_18998,N_17526,N_17561);
xor U18999 (N_18999,N_17431,N_17063);
nand U19000 (N_19000,N_18497,N_18749);
nor U19001 (N_19001,N_18371,N_18234);
and U19002 (N_19002,N_18925,N_18215);
and U19003 (N_19003,N_18722,N_18014);
or U19004 (N_19004,N_18112,N_18980);
nor U19005 (N_19005,N_18937,N_18914);
xor U19006 (N_19006,N_18872,N_18956);
and U19007 (N_19007,N_18150,N_18985);
and U19008 (N_19008,N_18965,N_18794);
and U19009 (N_19009,N_18069,N_18002);
xnor U19010 (N_19010,N_18630,N_18131);
nand U19011 (N_19011,N_18140,N_18336);
nand U19012 (N_19012,N_18922,N_18694);
or U19013 (N_19013,N_18175,N_18827);
nand U19014 (N_19014,N_18300,N_18455);
nand U19015 (N_19015,N_18538,N_18718);
or U19016 (N_19016,N_18037,N_18634);
xnor U19017 (N_19017,N_18829,N_18225);
or U19018 (N_19018,N_18022,N_18944);
nor U19019 (N_19019,N_18546,N_18589);
nand U19020 (N_19020,N_18159,N_18576);
nor U19021 (N_19021,N_18989,N_18657);
xnor U19022 (N_19022,N_18009,N_18063);
or U19023 (N_19023,N_18342,N_18543);
nor U19024 (N_19024,N_18427,N_18788);
nand U19025 (N_19025,N_18616,N_18291);
and U19026 (N_19026,N_18795,N_18001);
and U19027 (N_19027,N_18849,N_18417);
xnor U19028 (N_19028,N_18747,N_18835);
nor U19029 (N_19029,N_18414,N_18281);
nand U19030 (N_19030,N_18452,N_18902);
or U19031 (N_19031,N_18545,N_18519);
nand U19032 (N_19032,N_18400,N_18017);
and U19033 (N_19033,N_18242,N_18282);
nor U19034 (N_19034,N_18750,N_18223);
nand U19035 (N_19035,N_18510,N_18122);
or U19036 (N_19036,N_18712,N_18928);
nand U19037 (N_19037,N_18704,N_18803);
and U19038 (N_19038,N_18841,N_18528);
nand U19039 (N_19039,N_18777,N_18806);
xnor U19040 (N_19040,N_18461,N_18283);
nand U19041 (N_19041,N_18118,N_18278);
nor U19042 (N_19042,N_18953,N_18789);
nor U19043 (N_19043,N_18114,N_18912);
nand U19044 (N_19044,N_18854,N_18391);
xor U19045 (N_19045,N_18491,N_18678);
or U19046 (N_19046,N_18115,N_18309);
nor U19047 (N_19047,N_18144,N_18516);
xnor U19048 (N_19048,N_18015,N_18277);
or U19049 (N_19049,N_18745,N_18493);
nor U19050 (N_19050,N_18412,N_18683);
nand U19051 (N_19051,N_18020,N_18554);
xnor U19052 (N_19052,N_18329,N_18428);
nor U19053 (N_19053,N_18553,N_18601);
xor U19054 (N_19054,N_18062,N_18705);
nand U19055 (N_19055,N_18091,N_18586);
and U19056 (N_19056,N_18809,N_18116);
nor U19057 (N_19057,N_18056,N_18351);
nand U19058 (N_19058,N_18076,N_18097);
nor U19059 (N_19059,N_18879,N_18170);
nand U19060 (N_19060,N_18093,N_18903);
and U19061 (N_19061,N_18184,N_18326);
xor U19062 (N_19062,N_18172,N_18158);
or U19063 (N_19063,N_18167,N_18785);
nor U19064 (N_19064,N_18374,N_18688);
nand U19065 (N_19065,N_18540,N_18203);
and U19066 (N_19066,N_18018,N_18901);
nand U19067 (N_19067,N_18092,N_18462);
and U19068 (N_19068,N_18531,N_18924);
xor U19069 (N_19069,N_18617,N_18730);
or U19070 (N_19070,N_18422,N_18627);
xor U19071 (N_19071,N_18869,N_18366);
or U19072 (N_19072,N_18032,N_18075);
or U19073 (N_19073,N_18010,N_18209);
nor U19074 (N_19074,N_18890,N_18372);
nor U19075 (N_19075,N_18344,N_18232);
and U19076 (N_19076,N_18824,N_18111);
xnor U19077 (N_19077,N_18771,N_18684);
or U19078 (N_19078,N_18489,N_18844);
xor U19079 (N_19079,N_18068,N_18306);
nor U19080 (N_19080,N_18386,N_18620);
nand U19081 (N_19081,N_18907,N_18904);
xor U19082 (N_19082,N_18911,N_18316);
or U19083 (N_19083,N_18915,N_18072);
nor U19084 (N_19084,N_18436,N_18481);
nand U19085 (N_19085,N_18270,N_18542);
and U19086 (N_19086,N_18347,N_18446);
and U19087 (N_19087,N_18036,N_18752);
or U19088 (N_19088,N_18379,N_18966);
and U19089 (N_19089,N_18739,N_18641);
or U19090 (N_19090,N_18280,N_18467);
or U19091 (N_19091,N_18125,N_18363);
xnor U19092 (N_19092,N_18243,N_18143);
or U19093 (N_19093,N_18858,N_18130);
nand U19094 (N_19094,N_18043,N_18057);
or U19095 (N_19095,N_18052,N_18120);
nand U19096 (N_19096,N_18958,N_18050);
and U19097 (N_19097,N_18011,N_18706);
xnor U19098 (N_19098,N_18590,N_18474);
xor U19099 (N_19099,N_18898,N_18439);
or U19100 (N_19100,N_18210,N_18786);
nor U19101 (N_19101,N_18049,N_18679);
nand U19102 (N_19102,N_18707,N_18247);
nand U19103 (N_19103,N_18108,N_18725);
nor U19104 (N_19104,N_18358,N_18578);
nand U19105 (N_19105,N_18318,N_18146);
nor U19106 (N_19106,N_18486,N_18656);
nand U19107 (N_19107,N_18579,N_18463);
nor U19108 (N_19108,N_18887,N_18921);
xnor U19109 (N_19109,N_18698,N_18814);
nor U19110 (N_19110,N_18023,N_18896);
xor U19111 (N_19111,N_18064,N_18437);
or U19112 (N_19112,N_18830,N_18638);
and U19113 (N_19113,N_18867,N_18550);
and U19114 (N_19114,N_18834,N_18016);
nand U19115 (N_19115,N_18163,N_18496);
nor U19116 (N_19116,N_18339,N_18755);
or U19117 (N_19117,N_18449,N_18791);
and U19118 (N_19118,N_18645,N_18080);
xnor U19119 (N_19119,N_18539,N_18293);
xnor U19120 (N_19120,N_18848,N_18709);
nor U19121 (N_19121,N_18717,N_18744);
or U19122 (N_19122,N_18521,N_18605);
or U19123 (N_19123,N_18065,N_18674);
nor U19124 (N_19124,N_18876,N_18810);
or U19125 (N_19125,N_18622,N_18990);
nor U19126 (N_19126,N_18328,N_18945);
nand U19127 (N_19127,N_18799,N_18479);
xor U19128 (N_19128,N_18419,N_18581);
and U19129 (N_19129,N_18040,N_18792);
nand U19130 (N_19130,N_18136,N_18297);
xor U19131 (N_19131,N_18027,N_18310);
nor U19132 (N_19132,N_18758,N_18769);
xor U19133 (N_19133,N_18007,N_18754);
nand U19134 (N_19134,N_18950,N_18629);
nand U19135 (N_19135,N_18506,N_18190);
or U19136 (N_19136,N_18976,N_18729);
and U19137 (N_19137,N_18975,N_18171);
and U19138 (N_19138,N_18411,N_18337);
nand U19139 (N_19139,N_18299,N_18793);
nor U19140 (N_19140,N_18893,N_18853);
and U19141 (N_19141,N_18839,N_18689);
and U19142 (N_19142,N_18986,N_18024);
xor U19143 (N_19143,N_18659,N_18728);
xnor U19144 (N_19144,N_18384,N_18039);
or U19145 (N_19145,N_18443,N_18383);
nor U19146 (N_19146,N_18626,N_18089);
nand U19147 (N_19147,N_18602,N_18485);
or U19148 (N_19148,N_18646,N_18191);
or U19149 (N_19149,N_18587,N_18285);
or U19150 (N_19150,N_18327,N_18444);
nor U19151 (N_19151,N_18085,N_18425);
xor U19152 (N_19152,N_18984,N_18088);
and U19153 (N_19153,N_18940,N_18547);
nor U19154 (N_19154,N_18095,N_18987);
or U19155 (N_19155,N_18483,N_18889);
nand U19156 (N_19156,N_18644,N_18536);
xor U19157 (N_19157,N_18996,N_18224);
nand U19158 (N_19158,N_18708,N_18251);
nand U19159 (N_19159,N_18840,N_18783);
nor U19160 (N_19160,N_18660,N_18606);
xnor U19161 (N_19161,N_18238,N_18073);
and U19162 (N_19162,N_18222,N_18556);
and U19163 (N_19163,N_18932,N_18129);
or U19164 (N_19164,N_18857,N_18995);
xor U19165 (N_19165,N_18077,N_18677);
or U19166 (N_19166,N_18193,N_18256);
nor U19167 (N_19167,N_18811,N_18561);
or U19168 (N_19168,N_18367,N_18687);
xnor U19169 (N_19169,N_18059,N_18421);
nor U19170 (N_19170,N_18974,N_18655);
and U19171 (N_19171,N_18305,N_18868);
nand U19172 (N_19172,N_18906,N_18713);
or U19173 (N_19173,N_18537,N_18782);
or U19174 (N_19174,N_18200,N_18279);
nor U19175 (N_19175,N_18983,N_18774);
nor U19176 (N_19176,N_18658,N_18476);
and U19177 (N_19177,N_18507,N_18664);
and U19178 (N_19178,N_18760,N_18250);
nand U19179 (N_19179,N_18004,N_18322);
xor U19180 (N_19180,N_18737,N_18424);
nor U19181 (N_19181,N_18920,N_18923);
nand U19182 (N_19182,N_18308,N_18571);
or U19183 (N_19183,N_18354,N_18335);
nand U19184 (N_19184,N_18740,N_18632);
nor U19185 (N_19185,N_18820,N_18319);
xor U19186 (N_19186,N_18165,N_18153);
and U19187 (N_19187,N_18731,N_18535);
nand U19188 (N_19188,N_18727,N_18797);
or U19189 (N_19189,N_18380,N_18465);
nor U19190 (N_19190,N_18185,N_18218);
nand U19191 (N_19191,N_18784,N_18426);
nor U19192 (N_19192,N_18971,N_18487);
or U19193 (N_19193,N_18382,N_18375);
xor U19194 (N_19194,N_18913,N_18231);
xor U19195 (N_19195,N_18584,N_18842);
and U19196 (N_19196,N_18287,N_18407);
and U19197 (N_19197,N_18173,N_18388);
and U19198 (N_19198,N_18138,N_18880);
nand U19199 (N_19199,N_18307,N_18033);
and U19200 (N_19200,N_18636,N_18292);
nand U19201 (N_19201,N_18988,N_18441);
xnor U19202 (N_19202,N_18826,N_18034);
nand U19203 (N_19203,N_18759,N_18899);
or U19204 (N_19204,N_18315,N_18060);
and U19205 (N_19205,N_18770,N_18891);
and U19206 (N_19206,N_18523,N_18081);
nor U19207 (N_19207,N_18580,N_18952);
nor U19208 (N_19208,N_18653,N_18696);
or U19209 (N_19209,N_18863,N_18522);
xor U19210 (N_19210,N_18509,N_18503);
or U19211 (N_19211,N_18333,N_18457);
or U19212 (N_19212,N_18527,N_18753);
xnor U19213 (N_19213,N_18931,N_18262);
nand U19214 (N_19214,N_18877,N_18239);
nand U19215 (N_19215,N_18765,N_18711);
or U19216 (N_19216,N_18313,N_18202);
xor U19217 (N_19217,N_18330,N_18451);
xor U19218 (N_19218,N_18030,N_18403);
xnor U19219 (N_19219,N_18460,N_18997);
nor U19220 (N_19220,N_18357,N_18942);
nor U19221 (N_19221,N_18169,N_18423);
nor U19222 (N_19222,N_18926,N_18265);
xor U19223 (N_19223,N_18054,N_18373);
and U19224 (N_19224,N_18895,N_18948);
nor U19225 (N_19225,N_18733,N_18667);
or U19226 (N_19226,N_18723,N_18847);
nor U19227 (N_19227,N_18643,N_18416);
nand U19228 (N_19228,N_18756,N_18668);
nand U19229 (N_19229,N_18591,N_18544);
and U19230 (N_19230,N_18512,N_18045);
or U19231 (N_19231,N_18133,N_18669);
xnor U19232 (N_19232,N_18494,N_18048);
and U19233 (N_19233,N_18625,N_18181);
nand U19234 (N_19234,N_18078,N_18802);
and U19235 (N_19235,N_18177,N_18220);
or U19236 (N_19236,N_18410,N_18724);
nor U19237 (N_19237,N_18776,N_18343);
and U19238 (N_19238,N_18775,N_18480);
nand U19239 (N_19239,N_18505,N_18919);
nand U19240 (N_19240,N_18067,N_18324);
nor U19241 (N_19241,N_18355,N_18969);
nor U19242 (N_19242,N_18404,N_18126);
nor U19243 (N_19243,N_18087,N_18517);
xor U19244 (N_19244,N_18502,N_18151);
and U19245 (N_19245,N_18205,N_18935);
and U19246 (N_19246,N_18458,N_18703);
or U19247 (N_19247,N_18599,N_18495);
nand U19248 (N_19248,N_18716,N_18453);
xor U19249 (N_19249,N_18104,N_18398);
nor U19250 (N_19250,N_18066,N_18246);
nor U19251 (N_19251,N_18180,N_18325);
or U19252 (N_19252,N_18098,N_18888);
and U19253 (N_19253,N_18992,N_18003);
and U19254 (N_19254,N_18930,N_18255);
nor U19255 (N_19255,N_18000,N_18501);
nor U19256 (N_19256,N_18055,N_18160);
and U19257 (N_19257,N_18511,N_18764);
nand U19258 (N_19258,N_18141,N_18838);
nor U19259 (N_19259,N_18233,N_18440);
nand U19260 (N_19260,N_18697,N_18572);
nand U19261 (N_19261,N_18035,N_18148);
or U19262 (N_19262,N_18188,N_18096);
xor U19263 (N_19263,N_18102,N_18821);
xnor U19264 (N_19264,N_18947,N_18038);
or U19265 (N_19265,N_18442,N_18843);
or U19266 (N_19266,N_18135,N_18107);
or U19267 (N_19267,N_18909,N_18019);
nor U19268 (N_19268,N_18401,N_18473);
and U19269 (N_19269,N_18804,N_18615);
xnor U19270 (N_19270,N_18365,N_18435);
and U19271 (N_19271,N_18621,N_18445);
and U19272 (N_19272,N_18456,N_18204);
nand U19273 (N_19273,N_18682,N_18772);
xnor U19274 (N_19274,N_18533,N_18008);
nand U19275 (N_19275,N_18851,N_18781);
and U19276 (N_19276,N_18676,N_18377);
and U19277 (N_19277,N_18855,N_18530);
or U19278 (N_19278,N_18700,N_18999);
xnor U19279 (N_19279,N_18936,N_18642);
nand U19280 (N_19280,N_18680,N_18106);
nor U19281 (N_19281,N_18807,N_18113);
nand U19282 (N_19282,N_18047,N_18822);
xor U19283 (N_19283,N_18885,N_18800);
nand U19284 (N_19284,N_18870,N_18504);
nand U19285 (N_19285,N_18021,N_18475);
and U19286 (N_19286,N_18284,N_18272);
or U19287 (N_19287,N_18564,N_18156);
and U19288 (N_19288,N_18736,N_18562);
nand U19289 (N_19289,N_18860,N_18468);
nand U19290 (N_19290,N_18681,N_18397);
nor U19291 (N_19291,N_18525,N_18197);
nor U19292 (N_19292,N_18132,N_18084);
nand U19293 (N_19293,N_18303,N_18933);
nor U19294 (N_19294,N_18808,N_18236);
nand U19295 (N_19295,N_18083,N_18198);
nand U19296 (N_19296,N_18892,N_18690);
and U19297 (N_19297,N_18955,N_18492);
nor U19298 (N_19298,N_18735,N_18670);
xor U19299 (N_19299,N_18686,N_18127);
nor U19300 (N_19300,N_18402,N_18082);
or U19301 (N_19301,N_18046,N_18900);
nor U19302 (N_19302,N_18464,N_18345);
nand U19303 (N_19303,N_18273,N_18618);
nor U19304 (N_19304,N_18385,N_18026);
nand U19305 (N_19305,N_18058,N_18757);
nor U19306 (N_19306,N_18149,N_18429);
and U19307 (N_19307,N_18470,N_18370);
and U19308 (N_19308,N_18394,N_18268);
and U19309 (N_19309,N_18702,N_18179);
and U19310 (N_19310,N_18574,N_18661);
nor U19311 (N_19311,N_18662,N_18314);
and U19312 (N_19312,N_18552,N_18595);
xor U19313 (N_19313,N_18389,N_18418);
or U19314 (N_19314,N_18393,N_18378);
xor U19315 (N_19315,N_18099,N_18340);
xnor U19316 (N_19316,N_18420,N_18846);
xor U19317 (N_19317,N_18762,N_18189);
or U19318 (N_19318,N_18592,N_18360);
or U19319 (N_19319,N_18289,N_18332);
and U19320 (N_19320,N_18573,N_18852);
and U19321 (N_19321,N_18968,N_18128);
or U19322 (N_19322,N_18675,N_18356);
and U19323 (N_19323,N_18302,N_18430);
xor U19324 (N_19324,N_18548,N_18720);
nor U19325 (N_19325,N_18558,N_18886);
nor U19326 (N_19326,N_18152,N_18301);
xor U19327 (N_19327,N_18431,N_18031);
nor U19328 (N_19328,N_18350,N_18787);
nand U19329 (N_19329,N_18994,N_18652);
xnor U19330 (N_19330,N_18029,N_18226);
or U19331 (N_19331,N_18090,N_18448);
xor U19332 (N_19332,N_18593,N_18819);
nor U19333 (N_19333,N_18939,N_18836);
and U19334 (N_19334,N_18101,N_18219);
xnor U19335 (N_19335,N_18145,N_18195);
or U19336 (N_19336,N_18408,N_18732);
nor U19337 (N_19337,N_18353,N_18139);
and U19338 (N_19338,N_18815,N_18864);
xnor U19339 (N_19339,N_18905,N_18654);
nor U19340 (N_19340,N_18910,N_18610);
nor U19341 (N_19341,N_18244,N_18438);
xnor U19342 (N_19342,N_18364,N_18162);
nor U19343 (N_19343,N_18991,N_18390);
nor U19344 (N_19344,N_18498,N_18603);
xor U19345 (N_19345,N_18454,N_18254);
nand U19346 (N_19346,N_18977,N_18691);
or U19347 (N_19347,N_18155,N_18938);
and U19348 (N_19348,N_18798,N_18884);
and U19349 (N_19349,N_18714,N_18623);
or U19350 (N_19350,N_18563,N_18604);
nor U19351 (N_19351,N_18041,N_18500);
nand U19352 (N_19352,N_18568,N_18557);
xor U19353 (N_19353,N_18614,N_18981);
nand U19354 (N_19354,N_18883,N_18671);
or U19355 (N_19355,N_18274,N_18685);
nand U19356 (N_19356,N_18743,N_18582);
nor U19357 (N_19357,N_18192,N_18071);
or U19358 (N_19358,N_18628,N_18741);
or U19359 (N_19359,N_18751,N_18257);
xnor U19360 (N_19360,N_18134,N_18650);
and U19361 (N_19361,N_18142,N_18042);
and U19362 (N_19362,N_18918,N_18466);
nor U19363 (N_19363,N_18117,N_18478);
and U19364 (N_19364,N_18086,N_18212);
xor U19365 (N_19365,N_18790,N_18954);
nand U19366 (N_19366,N_18796,N_18432);
xnor U19367 (N_19367,N_18214,N_18359);
nor U19368 (N_19368,N_18154,N_18585);
and U19369 (N_19369,N_18813,N_18534);
xnor U19370 (N_19370,N_18979,N_18396);
nand U19371 (N_19371,N_18773,N_18253);
nand U19372 (N_19372,N_18817,N_18433);
xnor U19373 (N_19373,N_18006,N_18871);
and U19374 (N_19374,N_18611,N_18515);
or U19375 (N_19375,N_18882,N_18529);
nor U19376 (N_19376,N_18763,N_18249);
nor U19377 (N_19377,N_18946,N_18349);
xor U19378 (N_19378,N_18178,N_18105);
xor U19379 (N_19379,N_18013,N_18186);
nor U19380 (N_19380,N_18459,N_18213);
nor U19381 (N_19381,N_18241,N_18993);
and U19382 (N_19382,N_18633,N_18235);
and U19383 (N_19383,N_18321,N_18187);
and U19384 (N_19384,N_18508,N_18217);
xnor U19385 (N_19385,N_18121,N_18206);
nor U19386 (N_19386,N_18692,N_18701);
nand U19387 (N_19387,N_18594,N_18805);
nand U19388 (N_19388,N_18488,N_18894);
and U19389 (N_19389,N_18833,N_18588);
or U19390 (N_19390,N_18208,N_18779);
nor U19391 (N_19391,N_18298,N_18649);
xnor U19392 (N_19392,N_18673,N_18518);
nand U19393 (N_19393,N_18484,N_18028);
and U19394 (N_19394,N_18245,N_18577);
and U19395 (N_19395,N_18639,N_18295);
xor U19396 (N_19396,N_18334,N_18276);
and U19397 (N_19397,N_18941,N_18168);
and U19398 (N_19398,N_18881,N_18369);
xnor U19399 (N_19399,N_18477,N_18608);
or U19400 (N_19400,N_18267,N_18260);
nand U19401 (N_19401,N_18194,N_18166);
nor U19402 (N_19402,N_18695,N_18341);
nand U19403 (N_19403,N_18490,N_18978);
nor U19404 (N_19404,N_18828,N_18119);
or U19405 (N_19405,N_18856,N_18960);
nand U19406 (N_19406,N_18766,N_18575);
nand U19407 (N_19407,N_18312,N_18768);
nand U19408 (N_19408,N_18532,N_18271);
nand U19409 (N_19409,N_18699,N_18288);
nand U19410 (N_19410,N_18074,N_18216);
and U19411 (N_19411,N_18541,N_18053);
and U19412 (N_19412,N_18513,N_18823);
and U19413 (N_19413,N_18549,N_18998);
nor U19414 (N_19414,N_18612,N_18269);
nand U19415 (N_19415,N_18012,N_18304);
nand U19416 (N_19416,N_18103,N_18395);
nand U19417 (N_19417,N_18346,N_18780);
nor U19418 (N_19418,N_18051,N_18666);
or U19419 (N_19419,N_18818,N_18551);
nor U19420 (N_19420,N_18376,N_18286);
nor U19421 (N_19421,N_18647,N_18738);
or U19422 (N_19422,N_18970,N_18957);
nand U19423 (N_19423,N_18715,N_18294);
xor U19424 (N_19424,N_18296,N_18230);
and U19425 (N_19425,N_18381,N_18609);
and U19426 (N_19426,N_18927,N_18201);
or U19427 (N_19427,N_18710,N_18348);
or U19428 (N_19428,N_18266,N_18520);
nand U19429 (N_19429,N_18825,N_18259);
or U19430 (N_19430,N_18261,N_18959);
nor U19431 (N_19431,N_18472,N_18859);
nor U19432 (N_19432,N_18123,N_18812);
nor U19433 (N_19433,N_18157,N_18264);
xor U19434 (N_19434,N_18866,N_18311);
or U19435 (N_19435,N_18917,N_18228);
nor U19436 (N_19436,N_18607,N_18248);
xnor U19437 (N_19437,N_18837,N_18079);
and U19438 (N_19438,N_18962,N_18874);
xor U19439 (N_19439,N_18861,N_18361);
or U19440 (N_19440,N_18850,N_18450);
or U19441 (N_19441,N_18596,N_18005);
nand U19442 (N_19442,N_18631,N_18663);
nand U19443 (N_19443,N_18290,N_18409);
nor U19444 (N_19444,N_18164,N_18982);
nand U19445 (N_19445,N_18025,N_18597);
and U19446 (N_19446,N_18094,N_18275);
or U19447 (N_19447,N_18635,N_18832);
or U19448 (N_19448,N_18514,N_18405);
nor U19449 (N_19449,N_18352,N_18207);
nor U19450 (N_19450,N_18560,N_18229);
nand U19451 (N_19451,N_18964,N_18566);
xnor U19452 (N_19452,N_18044,N_18109);
nor U19453 (N_19453,N_18598,N_18967);
xor U19454 (N_19454,N_18845,N_18469);
or U19455 (N_19455,N_18471,N_18972);
xnor U19456 (N_19456,N_18567,N_18949);
nand U19457 (N_19457,N_18862,N_18211);
and U19458 (N_19458,N_18865,N_18387);
nor U19459 (N_19459,N_18482,N_18734);
or U19460 (N_19460,N_18406,N_18761);
or U19461 (N_19461,N_18110,N_18569);
or U19462 (N_19462,N_18137,N_18726);
and U19463 (N_19463,N_18651,N_18317);
or U19464 (N_19464,N_18100,N_18801);
nor U19465 (N_19465,N_18640,N_18331);
nand U19466 (N_19466,N_18672,N_18199);
nand U19467 (N_19467,N_18583,N_18499);
xor U19468 (N_19468,N_18320,N_18916);
nor U19469 (N_19469,N_18555,N_18767);
nand U19470 (N_19470,N_18943,N_18873);
xnor U19471 (N_19471,N_18748,N_18878);
nand U19472 (N_19472,N_18908,N_18196);
nor U19473 (N_19473,N_18721,N_18392);
nor U19474 (N_19474,N_18070,N_18600);
or U19475 (N_19475,N_18526,N_18746);
and U19476 (N_19476,N_18362,N_18934);
or U19477 (N_19477,N_18061,N_18434);
or U19478 (N_19478,N_18174,N_18619);
or U19479 (N_19479,N_18237,N_18624);
nand U19480 (N_19480,N_18565,N_18413);
xor U19481 (N_19481,N_18240,N_18875);
or U19482 (N_19482,N_18897,N_18637);
or U19483 (N_19483,N_18719,N_18252);
nor U19484 (N_19484,N_18323,N_18973);
nor U19485 (N_19485,N_18742,N_18447);
nor U19486 (N_19486,N_18183,N_18778);
nand U19487 (N_19487,N_18665,N_18147);
nand U19488 (N_19488,N_18221,N_18176);
or U19489 (N_19489,N_18124,N_18415);
nand U19490 (N_19490,N_18258,N_18613);
nor U19491 (N_19491,N_18648,N_18399);
nand U19492 (N_19492,N_18263,N_18182);
and U19493 (N_19493,N_18570,N_18559);
xnor U19494 (N_19494,N_18816,N_18831);
or U19495 (N_19495,N_18338,N_18693);
nand U19496 (N_19496,N_18963,N_18161);
or U19497 (N_19497,N_18961,N_18227);
and U19498 (N_19498,N_18929,N_18951);
xnor U19499 (N_19499,N_18368,N_18524);
and U19500 (N_19500,N_18132,N_18727);
xor U19501 (N_19501,N_18618,N_18085);
nor U19502 (N_19502,N_18513,N_18396);
xnor U19503 (N_19503,N_18709,N_18901);
or U19504 (N_19504,N_18567,N_18599);
and U19505 (N_19505,N_18376,N_18471);
nor U19506 (N_19506,N_18382,N_18663);
or U19507 (N_19507,N_18890,N_18892);
or U19508 (N_19508,N_18465,N_18883);
nand U19509 (N_19509,N_18356,N_18401);
nor U19510 (N_19510,N_18170,N_18571);
nand U19511 (N_19511,N_18871,N_18042);
nand U19512 (N_19512,N_18968,N_18648);
nor U19513 (N_19513,N_18683,N_18664);
nand U19514 (N_19514,N_18385,N_18896);
or U19515 (N_19515,N_18834,N_18531);
nor U19516 (N_19516,N_18438,N_18715);
xor U19517 (N_19517,N_18377,N_18636);
xor U19518 (N_19518,N_18045,N_18239);
or U19519 (N_19519,N_18391,N_18835);
xnor U19520 (N_19520,N_18167,N_18432);
xnor U19521 (N_19521,N_18359,N_18475);
nand U19522 (N_19522,N_18071,N_18874);
xor U19523 (N_19523,N_18521,N_18262);
xor U19524 (N_19524,N_18058,N_18035);
or U19525 (N_19525,N_18889,N_18188);
nand U19526 (N_19526,N_18179,N_18601);
or U19527 (N_19527,N_18677,N_18972);
and U19528 (N_19528,N_18713,N_18896);
nor U19529 (N_19529,N_18245,N_18686);
and U19530 (N_19530,N_18447,N_18564);
or U19531 (N_19531,N_18330,N_18635);
or U19532 (N_19532,N_18685,N_18923);
xor U19533 (N_19533,N_18597,N_18726);
xor U19534 (N_19534,N_18702,N_18292);
or U19535 (N_19535,N_18175,N_18497);
nor U19536 (N_19536,N_18737,N_18419);
and U19537 (N_19537,N_18526,N_18039);
nand U19538 (N_19538,N_18654,N_18396);
nand U19539 (N_19539,N_18641,N_18683);
nor U19540 (N_19540,N_18666,N_18354);
nand U19541 (N_19541,N_18949,N_18974);
nor U19542 (N_19542,N_18886,N_18581);
nand U19543 (N_19543,N_18807,N_18192);
xnor U19544 (N_19544,N_18062,N_18083);
nor U19545 (N_19545,N_18415,N_18802);
nand U19546 (N_19546,N_18821,N_18077);
nand U19547 (N_19547,N_18441,N_18657);
nor U19548 (N_19548,N_18995,N_18301);
nand U19549 (N_19549,N_18345,N_18538);
xor U19550 (N_19550,N_18494,N_18917);
xnor U19551 (N_19551,N_18959,N_18965);
nor U19552 (N_19552,N_18617,N_18695);
nor U19553 (N_19553,N_18375,N_18512);
xor U19554 (N_19554,N_18169,N_18287);
nand U19555 (N_19555,N_18676,N_18490);
and U19556 (N_19556,N_18361,N_18801);
and U19557 (N_19557,N_18943,N_18700);
xor U19558 (N_19558,N_18873,N_18099);
or U19559 (N_19559,N_18298,N_18949);
xnor U19560 (N_19560,N_18510,N_18952);
nor U19561 (N_19561,N_18566,N_18984);
and U19562 (N_19562,N_18746,N_18827);
xor U19563 (N_19563,N_18347,N_18659);
nor U19564 (N_19564,N_18310,N_18572);
xor U19565 (N_19565,N_18782,N_18718);
xnor U19566 (N_19566,N_18818,N_18064);
or U19567 (N_19567,N_18493,N_18356);
and U19568 (N_19568,N_18378,N_18560);
and U19569 (N_19569,N_18786,N_18145);
xor U19570 (N_19570,N_18036,N_18551);
and U19571 (N_19571,N_18993,N_18222);
and U19572 (N_19572,N_18471,N_18722);
nand U19573 (N_19573,N_18474,N_18973);
nor U19574 (N_19574,N_18136,N_18368);
or U19575 (N_19575,N_18669,N_18693);
or U19576 (N_19576,N_18495,N_18754);
and U19577 (N_19577,N_18253,N_18828);
or U19578 (N_19578,N_18112,N_18140);
nor U19579 (N_19579,N_18187,N_18817);
xnor U19580 (N_19580,N_18744,N_18815);
nor U19581 (N_19581,N_18252,N_18159);
nand U19582 (N_19582,N_18394,N_18222);
nor U19583 (N_19583,N_18693,N_18783);
nor U19584 (N_19584,N_18750,N_18960);
nor U19585 (N_19585,N_18122,N_18327);
and U19586 (N_19586,N_18002,N_18415);
nand U19587 (N_19587,N_18111,N_18837);
and U19588 (N_19588,N_18033,N_18612);
or U19589 (N_19589,N_18380,N_18696);
and U19590 (N_19590,N_18940,N_18403);
xnor U19591 (N_19591,N_18315,N_18899);
and U19592 (N_19592,N_18225,N_18346);
nand U19593 (N_19593,N_18391,N_18616);
nand U19594 (N_19594,N_18673,N_18132);
xnor U19595 (N_19595,N_18254,N_18141);
nand U19596 (N_19596,N_18630,N_18274);
nand U19597 (N_19597,N_18838,N_18516);
or U19598 (N_19598,N_18351,N_18092);
or U19599 (N_19599,N_18707,N_18209);
nand U19600 (N_19600,N_18895,N_18849);
nor U19601 (N_19601,N_18352,N_18065);
and U19602 (N_19602,N_18953,N_18839);
and U19603 (N_19603,N_18809,N_18550);
nand U19604 (N_19604,N_18367,N_18097);
nand U19605 (N_19605,N_18841,N_18951);
and U19606 (N_19606,N_18945,N_18743);
nand U19607 (N_19607,N_18374,N_18654);
and U19608 (N_19608,N_18541,N_18307);
or U19609 (N_19609,N_18515,N_18973);
and U19610 (N_19610,N_18749,N_18767);
or U19611 (N_19611,N_18955,N_18590);
or U19612 (N_19612,N_18354,N_18787);
nand U19613 (N_19613,N_18442,N_18554);
nand U19614 (N_19614,N_18708,N_18985);
and U19615 (N_19615,N_18263,N_18243);
xnor U19616 (N_19616,N_18335,N_18812);
and U19617 (N_19617,N_18743,N_18624);
or U19618 (N_19618,N_18006,N_18009);
nor U19619 (N_19619,N_18408,N_18175);
and U19620 (N_19620,N_18984,N_18093);
and U19621 (N_19621,N_18993,N_18141);
and U19622 (N_19622,N_18524,N_18646);
or U19623 (N_19623,N_18562,N_18116);
xnor U19624 (N_19624,N_18620,N_18977);
nor U19625 (N_19625,N_18092,N_18505);
or U19626 (N_19626,N_18113,N_18763);
nand U19627 (N_19627,N_18229,N_18159);
and U19628 (N_19628,N_18122,N_18739);
or U19629 (N_19629,N_18045,N_18153);
nor U19630 (N_19630,N_18742,N_18274);
xor U19631 (N_19631,N_18129,N_18617);
xnor U19632 (N_19632,N_18127,N_18183);
and U19633 (N_19633,N_18166,N_18519);
or U19634 (N_19634,N_18623,N_18971);
nor U19635 (N_19635,N_18658,N_18510);
and U19636 (N_19636,N_18042,N_18680);
xnor U19637 (N_19637,N_18472,N_18596);
nand U19638 (N_19638,N_18125,N_18661);
nor U19639 (N_19639,N_18145,N_18749);
and U19640 (N_19640,N_18281,N_18059);
and U19641 (N_19641,N_18986,N_18257);
and U19642 (N_19642,N_18591,N_18770);
or U19643 (N_19643,N_18640,N_18979);
or U19644 (N_19644,N_18358,N_18671);
nand U19645 (N_19645,N_18997,N_18276);
nand U19646 (N_19646,N_18788,N_18522);
nand U19647 (N_19647,N_18941,N_18795);
nand U19648 (N_19648,N_18660,N_18000);
nand U19649 (N_19649,N_18539,N_18014);
xor U19650 (N_19650,N_18980,N_18252);
nor U19651 (N_19651,N_18998,N_18278);
nor U19652 (N_19652,N_18165,N_18039);
or U19653 (N_19653,N_18388,N_18648);
or U19654 (N_19654,N_18697,N_18884);
nor U19655 (N_19655,N_18104,N_18314);
nor U19656 (N_19656,N_18776,N_18824);
nor U19657 (N_19657,N_18265,N_18351);
or U19658 (N_19658,N_18920,N_18672);
nand U19659 (N_19659,N_18449,N_18074);
nand U19660 (N_19660,N_18274,N_18493);
or U19661 (N_19661,N_18782,N_18445);
nor U19662 (N_19662,N_18244,N_18979);
and U19663 (N_19663,N_18185,N_18823);
and U19664 (N_19664,N_18934,N_18439);
or U19665 (N_19665,N_18752,N_18429);
nor U19666 (N_19666,N_18993,N_18348);
nand U19667 (N_19667,N_18886,N_18679);
xnor U19668 (N_19668,N_18528,N_18509);
or U19669 (N_19669,N_18231,N_18520);
nand U19670 (N_19670,N_18066,N_18393);
nor U19671 (N_19671,N_18435,N_18210);
and U19672 (N_19672,N_18966,N_18319);
xor U19673 (N_19673,N_18829,N_18450);
or U19674 (N_19674,N_18390,N_18901);
or U19675 (N_19675,N_18712,N_18829);
nor U19676 (N_19676,N_18779,N_18058);
nor U19677 (N_19677,N_18879,N_18751);
and U19678 (N_19678,N_18743,N_18971);
nand U19679 (N_19679,N_18766,N_18864);
nand U19680 (N_19680,N_18613,N_18005);
xnor U19681 (N_19681,N_18681,N_18904);
nor U19682 (N_19682,N_18639,N_18910);
xnor U19683 (N_19683,N_18257,N_18686);
nand U19684 (N_19684,N_18134,N_18957);
and U19685 (N_19685,N_18981,N_18269);
or U19686 (N_19686,N_18260,N_18873);
nand U19687 (N_19687,N_18922,N_18429);
or U19688 (N_19688,N_18602,N_18698);
xnor U19689 (N_19689,N_18445,N_18625);
and U19690 (N_19690,N_18767,N_18430);
nand U19691 (N_19691,N_18009,N_18805);
nand U19692 (N_19692,N_18649,N_18764);
xor U19693 (N_19693,N_18530,N_18376);
nor U19694 (N_19694,N_18520,N_18530);
nor U19695 (N_19695,N_18496,N_18324);
or U19696 (N_19696,N_18877,N_18221);
nand U19697 (N_19697,N_18311,N_18563);
xnor U19698 (N_19698,N_18856,N_18773);
nor U19699 (N_19699,N_18949,N_18101);
xor U19700 (N_19700,N_18030,N_18052);
xor U19701 (N_19701,N_18054,N_18840);
xor U19702 (N_19702,N_18265,N_18438);
nor U19703 (N_19703,N_18481,N_18307);
nor U19704 (N_19704,N_18962,N_18640);
or U19705 (N_19705,N_18365,N_18963);
xor U19706 (N_19706,N_18897,N_18962);
or U19707 (N_19707,N_18951,N_18367);
xnor U19708 (N_19708,N_18328,N_18044);
and U19709 (N_19709,N_18519,N_18859);
and U19710 (N_19710,N_18714,N_18255);
and U19711 (N_19711,N_18647,N_18111);
nand U19712 (N_19712,N_18988,N_18506);
or U19713 (N_19713,N_18471,N_18289);
nand U19714 (N_19714,N_18037,N_18511);
nor U19715 (N_19715,N_18352,N_18346);
nor U19716 (N_19716,N_18183,N_18957);
or U19717 (N_19717,N_18557,N_18174);
and U19718 (N_19718,N_18302,N_18208);
or U19719 (N_19719,N_18784,N_18012);
nand U19720 (N_19720,N_18956,N_18741);
or U19721 (N_19721,N_18013,N_18371);
or U19722 (N_19722,N_18062,N_18655);
xor U19723 (N_19723,N_18615,N_18649);
and U19724 (N_19724,N_18087,N_18148);
nand U19725 (N_19725,N_18250,N_18212);
nor U19726 (N_19726,N_18496,N_18111);
or U19727 (N_19727,N_18962,N_18360);
and U19728 (N_19728,N_18369,N_18288);
xor U19729 (N_19729,N_18101,N_18836);
and U19730 (N_19730,N_18009,N_18750);
nor U19731 (N_19731,N_18828,N_18695);
and U19732 (N_19732,N_18309,N_18761);
xnor U19733 (N_19733,N_18114,N_18838);
nor U19734 (N_19734,N_18542,N_18151);
nand U19735 (N_19735,N_18688,N_18247);
or U19736 (N_19736,N_18309,N_18812);
nor U19737 (N_19737,N_18487,N_18548);
nor U19738 (N_19738,N_18003,N_18567);
nand U19739 (N_19739,N_18584,N_18315);
or U19740 (N_19740,N_18748,N_18310);
or U19741 (N_19741,N_18430,N_18939);
and U19742 (N_19742,N_18176,N_18106);
and U19743 (N_19743,N_18956,N_18332);
and U19744 (N_19744,N_18616,N_18795);
xnor U19745 (N_19745,N_18194,N_18906);
or U19746 (N_19746,N_18204,N_18449);
nand U19747 (N_19747,N_18939,N_18111);
nor U19748 (N_19748,N_18480,N_18543);
nand U19749 (N_19749,N_18100,N_18580);
nor U19750 (N_19750,N_18022,N_18267);
or U19751 (N_19751,N_18349,N_18297);
and U19752 (N_19752,N_18625,N_18615);
nand U19753 (N_19753,N_18980,N_18204);
and U19754 (N_19754,N_18651,N_18793);
or U19755 (N_19755,N_18700,N_18632);
nand U19756 (N_19756,N_18344,N_18731);
nand U19757 (N_19757,N_18909,N_18320);
and U19758 (N_19758,N_18225,N_18042);
and U19759 (N_19759,N_18113,N_18032);
or U19760 (N_19760,N_18964,N_18907);
nor U19761 (N_19761,N_18789,N_18849);
nand U19762 (N_19762,N_18933,N_18980);
nand U19763 (N_19763,N_18070,N_18347);
xor U19764 (N_19764,N_18472,N_18118);
nor U19765 (N_19765,N_18177,N_18676);
nor U19766 (N_19766,N_18176,N_18083);
nor U19767 (N_19767,N_18213,N_18366);
and U19768 (N_19768,N_18009,N_18410);
and U19769 (N_19769,N_18723,N_18653);
nand U19770 (N_19770,N_18723,N_18604);
or U19771 (N_19771,N_18753,N_18587);
nor U19772 (N_19772,N_18678,N_18315);
and U19773 (N_19773,N_18854,N_18892);
nand U19774 (N_19774,N_18256,N_18851);
nor U19775 (N_19775,N_18021,N_18439);
xor U19776 (N_19776,N_18189,N_18583);
or U19777 (N_19777,N_18967,N_18729);
nand U19778 (N_19778,N_18397,N_18176);
xnor U19779 (N_19779,N_18262,N_18625);
or U19780 (N_19780,N_18286,N_18504);
and U19781 (N_19781,N_18019,N_18824);
and U19782 (N_19782,N_18459,N_18466);
or U19783 (N_19783,N_18363,N_18886);
nand U19784 (N_19784,N_18642,N_18695);
or U19785 (N_19785,N_18632,N_18836);
and U19786 (N_19786,N_18793,N_18131);
or U19787 (N_19787,N_18733,N_18872);
xor U19788 (N_19788,N_18984,N_18876);
nor U19789 (N_19789,N_18999,N_18260);
or U19790 (N_19790,N_18864,N_18783);
nor U19791 (N_19791,N_18447,N_18962);
or U19792 (N_19792,N_18198,N_18739);
nand U19793 (N_19793,N_18769,N_18892);
nand U19794 (N_19794,N_18584,N_18113);
or U19795 (N_19795,N_18538,N_18261);
or U19796 (N_19796,N_18093,N_18445);
and U19797 (N_19797,N_18126,N_18230);
nand U19798 (N_19798,N_18137,N_18173);
or U19799 (N_19799,N_18572,N_18033);
or U19800 (N_19800,N_18673,N_18416);
nand U19801 (N_19801,N_18355,N_18148);
nor U19802 (N_19802,N_18536,N_18641);
nand U19803 (N_19803,N_18826,N_18814);
xor U19804 (N_19804,N_18231,N_18280);
nor U19805 (N_19805,N_18741,N_18195);
nand U19806 (N_19806,N_18558,N_18638);
or U19807 (N_19807,N_18906,N_18282);
nor U19808 (N_19808,N_18642,N_18177);
or U19809 (N_19809,N_18865,N_18416);
or U19810 (N_19810,N_18273,N_18328);
xor U19811 (N_19811,N_18518,N_18457);
and U19812 (N_19812,N_18620,N_18489);
and U19813 (N_19813,N_18933,N_18307);
and U19814 (N_19814,N_18038,N_18002);
or U19815 (N_19815,N_18317,N_18959);
nor U19816 (N_19816,N_18850,N_18711);
or U19817 (N_19817,N_18031,N_18320);
or U19818 (N_19818,N_18635,N_18955);
or U19819 (N_19819,N_18973,N_18473);
nor U19820 (N_19820,N_18500,N_18712);
nor U19821 (N_19821,N_18825,N_18355);
nand U19822 (N_19822,N_18680,N_18437);
xor U19823 (N_19823,N_18315,N_18548);
nand U19824 (N_19824,N_18785,N_18332);
or U19825 (N_19825,N_18301,N_18286);
and U19826 (N_19826,N_18907,N_18201);
or U19827 (N_19827,N_18458,N_18960);
nor U19828 (N_19828,N_18649,N_18095);
or U19829 (N_19829,N_18685,N_18699);
xor U19830 (N_19830,N_18671,N_18432);
nor U19831 (N_19831,N_18555,N_18095);
nor U19832 (N_19832,N_18460,N_18257);
nor U19833 (N_19833,N_18663,N_18492);
and U19834 (N_19834,N_18892,N_18177);
or U19835 (N_19835,N_18063,N_18070);
and U19836 (N_19836,N_18925,N_18427);
nand U19837 (N_19837,N_18746,N_18799);
nor U19838 (N_19838,N_18505,N_18728);
nand U19839 (N_19839,N_18314,N_18821);
or U19840 (N_19840,N_18625,N_18838);
nor U19841 (N_19841,N_18520,N_18663);
or U19842 (N_19842,N_18391,N_18841);
nand U19843 (N_19843,N_18894,N_18133);
xor U19844 (N_19844,N_18832,N_18350);
or U19845 (N_19845,N_18214,N_18969);
and U19846 (N_19846,N_18377,N_18460);
xnor U19847 (N_19847,N_18538,N_18554);
xor U19848 (N_19848,N_18614,N_18766);
xnor U19849 (N_19849,N_18110,N_18611);
nand U19850 (N_19850,N_18583,N_18844);
nand U19851 (N_19851,N_18869,N_18440);
nand U19852 (N_19852,N_18079,N_18738);
xnor U19853 (N_19853,N_18975,N_18243);
or U19854 (N_19854,N_18683,N_18349);
nand U19855 (N_19855,N_18915,N_18307);
nor U19856 (N_19856,N_18156,N_18457);
or U19857 (N_19857,N_18474,N_18485);
nor U19858 (N_19858,N_18155,N_18287);
xnor U19859 (N_19859,N_18941,N_18934);
nor U19860 (N_19860,N_18900,N_18029);
nand U19861 (N_19861,N_18630,N_18572);
nor U19862 (N_19862,N_18760,N_18223);
and U19863 (N_19863,N_18908,N_18272);
nand U19864 (N_19864,N_18455,N_18607);
and U19865 (N_19865,N_18414,N_18688);
or U19866 (N_19866,N_18161,N_18397);
xor U19867 (N_19867,N_18610,N_18134);
xor U19868 (N_19868,N_18191,N_18796);
xnor U19869 (N_19869,N_18744,N_18766);
nand U19870 (N_19870,N_18375,N_18108);
and U19871 (N_19871,N_18324,N_18292);
xnor U19872 (N_19872,N_18728,N_18967);
nand U19873 (N_19873,N_18513,N_18761);
or U19874 (N_19874,N_18369,N_18910);
nor U19875 (N_19875,N_18955,N_18142);
xnor U19876 (N_19876,N_18469,N_18718);
or U19877 (N_19877,N_18036,N_18089);
or U19878 (N_19878,N_18240,N_18502);
or U19879 (N_19879,N_18309,N_18687);
and U19880 (N_19880,N_18023,N_18597);
nand U19881 (N_19881,N_18096,N_18945);
or U19882 (N_19882,N_18949,N_18917);
xnor U19883 (N_19883,N_18057,N_18020);
nor U19884 (N_19884,N_18482,N_18494);
and U19885 (N_19885,N_18658,N_18817);
nand U19886 (N_19886,N_18173,N_18154);
nand U19887 (N_19887,N_18742,N_18655);
nand U19888 (N_19888,N_18742,N_18276);
and U19889 (N_19889,N_18572,N_18142);
nor U19890 (N_19890,N_18021,N_18147);
and U19891 (N_19891,N_18472,N_18068);
nand U19892 (N_19892,N_18156,N_18561);
nor U19893 (N_19893,N_18634,N_18330);
nor U19894 (N_19894,N_18778,N_18075);
and U19895 (N_19895,N_18163,N_18612);
and U19896 (N_19896,N_18060,N_18748);
xor U19897 (N_19897,N_18080,N_18011);
and U19898 (N_19898,N_18514,N_18631);
nor U19899 (N_19899,N_18035,N_18878);
xor U19900 (N_19900,N_18561,N_18162);
xnor U19901 (N_19901,N_18664,N_18992);
or U19902 (N_19902,N_18314,N_18737);
and U19903 (N_19903,N_18642,N_18383);
nor U19904 (N_19904,N_18348,N_18199);
nor U19905 (N_19905,N_18807,N_18655);
nand U19906 (N_19906,N_18726,N_18206);
or U19907 (N_19907,N_18224,N_18475);
xor U19908 (N_19908,N_18597,N_18476);
xor U19909 (N_19909,N_18095,N_18073);
xor U19910 (N_19910,N_18679,N_18846);
nand U19911 (N_19911,N_18063,N_18663);
nand U19912 (N_19912,N_18420,N_18937);
nand U19913 (N_19913,N_18023,N_18923);
nor U19914 (N_19914,N_18891,N_18522);
or U19915 (N_19915,N_18930,N_18757);
or U19916 (N_19916,N_18247,N_18462);
xor U19917 (N_19917,N_18442,N_18248);
or U19918 (N_19918,N_18484,N_18834);
nand U19919 (N_19919,N_18515,N_18732);
or U19920 (N_19920,N_18416,N_18135);
or U19921 (N_19921,N_18284,N_18195);
or U19922 (N_19922,N_18263,N_18844);
nor U19923 (N_19923,N_18378,N_18831);
nor U19924 (N_19924,N_18357,N_18696);
nand U19925 (N_19925,N_18004,N_18529);
nor U19926 (N_19926,N_18409,N_18814);
nor U19927 (N_19927,N_18928,N_18797);
nand U19928 (N_19928,N_18024,N_18895);
xnor U19929 (N_19929,N_18602,N_18717);
nand U19930 (N_19930,N_18257,N_18827);
or U19931 (N_19931,N_18315,N_18838);
or U19932 (N_19932,N_18800,N_18913);
nand U19933 (N_19933,N_18170,N_18052);
or U19934 (N_19934,N_18083,N_18161);
nand U19935 (N_19935,N_18123,N_18348);
nor U19936 (N_19936,N_18188,N_18907);
nand U19937 (N_19937,N_18712,N_18298);
and U19938 (N_19938,N_18617,N_18986);
xor U19939 (N_19939,N_18504,N_18527);
nor U19940 (N_19940,N_18928,N_18011);
nor U19941 (N_19941,N_18737,N_18755);
or U19942 (N_19942,N_18178,N_18146);
and U19943 (N_19943,N_18765,N_18636);
nand U19944 (N_19944,N_18077,N_18179);
xor U19945 (N_19945,N_18891,N_18729);
nor U19946 (N_19946,N_18677,N_18740);
or U19947 (N_19947,N_18390,N_18444);
nor U19948 (N_19948,N_18773,N_18720);
and U19949 (N_19949,N_18980,N_18601);
or U19950 (N_19950,N_18312,N_18598);
or U19951 (N_19951,N_18905,N_18116);
and U19952 (N_19952,N_18915,N_18482);
nor U19953 (N_19953,N_18523,N_18104);
and U19954 (N_19954,N_18377,N_18678);
xor U19955 (N_19955,N_18285,N_18996);
nand U19956 (N_19956,N_18549,N_18825);
nand U19957 (N_19957,N_18605,N_18527);
nand U19958 (N_19958,N_18778,N_18781);
xor U19959 (N_19959,N_18195,N_18317);
and U19960 (N_19960,N_18974,N_18514);
and U19961 (N_19961,N_18003,N_18612);
and U19962 (N_19962,N_18745,N_18073);
nand U19963 (N_19963,N_18656,N_18552);
xnor U19964 (N_19964,N_18174,N_18220);
nand U19965 (N_19965,N_18528,N_18267);
nor U19966 (N_19966,N_18972,N_18655);
nand U19967 (N_19967,N_18977,N_18855);
or U19968 (N_19968,N_18916,N_18945);
xnor U19969 (N_19969,N_18012,N_18822);
or U19970 (N_19970,N_18106,N_18284);
and U19971 (N_19971,N_18736,N_18427);
or U19972 (N_19972,N_18754,N_18053);
or U19973 (N_19973,N_18983,N_18424);
or U19974 (N_19974,N_18222,N_18553);
and U19975 (N_19975,N_18654,N_18119);
nand U19976 (N_19976,N_18225,N_18664);
or U19977 (N_19977,N_18839,N_18454);
xnor U19978 (N_19978,N_18032,N_18745);
nand U19979 (N_19979,N_18413,N_18077);
and U19980 (N_19980,N_18802,N_18246);
or U19981 (N_19981,N_18552,N_18941);
nor U19982 (N_19982,N_18472,N_18694);
and U19983 (N_19983,N_18873,N_18505);
or U19984 (N_19984,N_18738,N_18781);
nor U19985 (N_19985,N_18779,N_18558);
or U19986 (N_19986,N_18764,N_18478);
xnor U19987 (N_19987,N_18263,N_18589);
xor U19988 (N_19988,N_18349,N_18678);
nand U19989 (N_19989,N_18068,N_18787);
nand U19990 (N_19990,N_18910,N_18199);
nor U19991 (N_19991,N_18805,N_18140);
xnor U19992 (N_19992,N_18390,N_18293);
and U19993 (N_19993,N_18342,N_18178);
nand U19994 (N_19994,N_18857,N_18021);
xor U19995 (N_19995,N_18431,N_18770);
and U19996 (N_19996,N_18318,N_18964);
or U19997 (N_19997,N_18349,N_18854);
nor U19998 (N_19998,N_18557,N_18932);
nor U19999 (N_19999,N_18546,N_18121);
or U20000 (N_20000,N_19847,N_19440);
nand U20001 (N_20001,N_19928,N_19115);
xor U20002 (N_20002,N_19237,N_19257);
or U20003 (N_20003,N_19932,N_19621);
and U20004 (N_20004,N_19233,N_19234);
nand U20005 (N_20005,N_19977,N_19147);
nor U20006 (N_20006,N_19341,N_19390);
and U20007 (N_20007,N_19904,N_19391);
and U20008 (N_20008,N_19017,N_19696);
nand U20009 (N_20009,N_19502,N_19172);
and U20010 (N_20010,N_19965,N_19357);
or U20011 (N_20011,N_19080,N_19191);
nor U20012 (N_20012,N_19458,N_19134);
or U20013 (N_20013,N_19307,N_19516);
and U20014 (N_20014,N_19765,N_19285);
nor U20015 (N_20015,N_19367,N_19102);
or U20016 (N_20016,N_19745,N_19418);
nor U20017 (N_20017,N_19706,N_19204);
and U20018 (N_20018,N_19700,N_19856);
nand U20019 (N_20019,N_19072,N_19784);
or U20020 (N_20020,N_19888,N_19301);
and U20021 (N_20021,N_19068,N_19826);
nand U20022 (N_20022,N_19135,N_19945);
and U20023 (N_20023,N_19279,N_19531);
xnor U20024 (N_20024,N_19109,N_19774);
nand U20025 (N_20025,N_19708,N_19808);
or U20026 (N_20026,N_19073,N_19805);
nand U20027 (N_20027,N_19771,N_19554);
xor U20028 (N_20028,N_19047,N_19840);
nor U20029 (N_20029,N_19255,N_19055);
xnor U20030 (N_20030,N_19915,N_19665);
or U20031 (N_20031,N_19356,N_19780);
and U20032 (N_20032,N_19354,N_19373);
xnor U20033 (N_20033,N_19087,N_19952);
and U20034 (N_20034,N_19836,N_19226);
nand U20035 (N_20035,N_19036,N_19295);
nand U20036 (N_20036,N_19327,N_19388);
xor U20037 (N_20037,N_19911,N_19930);
or U20038 (N_20038,N_19586,N_19697);
xnor U20039 (N_20039,N_19576,N_19180);
and U20040 (N_20040,N_19882,N_19743);
nand U20041 (N_20041,N_19997,N_19927);
xor U20042 (N_20042,N_19312,N_19564);
nor U20043 (N_20043,N_19719,N_19310);
or U20044 (N_20044,N_19528,N_19221);
xnor U20045 (N_20045,N_19013,N_19627);
or U20046 (N_20046,N_19566,N_19455);
nor U20047 (N_20047,N_19942,N_19283);
xor U20048 (N_20048,N_19416,N_19358);
nand U20049 (N_20049,N_19175,N_19355);
and U20050 (N_20050,N_19588,N_19287);
or U20051 (N_20051,N_19081,N_19173);
nor U20052 (N_20052,N_19262,N_19640);
or U20053 (N_20053,N_19452,N_19432);
nor U20054 (N_20054,N_19804,N_19251);
and U20055 (N_20055,N_19306,N_19832);
xor U20056 (N_20056,N_19595,N_19404);
or U20057 (N_20057,N_19485,N_19955);
nor U20058 (N_20058,N_19426,N_19843);
xnor U20059 (N_20059,N_19489,N_19508);
nor U20060 (N_20060,N_19905,N_19037);
xnor U20061 (N_20061,N_19145,N_19558);
and U20062 (N_20062,N_19764,N_19515);
or U20063 (N_20063,N_19641,N_19420);
and U20064 (N_20064,N_19596,N_19645);
nand U20065 (N_20065,N_19960,N_19325);
xor U20066 (N_20066,N_19095,N_19408);
nor U20067 (N_20067,N_19041,N_19166);
xnor U20068 (N_20068,N_19061,N_19230);
xnor U20069 (N_20069,N_19791,N_19031);
xor U20070 (N_20070,N_19304,N_19079);
nand U20071 (N_20071,N_19296,N_19948);
nor U20072 (N_20072,N_19660,N_19813);
or U20073 (N_20073,N_19735,N_19909);
and U20074 (N_20074,N_19239,N_19877);
xnor U20075 (N_20075,N_19857,N_19321);
xnor U20076 (N_20076,N_19574,N_19203);
xor U20077 (N_20077,N_19940,N_19323);
or U20078 (N_20078,N_19873,N_19028);
xor U20079 (N_20079,N_19365,N_19484);
nor U20080 (N_20080,N_19549,N_19620);
or U20081 (N_20081,N_19065,N_19991);
and U20082 (N_20082,N_19106,N_19579);
xor U20083 (N_20083,N_19842,N_19394);
and U20084 (N_20084,N_19683,N_19395);
xor U20085 (N_20085,N_19957,N_19985);
and U20086 (N_20086,N_19936,N_19693);
nor U20087 (N_20087,N_19529,N_19015);
xnor U20088 (N_20088,N_19199,N_19934);
and U20089 (N_20089,N_19274,N_19427);
nand U20090 (N_20090,N_19503,N_19205);
nand U20091 (N_20091,N_19319,N_19220);
nor U20092 (N_20092,N_19256,N_19371);
xnor U20093 (N_20093,N_19753,N_19801);
and U20094 (N_20094,N_19755,N_19012);
or U20095 (N_20095,N_19849,N_19639);
or U20096 (N_20096,N_19157,N_19907);
and U20097 (N_20097,N_19864,N_19286);
nand U20098 (N_20098,N_19309,N_19326);
nand U20099 (N_20099,N_19868,N_19789);
or U20100 (N_20100,N_19742,N_19439);
and U20101 (N_20101,N_19885,N_19751);
nand U20102 (N_20102,N_19786,N_19874);
nor U20103 (N_20103,N_19176,N_19889);
xnor U20104 (N_20104,N_19602,N_19214);
and U20105 (N_20105,N_19563,N_19430);
or U20106 (N_20106,N_19401,N_19605);
nand U20107 (N_20107,N_19634,N_19348);
and U20108 (N_20108,N_19225,N_19057);
xor U20109 (N_20109,N_19547,N_19591);
nand U20110 (N_20110,N_19510,N_19078);
xnor U20111 (N_20111,N_19402,N_19798);
nand U20112 (N_20112,N_19335,N_19378);
or U20113 (N_20113,N_19881,N_19763);
nand U20114 (N_20114,N_19520,N_19672);
nand U20115 (N_20115,N_19398,N_19974);
or U20116 (N_20116,N_19760,N_19730);
xor U20117 (N_20117,N_19681,N_19897);
nand U20118 (N_20118,N_19958,N_19436);
or U20119 (N_20119,N_19030,N_19623);
or U20120 (N_20120,N_19343,N_19916);
and U20121 (N_20121,N_19198,N_19463);
or U20122 (N_20122,N_19837,N_19071);
or U20123 (N_20123,N_19718,N_19263);
or U20124 (N_20124,N_19186,N_19662);
or U20125 (N_20125,N_19514,N_19770);
xnor U20126 (N_20126,N_19018,N_19497);
or U20127 (N_20127,N_19592,N_19034);
and U20128 (N_20128,N_19369,N_19494);
or U20129 (N_20129,N_19351,N_19601);
and U20130 (N_20130,N_19901,N_19224);
and U20131 (N_20131,N_19130,N_19112);
nand U20132 (N_20132,N_19195,N_19815);
nor U20133 (N_20133,N_19089,N_19350);
or U20134 (N_20134,N_19557,N_19773);
xor U20135 (N_20135,N_19535,N_19141);
xor U20136 (N_20136,N_19407,N_19025);
and U20137 (N_20137,N_19161,N_19121);
and U20138 (N_20138,N_19179,N_19118);
and U20139 (N_20139,N_19769,N_19260);
nand U20140 (N_20140,N_19893,N_19469);
nand U20141 (N_20141,N_19600,N_19336);
nor U20142 (N_20142,N_19984,N_19340);
or U20143 (N_20143,N_19655,N_19626);
and U20144 (N_20144,N_19707,N_19020);
or U20145 (N_20145,N_19069,N_19006);
xor U20146 (N_20146,N_19438,N_19537);
nand U20147 (N_20147,N_19562,N_19480);
xnor U20148 (N_20148,N_19527,N_19450);
and U20149 (N_20149,N_19154,N_19058);
xnor U20150 (N_20150,N_19261,N_19858);
nor U20151 (N_20151,N_19649,N_19242);
or U20152 (N_20152,N_19748,N_19419);
nor U20153 (N_20153,N_19216,N_19648);
nand U20154 (N_20154,N_19334,N_19787);
xor U20155 (N_20155,N_19616,N_19636);
or U20156 (N_20156,N_19010,N_19218);
nor U20157 (N_20157,N_19315,N_19617);
nand U20158 (N_20158,N_19859,N_19946);
or U20159 (N_20159,N_19076,N_19924);
or U20160 (N_20160,N_19680,N_19139);
and U20161 (N_20161,N_19133,N_19572);
or U20162 (N_20162,N_19425,N_19346);
or U20163 (N_20163,N_19604,N_19878);
or U20164 (N_20164,N_19146,N_19060);
and U20165 (N_20165,N_19184,N_19183);
and U20166 (N_20166,N_19377,N_19607);
or U20167 (N_20167,N_19059,N_19169);
and U20168 (N_20168,N_19249,N_19213);
xnor U20169 (N_20169,N_19011,N_19917);
xor U20170 (N_20170,N_19396,N_19935);
xnor U20171 (N_20171,N_19954,N_19713);
and U20172 (N_20172,N_19153,N_19642);
nor U20173 (N_20173,N_19293,N_19232);
nand U20174 (N_20174,N_19477,N_19202);
nor U20175 (N_20175,N_19875,N_19594);
nand U20176 (N_20176,N_19631,N_19125);
nand U20177 (N_20177,N_19568,N_19434);
nor U20178 (N_20178,N_19140,N_19435);
nand U20179 (N_20179,N_19509,N_19096);
or U20180 (N_20180,N_19189,N_19689);
nand U20181 (N_20181,N_19273,N_19611);
or U20182 (N_20182,N_19522,N_19381);
nand U20183 (N_20183,N_19539,N_19963);
xnor U20184 (N_20184,N_19701,N_19039);
xnor U20185 (N_20185,N_19375,N_19196);
xor U20186 (N_20186,N_19026,N_19585);
and U20187 (N_20187,N_19521,N_19698);
xnor U20188 (N_20188,N_19717,N_19953);
nor U20189 (N_20189,N_19559,N_19959);
nor U20190 (N_20190,N_19210,N_19488);
or U20191 (N_20191,N_19337,N_19448);
or U20192 (N_20192,N_19471,N_19867);
nor U20193 (N_20193,N_19542,N_19845);
or U20194 (N_20194,N_19148,N_19768);
nor U20195 (N_20195,N_19599,N_19684);
nor U20196 (N_20196,N_19070,N_19736);
xor U20197 (N_20197,N_19500,N_19227);
xnor U20198 (N_20198,N_19349,N_19454);
xor U20199 (N_20199,N_19785,N_19807);
nand U20200 (N_20200,N_19474,N_19284);
nor U20201 (N_20201,N_19368,N_19422);
nand U20202 (N_20202,N_19045,N_19086);
nor U20203 (N_20203,N_19160,N_19181);
nand U20204 (N_20204,N_19397,N_19062);
or U20205 (N_20205,N_19074,N_19264);
nand U20206 (N_20206,N_19229,N_19550);
nand U20207 (N_20207,N_19393,N_19099);
nand U20208 (N_20208,N_19551,N_19465);
nand U20209 (N_20209,N_19428,N_19362);
nor U20210 (N_20210,N_19519,N_19246);
and U20211 (N_20211,N_19120,N_19490);
or U20212 (N_20212,N_19788,N_19103);
nand U20213 (N_20213,N_19411,N_19051);
or U20214 (N_20214,N_19825,N_19444);
or U20215 (N_20215,N_19638,N_19912);
or U20216 (N_20216,N_19609,N_19906);
nor U20217 (N_20217,N_19322,N_19679);
or U20218 (N_20218,N_19667,N_19406);
xnor U20219 (N_20219,N_19548,N_19042);
xor U20220 (N_20220,N_19656,N_19910);
or U20221 (N_20221,N_19961,N_19248);
or U20222 (N_20222,N_19415,N_19282);
nor U20223 (N_20223,N_19253,N_19053);
nor U20224 (N_20224,N_19979,N_19704);
xnor U20225 (N_20225,N_19009,N_19048);
xor U20226 (N_20226,N_19598,N_19777);
xor U20227 (N_20227,N_19044,N_19654);
or U20228 (N_20228,N_19892,N_19270);
nand U20229 (N_20229,N_19676,N_19541);
xor U20230 (N_20230,N_19265,N_19811);
and U20231 (N_20231,N_19345,N_19333);
nand U20232 (N_20232,N_19491,N_19316);
xnor U20233 (N_20233,N_19721,N_19473);
nor U20234 (N_20234,N_19573,N_19302);
xor U20235 (N_20235,N_19806,N_19288);
or U20236 (N_20236,N_19215,N_19023);
xnor U20237 (N_20237,N_19986,N_19741);
xnor U20238 (N_20238,N_19466,N_19219);
nor U20239 (N_20239,N_19583,N_19479);
nor U20240 (N_20240,N_19207,N_19495);
and U20241 (N_20241,N_19459,N_19379);
nor U20242 (N_20242,N_19993,N_19240);
nor U20243 (N_20243,N_19839,N_19300);
xor U20244 (N_20244,N_19409,N_19744);
xnor U20245 (N_20245,N_19814,N_19913);
nor U20246 (N_20246,N_19685,N_19565);
and U20247 (N_20247,N_19259,N_19171);
nor U20248 (N_20248,N_19299,N_19890);
nor U20249 (N_20249,N_19113,N_19405);
nand U20250 (N_20250,N_19668,N_19949);
nand U20251 (N_20251,N_19339,N_19782);
and U20252 (N_20252,N_19518,N_19193);
nand U20253 (N_20253,N_19476,N_19413);
nor U20254 (N_20254,N_19824,N_19767);
nor U20255 (N_20255,N_19478,N_19200);
nor U20256 (N_20256,N_19794,N_19669);
and U20257 (N_20257,N_19117,N_19197);
or U20258 (N_20258,N_19005,N_19534);
xnor U20259 (N_20259,N_19383,N_19132);
nor U20260 (N_20260,N_19908,N_19482);
and U20261 (N_20261,N_19971,N_19486);
nand U20262 (N_20262,N_19329,N_19016);
or U20263 (N_20263,N_19855,N_19063);
or U20264 (N_20264,N_19029,N_19228);
nor U20265 (N_20265,N_19111,N_19084);
and U20266 (N_20266,N_19703,N_19483);
nor U20267 (N_20267,N_19746,N_19886);
or U20268 (N_20268,N_19725,N_19245);
or U20269 (N_20269,N_19964,N_19008);
and U20270 (N_20270,N_19313,N_19818);
xnor U20271 (N_20271,N_19553,N_19324);
nand U20272 (N_20272,N_19105,N_19795);
xnor U20273 (N_20273,N_19615,N_19833);
and U20274 (N_20274,N_19523,N_19000);
xnor U20275 (N_20275,N_19305,N_19691);
nor U20276 (N_20276,N_19569,N_19546);
and U20277 (N_20277,N_19809,N_19644);
nand U20278 (N_20278,N_19538,N_19457);
and U20279 (N_20279,N_19330,N_19575);
nor U20280 (N_20280,N_19046,N_19561);
nand U20281 (N_20281,N_19544,N_19116);
nand U20282 (N_20282,N_19525,N_19664);
xor U20283 (N_20283,N_19040,N_19066);
and U20284 (N_20284,N_19975,N_19290);
nor U20285 (N_20285,N_19374,N_19918);
and U20286 (N_20286,N_19762,N_19937);
nand U20287 (N_20287,N_19941,N_19727);
nor U20288 (N_20288,N_19268,N_19505);
nand U20289 (N_20289,N_19690,N_19820);
xor U20290 (N_20290,N_19570,N_19827);
nor U20291 (N_20291,N_19384,N_19077);
xor U20292 (N_20292,N_19281,N_19608);
nand U20293 (N_20293,N_19267,N_19841);
xnor U20294 (N_20294,N_19951,N_19156);
and U20295 (N_20295,N_19317,N_19332);
and U20296 (N_20296,N_19810,N_19075);
and U20297 (N_20297,N_19982,N_19555);
or U20298 (N_20298,N_19447,N_19054);
or U20299 (N_20299,N_19738,N_19775);
nor U20300 (N_20300,N_19272,N_19663);
nor U20301 (N_20301,N_19496,N_19159);
nor U20302 (N_20302,N_19709,N_19056);
and U20303 (N_20303,N_19919,N_19277);
xor U20304 (N_20304,N_19526,N_19817);
or U20305 (N_20305,N_19545,N_19035);
nand U20306 (N_20306,N_19097,N_19280);
xnor U20307 (N_20307,N_19728,N_19101);
xnor U20308 (N_20308,N_19128,N_19834);
xnor U20309 (N_20309,N_19123,N_19931);
nor U20310 (N_20310,N_19695,N_19914);
or U20311 (N_20311,N_19168,N_19619);
nand U20312 (N_20312,N_19923,N_19453);
nor U20313 (N_20313,N_19187,N_19734);
and U20314 (N_20314,N_19772,N_19580);
nand U20315 (N_20315,N_19694,N_19266);
nor U20316 (N_20316,N_19643,N_19819);
xnor U20317 (N_20317,N_19314,N_19410);
nand U20318 (N_20318,N_19678,N_19632);
nand U20319 (N_20319,N_19722,N_19122);
nand U20320 (N_20320,N_19587,N_19370);
and U20321 (N_20321,N_19297,N_19968);
nand U20322 (N_20322,N_19347,N_19441);
nand U20323 (N_20323,N_19143,N_19921);
nor U20324 (N_20324,N_19188,N_19876);
and U20325 (N_20325,N_19517,N_19567);
and U20326 (N_20326,N_19222,N_19387);
nor U20327 (N_20327,N_19581,N_19376);
nor U20328 (N_20328,N_19236,N_19790);
nand U20329 (N_20329,N_19978,N_19212);
xor U20330 (N_20330,N_19380,N_19699);
and U20331 (N_20331,N_19271,N_19726);
nor U20332 (N_20332,N_19666,N_19540);
and U20333 (N_20333,N_19019,N_19802);
or U20334 (N_20334,N_19038,N_19732);
nand U20335 (N_20335,N_19192,N_19468);
xor U20336 (N_20336,N_19812,N_19967);
or U20337 (N_20337,N_19114,N_19956);
nand U20338 (N_20338,N_19584,N_19331);
and U20339 (N_20339,N_19276,N_19994);
xnor U20340 (N_20340,N_19871,N_19758);
nor U20341 (N_20341,N_19129,N_19998);
xor U20342 (N_20342,N_19311,N_19163);
nand U20343 (N_20343,N_19150,N_19504);
nor U20344 (N_20344,N_19618,N_19032);
xor U20345 (N_20345,N_19606,N_19939);
xnor U20346 (N_20346,N_19646,N_19999);
nor U20347 (N_20347,N_19793,N_19710);
and U20348 (N_20348,N_19729,N_19137);
or U20349 (N_20349,N_19624,N_19896);
or U20350 (N_20350,N_19733,N_19254);
nand U20351 (N_20351,N_19671,N_19628);
nor U20352 (N_20352,N_19104,N_19711);
nand U20353 (N_20353,N_19844,N_19731);
and U20354 (N_20354,N_19823,N_19692);
or U20355 (N_20355,N_19593,N_19167);
and U20356 (N_20356,N_19661,N_19022);
or U20357 (N_20357,N_19962,N_19372);
or U20358 (N_20358,N_19759,N_19506);
nor U20359 (N_20359,N_19177,N_19902);
or U20360 (N_20360,N_19862,N_19001);
nor U20361 (N_20361,N_19828,N_19821);
nand U20362 (N_20362,N_19589,N_19138);
nor U20363 (N_20363,N_19152,N_19831);
xor U20364 (N_20364,N_19217,N_19647);
nor U20365 (N_20365,N_19501,N_19328);
and U20366 (N_20366,N_19714,N_19043);
nand U20367 (N_20367,N_19781,N_19400);
xnor U20368 (N_20368,N_19900,N_19498);
and U20369 (N_20369,N_19614,N_19988);
and U20370 (N_20370,N_19361,N_19470);
and U20371 (N_20371,N_19981,N_19512);
and U20372 (N_20372,N_19499,N_19652);
nor U20373 (N_20373,N_19423,N_19298);
nor U20374 (N_20374,N_19865,N_19869);
xnor U20375 (N_20375,N_19050,N_19792);
nor U20376 (N_20376,N_19543,N_19560);
and U20377 (N_20377,N_19674,N_19625);
and U20378 (N_20378,N_19850,N_19024);
nor U20379 (N_20379,N_19243,N_19158);
xor U20380 (N_20380,N_19052,N_19848);
xnor U20381 (N_20381,N_19208,N_19004);
xnor U20382 (N_20382,N_19947,N_19737);
xnor U20383 (N_20383,N_19278,N_19973);
nand U20384 (N_20384,N_19366,N_19092);
and U20385 (N_20385,N_19972,N_19461);
nand U20386 (N_20386,N_19492,N_19417);
nand U20387 (N_20387,N_19629,N_19863);
and U20388 (N_20388,N_19983,N_19872);
nand U20389 (N_20389,N_19223,N_19633);
or U20390 (N_20390,N_19637,N_19275);
nand U20391 (N_20391,N_19338,N_19883);
or U20392 (N_20392,N_19460,N_19211);
nor U20393 (N_20393,N_19846,N_19752);
nor U20394 (N_20394,N_19119,N_19318);
nand U20395 (N_20395,N_19635,N_19749);
or U20396 (N_20396,N_19320,N_19980);
or U20397 (N_20397,N_19144,N_19194);
and U20398 (N_20398,N_19630,N_19739);
or U20399 (N_20399,N_19100,N_19149);
or U20400 (N_20400,N_19238,N_19933);
nand U20401 (N_20401,N_19291,N_19651);
and U20402 (N_20402,N_19067,N_19590);
xnor U20403 (N_20403,N_19308,N_19724);
nand U20404 (N_20404,N_19613,N_19446);
nor U20405 (N_20405,N_19451,N_19235);
nand U20406 (N_20406,N_19088,N_19201);
xor U20407 (N_20407,N_19151,N_19090);
xnor U20408 (N_20408,N_19650,N_19880);
xnor U20409 (N_20409,N_19705,N_19481);
and U20410 (N_20410,N_19352,N_19155);
nand U20411 (N_20411,N_19162,N_19094);
xnor U20412 (N_20412,N_19110,N_19443);
and U20413 (N_20413,N_19344,N_19894);
nor U20414 (N_20414,N_19258,N_19206);
or U20415 (N_20415,N_19359,N_19852);
and U20416 (N_20416,N_19392,N_19449);
nor U20417 (N_20417,N_19966,N_19898);
xor U20418 (N_20418,N_19303,N_19174);
or U20419 (N_20419,N_19866,N_19757);
and U20420 (N_20420,N_19142,N_19269);
xor U20421 (N_20421,N_19577,N_19464);
nand U20422 (N_20422,N_19027,N_19712);
and U20423 (N_20423,N_19389,N_19603);
nand U20424 (N_20424,N_19926,N_19533);
xnor U20425 (N_20425,N_19552,N_19353);
and U20426 (N_20426,N_19870,N_19783);
nor U20427 (N_20427,N_19126,N_19879);
xnor U20428 (N_20428,N_19687,N_19950);
nand U20429 (N_20429,N_19475,N_19532);
nor U20430 (N_20430,N_19891,N_19385);
or U20431 (N_20431,N_19085,N_19970);
and U20432 (N_20432,N_19720,N_19424);
xnor U20433 (N_20433,N_19511,N_19688);
xor U20434 (N_20434,N_19131,N_19797);
and U20435 (N_20435,N_19838,N_19185);
and U20436 (N_20436,N_19677,N_19796);
xor U20437 (N_20437,N_19659,N_19250);
nor U20438 (N_20438,N_19530,N_19860);
nand U20439 (N_20439,N_19938,N_19002);
xnor U20440 (N_20440,N_19778,N_19456);
xnor U20441 (N_20441,N_19127,N_19107);
nand U20442 (N_20442,N_19612,N_19922);
or U20443 (N_20443,N_19412,N_19136);
and U20444 (N_20444,N_19445,N_19723);
nand U20445 (N_20445,N_19895,N_19433);
nand U20446 (N_20446,N_19920,N_19766);
nand U20447 (N_20447,N_19014,N_19247);
and U20448 (N_20448,N_19675,N_19083);
or U20449 (N_20449,N_19829,N_19761);
nand U20450 (N_20450,N_19033,N_19779);
nand U20451 (N_20451,N_19170,N_19442);
and U20452 (N_20452,N_19467,N_19657);
or U20453 (N_20453,N_19925,N_19610);
or U20454 (N_20454,N_19493,N_19754);
xor U20455 (N_20455,N_19976,N_19431);
nand U20456 (N_20456,N_19414,N_19231);
nor U20457 (N_20457,N_19990,N_19716);
and U20458 (N_20458,N_19429,N_19597);
or U20459 (N_20459,N_19462,N_19524);
nor U20460 (N_20460,N_19108,N_19244);
or U20461 (N_20461,N_19702,N_19289);
and U20462 (N_20462,N_19884,N_19252);
nor U20463 (N_20463,N_19472,N_19556);
nor U20464 (N_20464,N_19622,N_19209);
or U20465 (N_20465,N_19803,N_19756);
xor U20466 (N_20466,N_19178,N_19098);
or U20467 (N_20467,N_19835,N_19386);
nand U20468 (N_20468,N_19851,N_19021);
or U20469 (N_20469,N_19360,N_19507);
or U20470 (N_20470,N_19536,N_19673);
xor U20471 (N_20471,N_19403,N_19164);
nand U20472 (N_20472,N_19715,N_19853);
xnor U20473 (N_20473,N_19292,N_19987);
nor U20474 (N_20474,N_19091,N_19093);
nand U20475 (N_20475,N_19363,N_19682);
and U20476 (N_20476,N_19003,N_19943);
nand U20477 (N_20477,N_19653,N_19750);
nand U20478 (N_20478,N_19571,N_19740);
nor U20479 (N_20479,N_19241,N_19776);
or U20480 (N_20480,N_19995,N_19064);
nand U20481 (N_20481,N_19996,N_19899);
and U20482 (N_20482,N_19342,N_19421);
nand U20483 (N_20483,N_19049,N_19582);
xor U20484 (N_20484,N_19800,N_19944);
or U20485 (N_20485,N_19887,N_19989);
nor U20486 (N_20486,N_19382,N_19686);
xnor U20487 (N_20487,N_19854,N_19437);
xor U20488 (N_20488,N_19007,N_19992);
or U20489 (N_20489,N_19969,N_19082);
or U20490 (N_20490,N_19747,N_19861);
or U20491 (N_20491,N_19165,N_19182);
nand U20492 (N_20492,N_19364,N_19487);
and U20493 (N_20493,N_19190,N_19830);
xor U20494 (N_20494,N_19513,N_19294);
xor U20495 (N_20495,N_19124,N_19658);
nor U20496 (N_20496,N_19929,N_19670);
nand U20497 (N_20497,N_19799,N_19399);
xnor U20498 (N_20498,N_19816,N_19903);
xnor U20499 (N_20499,N_19822,N_19578);
or U20500 (N_20500,N_19748,N_19322);
xor U20501 (N_20501,N_19973,N_19038);
and U20502 (N_20502,N_19095,N_19049);
nor U20503 (N_20503,N_19456,N_19561);
or U20504 (N_20504,N_19782,N_19045);
and U20505 (N_20505,N_19707,N_19990);
and U20506 (N_20506,N_19740,N_19879);
or U20507 (N_20507,N_19718,N_19830);
xor U20508 (N_20508,N_19866,N_19783);
or U20509 (N_20509,N_19533,N_19471);
nand U20510 (N_20510,N_19070,N_19023);
and U20511 (N_20511,N_19251,N_19265);
and U20512 (N_20512,N_19483,N_19415);
nand U20513 (N_20513,N_19779,N_19145);
nor U20514 (N_20514,N_19334,N_19346);
nor U20515 (N_20515,N_19777,N_19402);
and U20516 (N_20516,N_19331,N_19005);
nand U20517 (N_20517,N_19545,N_19688);
nor U20518 (N_20518,N_19589,N_19414);
nor U20519 (N_20519,N_19340,N_19271);
xor U20520 (N_20520,N_19928,N_19502);
or U20521 (N_20521,N_19052,N_19417);
nand U20522 (N_20522,N_19521,N_19639);
nor U20523 (N_20523,N_19501,N_19084);
and U20524 (N_20524,N_19799,N_19902);
and U20525 (N_20525,N_19921,N_19965);
or U20526 (N_20526,N_19023,N_19512);
and U20527 (N_20527,N_19611,N_19099);
nor U20528 (N_20528,N_19885,N_19976);
and U20529 (N_20529,N_19071,N_19646);
xor U20530 (N_20530,N_19556,N_19617);
xnor U20531 (N_20531,N_19488,N_19555);
nor U20532 (N_20532,N_19816,N_19561);
and U20533 (N_20533,N_19336,N_19659);
nor U20534 (N_20534,N_19821,N_19811);
nand U20535 (N_20535,N_19582,N_19023);
nand U20536 (N_20536,N_19985,N_19721);
xor U20537 (N_20537,N_19915,N_19005);
xor U20538 (N_20538,N_19472,N_19167);
nand U20539 (N_20539,N_19497,N_19660);
xnor U20540 (N_20540,N_19990,N_19646);
nand U20541 (N_20541,N_19861,N_19893);
nand U20542 (N_20542,N_19777,N_19754);
and U20543 (N_20543,N_19624,N_19937);
xor U20544 (N_20544,N_19994,N_19262);
and U20545 (N_20545,N_19785,N_19134);
xnor U20546 (N_20546,N_19967,N_19424);
and U20547 (N_20547,N_19754,N_19522);
or U20548 (N_20548,N_19991,N_19123);
nand U20549 (N_20549,N_19131,N_19120);
nor U20550 (N_20550,N_19798,N_19320);
nor U20551 (N_20551,N_19287,N_19575);
nor U20552 (N_20552,N_19745,N_19520);
nand U20553 (N_20553,N_19277,N_19708);
nand U20554 (N_20554,N_19197,N_19650);
nor U20555 (N_20555,N_19396,N_19340);
nand U20556 (N_20556,N_19297,N_19623);
nor U20557 (N_20557,N_19853,N_19031);
nand U20558 (N_20558,N_19618,N_19139);
and U20559 (N_20559,N_19749,N_19762);
xnor U20560 (N_20560,N_19718,N_19139);
or U20561 (N_20561,N_19327,N_19577);
and U20562 (N_20562,N_19745,N_19815);
and U20563 (N_20563,N_19850,N_19193);
nor U20564 (N_20564,N_19420,N_19028);
nand U20565 (N_20565,N_19198,N_19074);
and U20566 (N_20566,N_19455,N_19365);
xnor U20567 (N_20567,N_19778,N_19069);
nand U20568 (N_20568,N_19610,N_19064);
xor U20569 (N_20569,N_19408,N_19409);
xor U20570 (N_20570,N_19673,N_19710);
and U20571 (N_20571,N_19120,N_19521);
xnor U20572 (N_20572,N_19890,N_19691);
nand U20573 (N_20573,N_19781,N_19156);
or U20574 (N_20574,N_19847,N_19256);
and U20575 (N_20575,N_19945,N_19070);
xor U20576 (N_20576,N_19779,N_19502);
and U20577 (N_20577,N_19922,N_19546);
nand U20578 (N_20578,N_19778,N_19184);
xnor U20579 (N_20579,N_19019,N_19796);
nand U20580 (N_20580,N_19127,N_19145);
or U20581 (N_20581,N_19101,N_19534);
nand U20582 (N_20582,N_19009,N_19229);
xor U20583 (N_20583,N_19745,N_19510);
nand U20584 (N_20584,N_19768,N_19156);
nor U20585 (N_20585,N_19856,N_19910);
or U20586 (N_20586,N_19633,N_19018);
or U20587 (N_20587,N_19243,N_19909);
nand U20588 (N_20588,N_19572,N_19974);
xor U20589 (N_20589,N_19776,N_19910);
nand U20590 (N_20590,N_19456,N_19679);
and U20591 (N_20591,N_19526,N_19599);
xor U20592 (N_20592,N_19119,N_19910);
nand U20593 (N_20593,N_19345,N_19656);
nor U20594 (N_20594,N_19578,N_19837);
or U20595 (N_20595,N_19598,N_19805);
and U20596 (N_20596,N_19560,N_19899);
xnor U20597 (N_20597,N_19981,N_19807);
and U20598 (N_20598,N_19825,N_19169);
nand U20599 (N_20599,N_19043,N_19798);
nand U20600 (N_20600,N_19397,N_19028);
and U20601 (N_20601,N_19388,N_19060);
nor U20602 (N_20602,N_19138,N_19687);
or U20603 (N_20603,N_19005,N_19581);
or U20604 (N_20604,N_19058,N_19855);
nand U20605 (N_20605,N_19790,N_19598);
xor U20606 (N_20606,N_19298,N_19073);
or U20607 (N_20607,N_19017,N_19805);
xnor U20608 (N_20608,N_19168,N_19342);
xnor U20609 (N_20609,N_19901,N_19327);
or U20610 (N_20610,N_19822,N_19207);
or U20611 (N_20611,N_19430,N_19992);
nand U20612 (N_20612,N_19889,N_19600);
or U20613 (N_20613,N_19504,N_19780);
nand U20614 (N_20614,N_19149,N_19821);
or U20615 (N_20615,N_19648,N_19960);
xor U20616 (N_20616,N_19958,N_19456);
or U20617 (N_20617,N_19182,N_19057);
and U20618 (N_20618,N_19889,N_19505);
nand U20619 (N_20619,N_19507,N_19198);
xor U20620 (N_20620,N_19325,N_19659);
nor U20621 (N_20621,N_19117,N_19243);
nand U20622 (N_20622,N_19644,N_19597);
nand U20623 (N_20623,N_19496,N_19032);
nor U20624 (N_20624,N_19689,N_19072);
or U20625 (N_20625,N_19060,N_19881);
nand U20626 (N_20626,N_19470,N_19379);
or U20627 (N_20627,N_19771,N_19954);
or U20628 (N_20628,N_19063,N_19042);
xor U20629 (N_20629,N_19713,N_19556);
and U20630 (N_20630,N_19487,N_19305);
nor U20631 (N_20631,N_19214,N_19625);
nor U20632 (N_20632,N_19898,N_19835);
xor U20633 (N_20633,N_19848,N_19016);
xor U20634 (N_20634,N_19265,N_19232);
and U20635 (N_20635,N_19787,N_19100);
or U20636 (N_20636,N_19017,N_19528);
nor U20637 (N_20637,N_19735,N_19988);
and U20638 (N_20638,N_19663,N_19070);
nand U20639 (N_20639,N_19767,N_19319);
nor U20640 (N_20640,N_19299,N_19003);
xnor U20641 (N_20641,N_19661,N_19197);
and U20642 (N_20642,N_19535,N_19636);
and U20643 (N_20643,N_19255,N_19554);
nor U20644 (N_20644,N_19230,N_19140);
and U20645 (N_20645,N_19845,N_19427);
nor U20646 (N_20646,N_19727,N_19804);
nor U20647 (N_20647,N_19578,N_19697);
or U20648 (N_20648,N_19801,N_19674);
and U20649 (N_20649,N_19769,N_19379);
xor U20650 (N_20650,N_19270,N_19931);
and U20651 (N_20651,N_19452,N_19467);
nand U20652 (N_20652,N_19923,N_19287);
xnor U20653 (N_20653,N_19462,N_19320);
xor U20654 (N_20654,N_19200,N_19898);
or U20655 (N_20655,N_19110,N_19109);
or U20656 (N_20656,N_19585,N_19450);
nand U20657 (N_20657,N_19527,N_19135);
nor U20658 (N_20658,N_19354,N_19669);
and U20659 (N_20659,N_19544,N_19826);
and U20660 (N_20660,N_19549,N_19722);
and U20661 (N_20661,N_19803,N_19162);
or U20662 (N_20662,N_19945,N_19881);
nand U20663 (N_20663,N_19443,N_19402);
nand U20664 (N_20664,N_19721,N_19451);
xor U20665 (N_20665,N_19957,N_19467);
nor U20666 (N_20666,N_19094,N_19185);
or U20667 (N_20667,N_19982,N_19318);
nor U20668 (N_20668,N_19136,N_19069);
nor U20669 (N_20669,N_19812,N_19188);
xor U20670 (N_20670,N_19665,N_19608);
xor U20671 (N_20671,N_19470,N_19133);
nand U20672 (N_20672,N_19715,N_19500);
or U20673 (N_20673,N_19053,N_19658);
and U20674 (N_20674,N_19069,N_19427);
or U20675 (N_20675,N_19080,N_19599);
and U20676 (N_20676,N_19144,N_19140);
or U20677 (N_20677,N_19478,N_19170);
or U20678 (N_20678,N_19804,N_19216);
or U20679 (N_20679,N_19176,N_19459);
and U20680 (N_20680,N_19589,N_19846);
xor U20681 (N_20681,N_19889,N_19652);
xor U20682 (N_20682,N_19823,N_19050);
and U20683 (N_20683,N_19027,N_19487);
or U20684 (N_20684,N_19203,N_19127);
nor U20685 (N_20685,N_19723,N_19066);
and U20686 (N_20686,N_19760,N_19320);
and U20687 (N_20687,N_19126,N_19026);
or U20688 (N_20688,N_19973,N_19369);
or U20689 (N_20689,N_19755,N_19920);
xnor U20690 (N_20690,N_19125,N_19092);
nor U20691 (N_20691,N_19530,N_19735);
or U20692 (N_20692,N_19969,N_19908);
nor U20693 (N_20693,N_19958,N_19438);
and U20694 (N_20694,N_19556,N_19772);
and U20695 (N_20695,N_19075,N_19067);
and U20696 (N_20696,N_19498,N_19500);
xor U20697 (N_20697,N_19209,N_19716);
and U20698 (N_20698,N_19728,N_19920);
and U20699 (N_20699,N_19267,N_19757);
and U20700 (N_20700,N_19722,N_19470);
xor U20701 (N_20701,N_19714,N_19515);
or U20702 (N_20702,N_19983,N_19417);
xor U20703 (N_20703,N_19516,N_19199);
and U20704 (N_20704,N_19439,N_19465);
and U20705 (N_20705,N_19175,N_19136);
xnor U20706 (N_20706,N_19992,N_19517);
nand U20707 (N_20707,N_19286,N_19291);
xor U20708 (N_20708,N_19160,N_19220);
and U20709 (N_20709,N_19471,N_19479);
and U20710 (N_20710,N_19931,N_19987);
nor U20711 (N_20711,N_19240,N_19569);
nand U20712 (N_20712,N_19305,N_19455);
xor U20713 (N_20713,N_19458,N_19942);
nor U20714 (N_20714,N_19189,N_19997);
or U20715 (N_20715,N_19823,N_19088);
nand U20716 (N_20716,N_19272,N_19530);
nand U20717 (N_20717,N_19683,N_19329);
or U20718 (N_20718,N_19373,N_19324);
or U20719 (N_20719,N_19316,N_19430);
or U20720 (N_20720,N_19676,N_19545);
or U20721 (N_20721,N_19307,N_19718);
or U20722 (N_20722,N_19637,N_19630);
xor U20723 (N_20723,N_19899,N_19014);
xnor U20724 (N_20724,N_19733,N_19120);
xor U20725 (N_20725,N_19198,N_19012);
nor U20726 (N_20726,N_19956,N_19659);
xnor U20727 (N_20727,N_19016,N_19022);
xnor U20728 (N_20728,N_19980,N_19029);
nor U20729 (N_20729,N_19167,N_19247);
nand U20730 (N_20730,N_19676,N_19804);
nand U20731 (N_20731,N_19173,N_19036);
and U20732 (N_20732,N_19085,N_19045);
nand U20733 (N_20733,N_19261,N_19472);
nor U20734 (N_20734,N_19753,N_19584);
nand U20735 (N_20735,N_19949,N_19815);
xnor U20736 (N_20736,N_19908,N_19216);
xnor U20737 (N_20737,N_19643,N_19457);
nor U20738 (N_20738,N_19418,N_19976);
nand U20739 (N_20739,N_19674,N_19142);
xor U20740 (N_20740,N_19308,N_19269);
xor U20741 (N_20741,N_19178,N_19390);
or U20742 (N_20742,N_19506,N_19656);
and U20743 (N_20743,N_19203,N_19884);
nor U20744 (N_20744,N_19604,N_19957);
and U20745 (N_20745,N_19652,N_19916);
xor U20746 (N_20746,N_19579,N_19675);
and U20747 (N_20747,N_19865,N_19768);
or U20748 (N_20748,N_19044,N_19525);
nand U20749 (N_20749,N_19101,N_19647);
nand U20750 (N_20750,N_19698,N_19195);
or U20751 (N_20751,N_19479,N_19896);
or U20752 (N_20752,N_19965,N_19430);
and U20753 (N_20753,N_19147,N_19113);
nor U20754 (N_20754,N_19923,N_19252);
and U20755 (N_20755,N_19840,N_19056);
nor U20756 (N_20756,N_19521,N_19601);
xor U20757 (N_20757,N_19069,N_19602);
xnor U20758 (N_20758,N_19560,N_19167);
and U20759 (N_20759,N_19574,N_19557);
and U20760 (N_20760,N_19716,N_19473);
nand U20761 (N_20761,N_19548,N_19077);
and U20762 (N_20762,N_19411,N_19255);
or U20763 (N_20763,N_19857,N_19278);
or U20764 (N_20764,N_19771,N_19171);
nor U20765 (N_20765,N_19910,N_19182);
or U20766 (N_20766,N_19476,N_19451);
xnor U20767 (N_20767,N_19102,N_19663);
and U20768 (N_20768,N_19821,N_19564);
nor U20769 (N_20769,N_19170,N_19381);
or U20770 (N_20770,N_19354,N_19380);
and U20771 (N_20771,N_19408,N_19706);
nor U20772 (N_20772,N_19022,N_19624);
xnor U20773 (N_20773,N_19227,N_19375);
nor U20774 (N_20774,N_19262,N_19443);
xor U20775 (N_20775,N_19125,N_19702);
or U20776 (N_20776,N_19937,N_19161);
or U20777 (N_20777,N_19876,N_19956);
nand U20778 (N_20778,N_19847,N_19781);
and U20779 (N_20779,N_19291,N_19599);
and U20780 (N_20780,N_19825,N_19348);
nor U20781 (N_20781,N_19570,N_19417);
and U20782 (N_20782,N_19449,N_19078);
and U20783 (N_20783,N_19468,N_19962);
nor U20784 (N_20784,N_19640,N_19866);
nor U20785 (N_20785,N_19833,N_19267);
nand U20786 (N_20786,N_19736,N_19261);
and U20787 (N_20787,N_19944,N_19336);
xnor U20788 (N_20788,N_19480,N_19326);
nor U20789 (N_20789,N_19521,N_19197);
nor U20790 (N_20790,N_19509,N_19831);
nor U20791 (N_20791,N_19167,N_19036);
xnor U20792 (N_20792,N_19812,N_19899);
nand U20793 (N_20793,N_19353,N_19942);
xnor U20794 (N_20794,N_19010,N_19302);
nor U20795 (N_20795,N_19093,N_19156);
nand U20796 (N_20796,N_19360,N_19461);
xor U20797 (N_20797,N_19748,N_19613);
nor U20798 (N_20798,N_19055,N_19281);
or U20799 (N_20799,N_19547,N_19740);
nand U20800 (N_20800,N_19724,N_19409);
or U20801 (N_20801,N_19762,N_19320);
nand U20802 (N_20802,N_19306,N_19009);
xnor U20803 (N_20803,N_19734,N_19213);
or U20804 (N_20804,N_19701,N_19242);
or U20805 (N_20805,N_19917,N_19649);
nand U20806 (N_20806,N_19628,N_19698);
or U20807 (N_20807,N_19619,N_19173);
nand U20808 (N_20808,N_19757,N_19005);
nand U20809 (N_20809,N_19344,N_19898);
or U20810 (N_20810,N_19584,N_19133);
nor U20811 (N_20811,N_19124,N_19378);
nor U20812 (N_20812,N_19843,N_19654);
or U20813 (N_20813,N_19982,N_19894);
nor U20814 (N_20814,N_19154,N_19981);
or U20815 (N_20815,N_19722,N_19217);
and U20816 (N_20816,N_19597,N_19091);
or U20817 (N_20817,N_19165,N_19973);
nand U20818 (N_20818,N_19548,N_19732);
nand U20819 (N_20819,N_19669,N_19097);
and U20820 (N_20820,N_19361,N_19520);
or U20821 (N_20821,N_19529,N_19047);
nand U20822 (N_20822,N_19591,N_19175);
or U20823 (N_20823,N_19733,N_19923);
xor U20824 (N_20824,N_19745,N_19499);
xor U20825 (N_20825,N_19801,N_19248);
nor U20826 (N_20826,N_19117,N_19529);
or U20827 (N_20827,N_19010,N_19921);
nand U20828 (N_20828,N_19717,N_19628);
nand U20829 (N_20829,N_19916,N_19928);
nand U20830 (N_20830,N_19004,N_19169);
xor U20831 (N_20831,N_19456,N_19739);
xnor U20832 (N_20832,N_19040,N_19300);
nor U20833 (N_20833,N_19415,N_19361);
nand U20834 (N_20834,N_19403,N_19917);
nand U20835 (N_20835,N_19887,N_19630);
and U20836 (N_20836,N_19505,N_19148);
nor U20837 (N_20837,N_19293,N_19239);
xor U20838 (N_20838,N_19360,N_19353);
nor U20839 (N_20839,N_19898,N_19373);
or U20840 (N_20840,N_19746,N_19380);
xnor U20841 (N_20841,N_19939,N_19995);
and U20842 (N_20842,N_19847,N_19945);
xnor U20843 (N_20843,N_19340,N_19504);
nand U20844 (N_20844,N_19046,N_19222);
nor U20845 (N_20845,N_19961,N_19291);
and U20846 (N_20846,N_19664,N_19371);
nor U20847 (N_20847,N_19461,N_19722);
and U20848 (N_20848,N_19674,N_19930);
nand U20849 (N_20849,N_19379,N_19306);
and U20850 (N_20850,N_19090,N_19392);
or U20851 (N_20851,N_19162,N_19079);
nor U20852 (N_20852,N_19333,N_19150);
or U20853 (N_20853,N_19482,N_19441);
and U20854 (N_20854,N_19912,N_19960);
and U20855 (N_20855,N_19302,N_19091);
xnor U20856 (N_20856,N_19031,N_19326);
and U20857 (N_20857,N_19779,N_19528);
or U20858 (N_20858,N_19926,N_19939);
nor U20859 (N_20859,N_19550,N_19670);
nand U20860 (N_20860,N_19124,N_19697);
or U20861 (N_20861,N_19839,N_19679);
or U20862 (N_20862,N_19224,N_19998);
or U20863 (N_20863,N_19598,N_19422);
nand U20864 (N_20864,N_19775,N_19732);
nor U20865 (N_20865,N_19808,N_19358);
nand U20866 (N_20866,N_19559,N_19508);
or U20867 (N_20867,N_19260,N_19032);
nand U20868 (N_20868,N_19572,N_19598);
and U20869 (N_20869,N_19568,N_19320);
nand U20870 (N_20870,N_19934,N_19075);
xnor U20871 (N_20871,N_19362,N_19866);
nor U20872 (N_20872,N_19673,N_19270);
nand U20873 (N_20873,N_19113,N_19510);
nor U20874 (N_20874,N_19451,N_19326);
nand U20875 (N_20875,N_19730,N_19054);
nor U20876 (N_20876,N_19664,N_19162);
or U20877 (N_20877,N_19114,N_19458);
or U20878 (N_20878,N_19883,N_19471);
nand U20879 (N_20879,N_19024,N_19481);
nand U20880 (N_20880,N_19182,N_19072);
nand U20881 (N_20881,N_19615,N_19332);
xor U20882 (N_20882,N_19480,N_19100);
nor U20883 (N_20883,N_19070,N_19404);
xnor U20884 (N_20884,N_19115,N_19830);
or U20885 (N_20885,N_19676,N_19666);
xor U20886 (N_20886,N_19106,N_19444);
xor U20887 (N_20887,N_19523,N_19721);
or U20888 (N_20888,N_19567,N_19383);
nor U20889 (N_20889,N_19893,N_19948);
nor U20890 (N_20890,N_19811,N_19613);
and U20891 (N_20891,N_19850,N_19746);
nor U20892 (N_20892,N_19671,N_19561);
nor U20893 (N_20893,N_19386,N_19075);
xor U20894 (N_20894,N_19401,N_19348);
or U20895 (N_20895,N_19722,N_19206);
xnor U20896 (N_20896,N_19703,N_19383);
and U20897 (N_20897,N_19343,N_19930);
and U20898 (N_20898,N_19101,N_19191);
or U20899 (N_20899,N_19320,N_19933);
and U20900 (N_20900,N_19939,N_19618);
nand U20901 (N_20901,N_19269,N_19608);
nor U20902 (N_20902,N_19502,N_19633);
xnor U20903 (N_20903,N_19674,N_19693);
nor U20904 (N_20904,N_19378,N_19826);
xnor U20905 (N_20905,N_19804,N_19737);
or U20906 (N_20906,N_19024,N_19713);
nor U20907 (N_20907,N_19139,N_19487);
or U20908 (N_20908,N_19361,N_19228);
xor U20909 (N_20909,N_19339,N_19269);
or U20910 (N_20910,N_19563,N_19615);
nor U20911 (N_20911,N_19290,N_19898);
nand U20912 (N_20912,N_19182,N_19343);
xor U20913 (N_20913,N_19966,N_19183);
or U20914 (N_20914,N_19122,N_19137);
or U20915 (N_20915,N_19482,N_19120);
nand U20916 (N_20916,N_19300,N_19881);
or U20917 (N_20917,N_19089,N_19026);
and U20918 (N_20918,N_19741,N_19569);
or U20919 (N_20919,N_19008,N_19796);
nand U20920 (N_20920,N_19671,N_19459);
xor U20921 (N_20921,N_19074,N_19975);
xor U20922 (N_20922,N_19747,N_19369);
nor U20923 (N_20923,N_19678,N_19259);
xor U20924 (N_20924,N_19430,N_19822);
xor U20925 (N_20925,N_19466,N_19690);
nor U20926 (N_20926,N_19709,N_19114);
nor U20927 (N_20927,N_19114,N_19500);
nand U20928 (N_20928,N_19161,N_19479);
or U20929 (N_20929,N_19469,N_19951);
nor U20930 (N_20930,N_19461,N_19347);
and U20931 (N_20931,N_19602,N_19814);
nand U20932 (N_20932,N_19703,N_19900);
and U20933 (N_20933,N_19347,N_19629);
xnor U20934 (N_20934,N_19159,N_19674);
or U20935 (N_20935,N_19819,N_19394);
xor U20936 (N_20936,N_19758,N_19570);
xnor U20937 (N_20937,N_19080,N_19512);
or U20938 (N_20938,N_19877,N_19519);
nor U20939 (N_20939,N_19024,N_19251);
nand U20940 (N_20940,N_19401,N_19949);
nand U20941 (N_20941,N_19143,N_19829);
or U20942 (N_20942,N_19743,N_19265);
and U20943 (N_20943,N_19846,N_19194);
and U20944 (N_20944,N_19059,N_19282);
and U20945 (N_20945,N_19266,N_19135);
and U20946 (N_20946,N_19773,N_19448);
or U20947 (N_20947,N_19985,N_19844);
xor U20948 (N_20948,N_19015,N_19326);
or U20949 (N_20949,N_19056,N_19278);
xor U20950 (N_20950,N_19524,N_19048);
xor U20951 (N_20951,N_19994,N_19596);
xor U20952 (N_20952,N_19106,N_19648);
xor U20953 (N_20953,N_19393,N_19791);
xnor U20954 (N_20954,N_19409,N_19044);
nor U20955 (N_20955,N_19516,N_19545);
nand U20956 (N_20956,N_19127,N_19522);
nor U20957 (N_20957,N_19618,N_19347);
or U20958 (N_20958,N_19300,N_19550);
or U20959 (N_20959,N_19391,N_19551);
nand U20960 (N_20960,N_19997,N_19854);
nand U20961 (N_20961,N_19665,N_19208);
nor U20962 (N_20962,N_19879,N_19502);
xnor U20963 (N_20963,N_19103,N_19738);
or U20964 (N_20964,N_19375,N_19022);
xor U20965 (N_20965,N_19018,N_19704);
nor U20966 (N_20966,N_19803,N_19222);
nor U20967 (N_20967,N_19510,N_19800);
xor U20968 (N_20968,N_19773,N_19830);
or U20969 (N_20969,N_19787,N_19939);
nor U20970 (N_20970,N_19708,N_19745);
nor U20971 (N_20971,N_19668,N_19166);
xnor U20972 (N_20972,N_19659,N_19136);
nand U20973 (N_20973,N_19646,N_19438);
or U20974 (N_20974,N_19146,N_19291);
nor U20975 (N_20975,N_19837,N_19796);
or U20976 (N_20976,N_19724,N_19141);
nor U20977 (N_20977,N_19530,N_19763);
and U20978 (N_20978,N_19303,N_19568);
nor U20979 (N_20979,N_19003,N_19133);
xnor U20980 (N_20980,N_19024,N_19712);
xnor U20981 (N_20981,N_19600,N_19065);
nand U20982 (N_20982,N_19000,N_19153);
nand U20983 (N_20983,N_19359,N_19102);
nand U20984 (N_20984,N_19586,N_19495);
and U20985 (N_20985,N_19254,N_19230);
or U20986 (N_20986,N_19096,N_19391);
xor U20987 (N_20987,N_19749,N_19616);
and U20988 (N_20988,N_19261,N_19220);
and U20989 (N_20989,N_19338,N_19417);
xor U20990 (N_20990,N_19500,N_19097);
nor U20991 (N_20991,N_19863,N_19393);
and U20992 (N_20992,N_19067,N_19773);
nor U20993 (N_20993,N_19572,N_19400);
nor U20994 (N_20994,N_19150,N_19852);
xnor U20995 (N_20995,N_19711,N_19889);
or U20996 (N_20996,N_19419,N_19616);
or U20997 (N_20997,N_19166,N_19314);
or U20998 (N_20998,N_19412,N_19941);
or U20999 (N_20999,N_19221,N_19442);
nand U21000 (N_21000,N_20974,N_20804);
nand U21001 (N_21001,N_20894,N_20347);
nand U21002 (N_21002,N_20095,N_20741);
nand U21003 (N_21003,N_20350,N_20850);
xnor U21004 (N_21004,N_20591,N_20487);
and U21005 (N_21005,N_20059,N_20885);
xor U21006 (N_21006,N_20392,N_20361);
xnor U21007 (N_21007,N_20299,N_20342);
nor U21008 (N_21008,N_20809,N_20817);
or U21009 (N_21009,N_20865,N_20620);
nand U21010 (N_21010,N_20933,N_20616);
and U21011 (N_21011,N_20096,N_20152);
and U21012 (N_21012,N_20601,N_20054);
xnor U21013 (N_21013,N_20679,N_20495);
or U21014 (N_21014,N_20563,N_20805);
and U21015 (N_21015,N_20860,N_20825);
or U21016 (N_21016,N_20357,N_20795);
xor U21017 (N_21017,N_20755,N_20611);
xnor U21018 (N_21018,N_20346,N_20649);
xor U21019 (N_21019,N_20390,N_20067);
xor U21020 (N_21020,N_20039,N_20723);
nand U21021 (N_21021,N_20635,N_20003);
or U21022 (N_21022,N_20638,N_20617);
nand U21023 (N_21023,N_20289,N_20184);
and U21024 (N_21024,N_20085,N_20694);
xnor U21025 (N_21025,N_20566,N_20125);
nor U21026 (N_21026,N_20109,N_20661);
nor U21027 (N_21027,N_20472,N_20092);
xnor U21028 (N_21028,N_20235,N_20510);
nand U21029 (N_21029,N_20997,N_20921);
nor U21030 (N_21030,N_20735,N_20791);
nor U21031 (N_21031,N_20405,N_20943);
and U21032 (N_21032,N_20721,N_20416);
nor U21033 (N_21033,N_20223,N_20808);
nand U21034 (N_21034,N_20952,N_20046);
nand U21035 (N_21035,N_20946,N_20282);
xor U21036 (N_21036,N_20882,N_20516);
xnor U21037 (N_21037,N_20760,N_20722);
xor U21038 (N_21038,N_20315,N_20270);
or U21039 (N_21039,N_20983,N_20904);
and U21040 (N_21040,N_20877,N_20603);
nor U21041 (N_21041,N_20041,N_20292);
xor U21042 (N_21042,N_20957,N_20806);
xor U21043 (N_21043,N_20160,N_20395);
and U21044 (N_21044,N_20064,N_20954);
or U21045 (N_21045,N_20536,N_20589);
xnor U21046 (N_21046,N_20705,N_20582);
and U21047 (N_21047,N_20686,N_20696);
and U21048 (N_21048,N_20440,N_20774);
or U21049 (N_21049,N_20720,N_20577);
or U21050 (N_21050,N_20258,N_20460);
nand U21051 (N_21051,N_20366,N_20135);
and U21052 (N_21052,N_20733,N_20984);
xnor U21053 (N_21053,N_20204,N_20783);
nor U21054 (N_21054,N_20917,N_20869);
xnor U21055 (N_21055,N_20622,N_20306);
nor U21056 (N_21056,N_20431,N_20560);
and U21057 (N_21057,N_20150,N_20540);
nor U21058 (N_21058,N_20961,N_20463);
xor U21059 (N_21059,N_20173,N_20631);
or U21060 (N_21060,N_20993,N_20290);
or U21061 (N_21061,N_20305,N_20313);
xor U21062 (N_21062,N_20280,N_20139);
and U21063 (N_21063,N_20834,N_20861);
nor U21064 (N_21064,N_20457,N_20134);
nand U21065 (N_21065,N_20147,N_20000);
nor U21066 (N_21066,N_20811,N_20537);
nor U21067 (N_21067,N_20142,N_20105);
and U21068 (N_21068,N_20345,N_20216);
and U21069 (N_21069,N_20454,N_20391);
nor U21070 (N_21070,N_20363,N_20272);
and U21071 (N_21071,N_20891,N_20940);
nor U21072 (N_21072,N_20951,N_20787);
and U21073 (N_21073,N_20883,N_20788);
nand U21074 (N_21074,N_20969,N_20584);
nor U21075 (N_21075,N_20596,N_20724);
xor U21076 (N_21076,N_20193,N_20473);
nor U21077 (N_21077,N_20364,N_20254);
xnor U21078 (N_21078,N_20352,N_20925);
nand U21079 (N_21079,N_20482,N_20518);
nand U21080 (N_21080,N_20101,N_20852);
nor U21081 (N_21081,N_20751,N_20358);
or U21082 (N_21082,N_20338,N_20077);
and U21083 (N_21083,N_20670,N_20878);
or U21084 (N_21084,N_20903,N_20653);
nor U21085 (N_21085,N_20428,N_20727);
nor U21086 (N_21086,N_20148,N_20189);
and U21087 (N_21087,N_20467,N_20091);
nor U21088 (N_21088,N_20221,N_20958);
or U21089 (N_21089,N_20180,N_20115);
xor U21090 (N_21090,N_20975,N_20005);
xor U21091 (N_21091,N_20406,N_20375);
nand U21092 (N_21092,N_20317,N_20422);
nor U21093 (N_21093,N_20504,N_20864);
nor U21094 (N_21094,N_20523,N_20511);
and U21095 (N_21095,N_20234,N_20253);
and U21096 (N_21096,N_20455,N_20063);
nor U21097 (N_21097,N_20826,N_20625);
nand U21098 (N_21098,N_20792,N_20771);
xnor U21099 (N_21099,N_20822,N_20075);
and U21100 (N_21100,N_20201,N_20621);
nor U21101 (N_21101,N_20079,N_20332);
nand U21102 (N_21102,N_20987,N_20161);
nand U21103 (N_21103,N_20785,N_20409);
and U21104 (N_21104,N_20146,N_20190);
xnor U21105 (N_21105,N_20572,N_20778);
xor U21106 (N_21106,N_20669,N_20384);
nor U21107 (N_21107,N_20261,N_20848);
nand U21108 (N_21108,N_20242,N_20123);
xnor U21109 (N_21109,N_20245,N_20595);
nor U21110 (N_21110,N_20074,N_20310);
or U21111 (N_21111,N_20509,N_20598);
or U21112 (N_21112,N_20828,N_20541);
nand U21113 (N_21113,N_20944,N_20704);
and U21114 (N_21114,N_20938,N_20592);
xnor U21115 (N_21115,N_20931,N_20586);
or U21116 (N_21116,N_20934,N_20047);
nor U21117 (N_21117,N_20073,N_20643);
and U21118 (N_21118,N_20626,N_20296);
or U21119 (N_21119,N_20329,N_20301);
xnor U21120 (N_21120,N_20320,N_20985);
or U21121 (N_21121,N_20965,N_20402);
xnor U21122 (N_21122,N_20374,N_20408);
or U21123 (N_21123,N_20496,N_20866);
xnor U21124 (N_21124,N_20027,N_20237);
xnor U21125 (N_21125,N_20627,N_20907);
xnor U21126 (N_21126,N_20750,N_20080);
and U21127 (N_21127,N_20973,N_20756);
xor U21128 (N_21128,N_20939,N_20702);
nor U21129 (N_21129,N_20126,N_20924);
nand U21130 (N_21130,N_20343,N_20008);
xor U21131 (N_21131,N_20248,N_20667);
xnor U21132 (N_21132,N_20775,N_20252);
and U21133 (N_21133,N_20102,N_20609);
nor U21134 (N_21134,N_20137,N_20200);
nand U21135 (N_21135,N_20437,N_20158);
nor U21136 (N_21136,N_20539,N_20976);
and U21137 (N_21137,N_20922,N_20094);
xnor U21138 (N_21138,N_20247,N_20678);
nor U21139 (N_21139,N_20240,N_20874);
or U21140 (N_21140,N_20881,N_20876);
nor U21141 (N_21141,N_20713,N_20155);
xor U21142 (N_21142,N_20862,N_20226);
nor U21143 (N_21143,N_20071,N_20318);
xnor U21144 (N_21144,N_20545,N_20830);
nand U21145 (N_21145,N_20297,N_20766);
xnor U21146 (N_21146,N_20819,N_20335);
nand U21147 (N_21147,N_20624,N_20024);
nand U21148 (N_21148,N_20082,N_20477);
xor U21149 (N_21149,N_20549,N_20485);
nand U21150 (N_21150,N_20948,N_20979);
and U21151 (N_21151,N_20859,N_20312);
and U21152 (N_21152,N_20311,N_20831);
and U21153 (N_21153,N_20953,N_20476);
nor U21154 (N_21154,N_20023,N_20418);
and U21155 (N_21155,N_20232,N_20475);
nand U21156 (N_21156,N_20793,N_20215);
nand U21157 (N_21157,N_20585,N_20579);
and U21158 (N_21158,N_20164,N_20530);
or U21159 (N_21159,N_20548,N_20857);
or U21160 (N_21160,N_20326,N_20786);
nand U21161 (N_21161,N_20656,N_20949);
or U21162 (N_21162,N_20749,N_20355);
nor U21163 (N_21163,N_20773,N_20174);
or U21164 (N_21164,N_20411,N_20647);
nor U21165 (N_21165,N_20991,N_20553);
nor U21166 (N_21166,N_20493,N_20203);
nand U21167 (N_21167,N_20729,N_20764);
nor U21168 (N_21168,N_20491,N_20657);
nor U21169 (N_21169,N_20707,N_20435);
nor U21170 (N_21170,N_20634,N_20262);
nand U21171 (N_21171,N_20370,N_20502);
nor U21172 (N_21172,N_20980,N_20651);
or U21173 (N_21173,N_20021,N_20851);
nor U21174 (N_21174,N_20165,N_20373);
and U21175 (N_21175,N_20765,N_20978);
nand U21176 (N_21176,N_20654,N_20918);
nand U21177 (N_21177,N_20644,N_20344);
nand U21178 (N_21178,N_20913,N_20932);
nand U21179 (N_21179,N_20562,N_20334);
and U21180 (N_21180,N_20176,N_20810);
xnor U21181 (N_21181,N_20479,N_20763);
xor U21182 (N_21182,N_20996,N_20725);
xnor U21183 (N_21183,N_20557,N_20167);
or U21184 (N_21184,N_20281,N_20593);
nor U21185 (N_21185,N_20693,N_20145);
nor U21186 (N_21186,N_20019,N_20381);
nand U21187 (N_21187,N_20841,N_20697);
xor U21188 (N_21188,N_20858,N_20849);
or U21189 (N_21189,N_20121,N_20066);
nand U21190 (N_21190,N_20149,N_20369);
and U21191 (N_21191,N_20856,N_20982);
nor U21192 (N_21192,N_20959,N_20923);
nor U21193 (N_21193,N_20905,N_20847);
nand U21194 (N_21194,N_20124,N_20655);
xnor U21195 (N_21195,N_20535,N_20829);
and U21196 (N_21196,N_20664,N_20555);
and U21197 (N_21197,N_20561,N_20719);
nand U21198 (N_21198,N_20612,N_20279);
xnor U21199 (N_21199,N_20056,N_20739);
nor U21200 (N_21200,N_20640,N_20425);
xor U21201 (N_21201,N_20525,N_20336);
nand U21202 (N_21202,N_20351,N_20010);
nor U21203 (N_21203,N_20183,N_20772);
nand U21204 (N_21204,N_20845,N_20886);
or U21205 (N_21205,N_20710,N_20768);
nand U21206 (N_21206,N_20945,N_20941);
nor U21207 (N_21207,N_20287,N_20636);
xor U21208 (N_21208,N_20439,N_20004);
nor U21209 (N_21209,N_20701,N_20218);
nor U21210 (N_21210,N_20875,N_20659);
xnor U21211 (N_21211,N_20711,N_20341);
nor U21212 (N_21212,N_20759,N_20846);
or U21213 (N_21213,N_20687,N_20058);
and U21214 (N_21214,N_20567,N_20323);
and U21215 (N_21215,N_20276,N_20111);
nor U21216 (N_21216,N_20520,N_20744);
and U21217 (N_21217,N_20259,N_20187);
and U21218 (N_21218,N_20674,N_20210);
or U21219 (N_21219,N_20527,N_20738);
nor U21220 (N_21220,N_20127,N_20412);
or U21221 (N_21221,N_20057,N_20802);
and U21222 (N_21222,N_20544,N_20515);
xor U21223 (N_21223,N_20602,N_20823);
nand U21224 (N_21224,N_20001,N_20486);
and U21225 (N_21225,N_20209,N_20090);
nor U21226 (N_21226,N_20295,N_20492);
or U21227 (N_21227,N_20742,N_20269);
nand U21228 (N_21228,N_20110,N_20257);
xor U21229 (N_21229,N_20188,N_20256);
and U21230 (N_21230,N_20162,N_20020);
or U21231 (N_21231,N_20587,N_20225);
and U21232 (N_21232,N_20947,N_20178);
xnor U21233 (N_21233,N_20608,N_20214);
xnor U21234 (N_21234,N_20445,N_20359);
and U21235 (N_21235,N_20995,N_20424);
nor U21236 (N_21236,N_20571,N_20196);
and U21237 (N_21237,N_20337,N_20827);
nor U21238 (N_21238,N_20458,N_20488);
and U21239 (N_21239,N_20497,N_20340);
and U21240 (N_21240,N_20716,N_20103);
nand U21241 (N_21241,N_20227,N_20906);
nand U21242 (N_21242,N_20330,N_20868);
xnor U21243 (N_21243,N_20112,N_20508);
xnor U21244 (N_21244,N_20100,N_20641);
nor U21245 (N_21245,N_20628,N_20506);
nor U21246 (N_21246,N_20842,N_20192);
xor U21247 (N_21247,N_20789,N_20986);
nor U21248 (N_21248,N_20503,N_20926);
xor U21249 (N_21249,N_20231,N_20388);
nand U21250 (N_21250,N_20185,N_20025);
nand U21251 (N_21251,N_20060,N_20360);
nand U21252 (N_21252,N_20229,N_20581);
nand U21253 (N_21253,N_20144,N_20767);
nor U21254 (N_21254,N_20154,N_20393);
nand U21255 (N_21255,N_20353,N_20519);
or U21256 (N_21256,N_20747,N_20444);
nor U21257 (N_21257,N_20386,N_20762);
and U21258 (N_21258,N_20662,N_20438);
nand U21259 (N_21259,N_20618,N_20998);
nand U21260 (N_21260,N_20956,N_20568);
nand U21261 (N_21261,N_20385,N_20513);
nor U21262 (N_21262,N_20052,N_20665);
nand U21263 (N_21263,N_20758,N_20228);
nand U21264 (N_21264,N_20970,N_20578);
nor U21265 (N_21265,N_20043,N_20029);
nor U21266 (N_21266,N_20050,N_20119);
nand U21267 (N_21267,N_20166,N_20597);
and U21268 (N_21268,N_20712,N_20106);
or U21269 (N_21269,N_20820,N_20576);
or U21270 (N_21270,N_20013,N_20348);
and U21271 (N_21271,N_20499,N_20081);
xnor U21272 (N_21272,N_20677,N_20920);
xnor U21273 (N_21273,N_20784,N_20919);
nor U21274 (N_21274,N_20465,N_20401);
nor U21275 (N_21275,N_20547,N_20414);
or U21276 (N_21276,N_20239,N_20500);
nand U21277 (N_21277,N_20265,N_20888);
and U21278 (N_21278,N_20302,N_20069);
xnor U21279 (N_21279,N_20378,N_20753);
nand U21280 (N_21280,N_20930,N_20610);
and U21281 (N_21281,N_20818,N_20521);
nand U21282 (N_21282,N_20117,N_20870);
xnor U21283 (N_21283,N_20086,N_20331);
and U21284 (N_21284,N_20794,N_20843);
xnor U21285 (N_21285,N_20615,N_20538);
or U21286 (N_21286,N_20404,N_20380);
xor U21287 (N_21287,N_20377,N_20140);
or U21288 (N_21288,N_20936,N_20650);
nand U21289 (N_21289,N_20098,N_20286);
nand U21290 (N_21290,N_20898,N_20087);
nor U21291 (N_21291,N_20706,N_20676);
or U21292 (N_21292,N_20994,N_20456);
and U21293 (N_21293,N_20078,N_20717);
nand U21294 (N_21294,N_20093,N_20194);
nand U21295 (N_21295,N_20195,N_20394);
xor U21296 (N_21296,N_20570,N_20604);
nand U21297 (N_21297,N_20423,N_20588);
or U21298 (N_21298,N_20104,N_20799);
nor U21299 (N_21299,N_20319,N_20011);
xnor U21300 (N_21300,N_20051,N_20143);
or U21301 (N_21301,N_20867,N_20880);
nor U21302 (N_21302,N_20040,N_20339);
xor U21303 (N_21303,N_20042,N_20734);
and U21304 (N_21304,N_20715,N_20614);
nor U21305 (N_21305,N_20977,N_20186);
or U21306 (N_21306,N_20895,N_20400);
xnor U21307 (N_21307,N_20448,N_20594);
xor U21308 (N_21308,N_20430,N_20322);
nand U21309 (N_21309,N_20801,N_20512);
or U21310 (N_21310,N_20800,N_20267);
nand U21311 (N_21311,N_20709,N_20745);
nor U21312 (N_21312,N_20084,N_20999);
xnor U21313 (N_21313,N_20835,N_20700);
or U21314 (N_21314,N_20033,N_20646);
xnor U21315 (N_21315,N_20559,N_20007);
xnor U21316 (N_21316,N_20893,N_20083);
xor U21317 (N_21317,N_20045,N_20554);
or U21318 (N_21318,N_20156,N_20372);
or U21319 (N_21319,N_20573,N_20220);
xor U21320 (N_21320,N_20892,N_20446);
nand U21321 (N_21321,N_20450,N_20871);
xnor U21322 (N_21322,N_20410,N_20207);
nor U21323 (N_21323,N_20447,N_20376);
nor U21324 (N_21324,N_20197,N_20908);
xor U21325 (N_21325,N_20246,N_20489);
nand U21326 (N_21326,N_20972,N_20097);
xor U21327 (N_21327,N_20403,N_20449);
nand U21328 (N_21328,N_20839,N_20556);
or U21329 (N_21329,N_20838,N_20927);
and U21330 (N_21330,N_20855,N_20451);
nor U21331 (N_21331,N_20249,N_20478);
and U21332 (N_21332,N_20757,N_20122);
or U21333 (N_21333,N_20470,N_20328);
nand U21334 (N_21334,N_20288,N_20990);
and U21335 (N_21335,N_20798,N_20837);
xnor U21336 (N_21336,N_20955,N_20580);
and U21337 (N_21337,N_20396,N_20133);
and U21338 (N_21338,N_20964,N_20191);
nand U21339 (N_21339,N_20528,N_20629);
or U21340 (N_21340,N_20534,N_20268);
and U21341 (N_21341,N_20217,N_20796);
and U21342 (N_21342,N_20006,N_20522);
xor U21343 (N_21343,N_20642,N_20550);
xnor U21344 (N_21344,N_20623,N_20663);
nor U21345 (N_21345,N_20212,N_20175);
xnor U21346 (N_21346,N_20131,N_20298);
and U21347 (N_21347,N_20872,N_20089);
nor U21348 (N_21348,N_20433,N_20365);
and U21349 (N_21349,N_20637,N_20718);
nand U21350 (N_21350,N_20264,N_20469);
nor U21351 (N_21351,N_20132,N_20675);
nor U21352 (N_21352,N_20420,N_20543);
nand U21353 (N_21353,N_20362,N_20030);
or U21354 (N_21354,N_20053,N_20206);
xnor U21355 (N_21355,N_20790,N_20630);
and U21356 (N_21356,N_20285,N_20699);
xnor U21357 (N_21357,N_20929,N_20564);
or U21358 (N_21358,N_20153,N_20708);
and U21359 (N_21359,N_20230,N_20896);
nor U21360 (N_21360,N_20014,N_20915);
xnor U21361 (N_21361,N_20278,N_20263);
xnor U21362 (N_21362,N_20068,N_20912);
nor U21363 (N_21363,N_20607,N_20099);
nand U21364 (N_21364,N_20483,N_20517);
and U21365 (N_21365,N_20909,N_20208);
nand U21366 (N_21366,N_20732,N_20224);
and U21367 (N_21367,N_20498,N_20038);
nor U21368 (N_21368,N_20356,N_20419);
and U21369 (N_21369,N_20128,N_20873);
and U21370 (N_21370,N_20325,N_20900);
nor U21371 (N_21371,N_20442,N_20389);
nand U21372 (N_21372,N_20379,N_20044);
or U21373 (N_21373,N_20432,N_20172);
nand U21374 (N_21374,N_20514,N_20816);
nor U21375 (N_21375,N_20928,N_20692);
xor U21376 (N_21376,N_20836,N_20303);
or U21377 (N_21377,N_20606,N_20202);
nor U21378 (N_21378,N_20022,N_20480);
and U21379 (N_21379,N_20076,N_20685);
and U21380 (N_21380,N_20660,N_20182);
and U21381 (N_21381,N_20695,N_20854);
xnor U21382 (N_21382,N_20652,N_20474);
xor U21383 (N_21383,N_20832,N_20383);
or U21384 (N_21384,N_20284,N_20690);
nor U21385 (N_21385,N_20777,N_20429);
nand U21386 (N_21386,N_20501,N_20198);
or U21387 (N_21387,N_20294,N_20782);
or U21388 (N_21388,N_20966,N_20118);
nand U21389 (N_21389,N_20464,N_20672);
and U21390 (N_21390,N_20552,N_20012);
nor U21391 (N_21391,N_20494,N_20397);
nand U21392 (N_21392,N_20989,N_20507);
nand U21393 (N_21393,N_20813,N_20682);
xor U21394 (N_21394,N_20002,N_20009);
and U21395 (N_21395,N_20436,N_20531);
nor U21396 (N_21396,N_20599,N_20236);
xor U21397 (N_21397,N_20901,N_20035);
xnor U21398 (N_21398,N_20426,N_20466);
and U21399 (N_21399,N_20277,N_20018);
nor U21400 (N_21400,N_20300,N_20316);
nor U21401 (N_21401,N_20484,N_20413);
xor U21402 (N_21402,N_20911,N_20714);
xnor U21403 (N_21403,N_20211,N_20748);
and U21404 (N_21404,N_20960,N_20417);
or U21405 (N_21405,N_20179,N_20461);
xor U21406 (N_21406,N_20910,N_20114);
nand U21407 (N_21407,N_20291,N_20890);
nand U21408 (N_21408,N_20671,N_20304);
nor U21409 (N_21409,N_20314,N_20251);
and U21410 (N_21410,N_20899,N_20736);
or U21411 (N_21411,N_20031,N_20061);
nor U21412 (N_21412,N_20250,N_20243);
and U21413 (N_21413,N_20434,N_20666);
or U21414 (N_21414,N_20307,N_20524);
nand U21415 (N_21415,N_20367,N_20689);
nor U21416 (N_21416,N_20797,N_20387);
and U21417 (N_21417,N_20632,N_20681);
xnor U21418 (N_21418,N_20684,N_20897);
or U21419 (N_21419,N_20971,N_20781);
or U21420 (N_21420,N_20407,N_20824);
nand U21421 (N_21421,N_20807,N_20551);
nand U21422 (N_21422,N_20780,N_20726);
nand U21423 (N_21423,N_20163,N_20935);
or U21424 (N_21424,N_20988,N_20222);
xnor U21425 (N_21425,N_20273,N_20761);
xnor U21426 (N_21426,N_20600,N_20181);
or U21427 (N_21427,N_20275,N_20481);
nand U21428 (N_21428,N_20968,N_20565);
or U21429 (N_21429,N_20130,N_20072);
xnor U21430 (N_21430,N_20271,N_20399);
and U21431 (N_21431,N_20887,N_20138);
xnor U21432 (N_21432,N_20583,N_20532);
or U21433 (N_21433,N_20136,N_20737);
nand U21434 (N_21434,N_20668,N_20613);
or U21435 (N_21435,N_20113,N_20863);
or U21436 (N_21436,N_20680,N_20177);
nand U21437 (N_21437,N_20371,N_20884);
xor U21438 (N_21438,N_20526,N_20992);
nor U21439 (N_21439,N_20441,N_20814);
xor U21440 (N_21440,N_20575,N_20648);
xnor U21441 (N_21441,N_20219,N_20468);
nand U21442 (N_21442,N_20633,N_20879);
or U21443 (N_21443,N_20116,N_20574);
xor U21444 (N_21444,N_20017,N_20619);
and U21445 (N_21445,N_20398,N_20168);
or U21446 (N_21446,N_20037,N_20902);
nand U21447 (N_21447,N_20108,N_20205);
or U21448 (N_21448,N_20238,N_20151);
xnor U21449 (N_21449,N_20505,N_20776);
xor U21450 (N_21450,N_20016,N_20062);
and U21451 (N_21451,N_20382,N_20889);
and U21452 (N_21452,N_20321,N_20769);
nor U21453 (N_21453,N_20260,N_20740);
and U21454 (N_21454,N_20213,N_20703);
xor U21455 (N_21455,N_20821,N_20658);
nor U21456 (N_21456,N_20490,N_20754);
and U21457 (N_21457,N_20569,N_20840);
xnor U21458 (N_21458,N_20274,N_20026);
nor U21459 (N_21459,N_20055,N_20645);
nor U21460 (N_21460,N_20255,N_20354);
or U21461 (N_21461,N_20770,N_20942);
nand U21462 (N_21462,N_20833,N_20752);
xor U21463 (N_21463,N_20981,N_20065);
nor U21464 (N_21464,N_20803,N_20032);
and U21465 (N_21465,N_20452,N_20471);
xor U21466 (N_21466,N_20036,N_20728);
and U21467 (N_21467,N_20293,N_20333);
xnor U21468 (N_21468,N_20558,N_20107);
nand U21469 (N_21469,N_20639,N_20327);
xor U21470 (N_21470,N_20048,N_20368);
and U21471 (N_21471,N_20141,N_20241);
or U21472 (N_21472,N_20746,N_20171);
xnor U21473 (N_21473,N_20590,N_20731);
xnor U21474 (N_21474,N_20421,N_20673);
and U21475 (N_21475,N_20967,N_20199);
xor U21476 (N_21476,N_20844,N_20815);
xor U21477 (N_21477,N_20743,N_20533);
or U21478 (N_21478,N_20170,N_20415);
nor U21479 (N_21479,N_20914,N_20812);
nand U21480 (N_21480,N_20049,N_20962);
xor U21481 (N_21481,N_20129,N_20088);
xor U21482 (N_21482,N_20542,N_20427);
nand U21483 (N_21483,N_20309,N_20698);
xnor U21484 (N_21484,N_20546,N_20683);
nand U21485 (N_21485,N_20034,N_20459);
or U21486 (N_21486,N_20916,N_20159);
and U21487 (N_21487,N_20937,N_20244);
nand U21488 (N_21488,N_20233,N_20730);
nand U21489 (N_21489,N_20070,N_20605);
xor U21490 (N_21490,N_20453,N_20169);
nor U21491 (N_21491,N_20462,N_20324);
xnor U21492 (N_21492,N_20853,N_20028);
or U21493 (N_21493,N_20688,N_20308);
nor U21494 (N_21494,N_20283,N_20529);
nor U21495 (N_21495,N_20120,N_20157);
xor U21496 (N_21496,N_20963,N_20779);
and U21497 (N_21497,N_20349,N_20443);
nand U21498 (N_21498,N_20015,N_20266);
and U21499 (N_21499,N_20691,N_20950);
nor U21500 (N_21500,N_20171,N_20559);
xnor U21501 (N_21501,N_20637,N_20925);
and U21502 (N_21502,N_20159,N_20824);
xor U21503 (N_21503,N_20915,N_20867);
nand U21504 (N_21504,N_20149,N_20446);
nand U21505 (N_21505,N_20700,N_20563);
nand U21506 (N_21506,N_20718,N_20183);
nor U21507 (N_21507,N_20452,N_20389);
or U21508 (N_21508,N_20588,N_20132);
nor U21509 (N_21509,N_20955,N_20311);
xor U21510 (N_21510,N_20117,N_20248);
xor U21511 (N_21511,N_20656,N_20902);
nor U21512 (N_21512,N_20174,N_20220);
nand U21513 (N_21513,N_20235,N_20491);
xnor U21514 (N_21514,N_20344,N_20970);
nand U21515 (N_21515,N_20500,N_20232);
nor U21516 (N_21516,N_20478,N_20967);
and U21517 (N_21517,N_20141,N_20550);
and U21518 (N_21518,N_20548,N_20530);
and U21519 (N_21519,N_20097,N_20553);
nand U21520 (N_21520,N_20961,N_20154);
xnor U21521 (N_21521,N_20795,N_20131);
nor U21522 (N_21522,N_20585,N_20664);
or U21523 (N_21523,N_20992,N_20569);
and U21524 (N_21524,N_20607,N_20008);
nor U21525 (N_21525,N_20950,N_20280);
xor U21526 (N_21526,N_20501,N_20296);
xor U21527 (N_21527,N_20520,N_20271);
nor U21528 (N_21528,N_20088,N_20501);
or U21529 (N_21529,N_20572,N_20275);
or U21530 (N_21530,N_20071,N_20864);
or U21531 (N_21531,N_20752,N_20309);
or U21532 (N_21532,N_20987,N_20070);
and U21533 (N_21533,N_20801,N_20999);
nor U21534 (N_21534,N_20441,N_20434);
nor U21535 (N_21535,N_20552,N_20942);
nand U21536 (N_21536,N_20923,N_20571);
xnor U21537 (N_21537,N_20837,N_20723);
and U21538 (N_21538,N_20698,N_20404);
xnor U21539 (N_21539,N_20703,N_20756);
nor U21540 (N_21540,N_20698,N_20657);
nor U21541 (N_21541,N_20175,N_20094);
or U21542 (N_21542,N_20421,N_20274);
and U21543 (N_21543,N_20254,N_20023);
or U21544 (N_21544,N_20904,N_20245);
nor U21545 (N_21545,N_20128,N_20855);
nor U21546 (N_21546,N_20959,N_20265);
nor U21547 (N_21547,N_20166,N_20210);
nand U21548 (N_21548,N_20456,N_20138);
xor U21549 (N_21549,N_20657,N_20433);
nand U21550 (N_21550,N_20583,N_20920);
or U21551 (N_21551,N_20429,N_20138);
and U21552 (N_21552,N_20298,N_20563);
nor U21553 (N_21553,N_20667,N_20183);
or U21554 (N_21554,N_20147,N_20103);
xor U21555 (N_21555,N_20152,N_20939);
nand U21556 (N_21556,N_20197,N_20575);
xor U21557 (N_21557,N_20534,N_20842);
and U21558 (N_21558,N_20870,N_20473);
and U21559 (N_21559,N_20155,N_20656);
nand U21560 (N_21560,N_20778,N_20239);
and U21561 (N_21561,N_20448,N_20472);
nand U21562 (N_21562,N_20347,N_20293);
nor U21563 (N_21563,N_20780,N_20596);
xnor U21564 (N_21564,N_20971,N_20380);
or U21565 (N_21565,N_20082,N_20777);
or U21566 (N_21566,N_20926,N_20629);
nand U21567 (N_21567,N_20856,N_20592);
xor U21568 (N_21568,N_20871,N_20547);
nand U21569 (N_21569,N_20766,N_20575);
or U21570 (N_21570,N_20077,N_20874);
nor U21571 (N_21571,N_20859,N_20180);
nand U21572 (N_21572,N_20381,N_20803);
and U21573 (N_21573,N_20396,N_20467);
or U21574 (N_21574,N_20730,N_20956);
xnor U21575 (N_21575,N_20997,N_20798);
nor U21576 (N_21576,N_20381,N_20192);
nor U21577 (N_21577,N_20158,N_20885);
or U21578 (N_21578,N_20663,N_20472);
or U21579 (N_21579,N_20456,N_20363);
and U21580 (N_21580,N_20812,N_20527);
xnor U21581 (N_21581,N_20153,N_20166);
nor U21582 (N_21582,N_20665,N_20912);
or U21583 (N_21583,N_20884,N_20082);
and U21584 (N_21584,N_20946,N_20176);
nand U21585 (N_21585,N_20341,N_20253);
and U21586 (N_21586,N_20629,N_20631);
and U21587 (N_21587,N_20791,N_20691);
xor U21588 (N_21588,N_20193,N_20031);
and U21589 (N_21589,N_20606,N_20500);
or U21590 (N_21590,N_20265,N_20994);
nor U21591 (N_21591,N_20728,N_20784);
nor U21592 (N_21592,N_20871,N_20663);
or U21593 (N_21593,N_20919,N_20559);
xnor U21594 (N_21594,N_20325,N_20320);
nor U21595 (N_21595,N_20964,N_20224);
xnor U21596 (N_21596,N_20835,N_20207);
xor U21597 (N_21597,N_20991,N_20399);
and U21598 (N_21598,N_20470,N_20267);
or U21599 (N_21599,N_20361,N_20405);
nand U21600 (N_21600,N_20736,N_20471);
nor U21601 (N_21601,N_20764,N_20498);
and U21602 (N_21602,N_20383,N_20528);
and U21603 (N_21603,N_20532,N_20544);
nand U21604 (N_21604,N_20133,N_20420);
nor U21605 (N_21605,N_20647,N_20505);
nand U21606 (N_21606,N_20302,N_20681);
or U21607 (N_21607,N_20557,N_20700);
nor U21608 (N_21608,N_20969,N_20820);
and U21609 (N_21609,N_20054,N_20844);
and U21610 (N_21610,N_20586,N_20263);
or U21611 (N_21611,N_20830,N_20858);
nor U21612 (N_21612,N_20656,N_20201);
nor U21613 (N_21613,N_20472,N_20209);
or U21614 (N_21614,N_20995,N_20251);
and U21615 (N_21615,N_20403,N_20727);
or U21616 (N_21616,N_20528,N_20396);
nand U21617 (N_21617,N_20711,N_20839);
nand U21618 (N_21618,N_20910,N_20715);
or U21619 (N_21619,N_20314,N_20416);
or U21620 (N_21620,N_20041,N_20727);
and U21621 (N_21621,N_20276,N_20869);
xor U21622 (N_21622,N_20953,N_20356);
nor U21623 (N_21623,N_20724,N_20677);
and U21624 (N_21624,N_20134,N_20220);
nand U21625 (N_21625,N_20490,N_20134);
nand U21626 (N_21626,N_20754,N_20175);
xnor U21627 (N_21627,N_20251,N_20802);
xor U21628 (N_21628,N_20037,N_20438);
or U21629 (N_21629,N_20177,N_20874);
xor U21630 (N_21630,N_20278,N_20452);
or U21631 (N_21631,N_20400,N_20781);
or U21632 (N_21632,N_20223,N_20290);
xor U21633 (N_21633,N_20366,N_20597);
nand U21634 (N_21634,N_20249,N_20863);
or U21635 (N_21635,N_20768,N_20973);
nand U21636 (N_21636,N_20725,N_20339);
nand U21637 (N_21637,N_20132,N_20643);
nand U21638 (N_21638,N_20861,N_20039);
nand U21639 (N_21639,N_20298,N_20759);
xor U21640 (N_21640,N_20142,N_20221);
and U21641 (N_21641,N_20745,N_20725);
or U21642 (N_21642,N_20924,N_20379);
xor U21643 (N_21643,N_20357,N_20859);
xnor U21644 (N_21644,N_20932,N_20431);
or U21645 (N_21645,N_20823,N_20859);
or U21646 (N_21646,N_20677,N_20941);
or U21647 (N_21647,N_20796,N_20525);
nor U21648 (N_21648,N_20155,N_20935);
nand U21649 (N_21649,N_20704,N_20728);
xor U21650 (N_21650,N_20036,N_20100);
or U21651 (N_21651,N_20682,N_20842);
xor U21652 (N_21652,N_20114,N_20421);
xor U21653 (N_21653,N_20222,N_20984);
nor U21654 (N_21654,N_20729,N_20573);
nor U21655 (N_21655,N_20823,N_20215);
and U21656 (N_21656,N_20760,N_20314);
nor U21657 (N_21657,N_20092,N_20062);
and U21658 (N_21658,N_20007,N_20129);
nor U21659 (N_21659,N_20352,N_20897);
nand U21660 (N_21660,N_20463,N_20785);
nand U21661 (N_21661,N_20363,N_20704);
xor U21662 (N_21662,N_20298,N_20541);
nand U21663 (N_21663,N_20833,N_20616);
or U21664 (N_21664,N_20569,N_20400);
nor U21665 (N_21665,N_20036,N_20019);
nand U21666 (N_21666,N_20318,N_20070);
or U21667 (N_21667,N_20103,N_20267);
nor U21668 (N_21668,N_20311,N_20932);
and U21669 (N_21669,N_20523,N_20252);
xnor U21670 (N_21670,N_20706,N_20854);
xnor U21671 (N_21671,N_20696,N_20357);
nand U21672 (N_21672,N_20203,N_20658);
xor U21673 (N_21673,N_20524,N_20182);
xnor U21674 (N_21674,N_20948,N_20689);
nand U21675 (N_21675,N_20943,N_20689);
nor U21676 (N_21676,N_20009,N_20805);
or U21677 (N_21677,N_20908,N_20346);
nand U21678 (N_21678,N_20458,N_20257);
and U21679 (N_21679,N_20170,N_20391);
and U21680 (N_21680,N_20890,N_20761);
nand U21681 (N_21681,N_20811,N_20612);
or U21682 (N_21682,N_20743,N_20804);
nor U21683 (N_21683,N_20928,N_20349);
nor U21684 (N_21684,N_20116,N_20162);
nand U21685 (N_21685,N_20151,N_20879);
nand U21686 (N_21686,N_20785,N_20437);
xor U21687 (N_21687,N_20603,N_20912);
xnor U21688 (N_21688,N_20600,N_20954);
nor U21689 (N_21689,N_20792,N_20244);
nand U21690 (N_21690,N_20992,N_20962);
or U21691 (N_21691,N_20820,N_20510);
nor U21692 (N_21692,N_20412,N_20792);
and U21693 (N_21693,N_20244,N_20381);
xnor U21694 (N_21694,N_20687,N_20432);
nand U21695 (N_21695,N_20088,N_20873);
or U21696 (N_21696,N_20232,N_20413);
nand U21697 (N_21697,N_20203,N_20339);
and U21698 (N_21698,N_20323,N_20103);
nand U21699 (N_21699,N_20653,N_20649);
xor U21700 (N_21700,N_20005,N_20192);
and U21701 (N_21701,N_20389,N_20675);
nor U21702 (N_21702,N_20735,N_20124);
or U21703 (N_21703,N_20724,N_20178);
or U21704 (N_21704,N_20723,N_20690);
nor U21705 (N_21705,N_20025,N_20537);
xor U21706 (N_21706,N_20465,N_20617);
and U21707 (N_21707,N_20393,N_20573);
and U21708 (N_21708,N_20479,N_20847);
and U21709 (N_21709,N_20094,N_20845);
nand U21710 (N_21710,N_20823,N_20656);
nor U21711 (N_21711,N_20789,N_20661);
nor U21712 (N_21712,N_20604,N_20252);
xnor U21713 (N_21713,N_20022,N_20355);
or U21714 (N_21714,N_20146,N_20417);
xnor U21715 (N_21715,N_20122,N_20147);
nor U21716 (N_21716,N_20547,N_20241);
and U21717 (N_21717,N_20589,N_20229);
and U21718 (N_21718,N_20097,N_20049);
or U21719 (N_21719,N_20323,N_20732);
nor U21720 (N_21720,N_20785,N_20883);
and U21721 (N_21721,N_20073,N_20658);
or U21722 (N_21722,N_20841,N_20995);
nor U21723 (N_21723,N_20347,N_20171);
xor U21724 (N_21724,N_20111,N_20937);
and U21725 (N_21725,N_20086,N_20130);
nand U21726 (N_21726,N_20480,N_20255);
xnor U21727 (N_21727,N_20118,N_20032);
nand U21728 (N_21728,N_20651,N_20797);
and U21729 (N_21729,N_20077,N_20358);
or U21730 (N_21730,N_20040,N_20468);
nor U21731 (N_21731,N_20987,N_20812);
xnor U21732 (N_21732,N_20286,N_20547);
xnor U21733 (N_21733,N_20676,N_20956);
xnor U21734 (N_21734,N_20023,N_20322);
or U21735 (N_21735,N_20609,N_20166);
or U21736 (N_21736,N_20469,N_20993);
xnor U21737 (N_21737,N_20857,N_20110);
nor U21738 (N_21738,N_20175,N_20916);
nor U21739 (N_21739,N_20345,N_20952);
nand U21740 (N_21740,N_20327,N_20505);
and U21741 (N_21741,N_20581,N_20791);
nor U21742 (N_21742,N_20334,N_20375);
or U21743 (N_21743,N_20863,N_20594);
or U21744 (N_21744,N_20273,N_20216);
xnor U21745 (N_21745,N_20879,N_20673);
and U21746 (N_21746,N_20855,N_20891);
or U21747 (N_21747,N_20709,N_20251);
or U21748 (N_21748,N_20258,N_20518);
and U21749 (N_21749,N_20780,N_20813);
and U21750 (N_21750,N_20429,N_20038);
nor U21751 (N_21751,N_20679,N_20343);
or U21752 (N_21752,N_20261,N_20869);
xor U21753 (N_21753,N_20827,N_20368);
and U21754 (N_21754,N_20964,N_20124);
and U21755 (N_21755,N_20310,N_20039);
or U21756 (N_21756,N_20697,N_20427);
nor U21757 (N_21757,N_20984,N_20059);
or U21758 (N_21758,N_20202,N_20074);
or U21759 (N_21759,N_20939,N_20434);
nor U21760 (N_21760,N_20999,N_20914);
xnor U21761 (N_21761,N_20137,N_20755);
nand U21762 (N_21762,N_20450,N_20259);
xor U21763 (N_21763,N_20296,N_20537);
or U21764 (N_21764,N_20941,N_20974);
and U21765 (N_21765,N_20249,N_20784);
nand U21766 (N_21766,N_20364,N_20594);
or U21767 (N_21767,N_20890,N_20919);
xor U21768 (N_21768,N_20046,N_20860);
or U21769 (N_21769,N_20950,N_20943);
xor U21770 (N_21770,N_20719,N_20569);
nand U21771 (N_21771,N_20431,N_20864);
xor U21772 (N_21772,N_20217,N_20210);
nand U21773 (N_21773,N_20189,N_20767);
or U21774 (N_21774,N_20974,N_20467);
or U21775 (N_21775,N_20939,N_20491);
xnor U21776 (N_21776,N_20153,N_20601);
xnor U21777 (N_21777,N_20488,N_20575);
nand U21778 (N_21778,N_20644,N_20414);
and U21779 (N_21779,N_20580,N_20488);
or U21780 (N_21780,N_20937,N_20817);
nor U21781 (N_21781,N_20867,N_20716);
or U21782 (N_21782,N_20771,N_20940);
or U21783 (N_21783,N_20074,N_20839);
nor U21784 (N_21784,N_20440,N_20871);
xnor U21785 (N_21785,N_20681,N_20129);
nand U21786 (N_21786,N_20198,N_20575);
xnor U21787 (N_21787,N_20216,N_20309);
or U21788 (N_21788,N_20943,N_20066);
xor U21789 (N_21789,N_20000,N_20609);
and U21790 (N_21790,N_20337,N_20380);
xnor U21791 (N_21791,N_20082,N_20303);
nor U21792 (N_21792,N_20415,N_20651);
nor U21793 (N_21793,N_20630,N_20528);
nor U21794 (N_21794,N_20949,N_20438);
or U21795 (N_21795,N_20271,N_20966);
and U21796 (N_21796,N_20560,N_20107);
nor U21797 (N_21797,N_20292,N_20417);
nand U21798 (N_21798,N_20642,N_20322);
and U21799 (N_21799,N_20930,N_20525);
nor U21800 (N_21800,N_20599,N_20771);
nor U21801 (N_21801,N_20806,N_20424);
or U21802 (N_21802,N_20821,N_20067);
xor U21803 (N_21803,N_20304,N_20279);
nand U21804 (N_21804,N_20653,N_20806);
nor U21805 (N_21805,N_20114,N_20923);
nor U21806 (N_21806,N_20112,N_20159);
or U21807 (N_21807,N_20987,N_20868);
and U21808 (N_21808,N_20771,N_20876);
nand U21809 (N_21809,N_20666,N_20924);
nor U21810 (N_21810,N_20513,N_20649);
xnor U21811 (N_21811,N_20388,N_20756);
and U21812 (N_21812,N_20373,N_20742);
or U21813 (N_21813,N_20935,N_20111);
nand U21814 (N_21814,N_20003,N_20946);
and U21815 (N_21815,N_20031,N_20862);
nor U21816 (N_21816,N_20897,N_20513);
and U21817 (N_21817,N_20199,N_20727);
nor U21818 (N_21818,N_20236,N_20407);
nand U21819 (N_21819,N_20617,N_20559);
nor U21820 (N_21820,N_20676,N_20973);
and U21821 (N_21821,N_20698,N_20364);
nor U21822 (N_21822,N_20222,N_20837);
or U21823 (N_21823,N_20434,N_20027);
xor U21824 (N_21824,N_20357,N_20583);
xnor U21825 (N_21825,N_20945,N_20969);
and U21826 (N_21826,N_20488,N_20263);
and U21827 (N_21827,N_20952,N_20108);
nor U21828 (N_21828,N_20062,N_20544);
xnor U21829 (N_21829,N_20698,N_20904);
xor U21830 (N_21830,N_20606,N_20542);
or U21831 (N_21831,N_20265,N_20277);
and U21832 (N_21832,N_20626,N_20563);
or U21833 (N_21833,N_20789,N_20879);
and U21834 (N_21834,N_20116,N_20303);
nand U21835 (N_21835,N_20909,N_20288);
nand U21836 (N_21836,N_20650,N_20576);
or U21837 (N_21837,N_20400,N_20605);
nor U21838 (N_21838,N_20365,N_20969);
xor U21839 (N_21839,N_20184,N_20876);
and U21840 (N_21840,N_20365,N_20883);
or U21841 (N_21841,N_20218,N_20015);
nor U21842 (N_21842,N_20235,N_20300);
nor U21843 (N_21843,N_20281,N_20999);
or U21844 (N_21844,N_20916,N_20262);
nand U21845 (N_21845,N_20349,N_20936);
and U21846 (N_21846,N_20063,N_20388);
nand U21847 (N_21847,N_20478,N_20577);
and U21848 (N_21848,N_20867,N_20996);
xor U21849 (N_21849,N_20500,N_20643);
xor U21850 (N_21850,N_20388,N_20895);
nand U21851 (N_21851,N_20778,N_20337);
xor U21852 (N_21852,N_20992,N_20414);
xnor U21853 (N_21853,N_20611,N_20645);
xor U21854 (N_21854,N_20082,N_20282);
or U21855 (N_21855,N_20673,N_20667);
xnor U21856 (N_21856,N_20257,N_20123);
nand U21857 (N_21857,N_20888,N_20708);
xnor U21858 (N_21858,N_20322,N_20676);
nor U21859 (N_21859,N_20711,N_20659);
or U21860 (N_21860,N_20211,N_20718);
nor U21861 (N_21861,N_20732,N_20018);
xor U21862 (N_21862,N_20313,N_20401);
or U21863 (N_21863,N_20949,N_20733);
nor U21864 (N_21864,N_20543,N_20421);
nand U21865 (N_21865,N_20082,N_20543);
and U21866 (N_21866,N_20702,N_20236);
or U21867 (N_21867,N_20336,N_20210);
xor U21868 (N_21868,N_20393,N_20234);
nand U21869 (N_21869,N_20666,N_20730);
or U21870 (N_21870,N_20962,N_20897);
nor U21871 (N_21871,N_20662,N_20977);
or U21872 (N_21872,N_20792,N_20119);
xnor U21873 (N_21873,N_20786,N_20076);
nand U21874 (N_21874,N_20482,N_20468);
nor U21875 (N_21875,N_20012,N_20778);
nor U21876 (N_21876,N_20637,N_20267);
xnor U21877 (N_21877,N_20074,N_20747);
nor U21878 (N_21878,N_20797,N_20264);
or U21879 (N_21879,N_20339,N_20120);
xnor U21880 (N_21880,N_20233,N_20291);
and U21881 (N_21881,N_20563,N_20269);
or U21882 (N_21882,N_20198,N_20260);
or U21883 (N_21883,N_20175,N_20584);
xor U21884 (N_21884,N_20239,N_20161);
or U21885 (N_21885,N_20857,N_20674);
nor U21886 (N_21886,N_20936,N_20867);
and U21887 (N_21887,N_20984,N_20259);
nor U21888 (N_21888,N_20786,N_20929);
xor U21889 (N_21889,N_20152,N_20995);
nand U21890 (N_21890,N_20966,N_20480);
xnor U21891 (N_21891,N_20760,N_20880);
nand U21892 (N_21892,N_20999,N_20130);
nor U21893 (N_21893,N_20405,N_20751);
and U21894 (N_21894,N_20283,N_20911);
nor U21895 (N_21895,N_20158,N_20443);
or U21896 (N_21896,N_20301,N_20807);
and U21897 (N_21897,N_20368,N_20156);
nor U21898 (N_21898,N_20995,N_20138);
nand U21899 (N_21899,N_20268,N_20391);
nand U21900 (N_21900,N_20696,N_20151);
or U21901 (N_21901,N_20145,N_20144);
nand U21902 (N_21902,N_20169,N_20673);
or U21903 (N_21903,N_20130,N_20433);
nand U21904 (N_21904,N_20117,N_20403);
or U21905 (N_21905,N_20297,N_20673);
xor U21906 (N_21906,N_20850,N_20038);
nand U21907 (N_21907,N_20723,N_20282);
nor U21908 (N_21908,N_20119,N_20059);
and U21909 (N_21909,N_20820,N_20130);
xor U21910 (N_21910,N_20464,N_20432);
nor U21911 (N_21911,N_20707,N_20108);
xnor U21912 (N_21912,N_20125,N_20446);
and U21913 (N_21913,N_20289,N_20781);
xnor U21914 (N_21914,N_20630,N_20339);
xor U21915 (N_21915,N_20762,N_20971);
or U21916 (N_21916,N_20636,N_20565);
nor U21917 (N_21917,N_20349,N_20925);
xnor U21918 (N_21918,N_20833,N_20534);
nor U21919 (N_21919,N_20125,N_20564);
or U21920 (N_21920,N_20990,N_20226);
nand U21921 (N_21921,N_20801,N_20297);
nand U21922 (N_21922,N_20503,N_20060);
nand U21923 (N_21923,N_20642,N_20818);
and U21924 (N_21924,N_20898,N_20985);
nand U21925 (N_21925,N_20510,N_20574);
xor U21926 (N_21926,N_20238,N_20605);
nand U21927 (N_21927,N_20143,N_20047);
or U21928 (N_21928,N_20570,N_20431);
or U21929 (N_21929,N_20153,N_20139);
nor U21930 (N_21930,N_20845,N_20791);
xor U21931 (N_21931,N_20609,N_20520);
and U21932 (N_21932,N_20364,N_20099);
nor U21933 (N_21933,N_20639,N_20782);
or U21934 (N_21934,N_20016,N_20624);
nand U21935 (N_21935,N_20600,N_20417);
or U21936 (N_21936,N_20668,N_20972);
nand U21937 (N_21937,N_20758,N_20078);
or U21938 (N_21938,N_20213,N_20167);
nor U21939 (N_21939,N_20332,N_20403);
or U21940 (N_21940,N_20417,N_20433);
xnor U21941 (N_21941,N_20718,N_20850);
nor U21942 (N_21942,N_20749,N_20557);
or U21943 (N_21943,N_20528,N_20486);
nor U21944 (N_21944,N_20730,N_20911);
and U21945 (N_21945,N_20075,N_20834);
and U21946 (N_21946,N_20587,N_20407);
or U21947 (N_21947,N_20924,N_20790);
xnor U21948 (N_21948,N_20731,N_20032);
or U21949 (N_21949,N_20825,N_20216);
xor U21950 (N_21950,N_20579,N_20611);
xnor U21951 (N_21951,N_20719,N_20711);
or U21952 (N_21952,N_20759,N_20133);
nand U21953 (N_21953,N_20628,N_20313);
nor U21954 (N_21954,N_20348,N_20851);
and U21955 (N_21955,N_20557,N_20423);
or U21956 (N_21956,N_20251,N_20645);
and U21957 (N_21957,N_20098,N_20255);
nand U21958 (N_21958,N_20560,N_20884);
and U21959 (N_21959,N_20735,N_20556);
or U21960 (N_21960,N_20203,N_20344);
or U21961 (N_21961,N_20177,N_20779);
nand U21962 (N_21962,N_20861,N_20174);
xnor U21963 (N_21963,N_20837,N_20260);
and U21964 (N_21964,N_20848,N_20009);
nand U21965 (N_21965,N_20444,N_20285);
or U21966 (N_21966,N_20205,N_20004);
nand U21967 (N_21967,N_20644,N_20533);
nor U21968 (N_21968,N_20059,N_20620);
and U21969 (N_21969,N_20499,N_20463);
or U21970 (N_21970,N_20811,N_20176);
and U21971 (N_21971,N_20037,N_20929);
and U21972 (N_21972,N_20099,N_20823);
and U21973 (N_21973,N_20343,N_20142);
and U21974 (N_21974,N_20998,N_20462);
nor U21975 (N_21975,N_20703,N_20078);
xor U21976 (N_21976,N_20604,N_20292);
xor U21977 (N_21977,N_20886,N_20932);
xor U21978 (N_21978,N_20276,N_20666);
nor U21979 (N_21979,N_20488,N_20348);
or U21980 (N_21980,N_20503,N_20983);
nand U21981 (N_21981,N_20845,N_20551);
and U21982 (N_21982,N_20828,N_20980);
nor U21983 (N_21983,N_20164,N_20100);
or U21984 (N_21984,N_20571,N_20036);
xor U21985 (N_21985,N_20930,N_20346);
xor U21986 (N_21986,N_20157,N_20124);
xnor U21987 (N_21987,N_20160,N_20612);
or U21988 (N_21988,N_20341,N_20510);
nand U21989 (N_21989,N_20857,N_20669);
nand U21990 (N_21990,N_20681,N_20695);
nand U21991 (N_21991,N_20785,N_20604);
and U21992 (N_21992,N_20265,N_20956);
and U21993 (N_21993,N_20452,N_20364);
and U21994 (N_21994,N_20264,N_20637);
and U21995 (N_21995,N_20310,N_20540);
nor U21996 (N_21996,N_20471,N_20394);
and U21997 (N_21997,N_20807,N_20253);
nand U21998 (N_21998,N_20697,N_20002);
or U21999 (N_21999,N_20426,N_20371);
xnor U22000 (N_22000,N_21962,N_21934);
nor U22001 (N_22001,N_21252,N_21900);
or U22002 (N_22002,N_21444,N_21313);
nor U22003 (N_22003,N_21331,N_21179);
xnor U22004 (N_22004,N_21165,N_21554);
and U22005 (N_22005,N_21149,N_21446);
xnor U22006 (N_22006,N_21615,N_21360);
nor U22007 (N_22007,N_21523,N_21792);
nor U22008 (N_22008,N_21551,N_21194);
or U22009 (N_22009,N_21354,N_21879);
nand U22010 (N_22010,N_21261,N_21238);
and U22011 (N_22011,N_21851,N_21706);
xnor U22012 (N_22012,N_21166,N_21480);
xor U22013 (N_22013,N_21545,N_21178);
xnor U22014 (N_22014,N_21002,N_21999);
nor U22015 (N_22015,N_21117,N_21952);
nand U22016 (N_22016,N_21373,N_21724);
and U22017 (N_22017,N_21870,N_21563);
xnor U22018 (N_22018,N_21335,N_21009);
xnor U22019 (N_22019,N_21232,N_21186);
or U22020 (N_22020,N_21182,N_21597);
or U22021 (N_22021,N_21134,N_21028);
or U22022 (N_22022,N_21422,N_21296);
xnor U22023 (N_22023,N_21547,N_21338);
or U22024 (N_22024,N_21702,N_21796);
and U22025 (N_22025,N_21124,N_21929);
nand U22026 (N_22026,N_21823,N_21483);
nand U22027 (N_22027,N_21986,N_21384);
nand U22028 (N_22028,N_21285,N_21287);
and U22029 (N_22029,N_21827,N_21522);
xor U22030 (N_22030,N_21111,N_21963);
nand U22031 (N_22031,N_21095,N_21618);
xor U22032 (N_22032,N_21072,N_21192);
and U22033 (N_22033,N_21731,N_21696);
or U22034 (N_22034,N_21803,N_21294);
xor U22035 (N_22035,N_21006,N_21251);
nand U22036 (N_22036,N_21040,N_21975);
nor U22037 (N_22037,N_21454,N_21121);
and U22038 (N_22038,N_21332,N_21498);
or U22039 (N_22039,N_21814,N_21998);
or U22040 (N_22040,N_21459,N_21381);
and U22041 (N_22041,N_21704,N_21090);
nor U22042 (N_22042,N_21966,N_21369);
and U22043 (N_22043,N_21687,N_21189);
or U22044 (N_22044,N_21712,N_21642);
nor U22045 (N_22045,N_21004,N_21030);
and U22046 (N_22046,N_21895,N_21118);
or U22047 (N_22047,N_21208,N_21160);
nor U22048 (N_22048,N_21525,N_21315);
nand U22049 (N_22049,N_21925,N_21809);
and U22050 (N_22050,N_21772,N_21861);
nor U22051 (N_22051,N_21484,N_21099);
xor U22052 (N_22052,N_21184,N_21911);
xor U22053 (N_22053,N_21461,N_21862);
xor U22054 (N_22054,N_21511,N_21056);
nor U22055 (N_22055,N_21539,N_21541);
nor U22056 (N_22056,N_21746,N_21938);
nor U22057 (N_22057,N_21964,N_21630);
or U22058 (N_22058,N_21295,N_21209);
xnor U22059 (N_22059,N_21005,N_21282);
and U22060 (N_22060,N_21932,N_21220);
nor U22061 (N_22061,N_21164,N_21361);
nor U22062 (N_22062,N_21349,N_21427);
nand U22063 (N_22063,N_21916,N_21265);
nor U22064 (N_22064,N_21123,N_21730);
nand U22065 (N_22065,N_21070,N_21061);
and U22066 (N_22066,N_21489,N_21799);
nand U22067 (N_22067,N_21626,N_21333);
xor U22068 (N_22068,N_21579,N_21717);
nand U22069 (N_22069,N_21752,N_21711);
xor U22070 (N_22070,N_21585,N_21259);
and U22071 (N_22071,N_21214,N_21413);
nor U22072 (N_22072,N_21695,N_21045);
and U22073 (N_22073,N_21927,N_21219);
nand U22074 (N_22074,N_21170,N_21949);
or U22075 (N_22075,N_21556,N_21302);
nand U22076 (N_22076,N_21364,N_21750);
xor U22077 (N_22077,N_21725,N_21942);
and U22078 (N_22078,N_21771,N_21253);
or U22079 (N_22079,N_21375,N_21041);
or U22080 (N_22080,N_21158,N_21866);
and U22081 (N_22081,N_21495,N_21403);
or U22082 (N_22082,N_21723,N_21212);
and U22083 (N_22083,N_21046,N_21091);
nor U22084 (N_22084,N_21671,N_21419);
nand U22085 (N_22085,N_21678,N_21007);
or U22086 (N_22086,N_21635,N_21255);
xor U22087 (N_22087,N_21292,N_21588);
or U22088 (N_22088,N_21162,N_21393);
nor U22089 (N_22089,N_21576,N_21574);
nor U22090 (N_22090,N_21137,N_21893);
nor U22091 (N_22091,N_21445,N_21082);
or U22092 (N_22092,N_21620,N_21339);
nand U22093 (N_22093,N_21698,N_21979);
or U22094 (N_22094,N_21264,N_21652);
or U22095 (N_22095,N_21584,N_21677);
nor U22096 (N_22096,N_21125,N_21863);
nand U22097 (N_22097,N_21318,N_21044);
and U22098 (N_22098,N_21751,N_21150);
nand U22099 (N_22099,N_21096,N_21831);
xnor U22100 (N_22100,N_21562,N_21856);
nand U22101 (N_22101,N_21634,N_21036);
nand U22102 (N_22102,N_21502,N_21146);
xor U22103 (N_22103,N_21719,N_21790);
nor U22104 (N_22104,N_21699,N_21303);
nor U22105 (N_22105,N_21992,N_21604);
and U22106 (N_22106,N_21055,N_21506);
xnor U22107 (N_22107,N_21376,N_21365);
and U22108 (N_22108,N_21367,N_21266);
or U22109 (N_22109,N_21016,N_21163);
or U22110 (N_22110,N_21518,N_21802);
or U22111 (N_22111,N_21819,N_21157);
xor U22112 (N_22112,N_21644,N_21936);
and U22113 (N_22113,N_21300,N_21305);
xnor U22114 (N_22114,N_21460,N_21756);
nand U22115 (N_22115,N_21434,N_21449);
and U22116 (N_22116,N_21477,N_21392);
nor U22117 (N_22117,N_21015,N_21472);
or U22118 (N_22118,N_21571,N_21793);
and U22119 (N_22119,N_21019,N_21269);
nor U22120 (N_22120,N_21279,N_21665);
and U22121 (N_22121,N_21476,N_21977);
xnor U22122 (N_22122,N_21374,N_21425);
nand U22123 (N_22123,N_21818,N_21967);
xnor U22124 (N_22124,N_21235,N_21071);
or U22125 (N_22125,N_21560,N_21878);
nand U22126 (N_22126,N_21749,N_21700);
or U22127 (N_22127,N_21093,N_21910);
or U22128 (N_22128,N_21097,N_21951);
and U22129 (N_22129,N_21216,N_21853);
or U22130 (N_22130,N_21815,N_21538);
or U22131 (N_22131,N_21281,N_21394);
or U22132 (N_22132,N_21196,N_21570);
nor U22133 (N_22133,N_21262,N_21778);
and U22134 (N_22134,N_21565,N_21410);
xnor U22135 (N_22135,N_21140,N_21894);
or U22136 (N_22136,N_21989,N_21116);
nand U22137 (N_22137,N_21453,N_21283);
and U22138 (N_22138,N_21368,N_21181);
or U22139 (N_22139,N_21325,N_21268);
nand U22140 (N_22140,N_21231,N_21693);
xnor U22141 (N_22141,N_21913,N_21222);
nor U22142 (N_22142,N_21583,N_21314);
xnor U22143 (N_22143,N_21600,N_21310);
xor U22144 (N_22144,N_21024,N_21548);
or U22145 (N_22145,N_21891,N_21138);
nand U22146 (N_22146,N_21038,N_21566);
xor U22147 (N_22147,N_21593,N_21785);
or U22148 (N_22148,N_21439,N_21844);
nand U22149 (N_22149,N_21464,N_21843);
and U22150 (N_22150,N_21256,N_21727);
xnor U22151 (N_22151,N_21039,N_21330);
nand U22152 (N_22152,N_21864,N_21397);
nor U22153 (N_22153,N_21985,N_21470);
nor U22154 (N_22154,N_21744,N_21976);
nand U22155 (N_22155,N_21766,N_21175);
nor U22156 (N_22156,N_21591,N_21546);
xnor U22157 (N_22157,N_21662,N_21807);
nor U22158 (N_22158,N_21120,N_21737);
or U22159 (N_22159,N_21567,N_21906);
xnor U22160 (N_22160,N_21504,N_21887);
and U22161 (N_22161,N_21892,N_21855);
nand U22162 (N_22162,N_21645,N_21564);
nor U22163 (N_22163,N_21580,N_21898);
and U22164 (N_22164,N_21277,N_21063);
nand U22165 (N_22165,N_21057,N_21648);
nand U22166 (N_22166,N_21743,N_21596);
and U22167 (N_22167,N_21904,N_21358);
xor U22168 (N_22168,N_21903,N_21107);
xor U22169 (N_22169,N_21833,N_21738);
xor U22170 (N_22170,N_21794,N_21681);
or U22171 (N_22171,N_21404,N_21025);
and U22172 (N_22172,N_21176,N_21488);
and U22173 (N_22173,N_21234,N_21399);
and U22174 (N_22174,N_21854,N_21380);
or U22175 (N_22175,N_21633,N_21774);
nand U22176 (N_22176,N_21608,N_21917);
nor U22177 (N_22177,N_21517,N_21048);
nand U22178 (N_22178,N_21215,N_21602);
and U22179 (N_22179,N_21312,N_21928);
nand U22180 (N_22180,N_21883,N_21968);
and U22181 (N_22181,N_21629,N_21379);
or U22182 (N_22182,N_21735,N_21617);
nand U22183 (N_22183,N_21027,N_21590);
xor U22184 (N_22184,N_21675,N_21202);
or U22185 (N_22185,N_21901,N_21466);
and U22186 (N_22186,N_21000,N_21837);
xnor U22187 (N_22187,N_21748,N_21406);
xor U22188 (N_22188,N_21961,N_21236);
xor U22189 (N_22189,N_21289,N_21508);
and U22190 (N_22190,N_21426,N_21156);
nor U22191 (N_22191,N_21616,N_21280);
nor U22192 (N_22192,N_21018,N_21653);
xor U22193 (N_22193,N_21153,N_21352);
or U22194 (N_22194,N_21243,N_21020);
and U22195 (N_22195,N_21142,N_21520);
nor U22196 (N_22196,N_21258,N_21346);
and U22197 (N_22197,N_21104,N_21185);
xor U22198 (N_22198,N_21919,N_21022);
nand U22199 (N_22199,N_21247,N_21801);
nor U22200 (N_22200,N_21415,N_21326);
nor U22201 (N_22201,N_21958,N_21143);
or U22202 (N_22202,N_21909,N_21159);
xnor U22203 (N_22203,N_21788,N_21713);
or U22204 (N_22204,N_21168,N_21612);
nor U22205 (N_22205,N_21848,N_21775);
xor U22206 (N_22206,N_21536,N_21356);
or U22207 (N_22207,N_21205,N_21284);
and U22208 (N_22208,N_21937,N_21797);
nor U22209 (N_22209,N_21047,N_21430);
xor U22210 (N_22210,N_21885,N_21921);
nand U22211 (N_22211,N_21126,N_21133);
xnor U22212 (N_22212,N_21290,N_21073);
or U22213 (N_22213,N_21011,N_21442);
or U22214 (N_22214,N_21941,N_21501);
or U22215 (N_22215,N_21776,N_21694);
or U22216 (N_22216,N_21553,N_21697);
nor U22217 (N_22217,N_21079,N_21327);
nand U22218 (N_22218,N_21759,N_21631);
nor U22219 (N_22219,N_21715,N_21703);
xor U22220 (N_22220,N_21709,N_21207);
or U22221 (N_22221,N_21824,N_21217);
xor U22222 (N_22222,N_21400,N_21203);
nand U22223 (N_22223,N_21667,N_21969);
or U22224 (N_22224,N_21198,N_21291);
nor U22225 (N_22225,N_21605,N_21533);
and U22226 (N_22226,N_21660,N_21573);
nand U22227 (N_22227,N_21328,N_21656);
and U22228 (N_22228,N_21119,N_21228);
or U22229 (N_22229,N_21761,N_21388);
and U22230 (N_22230,N_21940,N_21896);
or U22231 (N_22231,N_21514,N_21462);
nand U22232 (N_22232,N_21537,N_21492);
and U22233 (N_22233,N_21943,N_21524);
or U22234 (N_22234,N_21768,N_21263);
nand U22235 (N_22235,N_21211,N_21062);
nand U22236 (N_22236,N_21329,N_21347);
and U22237 (N_22237,N_21722,N_21147);
or U22238 (N_22238,N_21435,N_21603);
and U22239 (N_22239,N_21114,N_21650);
and U22240 (N_22240,N_21805,N_21569);
and U22241 (N_22241,N_21420,N_21859);
nor U22242 (N_22242,N_21884,N_21417);
nand U22243 (N_22243,N_21842,N_21069);
xnor U22244 (N_22244,N_21601,N_21270);
nor U22245 (N_22245,N_21075,N_21670);
nor U22246 (N_22246,N_21663,N_21475);
and U22247 (N_22247,N_21944,N_21353);
or U22248 (N_22248,N_21613,N_21486);
xnor U22249 (N_22249,N_21409,N_21915);
and U22250 (N_22250,N_21276,N_21307);
xnor U22251 (N_22251,N_21250,N_21920);
xnor U22252 (N_22252,N_21032,N_21619);
nand U22253 (N_22253,N_21254,N_21273);
xnor U22254 (N_22254,N_21177,N_21762);
nor U22255 (N_22255,N_21974,N_21973);
nor U22256 (N_22256,N_21197,N_21995);
or U22257 (N_22257,N_21960,N_21721);
xnor U22258 (N_22258,N_21780,N_21610);
nand U22259 (N_22259,N_21396,N_21609);
or U22260 (N_22260,N_21385,N_21688);
and U22261 (N_22261,N_21151,N_21306);
and U22262 (N_22262,N_21757,N_21267);
xnor U22263 (N_22263,N_21260,N_21233);
and U22264 (N_22264,N_21230,N_21463);
or U22265 (N_22265,N_21997,N_21543);
xnor U22266 (N_22266,N_21129,N_21053);
nand U22267 (N_22267,N_21414,N_21529);
xor U22268 (N_22268,N_21674,N_21043);
xor U22269 (N_22269,N_21206,N_21003);
nor U22270 (N_22270,N_21734,N_21383);
nor U22271 (N_22271,N_21589,N_21174);
nor U22272 (N_22272,N_21226,N_21431);
and U22273 (N_22273,N_21402,N_21786);
xnor U22274 (N_22274,N_21448,N_21673);
nand U22275 (N_22275,N_21391,N_21144);
and U22276 (N_22276,N_21691,N_21881);
xnor U22277 (N_22277,N_21077,N_21707);
or U22278 (N_22278,N_21363,N_21587);
nor U22279 (N_22279,N_21672,N_21437);
and U22280 (N_22280,N_21549,N_21485);
nand U22281 (N_22281,N_21922,N_21939);
nor U22282 (N_22282,N_21987,N_21804);
or U22283 (N_22283,N_21244,N_21741);
or U22284 (N_22284,N_21708,N_21646);
or U22285 (N_22285,N_21304,N_21732);
and U22286 (N_22286,N_21607,N_21516);
xnor U22287 (N_22287,N_21440,N_21808);
and U22288 (N_22288,N_21227,N_21865);
and U22289 (N_22289,N_21994,N_21828);
nor U22290 (N_22290,N_21013,N_21468);
nor U22291 (N_22291,N_21052,N_21078);
nand U22292 (N_22292,N_21760,N_21337);
and U22293 (N_22293,N_21873,N_21274);
or U22294 (N_22294,N_21647,N_21552);
nor U22295 (N_22295,N_21035,N_21301);
nor U22296 (N_22296,N_21297,N_21868);
or U22297 (N_22297,N_21481,N_21362);
or U22298 (N_22298,N_21850,N_21351);
xnor U22299 (N_22299,N_21320,N_21897);
or U22300 (N_22300,N_21763,N_21739);
nand U22301 (N_22301,N_21110,N_21640);
nor U22302 (N_22302,N_21953,N_21931);
nand U22303 (N_22303,N_21606,N_21578);
xnor U22304 (N_22304,N_21066,N_21990);
or U22305 (N_22305,N_21371,N_21218);
nand U22306 (N_22306,N_21658,N_21221);
and U22307 (N_22307,N_21372,N_21465);
nand U22308 (N_22308,N_21034,N_21272);
xnor U22309 (N_22309,N_21764,N_21542);
and U22310 (N_22310,N_21836,N_21503);
and U22311 (N_22311,N_21487,N_21581);
or U22312 (N_22312,N_21298,N_21201);
or U22313 (N_22313,N_21017,N_21886);
nand U22314 (N_22314,N_21458,N_21857);
and U22315 (N_22315,N_21594,N_21271);
and U22316 (N_22316,N_21237,N_21049);
xnor U22317 (N_22317,N_21135,N_21474);
or U22318 (N_22318,N_21187,N_21710);
nor U22319 (N_22319,N_21981,N_21521);
xnor U22320 (N_22320,N_21101,N_21154);
xor U22321 (N_22321,N_21935,N_21659);
or U22322 (N_22322,N_21342,N_21991);
nor U22323 (N_22323,N_21954,N_21195);
and U22324 (N_22324,N_21343,N_21692);
or U22325 (N_22325,N_21357,N_21102);
xnor U22326 (N_22326,N_21467,N_21872);
nand U22327 (N_22327,N_21544,N_21745);
and U22328 (N_22328,N_21145,N_21683);
or U22329 (N_22329,N_21155,N_21348);
xor U22330 (N_22330,N_21705,N_21782);
or U22331 (N_22331,N_21051,N_21497);
or U22332 (N_22332,N_21558,N_21507);
nand U22333 (N_22333,N_21905,N_21575);
nor U22334 (N_22334,N_21639,N_21889);
xnor U22335 (N_22335,N_21424,N_21317);
nand U22336 (N_22336,N_21914,N_21173);
or U22337 (N_22337,N_21638,N_21190);
nand U22338 (N_22338,N_21029,N_21065);
or U22339 (N_22339,N_21500,N_21847);
xor U22340 (N_22340,N_21867,N_21161);
or U22341 (N_22341,N_21088,N_21479);
or U22342 (N_22342,N_21664,N_21471);
and U22343 (N_22343,N_21682,N_21918);
nand U22344 (N_22344,N_21882,N_21433);
nor U22345 (N_22345,N_21770,N_21390);
nor U22346 (N_22346,N_21510,N_21685);
nor U22347 (N_22347,N_21115,N_21060);
or U22348 (N_22348,N_21334,N_21728);
nand U22349 (N_22349,N_21496,N_21996);
nand U22350 (N_22350,N_21316,N_21223);
xor U22351 (N_22351,N_21199,N_21628);
nor U22352 (N_22352,N_21740,N_21210);
and U22353 (N_22353,N_21655,N_21094);
xor U22354 (N_22354,N_21152,N_21299);
nor U22355 (N_22355,N_21686,N_21323);
nor U22356 (N_22356,N_21622,N_21846);
and U22357 (N_22357,N_21742,N_21395);
or U22358 (N_22358,N_21169,N_21971);
and U22359 (N_22359,N_21825,N_21447);
and U22360 (N_22360,N_21482,N_21311);
and U22361 (N_22361,N_21350,N_21319);
and U22362 (N_22362,N_21008,N_21451);
nor U22363 (N_22363,N_21528,N_21042);
nor U22364 (N_22364,N_21359,N_21001);
nand U22365 (N_22365,N_21183,N_21755);
nor U22366 (N_22366,N_21085,N_21515);
nand U22367 (N_22367,N_21172,N_21972);
or U22368 (N_22368,N_21241,N_21355);
and U22369 (N_22369,N_21436,N_21984);
and U22370 (N_22370,N_21758,N_21945);
and U22371 (N_22371,N_21200,N_21880);
nand U22372 (N_22372,N_21530,N_21970);
or U22373 (N_22373,N_21980,N_21534);
nand U22374 (N_22374,N_21509,N_21401);
and U22375 (N_22375,N_21012,N_21754);
xor U22376 (N_22376,N_21188,N_21816);
nand U22377 (N_22377,N_21614,N_21457);
xor U22378 (N_22378,N_21769,N_21108);
xnor U22379 (N_22379,N_21398,N_21240);
nor U22380 (N_22380,N_21010,N_21956);
and U22381 (N_22381,N_21838,N_21651);
or U22382 (N_22382,N_21561,N_21874);
nor U22383 (N_22383,N_21204,N_21643);
nand U22384 (N_22384,N_21926,N_21382);
nand U22385 (N_22385,N_21321,N_21054);
nand U22386 (N_22386,N_21781,N_21611);
nand U22387 (N_22387,N_21930,N_21733);
and U22388 (N_22388,N_21387,N_21021);
and U22389 (N_22389,N_21978,N_21888);
and U22390 (N_22390,N_21378,N_21167);
nand U22391 (N_22391,N_21679,N_21595);
and U22392 (N_22392,N_21806,N_21582);
xor U22393 (N_22393,N_21993,N_21257);
xor U22394 (N_22394,N_21798,N_21416);
or U22395 (N_22395,N_21813,N_21947);
nand U22396 (N_22396,N_21246,N_21491);
nand U22397 (N_22397,N_21418,N_21821);
or U22398 (N_22398,N_21869,N_21726);
nand U22399 (N_22399,N_21412,N_21127);
and U22400 (N_22400,N_21193,N_21014);
nand U22401 (N_22401,N_21624,N_21789);
nor U22402 (N_22402,N_21641,N_21852);
xor U22403 (N_22403,N_21113,N_21811);
and U22404 (N_22404,N_21109,N_21407);
and U22405 (N_22405,N_21309,N_21242);
xor U22406 (N_22406,N_21669,N_21141);
xor U22407 (N_22407,N_21950,N_21139);
or U22408 (N_22408,N_21820,N_21136);
nand U22409 (N_22409,N_21432,N_21983);
nor U22410 (N_22410,N_21627,N_21845);
or U22411 (N_22411,N_21288,N_21599);
nor U22412 (N_22412,N_21405,N_21948);
and U22413 (N_22413,N_21438,N_21103);
nand U22414 (N_22414,N_21858,N_21526);
and U22415 (N_22415,N_21493,N_21248);
xnor U22416 (N_22416,N_21690,N_21907);
nor U22417 (N_22417,N_21033,N_21224);
and U22418 (N_22418,N_21875,N_21191);
and U22419 (N_22419,N_21832,N_21512);
xnor U22420 (N_22420,N_21787,N_21171);
and U22421 (N_22421,N_21074,N_21747);
xor U22422 (N_22422,N_21598,N_21965);
or U22423 (N_22423,N_21666,N_21377);
nand U22424 (N_22424,N_21657,N_21822);
nor U22425 (N_22425,N_21701,N_21689);
and U22426 (N_22426,N_21540,N_21473);
and U22427 (N_22427,N_21621,N_21773);
xnor U22428 (N_22428,N_21668,N_21087);
and U22429 (N_22429,N_21982,N_21933);
xnor U22430 (N_22430,N_21112,N_21654);
nor U22431 (N_22431,N_21849,N_21084);
xor U22432 (N_22432,N_21322,N_21286);
nand U22433 (N_22433,N_21946,N_21527);
and U22434 (N_22434,N_21649,N_21389);
xor U22435 (N_22435,N_21469,N_21592);
or U22436 (N_22436,N_21455,N_21344);
nand U22437 (N_22437,N_21429,N_21059);
nor U22438 (N_22438,N_21083,N_21408);
xor U22439 (N_22439,N_21513,N_21988);
nand U22440 (N_22440,N_21637,N_21341);
nor U22441 (N_22441,N_21586,N_21278);
and U22442 (N_22442,N_21105,N_21089);
and U22443 (N_22443,N_21494,N_21092);
and U22444 (N_22444,N_21876,N_21568);
xnor U22445 (N_22445,N_21924,N_21718);
xnor U22446 (N_22446,N_21841,N_21490);
nand U22447 (N_22447,N_21531,N_21839);
and U22448 (N_22448,N_21275,N_21784);
and U22449 (N_22449,N_21908,N_21800);
nor U22450 (N_22450,N_21625,N_21577);
and U22451 (N_22451,N_21308,N_21148);
and U22452 (N_22452,N_21519,N_21676);
and U22453 (N_22453,N_21370,N_21661);
nand U22454 (N_22454,N_21064,N_21923);
and U22455 (N_22455,N_21450,N_21239);
or U22456 (N_22456,N_21213,N_21680);
and U22457 (N_22457,N_21428,N_21452);
or U22458 (N_22458,N_21421,N_21100);
nor U22459 (N_22459,N_21559,N_21058);
nand U22460 (N_22460,N_21031,N_21955);
nor U22461 (N_22461,N_21795,N_21765);
nand U22462 (N_22462,N_21249,N_21128);
nand U22463 (N_22463,N_21753,N_21081);
xnor U22464 (N_22464,N_21130,N_21899);
or U22465 (N_22465,N_21791,N_21779);
or U22466 (N_22466,N_21098,N_21817);
and U22467 (N_22467,N_21386,N_21826);
and U22468 (N_22468,N_21026,N_21037);
nand U22469 (N_22469,N_21871,N_21636);
nand U22470 (N_22470,N_21834,N_21877);
or U22471 (N_22471,N_21716,N_21912);
and U22472 (N_22472,N_21720,N_21443);
nor U22473 (N_22473,N_21535,N_21366);
or U22474 (N_22474,N_21729,N_21957);
nor U22475 (N_22475,N_21180,N_21840);
nand U22476 (N_22476,N_21835,N_21122);
or U22477 (N_22477,N_21767,N_21736);
nand U22478 (N_22478,N_21812,N_21810);
nand U22479 (N_22479,N_21068,N_21632);
and U22480 (N_22480,N_21456,N_21505);
or U22481 (N_22481,N_21714,N_21423);
nor U22482 (N_22482,N_21067,N_21829);
and U22483 (N_22483,N_21132,N_21890);
nand U22484 (N_22484,N_21557,N_21245);
and U22485 (N_22485,N_21080,N_21555);
xnor U22486 (N_22486,N_21345,N_21550);
nor U22487 (N_22487,N_21336,N_21229);
nand U22488 (N_22488,N_21293,N_21076);
and U22489 (N_22489,N_21572,N_21783);
xor U22490 (N_22490,N_21106,N_21050);
and U22491 (N_22491,N_21324,N_21411);
xor U22492 (N_22492,N_21131,N_21623);
and U22493 (N_22493,N_21830,N_21902);
and U22494 (N_22494,N_21340,N_21478);
or U22495 (N_22495,N_21532,N_21959);
and U22496 (N_22496,N_21441,N_21684);
or U22497 (N_22497,N_21023,N_21225);
and U22498 (N_22498,N_21499,N_21777);
nand U22499 (N_22499,N_21860,N_21086);
nand U22500 (N_22500,N_21626,N_21429);
and U22501 (N_22501,N_21967,N_21074);
xor U22502 (N_22502,N_21967,N_21533);
nor U22503 (N_22503,N_21021,N_21042);
nand U22504 (N_22504,N_21179,N_21051);
nand U22505 (N_22505,N_21335,N_21076);
nor U22506 (N_22506,N_21317,N_21761);
xor U22507 (N_22507,N_21117,N_21786);
xor U22508 (N_22508,N_21902,N_21120);
nor U22509 (N_22509,N_21053,N_21833);
xnor U22510 (N_22510,N_21727,N_21705);
xnor U22511 (N_22511,N_21658,N_21841);
or U22512 (N_22512,N_21956,N_21685);
nor U22513 (N_22513,N_21634,N_21980);
xnor U22514 (N_22514,N_21802,N_21701);
nand U22515 (N_22515,N_21938,N_21709);
or U22516 (N_22516,N_21763,N_21638);
or U22517 (N_22517,N_21902,N_21606);
nand U22518 (N_22518,N_21851,N_21197);
or U22519 (N_22519,N_21091,N_21872);
nand U22520 (N_22520,N_21229,N_21478);
nand U22521 (N_22521,N_21784,N_21688);
or U22522 (N_22522,N_21166,N_21959);
xor U22523 (N_22523,N_21930,N_21280);
or U22524 (N_22524,N_21471,N_21686);
or U22525 (N_22525,N_21510,N_21330);
xor U22526 (N_22526,N_21317,N_21721);
nor U22527 (N_22527,N_21530,N_21236);
nor U22528 (N_22528,N_21622,N_21943);
nand U22529 (N_22529,N_21052,N_21997);
or U22530 (N_22530,N_21074,N_21815);
xnor U22531 (N_22531,N_21926,N_21481);
xnor U22532 (N_22532,N_21850,N_21285);
nor U22533 (N_22533,N_21123,N_21896);
and U22534 (N_22534,N_21984,N_21299);
nand U22535 (N_22535,N_21582,N_21464);
nor U22536 (N_22536,N_21420,N_21340);
nor U22537 (N_22537,N_21276,N_21928);
and U22538 (N_22538,N_21688,N_21970);
xor U22539 (N_22539,N_21962,N_21674);
nand U22540 (N_22540,N_21101,N_21452);
nand U22541 (N_22541,N_21042,N_21685);
nor U22542 (N_22542,N_21462,N_21134);
nor U22543 (N_22543,N_21355,N_21906);
nand U22544 (N_22544,N_21948,N_21988);
xnor U22545 (N_22545,N_21474,N_21866);
xor U22546 (N_22546,N_21495,N_21795);
xnor U22547 (N_22547,N_21627,N_21448);
xnor U22548 (N_22548,N_21353,N_21473);
nand U22549 (N_22549,N_21651,N_21796);
xor U22550 (N_22550,N_21260,N_21124);
and U22551 (N_22551,N_21106,N_21159);
or U22552 (N_22552,N_21439,N_21651);
or U22553 (N_22553,N_21195,N_21713);
or U22554 (N_22554,N_21455,N_21942);
nand U22555 (N_22555,N_21101,N_21196);
and U22556 (N_22556,N_21404,N_21135);
and U22557 (N_22557,N_21828,N_21012);
xnor U22558 (N_22558,N_21579,N_21154);
xnor U22559 (N_22559,N_21641,N_21986);
nor U22560 (N_22560,N_21542,N_21927);
xnor U22561 (N_22561,N_21687,N_21806);
xnor U22562 (N_22562,N_21805,N_21204);
and U22563 (N_22563,N_21337,N_21460);
nand U22564 (N_22564,N_21873,N_21518);
and U22565 (N_22565,N_21494,N_21926);
or U22566 (N_22566,N_21300,N_21609);
xnor U22567 (N_22567,N_21535,N_21453);
nand U22568 (N_22568,N_21155,N_21833);
nor U22569 (N_22569,N_21304,N_21521);
nor U22570 (N_22570,N_21799,N_21220);
and U22571 (N_22571,N_21861,N_21541);
nor U22572 (N_22572,N_21570,N_21432);
nand U22573 (N_22573,N_21490,N_21804);
xor U22574 (N_22574,N_21466,N_21875);
or U22575 (N_22575,N_21635,N_21049);
xor U22576 (N_22576,N_21932,N_21359);
and U22577 (N_22577,N_21264,N_21667);
and U22578 (N_22578,N_21840,N_21206);
or U22579 (N_22579,N_21999,N_21495);
or U22580 (N_22580,N_21977,N_21245);
or U22581 (N_22581,N_21487,N_21901);
nor U22582 (N_22582,N_21935,N_21233);
nand U22583 (N_22583,N_21619,N_21949);
and U22584 (N_22584,N_21756,N_21484);
and U22585 (N_22585,N_21821,N_21878);
nor U22586 (N_22586,N_21999,N_21275);
nand U22587 (N_22587,N_21551,N_21655);
and U22588 (N_22588,N_21833,N_21283);
nor U22589 (N_22589,N_21478,N_21858);
and U22590 (N_22590,N_21533,N_21257);
nor U22591 (N_22591,N_21355,N_21572);
and U22592 (N_22592,N_21135,N_21582);
and U22593 (N_22593,N_21425,N_21056);
nand U22594 (N_22594,N_21924,N_21677);
and U22595 (N_22595,N_21947,N_21365);
xnor U22596 (N_22596,N_21207,N_21655);
and U22597 (N_22597,N_21076,N_21700);
xor U22598 (N_22598,N_21232,N_21717);
or U22599 (N_22599,N_21611,N_21001);
and U22600 (N_22600,N_21016,N_21270);
and U22601 (N_22601,N_21313,N_21884);
xnor U22602 (N_22602,N_21849,N_21829);
or U22603 (N_22603,N_21795,N_21564);
or U22604 (N_22604,N_21328,N_21470);
or U22605 (N_22605,N_21277,N_21571);
nor U22606 (N_22606,N_21995,N_21812);
or U22607 (N_22607,N_21353,N_21319);
xnor U22608 (N_22608,N_21421,N_21970);
xnor U22609 (N_22609,N_21972,N_21299);
nand U22610 (N_22610,N_21448,N_21023);
or U22611 (N_22611,N_21896,N_21324);
or U22612 (N_22612,N_21153,N_21105);
nor U22613 (N_22613,N_21963,N_21339);
or U22614 (N_22614,N_21406,N_21137);
nor U22615 (N_22615,N_21609,N_21504);
nor U22616 (N_22616,N_21254,N_21317);
xnor U22617 (N_22617,N_21714,N_21770);
xor U22618 (N_22618,N_21688,N_21972);
nor U22619 (N_22619,N_21083,N_21165);
nand U22620 (N_22620,N_21244,N_21304);
xnor U22621 (N_22621,N_21751,N_21259);
nor U22622 (N_22622,N_21778,N_21470);
nor U22623 (N_22623,N_21812,N_21754);
and U22624 (N_22624,N_21455,N_21811);
xor U22625 (N_22625,N_21579,N_21278);
or U22626 (N_22626,N_21224,N_21649);
and U22627 (N_22627,N_21548,N_21756);
or U22628 (N_22628,N_21868,N_21173);
nor U22629 (N_22629,N_21322,N_21633);
nor U22630 (N_22630,N_21064,N_21496);
nor U22631 (N_22631,N_21046,N_21280);
or U22632 (N_22632,N_21088,N_21391);
nor U22633 (N_22633,N_21488,N_21832);
nand U22634 (N_22634,N_21254,N_21301);
nor U22635 (N_22635,N_21160,N_21262);
nor U22636 (N_22636,N_21463,N_21749);
nor U22637 (N_22637,N_21459,N_21314);
nand U22638 (N_22638,N_21815,N_21685);
and U22639 (N_22639,N_21830,N_21027);
xnor U22640 (N_22640,N_21821,N_21057);
and U22641 (N_22641,N_21667,N_21049);
nor U22642 (N_22642,N_21041,N_21252);
nand U22643 (N_22643,N_21313,N_21845);
and U22644 (N_22644,N_21453,N_21331);
or U22645 (N_22645,N_21690,N_21891);
nor U22646 (N_22646,N_21458,N_21009);
nor U22647 (N_22647,N_21069,N_21810);
nand U22648 (N_22648,N_21928,N_21599);
and U22649 (N_22649,N_21464,N_21651);
and U22650 (N_22650,N_21383,N_21573);
nor U22651 (N_22651,N_21742,N_21893);
nor U22652 (N_22652,N_21560,N_21783);
nor U22653 (N_22653,N_21311,N_21858);
nor U22654 (N_22654,N_21290,N_21768);
nand U22655 (N_22655,N_21810,N_21771);
xor U22656 (N_22656,N_21414,N_21738);
xnor U22657 (N_22657,N_21244,N_21825);
or U22658 (N_22658,N_21585,N_21523);
and U22659 (N_22659,N_21555,N_21326);
or U22660 (N_22660,N_21788,N_21164);
nor U22661 (N_22661,N_21623,N_21694);
or U22662 (N_22662,N_21469,N_21307);
or U22663 (N_22663,N_21065,N_21975);
or U22664 (N_22664,N_21300,N_21227);
xnor U22665 (N_22665,N_21283,N_21151);
or U22666 (N_22666,N_21069,N_21731);
or U22667 (N_22667,N_21695,N_21799);
and U22668 (N_22668,N_21816,N_21736);
or U22669 (N_22669,N_21347,N_21133);
and U22670 (N_22670,N_21651,N_21242);
nand U22671 (N_22671,N_21861,N_21527);
or U22672 (N_22672,N_21200,N_21842);
nor U22673 (N_22673,N_21075,N_21993);
xor U22674 (N_22674,N_21472,N_21808);
xor U22675 (N_22675,N_21022,N_21639);
nand U22676 (N_22676,N_21622,N_21031);
or U22677 (N_22677,N_21819,N_21296);
and U22678 (N_22678,N_21787,N_21620);
nand U22679 (N_22679,N_21771,N_21676);
nor U22680 (N_22680,N_21453,N_21602);
nor U22681 (N_22681,N_21875,N_21258);
or U22682 (N_22682,N_21228,N_21354);
or U22683 (N_22683,N_21434,N_21558);
nand U22684 (N_22684,N_21747,N_21239);
and U22685 (N_22685,N_21326,N_21911);
or U22686 (N_22686,N_21113,N_21570);
nor U22687 (N_22687,N_21928,N_21651);
xor U22688 (N_22688,N_21824,N_21790);
nor U22689 (N_22689,N_21750,N_21385);
xnor U22690 (N_22690,N_21352,N_21524);
xnor U22691 (N_22691,N_21604,N_21502);
xnor U22692 (N_22692,N_21690,N_21403);
nand U22693 (N_22693,N_21206,N_21997);
nand U22694 (N_22694,N_21792,N_21676);
xor U22695 (N_22695,N_21805,N_21495);
nand U22696 (N_22696,N_21501,N_21226);
nand U22697 (N_22697,N_21260,N_21057);
nand U22698 (N_22698,N_21881,N_21218);
xnor U22699 (N_22699,N_21329,N_21134);
xnor U22700 (N_22700,N_21283,N_21499);
xor U22701 (N_22701,N_21349,N_21789);
nand U22702 (N_22702,N_21253,N_21615);
nor U22703 (N_22703,N_21702,N_21168);
or U22704 (N_22704,N_21548,N_21653);
nor U22705 (N_22705,N_21384,N_21156);
xnor U22706 (N_22706,N_21275,N_21549);
xor U22707 (N_22707,N_21789,N_21724);
nand U22708 (N_22708,N_21363,N_21015);
nor U22709 (N_22709,N_21917,N_21628);
nor U22710 (N_22710,N_21400,N_21045);
and U22711 (N_22711,N_21046,N_21761);
and U22712 (N_22712,N_21978,N_21673);
xnor U22713 (N_22713,N_21812,N_21885);
or U22714 (N_22714,N_21405,N_21233);
xor U22715 (N_22715,N_21953,N_21250);
xnor U22716 (N_22716,N_21450,N_21542);
nor U22717 (N_22717,N_21348,N_21606);
nand U22718 (N_22718,N_21743,N_21837);
or U22719 (N_22719,N_21246,N_21110);
nand U22720 (N_22720,N_21588,N_21266);
nand U22721 (N_22721,N_21923,N_21056);
xor U22722 (N_22722,N_21193,N_21168);
nor U22723 (N_22723,N_21434,N_21342);
and U22724 (N_22724,N_21779,N_21018);
or U22725 (N_22725,N_21428,N_21451);
nand U22726 (N_22726,N_21901,N_21678);
and U22727 (N_22727,N_21602,N_21997);
nor U22728 (N_22728,N_21004,N_21897);
or U22729 (N_22729,N_21473,N_21866);
nand U22730 (N_22730,N_21455,N_21479);
nand U22731 (N_22731,N_21516,N_21101);
xnor U22732 (N_22732,N_21484,N_21026);
nor U22733 (N_22733,N_21675,N_21273);
and U22734 (N_22734,N_21533,N_21730);
or U22735 (N_22735,N_21947,N_21501);
or U22736 (N_22736,N_21464,N_21188);
nand U22737 (N_22737,N_21226,N_21920);
nand U22738 (N_22738,N_21158,N_21997);
nand U22739 (N_22739,N_21059,N_21537);
nor U22740 (N_22740,N_21753,N_21143);
xnor U22741 (N_22741,N_21759,N_21371);
or U22742 (N_22742,N_21800,N_21518);
and U22743 (N_22743,N_21840,N_21482);
and U22744 (N_22744,N_21886,N_21426);
and U22745 (N_22745,N_21807,N_21962);
nor U22746 (N_22746,N_21655,N_21886);
xnor U22747 (N_22747,N_21002,N_21798);
xor U22748 (N_22748,N_21647,N_21686);
or U22749 (N_22749,N_21545,N_21078);
xor U22750 (N_22750,N_21281,N_21555);
nor U22751 (N_22751,N_21861,N_21202);
or U22752 (N_22752,N_21233,N_21396);
xnor U22753 (N_22753,N_21579,N_21845);
or U22754 (N_22754,N_21828,N_21968);
xnor U22755 (N_22755,N_21440,N_21668);
or U22756 (N_22756,N_21528,N_21580);
nor U22757 (N_22757,N_21029,N_21596);
xnor U22758 (N_22758,N_21491,N_21336);
or U22759 (N_22759,N_21411,N_21312);
nand U22760 (N_22760,N_21813,N_21916);
xnor U22761 (N_22761,N_21437,N_21681);
or U22762 (N_22762,N_21033,N_21572);
nand U22763 (N_22763,N_21449,N_21922);
or U22764 (N_22764,N_21785,N_21660);
nand U22765 (N_22765,N_21861,N_21935);
or U22766 (N_22766,N_21711,N_21505);
and U22767 (N_22767,N_21763,N_21176);
xnor U22768 (N_22768,N_21049,N_21763);
nor U22769 (N_22769,N_21458,N_21383);
xnor U22770 (N_22770,N_21745,N_21608);
or U22771 (N_22771,N_21988,N_21217);
or U22772 (N_22772,N_21329,N_21288);
xor U22773 (N_22773,N_21227,N_21100);
nand U22774 (N_22774,N_21621,N_21367);
or U22775 (N_22775,N_21084,N_21388);
or U22776 (N_22776,N_21659,N_21725);
or U22777 (N_22777,N_21039,N_21093);
xor U22778 (N_22778,N_21318,N_21383);
or U22779 (N_22779,N_21933,N_21818);
nor U22780 (N_22780,N_21906,N_21186);
nor U22781 (N_22781,N_21715,N_21388);
or U22782 (N_22782,N_21047,N_21552);
nor U22783 (N_22783,N_21887,N_21415);
or U22784 (N_22784,N_21722,N_21086);
nor U22785 (N_22785,N_21757,N_21939);
nand U22786 (N_22786,N_21827,N_21499);
xnor U22787 (N_22787,N_21710,N_21202);
or U22788 (N_22788,N_21470,N_21627);
or U22789 (N_22789,N_21462,N_21781);
nand U22790 (N_22790,N_21163,N_21608);
nor U22791 (N_22791,N_21255,N_21753);
nor U22792 (N_22792,N_21068,N_21240);
and U22793 (N_22793,N_21081,N_21833);
and U22794 (N_22794,N_21936,N_21180);
xor U22795 (N_22795,N_21610,N_21294);
nand U22796 (N_22796,N_21094,N_21268);
or U22797 (N_22797,N_21169,N_21115);
xor U22798 (N_22798,N_21142,N_21846);
nand U22799 (N_22799,N_21594,N_21504);
nand U22800 (N_22800,N_21698,N_21107);
nor U22801 (N_22801,N_21529,N_21178);
and U22802 (N_22802,N_21523,N_21161);
and U22803 (N_22803,N_21003,N_21609);
or U22804 (N_22804,N_21990,N_21420);
nor U22805 (N_22805,N_21551,N_21366);
and U22806 (N_22806,N_21311,N_21999);
nor U22807 (N_22807,N_21504,N_21064);
xnor U22808 (N_22808,N_21231,N_21568);
and U22809 (N_22809,N_21765,N_21591);
nor U22810 (N_22810,N_21384,N_21798);
xor U22811 (N_22811,N_21949,N_21825);
xor U22812 (N_22812,N_21749,N_21335);
nor U22813 (N_22813,N_21613,N_21264);
and U22814 (N_22814,N_21160,N_21650);
nand U22815 (N_22815,N_21260,N_21550);
xor U22816 (N_22816,N_21437,N_21754);
and U22817 (N_22817,N_21133,N_21470);
or U22818 (N_22818,N_21070,N_21793);
nand U22819 (N_22819,N_21711,N_21166);
nand U22820 (N_22820,N_21983,N_21724);
nand U22821 (N_22821,N_21789,N_21058);
nor U22822 (N_22822,N_21006,N_21204);
nand U22823 (N_22823,N_21463,N_21736);
nor U22824 (N_22824,N_21378,N_21050);
and U22825 (N_22825,N_21445,N_21848);
nand U22826 (N_22826,N_21041,N_21049);
nor U22827 (N_22827,N_21017,N_21340);
xnor U22828 (N_22828,N_21729,N_21696);
xnor U22829 (N_22829,N_21369,N_21901);
nor U22830 (N_22830,N_21747,N_21305);
and U22831 (N_22831,N_21046,N_21419);
nor U22832 (N_22832,N_21672,N_21548);
nand U22833 (N_22833,N_21729,N_21752);
nand U22834 (N_22834,N_21125,N_21251);
nand U22835 (N_22835,N_21438,N_21328);
nor U22836 (N_22836,N_21477,N_21942);
and U22837 (N_22837,N_21125,N_21561);
xnor U22838 (N_22838,N_21139,N_21456);
or U22839 (N_22839,N_21254,N_21753);
or U22840 (N_22840,N_21403,N_21496);
and U22841 (N_22841,N_21520,N_21850);
xnor U22842 (N_22842,N_21868,N_21822);
nand U22843 (N_22843,N_21294,N_21912);
and U22844 (N_22844,N_21667,N_21113);
xnor U22845 (N_22845,N_21017,N_21468);
and U22846 (N_22846,N_21465,N_21859);
nor U22847 (N_22847,N_21774,N_21919);
xnor U22848 (N_22848,N_21610,N_21469);
and U22849 (N_22849,N_21270,N_21584);
xor U22850 (N_22850,N_21616,N_21045);
xor U22851 (N_22851,N_21713,N_21280);
or U22852 (N_22852,N_21630,N_21743);
xnor U22853 (N_22853,N_21323,N_21017);
and U22854 (N_22854,N_21053,N_21098);
or U22855 (N_22855,N_21449,N_21161);
or U22856 (N_22856,N_21356,N_21016);
xor U22857 (N_22857,N_21654,N_21165);
or U22858 (N_22858,N_21961,N_21121);
nor U22859 (N_22859,N_21225,N_21891);
or U22860 (N_22860,N_21996,N_21063);
nand U22861 (N_22861,N_21404,N_21641);
nor U22862 (N_22862,N_21408,N_21738);
or U22863 (N_22863,N_21706,N_21033);
and U22864 (N_22864,N_21241,N_21048);
and U22865 (N_22865,N_21278,N_21470);
or U22866 (N_22866,N_21221,N_21299);
nand U22867 (N_22867,N_21251,N_21626);
or U22868 (N_22868,N_21530,N_21148);
and U22869 (N_22869,N_21738,N_21016);
or U22870 (N_22870,N_21900,N_21726);
xor U22871 (N_22871,N_21020,N_21259);
nor U22872 (N_22872,N_21512,N_21684);
or U22873 (N_22873,N_21888,N_21619);
nor U22874 (N_22874,N_21387,N_21909);
xnor U22875 (N_22875,N_21658,N_21772);
xor U22876 (N_22876,N_21152,N_21836);
and U22877 (N_22877,N_21267,N_21925);
xor U22878 (N_22878,N_21241,N_21315);
and U22879 (N_22879,N_21139,N_21386);
or U22880 (N_22880,N_21563,N_21194);
xor U22881 (N_22881,N_21696,N_21454);
xor U22882 (N_22882,N_21393,N_21355);
nor U22883 (N_22883,N_21011,N_21582);
xor U22884 (N_22884,N_21875,N_21452);
nand U22885 (N_22885,N_21612,N_21407);
xor U22886 (N_22886,N_21479,N_21407);
or U22887 (N_22887,N_21297,N_21800);
xor U22888 (N_22888,N_21467,N_21237);
and U22889 (N_22889,N_21249,N_21710);
or U22890 (N_22890,N_21325,N_21817);
and U22891 (N_22891,N_21121,N_21753);
or U22892 (N_22892,N_21893,N_21251);
nand U22893 (N_22893,N_21692,N_21048);
nor U22894 (N_22894,N_21985,N_21889);
or U22895 (N_22895,N_21577,N_21486);
nand U22896 (N_22896,N_21534,N_21799);
nor U22897 (N_22897,N_21383,N_21496);
nand U22898 (N_22898,N_21472,N_21278);
xor U22899 (N_22899,N_21671,N_21527);
and U22900 (N_22900,N_21601,N_21796);
nand U22901 (N_22901,N_21051,N_21324);
nor U22902 (N_22902,N_21209,N_21720);
nand U22903 (N_22903,N_21322,N_21464);
xnor U22904 (N_22904,N_21147,N_21739);
or U22905 (N_22905,N_21800,N_21954);
or U22906 (N_22906,N_21012,N_21358);
or U22907 (N_22907,N_21197,N_21700);
or U22908 (N_22908,N_21005,N_21811);
nor U22909 (N_22909,N_21970,N_21904);
xor U22910 (N_22910,N_21317,N_21664);
and U22911 (N_22911,N_21592,N_21813);
and U22912 (N_22912,N_21361,N_21956);
nand U22913 (N_22913,N_21717,N_21414);
nand U22914 (N_22914,N_21812,N_21524);
nand U22915 (N_22915,N_21947,N_21509);
or U22916 (N_22916,N_21094,N_21354);
nor U22917 (N_22917,N_21637,N_21811);
nand U22918 (N_22918,N_21409,N_21994);
nand U22919 (N_22919,N_21881,N_21550);
nor U22920 (N_22920,N_21614,N_21459);
and U22921 (N_22921,N_21436,N_21304);
and U22922 (N_22922,N_21572,N_21815);
or U22923 (N_22923,N_21394,N_21304);
xor U22924 (N_22924,N_21125,N_21461);
and U22925 (N_22925,N_21351,N_21135);
and U22926 (N_22926,N_21193,N_21106);
or U22927 (N_22927,N_21899,N_21433);
or U22928 (N_22928,N_21554,N_21066);
xor U22929 (N_22929,N_21261,N_21044);
nor U22930 (N_22930,N_21413,N_21906);
and U22931 (N_22931,N_21697,N_21101);
nand U22932 (N_22932,N_21924,N_21703);
or U22933 (N_22933,N_21708,N_21787);
xor U22934 (N_22934,N_21833,N_21131);
and U22935 (N_22935,N_21384,N_21891);
nor U22936 (N_22936,N_21177,N_21018);
nor U22937 (N_22937,N_21689,N_21755);
and U22938 (N_22938,N_21416,N_21364);
xor U22939 (N_22939,N_21276,N_21805);
xor U22940 (N_22940,N_21691,N_21402);
xnor U22941 (N_22941,N_21625,N_21193);
and U22942 (N_22942,N_21634,N_21076);
xnor U22943 (N_22943,N_21545,N_21921);
nor U22944 (N_22944,N_21397,N_21394);
and U22945 (N_22945,N_21180,N_21645);
nand U22946 (N_22946,N_21669,N_21289);
xor U22947 (N_22947,N_21384,N_21052);
and U22948 (N_22948,N_21525,N_21506);
nor U22949 (N_22949,N_21761,N_21844);
or U22950 (N_22950,N_21548,N_21691);
xor U22951 (N_22951,N_21710,N_21550);
or U22952 (N_22952,N_21917,N_21835);
nand U22953 (N_22953,N_21033,N_21839);
and U22954 (N_22954,N_21154,N_21176);
and U22955 (N_22955,N_21071,N_21420);
nand U22956 (N_22956,N_21135,N_21596);
and U22957 (N_22957,N_21475,N_21553);
or U22958 (N_22958,N_21052,N_21904);
xor U22959 (N_22959,N_21975,N_21490);
nand U22960 (N_22960,N_21845,N_21473);
nand U22961 (N_22961,N_21961,N_21650);
nand U22962 (N_22962,N_21499,N_21293);
and U22963 (N_22963,N_21799,N_21283);
xnor U22964 (N_22964,N_21891,N_21450);
nor U22965 (N_22965,N_21370,N_21138);
and U22966 (N_22966,N_21365,N_21470);
nand U22967 (N_22967,N_21159,N_21620);
or U22968 (N_22968,N_21741,N_21034);
nor U22969 (N_22969,N_21378,N_21076);
or U22970 (N_22970,N_21505,N_21431);
nor U22971 (N_22971,N_21585,N_21127);
xor U22972 (N_22972,N_21038,N_21874);
and U22973 (N_22973,N_21199,N_21676);
nand U22974 (N_22974,N_21343,N_21077);
xnor U22975 (N_22975,N_21649,N_21351);
nand U22976 (N_22976,N_21754,N_21304);
nor U22977 (N_22977,N_21927,N_21915);
or U22978 (N_22978,N_21877,N_21125);
or U22979 (N_22979,N_21863,N_21970);
and U22980 (N_22980,N_21074,N_21725);
or U22981 (N_22981,N_21307,N_21554);
and U22982 (N_22982,N_21756,N_21626);
xor U22983 (N_22983,N_21899,N_21127);
nor U22984 (N_22984,N_21841,N_21373);
and U22985 (N_22985,N_21280,N_21213);
xor U22986 (N_22986,N_21374,N_21051);
nand U22987 (N_22987,N_21604,N_21925);
xor U22988 (N_22988,N_21742,N_21206);
nand U22989 (N_22989,N_21293,N_21861);
nand U22990 (N_22990,N_21596,N_21449);
nand U22991 (N_22991,N_21621,N_21208);
nand U22992 (N_22992,N_21534,N_21225);
nand U22993 (N_22993,N_21225,N_21447);
nand U22994 (N_22994,N_21864,N_21610);
xnor U22995 (N_22995,N_21738,N_21936);
xor U22996 (N_22996,N_21070,N_21903);
and U22997 (N_22997,N_21414,N_21528);
nand U22998 (N_22998,N_21176,N_21224);
nand U22999 (N_22999,N_21031,N_21672);
nand U23000 (N_23000,N_22460,N_22236);
nand U23001 (N_23001,N_22938,N_22175);
nand U23002 (N_23002,N_22441,N_22385);
xnor U23003 (N_23003,N_22398,N_22926);
or U23004 (N_23004,N_22307,N_22140);
and U23005 (N_23005,N_22717,N_22509);
and U23006 (N_23006,N_22574,N_22208);
xnor U23007 (N_23007,N_22279,N_22686);
nand U23008 (N_23008,N_22377,N_22586);
or U23009 (N_23009,N_22751,N_22759);
or U23010 (N_23010,N_22654,N_22418);
xnor U23011 (N_23011,N_22263,N_22795);
nor U23012 (N_23012,N_22476,N_22810);
and U23013 (N_23013,N_22115,N_22295);
xnor U23014 (N_23014,N_22281,N_22419);
or U23015 (N_23015,N_22846,N_22044);
nand U23016 (N_23016,N_22904,N_22943);
xnor U23017 (N_23017,N_22864,N_22312);
and U23018 (N_23018,N_22134,N_22556);
nand U23019 (N_23019,N_22318,N_22296);
nor U23020 (N_23020,N_22786,N_22611);
nor U23021 (N_23021,N_22701,N_22257);
nor U23022 (N_23022,N_22655,N_22600);
nand U23023 (N_23023,N_22968,N_22821);
and U23024 (N_23024,N_22889,N_22231);
nor U23025 (N_23025,N_22573,N_22401);
nor U23026 (N_23026,N_22760,N_22414);
or U23027 (N_23027,N_22519,N_22400);
and U23028 (N_23028,N_22188,N_22748);
or U23029 (N_23029,N_22100,N_22771);
xor U23030 (N_23030,N_22709,N_22205);
or U23031 (N_23031,N_22011,N_22851);
or U23032 (N_23032,N_22526,N_22841);
xor U23033 (N_23033,N_22991,N_22733);
nand U23034 (N_23034,N_22110,N_22329);
nor U23035 (N_23035,N_22156,N_22308);
and U23036 (N_23036,N_22314,N_22206);
nand U23037 (N_23037,N_22497,N_22054);
and U23038 (N_23038,N_22708,N_22066);
nor U23039 (N_23039,N_22085,N_22446);
xor U23040 (N_23040,N_22320,N_22478);
nand U23041 (N_23041,N_22728,N_22641);
and U23042 (N_23042,N_22808,N_22809);
nor U23043 (N_23043,N_22690,N_22051);
or U23044 (N_23044,N_22700,N_22982);
and U23045 (N_23045,N_22038,N_22812);
xor U23046 (N_23046,N_22373,N_22958);
and U23047 (N_23047,N_22006,N_22094);
or U23048 (N_23048,N_22456,N_22683);
and U23049 (N_23049,N_22029,N_22592);
xor U23050 (N_23050,N_22356,N_22956);
nand U23051 (N_23051,N_22921,N_22613);
and U23052 (N_23052,N_22363,N_22089);
xor U23053 (N_23053,N_22661,N_22726);
nand U23054 (N_23054,N_22932,N_22033);
or U23055 (N_23055,N_22510,N_22292);
nand U23056 (N_23056,N_22560,N_22002);
or U23057 (N_23057,N_22822,N_22407);
and U23058 (N_23058,N_22855,N_22170);
nand U23059 (N_23059,N_22537,N_22350);
xor U23060 (N_23060,N_22805,N_22757);
xnor U23061 (N_23061,N_22157,N_22668);
xnor U23062 (N_23062,N_22250,N_22025);
xnor U23063 (N_23063,N_22732,N_22463);
xnor U23064 (N_23064,N_22590,N_22234);
nand U23065 (N_23065,N_22343,N_22713);
nand U23066 (N_23066,N_22610,N_22857);
nor U23067 (N_23067,N_22939,N_22685);
xor U23068 (N_23068,N_22076,N_22505);
or U23069 (N_23069,N_22397,N_22238);
nand U23070 (N_23070,N_22702,N_22266);
xnor U23071 (N_23071,N_22918,N_22435);
or U23072 (N_23072,N_22718,N_22079);
nor U23073 (N_23073,N_22313,N_22890);
nor U23074 (N_23074,N_22642,N_22349);
and U23075 (N_23075,N_22167,N_22545);
nand U23076 (N_23076,N_22255,N_22549);
nand U23077 (N_23077,N_22133,N_22737);
or U23078 (N_23078,N_22269,N_22354);
or U23079 (N_23079,N_22249,N_22622);
nand U23080 (N_23080,N_22251,N_22597);
or U23081 (N_23081,N_22352,N_22226);
nor U23082 (N_23082,N_22376,N_22301);
nand U23083 (N_23083,N_22430,N_22983);
nor U23084 (N_23084,N_22372,N_22587);
nor U23085 (N_23085,N_22999,N_22146);
nand U23086 (N_23086,N_22950,N_22941);
nor U23087 (N_23087,N_22520,N_22826);
nand U23088 (N_23088,N_22962,N_22863);
or U23089 (N_23089,N_22384,N_22707);
nor U23090 (N_23090,N_22436,N_22780);
and U23091 (N_23091,N_22224,N_22288);
or U23092 (N_23092,N_22050,N_22582);
nor U23093 (N_23093,N_22432,N_22862);
and U23094 (N_23094,N_22525,N_22636);
nand U23095 (N_23095,N_22274,N_22694);
or U23096 (N_23096,N_22619,N_22210);
nand U23097 (N_23097,N_22114,N_22498);
or U23098 (N_23098,N_22504,N_22843);
or U23099 (N_23099,N_22433,N_22179);
nor U23100 (N_23100,N_22811,N_22682);
or U23101 (N_23101,N_22596,N_22163);
nand U23102 (N_23102,N_22286,N_22328);
nor U23103 (N_23103,N_22754,N_22945);
and U23104 (N_23104,N_22989,N_22070);
nand U23105 (N_23105,N_22413,N_22680);
and U23106 (N_23106,N_22217,N_22866);
nand U23107 (N_23107,N_22098,N_22792);
nor U23108 (N_23108,N_22230,N_22233);
nor U23109 (N_23109,N_22874,N_22987);
and U23110 (N_23110,N_22067,N_22566);
nand U23111 (N_23111,N_22145,N_22727);
xor U23112 (N_23112,N_22333,N_22053);
nand U23113 (N_23113,N_22192,N_22195);
xor U23114 (N_23114,N_22532,N_22039);
and U23115 (N_23115,N_22720,N_22593);
or U23116 (N_23116,N_22062,N_22302);
nand U23117 (N_23117,N_22201,N_22896);
or U23118 (N_23118,N_22045,N_22993);
and U23119 (N_23119,N_22297,N_22577);
and U23120 (N_23120,N_22036,N_22640);
and U23121 (N_23121,N_22730,N_22305);
xor U23122 (N_23122,N_22187,N_22180);
nand U23123 (N_23123,N_22660,N_22511);
nand U23124 (N_23124,N_22567,N_22755);
or U23125 (N_23125,N_22130,N_22850);
or U23126 (N_23126,N_22774,N_22239);
nand U23127 (N_23127,N_22341,N_22802);
or U23128 (N_23128,N_22023,N_22469);
nor U23129 (N_23129,N_22174,N_22221);
nor U23130 (N_23130,N_22309,N_22304);
nor U23131 (N_23131,N_22834,N_22182);
and U23132 (N_23132,N_22193,N_22656);
xnor U23133 (N_23133,N_22606,N_22670);
nand U23134 (N_23134,N_22688,N_22824);
nand U23135 (N_23135,N_22220,N_22643);
and U23136 (N_23136,N_22876,N_22366);
nor U23137 (N_23137,N_22798,N_22598);
and U23138 (N_23138,N_22984,N_22061);
nor U23139 (N_23139,N_22064,N_22589);
or U23140 (N_23140,N_22796,N_22458);
xnor U23141 (N_23141,N_22628,N_22813);
or U23142 (N_23142,N_22514,N_22695);
or U23143 (N_23143,N_22554,N_22471);
xor U23144 (N_23144,N_22770,N_22767);
nand U23145 (N_23145,N_22595,N_22340);
nor U23146 (N_23146,N_22937,N_22990);
nor U23147 (N_23147,N_22823,N_22629);
nor U23148 (N_23148,N_22369,N_22888);
nor U23149 (N_23149,N_22922,N_22090);
and U23150 (N_23150,N_22472,N_22247);
nand U23151 (N_23151,N_22368,N_22576);
nor U23152 (N_23152,N_22764,N_22900);
and U23153 (N_23153,N_22522,N_22513);
and U23154 (N_23154,N_22898,N_22048);
nand U23155 (N_23155,N_22042,N_22976);
xnor U23156 (N_23156,N_22164,N_22957);
or U23157 (N_23157,N_22552,N_22705);
nand U23158 (N_23158,N_22691,N_22998);
and U23159 (N_23159,N_22992,N_22663);
xor U23160 (N_23160,N_22000,N_22551);
or U23161 (N_23161,N_22365,N_22158);
xnor U23162 (N_23162,N_22814,N_22410);
xnor U23163 (N_23163,N_22283,N_22264);
nor U23164 (N_23164,N_22734,N_22262);
xnor U23165 (N_23165,N_22388,N_22014);
nand U23166 (N_23166,N_22944,N_22789);
xor U23167 (N_23167,N_22781,N_22964);
or U23168 (N_23168,N_22417,N_22241);
and U23169 (N_23169,N_22583,N_22387);
and U23170 (N_23170,N_22666,N_22785);
nor U23171 (N_23171,N_22126,N_22801);
and U23172 (N_23172,N_22607,N_22121);
or U23173 (N_23173,N_22165,N_22972);
nor U23174 (N_23174,N_22246,N_22731);
or U23175 (N_23175,N_22591,N_22617);
xor U23176 (N_23176,N_22651,N_22844);
xnor U23177 (N_23177,N_22920,N_22563);
nand U23178 (N_23178,N_22854,N_22547);
and U23179 (N_23179,N_22815,N_22123);
and U23180 (N_23180,N_22111,N_22877);
and U23181 (N_23181,N_22893,N_22750);
or U23182 (N_23182,N_22203,N_22016);
or U23183 (N_23183,N_22390,N_22829);
nand U23184 (N_23184,N_22049,N_22151);
nor U23185 (N_23185,N_22618,N_22060);
and U23186 (N_23186,N_22806,N_22621);
or U23187 (N_23187,N_22746,N_22449);
or U23188 (N_23188,N_22706,N_22996);
nand U23189 (N_23189,N_22544,N_22259);
nand U23190 (N_23190,N_22367,N_22847);
or U23191 (N_23191,N_22323,N_22970);
nand U23192 (N_23192,N_22204,N_22040);
nand U23193 (N_23193,N_22483,N_22882);
nor U23194 (N_23194,N_22773,N_22183);
xor U23195 (N_23195,N_22873,N_22612);
nor U23196 (N_23196,N_22927,N_22104);
and U23197 (N_23197,N_22625,N_22272);
xnor U23198 (N_23198,N_22946,N_22459);
or U23199 (N_23199,N_22742,N_22389);
nor U23200 (N_23200,N_22059,N_22434);
and U23201 (N_23201,N_22977,N_22645);
nor U23202 (N_23202,N_22819,N_22339);
xnor U23203 (N_23203,N_22176,N_22171);
and U23204 (N_23204,N_22845,N_22277);
nand U23205 (N_23205,N_22797,N_22495);
nor U23206 (N_23206,N_22561,N_22298);
nand U23207 (N_23207,N_22777,N_22490);
or U23208 (N_23208,N_22667,N_22258);
xor U23209 (N_23209,N_22923,N_22428);
nand U23210 (N_23210,N_22093,N_22268);
xnor U23211 (N_23211,N_22639,N_22679);
or U23212 (N_23212,N_22934,N_22530);
or U23213 (N_23213,N_22485,N_22744);
or U23214 (N_23214,N_22959,N_22697);
or U23215 (N_23215,N_22482,N_22055);
and U23216 (N_23216,N_22256,N_22439);
nand U23217 (N_23217,N_22539,N_22335);
or U23218 (N_23218,N_22191,N_22570);
xnor U23219 (N_23219,N_22300,N_22196);
xor U23220 (N_23220,N_22528,N_22886);
xnor U23221 (N_23221,N_22396,N_22883);
or U23222 (N_23222,N_22803,N_22360);
nand U23223 (N_23223,N_22658,N_22383);
nand U23224 (N_23224,N_22440,N_22173);
xor U23225 (N_23225,N_22327,N_22101);
nor U23226 (N_23226,N_22020,N_22738);
nor U23227 (N_23227,N_22106,N_22536);
and U23228 (N_23228,N_22800,N_22034);
xnor U23229 (N_23229,N_22316,N_22672);
nand U23230 (N_23230,N_22955,N_22649);
or U23231 (N_23231,N_22489,N_22132);
nor U23232 (N_23232,N_22169,N_22491);
nand U23233 (N_23233,N_22626,N_22779);
nor U23234 (N_23234,N_22588,N_22310);
nor U23235 (N_23235,N_22897,N_22077);
nor U23236 (N_23236,N_22065,N_22529);
nand U23237 (N_23237,N_22159,N_22144);
or U23238 (N_23238,N_22963,N_22985);
and U23239 (N_23239,N_22075,N_22739);
xnor U23240 (N_23240,N_22382,N_22531);
xor U23241 (N_23241,N_22185,N_22475);
or U23242 (N_23242,N_22931,N_22161);
xnor U23243 (N_23243,N_22899,N_22867);
xnor U23244 (N_23244,N_22892,N_22839);
xor U23245 (N_23245,N_22571,N_22411);
nand U23246 (N_23246,N_22409,N_22102);
nor U23247 (N_23247,N_22326,N_22222);
and U23248 (N_23248,N_22580,N_22517);
and U23249 (N_23249,N_22692,N_22481);
or U23250 (N_23250,N_22008,N_22166);
xnor U23251 (N_23251,N_22515,N_22142);
or U23252 (N_23252,N_22860,N_22758);
nand U23253 (N_23253,N_22568,N_22056);
nand U23254 (N_23254,N_22214,N_22678);
and U23255 (N_23255,N_22450,N_22153);
or U23256 (N_23256,N_22470,N_22474);
nand U23257 (N_23257,N_22452,N_22324);
nand U23258 (N_23258,N_22148,N_22558);
xnor U23259 (N_23259,N_22125,N_22858);
xnor U23260 (N_23260,N_22046,N_22729);
nand U23261 (N_23261,N_22884,N_22135);
and U23262 (N_23262,N_22951,N_22374);
or U23263 (N_23263,N_22769,N_22361);
nor U23264 (N_23264,N_22351,N_22585);
nor U23265 (N_23265,N_22437,N_22399);
nand U23266 (N_23266,N_22825,N_22914);
nand U23267 (N_23267,N_22870,N_22788);
nor U23268 (N_23268,N_22083,N_22453);
or U23269 (N_23269,N_22007,N_22724);
and U23270 (N_23270,N_22357,N_22630);
nor U23271 (N_23271,N_22448,N_22493);
xor U23272 (N_23272,N_22865,N_22548);
nand U23273 (N_23273,N_22784,N_22712);
nor U23274 (N_23274,N_22395,N_22928);
xor U23275 (N_23275,N_22451,N_22019);
or U23276 (N_23276,N_22122,N_22534);
nand U23277 (N_23277,N_22457,N_22391);
nand U23278 (N_23278,N_22464,N_22403);
nor U23279 (N_23279,N_22979,N_22186);
or U23280 (N_23280,N_22852,N_22081);
and U23281 (N_23281,N_22714,N_22917);
or U23282 (N_23282,N_22290,N_22232);
nor U23283 (N_23283,N_22035,N_22930);
and U23284 (N_23284,N_22253,N_22868);
nand U23285 (N_23285,N_22856,N_22503);
xnor U23286 (N_23286,N_22572,N_22778);
or U23287 (N_23287,N_22671,N_22026);
nor U23288 (N_23288,N_22276,N_22632);
nor U23289 (N_23289,N_22794,N_22078);
nand U23290 (N_23290,N_22325,N_22080);
or U23291 (N_23291,N_22404,N_22118);
nor U23292 (N_23292,N_22791,N_22096);
nor U23293 (N_23293,N_22355,N_22961);
nand U23294 (N_23294,N_22228,N_22753);
nand U23295 (N_23295,N_22252,N_22915);
or U23296 (N_23296,N_22669,N_22995);
nand U23297 (N_23297,N_22909,N_22512);
nor U23298 (N_23298,N_22108,N_22541);
or U23299 (N_23299,N_22480,N_22107);
or U23300 (N_23300,N_22994,N_22535);
and U23301 (N_23301,N_22675,N_22664);
nand U23302 (N_23302,N_22105,N_22074);
and U23303 (N_23303,N_22527,N_22848);
xnor U23304 (N_23304,N_22665,N_22240);
or U23305 (N_23305,N_22202,N_22068);
nor U23306 (N_23306,N_22837,N_22037);
nand U23307 (N_23307,N_22698,N_22901);
xnor U23308 (N_23308,N_22947,N_22584);
xor U23309 (N_23309,N_22386,N_22147);
and U23310 (N_23310,N_22129,N_22935);
nor U23311 (N_23311,N_22421,N_22199);
xor U23312 (N_23312,N_22141,N_22684);
xor U23313 (N_23313,N_22378,N_22562);
nand U23314 (N_23314,N_22427,N_22542);
nor U23315 (N_23315,N_22334,N_22816);
nand U23316 (N_23316,N_22523,N_22178);
and U23317 (N_23317,N_22557,N_22223);
and U23318 (N_23318,N_22971,N_22502);
nor U23319 (N_23319,N_22902,N_22818);
and U23320 (N_23320,N_22088,N_22218);
nand U23321 (N_23321,N_22879,N_22681);
or U23322 (N_23322,N_22136,N_22980);
and U23323 (N_23323,N_22337,N_22905);
nand U23324 (N_23324,N_22910,N_22124);
or U23325 (N_23325,N_22776,N_22763);
nor U23326 (N_23326,N_22948,N_22652);
and U23327 (N_23327,N_22673,N_22756);
or U23328 (N_23328,N_22689,N_22952);
nand U23329 (N_23329,N_22859,N_22315);
nand U23330 (N_23330,N_22346,N_22086);
nor U23331 (N_23331,N_22416,N_22719);
and U23332 (N_23332,N_22082,N_22913);
xor U23333 (N_23333,N_22285,N_22975);
nand U23334 (N_23334,N_22650,N_22092);
and U23335 (N_23335,N_22594,N_22782);
nand U23336 (N_23336,N_22431,N_22677);
xor U23337 (N_23337,N_22412,N_22986);
and U23338 (N_23338,N_22659,N_22321);
nand U23339 (N_23339,N_22380,N_22965);
and U23340 (N_23340,N_22209,N_22745);
and U23341 (N_23341,N_22072,N_22559);
and U23342 (N_23342,N_22775,N_22402);
and U23343 (N_23343,N_22112,N_22500);
xor U23344 (N_23344,N_22287,N_22762);
and U23345 (N_23345,N_22916,N_22332);
nor U23346 (N_23346,N_22703,N_22942);
xor U23347 (N_23347,N_22137,N_22790);
nor U23348 (N_23348,N_22393,N_22603);
xor U23349 (N_23349,N_22506,N_22735);
xor U23350 (N_23350,N_22152,N_22197);
nand U23351 (N_23351,N_22479,N_22198);
xnor U23352 (N_23352,N_22027,N_22270);
or U23353 (N_23353,N_22271,N_22827);
and U23354 (N_23354,N_22575,N_22211);
xor U23355 (N_23355,N_22408,N_22605);
and U23356 (N_23356,N_22891,N_22415);
or U23357 (N_23357,N_22336,N_22492);
nor U23358 (N_23358,N_22017,N_22954);
nand U23359 (N_23359,N_22477,N_22445);
nand U23360 (N_23360,N_22553,N_22465);
and U23361 (N_23361,N_22978,N_22229);
or U23362 (N_23362,N_22973,N_22009);
xnor U23363 (N_23363,N_22631,N_22524);
nand U23364 (N_23364,N_22265,N_22216);
nor U23365 (N_23365,N_22820,N_22189);
xor U23366 (N_23366,N_22429,N_22420);
nand U23367 (N_23367,N_22501,N_22743);
and U23368 (N_23368,N_22087,N_22494);
and U23369 (N_23369,N_22616,N_22073);
or U23370 (N_23370,N_22836,N_22364);
xnor U23371 (N_23371,N_22245,N_22496);
and U23372 (N_23372,N_22190,N_22103);
nand U23373 (N_23373,N_22127,N_22444);
xnor U23374 (N_23374,N_22725,N_22370);
nor U23375 (N_23375,N_22488,N_22338);
nand U23376 (N_23376,N_22097,N_22024);
and U23377 (N_23377,N_22172,N_22131);
xnor U23378 (N_23378,N_22261,N_22242);
or U23379 (N_23379,N_22840,N_22615);
nor U23380 (N_23380,N_22022,N_22853);
nor U23381 (N_23381,N_22306,N_22162);
nand U23382 (N_23382,N_22711,N_22828);
xnor U23383 (N_23383,N_22181,N_22212);
and U23384 (N_23384,N_22768,N_22555);
nor U23385 (N_23385,N_22284,N_22267);
and U23386 (N_23386,N_22138,N_22521);
xnor U23387 (N_23387,N_22113,N_22322);
nor U23388 (N_23388,N_22468,N_22653);
nor U23389 (N_23389,N_22215,N_22069);
or U23390 (N_23390,N_22330,N_22507);
xor U23391 (N_23391,N_22740,N_22254);
xnor U23392 (N_23392,N_22235,N_22379);
or U23393 (N_23393,N_22299,N_22752);
nand U23394 (N_23394,N_22486,N_22878);
nand U23395 (N_23395,N_22150,N_22969);
nor U23396 (N_23396,N_22154,N_22487);
nand U23397 (N_23397,N_22331,N_22273);
xor U23398 (N_23398,N_22736,N_22143);
or U23399 (N_23399,N_22359,N_22614);
and U23400 (N_23400,N_22648,N_22120);
xor U23401 (N_23401,N_22831,N_22637);
nor U23402 (N_23402,N_22516,N_22319);
xnor U23403 (N_23403,N_22581,N_22289);
nor U23404 (N_23404,N_22375,N_22084);
and U23405 (N_23405,N_22043,N_22012);
or U23406 (N_23406,N_22461,N_22005);
nand U23407 (N_23407,N_22518,N_22538);
and U23408 (N_23408,N_22194,N_22647);
nor U23409 (N_23409,N_22294,N_22721);
xor U23410 (N_23410,N_22003,N_22894);
nor U23411 (N_23411,N_22244,N_22031);
or U23412 (N_23412,N_22787,N_22508);
or U23413 (N_23413,N_22696,N_22422);
nand U23414 (N_23414,N_22392,N_22041);
and U23415 (N_23415,N_22579,N_22057);
nor U23416 (N_23416,N_22311,N_22177);
or U23417 (N_23417,N_22908,N_22071);
xor U23418 (N_23418,N_22347,N_22936);
or U23419 (N_23419,N_22010,N_22772);
xor U23420 (N_23420,N_22715,N_22747);
nand U23421 (N_23421,N_22749,N_22109);
and U23422 (N_23422,N_22499,N_22345);
nor U23423 (N_23423,N_22293,N_22869);
xnor U23424 (N_23424,N_22353,N_22063);
nor U23425 (N_23425,N_22207,N_22635);
or U23426 (N_23426,N_22966,N_22447);
nand U23427 (N_23427,N_22362,N_22912);
or U23428 (N_23428,N_22032,N_22282);
nand U23429 (N_23429,N_22633,N_22716);
nand U23430 (N_23430,N_22793,N_22213);
nand U23431 (N_23431,N_22454,N_22168);
xor U23432 (N_23432,N_22533,N_22833);
or U23433 (N_23433,N_22004,N_22644);
or U23434 (N_23434,N_22015,N_22394);
nor U23435 (N_23435,N_22885,N_22949);
nor U23436 (N_23436,N_22455,N_22624);
xnor U23437 (N_23437,N_22047,N_22783);
nand U23438 (N_23438,N_22139,N_22443);
nand U23439 (N_23439,N_22358,N_22602);
and U23440 (N_23440,N_22807,N_22906);
xnor U23441 (N_23441,N_22838,N_22371);
or U23442 (N_23442,N_22462,N_22280);
or U23443 (N_23443,N_22835,N_22929);
xnor U23444 (N_23444,N_22881,N_22704);
and U23445 (N_23445,N_22275,N_22540);
xnor U23446 (N_23446,N_22662,N_22546);
and U23447 (N_23447,N_22875,N_22799);
nor U23448 (N_23448,N_22674,N_22342);
and U23449 (N_23449,N_22861,N_22687);
xnor U23450 (N_23450,N_22933,N_22710);
nor U23451 (N_23451,N_22200,N_22099);
or U23452 (N_23452,N_22699,N_22237);
or U23453 (N_23453,N_22030,N_22423);
nor U23454 (N_23454,N_22638,N_22473);
and U23455 (N_23455,N_22128,N_22953);
nor U23456 (N_23456,N_22627,N_22601);
nand U23457 (N_23457,N_22058,N_22438);
xnor U23458 (N_23458,N_22849,N_22609);
or U23459 (N_23459,N_22895,N_22550);
and U23460 (N_23460,N_22832,N_22722);
or U23461 (N_23461,N_22381,N_22543);
xnor U23462 (N_23462,N_22013,N_22997);
nand U23463 (N_23463,N_22569,N_22317);
and U23464 (N_23464,N_22028,N_22565);
xor U23465 (N_23465,N_22903,N_22911);
and U23466 (N_23466,N_22243,N_22425);
and U23467 (N_23467,N_22260,N_22091);
nand U23468 (N_23468,N_22871,N_22466);
xnor U23469 (N_23469,N_22227,N_22817);
nand U23470 (N_23470,N_22623,N_22303);
nand U23471 (N_23471,N_22761,N_22406);
nand U23472 (N_23472,N_22117,N_22620);
or U23473 (N_23473,N_22960,N_22155);
xnor U23474 (N_23474,N_22052,N_22974);
and U23475 (N_23475,N_22225,N_22467);
nand U23476 (N_23476,N_22657,N_22907);
xnor U23477 (N_23477,N_22676,N_22442);
and U23478 (N_23478,N_22981,N_22741);
nand U23479 (N_23479,N_22604,N_22646);
nand U23480 (N_23480,N_22001,N_22693);
or U23481 (N_23481,N_22925,N_22924);
xnor U23482 (N_23482,N_22149,N_22564);
xor U23483 (N_23483,N_22599,N_22804);
nor U23484 (N_23484,N_22872,N_22608);
nand U23485 (N_23485,N_22021,N_22484);
nor U23486 (N_23486,N_22634,N_22116);
or U23487 (N_23487,N_22348,N_22967);
and U23488 (N_23488,N_22095,N_22405);
xor U23489 (N_23489,N_22880,N_22426);
nor U23490 (N_23490,N_22119,N_22578);
or U23491 (N_23491,N_22940,N_22424);
and U23492 (N_23492,N_22160,N_22842);
nor U23493 (N_23493,N_22988,N_22887);
xnor U23494 (N_23494,N_22291,N_22219);
nand U23495 (N_23495,N_22766,N_22248);
nor U23496 (N_23496,N_22018,N_22765);
xor U23497 (N_23497,N_22278,N_22830);
nand U23498 (N_23498,N_22919,N_22723);
nand U23499 (N_23499,N_22184,N_22344);
xnor U23500 (N_23500,N_22812,N_22022);
and U23501 (N_23501,N_22800,N_22191);
nor U23502 (N_23502,N_22280,N_22326);
xnor U23503 (N_23503,N_22466,N_22490);
nand U23504 (N_23504,N_22779,N_22947);
nand U23505 (N_23505,N_22341,N_22866);
nor U23506 (N_23506,N_22080,N_22845);
or U23507 (N_23507,N_22721,N_22558);
and U23508 (N_23508,N_22820,N_22783);
xor U23509 (N_23509,N_22042,N_22530);
nand U23510 (N_23510,N_22943,N_22237);
nor U23511 (N_23511,N_22649,N_22706);
nor U23512 (N_23512,N_22875,N_22098);
and U23513 (N_23513,N_22486,N_22139);
or U23514 (N_23514,N_22339,N_22962);
or U23515 (N_23515,N_22692,N_22016);
or U23516 (N_23516,N_22891,N_22334);
nor U23517 (N_23517,N_22063,N_22858);
xor U23518 (N_23518,N_22376,N_22773);
and U23519 (N_23519,N_22843,N_22789);
nor U23520 (N_23520,N_22174,N_22348);
nor U23521 (N_23521,N_22617,N_22117);
nand U23522 (N_23522,N_22364,N_22948);
nor U23523 (N_23523,N_22618,N_22820);
nor U23524 (N_23524,N_22010,N_22742);
and U23525 (N_23525,N_22890,N_22286);
xnor U23526 (N_23526,N_22163,N_22105);
xor U23527 (N_23527,N_22626,N_22493);
nor U23528 (N_23528,N_22446,N_22634);
nor U23529 (N_23529,N_22995,N_22511);
nand U23530 (N_23530,N_22490,N_22841);
or U23531 (N_23531,N_22418,N_22279);
or U23532 (N_23532,N_22448,N_22818);
and U23533 (N_23533,N_22747,N_22803);
nand U23534 (N_23534,N_22435,N_22573);
nor U23535 (N_23535,N_22046,N_22331);
or U23536 (N_23536,N_22831,N_22853);
nand U23537 (N_23537,N_22807,N_22674);
xnor U23538 (N_23538,N_22973,N_22044);
nor U23539 (N_23539,N_22720,N_22592);
nor U23540 (N_23540,N_22601,N_22744);
nor U23541 (N_23541,N_22996,N_22514);
nor U23542 (N_23542,N_22717,N_22488);
and U23543 (N_23543,N_22698,N_22810);
nand U23544 (N_23544,N_22538,N_22754);
nor U23545 (N_23545,N_22940,N_22194);
or U23546 (N_23546,N_22702,N_22263);
nor U23547 (N_23547,N_22716,N_22116);
nor U23548 (N_23548,N_22495,N_22136);
xnor U23549 (N_23549,N_22989,N_22185);
nor U23550 (N_23550,N_22772,N_22609);
or U23551 (N_23551,N_22611,N_22252);
xor U23552 (N_23552,N_22643,N_22159);
or U23553 (N_23553,N_22698,N_22537);
or U23554 (N_23554,N_22605,N_22046);
nor U23555 (N_23555,N_22947,N_22863);
nor U23556 (N_23556,N_22779,N_22249);
nor U23557 (N_23557,N_22537,N_22876);
xnor U23558 (N_23558,N_22277,N_22203);
nand U23559 (N_23559,N_22273,N_22747);
or U23560 (N_23560,N_22305,N_22937);
nand U23561 (N_23561,N_22341,N_22509);
and U23562 (N_23562,N_22245,N_22352);
and U23563 (N_23563,N_22904,N_22969);
nor U23564 (N_23564,N_22203,N_22190);
or U23565 (N_23565,N_22782,N_22436);
nand U23566 (N_23566,N_22741,N_22214);
nor U23567 (N_23567,N_22610,N_22564);
xor U23568 (N_23568,N_22673,N_22881);
xor U23569 (N_23569,N_22453,N_22466);
and U23570 (N_23570,N_22323,N_22065);
xnor U23571 (N_23571,N_22078,N_22213);
or U23572 (N_23572,N_22129,N_22933);
and U23573 (N_23573,N_22598,N_22979);
and U23574 (N_23574,N_22236,N_22941);
and U23575 (N_23575,N_22671,N_22079);
nor U23576 (N_23576,N_22727,N_22584);
nor U23577 (N_23577,N_22976,N_22177);
or U23578 (N_23578,N_22968,N_22032);
nor U23579 (N_23579,N_22070,N_22616);
and U23580 (N_23580,N_22162,N_22000);
or U23581 (N_23581,N_22563,N_22688);
nor U23582 (N_23582,N_22741,N_22885);
and U23583 (N_23583,N_22389,N_22074);
or U23584 (N_23584,N_22137,N_22048);
nand U23585 (N_23585,N_22705,N_22473);
nand U23586 (N_23586,N_22612,N_22105);
nand U23587 (N_23587,N_22811,N_22836);
nor U23588 (N_23588,N_22559,N_22968);
and U23589 (N_23589,N_22393,N_22688);
nand U23590 (N_23590,N_22994,N_22009);
or U23591 (N_23591,N_22816,N_22239);
xnor U23592 (N_23592,N_22676,N_22718);
nor U23593 (N_23593,N_22552,N_22523);
and U23594 (N_23594,N_22932,N_22376);
nor U23595 (N_23595,N_22077,N_22289);
xnor U23596 (N_23596,N_22303,N_22361);
nor U23597 (N_23597,N_22453,N_22370);
nand U23598 (N_23598,N_22129,N_22293);
nand U23599 (N_23599,N_22008,N_22668);
and U23600 (N_23600,N_22847,N_22969);
and U23601 (N_23601,N_22572,N_22330);
nand U23602 (N_23602,N_22498,N_22166);
or U23603 (N_23603,N_22811,N_22540);
nor U23604 (N_23604,N_22489,N_22683);
or U23605 (N_23605,N_22664,N_22902);
nor U23606 (N_23606,N_22105,N_22241);
and U23607 (N_23607,N_22417,N_22523);
and U23608 (N_23608,N_22584,N_22291);
nor U23609 (N_23609,N_22488,N_22510);
xnor U23610 (N_23610,N_22868,N_22124);
xor U23611 (N_23611,N_22472,N_22468);
nand U23612 (N_23612,N_22828,N_22585);
nor U23613 (N_23613,N_22021,N_22397);
and U23614 (N_23614,N_22814,N_22981);
nor U23615 (N_23615,N_22514,N_22785);
and U23616 (N_23616,N_22924,N_22939);
or U23617 (N_23617,N_22984,N_22174);
or U23618 (N_23618,N_22076,N_22156);
nand U23619 (N_23619,N_22248,N_22200);
nor U23620 (N_23620,N_22615,N_22892);
and U23621 (N_23621,N_22369,N_22027);
nand U23622 (N_23622,N_22061,N_22236);
nand U23623 (N_23623,N_22353,N_22881);
or U23624 (N_23624,N_22119,N_22909);
and U23625 (N_23625,N_22226,N_22985);
or U23626 (N_23626,N_22439,N_22584);
nand U23627 (N_23627,N_22576,N_22614);
and U23628 (N_23628,N_22133,N_22695);
nor U23629 (N_23629,N_22500,N_22328);
or U23630 (N_23630,N_22438,N_22123);
or U23631 (N_23631,N_22036,N_22547);
or U23632 (N_23632,N_22041,N_22386);
nand U23633 (N_23633,N_22440,N_22828);
xor U23634 (N_23634,N_22496,N_22432);
nand U23635 (N_23635,N_22216,N_22271);
and U23636 (N_23636,N_22533,N_22525);
and U23637 (N_23637,N_22807,N_22932);
xnor U23638 (N_23638,N_22274,N_22304);
xor U23639 (N_23639,N_22641,N_22532);
xnor U23640 (N_23640,N_22178,N_22479);
and U23641 (N_23641,N_22220,N_22664);
or U23642 (N_23642,N_22056,N_22121);
or U23643 (N_23643,N_22638,N_22624);
nand U23644 (N_23644,N_22169,N_22605);
and U23645 (N_23645,N_22782,N_22708);
and U23646 (N_23646,N_22894,N_22306);
or U23647 (N_23647,N_22216,N_22666);
xor U23648 (N_23648,N_22348,N_22903);
nor U23649 (N_23649,N_22987,N_22530);
nor U23650 (N_23650,N_22031,N_22812);
and U23651 (N_23651,N_22403,N_22939);
nor U23652 (N_23652,N_22972,N_22737);
and U23653 (N_23653,N_22226,N_22759);
and U23654 (N_23654,N_22806,N_22632);
xor U23655 (N_23655,N_22862,N_22254);
nand U23656 (N_23656,N_22185,N_22151);
xor U23657 (N_23657,N_22499,N_22647);
and U23658 (N_23658,N_22984,N_22118);
and U23659 (N_23659,N_22513,N_22887);
nor U23660 (N_23660,N_22597,N_22751);
xor U23661 (N_23661,N_22166,N_22377);
nor U23662 (N_23662,N_22503,N_22317);
and U23663 (N_23663,N_22314,N_22094);
nand U23664 (N_23664,N_22148,N_22810);
and U23665 (N_23665,N_22311,N_22812);
xnor U23666 (N_23666,N_22302,N_22908);
nand U23667 (N_23667,N_22880,N_22788);
and U23668 (N_23668,N_22117,N_22758);
and U23669 (N_23669,N_22585,N_22055);
or U23670 (N_23670,N_22193,N_22964);
or U23671 (N_23671,N_22920,N_22410);
and U23672 (N_23672,N_22140,N_22024);
nor U23673 (N_23673,N_22380,N_22716);
nor U23674 (N_23674,N_22618,N_22747);
xor U23675 (N_23675,N_22889,N_22258);
or U23676 (N_23676,N_22227,N_22771);
nand U23677 (N_23677,N_22913,N_22609);
xor U23678 (N_23678,N_22831,N_22624);
nand U23679 (N_23679,N_22340,N_22533);
nand U23680 (N_23680,N_22084,N_22759);
nand U23681 (N_23681,N_22985,N_22499);
or U23682 (N_23682,N_22542,N_22901);
xor U23683 (N_23683,N_22718,N_22202);
and U23684 (N_23684,N_22936,N_22399);
and U23685 (N_23685,N_22257,N_22036);
nor U23686 (N_23686,N_22200,N_22464);
nor U23687 (N_23687,N_22871,N_22823);
or U23688 (N_23688,N_22246,N_22053);
and U23689 (N_23689,N_22420,N_22556);
and U23690 (N_23690,N_22385,N_22103);
or U23691 (N_23691,N_22430,N_22153);
and U23692 (N_23692,N_22868,N_22447);
and U23693 (N_23693,N_22018,N_22515);
or U23694 (N_23694,N_22734,N_22231);
or U23695 (N_23695,N_22110,N_22754);
and U23696 (N_23696,N_22394,N_22697);
and U23697 (N_23697,N_22359,N_22117);
and U23698 (N_23698,N_22251,N_22788);
or U23699 (N_23699,N_22078,N_22535);
and U23700 (N_23700,N_22043,N_22758);
and U23701 (N_23701,N_22789,N_22137);
xnor U23702 (N_23702,N_22240,N_22928);
xnor U23703 (N_23703,N_22408,N_22995);
nor U23704 (N_23704,N_22663,N_22499);
or U23705 (N_23705,N_22851,N_22017);
xnor U23706 (N_23706,N_22699,N_22080);
nand U23707 (N_23707,N_22030,N_22082);
xor U23708 (N_23708,N_22835,N_22149);
nand U23709 (N_23709,N_22358,N_22799);
and U23710 (N_23710,N_22882,N_22755);
nand U23711 (N_23711,N_22842,N_22068);
nor U23712 (N_23712,N_22942,N_22428);
xor U23713 (N_23713,N_22066,N_22802);
nand U23714 (N_23714,N_22172,N_22207);
nand U23715 (N_23715,N_22694,N_22151);
and U23716 (N_23716,N_22211,N_22253);
xor U23717 (N_23717,N_22259,N_22743);
xnor U23718 (N_23718,N_22843,N_22579);
nand U23719 (N_23719,N_22424,N_22628);
or U23720 (N_23720,N_22818,N_22754);
nor U23721 (N_23721,N_22117,N_22261);
xnor U23722 (N_23722,N_22629,N_22453);
or U23723 (N_23723,N_22197,N_22110);
xor U23724 (N_23724,N_22355,N_22811);
nand U23725 (N_23725,N_22997,N_22157);
nand U23726 (N_23726,N_22904,N_22196);
or U23727 (N_23727,N_22341,N_22398);
and U23728 (N_23728,N_22934,N_22410);
or U23729 (N_23729,N_22427,N_22162);
nand U23730 (N_23730,N_22315,N_22638);
xor U23731 (N_23731,N_22616,N_22555);
nand U23732 (N_23732,N_22219,N_22167);
nand U23733 (N_23733,N_22015,N_22296);
and U23734 (N_23734,N_22435,N_22571);
nor U23735 (N_23735,N_22742,N_22260);
nor U23736 (N_23736,N_22517,N_22352);
nor U23737 (N_23737,N_22286,N_22312);
xor U23738 (N_23738,N_22753,N_22802);
nand U23739 (N_23739,N_22787,N_22956);
nand U23740 (N_23740,N_22177,N_22339);
and U23741 (N_23741,N_22725,N_22637);
and U23742 (N_23742,N_22428,N_22614);
nor U23743 (N_23743,N_22068,N_22843);
nor U23744 (N_23744,N_22567,N_22369);
or U23745 (N_23745,N_22512,N_22266);
nor U23746 (N_23746,N_22289,N_22076);
and U23747 (N_23747,N_22459,N_22662);
and U23748 (N_23748,N_22532,N_22105);
nor U23749 (N_23749,N_22546,N_22379);
and U23750 (N_23750,N_22508,N_22889);
and U23751 (N_23751,N_22871,N_22172);
xor U23752 (N_23752,N_22709,N_22801);
xnor U23753 (N_23753,N_22089,N_22340);
or U23754 (N_23754,N_22019,N_22274);
or U23755 (N_23755,N_22497,N_22588);
nor U23756 (N_23756,N_22877,N_22532);
nor U23757 (N_23757,N_22844,N_22951);
xnor U23758 (N_23758,N_22743,N_22490);
nor U23759 (N_23759,N_22955,N_22204);
xnor U23760 (N_23760,N_22906,N_22354);
and U23761 (N_23761,N_22596,N_22255);
or U23762 (N_23762,N_22428,N_22030);
nand U23763 (N_23763,N_22981,N_22616);
nand U23764 (N_23764,N_22370,N_22742);
nand U23765 (N_23765,N_22751,N_22890);
nor U23766 (N_23766,N_22562,N_22518);
nor U23767 (N_23767,N_22342,N_22847);
and U23768 (N_23768,N_22415,N_22137);
and U23769 (N_23769,N_22853,N_22282);
or U23770 (N_23770,N_22187,N_22181);
and U23771 (N_23771,N_22136,N_22343);
xor U23772 (N_23772,N_22318,N_22518);
nor U23773 (N_23773,N_22747,N_22918);
or U23774 (N_23774,N_22497,N_22498);
nor U23775 (N_23775,N_22826,N_22927);
and U23776 (N_23776,N_22816,N_22724);
xor U23777 (N_23777,N_22250,N_22393);
and U23778 (N_23778,N_22813,N_22636);
nand U23779 (N_23779,N_22789,N_22828);
xnor U23780 (N_23780,N_22379,N_22221);
or U23781 (N_23781,N_22517,N_22726);
nor U23782 (N_23782,N_22919,N_22167);
nor U23783 (N_23783,N_22176,N_22174);
or U23784 (N_23784,N_22459,N_22838);
xor U23785 (N_23785,N_22496,N_22939);
nand U23786 (N_23786,N_22818,N_22968);
xnor U23787 (N_23787,N_22355,N_22541);
xnor U23788 (N_23788,N_22697,N_22367);
and U23789 (N_23789,N_22826,N_22349);
xnor U23790 (N_23790,N_22839,N_22158);
or U23791 (N_23791,N_22356,N_22609);
and U23792 (N_23792,N_22263,N_22843);
or U23793 (N_23793,N_22404,N_22755);
nand U23794 (N_23794,N_22187,N_22776);
nand U23795 (N_23795,N_22953,N_22007);
xor U23796 (N_23796,N_22100,N_22028);
xnor U23797 (N_23797,N_22264,N_22246);
nand U23798 (N_23798,N_22946,N_22167);
or U23799 (N_23799,N_22635,N_22532);
and U23800 (N_23800,N_22911,N_22671);
or U23801 (N_23801,N_22853,N_22206);
nand U23802 (N_23802,N_22380,N_22563);
nor U23803 (N_23803,N_22574,N_22024);
nand U23804 (N_23804,N_22063,N_22609);
or U23805 (N_23805,N_22026,N_22859);
nor U23806 (N_23806,N_22636,N_22728);
or U23807 (N_23807,N_22536,N_22259);
nor U23808 (N_23808,N_22788,N_22184);
nand U23809 (N_23809,N_22536,N_22353);
or U23810 (N_23810,N_22709,N_22611);
or U23811 (N_23811,N_22565,N_22310);
or U23812 (N_23812,N_22833,N_22832);
and U23813 (N_23813,N_22193,N_22119);
and U23814 (N_23814,N_22257,N_22145);
or U23815 (N_23815,N_22106,N_22970);
or U23816 (N_23816,N_22629,N_22294);
nor U23817 (N_23817,N_22957,N_22384);
xor U23818 (N_23818,N_22697,N_22818);
or U23819 (N_23819,N_22421,N_22100);
nor U23820 (N_23820,N_22920,N_22806);
nor U23821 (N_23821,N_22931,N_22353);
and U23822 (N_23822,N_22709,N_22587);
and U23823 (N_23823,N_22361,N_22796);
and U23824 (N_23824,N_22255,N_22554);
xnor U23825 (N_23825,N_22489,N_22619);
nor U23826 (N_23826,N_22441,N_22799);
or U23827 (N_23827,N_22663,N_22080);
or U23828 (N_23828,N_22849,N_22024);
or U23829 (N_23829,N_22977,N_22460);
and U23830 (N_23830,N_22550,N_22435);
nor U23831 (N_23831,N_22152,N_22941);
nor U23832 (N_23832,N_22578,N_22736);
and U23833 (N_23833,N_22840,N_22240);
nand U23834 (N_23834,N_22872,N_22485);
and U23835 (N_23835,N_22409,N_22662);
nor U23836 (N_23836,N_22795,N_22021);
and U23837 (N_23837,N_22895,N_22278);
or U23838 (N_23838,N_22072,N_22038);
or U23839 (N_23839,N_22024,N_22606);
nor U23840 (N_23840,N_22647,N_22332);
and U23841 (N_23841,N_22124,N_22175);
nor U23842 (N_23842,N_22350,N_22079);
xnor U23843 (N_23843,N_22392,N_22420);
and U23844 (N_23844,N_22219,N_22405);
nor U23845 (N_23845,N_22428,N_22366);
nand U23846 (N_23846,N_22329,N_22753);
xor U23847 (N_23847,N_22246,N_22753);
and U23848 (N_23848,N_22717,N_22780);
or U23849 (N_23849,N_22071,N_22976);
or U23850 (N_23850,N_22012,N_22751);
xnor U23851 (N_23851,N_22669,N_22864);
and U23852 (N_23852,N_22736,N_22318);
nor U23853 (N_23853,N_22655,N_22438);
nor U23854 (N_23854,N_22753,N_22798);
xnor U23855 (N_23855,N_22069,N_22452);
nor U23856 (N_23856,N_22771,N_22486);
or U23857 (N_23857,N_22732,N_22062);
or U23858 (N_23858,N_22148,N_22248);
and U23859 (N_23859,N_22049,N_22788);
and U23860 (N_23860,N_22134,N_22426);
nor U23861 (N_23861,N_22141,N_22596);
xor U23862 (N_23862,N_22382,N_22008);
xnor U23863 (N_23863,N_22055,N_22584);
nand U23864 (N_23864,N_22619,N_22971);
and U23865 (N_23865,N_22138,N_22999);
nor U23866 (N_23866,N_22066,N_22649);
xnor U23867 (N_23867,N_22537,N_22283);
or U23868 (N_23868,N_22198,N_22553);
nor U23869 (N_23869,N_22080,N_22848);
or U23870 (N_23870,N_22343,N_22108);
xnor U23871 (N_23871,N_22851,N_22567);
or U23872 (N_23872,N_22841,N_22520);
and U23873 (N_23873,N_22311,N_22713);
nor U23874 (N_23874,N_22777,N_22906);
or U23875 (N_23875,N_22569,N_22778);
nor U23876 (N_23876,N_22248,N_22240);
and U23877 (N_23877,N_22758,N_22602);
or U23878 (N_23878,N_22439,N_22262);
or U23879 (N_23879,N_22931,N_22299);
or U23880 (N_23880,N_22212,N_22783);
nand U23881 (N_23881,N_22085,N_22169);
and U23882 (N_23882,N_22491,N_22488);
nand U23883 (N_23883,N_22904,N_22973);
or U23884 (N_23884,N_22132,N_22010);
nand U23885 (N_23885,N_22650,N_22915);
nand U23886 (N_23886,N_22896,N_22389);
nor U23887 (N_23887,N_22726,N_22826);
nor U23888 (N_23888,N_22086,N_22776);
and U23889 (N_23889,N_22406,N_22494);
or U23890 (N_23890,N_22329,N_22136);
or U23891 (N_23891,N_22461,N_22206);
or U23892 (N_23892,N_22012,N_22413);
and U23893 (N_23893,N_22327,N_22522);
and U23894 (N_23894,N_22852,N_22338);
and U23895 (N_23895,N_22601,N_22135);
or U23896 (N_23896,N_22467,N_22751);
or U23897 (N_23897,N_22666,N_22784);
or U23898 (N_23898,N_22689,N_22614);
or U23899 (N_23899,N_22000,N_22070);
nor U23900 (N_23900,N_22820,N_22209);
and U23901 (N_23901,N_22185,N_22000);
nor U23902 (N_23902,N_22332,N_22212);
nor U23903 (N_23903,N_22068,N_22148);
xnor U23904 (N_23904,N_22603,N_22277);
nand U23905 (N_23905,N_22024,N_22804);
nor U23906 (N_23906,N_22138,N_22452);
xor U23907 (N_23907,N_22718,N_22832);
and U23908 (N_23908,N_22356,N_22392);
nor U23909 (N_23909,N_22396,N_22854);
nand U23910 (N_23910,N_22218,N_22067);
xor U23911 (N_23911,N_22977,N_22699);
xnor U23912 (N_23912,N_22203,N_22576);
and U23913 (N_23913,N_22957,N_22267);
nor U23914 (N_23914,N_22302,N_22518);
nor U23915 (N_23915,N_22738,N_22679);
nand U23916 (N_23916,N_22025,N_22543);
xnor U23917 (N_23917,N_22551,N_22217);
or U23918 (N_23918,N_22005,N_22223);
nand U23919 (N_23919,N_22418,N_22376);
or U23920 (N_23920,N_22312,N_22545);
nand U23921 (N_23921,N_22489,N_22381);
nand U23922 (N_23922,N_22269,N_22150);
or U23923 (N_23923,N_22506,N_22771);
or U23924 (N_23924,N_22861,N_22130);
nand U23925 (N_23925,N_22664,N_22095);
nor U23926 (N_23926,N_22727,N_22842);
or U23927 (N_23927,N_22053,N_22607);
and U23928 (N_23928,N_22171,N_22133);
and U23929 (N_23929,N_22271,N_22077);
or U23930 (N_23930,N_22037,N_22941);
and U23931 (N_23931,N_22668,N_22454);
xnor U23932 (N_23932,N_22097,N_22191);
xor U23933 (N_23933,N_22628,N_22653);
and U23934 (N_23934,N_22097,N_22393);
and U23935 (N_23935,N_22829,N_22958);
and U23936 (N_23936,N_22495,N_22189);
xor U23937 (N_23937,N_22520,N_22890);
and U23938 (N_23938,N_22761,N_22165);
xnor U23939 (N_23939,N_22869,N_22096);
xnor U23940 (N_23940,N_22869,N_22363);
nor U23941 (N_23941,N_22353,N_22908);
and U23942 (N_23942,N_22902,N_22165);
nor U23943 (N_23943,N_22344,N_22580);
nor U23944 (N_23944,N_22889,N_22957);
xor U23945 (N_23945,N_22749,N_22457);
and U23946 (N_23946,N_22497,N_22787);
xnor U23947 (N_23947,N_22643,N_22870);
and U23948 (N_23948,N_22560,N_22651);
nor U23949 (N_23949,N_22442,N_22545);
and U23950 (N_23950,N_22524,N_22566);
nand U23951 (N_23951,N_22410,N_22627);
or U23952 (N_23952,N_22423,N_22398);
nand U23953 (N_23953,N_22694,N_22126);
nand U23954 (N_23954,N_22291,N_22211);
nor U23955 (N_23955,N_22522,N_22945);
xor U23956 (N_23956,N_22328,N_22982);
or U23957 (N_23957,N_22723,N_22016);
xnor U23958 (N_23958,N_22730,N_22957);
nand U23959 (N_23959,N_22302,N_22093);
nand U23960 (N_23960,N_22509,N_22694);
nor U23961 (N_23961,N_22472,N_22397);
nand U23962 (N_23962,N_22728,N_22398);
xnor U23963 (N_23963,N_22498,N_22769);
nand U23964 (N_23964,N_22438,N_22513);
nand U23965 (N_23965,N_22505,N_22743);
or U23966 (N_23966,N_22204,N_22475);
nand U23967 (N_23967,N_22976,N_22532);
nand U23968 (N_23968,N_22753,N_22128);
nand U23969 (N_23969,N_22056,N_22188);
or U23970 (N_23970,N_22164,N_22383);
and U23971 (N_23971,N_22642,N_22362);
nand U23972 (N_23972,N_22721,N_22891);
nand U23973 (N_23973,N_22922,N_22752);
or U23974 (N_23974,N_22506,N_22682);
xor U23975 (N_23975,N_22099,N_22424);
nand U23976 (N_23976,N_22697,N_22744);
and U23977 (N_23977,N_22204,N_22515);
or U23978 (N_23978,N_22605,N_22083);
nor U23979 (N_23979,N_22822,N_22855);
and U23980 (N_23980,N_22228,N_22746);
xnor U23981 (N_23981,N_22205,N_22441);
and U23982 (N_23982,N_22799,N_22250);
or U23983 (N_23983,N_22554,N_22791);
or U23984 (N_23984,N_22604,N_22417);
or U23985 (N_23985,N_22693,N_22709);
nand U23986 (N_23986,N_22574,N_22168);
and U23987 (N_23987,N_22429,N_22254);
or U23988 (N_23988,N_22618,N_22293);
nand U23989 (N_23989,N_22419,N_22399);
nor U23990 (N_23990,N_22316,N_22796);
nor U23991 (N_23991,N_22396,N_22973);
nor U23992 (N_23992,N_22701,N_22605);
nor U23993 (N_23993,N_22299,N_22970);
nor U23994 (N_23994,N_22091,N_22988);
or U23995 (N_23995,N_22751,N_22830);
or U23996 (N_23996,N_22615,N_22106);
xnor U23997 (N_23997,N_22741,N_22890);
nor U23998 (N_23998,N_22176,N_22657);
and U23999 (N_23999,N_22614,N_22734);
xnor U24000 (N_24000,N_23316,N_23380);
nor U24001 (N_24001,N_23008,N_23466);
nand U24002 (N_24002,N_23113,N_23818);
and U24003 (N_24003,N_23475,N_23406);
nor U24004 (N_24004,N_23399,N_23169);
nor U24005 (N_24005,N_23245,N_23176);
or U24006 (N_24006,N_23044,N_23618);
xnor U24007 (N_24007,N_23200,N_23847);
xor U24008 (N_24008,N_23971,N_23908);
nor U24009 (N_24009,N_23518,N_23923);
nor U24010 (N_24010,N_23440,N_23034);
nand U24011 (N_24011,N_23048,N_23275);
xnor U24012 (N_24012,N_23080,N_23456);
and U24013 (N_24013,N_23804,N_23589);
nor U24014 (N_24014,N_23712,N_23092);
and U24015 (N_24015,N_23689,N_23401);
or U24016 (N_24016,N_23747,N_23797);
nor U24017 (N_24017,N_23723,N_23094);
nand U24018 (N_24018,N_23108,N_23991);
nor U24019 (N_24019,N_23248,N_23887);
nor U24020 (N_24020,N_23769,N_23358);
xnor U24021 (N_24021,N_23146,N_23751);
nand U24022 (N_24022,N_23820,N_23356);
xnor U24023 (N_24023,N_23251,N_23269);
nand U24024 (N_24024,N_23821,N_23650);
nor U24025 (N_24025,N_23542,N_23907);
or U24026 (N_24026,N_23594,N_23533);
nor U24027 (N_24027,N_23919,N_23615);
and U24028 (N_24028,N_23564,N_23732);
nor U24029 (N_24029,N_23695,N_23610);
xor U24030 (N_24030,N_23521,N_23304);
nand U24031 (N_24031,N_23525,N_23089);
nand U24032 (N_24032,N_23881,N_23026);
and U24033 (N_24033,N_23928,N_23306);
or U24034 (N_24034,N_23760,N_23943);
nand U24035 (N_24035,N_23672,N_23052);
and U24036 (N_24036,N_23683,N_23260);
nand U24037 (N_24037,N_23295,N_23903);
xnor U24038 (N_24038,N_23174,N_23638);
xor U24039 (N_24039,N_23381,N_23411);
nor U24040 (N_24040,N_23229,N_23460);
and U24041 (N_24041,N_23485,N_23942);
xnor U24042 (N_24042,N_23920,N_23081);
nand U24043 (N_24043,N_23163,N_23735);
and U24044 (N_24044,N_23710,N_23540);
nand U24045 (N_24045,N_23344,N_23425);
nor U24046 (N_24046,N_23022,N_23532);
and U24047 (N_24047,N_23974,N_23167);
nand U24048 (N_24048,N_23509,N_23230);
or U24049 (N_24049,N_23668,N_23550);
nor U24050 (N_24050,N_23020,N_23177);
and U24051 (N_24051,N_23010,N_23256);
and U24052 (N_24052,N_23310,N_23617);
nand U24053 (N_24053,N_23687,N_23038);
nor U24054 (N_24054,N_23368,N_23072);
and U24055 (N_24055,N_23927,N_23083);
nor U24056 (N_24056,N_23675,N_23470);
xnor U24057 (N_24057,N_23829,N_23995);
xor U24058 (N_24058,N_23205,N_23603);
nor U24059 (N_24059,N_23472,N_23294);
or U24060 (N_24060,N_23395,N_23292);
xnor U24061 (N_24061,N_23711,N_23051);
nor U24062 (N_24062,N_23186,N_23671);
xnor U24063 (N_24063,N_23071,N_23377);
nand U24064 (N_24064,N_23916,N_23910);
or U24065 (N_24065,N_23115,N_23501);
nor U24066 (N_24066,N_23773,N_23794);
xnor U24067 (N_24067,N_23311,N_23076);
or U24068 (N_24068,N_23741,N_23299);
and U24069 (N_24069,N_23001,N_23599);
and U24070 (N_24070,N_23144,N_23369);
or U24071 (N_24071,N_23544,N_23152);
nand U24072 (N_24072,N_23236,N_23447);
xnor U24073 (N_24073,N_23692,N_23165);
and U24074 (N_24074,N_23983,N_23779);
xor U24075 (N_24075,N_23998,N_23491);
or U24076 (N_24076,N_23187,N_23562);
nand U24077 (N_24077,N_23255,N_23137);
nand U24078 (N_24078,N_23517,N_23379);
nand U24079 (N_24079,N_23280,N_23097);
nand U24080 (N_24080,N_23288,N_23850);
and U24081 (N_24081,N_23351,N_23538);
xor U24082 (N_24082,N_23590,N_23558);
nor U24083 (N_24083,N_23678,N_23098);
or U24084 (N_24084,N_23309,N_23028);
nor U24085 (N_24085,N_23270,N_23947);
xor U24086 (N_24086,N_23597,N_23627);
xor U24087 (N_24087,N_23832,N_23331);
nand U24088 (N_24088,N_23053,N_23366);
nor U24089 (N_24089,N_23359,N_23272);
xnor U24090 (N_24090,N_23107,N_23463);
or U24091 (N_24091,N_23824,N_23465);
and U24092 (N_24092,N_23863,N_23082);
or U24093 (N_24093,N_23748,N_23003);
and U24094 (N_24094,N_23009,N_23816);
nand U24095 (N_24095,N_23516,N_23583);
nor U24096 (N_24096,N_23807,N_23729);
and U24097 (N_24097,N_23731,N_23030);
nand U24098 (N_24098,N_23029,N_23625);
xnor U24099 (N_24099,N_23147,N_23823);
nor U24100 (N_24100,N_23314,N_23375);
nor U24101 (N_24101,N_23159,N_23642);
nand U24102 (N_24102,N_23874,N_23450);
nand U24103 (N_24103,N_23244,N_23233);
nor U24104 (N_24104,N_23720,N_23464);
xor U24105 (N_24105,N_23041,N_23857);
xnor U24106 (N_24106,N_23855,N_23911);
xor U24107 (N_24107,N_23803,N_23252);
and U24108 (N_24108,N_23204,N_23702);
nor U24109 (N_24109,N_23981,N_23929);
and U24110 (N_24110,N_23969,N_23070);
and U24111 (N_24111,N_23812,N_23962);
nand U24112 (N_24112,N_23452,N_23116);
xor U24113 (N_24113,N_23324,N_23524);
and U24114 (N_24114,N_23700,N_23035);
nand U24115 (N_24115,N_23944,N_23705);
nand U24116 (N_24116,N_23964,N_23017);
or U24117 (N_24117,N_23922,N_23199);
or U24118 (N_24118,N_23750,N_23960);
nor U24119 (N_24119,N_23125,N_23914);
or U24120 (N_24120,N_23455,N_23905);
xnor U24121 (N_24121,N_23537,N_23242);
xor U24122 (N_24122,N_23561,N_23132);
xnor U24123 (N_24123,N_23011,N_23254);
and U24124 (N_24124,N_23577,N_23523);
or U24125 (N_24125,N_23828,N_23334);
xor U24126 (N_24126,N_23303,N_23527);
or U24127 (N_24127,N_23579,N_23228);
or U24128 (N_24128,N_23873,N_23197);
nor U24129 (N_24129,N_23099,N_23541);
and U24130 (N_24130,N_23640,N_23000);
and U24131 (N_24131,N_23154,N_23612);
and U24132 (N_24132,N_23774,N_23481);
or U24133 (N_24133,N_23293,N_23067);
xnor U24134 (N_24134,N_23392,N_23933);
xnor U24135 (N_24135,N_23586,N_23184);
nor U24136 (N_24136,N_23234,N_23364);
xnor U24137 (N_24137,N_23383,N_23047);
nand U24138 (N_24138,N_23024,N_23755);
nand U24139 (N_24139,N_23600,N_23085);
nand U24140 (N_24140,N_23330,N_23609);
and U24141 (N_24141,N_23906,N_23802);
or U24142 (N_24142,N_23385,N_23734);
nand U24143 (N_24143,N_23993,N_23637);
nor U24144 (N_24144,N_23814,N_23339);
nand U24145 (N_24145,N_23241,N_23882);
xor U24146 (N_24146,N_23461,N_23346);
xnor U24147 (N_24147,N_23651,N_23396);
nand U24148 (N_24148,N_23208,N_23939);
nor U24149 (N_24149,N_23694,N_23374);
nand U24150 (N_24150,N_23247,N_23635);
nor U24151 (N_24151,N_23831,N_23834);
nand U24152 (N_24152,N_23511,N_23063);
nand U24153 (N_24153,N_23110,N_23614);
nor U24154 (N_24154,N_23124,N_23982);
xnor U24155 (N_24155,N_23219,N_23681);
xnor U24156 (N_24156,N_23393,N_23179);
xor U24157 (N_24157,N_23646,N_23736);
and U24158 (N_24158,N_23183,N_23566);
and U24159 (N_24159,N_23046,N_23508);
nor U24160 (N_24160,N_23210,N_23231);
nor U24161 (N_24161,N_23037,N_23663);
nand U24162 (N_24162,N_23345,N_23434);
or U24163 (N_24163,N_23768,N_23168);
and U24164 (N_24164,N_23556,N_23900);
xnor U24165 (N_24165,N_23134,N_23058);
or U24166 (N_24166,N_23634,N_23135);
nor U24167 (N_24167,N_23826,N_23648);
xor U24168 (N_24168,N_23415,N_23622);
nor U24169 (N_24169,N_23567,N_23340);
nor U24170 (N_24170,N_23502,N_23601);
and U24171 (N_24171,N_23665,N_23250);
or U24172 (N_24172,N_23496,N_23512);
nand U24173 (N_24173,N_23438,N_23505);
nor U24174 (N_24174,N_23221,N_23764);
nand U24175 (N_24175,N_23825,N_23235);
nand U24176 (N_24176,N_23361,N_23321);
or U24177 (N_24177,N_23921,N_23238);
xor U24178 (N_24178,N_23817,N_23422);
or U24179 (N_24179,N_23867,N_23613);
nor U24180 (N_24180,N_23936,N_23019);
xor U24181 (N_24181,N_23387,N_23431);
or U24182 (N_24182,N_23077,N_23068);
and U24183 (N_24183,N_23569,N_23018);
nor U24184 (N_24184,N_23087,N_23467);
nor U24185 (N_24185,N_23519,N_23428);
nand U24186 (N_24186,N_23468,N_23106);
nand U24187 (N_24187,N_23102,N_23909);
and U24188 (N_24188,N_23746,N_23273);
nor U24189 (N_24189,N_23996,N_23363);
nor U24190 (N_24190,N_23598,N_23480);
nand U24191 (N_24191,N_23979,N_23931);
or U24192 (N_24192,N_23155,N_23386);
xor U24193 (N_24193,N_23770,N_23565);
nor U24194 (N_24194,N_23477,N_23941);
or U24195 (N_24195,N_23448,N_23439);
nor U24196 (N_24196,N_23629,N_23858);
or U24197 (N_24197,N_23782,N_23126);
xor U24198 (N_24198,N_23259,N_23785);
xnor U24199 (N_24199,N_23877,N_23660);
xor U24200 (N_24200,N_23957,N_23840);
or U24201 (N_24201,N_23062,N_23693);
and U24202 (N_24202,N_23582,N_23984);
xnor U24203 (N_24203,N_23086,N_23889);
nand U24204 (N_24204,N_23326,N_23657);
nand U24205 (N_24205,N_23655,N_23917);
and U24206 (N_24206,N_23454,N_23551);
and U24207 (N_24207,N_23703,N_23185);
nor U24208 (N_24208,N_23194,N_23066);
or U24209 (N_24209,N_23285,N_23193);
and U24210 (N_24210,N_23503,N_23967);
xor U24211 (N_24211,N_23362,N_23446);
and U24212 (N_24212,N_23459,N_23312);
nor U24213 (N_24213,N_23725,N_23261);
and U24214 (N_24214,N_23726,N_23716);
or U24215 (N_24215,N_23975,N_23243);
nor U24216 (N_24216,N_23557,N_23654);
xor U24217 (N_24217,N_23105,N_23658);
and U24218 (N_24218,N_23198,N_23427);
and U24219 (N_24219,N_23056,N_23253);
xnor U24220 (N_24220,N_23320,N_23898);
xnor U24221 (N_24221,N_23913,N_23435);
or U24222 (N_24222,N_23227,N_23699);
xnor U24223 (N_24223,N_23781,N_23278);
xor U24224 (N_24224,N_23333,N_23581);
or U24225 (N_24225,N_23656,N_23886);
nor U24226 (N_24226,N_23758,N_23684);
and U24227 (N_24227,N_23948,N_23645);
nand U24228 (N_24228,N_23783,N_23103);
nor U24229 (N_24229,N_23878,N_23265);
and U24230 (N_24230,N_23515,N_23189);
or U24231 (N_24231,N_23968,N_23584);
or U24232 (N_24232,N_23997,N_23739);
nand U24233 (N_24233,N_23170,N_23350);
nor U24234 (N_24234,N_23045,N_23043);
nand U24235 (N_24235,N_23871,N_23765);
nor U24236 (N_24236,N_23894,N_23372);
xnor U24237 (N_24237,N_23520,N_23707);
or U24238 (N_24238,N_23271,N_23553);
and U24239 (N_24239,N_23360,N_23282);
and U24240 (N_24240,N_23891,N_23930);
or U24241 (N_24241,N_23757,N_23950);
or U24242 (N_24242,N_23813,N_23940);
and U24243 (N_24243,N_23192,N_23506);
and U24244 (N_24244,N_23182,N_23397);
and U24245 (N_24245,N_23213,N_23141);
and U24246 (N_24246,N_23493,N_23611);
or U24247 (N_24247,N_23514,N_23389);
xor U24248 (N_24248,N_23206,N_23596);
or U24249 (N_24249,N_23109,N_23639);
nand U24250 (N_24250,N_23780,N_23258);
nor U24251 (N_24251,N_23535,N_23744);
xnor U24252 (N_24252,N_23162,N_23059);
xor U24253 (N_24253,N_23680,N_23897);
nor U24254 (N_24254,N_23420,N_23970);
nor U24255 (N_24255,N_23737,N_23845);
xnor U24256 (N_24256,N_23628,N_23846);
and U24257 (N_24257,N_23578,N_23136);
or U24258 (N_24258,N_23343,N_23093);
or U24259 (N_24259,N_23322,N_23139);
xnor U24260 (N_24260,N_23216,N_23268);
xor U24261 (N_24261,N_23133,N_23257);
nor U24262 (N_24262,N_23423,N_23078);
or U24263 (N_24263,N_23490,N_23547);
or U24264 (N_24264,N_23698,N_23895);
xnor U24265 (N_24265,N_23959,N_23743);
and U24266 (N_24266,N_23025,N_23786);
nor U24267 (N_24267,N_23837,N_23088);
and U24268 (N_24268,N_23408,N_23100);
or U24269 (N_24269,N_23302,N_23573);
and U24270 (N_24270,N_23403,N_23761);
or U24271 (N_24271,N_23354,N_23706);
or U24272 (N_24272,N_23752,N_23795);
or U24273 (N_24273,N_23417,N_23652);
and U24274 (N_24274,N_23669,N_23549);
nor U24275 (N_24275,N_23203,N_23277);
xnor U24276 (N_24276,N_23801,N_23483);
and U24277 (N_24277,N_23178,N_23872);
nor U24278 (N_24278,N_23153,N_23307);
nand U24279 (N_24279,N_23559,N_23842);
nor U24280 (N_24280,N_23064,N_23575);
nand U24281 (N_24281,N_23819,N_23457);
and U24282 (N_24282,N_23370,N_23954);
nor U24283 (N_24283,N_23091,N_23545);
nor U24284 (N_24284,N_23436,N_23649);
and U24285 (N_24285,N_23902,N_23543);
or U24286 (N_24286,N_23958,N_23745);
nand U24287 (N_24287,N_23787,N_23171);
or U24288 (N_24288,N_23384,N_23714);
nand U24289 (N_24289,N_23836,N_23632);
or U24290 (N_24290,N_23955,N_23104);
nand U24291 (N_24291,N_23050,N_23497);
nand U24292 (N_24292,N_23851,N_23337);
nand U24293 (N_24293,N_23014,N_23718);
or U24294 (N_24294,N_23572,N_23479);
nor U24295 (N_24295,N_23095,N_23191);
and U24296 (N_24296,N_23484,N_23934);
nor U24297 (N_24297,N_23976,N_23643);
nor U24298 (N_24298,N_23588,N_23027);
and U24299 (N_24299,N_23937,N_23398);
xnor U24300 (N_24300,N_23945,N_23555);
nor U24301 (N_24301,N_23342,N_23724);
and U24302 (N_24302,N_23890,N_23410);
and U24303 (N_24303,N_23195,N_23462);
nor U24304 (N_24304,N_23209,N_23616);
nor U24305 (N_24305,N_23513,N_23861);
nor U24306 (N_24306,N_23901,N_23042);
or U24307 (N_24307,N_23719,N_23630);
and U24308 (N_24308,N_23951,N_23978);
nor U24309 (N_24309,N_23373,N_23591);
nor U24310 (N_24310,N_23328,N_23054);
or U24311 (N_24311,N_23560,N_23722);
xnor U24312 (N_24312,N_23138,N_23388);
nand U24313 (N_24313,N_23987,N_23666);
and U24314 (N_24314,N_23130,N_23778);
nand U24315 (N_24315,N_23114,N_23140);
or U24316 (N_24316,N_23691,N_23033);
nor U24317 (N_24317,N_23430,N_23500);
or U24318 (N_24318,N_23528,N_23529);
and U24319 (N_24319,N_23469,N_23868);
or U24320 (N_24320,N_23738,N_23604);
and U24321 (N_24321,N_23507,N_23756);
and U24322 (N_24322,N_23433,N_23232);
and U24323 (N_24323,N_23414,N_23266);
and U24324 (N_24324,N_23355,N_23784);
xnor U24325 (N_24325,N_23742,N_23246);
xor U24326 (N_24326,N_23548,N_23166);
xnor U24327 (N_24327,N_23471,N_23992);
or U24328 (N_24328,N_23498,N_23437);
and U24329 (N_24329,N_23158,N_23021);
xnor U24330 (N_24330,N_23161,N_23443);
and U24331 (N_24331,N_23214,N_23036);
xor U24332 (N_24332,N_23237,N_23129);
or U24333 (N_24333,N_23202,N_23365);
and U24334 (N_24334,N_23055,N_23290);
or U24335 (N_24335,N_23404,N_23715);
xnor U24336 (N_24336,N_23990,N_23988);
nand U24337 (N_24337,N_23218,N_23090);
nor U24338 (N_24338,N_23016,N_23965);
or U24339 (N_24339,N_23156,N_23674);
and U24340 (N_24340,N_23686,N_23754);
and U24341 (N_24341,N_23626,N_23806);
or U24342 (N_24342,N_23220,N_23069);
and U24343 (N_24343,N_23977,N_23039);
and U24344 (N_24344,N_23763,N_23262);
nor U24345 (N_24345,N_23402,N_23127);
and U24346 (N_24346,N_23932,N_23859);
or U24347 (N_24347,N_23151,N_23790);
or U24348 (N_24348,N_23989,N_23673);
or U24349 (N_24349,N_23224,N_23117);
or U24350 (N_24350,N_23486,N_23608);
and U24351 (N_24351,N_23510,N_23264);
nand U24352 (N_24352,N_23972,N_23717);
xor U24353 (N_24353,N_23865,N_23031);
nor U24354 (N_24354,N_23487,N_23904);
nor U24355 (N_24355,N_23662,N_23349);
and U24356 (N_24356,N_23444,N_23776);
and U24357 (N_24357,N_23201,N_23180);
and U24358 (N_24358,N_23376,N_23587);
or U24359 (N_24359,N_23313,N_23606);
nand U24360 (N_24360,N_23263,N_23876);
and U24361 (N_24361,N_23833,N_23841);
nor U24362 (N_24362,N_23864,N_23329);
nand U24363 (N_24363,N_23593,N_23323);
nand U24364 (N_24364,N_23869,N_23429);
nand U24365 (N_24365,N_23727,N_23796);
or U24366 (N_24366,N_23585,N_23623);
nand U24367 (N_24367,N_23994,N_23286);
nor U24368 (N_24368,N_23488,N_23912);
xnor U24369 (N_24369,N_23570,N_23005);
and U24370 (N_24370,N_23844,N_23338);
nand U24371 (N_24371,N_23451,N_23418);
nand U24372 (N_24372,N_23679,N_23647);
nand U24373 (N_24373,N_23644,N_23061);
nor U24374 (N_24374,N_23862,N_23074);
or U24375 (N_24375,N_23495,N_23341);
or U24376 (N_24376,N_23300,N_23664);
xor U24377 (N_24377,N_23296,N_23677);
nand U24378 (N_24378,N_23308,N_23453);
xnor U24379 (N_24379,N_23442,N_23670);
xnor U24380 (N_24380,N_23407,N_23838);
nor U24381 (N_24381,N_23297,N_23196);
xor U24382 (N_24382,N_23499,N_23676);
nor U24383 (N_24383,N_23822,N_23875);
nor U24384 (N_24384,N_23605,N_23318);
and U24385 (N_24385,N_23118,N_23696);
nand U24386 (N_24386,N_23766,N_23641);
nor U24387 (N_24387,N_23708,N_23883);
or U24388 (N_24388,N_23534,N_23409);
or U24389 (N_24389,N_23815,N_23225);
nand U24390 (N_24390,N_23592,N_23697);
and U24391 (N_24391,N_23949,N_23073);
nor U24392 (N_24392,N_23504,N_23574);
or U24393 (N_24393,N_23412,N_23283);
nor U24394 (N_24394,N_23685,N_23854);
xnor U24395 (N_24395,N_23421,N_23327);
and U24396 (N_24396,N_23682,N_23771);
nor U24397 (N_24397,N_23172,N_23382);
xor U24398 (N_24398,N_23175,N_23419);
nor U24399 (N_24399,N_23536,N_23805);
nor U24400 (N_24400,N_23624,N_23935);
nor U24401 (N_24401,N_23284,N_23653);
or U24402 (N_24402,N_23733,N_23449);
xor U24403 (N_24403,N_23704,N_23777);
xor U24404 (N_24404,N_23728,N_23986);
nand U24405 (N_24405,N_23870,N_23860);
and U24406 (N_24406,N_23966,N_23999);
xor U24407 (N_24407,N_23849,N_23848);
nand U24408 (N_24408,N_23226,N_23075);
nand U24409 (N_24409,N_23367,N_23791);
nor U24410 (N_24410,N_23289,N_23123);
nand U24411 (N_24411,N_23985,N_23004);
or U24412 (N_24412,N_23918,N_23276);
and U24413 (N_24413,N_23753,N_23852);
nor U24414 (N_24414,N_23079,N_23032);
xor U24415 (N_24415,N_23274,N_23347);
nor U24416 (N_24416,N_23239,N_23150);
and U24417 (N_24417,N_23980,N_23607);
nand U24418 (N_24418,N_23602,N_23145);
or U24419 (N_24419,N_23298,N_23223);
or U24420 (N_24420,N_23925,N_23762);
nor U24421 (N_24421,N_23554,N_23291);
nand U24422 (N_24422,N_23121,N_23926);
or U24423 (N_24423,N_23489,N_23482);
xnor U24424 (N_24424,N_23946,N_23580);
xnor U24425 (N_24425,N_23040,N_23207);
or U24426 (N_24426,N_23149,N_23798);
xor U24427 (N_24427,N_23810,N_23631);
xor U24428 (N_24428,N_23952,N_23181);
and U24429 (N_24429,N_23305,N_23101);
nor U24430 (N_24430,N_23267,N_23661);
nand U24431 (N_24431,N_23458,N_23432);
nand U24432 (N_24432,N_23494,N_23119);
or U24433 (N_24433,N_23963,N_23122);
and U24434 (N_24434,N_23839,N_23476);
and U24435 (N_24435,N_23530,N_23473);
and U24436 (N_24436,N_23315,N_23281);
nor U24437 (N_24437,N_23002,N_23120);
nand U24438 (N_24438,N_23893,N_23357);
xor U24439 (N_24439,N_23348,N_23390);
nand U24440 (N_24440,N_23853,N_23287);
or U24441 (N_24441,N_23827,N_23249);
nand U24442 (N_24442,N_23740,N_23730);
and U24443 (N_24443,N_23636,N_23809);
nor U24444 (N_24444,N_23709,N_23478);
xor U24445 (N_24445,N_23128,N_23015);
xor U24446 (N_24446,N_23563,N_23400);
nor U24447 (N_24447,N_23424,N_23788);
or U24448 (N_24448,N_23353,N_23416);
or U24449 (N_24449,N_23336,N_23866);
or U24450 (N_24450,N_23749,N_23633);
nand U24451 (N_24451,N_23441,N_23688);
nor U24452 (N_24452,N_23884,N_23317);
xor U24453 (N_24453,N_23799,N_23539);
and U24454 (N_24454,N_23474,N_23595);
nor U24455 (N_24455,N_23173,N_23405);
nor U24456 (N_24456,N_23793,N_23157);
or U24457 (N_24457,N_23160,N_23049);
and U24458 (N_24458,N_23084,N_23531);
nand U24459 (N_24459,N_23885,N_23843);
or U24460 (N_24460,N_23222,N_23759);
nor U24461 (N_24461,N_23690,N_23013);
nor U24462 (N_24462,N_23888,N_23143);
nor U24463 (N_24463,N_23619,N_23023);
xnor U24464 (N_24464,N_23332,N_23352);
or U24465 (N_24465,N_23571,N_23856);
xor U24466 (N_24466,N_23112,N_23811);
xnor U24467 (N_24467,N_23060,N_23335);
nand U24468 (N_24468,N_23096,N_23279);
or U24469 (N_24469,N_23667,N_23142);
nand U24470 (N_24470,N_23879,N_23552);
nor U24471 (N_24471,N_23492,N_23426);
nor U24472 (N_24472,N_23659,N_23808);
nor U24473 (N_24473,N_23924,N_23789);
xor U24474 (N_24474,N_23215,N_23938);
and U24475 (N_24475,N_23713,N_23892);
nor U24476 (N_24476,N_23775,N_23148);
nand U24477 (N_24477,N_23131,N_23445);
nand U24478 (N_24478,N_23012,N_23772);
nor U24479 (N_24479,N_23188,N_23546);
nand U24480 (N_24480,N_23568,N_23961);
xnor U24481 (N_24481,N_23371,N_23896);
and U24482 (N_24482,N_23413,N_23830);
nand U24483 (N_24483,N_23211,N_23006);
nand U24484 (N_24484,N_23956,N_23800);
nor U24485 (N_24485,N_23899,N_23973);
nand U24486 (N_24486,N_23792,N_23319);
and U24487 (N_24487,N_23394,N_23391);
and U24488 (N_24488,N_23057,N_23721);
or U24489 (N_24489,N_23767,N_23240);
and U24490 (N_24490,N_23378,N_23111);
nor U24491 (N_24491,N_23701,N_23217);
nor U24492 (N_24492,N_23301,N_23953);
and U24493 (N_24493,N_23620,N_23621);
xnor U24494 (N_24494,N_23880,N_23065);
xor U24495 (N_24495,N_23212,N_23164);
or U24496 (N_24496,N_23915,N_23576);
or U24497 (N_24497,N_23190,N_23007);
nand U24498 (N_24498,N_23325,N_23522);
nor U24499 (N_24499,N_23835,N_23526);
xor U24500 (N_24500,N_23798,N_23646);
nor U24501 (N_24501,N_23053,N_23090);
nor U24502 (N_24502,N_23482,N_23830);
xnor U24503 (N_24503,N_23901,N_23503);
nand U24504 (N_24504,N_23317,N_23650);
or U24505 (N_24505,N_23354,N_23268);
nand U24506 (N_24506,N_23437,N_23740);
and U24507 (N_24507,N_23706,N_23098);
and U24508 (N_24508,N_23677,N_23619);
xnor U24509 (N_24509,N_23543,N_23782);
or U24510 (N_24510,N_23727,N_23283);
or U24511 (N_24511,N_23278,N_23259);
nor U24512 (N_24512,N_23756,N_23688);
and U24513 (N_24513,N_23301,N_23622);
nor U24514 (N_24514,N_23736,N_23910);
nor U24515 (N_24515,N_23072,N_23201);
and U24516 (N_24516,N_23152,N_23524);
and U24517 (N_24517,N_23287,N_23366);
xnor U24518 (N_24518,N_23797,N_23352);
or U24519 (N_24519,N_23669,N_23429);
xor U24520 (N_24520,N_23306,N_23229);
or U24521 (N_24521,N_23332,N_23282);
nand U24522 (N_24522,N_23372,N_23928);
nand U24523 (N_24523,N_23079,N_23571);
nand U24524 (N_24524,N_23531,N_23568);
nor U24525 (N_24525,N_23412,N_23759);
and U24526 (N_24526,N_23158,N_23943);
xnor U24527 (N_24527,N_23603,N_23003);
and U24528 (N_24528,N_23139,N_23550);
and U24529 (N_24529,N_23452,N_23019);
xor U24530 (N_24530,N_23863,N_23430);
and U24531 (N_24531,N_23557,N_23930);
nand U24532 (N_24532,N_23161,N_23699);
or U24533 (N_24533,N_23502,N_23028);
xor U24534 (N_24534,N_23745,N_23016);
nand U24535 (N_24535,N_23931,N_23492);
xor U24536 (N_24536,N_23791,N_23432);
or U24537 (N_24537,N_23266,N_23790);
or U24538 (N_24538,N_23282,N_23137);
and U24539 (N_24539,N_23383,N_23779);
xor U24540 (N_24540,N_23965,N_23791);
nor U24541 (N_24541,N_23377,N_23883);
nand U24542 (N_24542,N_23771,N_23698);
nor U24543 (N_24543,N_23822,N_23559);
or U24544 (N_24544,N_23236,N_23396);
nor U24545 (N_24545,N_23839,N_23609);
nor U24546 (N_24546,N_23445,N_23225);
xnor U24547 (N_24547,N_23546,N_23153);
xnor U24548 (N_24548,N_23387,N_23839);
xnor U24549 (N_24549,N_23192,N_23171);
xnor U24550 (N_24550,N_23750,N_23402);
nand U24551 (N_24551,N_23367,N_23635);
nor U24552 (N_24552,N_23512,N_23180);
and U24553 (N_24553,N_23123,N_23836);
nand U24554 (N_24554,N_23417,N_23918);
nand U24555 (N_24555,N_23561,N_23327);
and U24556 (N_24556,N_23190,N_23338);
nand U24557 (N_24557,N_23494,N_23332);
nor U24558 (N_24558,N_23378,N_23907);
xnor U24559 (N_24559,N_23262,N_23259);
xor U24560 (N_24560,N_23982,N_23866);
nand U24561 (N_24561,N_23016,N_23469);
and U24562 (N_24562,N_23686,N_23065);
xnor U24563 (N_24563,N_23591,N_23464);
nor U24564 (N_24564,N_23199,N_23935);
nand U24565 (N_24565,N_23196,N_23746);
nor U24566 (N_24566,N_23271,N_23324);
and U24567 (N_24567,N_23374,N_23279);
nor U24568 (N_24568,N_23197,N_23794);
xnor U24569 (N_24569,N_23449,N_23967);
xnor U24570 (N_24570,N_23396,N_23683);
nand U24571 (N_24571,N_23485,N_23914);
and U24572 (N_24572,N_23861,N_23491);
or U24573 (N_24573,N_23354,N_23257);
xor U24574 (N_24574,N_23450,N_23497);
nand U24575 (N_24575,N_23165,N_23646);
nor U24576 (N_24576,N_23142,N_23332);
or U24577 (N_24577,N_23909,N_23977);
and U24578 (N_24578,N_23473,N_23391);
nor U24579 (N_24579,N_23921,N_23546);
and U24580 (N_24580,N_23428,N_23436);
xor U24581 (N_24581,N_23983,N_23764);
and U24582 (N_24582,N_23947,N_23104);
nand U24583 (N_24583,N_23178,N_23516);
xnor U24584 (N_24584,N_23672,N_23734);
nor U24585 (N_24585,N_23311,N_23184);
nor U24586 (N_24586,N_23175,N_23423);
nor U24587 (N_24587,N_23659,N_23804);
nor U24588 (N_24588,N_23142,N_23891);
xnor U24589 (N_24589,N_23230,N_23534);
xor U24590 (N_24590,N_23926,N_23556);
nand U24591 (N_24591,N_23811,N_23058);
and U24592 (N_24592,N_23245,N_23970);
xnor U24593 (N_24593,N_23410,N_23373);
and U24594 (N_24594,N_23693,N_23292);
or U24595 (N_24595,N_23389,N_23354);
nor U24596 (N_24596,N_23457,N_23116);
and U24597 (N_24597,N_23132,N_23424);
xor U24598 (N_24598,N_23038,N_23411);
nor U24599 (N_24599,N_23147,N_23122);
xnor U24600 (N_24600,N_23185,N_23652);
and U24601 (N_24601,N_23848,N_23424);
and U24602 (N_24602,N_23823,N_23988);
nor U24603 (N_24603,N_23490,N_23328);
and U24604 (N_24604,N_23811,N_23953);
nor U24605 (N_24605,N_23196,N_23995);
nor U24606 (N_24606,N_23104,N_23952);
nand U24607 (N_24607,N_23522,N_23509);
xor U24608 (N_24608,N_23363,N_23534);
or U24609 (N_24609,N_23747,N_23973);
nor U24610 (N_24610,N_23463,N_23145);
or U24611 (N_24611,N_23998,N_23873);
or U24612 (N_24612,N_23850,N_23590);
xnor U24613 (N_24613,N_23431,N_23080);
nor U24614 (N_24614,N_23356,N_23196);
nor U24615 (N_24615,N_23268,N_23195);
nand U24616 (N_24616,N_23169,N_23228);
nor U24617 (N_24617,N_23420,N_23051);
or U24618 (N_24618,N_23743,N_23882);
nand U24619 (N_24619,N_23357,N_23719);
xor U24620 (N_24620,N_23740,N_23131);
nand U24621 (N_24621,N_23025,N_23227);
or U24622 (N_24622,N_23292,N_23560);
nor U24623 (N_24623,N_23510,N_23078);
nor U24624 (N_24624,N_23085,N_23661);
nor U24625 (N_24625,N_23537,N_23997);
nor U24626 (N_24626,N_23353,N_23557);
or U24627 (N_24627,N_23745,N_23908);
or U24628 (N_24628,N_23132,N_23194);
or U24629 (N_24629,N_23821,N_23331);
xor U24630 (N_24630,N_23778,N_23649);
or U24631 (N_24631,N_23832,N_23001);
or U24632 (N_24632,N_23669,N_23060);
or U24633 (N_24633,N_23420,N_23745);
nor U24634 (N_24634,N_23843,N_23584);
nand U24635 (N_24635,N_23489,N_23680);
or U24636 (N_24636,N_23552,N_23236);
nand U24637 (N_24637,N_23235,N_23291);
or U24638 (N_24638,N_23986,N_23674);
nor U24639 (N_24639,N_23025,N_23990);
xor U24640 (N_24640,N_23594,N_23469);
nand U24641 (N_24641,N_23483,N_23405);
nand U24642 (N_24642,N_23304,N_23611);
nand U24643 (N_24643,N_23142,N_23698);
or U24644 (N_24644,N_23728,N_23485);
nand U24645 (N_24645,N_23813,N_23801);
nand U24646 (N_24646,N_23270,N_23877);
and U24647 (N_24647,N_23001,N_23631);
and U24648 (N_24648,N_23870,N_23923);
and U24649 (N_24649,N_23514,N_23076);
and U24650 (N_24650,N_23156,N_23754);
or U24651 (N_24651,N_23930,N_23031);
or U24652 (N_24652,N_23084,N_23562);
nor U24653 (N_24653,N_23747,N_23717);
nand U24654 (N_24654,N_23707,N_23571);
xnor U24655 (N_24655,N_23313,N_23553);
and U24656 (N_24656,N_23645,N_23375);
and U24657 (N_24657,N_23691,N_23159);
xor U24658 (N_24658,N_23758,N_23935);
or U24659 (N_24659,N_23829,N_23333);
nand U24660 (N_24660,N_23810,N_23825);
or U24661 (N_24661,N_23066,N_23462);
and U24662 (N_24662,N_23523,N_23738);
and U24663 (N_24663,N_23798,N_23452);
nand U24664 (N_24664,N_23483,N_23847);
or U24665 (N_24665,N_23076,N_23015);
or U24666 (N_24666,N_23554,N_23804);
nand U24667 (N_24667,N_23676,N_23933);
nand U24668 (N_24668,N_23437,N_23165);
and U24669 (N_24669,N_23642,N_23181);
nand U24670 (N_24670,N_23936,N_23825);
xor U24671 (N_24671,N_23567,N_23333);
xor U24672 (N_24672,N_23263,N_23345);
nand U24673 (N_24673,N_23337,N_23571);
nor U24674 (N_24674,N_23904,N_23958);
nor U24675 (N_24675,N_23286,N_23901);
nor U24676 (N_24676,N_23658,N_23686);
or U24677 (N_24677,N_23999,N_23742);
and U24678 (N_24678,N_23178,N_23783);
xnor U24679 (N_24679,N_23617,N_23499);
or U24680 (N_24680,N_23413,N_23746);
and U24681 (N_24681,N_23063,N_23733);
and U24682 (N_24682,N_23174,N_23274);
and U24683 (N_24683,N_23953,N_23990);
or U24684 (N_24684,N_23263,N_23126);
xnor U24685 (N_24685,N_23608,N_23142);
and U24686 (N_24686,N_23310,N_23734);
xnor U24687 (N_24687,N_23693,N_23664);
or U24688 (N_24688,N_23146,N_23427);
nand U24689 (N_24689,N_23150,N_23572);
or U24690 (N_24690,N_23760,N_23617);
nand U24691 (N_24691,N_23949,N_23331);
or U24692 (N_24692,N_23364,N_23317);
nand U24693 (N_24693,N_23863,N_23265);
or U24694 (N_24694,N_23496,N_23556);
xor U24695 (N_24695,N_23297,N_23275);
xor U24696 (N_24696,N_23707,N_23884);
and U24697 (N_24697,N_23041,N_23941);
or U24698 (N_24698,N_23578,N_23633);
and U24699 (N_24699,N_23749,N_23925);
or U24700 (N_24700,N_23150,N_23554);
nor U24701 (N_24701,N_23201,N_23911);
nor U24702 (N_24702,N_23798,N_23466);
xor U24703 (N_24703,N_23969,N_23103);
xor U24704 (N_24704,N_23281,N_23125);
nor U24705 (N_24705,N_23625,N_23014);
nand U24706 (N_24706,N_23964,N_23792);
and U24707 (N_24707,N_23589,N_23866);
or U24708 (N_24708,N_23444,N_23027);
and U24709 (N_24709,N_23414,N_23321);
or U24710 (N_24710,N_23141,N_23042);
nor U24711 (N_24711,N_23526,N_23677);
or U24712 (N_24712,N_23737,N_23438);
nand U24713 (N_24713,N_23876,N_23641);
or U24714 (N_24714,N_23700,N_23394);
nand U24715 (N_24715,N_23258,N_23856);
xor U24716 (N_24716,N_23610,N_23360);
or U24717 (N_24717,N_23115,N_23304);
and U24718 (N_24718,N_23697,N_23969);
xnor U24719 (N_24719,N_23843,N_23754);
nand U24720 (N_24720,N_23345,N_23447);
or U24721 (N_24721,N_23554,N_23708);
and U24722 (N_24722,N_23614,N_23887);
or U24723 (N_24723,N_23085,N_23002);
or U24724 (N_24724,N_23741,N_23002);
nand U24725 (N_24725,N_23360,N_23944);
nor U24726 (N_24726,N_23751,N_23329);
or U24727 (N_24727,N_23948,N_23564);
nor U24728 (N_24728,N_23862,N_23224);
and U24729 (N_24729,N_23590,N_23135);
xnor U24730 (N_24730,N_23915,N_23429);
xor U24731 (N_24731,N_23921,N_23887);
or U24732 (N_24732,N_23996,N_23524);
nor U24733 (N_24733,N_23491,N_23785);
or U24734 (N_24734,N_23817,N_23008);
nor U24735 (N_24735,N_23645,N_23231);
or U24736 (N_24736,N_23989,N_23187);
or U24737 (N_24737,N_23501,N_23680);
nor U24738 (N_24738,N_23541,N_23833);
xor U24739 (N_24739,N_23788,N_23479);
nand U24740 (N_24740,N_23848,N_23257);
xor U24741 (N_24741,N_23219,N_23232);
nand U24742 (N_24742,N_23683,N_23250);
nor U24743 (N_24743,N_23816,N_23113);
or U24744 (N_24744,N_23654,N_23034);
and U24745 (N_24745,N_23577,N_23009);
and U24746 (N_24746,N_23767,N_23880);
xor U24747 (N_24747,N_23400,N_23452);
xnor U24748 (N_24748,N_23186,N_23271);
or U24749 (N_24749,N_23375,N_23835);
nor U24750 (N_24750,N_23313,N_23358);
nor U24751 (N_24751,N_23912,N_23160);
xnor U24752 (N_24752,N_23775,N_23888);
nor U24753 (N_24753,N_23253,N_23493);
and U24754 (N_24754,N_23712,N_23925);
nand U24755 (N_24755,N_23345,N_23629);
nor U24756 (N_24756,N_23526,N_23397);
nor U24757 (N_24757,N_23353,N_23765);
xor U24758 (N_24758,N_23747,N_23207);
xnor U24759 (N_24759,N_23086,N_23214);
nand U24760 (N_24760,N_23151,N_23545);
nor U24761 (N_24761,N_23252,N_23255);
and U24762 (N_24762,N_23660,N_23851);
and U24763 (N_24763,N_23419,N_23749);
xor U24764 (N_24764,N_23444,N_23996);
xnor U24765 (N_24765,N_23941,N_23162);
nand U24766 (N_24766,N_23849,N_23091);
nand U24767 (N_24767,N_23311,N_23325);
nand U24768 (N_24768,N_23036,N_23147);
or U24769 (N_24769,N_23747,N_23485);
nand U24770 (N_24770,N_23690,N_23711);
or U24771 (N_24771,N_23750,N_23272);
or U24772 (N_24772,N_23460,N_23060);
nor U24773 (N_24773,N_23798,N_23590);
xor U24774 (N_24774,N_23927,N_23205);
or U24775 (N_24775,N_23670,N_23844);
nand U24776 (N_24776,N_23607,N_23090);
and U24777 (N_24777,N_23631,N_23827);
and U24778 (N_24778,N_23484,N_23719);
nand U24779 (N_24779,N_23187,N_23711);
or U24780 (N_24780,N_23485,N_23548);
nor U24781 (N_24781,N_23900,N_23056);
xor U24782 (N_24782,N_23202,N_23465);
xor U24783 (N_24783,N_23134,N_23630);
nand U24784 (N_24784,N_23268,N_23314);
and U24785 (N_24785,N_23583,N_23448);
or U24786 (N_24786,N_23586,N_23609);
nor U24787 (N_24787,N_23838,N_23978);
and U24788 (N_24788,N_23879,N_23605);
xnor U24789 (N_24789,N_23650,N_23579);
nor U24790 (N_24790,N_23329,N_23359);
nor U24791 (N_24791,N_23920,N_23030);
and U24792 (N_24792,N_23321,N_23709);
and U24793 (N_24793,N_23417,N_23545);
nand U24794 (N_24794,N_23961,N_23039);
or U24795 (N_24795,N_23893,N_23365);
and U24796 (N_24796,N_23550,N_23019);
nor U24797 (N_24797,N_23507,N_23405);
or U24798 (N_24798,N_23650,N_23497);
or U24799 (N_24799,N_23630,N_23517);
and U24800 (N_24800,N_23509,N_23949);
xor U24801 (N_24801,N_23570,N_23132);
xnor U24802 (N_24802,N_23652,N_23934);
nand U24803 (N_24803,N_23861,N_23856);
and U24804 (N_24804,N_23346,N_23354);
xnor U24805 (N_24805,N_23976,N_23075);
or U24806 (N_24806,N_23789,N_23610);
and U24807 (N_24807,N_23092,N_23107);
or U24808 (N_24808,N_23561,N_23533);
nand U24809 (N_24809,N_23841,N_23993);
or U24810 (N_24810,N_23944,N_23827);
nand U24811 (N_24811,N_23598,N_23288);
and U24812 (N_24812,N_23616,N_23214);
or U24813 (N_24813,N_23657,N_23647);
xnor U24814 (N_24814,N_23910,N_23321);
and U24815 (N_24815,N_23372,N_23915);
nand U24816 (N_24816,N_23652,N_23444);
xor U24817 (N_24817,N_23500,N_23676);
nor U24818 (N_24818,N_23429,N_23542);
xnor U24819 (N_24819,N_23486,N_23892);
and U24820 (N_24820,N_23212,N_23824);
or U24821 (N_24821,N_23710,N_23169);
nand U24822 (N_24822,N_23376,N_23820);
nor U24823 (N_24823,N_23805,N_23032);
nand U24824 (N_24824,N_23269,N_23934);
nor U24825 (N_24825,N_23804,N_23408);
nor U24826 (N_24826,N_23349,N_23215);
nor U24827 (N_24827,N_23966,N_23667);
nor U24828 (N_24828,N_23665,N_23311);
xor U24829 (N_24829,N_23922,N_23899);
or U24830 (N_24830,N_23580,N_23456);
or U24831 (N_24831,N_23542,N_23799);
nand U24832 (N_24832,N_23502,N_23826);
or U24833 (N_24833,N_23899,N_23845);
nor U24834 (N_24834,N_23256,N_23377);
xnor U24835 (N_24835,N_23338,N_23074);
and U24836 (N_24836,N_23039,N_23625);
nand U24837 (N_24837,N_23964,N_23074);
nor U24838 (N_24838,N_23005,N_23220);
and U24839 (N_24839,N_23752,N_23239);
or U24840 (N_24840,N_23654,N_23088);
nor U24841 (N_24841,N_23369,N_23481);
and U24842 (N_24842,N_23549,N_23810);
and U24843 (N_24843,N_23394,N_23557);
xor U24844 (N_24844,N_23466,N_23591);
xnor U24845 (N_24845,N_23472,N_23770);
xnor U24846 (N_24846,N_23580,N_23102);
and U24847 (N_24847,N_23465,N_23997);
or U24848 (N_24848,N_23655,N_23428);
xnor U24849 (N_24849,N_23648,N_23983);
nand U24850 (N_24850,N_23747,N_23263);
nor U24851 (N_24851,N_23481,N_23928);
nor U24852 (N_24852,N_23725,N_23656);
or U24853 (N_24853,N_23666,N_23339);
nand U24854 (N_24854,N_23365,N_23906);
nor U24855 (N_24855,N_23471,N_23634);
or U24856 (N_24856,N_23484,N_23931);
or U24857 (N_24857,N_23430,N_23613);
nor U24858 (N_24858,N_23598,N_23658);
or U24859 (N_24859,N_23577,N_23183);
xnor U24860 (N_24860,N_23133,N_23529);
nor U24861 (N_24861,N_23069,N_23506);
nand U24862 (N_24862,N_23413,N_23146);
nor U24863 (N_24863,N_23042,N_23129);
xor U24864 (N_24864,N_23018,N_23237);
xor U24865 (N_24865,N_23470,N_23567);
xor U24866 (N_24866,N_23922,N_23118);
nor U24867 (N_24867,N_23624,N_23733);
or U24868 (N_24868,N_23458,N_23380);
or U24869 (N_24869,N_23566,N_23960);
nand U24870 (N_24870,N_23544,N_23616);
or U24871 (N_24871,N_23202,N_23798);
or U24872 (N_24872,N_23653,N_23127);
or U24873 (N_24873,N_23320,N_23259);
nand U24874 (N_24874,N_23033,N_23599);
xnor U24875 (N_24875,N_23588,N_23993);
nand U24876 (N_24876,N_23018,N_23917);
nor U24877 (N_24877,N_23118,N_23339);
and U24878 (N_24878,N_23887,N_23176);
nand U24879 (N_24879,N_23149,N_23298);
or U24880 (N_24880,N_23401,N_23416);
and U24881 (N_24881,N_23352,N_23279);
and U24882 (N_24882,N_23124,N_23706);
nor U24883 (N_24883,N_23549,N_23012);
xnor U24884 (N_24884,N_23270,N_23511);
and U24885 (N_24885,N_23060,N_23320);
xnor U24886 (N_24886,N_23992,N_23392);
or U24887 (N_24887,N_23091,N_23181);
or U24888 (N_24888,N_23495,N_23841);
or U24889 (N_24889,N_23039,N_23465);
nor U24890 (N_24890,N_23733,N_23619);
or U24891 (N_24891,N_23312,N_23766);
nand U24892 (N_24892,N_23560,N_23273);
xnor U24893 (N_24893,N_23143,N_23907);
or U24894 (N_24894,N_23179,N_23629);
and U24895 (N_24895,N_23949,N_23193);
xor U24896 (N_24896,N_23348,N_23900);
nor U24897 (N_24897,N_23693,N_23247);
and U24898 (N_24898,N_23624,N_23281);
or U24899 (N_24899,N_23587,N_23616);
xor U24900 (N_24900,N_23849,N_23783);
and U24901 (N_24901,N_23021,N_23703);
or U24902 (N_24902,N_23894,N_23125);
nand U24903 (N_24903,N_23555,N_23484);
or U24904 (N_24904,N_23942,N_23486);
nand U24905 (N_24905,N_23454,N_23498);
nor U24906 (N_24906,N_23119,N_23160);
or U24907 (N_24907,N_23277,N_23720);
or U24908 (N_24908,N_23192,N_23312);
and U24909 (N_24909,N_23938,N_23548);
nand U24910 (N_24910,N_23962,N_23065);
nand U24911 (N_24911,N_23988,N_23270);
xnor U24912 (N_24912,N_23072,N_23722);
or U24913 (N_24913,N_23285,N_23077);
or U24914 (N_24914,N_23831,N_23879);
nor U24915 (N_24915,N_23118,N_23681);
and U24916 (N_24916,N_23320,N_23035);
xnor U24917 (N_24917,N_23791,N_23040);
nor U24918 (N_24918,N_23474,N_23957);
and U24919 (N_24919,N_23798,N_23510);
or U24920 (N_24920,N_23293,N_23037);
or U24921 (N_24921,N_23160,N_23597);
or U24922 (N_24922,N_23728,N_23112);
nand U24923 (N_24923,N_23979,N_23715);
xor U24924 (N_24924,N_23824,N_23067);
and U24925 (N_24925,N_23147,N_23542);
nand U24926 (N_24926,N_23299,N_23695);
xor U24927 (N_24927,N_23718,N_23956);
xnor U24928 (N_24928,N_23876,N_23433);
nand U24929 (N_24929,N_23912,N_23829);
or U24930 (N_24930,N_23284,N_23730);
nor U24931 (N_24931,N_23397,N_23662);
nor U24932 (N_24932,N_23200,N_23882);
nand U24933 (N_24933,N_23270,N_23334);
and U24934 (N_24934,N_23238,N_23433);
and U24935 (N_24935,N_23370,N_23357);
nand U24936 (N_24936,N_23784,N_23287);
or U24937 (N_24937,N_23516,N_23588);
or U24938 (N_24938,N_23106,N_23954);
and U24939 (N_24939,N_23586,N_23690);
nand U24940 (N_24940,N_23651,N_23249);
xor U24941 (N_24941,N_23907,N_23260);
nor U24942 (N_24942,N_23121,N_23799);
nor U24943 (N_24943,N_23309,N_23788);
or U24944 (N_24944,N_23281,N_23081);
or U24945 (N_24945,N_23994,N_23021);
nand U24946 (N_24946,N_23407,N_23498);
and U24947 (N_24947,N_23989,N_23347);
xor U24948 (N_24948,N_23651,N_23657);
nand U24949 (N_24949,N_23689,N_23072);
nor U24950 (N_24950,N_23077,N_23337);
xor U24951 (N_24951,N_23312,N_23834);
nand U24952 (N_24952,N_23086,N_23363);
nand U24953 (N_24953,N_23587,N_23735);
and U24954 (N_24954,N_23022,N_23226);
or U24955 (N_24955,N_23009,N_23753);
or U24956 (N_24956,N_23224,N_23328);
xnor U24957 (N_24957,N_23498,N_23790);
and U24958 (N_24958,N_23115,N_23349);
xor U24959 (N_24959,N_23825,N_23900);
nand U24960 (N_24960,N_23135,N_23812);
or U24961 (N_24961,N_23341,N_23875);
and U24962 (N_24962,N_23300,N_23027);
and U24963 (N_24963,N_23186,N_23918);
and U24964 (N_24964,N_23439,N_23745);
nand U24965 (N_24965,N_23162,N_23830);
nor U24966 (N_24966,N_23037,N_23189);
nand U24967 (N_24967,N_23864,N_23868);
nand U24968 (N_24968,N_23832,N_23679);
nor U24969 (N_24969,N_23447,N_23672);
and U24970 (N_24970,N_23330,N_23293);
xnor U24971 (N_24971,N_23443,N_23594);
nor U24972 (N_24972,N_23951,N_23878);
and U24973 (N_24973,N_23842,N_23353);
or U24974 (N_24974,N_23750,N_23422);
xnor U24975 (N_24975,N_23363,N_23465);
and U24976 (N_24976,N_23162,N_23882);
or U24977 (N_24977,N_23463,N_23844);
or U24978 (N_24978,N_23105,N_23220);
or U24979 (N_24979,N_23797,N_23887);
nor U24980 (N_24980,N_23766,N_23613);
nor U24981 (N_24981,N_23530,N_23927);
or U24982 (N_24982,N_23446,N_23971);
nand U24983 (N_24983,N_23890,N_23321);
nor U24984 (N_24984,N_23237,N_23501);
or U24985 (N_24985,N_23752,N_23323);
xnor U24986 (N_24986,N_23541,N_23023);
and U24987 (N_24987,N_23749,N_23969);
or U24988 (N_24988,N_23673,N_23919);
nor U24989 (N_24989,N_23113,N_23885);
nand U24990 (N_24990,N_23728,N_23629);
or U24991 (N_24991,N_23950,N_23450);
or U24992 (N_24992,N_23329,N_23196);
and U24993 (N_24993,N_23909,N_23823);
xnor U24994 (N_24994,N_23334,N_23095);
nor U24995 (N_24995,N_23548,N_23919);
nand U24996 (N_24996,N_23943,N_23629);
or U24997 (N_24997,N_23808,N_23008);
xnor U24998 (N_24998,N_23204,N_23742);
nor U24999 (N_24999,N_23422,N_23134);
nor UO_0 (O_0,N_24637,N_24424);
or UO_1 (O_1,N_24951,N_24200);
nor UO_2 (O_2,N_24716,N_24724);
nor UO_3 (O_3,N_24139,N_24158);
xor UO_4 (O_4,N_24109,N_24731);
or UO_5 (O_5,N_24062,N_24782);
or UO_6 (O_6,N_24331,N_24334);
or UO_7 (O_7,N_24464,N_24524);
or UO_8 (O_8,N_24214,N_24642);
nand UO_9 (O_9,N_24674,N_24182);
or UO_10 (O_10,N_24603,N_24579);
nor UO_11 (O_11,N_24791,N_24426);
nor UO_12 (O_12,N_24238,N_24680);
and UO_13 (O_13,N_24557,N_24648);
or UO_14 (O_14,N_24735,N_24953);
or UO_15 (O_15,N_24169,N_24691);
xnor UO_16 (O_16,N_24373,N_24185);
and UO_17 (O_17,N_24552,N_24818);
nor UO_18 (O_18,N_24343,N_24313);
nand UO_19 (O_19,N_24743,N_24228);
xor UO_20 (O_20,N_24055,N_24624);
and UO_21 (O_21,N_24088,N_24744);
xnor UO_22 (O_22,N_24177,N_24606);
and UO_23 (O_23,N_24151,N_24201);
and UO_24 (O_24,N_24895,N_24004);
or UO_25 (O_25,N_24053,N_24254);
and UO_26 (O_26,N_24502,N_24758);
xnor UO_27 (O_27,N_24654,N_24755);
nor UO_28 (O_28,N_24243,N_24087);
and UO_29 (O_29,N_24460,N_24415);
or UO_30 (O_30,N_24417,N_24566);
and UO_31 (O_31,N_24276,N_24248);
nand UO_32 (O_32,N_24006,N_24107);
nand UO_33 (O_33,N_24193,N_24310);
xor UO_34 (O_34,N_24131,N_24303);
nor UO_35 (O_35,N_24116,N_24099);
and UO_36 (O_36,N_24455,N_24219);
nand UO_37 (O_37,N_24007,N_24033);
nor UO_38 (O_38,N_24696,N_24129);
and UO_39 (O_39,N_24340,N_24559);
xor UO_40 (O_40,N_24932,N_24242);
nor UO_41 (O_41,N_24757,N_24555);
or UO_42 (O_42,N_24583,N_24830);
xor UO_43 (O_43,N_24488,N_24599);
nand UO_44 (O_44,N_24686,N_24480);
and UO_45 (O_45,N_24647,N_24733);
and UO_46 (O_46,N_24610,N_24281);
xnor UO_47 (O_47,N_24876,N_24278);
nor UO_48 (O_48,N_24536,N_24473);
nor UO_49 (O_49,N_24096,N_24226);
nand UO_50 (O_50,N_24233,N_24991);
xnor UO_51 (O_51,N_24086,N_24689);
nor UO_52 (O_52,N_24285,N_24710);
or UO_53 (O_53,N_24292,N_24179);
and UO_54 (O_54,N_24589,N_24130);
and UO_55 (O_55,N_24511,N_24348);
nand UO_56 (O_56,N_24788,N_24543);
nand UO_57 (O_57,N_24512,N_24585);
or UO_58 (O_58,N_24629,N_24225);
or UO_59 (O_59,N_24355,N_24938);
and UO_60 (O_60,N_24410,N_24890);
nand UO_61 (O_61,N_24282,N_24018);
nand UO_62 (O_62,N_24732,N_24723);
nand UO_63 (O_63,N_24729,N_24548);
nand UO_64 (O_64,N_24220,N_24100);
or UO_65 (O_65,N_24261,N_24305);
nand UO_66 (O_66,N_24293,N_24061);
xnor UO_67 (O_67,N_24121,N_24759);
and UO_68 (O_68,N_24841,N_24534);
and UO_69 (O_69,N_24584,N_24860);
or UO_70 (O_70,N_24409,N_24257);
nor UO_71 (O_71,N_24582,N_24102);
nor UO_72 (O_72,N_24147,N_24598);
nand UO_73 (O_73,N_24304,N_24259);
nor UO_74 (O_74,N_24880,N_24056);
nor UO_75 (O_75,N_24077,N_24519);
or UO_76 (O_76,N_24864,N_24644);
or UO_77 (O_77,N_24835,N_24527);
nand UO_78 (O_78,N_24176,N_24943);
nor UO_79 (O_79,N_24207,N_24309);
nor UO_80 (O_80,N_24105,N_24707);
or UO_81 (O_81,N_24588,N_24814);
or UO_82 (O_82,N_24518,N_24790);
or UO_83 (O_83,N_24150,N_24989);
xor UO_84 (O_84,N_24580,N_24154);
or UO_85 (O_85,N_24453,N_24471);
nor UO_86 (O_86,N_24551,N_24926);
nor UO_87 (O_87,N_24294,N_24570);
and UO_88 (O_88,N_24153,N_24302);
or UO_89 (O_89,N_24851,N_24380);
nor UO_90 (O_90,N_24134,N_24652);
and UO_91 (O_91,N_24392,N_24274);
xor UO_92 (O_92,N_24927,N_24314);
or UO_93 (O_93,N_24015,N_24052);
or UO_94 (O_94,N_24019,N_24117);
nand UO_95 (O_95,N_24683,N_24012);
nand UO_96 (O_96,N_24358,N_24118);
or UO_97 (O_97,N_24626,N_24039);
nand UO_98 (O_98,N_24605,N_24047);
xor UO_99 (O_99,N_24965,N_24336);
nor UO_100 (O_100,N_24553,N_24907);
xnor UO_101 (O_101,N_24750,N_24327);
and UO_102 (O_102,N_24670,N_24229);
xnor UO_103 (O_103,N_24796,N_24715);
nand UO_104 (O_104,N_24523,N_24458);
xnor UO_105 (O_105,N_24486,N_24379);
xnor UO_106 (O_106,N_24526,N_24738);
xnor UO_107 (O_107,N_24429,N_24323);
xor UO_108 (O_108,N_24998,N_24959);
and UO_109 (O_109,N_24065,N_24677);
or UO_110 (O_110,N_24060,N_24896);
xor UO_111 (O_111,N_24402,N_24728);
xor UO_112 (O_112,N_24970,N_24741);
or UO_113 (O_113,N_24122,N_24885);
xor UO_114 (O_114,N_24048,N_24252);
nor UO_115 (O_115,N_24714,N_24345);
nor UO_116 (O_116,N_24479,N_24073);
and UO_117 (O_117,N_24337,N_24286);
xor UO_118 (O_118,N_24571,N_24978);
nand UO_119 (O_119,N_24936,N_24993);
nor UO_120 (O_120,N_24772,N_24263);
or UO_121 (O_121,N_24525,N_24298);
or UO_122 (O_122,N_24789,N_24399);
and UO_123 (O_123,N_24645,N_24866);
or UO_124 (O_124,N_24808,N_24217);
nor UO_125 (O_125,N_24316,N_24847);
xnor UO_126 (O_126,N_24240,N_24776);
and UO_127 (O_127,N_24903,N_24187);
xnor UO_128 (O_128,N_24522,N_24889);
or UO_129 (O_129,N_24563,N_24204);
xnor UO_130 (O_130,N_24748,N_24668);
nand UO_131 (O_131,N_24747,N_24958);
nand UO_132 (O_132,N_24416,N_24403);
or UO_133 (O_133,N_24195,N_24875);
or UO_134 (O_134,N_24465,N_24940);
or UO_135 (O_135,N_24820,N_24308);
and UO_136 (O_136,N_24492,N_24752);
xnor UO_137 (O_137,N_24126,N_24597);
xor UO_138 (O_138,N_24300,N_24886);
nor UO_139 (O_139,N_24663,N_24699);
nand UO_140 (O_140,N_24690,N_24974);
nor UO_141 (O_141,N_24547,N_24350);
xnor UO_142 (O_142,N_24203,N_24725);
or UO_143 (O_143,N_24858,N_24709);
xor UO_144 (O_144,N_24095,N_24852);
nand UO_145 (O_145,N_24844,N_24838);
or UO_146 (O_146,N_24024,N_24608);
or UO_147 (O_147,N_24985,N_24009);
and UO_148 (O_148,N_24171,N_24956);
xnor UO_149 (O_149,N_24786,N_24672);
and UO_150 (O_150,N_24156,N_24070);
xnor UO_151 (O_151,N_24110,N_24250);
and UO_152 (O_152,N_24387,N_24516);
nand UO_153 (O_153,N_24661,N_24028);
nand UO_154 (O_154,N_24863,N_24344);
nor UO_155 (O_155,N_24658,N_24255);
nand UO_156 (O_156,N_24166,N_24705);
nor UO_157 (O_157,N_24703,N_24478);
and UO_158 (O_158,N_24135,N_24635);
and UO_159 (O_159,N_24448,N_24010);
or UO_160 (O_160,N_24942,N_24438);
or UO_161 (O_161,N_24587,N_24155);
or UO_162 (O_162,N_24720,N_24262);
and UO_163 (O_163,N_24237,N_24990);
xor UO_164 (O_164,N_24627,N_24630);
nand UO_165 (O_165,N_24421,N_24325);
and UO_166 (O_166,N_24470,N_24769);
nor UO_167 (O_167,N_24374,N_24422);
or UO_168 (O_168,N_24961,N_24829);
nand UO_169 (O_169,N_24981,N_24142);
xnor UO_170 (O_170,N_24036,N_24817);
nor UO_171 (O_171,N_24545,N_24873);
or UO_172 (O_172,N_24919,N_24020);
nand UO_173 (O_173,N_24489,N_24145);
and UO_174 (O_174,N_24490,N_24218);
nor UO_175 (O_175,N_24430,N_24827);
xnor UO_176 (O_176,N_24454,N_24602);
and UO_177 (O_177,N_24538,N_24550);
xnor UO_178 (O_178,N_24591,N_24939);
xnor UO_179 (O_179,N_24022,N_24681);
xnor UO_180 (O_180,N_24918,N_24045);
nor UO_181 (O_181,N_24870,N_24666);
and UO_182 (O_182,N_24468,N_24891);
or UO_183 (O_183,N_24026,N_24013);
nand UO_184 (O_184,N_24042,N_24211);
or UO_185 (O_185,N_24862,N_24495);
or UO_186 (O_186,N_24955,N_24208);
or UO_187 (O_187,N_24616,N_24562);
xnor UO_188 (O_188,N_24832,N_24071);
xor UO_189 (O_189,N_24722,N_24567);
nand UO_190 (O_190,N_24843,N_24299);
nor UO_191 (O_191,N_24418,N_24290);
and UO_192 (O_192,N_24157,N_24655);
nand UO_193 (O_193,N_24615,N_24797);
nand UO_194 (O_194,N_24330,N_24698);
or UO_195 (O_195,N_24520,N_24718);
or UO_196 (O_196,N_24123,N_24848);
xnor UO_197 (O_197,N_24329,N_24877);
nor UO_198 (O_198,N_24914,N_24452);
nand UO_199 (O_199,N_24785,N_24834);
xor UO_200 (O_200,N_24349,N_24819);
or UO_201 (O_201,N_24030,N_24143);
or UO_202 (O_202,N_24287,N_24528);
xnor UO_203 (O_203,N_24736,N_24529);
xor UO_204 (O_204,N_24114,N_24979);
nor UO_205 (O_205,N_24081,N_24572);
xnor UO_206 (O_206,N_24364,N_24702);
and UO_207 (O_207,N_24717,N_24692);
or UO_208 (O_208,N_24920,N_24236);
nor UO_209 (O_209,N_24186,N_24879);
and UO_210 (O_210,N_24641,N_24427);
xnor UO_211 (O_211,N_24215,N_24172);
nor UO_212 (O_212,N_24678,N_24335);
and UO_213 (O_213,N_24771,N_24366);
and UO_214 (O_214,N_24106,N_24962);
nor UO_215 (O_215,N_24569,N_24221);
nand UO_216 (O_216,N_24206,N_24230);
xnor UO_217 (O_217,N_24734,N_24016);
xor UO_218 (O_218,N_24390,N_24662);
or UO_219 (O_219,N_24108,N_24167);
or UO_220 (O_220,N_24777,N_24173);
nand UO_221 (O_221,N_24398,N_24017);
or UO_222 (O_222,N_24611,N_24934);
xnor UO_223 (O_223,N_24513,N_24533);
nand UO_224 (O_224,N_24191,N_24685);
xnor UO_225 (O_225,N_24368,N_24556);
nor UO_226 (O_226,N_24800,N_24887);
or UO_227 (O_227,N_24425,N_24963);
or UO_228 (O_228,N_24216,N_24499);
nor UO_229 (O_229,N_24778,N_24968);
nor UO_230 (O_230,N_24174,N_24804);
or UO_231 (O_231,N_24450,N_24621);
nor UO_232 (O_232,N_24811,N_24531);
or UO_233 (O_233,N_24894,N_24609);
xnor UO_234 (O_234,N_24952,N_24651);
xnor UO_235 (O_235,N_24183,N_24011);
nand UO_236 (O_236,N_24631,N_24269);
and UO_237 (O_237,N_24745,N_24423);
xnor UO_238 (O_238,N_24124,N_24833);
or UO_239 (O_239,N_24083,N_24377);
or UO_240 (O_240,N_24754,N_24049);
nor UO_241 (O_241,N_24773,N_24136);
or UO_242 (O_242,N_24023,N_24224);
nand UO_243 (O_243,N_24456,N_24370);
nand UO_244 (O_244,N_24359,N_24872);
and UO_245 (O_245,N_24202,N_24823);
nor UO_246 (O_246,N_24498,N_24069);
or UO_247 (O_247,N_24669,N_24035);
nand UO_248 (O_248,N_24266,N_24021);
nor UO_249 (O_249,N_24149,N_24138);
nor UO_250 (O_250,N_24600,N_24044);
and UO_251 (O_251,N_24535,N_24002);
and UO_252 (O_252,N_24477,N_24483);
nor UO_253 (O_253,N_24072,N_24439);
xor UO_254 (O_254,N_24446,N_24148);
and UO_255 (O_255,N_24988,N_24507);
and UO_256 (O_256,N_24144,N_24950);
and UO_257 (O_257,N_24159,N_24311);
or UO_258 (O_258,N_24029,N_24774);
xor UO_259 (O_259,N_24500,N_24270);
nor UO_260 (O_260,N_24251,N_24892);
xnor UO_261 (O_261,N_24924,N_24175);
and UO_262 (O_262,N_24713,N_24063);
or UO_263 (O_263,N_24840,N_24941);
nor UO_264 (O_264,N_24098,N_24394);
xor UO_265 (O_265,N_24494,N_24781);
or UO_266 (O_266,N_24431,N_24319);
nor UO_267 (O_267,N_24120,N_24997);
nand UO_268 (O_268,N_24068,N_24440);
or UO_269 (O_269,N_24893,N_24813);
and UO_270 (O_270,N_24901,N_24493);
xnor UO_271 (O_271,N_24568,N_24501);
xnor UO_272 (O_272,N_24405,N_24103);
xor UO_273 (O_273,N_24184,N_24372);
nand UO_274 (O_274,N_24265,N_24937);
nor UO_275 (O_275,N_24321,N_24161);
nor UO_276 (O_276,N_24764,N_24592);
nor UO_277 (O_277,N_24697,N_24613);
nor UO_278 (O_278,N_24104,N_24995);
nand UO_279 (O_279,N_24196,N_24090);
nand UO_280 (O_280,N_24256,N_24246);
nor UO_281 (O_281,N_24816,N_24982);
xor UO_282 (O_282,N_24910,N_24444);
and UO_283 (O_283,N_24595,N_24761);
nand UO_284 (O_284,N_24646,N_24354);
nor UO_285 (O_285,N_24442,N_24428);
nor UO_286 (O_286,N_24854,N_24869);
xnor UO_287 (O_287,N_24280,N_24971);
or UO_288 (O_288,N_24622,N_24760);
xor UO_289 (O_289,N_24317,N_24980);
nor UO_290 (O_290,N_24115,N_24165);
xor UO_291 (O_291,N_24593,N_24451);
nand UO_292 (O_292,N_24730,N_24544);
and UO_293 (O_293,N_24649,N_24882);
nand UO_294 (O_294,N_24180,N_24521);
nand UO_295 (O_295,N_24333,N_24235);
xnor UO_296 (O_296,N_24362,N_24874);
xnor UO_297 (O_297,N_24917,N_24043);
and UO_298 (O_298,N_24815,N_24381);
nor UO_299 (O_299,N_24515,N_24849);
and UO_300 (O_300,N_24753,N_24388);
and UO_301 (O_301,N_24749,N_24393);
and UO_302 (O_302,N_24828,N_24638);
nand UO_303 (O_303,N_24085,N_24911);
and UO_304 (O_304,N_24633,N_24667);
xor UO_305 (O_305,N_24284,N_24945);
nand UO_306 (O_306,N_24227,N_24435);
nand UO_307 (O_307,N_24821,N_24487);
nand UO_308 (O_308,N_24482,N_24315);
xor UO_309 (O_309,N_24897,N_24966);
xor UO_310 (O_310,N_24969,N_24532);
xnor UO_311 (O_311,N_24565,N_24855);
xnor UO_312 (O_312,N_24058,N_24367);
and UO_313 (O_313,N_24443,N_24283);
xor UO_314 (O_314,N_24767,N_24798);
nor UO_315 (O_315,N_24682,N_24857);
nor UO_316 (O_316,N_24384,N_24922);
and UO_317 (O_317,N_24967,N_24375);
nor UO_318 (O_318,N_24389,N_24484);
nor UO_319 (O_319,N_24701,N_24825);
xor UO_320 (O_320,N_24436,N_24000);
or UO_321 (O_321,N_24931,N_24719);
nor UO_322 (O_322,N_24476,N_24619);
and UO_323 (O_323,N_24809,N_24558);
xor UO_324 (O_324,N_24996,N_24365);
or UO_325 (O_325,N_24322,N_24383);
or UO_326 (O_326,N_24742,N_24306);
nand UO_327 (O_327,N_24496,N_24594);
nor UO_328 (O_328,N_24222,N_24093);
nand UO_329 (O_329,N_24168,N_24746);
nand UO_330 (O_330,N_24008,N_24395);
nand UO_331 (O_331,N_24445,N_24244);
or UO_332 (O_332,N_24210,N_24064);
xor UO_333 (O_333,N_24092,N_24923);
or UO_334 (O_334,N_24360,N_24868);
and UO_335 (O_335,N_24846,N_24091);
nand UO_336 (O_336,N_24295,N_24067);
xor UO_337 (O_337,N_24101,N_24141);
nand UO_338 (O_338,N_24768,N_24447);
nand UO_339 (O_339,N_24080,N_24801);
nor UO_340 (O_340,N_24462,N_24721);
or UO_341 (O_341,N_24904,N_24051);
or UO_342 (O_342,N_24999,N_24273);
or UO_343 (O_343,N_24653,N_24260);
or UO_344 (O_344,N_24947,N_24059);
or UO_345 (O_345,N_24657,N_24539);
nand UO_346 (O_346,N_24188,N_24032);
or UO_347 (O_347,N_24839,N_24112);
xor UO_348 (O_348,N_24906,N_24170);
nand UO_349 (O_349,N_24472,N_24933);
nor UO_350 (O_350,N_24277,N_24807);
xnor UO_351 (O_351,N_24793,N_24137);
and UO_352 (O_352,N_24419,N_24756);
xnor UO_353 (O_353,N_24089,N_24400);
and UO_354 (O_354,N_24842,N_24806);
and UO_355 (O_355,N_24695,N_24604);
and UO_356 (O_356,N_24614,N_24612);
nand UO_357 (O_357,N_24915,N_24671);
nand UO_358 (O_358,N_24617,N_24412);
nand UO_359 (O_359,N_24296,N_24312);
nor UO_360 (O_360,N_24510,N_24034);
and UO_361 (O_361,N_24643,N_24461);
nor UO_362 (O_362,N_24066,N_24706);
xor UO_363 (O_363,N_24027,N_24025);
xnor UO_364 (O_364,N_24795,N_24618);
or UO_365 (O_365,N_24656,N_24948);
xnor UO_366 (O_366,N_24766,N_24075);
and UO_367 (O_367,N_24930,N_24128);
nor UO_368 (O_368,N_24258,N_24659);
xor UO_369 (O_369,N_24094,N_24577);
xnor UO_370 (O_370,N_24992,N_24765);
nor UO_371 (O_371,N_24113,N_24332);
and UO_372 (O_372,N_24459,N_24382);
nor UO_373 (O_373,N_24057,N_24783);
nand UO_374 (O_374,N_24132,N_24625);
or UO_375 (O_375,N_24822,N_24537);
and UO_376 (O_376,N_24046,N_24983);
nand UO_377 (O_377,N_24779,N_24223);
nor UO_378 (O_378,N_24181,N_24209);
and UO_379 (O_379,N_24506,N_24883);
or UO_380 (O_380,N_24178,N_24636);
nand UO_381 (O_381,N_24975,N_24038);
or UO_382 (O_382,N_24576,N_24560);
nor UO_383 (O_383,N_24420,N_24554);
or UO_384 (O_384,N_24687,N_24639);
nand UO_385 (O_385,N_24245,N_24711);
and UO_386 (O_386,N_24197,N_24307);
or UO_387 (O_387,N_24908,N_24198);
xnor UO_388 (O_388,N_24799,N_24751);
or UO_389 (O_389,N_24386,N_24632);
and UO_390 (O_390,N_24688,N_24014);
nand UO_391 (O_391,N_24469,N_24546);
nand UO_392 (O_392,N_24984,N_24272);
and UO_393 (O_393,N_24378,N_24739);
xor UO_394 (O_394,N_24407,N_24318);
and UO_395 (O_395,N_24954,N_24964);
nor UO_396 (O_396,N_24347,N_24865);
or UO_397 (O_397,N_24385,N_24912);
nor UO_398 (O_398,N_24628,N_24003);
nor UO_399 (O_399,N_24623,N_24291);
xor UO_400 (O_400,N_24737,N_24794);
xor UO_401 (O_401,N_24935,N_24867);
and UO_402 (O_402,N_24054,N_24530);
and UO_403 (O_403,N_24700,N_24665);
nor UO_404 (O_404,N_24346,N_24376);
and UO_405 (O_405,N_24212,N_24727);
xor UO_406 (O_406,N_24944,N_24900);
or UO_407 (O_407,N_24726,N_24986);
nand UO_408 (O_408,N_24859,N_24925);
nand UO_409 (O_409,N_24084,N_24660);
nand UO_410 (O_410,N_24960,N_24780);
xnor UO_411 (O_411,N_24357,N_24005);
or UO_412 (O_412,N_24957,N_24973);
and UO_413 (O_413,N_24271,N_24239);
and UO_414 (O_414,N_24850,N_24561);
nor UO_415 (O_415,N_24152,N_24921);
xnor UO_416 (O_416,N_24987,N_24119);
and UO_417 (O_417,N_24856,N_24397);
nand UO_418 (O_418,N_24762,N_24485);
and UO_419 (O_419,N_24342,N_24232);
or UO_420 (O_420,N_24491,N_24297);
nand UO_421 (O_421,N_24845,N_24481);
and UO_422 (O_422,N_24837,N_24763);
and UO_423 (O_423,N_24467,N_24404);
or UO_424 (O_424,N_24163,N_24508);
xnor UO_425 (O_425,N_24916,N_24573);
nor UO_426 (O_426,N_24497,N_24884);
nor UO_427 (O_427,N_24503,N_24275);
and UO_428 (O_428,N_24433,N_24474);
or UO_429 (O_429,N_24434,N_24871);
or UO_430 (O_430,N_24338,N_24740);
nand UO_431 (O_431,N_24929,N_24601);
nor UO_432 (O_432,N_24363,N_24127);
nand UO_433 (O_433,N_24810,N_24812);
nor UO_434 (O_434,N_24457,N_24339);
and UO_435 (O_435,N_24205,N_24432);
nor UO_436 (O_436,N_24712,N_24898);
or UO_437 (O_437,N_24162,N_24268);
nand UO_438 (O_438,N_24775,N_24082);
nand UO_439 (O_439,N_24231,N_24463);
xnor UO_440 (O_440,N_24356,N_24040);
nand UO_441 (O_441,N_24192,N_24234);
and UO_442 (O_442,N_24074,N_24352);
or UO_443 (O_443,N_24902,N_24437);
nor UO_444 (O_444,N_24972,N_24041);
nand UO_445 (O_445,N_24111,N_24140);
or UO_446 (O_446,N_24078,N_24351);
xnor UO_447 (O_447,N_24640,N_24289);
and UO_448 (O_448,N_24001,N_24684);
nor UO_449 (O_449,N_24946,N_24301);
or UO_450 (O_450,N_24792,N_24586);
nand UO_451 (O_451,N_24578,N_24575);
and UO_452 (O_452,N_24802,N_24320);
xor UO_453 (O_453,N_24194,N_24160);
nor UO_454 (O_454,N_24353,N_24596);
and UO_455 (O_455,N_24590,N_24694);
or UO_456 (O_456,N_24878,N_24213);
nor UO_457 (O_457,N_24441,N_24475);
nand UO_458 (O_458,N_24803,N_24391);
and UO_459 (O_459,N_24133,N_24564);
and UO_460 (O_460,N_24037,N_24634);
or UO_461 (O_461,N_24977,N_24414);
xor UO_462 (O_462,N_24976,N_24831);
nand UO_463 (O_463,N_24264,N_24267);
nor UO_464 (O_464,N_24411,N_24199);
and UO_465 (O_465,N_24836,N_24581);
and UO_466 (O_466,N_24704,N_24861);
xor UO_467 (O_467,N_24241,N_24324);
nand UO_468 (O_468,N_24881,N_24664);
nand UO_469 (O_469,N_24371,N_24189);
xnor UO_470 (O_470,N_24909,N_24899);
and UO_471 (O_471,N_24369,N_24288);
or UO_472 (O_472,N_24514,N_24824);
or UO_473 (O_473,N_24050,N_24505);
xor UO_474 (O_474,N_24517,N_24253);
or UO_475 (O_475,N_24328,N_24249);
and UO_476 (O_476,N_24408,N_24650);
or UO_477 (O_477,N_24466,N_24361);
or UO_478 (O_478,N_24949,N_24449);
and UO_479 (O_479,N_24190,N_24125);
nand UO_480 (O_480,N_24787,N_24574);
nand UO_481 (O_481,N_24994,N_24279);
nand UO_482 (O_482,N_24541,N_24905);
xor UO_483 (O_483,N_24675,N_24031);
or UO_484 (O_484,N_24888,N_24784);
nand UO_485 (O_485,N_24326,N_24247);
nor UO_486 (O_486,N_24549,N_24805);
or UO_487 (O_487,N_24913,N_24164);
nor UO_488 (O_488,N_24401,N_24079);
or UO_489 (O_489,N_24540,N_24770);
xnor UO_490 (O_490,N_24673,N_24693);
xor UO_491 (O_491,N_24076,N_24679);
and UO_492 (O_492,N_24826,N_24676);
and UO_493 (O_493,N_24542,N_24341);
and UO_494 (O_494,N_24607,N_24853);
xnor UO_495 (O_495,N_24097,N_24406);
xor UO_496 (O_496,N_24504,N_24708);
nor UO_497 (O_497,N_24620,N_24396);
xor UO_498 (O_498,N_24413,N_24146);
xnor UO_499 (O_499,N_24928,N_24509);
or UO_500 (O_500,N_24254,N_24626);
and UO_501 (O_501,N_24894,N_24716);
xnor UO_502 (O_502,N_24238,N_24525);
or UO_503 (O_503,N_24853,N_24229);
nor UO_504 (O_504,N_24365,N_24363);
nand UO_505 (O_505,N_24484,N_24915);
and UO_506 (O_506,N_24646,N_24195);
and UO_507 (O_507,N_24453,N_24954);
nand UO_508 (O_508,N_24757,N_24114);
nand UO_509 (O_509,N_24573,N_24031);
nand UO_510 (O_510,N_24253,N_24910);
nor UO_511 (O_511,N_24041,N_24839);
nand UO_512 (O_512,N_24067,N_24124);
and UO_513 (O_513,N_24650,N_24251);
or UO_514 (O_514,N_24782,N_24549);
xnor UO_515 (O_515,N_24343,N_24797);
nand UO_516 (O_516,N_24586,N_24972);
and UO_517 (O_517,N_24454,N_24373);
and UO_518 (O_518,N_24237,N_24023);
or UO_519 (O_519,N_24719,N_24668);
xnor UO_520 (O_520,N_24090,N_24988);
or UO_521 (O_521,N_24909,N_24218);
nand UO_522 (O_522,N_24891,N_24174);
or UO_523 (O_523,N_24986,N_24576);
nor UO_524 (O_524,N_24713,N_24353);
or UO_525 (O_525,N_24406,N_24383);
nand UO_526 (O_526,N_24610,N_24286);
xor UO_527 (O_527,N_24817,N_24076);
or UO_528 (O_528,N_24416,N_24463);
nand UO_529 (O_529,N_24635,N_24418);
nand UO_530 (O_530,N_24993,N_24531);
nand UO_531 (O_531,N_24037,N_24832);
nor UO_532 (O_532,N_24920,N_24623);
xor UO_533 (O_533,N_24365,N_24342);
or UO_534 (O_534,N_24741,N_24405);
and UO_535 (O_535,N_24587,N_24507);
or UO_536 (O_536,N_24818,N_24932);
nor UO_537 (O_537,N_24416,N_24189);
and UO_538 (O_538,N_24094,N_24488);
and UO_539 (O_539,N_24919,N_24335);
nor UO_540 (O_540,N_24316,N_24133);
or UO_541 (O_541,N_24734,N_24844);
and UO_542 (O_542,N_24763,N_24883);
or UO_543 (O_543,N_24411,N_24251);
nor UO_544 (O_544,N_24762,N_24193);
and UO_545 (O_545,N_24176,N_24338);
nor UO_546 (O_546,N_24225,N_24199);
or UO_547 (O_547,N_24844,N_24686);
and UO_548 (O_548,N_24849,N_24339);
nand UO_549 (O_549,N_24064,N_24336);
or UO_550 (O_550,N_24711,N_24359);
or UO_551 (O_551,N_24569,N_24519);
nor UO_552 (O_552,N_24093,N_24911);
xor UO_553 (O_553,N_24780,N_24129);
nor UO_554 (O_554,N_24874,N_24538);
and UO_555 (O_555,N_24636,N_24689);
or UO_556 (O_556,N_24819,N_24983);
nor UO_557 (O_557,N_24100,N_24223);
and UO_558 (O_558,N_24530,N_24669);
and UO_559 (O_559,N_24582,N_24205);
nor UO_560 (O_560,N_24241,N_24773);
nor UO_561 (O_561,N_24160,N_24137);
or UO_562 (O_562,N_24011,N_24214);
nand UO_563 (O_563,N_24311,N_24721);
xor UO_564 (O_564,N_24218,N_24784);
nand UO_565 (O_565,N_24737,N_24357);
or UO_566 (O_566,N_24905,N_24136);
and UO_567 (O_567,N_24059,N_24317);
nand UO_568 (O_568,N_24788,N_24642);
xnor UO_569 (O_569,N_24198,N_24118);
nor UO_570 (O_570,N_24818,N_24726);
nor UO_571 (O_571,N_24874,N_24967);
nand UO_572 (O_572,N_24110,N_24970);
nor UO_573 (O_573,N_24756,N_24138);
nand UO_574 (O_574,N_24223,N_24910);
and UO_575 (O_575,N_24709,N_24414);
nand UO_576 (O_576,N_24141,N_24755);
and UO_577 (O_577,N_24093,N_24565);
xnor UO_578 (O_578,N_24116,N_24819);
and UO_579 (O_579,N_24147,N_24145);
xnor UO_580 (O_580,N_24775,N_24317);
nand UO_581 (O_581,N_24728,N_24841);
or UO_582 (O_582,N_24314,N_24709);
nor UO_583 (O_583,N_24685,N_24789);
or UO_584 (O_584,N_24431,N_24656);
and UO_585 (O_585,N_24701,N_24305);
xnor UO_586 (O_586,N_24815,N_24527);
xnor UO_587 (O_587,N_24917,N_24615);
and UO_588 (O_588,N_24126,N_24233);
nand UO_589 (O_589,N_24148,N_24335);
or UO_590 (O_590,N_24419,N_24467);
xor UO_591 (O_591,N_24385,N_24786);
nand UO_592 (O_592,N_24522,N_24246);
xor UO_593 (O_593,N_24543,N_24694);
xor UO_594 (O_594,N_24593,N_24181);
or UO_595 (O_595,N_24263,N_24106);
nand UO_596 (O_596,N_24660,N_24495);
nand UO_597 (O_597,N_24190,N_24176);
and UO_598 (O_598,N_24982,N_24936);
and UO_599 (O_599,N_24292,N_24191);
nor UO_600 (O_600,N_24325,N_24670);
nor UO_601 (O_601,N_24433,N_24068);
or UO_602 (O_602,N_24735,N_24983);
or UO_603 (O_603,N_24196,N_24446);
xnor UO_604 (O_604,N_24929,N_24612);
and UO_605 (O_605,N_24762,N_24701);
and UO_606 (O_606,N_24098,N_24318);
and UO_607 (O_607,N_24560,N_24991);
and UO_608 (O_608,N_24254,N_24795);
nand UO_609 (O_609,N_24154,N_24590);
and UO_610 (O_610,N_24050,N_24798);
nand UO_611 (O_611,N_24923,N_24592);
nor UO_612 (O_612,N_24939,N_24422);
xor UO_613 (O_613,N_24558,N_24284);
nor UO_614 (O_614,N_24510,N_24659);
nand UO_615 (O_615,N_24051,N_24188);
nor UO_616 (O_616,N_24519,N_24743);
nand UO_617 (O_617,N_24024,N_24070);
nor UO_618 (O_618,N_24642,N_24124);
or UO_619 (O_619,N_24218,N_24223);
and UO_620 (O_620,N_24678,N_24041);
or UO_621 (O_621,N_24493,N_24550);
and UO_622 (O_622,N_24834,N_24685);
xnor UO_623 (O_623,N_24497,N_24516);
and UO_624 (O_624,N_24727,N_24229);
xor UO_625 (O_625,N_24756,N_24206);
xor UO_626 (O_626,N_24669,N_24867);
xnor UO_627 (O_627,N_24182,N_24885);
nor UO_628 (O_628,N_24708,N_24565);
nor UO_629 (O_629,N_24718,N_24690);
and UO_630 (O_630,N_24117,N_24974);
nor UO_631 (O_631,N_24051,N_24771);
or UO_632 (O_632,N_24089,N_24344);
and UO_633 (O_633,N_24457,N_24367);
nor UO_634 (O_634,N_24956,N_24066);
nand UO_635 (O_635,N_24690,N_24993);
or UO_636 (O_636,N_24086,N_24939);
nor UO_637 (O_637,N_24911,N_24737);
or UO_638 (O_638,N_24915,N_24119);
xnor UO_639 (O_639,N_24176,N_24934);
xor UO_640 (O_640,N_24953,N_24348);
nand UO_641 (O_641,N_24580,N_24748);
nor UO_642 (O_642,N_24455,N_24794);
nor UO_643 (O_643,N_24740,N_24836);
and UO_644 (O_644,N_24981,N_24466);
nor UO_645 (O_645,N_24599,N_24603);
nand UO_646 (O_646,N_24504,N_24883);
or UO_647 (O_647,N_24693,N_24366);
or UO_648 (O_648,N_24792,N_24475);
or UO_649 (O_649,N_24522,N_24569);
xor UO_650 (O_650,N_24497,N_24267);
and UO_651 (O_651,N_24027,N_24473);
nand UO_652 (O_652,N_24743,N_24608);
or UO_653 (O_653,N_24949,N_24895);
and UO_654 (O_654,N_24525,N_24150);
xnor UO_655 (O_655,N_24391,N_24487);
xnor UO_656 (O_656,N_24230,N_24415);
and UO_657 (O_657,N_24213,N_24205);
xnor UO_658 (O_658,N_24691,N_24051);
nor UO_659 (O_659,N_24770,N_24895);
nor UO_660 (O_660,N_24765,N_24890);
or UO_661 (O_661,N_24332,N_24931);
xnor UO_662 (O_662,N_24009,N_24493);
nand UO_663 (O_663,N_24310,N_24323);
nor UO_664 (O_664,N_24502,N_24432);
and UO_665 (O_665,N_24561,N_24713);
or UO_666 (O_666,N_24762,N_24341);
nand UO_667 (O_667,N_24015,N_24498);
nor UO_668 (O_668,N_24655,N_24642);
xor UO_669 (O_669,N_24660,N_24858);
nor UO_670 (O_670,N_24301,N_24196);
xnor UO_671 (O_671,N_24399,N_24877);
nand UO_672 (O_672,N_24541,N_24612);
or UO_673 (O_673,N_24299,N_24856);
xor UO_674 (O_674,N_24388,N_24482);
and UO_675 (O_675,N_24548,N_24421);
nand UO_676 (O_676,N_24535,N_24970);
and UO_677 (O_677,N_24604,N_24894);
xnor UO_678 (O_678,N_24665,N_24618);
nor UO_679 (O_679,N_24695,N_24574);
xor UO_680 (O_680,N_24630,N_24931);
xnor UO_681 (O_681,N_24468,N_24238);
or UO_682 (O_682,N_24393,N_24281);
and UO_683 (O_683,N_24780,N_24375);
nand UO_684 (O_684,N_24148,N_24465);
nand UO_685 (O_685,N_24907,N_24352);
nand UO_686 (O_686,N_24017,N_24712);
nor UO_687 (O_687,N_24111,N_24210);
and UO_688 (O_688,N_24259,N_24663);
xnor UO_689 (O_689,N_24189,N_24757);
and UO_690 (O_690,N_24133,N_24299);
or UO_691 (O_691,N_24985,N_24861);
nand UO_692 (O_692,N_24284,N_24221);
or UO_693 (O_693,N_24654,N_24647);
nor UO_694 (O_694,N_24487,N_24298);
xnor UO_695 (O_695,N_24184,N_24649);
or UO_696 (O_696,N_24399,N_24311);
xnor UO_697 (O_697,N_24955,N_24554);
and UO_698 (O_698,N_24627,N_24064);
nand UO_699 (O_699,N_24086,N_24710);
or UO_700 (O_700,N_24734,N_24930);
or UO_701 (O_701,N_24507,N_24039);
xor UO_702 (O_702,N_24834,N_24381);
xnor UO_703 (O_703,N_24622,N_24159);
and UO_704 (O_704,N_24750,N_24234);
or UO_705 (O_705,N_24288,N_24988);
nor UO_706 (O_706,N_24755,N_24020);
xnor UO_707 (O_707,N_24004,N_24752);
and UO_708 (O_708,N_24655,N_24136);
and UO_709 (O_709,N_24725,N_24103);
nand UO_710 (O_710,N_24558,N_24752);
and UO_711 (O_711,N_24498,N_24501);
or UO_712 (O_712,N_24314,N_24256);
and UO_713 (O_713,N_24306,N_24510);
and UO_714 (O_714,N_24335,N_24224);
and UO_715 (O_715,N_24684,N_24798);
nand UO_716 (O_716,N_24794,N_24626);
nand UO_717 (O_717,N_24711,N_24200);
or UO_718 (O_718,N_24534,N_24911);
or UO_719 (O_719,N_24478,N_24943);
nand UO_720 (O_720,N_24689,N_24504);
and UO_721 (O_721,N_24533,N_24566);
xor UO_722 (O_722,N_24406,N_24012);
xnor UO_723 (O_723,N_24293,N_24968);
nand UO_724 (O_724,N_24204,N_24519);
nor UO_725 (O_725,N_24243,N_24319);
or UO_726 (O_726,N_24321,N_24847);
and UO_727 (O_727,N_24032,N_24975);
or UO_728 (O_728,N_24711,N_24840);
xnor UO_729 (O_729,N_24143,N_24574);
nor UO_730 (O_730,N_24125,N_24483);
xnor UO_731 (O_731,N_24410,N_24124);
nand UO_732 (O_732,N_24595,N_24520);
xor UO_733 (O_733,N_24188,N_24219);
nor UO_734 (O_734,N_24690,N_24106);
nand UO_735 (O_735,N_24377,N_24830);
or UO_736 (O_736,N_24099,N_24294);
xnor UO_737 (O_737,N_24942,N_24450);
nand UO_738 (O_738,N_24312,N_24009);
or UO_739 (O_739,N_24934,N_24827);
nand UO_740 (O_740,N_24488,N_24584);
xor UO_741 (O_741,N_24137,N_24769);
nand UO_742 (O_742,N_24808,N_24034);
and UO_743 (O_743,N_24167,N_24352);
nor UO_744 (O_744,N_24614,N_24469);
nor UO_745 (O_745,N_24969,N_24940);
nor UO_746 (O_746,N_24971,N_24408);
nand UO_747 (O_747,N_24440,N_24860);
nand UO_748 (O_748,N_24452,N_24538);
nor UO_749 (O_749,N_24734,N_24129);
or UO_750 (O_750,N_24886,N_24307);
xnor UO_751 (O_751,N_24685,N_24523);
xnor UO_752 (O_752,N_24744,N_24659);
and UO_753 (O_753,N_24384,N_24744);
xor UO_754 (O_754,N_24125,N_24003);
and UO_755 (O_755,N_24156,N_24328);
nor UO_756 (O_756,N_24705,N_24469);
nor UO_757 (O_757,N_24353,N_24414);
and UO_758 (O_758,N_24617,N_24493);
and UO_759 (O_759,N_24803,N_24508);
xor UO_760 (O_760,N_24135,N_24720);
or UO_761 (O_761,N_24030,N_24396);
nor UO_762 (O_762,N_24629,N_24543);
nand UO_763 (O_763,N_24641,N_24719);
nor UO_764 (O_764,N_24945,N_24750);
and UO_765 (O_765,N_24276,N_24709);
nor UO_766 (O_766,N_24128,N_24938);
and UO_767 (O_767,N_24612,N_24307);
nor UO_768 (O_768,N_24795,N_24609);
xnor UO_769 (O_769,N_24845,N_24790);
or UO_770 (O_770,N_24771,N_24847);
xnor UO_771 (O_771,N_24324,N_24518);
or UO_772 (O_772,N_24506,N_24497);
nand UO_773 (O_773,N_24158,N_24111);
nor UO_774 (O_774,N_24815,N_24021);
nand UO_775 (O_775,N_24744,N_24865);
nand UO_776 (O_776,N_24638,N_24418);
and UO_777 (O_777,N_24627,N_24323);
or UO_778 (O_778,N_24723,N_24166);
xnor UO_779 (O_779,N_24452,N_24868);
nor UO_780 (O_780,N_24027,N_24498);
xnor UO_781 (O_781,N_24005,N_24470);
nor UO_782 (O_782,N_24598,N_24031);
nand UO_783 (O_783,N_24474,N_24858);
and UO_784 (O_784,N_24659,N_24315);
xor UO_785 (O_785,N_24034,N_24138);
and UO_786 (O_786,N_24703,N_24386);
nor UO_787 (O_787,N_24562,N_24831);
or UO_788 (O_788,N_24891,N_24331);
xor UO_789 (O_789,N_24826,N_24524);
nor UO_790 (O_790,N_24384,N_24175);
or UO_791 (O_791,N_24839,N_24266);
xnor UO_792 (O_792,N_24412,N_24111);
and UO_793 (O_793,N_24722,N_24820);
xor UO_794 (O_794,N_24769,N_24060);
nor UO_795 (O_795,N_24266,N_24621);
or UO_796 (O_796,N_24540,N_24065);
nand UO_797 (O_797,N_24540,N_24361);
xnor UO_798 (O_798,N_24906,N_24254);
xnor UO_799 (O_799,N_24344,N_24916);
nand UO_800 (O_800,N_24630,N_24107);
nand UO_801 (O_801,N_24884,N_24093);
nand UO_802 (O_802,N_24136,N_24144);
nand UO_803 (O_803,N_24988,N_24669);
xor UO_804 (O_804,N_24642,N_24966);
xor UO_805 (O_805,N_24176,N_24040);
nand UO_806 (O_806,N_24119,N_24317);
or UO_807 (O_807,N_24208,N_24071);
nor UO_808 (O_808,N_24232,N_24664);
nand UO_809 (O_809,N_24195,N_24965);
nand UO_810 (O_810,N_24582,N_24328);
and UO_811 (O_811,N_24738,N_24791);
and UO_812 (O_812,N_24877,N_24342);
nand UO_813 (O_813,N_24738,N_24390);
nor UO_814 (O_814,N_24107,N_24956);
and UO_815 (O_815,N_24015,N_24261);
and UO_816 (O_816,N_24200,N_24842);
and UO_817 (O_817,N_24854,N_24517);
nor UO_818 (O_818,N_24407,N_24425);
nand UO_819 (O_819,N_24664,N_24815);
xnor UO_820 (O_820,N_24202,N_24827);
xor UO_821 (O_821,N_24541,N_24598);
or UO_822 (O_822,N_24982,N_24751);
xnor UO_823 (O_823,N_24212,N_24600);
nor UO_824 (O_824,N_24704,N_24947);
xor UO_825 (O_825,N_24010,N_24708);
nor UO_826 (O_826,N_24292,N_24368);
or UO_827 (O_827,N_24080,N_24050);
xnor UO_828 (O_828,N_24977,N_24725);
and UO_829 (O_829,N_24829,N_24052);
and UO_830 (O_830,N_24242,N_24509);
and UO_831 (O_831,N_24362,N_24037);
or UO_832 (O_832,N_24806,N_24210);
nor UO_833 (O_833,N_24375,N_24577);
or UO_834 (O_834,N_24480,N_24100);
xor UO_835 (O_835,N_24016,N_24534);
nor UO_836 (O_836,N_24374,N_24671);
and UO_837 (O_837,N_24904,N_24581);
nand UO_838 (O_838,N_24598,N_24088);
nand UO_839 (O_839,N_24278,N_24032);
nand UO_840 (O_840,N_24457,N_24850);
nand UO_841 (O_841,N_24829,N_24995);
nand UO_842 (O_842,N_24915,N_24705);
or UO_843 (O_843,N_24576,N_24032);
xor UO_844 (O_844,N_24671,N_24568);
xnor UO_845 (O_845,N_24830,N_24603);
xnor UO_846 (O_846,N_24146,N_24429);
nand UO_847 (O_847,N_24911,N_24379);
xor UO_848 (O_848,N_24336,N_24068);
and UO_849 (O_849,N_24164,N_24421);
nor UO_850 (O_850,N_24597,N_24247);
nor UO_851 (O_851,N_24810,N_24735);
nor UO_852 (O_852,N_24417,N_24814);
xor UO_853 (O_853,N_24855,N_24498);
or UO_854 (O_854,N_24200,N_24199);
and UO_855 (O_855,N_24958,N_24366);
nand UO_856 (O_856,N_24186,N_24473);
xor UO_857 (O_857,N_24300,N_24816);
and UO_858 (O_858,N_24956,N_24472);
nor UO_859 (O_859,N_24545,N_24959);
nor UO_860 (O_860,N_24348,N_24337);
and UO_861 (O_861,N_24510,N_24680);
and UO_862 (O_862,N_24051,N_24826);
or UO_863 (O_863,N_24877,N_24814);
nor UO_864 (O_864,N_24102,N_24197);
nand UO_865 (O_865,N_24227,N_24806);
and UO_866 (O_866,N_24256,N_24929);
and UO_867 (O_867,N_24914,N_24311);
or UO_868 (O_868,N_24841,N_24334);
nor UO_869 (O_869,N_24026,N_24659);
nand UO_870 (O_870,N_24136,N_24718);
nand UO_871 (O_871,N_24050,N_24962);
and UO_872 (O_872,N_24386,N_24192);
xnor UO_873 (O_873,N_24945,N_24505);
or UO_874 (O_874,N_24250,N_24266);
or UO_875 (O_875,N_24801,N_24358);
nor UO_876 (O_876,N_24951,N_24333);
and UO_877 (O_877,N_24136,N_24431);
nand UO_878 (O_878,N_24415,N_24609);
nor UO_879 (O_879,N_24295,N_24620);
and UO_880 (O_880,N_24961,N_24620);
nor UO_881 (O_881,N_24816,N_24159);
nand UO_882 (O_882,N_24531,N_24795);
and UO_883 (O_883,N_24756,N_24651);
and UO_884 (O_884,N_24443,N_24099);
nand UO_885 (O_885,N_24148,N_24580);
nand UO_886 (O_886,N_24727,N_24348);
or UO_887 (O_887,N_24689,N_24867);
xor UO_888 (O_888,N_24806,N_24001);
xnor UO_889 (O_889,N_24487,N_24365);
nor UO_890 (O_890,N_24960,N_24077);
nor UO_891 (O_891,N_24089,N_24598);
nand UO_892 (O_892,N_24247,N_24492);
nand UO_893 (O_893,N_24498,N_24205);
and UO_894 (O_894,N_24885,N_24860);
nand UO_895 (O_895,N_24067,N_24573);
or UO_896 (O_896,N_24180,N_24247);
xnor UO_897 (O_897,N_24635,N_24146);
and UO_898 (O_898,N_24163,N_24473);
xor UO_899 (O_899,N_24513,N_24591);
or UO_900 (O_900,N_24759,N_24249);
nor UO_901 (O_901,N_24614,N_24146);
nand UO_902 (O_902,N_24346,N_24081);
and UO_903 (O_903,N_24494,N_24636);
nor UO_904 (O_904,N_24510,N_24505);
nor UO_905 (O_905,N_24056,N_24785);
nor UO_906 (O_906,N_24216,N_24844);
xnor UO_907 (O_907,N_24349,N_24253);
nor UO_908 (O_908,N_24544,N_24744);
nand UO_909 (O_909,N_24812,N_24360);
or UO_910 (O_910,N_24001,N_24917);
xnor UO_911 (O_911,N_24221,N_24823);
or UO_912 (O_912,N_24753,N_24223);
or UO_913 (O_913,N_24396,N_24917);
nor UO_914 (O_914,N_24501,N_24639);
xor UO_915 (O_915,N_24949,N_24745);
and UO_916 (O_916,N_24626,N_24652);
and UO_917 (O_917,N_24180,N_24382);
and UO_918 (O_918,N_24242,N_24092);
nor UO_919 (O_919,N_24890,N_24307);
xnor UO_920 (O_920,N_24059,N_24489);
xor UO_921 (O_921,N_24004,N_24591);
nor UO_922 (O_922,N_24209,N_24604);
or UO_923 (O_923,N_24462,N_24013);
nor UO_924 (O_924,N_24482,N_24737);
nor UO_925 (O_925,N_24687,N_24983);
nor UO_926 (O_926,N_24200,N_24765);
xnor UO_927 (O_927,N_24312,N_24910);
or UO_928 (O_928,N_24425,N_24967);
nand UO_929 (O_929,N_24006,N_24686);
nor UO_930 (O_930,N_24851,N_24507);
xnor UO_931 (O_931,N_24843,N_24741);
or UO_932 (O_932,N_24111,N_24046);
and UO_933 (O_933,N_24392,N_24747);
nor UO_934 (O_934,N_24408,N_24595);
nand UO_935 (O_935,N_24803,N_24380);
or UO_936 (O_936,N_24850,N_24739);
nor UO_937 (O_937,N_24952,N_24913);
nand UO_938 (O_938,N_24996,N_24156);
nor UO_939 (O_939,N_24998,N_24400);
xnor UO_940 (O_940,N_24827,N_24387);
nand UO_941 (O_941,N_24653,N_24488);
or UO_942 (O_942,N_24516,N_24450);
nand UO_943 (O_943,N_24508,N_24939);
nand UO_944 (O_944,N_24917,N_24299);
nor UO_945 (O_945,N_24151,N_24394);
and UO_946 (O_946,N_24037,N_24001);
nor UO_947 (O_947,N_24787,N_24486);
and UO_948 (O_948,N_24658,N_24933);
xor UO_949 (O_949,N_24151,N_24871);
or UO_950 (O_950,N_24301,N_24191);
nor UO_951 (O_951,N_24273,N_24050);
and UO_952 (O_952,N_24064,N_24993);
or UO_953 (O_953,N_24241,N_24523);
or UO_954 (O_954,N_24403,N_24407);
nor UO_955 (O_955,N_24136,N_24289);
xor UO_956 (O_956,N_24134,N_24688);
or UO_957 (O_957,N_24389,N_24179);
xnor UO_958 (O_958,N_24198,N_24497);
xor UO_959 (O_959,N_24996,N_24771);
and UO_960 (O_960,N_24604,N_24482);
and UO_961 (O_961,N_24951,N_24522);
nand UO_962 (O_962,N_24856,N_24352);
and UO_963 (O_963,N_24203,N_24371);
nand UO_964 (O_964,N_24739,N_24214);
or UO_965 (O_965,N_24618,N_24112);
and UO_966 (O_966,N_24792,N_24595);
nor UO_967 (O_967,N_24660,N_24539);
nand UO_968 (O_968,N_24970,N_24255);
or UO_969 (O_969,N_24692,N_24580);
nor UO_970 (O_970,N_24039,N_24111);
and UO_971 (O_971,N_24919,N_24050);
nor UO_972 (O_972,N_24480,N_24300);
and UO_973 (O_973,N_24992,N_24566);
and UO_974 (O_974,N_24959,N_24645);
and UO_975 (O_975,N_24871,N_24478);
nand UO_976 (O_976,N_24718,N_24441);
or UO_977 (O_977,N_24415,N_24534);
nand UO_978 (O_978,N_24986,N_24968);
nand UO_979 (O_979,N_24314,N_24265);
nor UO_980 (O_980,N_24432,N_24099);
xor UO_981 (O_981,N_24949,N_24723);
and UO_982 (O_982,N_24353,N_24675);
and UO_983 (O_983,N_24465,N_24537);
and UO_984 (O_984,N_24669,N_24217);
nand UO_985 (O_985,N_24180,N_24852);
xnor UO_986 (O_986,N_24641,N_24959);
and UO_987 (O_987,N_24447,N_24180);
nor UO_988 (O_988,N_24124,N_24607);
or UO_989 (O_989,N_24893,N_24892);
nand UO_990 (O_990,N_24632,N_24143);
and UO_991 (O_991,N_24203,N_24560);
xor UO_992 (O_992,N_24412,N_24791);
nor UO_993 (O_993,N_24643,N_24890);
nor UO_994 (O_994,N_24528,N_24747);
nor UO_995 (O_995,N_24531,N_24770);
xor UO_996 (O_996,N_24323,N_24379);
and UO_997 (O_997,N_24931,N_24554);
and UO_998 (O_998,N_24589,N_24261);
or UO_999 (O_999,N_24661,N_24550);
nand UO_1000 (O_1000,N_24856,N_24671);
and UO_1001 (O_1001,N_24215,N_24316);
nand UO_1002 (O_1002,N_24573,N_24220);
and UO_1003 (O_1003,N_24684,N_24916);
nor UO_1004 (O_1004,N_24311,N_24848);
nand UO_1005 (O_1005,N_24814,N_24087);
or UO_1006 (O_1006,N_24310,N_24542);
and UO_1007 (O_1007,N_24592,N_24778);
nor UO_1008 (O_1008,N_24674,N_24880);
nand UO_1009 (O_1009,N_24847,N_24036);
and UO_1010 (O_1010,N_24697,N_24090);
xnor UO_1011 (O_1011,N_24954,N_24427);
and UO_1012 (O_1012,N_24094,N_24966);
xnor UO_1013 (O_1013,N_24497,N_24558);
nor UO_1014 (O_1014,N_24716,N_24286);
or UO_1015 (O_1015,N_24823,N_24201);
nand UO_1016 (O_1016,N_24815,N_24504);
nor UO_1017 (O_1017,N_24935,N_24335);
nor UO_1018 (O_1018,N_24763,N_24192);
and UO_1019 (O_1019,N_24591,N_24823);
nand UO_1020 (O_1020,N_24449,N_24148);
nor UO_1021 (O_1021,N_24193,N_24871);
nand UO_1022 (O_1022,N_24556,N_24876);
or UO_1023 (O_1023,N_24754,N_24016);
and UO_1024 (O_1024,N_24422,N_24931);
or UO_1025 (O_1025,N_24096,N_24292);
nand UO_1026 (O_1026,N_24163,N_24095);
nand UO_1027 (O_1027,N_24138,N_24447);
and UO_1028 (O_1028,N_24539,N_24241);
and UO_1029 (O_1029,N_24244,N_24462);
and UO_1030 (O_1030,N_24318,N_24585);
nand UO_1031 (O_1031,N_24366,N_24989);
and UO_1032 (O_1032,N_24775,N_24125);
or UO_1033 (O_1033,N_24121,N_24403);
nand UO_1034 (O_1034,N_24244,N_24379);
or UO_1035 (O_1035,N_24718,N_24482);
xor UO_1036 (O_1036,N_24960,N_24542);
nor UO_1037 (O_1037,N_24603,N_24351);
xor UO_1038 (O_1038,N_24704,N_24439);
xor UO_1039 (O_1039,N_24570,N_24569);
and UO_1040 (O_1040,N_24912,N_24457);
nand UO_1041 (O_1041,N_24142,N_24081);
nand UO_1042 (O_1042,N_24084,N_24636);
and UO_1043 (O_1043,N_24015,N_24531);
or UO_1044 (O_1044,N_24435,N_24432);
nor UO_1045 (O_1045,N_24954,N_24797);
xnor UO_1046 (O_1046,N_24949,N_24781);
xnor UO_1047 (O_1047,N_24682,N_24382);
nand UO_1048 (O_1048,N_24577,N_24883);
nand UO_1049 (O_1049,N_24562,N_24447);
and UO_1050 (O_1050,N_24752,N_24457);
xor UO_1051 (O_1051,N_24331,N_24709);
xnor UO_1052 (O_1052,N_24524,N_24316);
or UO_1053 (O_1053,N_24526,N_24816);
and UO_1054 (O_1054,N_24668,N_24052);
xor UO_1055 (O_1055,N_24086,N_24406);
or UO_1056 (O_1056,N_24212,N_24442);
and UO_1057 (O_1057,N_24873,N_24697);
or UO_1058 (O_1058,N_24115,N_24343);
nand UO_1059 (O_1059,N_24794,N_24931);
nor UO_1060 (O_1060,N_24934,N_24647);
or UO_1061 (O_1061,N_24009,N_24302);
xnor UO_1062 (O_1062,N_24177,N_24782);
nor UO_1063 (O_1063,N_24631,N_24969);
xor UO_1064 (O_1064,N_24455,N_24246);
and UO_1065 (O_1065,N_24334,N_24457);
nor UO_1066 (O_1066,N_24845,N_24680);
and UO_1067 (O_1067,N_24609,N_24499);
xnor UO_1068 (O_1068,N_24784,N_24471);
nand UO_1069 (O_1069,N_24295,N_24502);
xor UO_1070 (O_1070,N_24142,N_24250);
nor UO_1071 (O_1071,N_24471,N_24849);
or UO_1072 (O_1072,N_24710,N_24369);
nand UO_1073 (O_1073,N_24563,N_24898);
and UO_1074 (O_1074,N_24203,N_24794);
nand UO_1075 (O_1075,N_24461,N_24249);
and UO_1076 (O_1076,N_24472,N_24920);
or UO_1077 (O_1077,N_24045,N_24522);
nor UO_1078 (O_1078,N_24003,N_24142);
or UO_1079 (O_1079,N_24724,N_24645);
nand UO_1080 (O_1080,N_24265,N_24129);
xnor UO_1081 (O_1081,N_24802,N_24567);
and UO_1082 (O_1082,N_24510,N_24846);
nand UO_1083 (O_1083,N_24279,N_24032);
nand UO_1084 (O_1084,N_24770,N_24284);
nor UO_1085 (O_1085,N_24142,N_24673);
nand UO_1086 (O_1086,N_24267,N_24386);
or UO_1087 (O_1087,N_24853,N_24336);
or UO_1088 (O_1088,N_24859,N_24508);
xnor UO_1089 (O_1089,N_24352,N_24676);
or UO_1090 (O_1090,N_24276,N_24205);
xor UO_1091 (O_1091,N_24914,N_24110);
xnor UO_1092 (O_1092,N_24313,N_24021);
and UO_1093 (O_1093,N_24234,N_24713);
or UO_1094 (O_1094,N_24746,N_24533);
nand UO_1095 (O_1095,N_24213,N_24322);
nand UO_1096 (O_1096,N_24050,N_24547);
and UO_1097 (O_1097,N_24363,N_24209);
or UO_1098 (O_1098,N_24368,N_24719);
xnor UO_1099 (O_1099,N_24546,N_24292);
nor UO_1100 (O_1100,N_24158,N_24130);
nor UO_1101 (O_1101,N_24815,N_24786);
xnor UO_1102 (O_1102,N_24808,N_24148);
nor UO_1103 (O_1103,N_24595,N_24027);
xnor UO_1104 (O_1104,N_24803,N_24982);
or UO_1105 (O_1105,N_24552,N_24342);
xnor UO_1106 (O_1106,N_24067,N_24209);
xnor UO_1107 (O_1107,N_24590,N_24301);
nor UO_1108 (O_1108,N_24524,N_24219);
xor UO_1109 (O_1109,N_24886,N_24976);
nor UO_1110 (O_1110,N_24009,N_24569);
and UO_1111 (O_1111,N_24338,N_24741);
nor UO_1112 (O_1112,N_24906,N_24191);
or UO_1113 (O_1113,N_24479,N_24460);
nand UO_1114 (O_1114,N_24690,N_24567);
and UO_1115 (O_1115,N_24511,N_24407);
nor UO_1116 (O_1116,N_24594,N_24610);
nor UO_1117 (O_1117,N_24493,N_24456);
xnor UO_1118 (O_1118,N_24539,N_24734);
nor UO_1119 (O_1119,N_24482,N_24887);
or UO_1120 (O_1120,N_24915,N_24092);
or UO_1121 (O_1121,N_24109,N_24658);
xnor UO_1122 (O_1122,N_24973,N_24058);
nor UO_1123 (O_1123,N_24452,N_24483);
or UO_1124 (O_1124,N_24253,N_24120);
xor UO_1125 (O_1125,N_24071,N_24920);
nand UO_1126 (O_1126,N_24161,N_24983);
nand UO_1127 (O_1127,N_24423,N_24005);
nand UO_1128 (O_1128,N_24774,N_24942);
and UO_1129 (O_1129,N_24876,N_24361);
nand UO_1130 (O_1130,N_24020,N_24288);
xor UO_1131 (O_1131,N_24912,N_24838);
nand UO_1132 (O_1132,N_24143,N_24269);
nand UO_1133 (O_1133,N_24139,N_24580);
xnor UO_1134 (O_1134,N_24062,N_24024);
xor UO_1135 (O_1135,N_24022,N_24793);
nor UO_1136 (O_1136,N_24975,N_24953);
nand UO_1137 (O_1137,N_24442,N_24720);
nor UO_1138 (O_1138,N_24349,N_24501);
xor UO_1139 (O_1139,N_24316,N_24251);
and UO_1140 (O_1140,N_24351,N_24975);
xnor UO_1141 (O_1141,N_24779,N_24340);
nor UO_1142 (O_1142,N_24714,N_24461);
xor UO_1143 (O_1143,N_24103,N_24186);
and UO_1144 (O_1144,N_24926,N_24444);
or UO_1145 (O_1145,N_24038,N_24363);
xnor UO_1146 (O_1146,N_24216,N_24897);
nand UO_1147 (O_1147,N_24774,N_24979);
nand UO_1148 (O_1148,N_24353,N_24678);
xor UO_1149 (O_1149,N_24282,N_24270);
and UO_1150 (O_1150,N_24574,N_24322);
nor UO_1151 (O_1151,N_24736,N_24596);
nor UO_1152 (O_1152,N_24173,N_24793);
xor UO_1153 (O_1153,N_24331,N_24062);
nand UO_1154 (O_1154,N_24794,N_24533);
or UO_1155 (O_1155,N_24435,N_24727);
nor UO_1156 (O_1156,N_24177,N_24174);
nor UO_1157 (O_1157,N_24291,N_24321);
nor UO_1158 (O_1158,N_24228,N_24982);
or UO_1159 (O_1159,N_24043,N_24364);
or UO_1160 (O_1160,N_24100,N_24963);
xnor UO_1161 (O_1161,N_24008,N_24243);
nor UO_1162 (O_1162,N_24682,N_24749);
and UO_1163 (O_1163,N_24728,N_24390);
nand UO_1164 (O_1164,N_24713,N_24989);
nand UO_1165 (O_1165,N_24430,N_24863);
or UO_1166 (O_1166,N_24409,N_24639);
nand UO_1167 (O_1167,N_24167,N_24720);
nor UO_1168 (O_1168,N_24908,N_24061);
and UO_1169 (O_1169,N_24945,N_24805);
nor UO_1170 (O_1170,N_24561,N_24867);
nor UO_1171 (O_1171,N_24045,N_24902);
xnor UO_1172 (O_1172,N_24373,N_24617);
nand UO_1173 (O_1173,N_24064,N_24774);
nand UO_1174 (O_1174,N_24322,N_24850);
xnor UO_1175 (O_1175,N_24010,N_24932);
or UO_1176 (O_1176,N_24458,N_24718);
xor UO_1177 (O_1177,N_24341,N_24695);
xor UO_1178 (O_1178,N_24664,N_24597);
or UO_1179 (O_1179,N_24391,N_24495);
and UO_1180 (O_1180,N_24466,N_24463);
or UO_1181 (O_1181,N_24411,N_24516);
nor UO_1182 (O_1182,N_24088,N_24013);
nand UO_1183 (O_1183,N_24066,N_24001);
xnor UO_1184 (O_1184,N_24181,N_24447);
xnor UO_1185 (O_1185,N_24625,N_24140);
nand UO_1186 (O_1186,N_24507,N_24700);
or UO_1187 (O_1187,N_24681,N_24941);
or UO_1188 (O_1188,N_24704,N_24235);
or UO_1189 (O_1189,N_24002,N_24318);
xor UO_1190 (O_1190,N_24343,N_24009);
nand UO_1191 (O_1191,N_24358,N_24731);
nand UO_1192 (O_1192,N_24528,N_24818);
nor UO_1193 (O_1193,N_24044,N_24167);
nor UO_1194 (O_1194,N_24327,N_24581);
and UO_1195 (O_1195,N_24937,N_24500);
nand UO_1196 (O_1196,N_24282,N_24188);
or UO_1197 (O_1197,N_24198,N_24863);
and UO_1198 (O_1198,N_24635,N_24401);
or UO_1199 (O_1199,N_24601,N_24556);
nand UO_1200 (O_1200,N_24075,N_24647);
or UO_1201 (O_1201,N_24644,N_24789);
and UO_1202 (O_1202,N_24340,N_24189);
nand UO_1203 (O_1203,N_24178,N_24917);
xnor UO_1204 (O_1204,N_24126,N_24034);
or UO_1205 (O_1205,N_24632,N_24933);
xor UO_1206 (O_1206,N_24687,N_24601);
or UO_1207 (O_1207,N_24201,N_24630);
and UO_1208 (O_1208,N_24794,N_24441);
nor UO_1209 (O_1209,N_24944,N_24555);
and UO_1210 (O_1210,N_24825,N_24990);
nor UO_1211 (O_1211,N_24206,N_24762);
xnor UO_1212 (O_1212,N_24088,N_24586);
nor UO_1213 (O_1213,N_24169,N_24179);
nand UO_1214 (O_1214,N_24105,N_24750);
xnor UO_1215 (O_1215,N_24858,N_24917);
xor UO_1216 (O_1216,N_24207,N_24310);
or UO_1217 (O_1217,N_24335,N_24373);
and UO_1218 (O_1218,N_24222,N_24798);
or UO_1219 (O_1219,N_24792,N_24250);
nand UO_1220 (O_1220,N_24312,N_24149);
nand UO_1221 (O_1221,N_24646,N_24053);
nor UO_1222 (O_1222,N_24039,N_24988);
or UO_1223 (O_1223,N_24913,N_24918);
xor UO_1224 (O_1224,N_24007,N_24417);
nor UO_1225 (O_1225,N_24387,N_24574);
or UO_1226 (O_1226,N_24913,N_24229);
xor UO_1227 (O_1227,N_24470,N_24963);
xnor UO_1228 (O_1228,N_24766,N_24189);
nor UO_1229 (O_1229,N_24128,N_24820);
xnor UO_1230 (O_1230,N_24552,N_24127);
nor UO_1231 (O_1231,N_24279,N_24788);
and UO_1232 (O_1232,N_24701,N_24198);
nand UO_1233 (O_1233,N_24332,N_24351);
nand UO_1234 (O_1234,N_24531,N_24592);
or UO_1235 (O_1235,N_24898,N_24596);
and UO_1236 (O_1236,N_24339,N_24206);
and UO_1237 (O_1237,N_24911,N_24693);
or UO_1238 (O_1238,N_24834,N_24172);
xor UO_1239 (O_1239,N_24735,N_24275);
xnor UO_1240 (O_1240,N_24770,N_24108);
or UO_1241 (O_1241,N_24715,N_24724);
or UO_1242 (O_1242,N_24621,N_24018);
nor UO_1243 (O_1243,N_24593,N_24481);
xor UO_1244 (O_1244,N_24762,N_24235);
or UO_1245 (O_1245,N_24181,N_24934);
nor UO_1246 (O_1246,N_24588,N_24677);
and UO_1247 (O_1247,N_24082,N_24403);
and UO_1248 (O_1248,N_24889,N_24359);
and UO_1249 (O_1249,N_24294,N_24393);
and UO_1250 (O_1250,N_24157,N_24771);
nand UO_1251 (O_1251,N_24229,N_24759);
or UO_1252 (O_1252,N_24546,N_24260);
nand UO_1253 (O_1253,N_24460,N_24677);
and UO_1254 (O_1254,N_24566,N_24311);
nand UO_1255 (O_1255,N_24930,N_24967);
nand UO_1256 (O_1256,N_24180,N_24464);
nand UO_1257 (O_1257,N_24806,N_24449);
nor UO_1258 (O_1258,N_24980,N_24017);
nor UO_1259 (O_1259,N_24718,N_24276);
xor UO_1260 (O_1260,N_24767,N_24547);
or UO_1261 (O_1261,N_24626,N_24123);
or UO_1262 (O_1262,N_24615,N_24061);
and UO_1263 (O_1263,N_24018,N_24581);
or UO_1264 (O_1264,N_24565,N_24526);
xnor UO_1265 (O_1265,N_24259,N_24891);
xor UO_1266 (O_1266,N_24173,N_24469);
or UO_1267 (O_1267,N_24227,N_24413);
or UO_1268 (O_1268,N_24306,N_24410);
nand UO_1269 (O_1269,N_24555,N_24880);
nor UO_1270 (O_1270,N_24392,N_24806);
nand UO_1271 (O_1271,N_24193,N_24406);
nand UO_1272 (O_1272,N_24542,N_24723);
nor UO_1273 (O_1273,N_24563,N_24603);
or UO_1274 (O_1274,N_24998,N_24631);
or UO_1275 (O_1275,N_24963,N_24438);
and UO_1276 (O_1276,N_24606,N_24725);
or UO_1277 (O_1277,N_24511,N_24496);
or UO_1278 (O_1278,N_24894,N_24881);
or UO_1279 (O_1279,N_24101,N_24473);
and UO_1280 (O_1280,N_24626,N_24262);
and UO_1281 (O_1281,N_24524,N_24754);
and UO_1282 (O_1282,N_24563,N_24275);
nand UO_1283 (O_1283,N_24307,N_24536);
nand UO_1284 (O_1284,N_24669,N_24126);
nor UO_1285 (O_1285,N_24155,N_24431);
nand UO_1286 (O_1286,N_24137,N_24366);
and UO_1287 (O_1287,N_24323,N_24653);
and UO_1288 (O_1288,N_24583,N_24129);
nor UO_1289 (O_1289,N_24333,N_24708);
or UO_1290 (O_1290,N_24609,N_24047);
nor UO_1291 (O_1291,N_24338,N_24714);
and UO_1292 (O_1292,N_24204,N_24723);
and UO_1293 (O_1293,N_24269,N_24287);
and UO_1294 (O_1294,N_24328,N_24609);
nand UO_1295 (O_1295,N_24397,N_24003);
nor UO_1296 (O_1296,N_24379,N_24448);
and UO_1297 (O_1297,N_24424,N_24556);
xnor UO_1298 (O_1298,N_24453,N_24018);
nand UO_1299 (O_1299,N_24231,N_24485);
and UO_1300 (O_1300,N_24084,N_24434);
or UO_1301 (O_1301,N_24936,N_24232);
xnor UO_1302 (O_1302,N_24136,N_24482);
nor UO_1303 (O_1303,N_24429,N_24299);
xnor UO_1304 (O_1304,N_24782,N_24543);
nand UO_1305 (O_1305,N_24863,N_24127);
nor UO_1306 (O_1306,N_24546,N_24806);
nand UO_1307 (O_1307,N_24636,N_24403);
nor UO_1308 (O_1308,N_24361,N_24539);
nand UO_1309 (O_1309,N_24637,N_24734);
nand UO_1310 (O_1310,N_24599,N_24836);
and UO_1311 (O_1311,N_24968,N_24935);
nor UO_1312 (O_1312,N_24012,N_24446);
nor UO_1313 (O_1313,N_24925,N_24244);
nor UO_1314 (O_1314,N_24335,N_24223);
xor UO_1315 (O_1315,N_24574,N_24952);
xnor UO_1316 (O_1316,N_24303,N_24847);
nand UO_1317 (O_1317,N_24180,N_24939);
xnor UO_1318 (O_1318,N_24219,N_24319);
nor UO_1319 (O_1319,N_24910,N_24077);
xnor UO_1320 (O_1320,N_24549,N_24878);
nand UO_1321 (O_1321,N_24391,N_24083);
xor UO_1322 (O_1322,N_24969,N_24884);
and UO_1323 (O_1323,N_24657,N_24950);
and UO_1324 (O_1324,N_24320,N_24863);
xnor UO_1325 (O_1325,N_24478,N_24681);
and UO_1326 (O_1326,N_24501,N_24916);
xnor UO_1327 (O_1327,N_24148,N_24137);
nand UO_1328 (O_1328,N_24838,N_24651);
nand UO_1329 (O_1329,N_24498,N_24937);
nand UO_1330 (O_1330,N_24627,N_24752);
nor UO_1331 (O_1331,N_24462,N_24200);
nand UO_1332 (O_1332,N_24374,N_24228);
nand UO_1333 (O_1333,N_24487,N_24739);
xor UO_1334 (O_1334,N_24100,N_24189);
and UO_1335 (O_1335,N_24427,N_24932);
nand UO_1336 (O_1336,N_24102,N_24329);
and UO_1337 (O_1337,N_24835,N_24201);
nor UO_1338 (O_1338,N_24779,N_24326);
nor UO_1339 (O_1339,N_24071,N_24165);
nor UO_1340 (O_1340,N_24953,N_24146);
nand UO_1341 (O_1341,N_24177,N_24233);
nand UO_1342 (O_1342,N_24100,N_24240);
xnor UO_1343 (O_1343,N_24931,N_24414);
or UO_1344 (O_1344,N_24531,N_24835);
and UO_1345 (O_1345,N_24478,N_24696);
and UO_1346 (O_1346,N_24374,N_24681);
nor UO_1347 (O_1347,N_24634,N_24826);
nand UO_1348 (O_1348,N_24429,N_24280);
or UO_1349 (O_1349,N_24513,N_24357);
nor UO_1350 (O_1350,N_24504,N_24313);
xor UO_1351 (O_1351,N_24186,N_24158);
nand UO_1352 (O_1352,N_24454,N_24975);
xnor UO_1353 (O_1353,N_24699,N_24655);
xnor UO_1354 (O_1354,N_24784,N_24499);
and UO_1355 (O_1355,N_24680,N_24740);
or UO_1356 (O_1356,N_24184,N_24227);
nand UO_1357 (O_1357,N_24863,N_24428);
xor UO_1358 (O_1358,N_24387,N_24195);
or UO_1359 (O_1359,N_24659,N_24943);
or UO_1360 (O_1360,N_24236,N_24474);
nor UO_1361 (O_1361,N_24756,N_24122);
nor UO_1362 (O_1362,N_24207,N_24937);
or UO_1363 (O_1363,N_24802,N_24902);
xnor UO_1364 (O_1364,N_24104,N_24740);
nor UO_1365 (O_1365,N_24719,N_24764);
nor UO_1366 (O_1366,N_24712,N_24704);
xnor UO_1367 (O_1367,N_24656,N_24022);
nor UO_1368 (O_1368,N_24288,N_24168);
nand UO_1369 (O_1369,N_24482,N_24944);
and UO_1370 (O_1370,N_24713,N_24885);
xor UO_1371 (O_1371,N_24556,N_24028);
xnor UO_1372 (O_1372,N_24472,N_24046);
and UO_1373 (O_1373,N_24039,N_24347);
and UO_1374 (O_1374,N_24913,N_24698);
and UO_1375 (O_1375,N_24177,N_24514);
xnor UO_1376 (O_1376,N_24415,N_24388);
or UO_1377 (O_1377,N_24235,N_24711);
and UO_1378 (O_1378,N_24404,N_24470);
and UO_1379 (O_1379,N_24196,N_24938);
or UO_1380 (O_1380,N_24337,N_24080);
or UO_1381 (O_1381,N_24714,N_24152);
xor UO_1382 (O_1382,N_24483,N_24267);
nand UO_1383 (O_1383,N_24883,N_24324);
xor UO_1384 (O_1384,N_24827,N_24548);
xor UO_1385 (O_1385,N_24353,N_24375);
nand UO_1386 (O_1386,N_24230,N_24037);
nor UO_1387 (O_1387,N_24814,N_24789);
nor UO_1388 (O_1388,N_24287,N_24848);
nand UO_1389 (O_1389,N_24517,N_24669);
nand UO_1390 (O_1390,N_24680,N_24362);
nand UO_1391 (O_1391,N_24364,N_24897);
nor UO_1392 (O_1392,N_24411,N_24656);
or UO_1393 (O_1393,N_24897,N_24291);
nor UO_1394 (O_1394,N_24180,N_24086);
nor UO_1395 (O_1395,N_24397,N_24500);
nand UO_1396 (O_1396,N_24010,N_24476);
nor UO_1397 (O_1397,N_24472,N_24819);
and UO_1398 (O_1398,N_24048,N_24574);
xnor UO_1399 (O_1399,N_24414,N_24820);
xnor UO_1400 (O_1400,N_24812,N_24550);
and UO_1401 (O_1401,N_24838,N_24292);
or UO_1402 (O_1402,N_24718,N_24772);
xor UO_1403 (O_1403,N_24284,N_24251);
xor UO_1404 (O_1404,N_24843,N_24895);
xor UO_1405 (O_1405,N_24503,N_24909);
or UO_1406 (O_1406,N_24475,N_24772);
xor UO_1407 (O_1407,N_24284,N_24920);
nor UO_1408 (O_1408,N_24164,N_24078);
xnor UO_1409 (O_1409,N_24158,N_24062);
or UO_1410 (O_1410,N_24368,N_24073);
nand UO_1411 (O_1411,N_24467,N_24545);
nand UO_1412 (O_1412,N_24677,N_24670);
or UO_1413 (O_1413,N_24731,N_24552);
xnor UO_1414 (O_1414,N_24281,N_24419);
nor UO_1415 (O_1415,N_24575,N_24353);
nor UO_1416 (O_1416,N_24984,N_24647);
and UO_1417 (O_1417,N_24922,N_24995);
nor UO_1418 (O_1418,N_24764,N_24511);
and UO_1419 (O_1419,N_24973,N_24373);
xnor UO_1420 (O_1420,N_24805,N_24714);
or UO_1421 (O_1421,N_24777,N_24037);
and UO_1422 (O_1422,N_24352,N_24123);
xor UO_1423 (O_1423,N_24406,N_24705);
and UO_1424 (O_1424,N_24910,N_24748);
nand UO_1425 (O_1425,N_24918,N_24267);
nand UO_1426 (O_1426,N_24356,N_24361);
or UO_1427 (O_1427,N_24761,N_24502);
nand UO_1428 (O_1428,N_24925,N_24612);
nor UO_1429 (O_1429,N_24188,N_24445);
and UO_1430 (O_1430,N_24151,N_24289);
and UO_1431 (O_1431,N_24602,N_24521);
and UO_1432 (O_1432,N_24318,N_24678);
nand UO_1433 (O_1433,N_24195,N_24781);
and UO_1434 (O_1434,N_24251,N_24240);
or UO_1435 (O_1435,N_24946,N_24753);
or UO_1436 (O_1436,N_24147,N_24020);
or UO_1437 (O_1437,N_24422,N_24109);
xor UO_1438 (O_1438,N_24237,N_24380);
nand UO_1439 (O_1439,N_24483,N_24771);
and UO_1440 (O_1440,N_24177,N_24348);
nand UO_1441 (O_1441,N_24035,N_24967);
xor UO_1442 (O_1442,N_24579,N_24334);
nand UO_1443 (O_1443,N_24900,N_24359);
or UO_1444 (O_1444,N_24737,N_24292);
or UO_1445 (O_1445,N_24951,N_24768);
or UO_1446 (O_1446,N_24465,N_24759);
and UO_1447 (O_1447,N_24885,N_24292);
nor UO_1448 (O_1448,N_24848,N_24879);
xnor UO_1449 (O_1449,N_24755,N_24900);
xnor UO_1450 (O_1450,N_24864,N_24055);
nor UO_1451 (O_1451,N_24860,N_24652);
nand UO_1452 (O_1452,N_24169,N_24819);
or UO_1453 (O_1453,N_24586,N_24535);
and UO_1454 (O_1454,N_24340,N_24918);
nor UO_1455 (O_1455,N_24092,N_24826);
nand UO_1456 (O_1456,N_24930,N_24409);
xor UO_1457 (O_1457,N_24479,N_24409);
nor UO_1458 (O_1458,N_24948,N_24987);
or UO_1459 (O_1459,N_24786,N_24063);
nand UO_1460 (O_1460,N_24762,N_24129);
or UO_1461 (O_1461,N_24557,N_24036);
xor UO_1462 (O_1462,N_24967,N_24802);
and UO_1463 (O_1463,N_24688,N_24174);
nand UO_1464 (O_1464,N_24275,N_24964);
or UO_1465 (O_1465,N_24132,N_24761);
and UO_1466 (O_1466,N_24435,N_24716);
and UO_1467 (O_1467,N_24789,N_24614);
and UO_1468 (O_1468,N_24905,N_24463);
or UO_1469 (O_1469,N_24426,N_24844);
xor UO_1470 (O_1470,N_24630,N_24189);
or UO_1471 (O_1471,N_24716,N_24091);
or UO_1472 (O_1472,N_24660,N_24635);
and UO_1473 (O_1473,N_24616,N_24309);
xnor UO_1474 (O_1474,N_24965,N_24011);
xnor UO_1475 (O_1475,N_24235,N_24791);
or UO_1476 (O_1476,N_24423,N_24064);
or UO_1477 (O_1477,N_24278,N_24791);
xor UO_1478 (O_1478,N_24441,N_24416);
and UO_1479 (O_1479,N_24295,N_24608);
and UO_1480 (O_1480,N_24180,N_24378);
nand UO_1481 (O_1481,N_24570,N_24262);
and UO_1482 (O_1482,N_24888,N_24873);
xnor UO_1483 (O_1483,N_24564,N_24057);
or UO_1484 (O_1484,N_24940,N_24422);
nand UO_1485 (O_1485,N_24753,N_24210);
xnor UO_1486 (O_1486,N_24059,N_24395);
or UO_1487 (O_1487,N_24115,N_24383);
nor UO_1488 (O_1488,N_24989,N_24932);
nor UO_1489 (O_1489,N_24770,N_24401);
nand UO_1490 (O_1490,N_24980,N_24715);
and UO_1491 (O_1491,N_24437,N_24608);
xor UO_1492 (O_1492,N_24463,N_24899);
nor UO_1493 (O_1493,N_24593,N_24602);
nand UO_1494 (O_1494,N_24094,N_24336);
and UO_1495 (O_1495,N_24775,N_24234);
nor UO_1496 (O_1496,N_24762,N_24220);
or UO_1497 (O_1497,N_24066,N_24045);
nor UO_1498 (O_1498,N_24494,N_24354);
or UO_1499 (O_1499,N_24662,N_24365);
and UO_1500 (O_1500,N_24563,N_24994);
or UO_1501 (O_1501,N_24775,N_24564);
nor UO_1502 (O_1502,N_24564,N_24760);
or UO_1503 (O_1503,N_24782,N_24771);
nor UO_1504 (O_1504,N_24046,N_24446);
or UO_1505 (O_1505,N_24478,N_24170);
xnor UO_1506 (O_1506,N_24411,N_24201);
xor UO_1507 (O_1507,N_24483,N_24182);
and UO_1508 (O_1508,N_24020,N_24596);
or UO_1509 (O_1509,N_24412,N_24848);
nand UO_1510 (O_1510,N_24222,N_24442);
and UO_1511 (O_1511,N_24271,N_24558);
nor UO_1512 (O_1512,N_24873,N_24220);
xnor UO_1513 (O_1513,N_24563,N_24614);
and UO_1514 (O_1514,N_24838,N_24081);
and UO_1515 (O_1515,N_24722,N_24996);
and UO_1516 (O_1516,N_24495,N_24254);
xor UO_1517 (O_1517,N_24896,N_24237);
nor UO_1518 (O_1518,N_24457,N_24840);
or UO_1519 (O_1519,N_24916,N_24601);
and UO_1520 (O_1520,N_24111,N_24038);
nand UO_1521 (O_1521,N_24474,N_24010);
nor UO_1522 (O_1522,N_24232,N_24388);
nand UO_1523 (O_1523,N_24824,N_24205);
and UO_1524 (O_1524,N_24808,N_24393);
or UO_1525 (O_1525,N_24023,N_24598);
xnor UO_1526 (O_1526,N_24965,N_24833);
and UO_1527 (O_1527,N_24328,N_24474);
nor UO_1528 (O_1528,N_24475,N_24043);
and UO_1529 (O_1529,N_24389,N_24986);
xor UO_1530 (O_1530,N_24021,N_24495);
nand UO_1531 (O_1531,N_24308,N_24499);
xor UO_1532 (O_1532,N_24022,N_24527);
xor UO_1533 (O_1533,N_24107,N_24256);
xnor UO_1534 (O_1534,N_24581,N_24876);
nand UO_1535 (O_1535,N_24564,N_24848);
and UO_1536 (O_1536,N_24369,N_24101);
or UO_1537 (O_1537,N_24790,N_24165);
nand UO_1538 (O_1538,N_24915,N_24153);
and UO_1539 (O_1539,N_24417,N_24552);
or UO_1540 (O_1540,N_24560,N_24723);
and UO_1541 (O_1541,N_24136,N_24841);
or UO_1542 (O_1542,N_24381,N_24661);
xnor UO_1543 (O_1543,N_24632,N_24670);
nor UO_1544 (O_1544,N_24385,N_24664);
nand UO_1545 (O_1545,N_24644,N_24373);
xor UO_1546 (O_1546,N_24236,N_24705);
and UO_1547 (O_1547,N_24812,N_24591);
xnor UO_1548 (O_1548,N_24952,N_24152);
xor UO_1549 (O_1549,N_24863,N_24130);
nand UO_1550 (O_1550,N_24503,N_24253);
nand UO_1551 (O_1551,N_24684,N_24509);
and UO_1552 (O_1552,N_24964,N_24073);
nor UO_1553 (O_1553,N_24145,N_24853);
nor UO_1554 (O_1554,N_24659,N_24886);
or UO_1555 (O_1555,N_24878,N_24437);
xnor UO_1556 (O_1556,N_24192,N_24523);
and UO_1557 (O_1557,N_24066,N_24666);
or UO_1558 (O_1558,N_24324,N_24905);
nor UO_1559 (O_1559,N_24476,N_24514);
nor UO_1560 (O_1560,N_24519,N_24457);
nor UO_1561 (O_1561,N_24650,N_24768);
nand UO_1562 (O_1562,N_24029,N_24569);
and UO_1563 (O_1563,N_24825,N_24592);
xnor UO_1564 (O_1564,N_24483,N_24472);
or UO_1565 (O_1565,N_24983,N_24193);
nand UO_1566 (O_1566,N_24526,N_24106);
xor UO_1567 (O_1567,N_24461,N_24363);
and UO_1568 (O_1568,N_24358,N_24441);
xnor UO_1569 (O_1569,N_24161,N_24658);
xnor UO_1570 (O_1570,N_24109,N_24808);
and UO_1571 (O_1571,N_24410,N_24738);
or UO_1572 (O_1572,N_24408,N_24315);
xnor UO_1573 (O_1573,N_24295,N_24634);
xor UO_1574 (O_1574,N_24796,N_24885);
and UO_1575 (O_1575,N_24525,N_24855);
nand UO_1576 (O_1576,N_24230,N_24797);
or UO_1577 (O_1577,N_24163,N_24956);
xor UO_1578 (O_1578,N_24407,N_24059);
xnor UO_1579 (O_1579,N_24449,N_24777);
nor UO_1580 (O_1580,N_24477,N_24518);
or UO_1581 (O_1581,N_24984,N_24410);
nor UO_1582 (O_1582,N_24555,N_24484);
nor UO_1583 (O_1583,N_24394,N_24769);
nor UO_1584 (O_1584,N_24051,N_24796);
and UO_1585 (O_1585,N_24410,N_24150);
nand UO_1586 (O_1586,N_24199,N_24311);
and UO_1587 (O_1587,N_24251,N_24455);
nor UO_1588 (O_1588,N_24054,N_24992);
nor UO_1589 (O_1589,N_24839,N_24794);
and UO_1590 (O_1590,N_24077,N_24847);
nor UO_1591 (O_1591,N_24926,N_24370);
nand UO_1592 (O_1592,N_24976,N_24300);
nand UO_1593 (O_1593,N_24410,N_24718);
nor UO_1594 (O_1594,N_24226,N_24378);
nand UO_1595 (O_1595,N_24738,N_24535);
and UO_1596 (O_1596,N_24859,N_24849);
and UO_1597 (O_1597,N_24673,N_24125);
and UO_1598 (O_1598,N_24945,N_24795);
nor UO_1599 (O_1599,N_24359,N_24057);
nor UO_1600 (O_1600,N_24055,N_24147);
xnor UO_1601 (O_1601,N_24443,N_24032);
nor UO_1602 (O_1602,N_24731,N_24637);
or UO_1603 (O_1603,N_24772,N_24031);
nor UO_1604 (O_1604,N_24976,N_24630);
xnor UO_1605 (O_1605,N_24452,N_24560);
nand UO_1606 (O_1606,N_24718,N_24825);
and UO_1607 (O_1607,N_24314,N_24106);
and UO_1608 (O_1608,N_24118,N_24928);
and UO_1609 (O_1609,N_24931,N_24413);
xor UO_1610 (O_1610,N_24049,N_24636);
and UO_1611 (O_1611,N_24100,N_24032);
xnor UO_1612 (O_1612,N_24775,N_24984);
and UO_1613 (O_1613,N_24135,N_24916);
xnor UO_1614 (O_1614,N_24293,N_24994);
nand UO_1615 (O_1615,N_24500,N_24141);
or UO_1616 (O_1616,N_24794,N_24974);
nor UO_1617 (O_1617,N_24722,N_24746);
and UO_1618 (O_1618,N_24814,N_24890);
and UO_1619 (O_1619,N_24343,N_24110);
nor UO_1620 (O_1620,N_24061,N_24437);
and UO_1621 (O_1621,N_24136,N_24960);
and UO_1622 (O_1622,N_24355,N_24319);
nand UO_1623 (O_1623,N_24898,N_24593);
nor UO_1624 (O_1624,N_24006,N_24698);
xor UO_1625 (O_1625,N_24275,N_24083);
nand UO_1626 (O_1626,N_24176,N_24591);
nand UO_1627 (O_1627,N_24584,N_24504);
nor UO_1628 (O_1628,N_24834,N_24950);
or UO_1629 (O_1629,N_24670,N_24995);
xnor UO_1630 (O_1630,N_24752,N_24450);
xor UO_1631 (O_1631,N_24301,N_24304);
and UO_1632 (O_1632,N_24586,N_24751);
and UO_1633 (O_1633,N_24400,N_24565);
nand UO_1634 (O_1634,N_24633,N_24867);
nand UO_1635 (O_1635,N_24196,N_24715);
xor UO_1636 (O_1636,N_24294,N_24422);
nor UO_1637 (O_1637,N_24861,N_24377);
nor UO_1638 (O_1638,N_24054,N_24124);
nor UO_1639 (O_1639,N_24750,N_24569);
nor UO_1640 (O_1640,N_24491,N_24498);
xor UO_1641 (O_1641,N_24777,N_24292);
and UO_1642 (O_1642,N_24516,N_24367);
or UO_1643 (O_1643,N_24261,N_24166);
or UO_1644 (O_1644,N_24534,N_24036);
or UO_1645 (O_1645,N_24605,N_24526);
xnor UO_1646 (O_1646,N_24892,N_24162);
nand UO_1647 (O_1647,N_24743,N_24270);
nand UO_1648 (O_1648,N_24387,N_24847);
nor UO_1649 (O_1649,N_24641,N_24507);
or UO_1650 (O_1650,N_24742,N_24662);
or UO_1651 (O_1651,N_24900,N_24109);
and UO_1652 (O_1652,N_24274,N_24061);
or UO_1653 (O_1653,N_24358,N_24686);
or UO_1654 (O_1654,N_24457,N_24748);
nand UO_1655 (O_1655,N_24080,N_24268);
and UO_1656 (O_1656,N_24933,N_24538);
nor UO_1657 (O_1657,N_24179,N_24606);
or UO_1658 (O_1658,N_24738,N_24796);
and UO_1659 (O_1659,N_24089,N_24669);
xor UO_1660 (O_1660,N_24786,N_24978);
nor UO_1661 (O_1661,N_24279,N_24331);
nor UO_1662 (O_1662,N_24735,N_24692);
nand UO_1663 (O_1663,N_24940,N_24485);
and UO_1664 (O_1664,N_24075,N_24555);
nand UO_1665 (O_1665,N_24523,N_24959);
xnor UO_1666 (O_1666,N_24112,N_24752);
nor UO_1667 (O_1667,N_24797,N_24011);
xor UO_1668 (O_1668,N_24049,N_24278);
nand UO_1669 (O_1669,N_24431,N_24075);
xor UO_1670 (O_1670,N_24256,N_24698);
and UO_1671 (O_1671,N_24353,N_24643);
and UO_1672 (O_1672,N_24389,N_24416);
and UO_1673 (O_1673,N_24138,N_24522);
or UO_1674 (O_1674,N_24250,N_24066);
and UO_1675 (O_1675,N_24110,N_24081);
nor UO_1676 (O_1676,N_24993,N_24466);
nor UO_1677 (O_1677,N_24162,N_24225);
xor UO_1678 (O_1678,N_24672,N_24469);
or UO_1679 (O_1679,N_24570,N_24441);
nand UO_1680 (O_1680,N_24835,N_24384);
xnor UO_1681 (O_1681,N_24903,N_24218);
nor UO_1682 (O_1682,N_24319,N_24954);
xor UO_1683 (O_1683,N_24180,N_24813);
and UO_1684 (O_1684,N_24858,N_24326);
nor UO_1685 (O_1685,N_24310,N_24070);
xnor UO_1686 (O_1686,N_24647,N_24339);
xnor UO_1687 (O_1687,N_24343,N_24338);
nand UO_1688 (O_1688,N_24318,N_24311);
nor UO_1689 (O_1689,N_24108,N_24431);
nor UO_1690 (O_1690,N_24359,N_24981);
xnor UO_1691 (O_1691,N_24544,N_24515);
or UO_1692 (O_1692,N_24786,N_24179);
nand UO_1693 (O_1693,N_24348,N_24643);
nand UO_1694 (O_1694,N_24555,N_24056);
and UO_1695 (O_1695,N_24168,N_24796);
and UO_1696 (O_1696,N_24267,N_24997);
or UO_1697 (O_1697,N_24845,N_24073);
nor UO_1698 (O_1698,N_24612,N_24026);
nor UO_1699 (O_1699,N_24928,N_24435);
xor UO_1700 (O_1700,N_24025,N_24575);
and UO_1701 (O_1701,N_24897,N_24137);
nand UO_1702 (O_1702,N_24079,N_24746);
and UO_1703 (O_1703,N_24956,N_24902);
nor UO_1704 (O_1704,N_24325,N_24713);
nand UO_1705 (O_1705,N_24865,N_24868);
and UO_1706 (O_1706,N_24572,N_24904);
and UO_1707 (O_1707,N_24584,N_24568);
nor UO_1708 (O_1708,N_24496,N_24217);
xnor UO_1709 (O_1709,N_24277,N_24489);
and UO_1710 (O_1710,N_24502,N_24042);
xor UO_1711 (O_1711,N_24692,N_24043);
and UO_1712 (O_1712,N_24964,N_24638);
nand UO_1713 (O_1713,N_24316,N_24967);
nand UO_1714 (O_1714,N_24238,N_24426);
or UO_1715 (O_1715,N_24788,N_24283);
or UO_1716 (O_1716,N_24531,N_24529);
xor UO_1717 (O_1717,N_24232,N_24178);
nand UO_1718 (O_1718,N_24713,N_24082);
xnor UO_1719 (O_1719,N_24583,N_24426);
and UO_1720 (O_1720,N_24715,N_24383);
xnor UO_1721 (O_1721,N_24338,N_24055);
nand UO_1722 (O_1722,N_24155,N_24745);
and UO_1723 (O_1723,N_24601,N_24259);
nor UO_1724 (O_1724,N_24195,N_24397);
and UO_1725 (O_1725,N_24023,N_24665);
or UO_1726 (O_1726,N_24085,N_24407);
nand UO_1727 (O_1727,N_24580,N_24672);
and UO_1728 (O_1728,N_24790,N_24807);
and UO_1729 (O_1729,N_24857,N_24153);
nand UO_1730 (O_1730,N_24917,N_24269);
nor UO_1731 (O_1731,N_24968,N_24031);
nand UO_1732 (O_1732,N_24346,N_24088);
and UO_1733 (O_1733,N_24111,N_24282);
nor UO_1734 (O_1734,N_24901,N_24799);
or UO_1735 (O_1735,N_24966,N_24020);
nand UO_1736 (O_1736,N_24164,N_24740);
or UO_1737 (O_1737,N_24611,N_24867);
or UO_1738 (O_1738,N_24774,N_24933);
and UO_1739 (O_1739,N_24563,N_24371);
or UO_1740 (O_1740,N_24345,N_24504);
or UO_1741 (O_1741,N_24010,N_24509);
and UO_1742 (O_1742,N_24854,N_24137);
or UO_1743 (O_1743,N_24755,N_24097);
nor UO_1744 (O_1744,N_24714,N_24755);
nor UO_1745 (O_1745,N_24421,N_24041);
and UO_1746 (O_1746,N_24442,N_24778);
and UO_1747 (O_1747,N_24993,N_24496);
and UO_1748 (O_1748,N_24290,N_24714);
and UO_1749 (O_1749,N_24886,N_24844);
or UO_1750 (O_1750,N_24229,N_24894);
nor UO_1751 (O_1751,N_24057,N_24897);
or UO_1752 (O_1752,N_24791,N_24523);
nor UO_1753 (O_1753,N_24924,N_24371);
nand UO_1754 (O_1754,N_24174,N_24462);
nand UO_1755 (O_1755,N_24720,N_24600);
nor UO_1756 (O_1756,N_24223,N_24829);
nor UO_1757 (O_1757,N_24882,N_24510);
or UO_1758 (O_1758,N_24252,N_24129);
xor UO_1759 (O_1759,N_24072,N_24715);
or UO_1760 (O_1760,N_24127,N_24564);
nand UO_1761 (O_1761,N_24457,N_24598);
nand UO_1762 (O_1762,N_24969,N_24214);
nand UO_1763 (O_1763,N_24186,N_24499);
nor UO_1764 (O_1764,N_24652,N_24737);
xnor UO_1765 (O_1765,N_24627,N_24507);
and UO_1766 (O_1766,N_24915,N_24367);
or UO_1767 (O_1767,N_24881,N_24795);
xnor UO_1768 (O_1768,N_24463,N_24957);
and UO_1769 (O_1769,N_24165,N_24119);
xor UO_1770 (O_1770,N_24366,N_24683);
nor UO_1771 (O_1771,N_24476,N_24778);
and UO_1772 (O_1772,N_24327,N_24376);
nand UO_1773 (O_1773,N_24735,N_24080);
nor UO_1774 (O_1774,N_24844,N_24320);
xor UO_1775 (O_1775,N_24683,N_24049);
nand UO_1776 (O_1776,N_24926,N_24837);
nor UO_1777 (O_1777,N_24096,N_24296);
or UO_1778 (O_1778,N_24096,N_24746);
nand UO_1779 (O_1779,N_24408,N_24743);
xor UO_1780 (O_1780,N_24493,N_24379);
and UO_1781 (O_1781,N_24863,N_24304);
nor UO_1782 (O_1782,N_24554,N_24986);
xnor UO_1783 (O_1783,N_24152,N_24536);
nand UO_1784 (O_1784,N_24618,N_24049);
nand UO_1785 (O_1785,N_24698,N_24775);
or UO_1786 (O_1786,N_24384,N_24121);
nor UO_1787 (O_1787,N_24171,N_24727);
nor UO_1788 (O_1788,N_24775,N_24290);
nor UO_1789 (O_1789,N_24388,N_24870);
nor UO_1790 (O_1790,N_24063,N_24851);
nor UO_1791 (O_1791,N_24221,N_24988);
nand UO_1792 (O_1792,N_24864,N_24467);
xor UO_1793 (O_1793,N_24667,N_24632);
or UO_1794 (O_1794,N_24057,N_24747);
and UO_1795 (O_1795,N_24747,N_24630);
nor UO_1796 (O_1796,N_24441,N_24880);
nor UO_1797 (O_1797,N_24031,N_24673);
and UO_1798 (O_1798,N_24824,N_24986);
and UO_1799 (O_1799,N_24103,N_24684);
nor UO_1800 (O_1800,N_24254,N_24719);
or UO_1801 (O_1801,N_24027,N_24460);
or UO_1802 (O_1802,N_24670,N_24386);
nand UO_1803 (O_1803,N_24612,N_24704);
and UO_1804 (O_1804,N_24896,N_24372);
xor UO_1805 (O_1805,N_24495,N_24692);
xnor UO_1806 (O_1806,N_24524,N_24843);
or UO_1807 (O_1807,N_24018,N_24855);
or UO_1808 (O_1808,N_24463,N_24603);
nand UO_1809 (O_1809,N_24305,N_24404);
and UO_1810 (O_1810,N_24878,N_24936);
and UO_1811 (O_1811,N_24158,N_24441);
or UO_1812 (O_1812,N_24788,N_24697);
nand UO_1813 (O_1813,N_24153,N_24591);
and UO_1814 (O_1814,N_24784,N_24814);
and UO_1815 (O_1815,N_24239,N_24571);
or UO_1816 (O_1816,N_24490,N_24888);
or UO_1817 (O_1817,N_24984,N_24522);
and UO_1818 (O_1818,N_24693,N_24758);
or UO_1819 (O_1819,N_24892,N_24982);
and UO_1820 (O_1820,N_24364,N_24827);
nand UO_1821 (O_1821,N_24517,N_24485);
and UO_1822 (O_1822,N_24456,N_24819);
xor UO_1823 (O_1823,N_24087,N_24709);
and UO_1824 (O_1824,N_24496,N_24875);
and UO_1825 (O_1825,N_24008,N_24310);
and UO_1826 (O_1826,N_24569,N_24298);
nor UO_1827 (O_1827,N_24809,N_24889);
nand UO_1828 (O_1828,N_24069,N_24931);
or UO_1829 (O_1829,N_24654,N_24198);
xnor UO_1830 (O_1830,N_24539,N_24166);
and UO_1831 (O_1831,N_24896,N_24239);
xor UO_1832 (O_1832,N_24231,N_24550);
and UO_1833 (O_1833,N_24322,N_24408);
nor UO_1834 (O_1834,N_24173,N_24763);
and UO_1835 (O_1835,N_24897,N_24692);
xor UO_1836 (O_1836,N_24472,N_24861);
nand UO_1837 (O_1837,N_24368,N_24251);
and UO_1838 (O_1838,N_24443,N_24472);
nand UO_1839 (O_1839,N_24658,N_24489);
xnor UO_1840 (O_1840,N_24239,N_24962);
and UO_1841 (O_1841,N_24334,N_24722);
and UO_1842 (O_1842,N_24050,N_24151);
nand UO_1843 (O_1843,N_24427,N_24436);
xnor UO_1844 (O_1844,N_24201,N_24922);
and UO_1845 (O_1845,N_24916,N_24160);
nand UO_1846 (O_1846,N_24231,N_24012);
xor UO_1847 (O_1847,N_24204,N_24415);
nand UO_1848 (O_1848,N_24335,N_24317);
nor UO_1849 (O_1849,N_24781,N_24197);
or UO_1850 (O_1850,N_24456,N_24644);
xnor UO_1851 (O_1851,N_24975,N_24469);
and UO_1852 (O_1852,N_24417,N_24435);
nand UO_1853 (O_1853,N_24849,N_24421);
nor UO_1854 (O_1854,N_24150,N_24242);
nor UO_1855 (O_1855,N_24679,N_24471);
xnor UO_1856 (O_1856,N_24097,N_24695);
nor UO_1857 (O_1857,N_24194,N_24163);
nand UO_1858 (O_1858,N_24982,N_24786);
xor UO_1859 (O_1859,N_24975,N_24233);
or UO_1860 (O_1860,N_24493,N_24220);
xnor UO_1861 (O_1861,N_24441,N_24410);
nand UO_1862 (O_1862,N_24635,N_24550);
xor UO_1863 (O_1863,N_24788,N_24382);
nand UO_1864 (O_1864,N_24708,N_24047);
or UO_1865 (O_1865,N_24427,N_24762);
nand UO_1866 (O_1866,N_24495,N_24917);
or UO_1867 (O_1867,N_24864,N_24166);
nor UO_1868 (O_1868,N_24294,N_24129);
xnor UO_1869 (O_1869,N_24004,N_24075);
nand UO_1870 (O_1870,N_24207,N_24788);
nand UO_1871 (O_1871,N_24701,N_24523);
nand UO_1872 (O_1872,N_24584,N_24250);
and UO_1873 (O_1873,N_24410,N_24836);
xnor UO_1874 (O_1874,N_24941,N_24015);
nor UO_1875 (O_1875,N_24996,N_24484);
nor UO_1876 (O_1876,N_24932,N_24715);
and UO_1877 (O_1877,N_24974,N_24676);
xnor UO_1878 (O_1878,N_24500,N_24571);
and UO_1879 (O_1879,N_24951,N_24529);
and UO_1880 (O_1880,N_24883,N_24540);
xor UO_1881 (O_1881,N_24036,N_24406);
and UO_1882 (O_1882,N_24528,N_24738);
or UO_1883 (O_1883,N_24785,N_24303);
xnor UO_1884 (O_1884,N_24550,N_24072);
and UO_1885 (O_1885,N_24130,N_24013);
nor UO_1886 (O_1886,N_24417,N_24125);
xor UO_1887 (O_1887,N_24038,N_24410);
or UO_1888 (O_1888,N_24574,N_24501);
and UO_1889 (O_1889,N_24252,N_24168);
or UO_1890 (O_1890,N_24717,N_24635);
or UO_1891 (O_1891,N_24399,N_24329);
nor UO_1892 (O_1892,N_24446,N_24853);
or UO_1893 (O_1893,N_24922,N_24958);
nand UO_1894 (O_1894,N_24327,N_24203);
nor UO_1895 (O_1895,N_24033,N_24462);
or UO_1896 (O_1896,N_24080,N_24366);
or UO_1897 (O_1897,N_24700,N_24875);
nor UO_1898 (O_1898,N_24067,N_24975);
xor UO_1899 (O_1899,N_24747,N_24809);
and UO_1900 (O_1900,N_24572,N_24619);
or UO_1901 (O_1901,N_24083,N_24858);
nand UO_1902 (O_1902,N_24081,N_24187);
or UO_1903 (O_1903,N_24145,N_24786);
and UO_1904 (O_1904,N_24737,N_24511);
nor UO_1905 (O_1905,N_24949,N_24529);
xnor UO_1906 (O_1906,N_24864,N_24057);
and UO_1907 (O_1907,N_24350,N_24834);
and UO_1908 (O_1908,N_24838,N_24719);
nand UO_1909 (O_1909,N_24368,N_24933);
nand UO_1910 (O_1910,N_24965,N_24670);
nand UO_1911 (O_1911,N_24637,N_24169);
or UO_1912 (O_1912,N_24353,N_24890);
or UO_1913 (O_1913,N_24142,N_24030);
and UO_1914 (O_1914,N_24416,N_24374);
and UO_1915 (O_1915,N_24545,N_24838);
nand UO_1916 (O_1916,N_24110,N_24934);
xnor UO_1917 (O_1917,N_24534,N_24900);
nor UO_1918 (O_1918,N_24691,N_24410);
nor UO_1919 (O_1919,N_24738,N_24803);
nand UO_1920 (O_1920,N_24432,N_24373);
or UO_1921 (O_1921,N_24527,N_24054);
or UO_1922 (O_1922,N_24124,N_24668);
nor UO_1923 (O_1923,N_24905,N_24161);
and UO_1924 (O_1924,N_24796,N_24960);
nand UO_1925 (O_1925,N_24400,N_24526);
xor UO_1926 (O_1926,N_24047,N_24137);
and UO_1927 (O_1927,N_24984,N_24686);
nor UO_1928 (O_1928,N_24693,N_24215);
or UO_1929 (O_1929,N_24450,N_24724);
and UO_1930 (O_1930,N_24253,N_24800);
nor UO_1931 (O_1931,N_24854,N_24589);
or UO_1932 (O_1932,N_24675,N_24602);
nand UO_1933 (O_1933,N_24384,N_24723);
xnor UO_1934 (O_1934,N_24466,N_24606);
or UO_1935 (O_1935,N_24032,N_24014);
nor UO_1936 (O_1936,N_24668,N_24654);
nand UO_1937 (O_1937,N_24583,N_24739);
nand UO_1938 (O_1938,N_24389,N_24976);
or UO_1939 (O_1939,N_24632,N_24756);
nand UO_1940 (O_1940,N_24227,N_24147);
or UO_1941 (O_1941,N_24195,N_24183);
nor UO_1942 (O_1942,N_24372,N_24755);
xor UO_1943 (O_1943,N_24748,N_24877);
or UO_1944 (O_1944,N_24599,N_24879);
and UO_1945 (O_1945,N_24553,N_24590);
xnor UO_1946 (O_1946,N_24609,N_24654);
and UO_1947 (O_1947,N_24851,N_24377);
nor UO_1948 (O_1948,N_24734,N_24017);
and UO_1949 (O_1949,N_24661,N_24163);
xnor UO_1950 (O_1950,N_24212,N_24040);
xor UO_1951 (O_1951,N_24468,N_24633);
or UO_1952 (O_1952,N_24498,N_24677);
nor UO_1953 (O_1953,N_24801,N_24290);
nor UO_1954 (O_1954,N_24820,N_24014);
and UO_1955 (O_1955,N_24416,N_24777);
and UO_1956 (O_1956,N_24499,N_24846);
nor UO_1957 (O_1957,N_24741,N_24910);
nor UO_1958 (O_1958,N_24426,N_24382);
nor UO_1959 (O_1959,N_24436,N_24349);
and UO_1960 (O_1960,N_24186,N_24744);
nor UO_1961 (O_1961,N_24254,N_24139);
nand UO_1962 (O_1962,N_24444,N_24424);
nand UO_1963 (O_1963,N_24200,N_24221);
nor UO_1964 (O_1964,N_24235,N_24860);
nand UO_1965 (O_1965,N_24773,N_24946);
or UO_1966 (O_1966,N_24400,N_24323);
and UO_1967 (O_1967,N_24116,N_24640);
and UO_1968 (O_1968,N_24236,N_24348);
nand UO_1969 (O_1969,N_24607,N_24867);
nor UO_1970 (O_1970,N_24483,N_24475);
and UO_1971 (O_1971,N_24071,N_24100);
nand UO_1972 (O_1972,N_24954,N_24946);
xor UO_1973 (O_1973,N_24470,N_24788);
nor UO_1974 (O_1974,N_24563,N_24754);
xnor UO_1975 (O_1975,N_24208,N_24284);
nand UO_1976 (O_1976,N_24272,N_24618);
nand UO_1977 (O_1977,N_24988,N_24859);
nand UO_1978 (O_1978,N_24982,N_24040);
xor UO_1979 (O_1979,N_24966,N_24229);
or UO_1980 (O_1980,N_24483,N_24101);
or UO_1981 (O_1981,N_24195,N_24898);
nand UO_1982 (O_1982,N_24363,N_24241);
nand UO_1983 (O_1983,N_24756,N_24236);
and UO_1984 (O_1984,N_24237,N_24089);
or UO_1985 (O_1985,N_24897,N_24488);
nand UO_1986 (O_1986,N_24710,N_24116);
and UO_1987 (O_1987,N_24048,N_24056);
nand UO_1988 (O_1988,N_24338,N_24307);
and UO_1989 (O_1989,N_24003,N_24365);
nand UO_1990 (O_1990,N_24770,N_24339);
nor UO_1991 (O_1991,N_24051,N_24032);
or UO_1992 (O_1992,N_24413,N_24876);
xnor UO_1993 (O_1993,N_24727,N_24316);
nor UO_1994 (O_1994,N_24132,N_24854);
nor UO_1995 (O_1995,N_24515,N_24563);
nor UO_1996 (O_1996,N_24219,N_24588);
or UO_1997 (O_1997,N_24930,N_24400);
nand UO_1998 (O_1998,N_24812,N_24668);
nand UO_1999 (O_1999,N_24132,N_24407);
xnor UO_2000 (O_2000,N_24426,N_24949);
nand UO_2001 (O_2001,N_24448,N_24651);
and UO_2002 (O_2002,N_24722,N_24455);
xor UO_2003 (O_2003,N_24509,N_24735);
and UO_2004 (O_2004,N_24365,N_24912);
nand UO_2005 (O_2005,N_24652,N_24578);
and UO_2006 (O_2006,N_24181,N_24507);
or UO_2007 (O_2007,N_24035,N_24267);
and UO_2008 (O_2008,N_24281,N_24348);
or UO_2009 (O_2009,N_24236,N_24063);
and UO_2010 (O_2010,N_24414,N_24040);
nor UO_2011 (O_2011,N_24625,N_24337);
nand UO_2012 (O_2012,N_24300,N_24597);
xor UO_2013 (O_2013,N_24105,N_24352);
xor UO_2014 (O_2014,N_24040,N_24236);
and UO_2015 (O_2015,N_24821,N_24858);
xnor UO_2016 (O_2016,N_24492,N_24239);
or UO_2017 (O_2017,N_24255,N_24554);
or UO_2018 (O_2018,N_24357,N_24319);
xnor UO_2019 (O_2019,N_24948,N_24575);
and UO_2020 (O_2020,N_24838,N_24939);
and UO_2021 (O_2021,N_24033,N_24954);
nand UO_2022 (O_2022,N_24228,N_24955);
xor UO_2023 (O_2023,N_24964,N_24586);
nand UO_2024 (O_2024,N_24150,N_24101);
nor UO_2025 (O_2025,N_24357,N_24312);
xnor UO_2026 (O_2026,N_24447,N_24607);
and UO_2027 (O_2027,N_24425,N_24140);
or UO_2028 (O_2028,N_24742,N_24384);
nand UO_2029 (O_2029,N_24665,N_24395);
or UO_2030 (O_2030,N_24573,N_24560);
nor UO_2031 (O_2031,N_24615,N_24561);
nand UO_2032 (O_2032,N_24176,N_24239);
and UO_2033 (O_2033,N_24889,N_24077);
and UO_2034 (O_2034,N_24283,N_24063);
and UO_2035 (O_2035,N_24758,N_24822);
and UO_2036 (O_2036,N_24910,N_24564);
xor UO_2037 (O_2037,N_24576,N_24539);
or UO_2038 (O_2038,N_24869,N_24615);
nand UO_2039 (O_2039,N_24850,N_24714);
xnor UO_2040 (O_2040,N_24008,N_24471);
or UO_2041 (O_2041,N_24700,N_24482);
nand UO_2042 (O_2042,N_24803,N_24927);
nand UO_2043 (O_2043,N_24973,N_24846);
nand UO_2044 (O_2044,N_24286,N_24755);
nand UO_2045 (O_2045,N_24790,N_24357);
xor UO_2046 (O_2046,N_24586,N_24844);
nand UO_2047 (O_2047,N_24387,N_24784);
or UO_2048 (O_2048,N_24215,N_24988);
and UO_2049 (O_2049,N_24210,N_24848);
xor UO_2050 (O_2050,N_24347,N_24131);
and UO_2051 (O_2051,N_24066,N_24221);
nor UO_2052 (O_2052,N_24196,N_24799);
xnor UO_2053 (O_2053,N_24169,N_24103);
or UO_2054 (O_2054,N_24949,N_24307);
xor UO_2055 (O_2055,N_24388,N_24469);
nor UO_2056 (O_2056,N_24590,N_24045);
and UO_2057 (O_2057,N_24317,N_24807);
xor UO_2058 (O_2058,N_24595,N_24002);
and UO_2059 (O_2059,N_24751,N_24879);
nor UO_2060 (O_2060,N_24615,N_24851);
xnor UO_2061 (O_2061,N_24976,N_24182);
nor UO_2062 (O_2062,N_24290,N_24194);
xnor UO_2063 (O_2063,N_24923,N_24390);
xnor UO_2064 (O_2064,N_24655,N_24788);
or UO_2065 (O_2065,N_24457,N_24286);
nor UO_2066 (O_2066,N_24895,N_24432);
or UO_2067 (O_2067,N_24034,N_24252);
or UO_2068 (O_2068,N_24346,N_24825);
nand UO_2069 (O_2069,N_24121,N_24842);
and UO_2070 (O_2070,N_24103,N_24100);
and UO_2071 (O_2071,N_24867,N_24969);
or UO_2072 (O_2072,N_24827,N_24309);
nand UO_2073 (O_2073,N_24793,N_24672);
nand UO_2074 (O_2074,N_24537,N_24975);
and UO_2075 (O_2075,N_24787,N_24087);
and UO_2076 (O_2076,N_24561,N_24633);
nor UO_2077 (O_2077,N_24910,N_24066);
or UO_2078 (O_2078,N_24209,N_24502);
xor UO_2079 (O_2079,N_24537,N_24016);
xnor UO_2080 (O_2080,N_24212,N_24572);
nor UO_2081 (O_2081,N_24392,N_24677);
and UO_2082 (O_2082,N_24418,N_24882);
nand UO_2083 (O_2083,N_24497,N_24679);
nand UO_2084 (O_2084,N_24220,N_24814);
and UO_2085 (O_2085,N_24671,N_24960);
and UO_2086 (O_2086,N_24653,N_24925);
nor UO_2087 (O_2087,N_24131,N_24326);
or UO_2088 (O_2088,N_24827,N_24112);
or UO_2089 (O_2089,N_24644,N_24118);
nand UO_2090 (O_2090,N_24474,N_24399);
nor UO_2091 (O_2091,N_24201,N_24396);
or UO_2092 (O_2092,N_24005,N_24002);
nor UO_2093 (O_2093,N_24924,N_24419);
nor UO_2094 (O_2094,N_24292,N_24840);
xnor UO_2095 (O_2095,N_24142,N_24838);
nand UO_2096 (O_2096,N_24381,N_24832);
and UO_2097 (O_2097,N_24740,N_24271);
xnor UO_2098 (O_2098,N_24982,N_24724);
xnor UO_2099 (O_2099,N_24392,N_24812);
or UO_2100 (O_2100,N_24979,N_24270);
or UO_2101 (O_2101,N_24791,N_24483);
or UO_2102 (O_2102,N_24175,N_24507);
and UO_2103 (O_2103,N_24836,N_24788);
nor UO_2104 (O_2104,N_24725,N_24337);
xnor UO_2105 (O_2105,N_24803,N_24525);
nor UO_2106 (O_2106,N_24898,N_24603);
or UO_2107 (O_2107,N_24719,N_24015);
nor UO_2108 (O_2108,N_24626,N_24111);
nor UO_2109 (O_2109,N_24013,N_24775);
nand UO_2110 (O_2110,N_24955,N_24512);
xnor UO_2111 (O_2111,N_24348,N_24289);
xnor UO_2112 (O_2112,N_24651,N_24940);
nand UO_2113 (O_2113,N_24277,N_24552);
xor UO_2114 (O_2114,N_24553,N_24656);
nand UO_2115 (O_2115,N_24464,N_24812);
and UO_2116 (O_2116,N_24768,N_24550);
xnor UO_2117 (O_2117,N_24368,N_24988);
or UO_2118 (O_2118,N_24720,N_24981);
or UO_2119 (O_2119,N_24486,N_24294);
xor UO_2120 (O_2120,N_24877,N_24409);
xnor UO_2121 (O_2121,N_24369,N_24978);
and UO_2122 (O_2122,N_24765,N_24364);
nand UO_2123 (O_2123,N_24184,N_24012);
or UO_2124 (O_2124,N_24895,N_24242);
and UO_2125 (O_2125,N_24191,N_24663);
or UO_2126 (O_2126,N_24303,N_24146);
or UO_2127 (O_2127,N_24094,N_24406);
nand UO_2128 (O_2128,N_24367,N_24882);
xor UO_2129 (O_2129,N_24273,N_24903);
nand UO_2130 (O_2130,N_24450,N_24472);
xor UO_2131 (O_2131,N_24762,N_24187);
or UO_2132 (O_2132,N_24651,N_24036);
nor UO_2133 (O_2133,N_24102,N_24001);
nor UO_2134 (O_2134,N_24017,N_24503);
and UO_2135 (O_2135,N_24643,N_24999);
nand UO_2136 (O_2136,N_24490,N_24500);
or UO_2137 (O_2137,N_24090,N_24989);
nor UO_2138 (O_2138,N_24456,N_24766);
nand UO_2139 (O_2139,N_24873,N_24826);
nor UO_2140 (O_2140,N_24038,N_24664);
nand UO_2141 (O_2141,N_24938,N_24936);
nand UO_2142 (O_2142,N_24633,N_24337);
nand UO_2143 (O_2143,N_24042,N_24579);
or UO_2144 (O_2144,N_24639,N_24095);
nand UO_2145 (O_2145,N_24773,N_24736);
and UO_2146 (O_2146,N_24663,N_24694);
and UO_2147 (O_2147,N_24267,N_24498);
nand UO_2148 (O_2148,N_24269,N_24648);
xnor UO_2149 (O_2149,N_24510,N_24614);
xor UO_2150 (O_2150,N_24644,N_24211);
nand UO_2151 (O_2151,N_24033,N_24877);
xnor UO_2152 (O_2152,N_24841,N_24678);
nand UO_2153 (O_2153,N_24797,N_24081);
nand UO_2154 (O_2154,N_24085,N_24143);
nand UO_2155 (O_2155,N_24825,N_24616);
and UO_2156 (O_2156,N_24277,N_24276);
xnor UO_2157 (O_2157,N_24310,N_24013);
nor UO_2158 (O_2158,N_24694,N_24757);
and UO_2159 (O_2159,N_24996,N_24678);
nand UO_2160 (O_2160,N_24114,N_24578);
xnor UO_2161 (O_2161,N_24675,N_24664);
xnor UO_2162 (O_2162,N_24788,N_24271);
xor UO_2163 (O_2163,N_24300,N_24395);
xnor UO_2164 (O_2164,N_24069,N_24247);
or UO_2165 (O_2165,N_24830,N_24223);
nand UO_2166 (O_2166,N_24140,N_24212);
and UO_2167 (O_2167,N_24605,N_24676);
and UO_2168 (O_2168,N_24653,N_24388);
nand UO_2169 (O_2169,N_24736,N_24549);
nor UO_2170 (O_2170,N_24192,N_24068);
nor UO_2171 (O_2171,N_24149,N_24290);
nand UO_2172 (O_2172,N_24883,N_24762);
nor UO_2173 (O_2173,N_24311,N_24406);
and UO_2174 (O_2174,N_24577,N_24247);
or UO_2175 (O_2175,N_24624,N_24861);
nand UO_2176 (O_2176,N_24169,N_24739);
or UO_2177 (O_2177,N_24231,N_24828);
nor UO_2178 (O_2178,N_24143,N_24188);
xor UO_2179 (O_2179,N_24765,N_24646);
or UO_2180 (O_2180,N_24601,N_24758);
and UO_2181 (O_2181,N_24408,N_24794);
and UO_2182 (O_2182,N_24096,N_24375);
nor UO_2183 (O_2183,N_24758,N_24623);
xor UO_2184 (O_2184,N_24687,N_24102);
or UO_2185 (O_2185,N_24515,N_24457);
nand UO_2186 (O_2186,N_24648,N_24563);
and UO_2187 (O_2187,N_24719,N_24341);
and UO_2188 (O_2188,N_24326,N_24666);
nor UO_2189 (O_2189,N_24420,N_24522);
nand UO_2190 (O_2190,N_24785,N_24675);
or UO_2191 (O_2191,N_24272,N_24626);
xor UO_2192 (O_2192,N_24301,N_24710);
nand UO_2193 (O_2193,N_24238,N_24604);
or UO_2194 (O_2194,N_24178,N_24756);
or UO_2195 (O_2195,N_24220,N_24933);
nand UO_2196 (O_2196,N_24135,N_24386);
nand UO_2197 (O_2197,N_24020,N_24999);
or UO_2198 (O_2198,N_24941,N_24290);
nand UO_2199 (O_2199,N_24216,N_24525);
or UO_2200 (O_2200,N_24520,N_24175);
xor UO_2201 (O_2201,N_24898,N_24064);
or UO_2202 (O_2202,N_24666,N_24909);
or UO_2203 (O_2203,N_24357,N_24457);
xor UO_2204 (O_2204,N_24742,N_24599);
nand UO_2205 (O_2205,N_24441,N_24090);
nand UO_2206 (O_2206,N_24974,N_24108);
nor UO_2207 (O_2207,N_24397,N_24794);
xnor UO_2208 (O_2208,N_24936,N_24828);
nand UO_2209 (O_2209,N_24659,N_24282);
xor UO_2210 (O_2210,N_24060,N_24696);
and UO_2211 (O_2211,N_24773,N_24913);
xnor UO_2212 (O_2212,N_24916,N_24491);
nand UO_2213 (O_2213,N_24038,N_24858);
or UO_2214 (O_2214,N_24652,N_24666);
or UO_2215 (O_2215,N_24501,N_24667);
and UO_2216 (O_2216,N_24526,N_24607);
nor UO_2217 (O_2217,N_24718,N_24665);
nand UO_2218 (O_2218,N_24312,N_24120);
nand UO_2219 (O_2219,N_24247,N_24176);
xor UO_2220 (O_2220,N_24020,N_24649);
nor UO_2221 (O_2221,N_24717,N_24332);
or UO_2222 (O_2222,N_24567,N_24835);
and UO_2223 (O_2223,N_24179,N_24063);
xnor UO_2224 (O_2224,N_24470,N_24502);
nand UO_2225 (O_2225,N_24013,N_24401);
and UO_2226 (O_2226,N_24314,N_24139);
xnor UO_2227 (O_2227,N_24211,N_24587);
nand UO_2228 (O_2228,N_24798,N_24302);
nand UO_2229 (O_2229,N_24652,N_24994);
nor UO_2230 (O_2230,N_24002,N_24854);
nand UO_2231 (O_2231,N_24171,N_24183);
xnor UO_2232 (O_2232,N_24706,N_24786);
and UO_2233 (O_2233,N_24858,N_24426);
nor UO_2234 (O_2234,N_24682,N_24528);
nor UO_2235 (O_2235,N_24347,N_24566);
or UO_2236 (O_2236,N_24640,N_24533);
or UO_2237 (O_2237,N_24142,N_24718);
nor UO_2238 (O_2238,N_24035,N_24620);
xnor UO_2239 (O_2239,N_24489,N_24330);
and UO_2240 (O_2240,N_24110,N_24553);
nand UO_2241 (O_2241,N_24444,N_24209);
xor UO_2242 (O_2242,N_24779,N_24160);
nand UO_2243 (O_2243,N_24627,N_24958);
nor UO_2244 (O_2244,N_24170,N_24555);
xnor UO_2245 (O_2245,N_24255,N_24862);
or UO_2246 (O_2246,N_24180,N_24076);
or UO_2247 (O_2247,N_24983,N_24715);
xor UO_2248 (O_2248,N_24944,N_24800);
nand UO_2249 (O_2249,N_24217,N_24992);
or UO_2250 (O_2250,N_24715,N_24050);
or UO_2251 (O_2251,N_24994,N_24767);
xor UO_2252 (O_2252,N_24993,N_24412);
nand UO_2253 (O_2253,N_24656,N_24207);
nor UO_2254 (O_2254,N_24556,N_24706);
or UO_2255 (O_2255,N_24230,N_24689);
nand UO_2256 (O_2256,N_24400,N_24669);
nand UO_2257 (O_2257,N_24940,N_24116);
nor UO_2258 (O_2258,N_24145,N_24751);
nor UO_2259 (O_2259,N_24986,N_24039);
nor UO_2260 (O_2260,N_24340,N_24434);
nand UO_2261 (O_2261,N_24221,N_24279);
or UO_2262 (O_2262,N_24753,N_24311);
and UO_2263 (O_2263,N_24340,N_24448);
nand UO_2264 (O_2264,N_24923,N_24060);
and UO_2265 (O_2265,N_24514,N_24152);
xnor UO_2266 (O_2266,N_24617,N_24247);
xor UO_2267 (O_2267,N_24957,N_24596);
nor UO_2268 (O_2268,N_24793,N_24647);
and UO_2269 (O_2269,N_24530,N_24733);
and UO_2270 (O_2270,N_24152,N_24388);
and UO_2271 (O_2271,N_24178,N_24597);
nor UO_2272 (O_2272,N_24210,N_24123);
nor UO_2273 (O_2273,N_24753,N_24474);
nand UO_2274 (O_2274,N_24991,N_24254);
nand UO_2275 (O_2275,N_24821,N_24418);
or UO_2276 (O_2276,N_24296,N_24365);
xnor UO_2277 (O_2277,N_24029,N_24512);
and UO_2278 (O_2278,N_24338,N_24917);
nand UO_2279 (O_2279,N_24958,N_24482);
xnor UO_2280 (O_2280,N_24192,N_24795);
and UO_2281 (O_2281,N_24011,N_24740);
and UO_2282 (O_2282,N_24526,N_24388);
nor UO_2283 (O_2283,N_24634,N_24338);
nor UO_2284 (O_2284,N_24368,N_24118);
xor UO_2285 (O_2285,N_24441,N_24164);
xnor UO_2286 (O_2286,N_24250,N_24824);
and UO_2287 (O_2287,N_24431,N_24800);
nor UO_2288 (O_2288,N_24689,N_24427);
and UO_2289 (O_2289,N_24078,N_24969);
nor UO_2290 (O_2290,N_24984,N_24924);
xor UO_2291 (O_2291,N_24929,N_24719);
nor UO_2292 (O_2292,N_24913,N_24814);
xnor UO_2293 (O_2293,N_24022,N_24244);
or UO_2294 (O_2294,N_24811,N_24899);
nor UO_2295 (O_2295,N_24219,N_24353);
or UO_2296 (O_2296,N_24638,N_24442);
and UO_2297 (O_2297,N_24558,N_24589);
xor UO_2298 (O_2298,N_24893,N_24394);
nand UO_2299 (O_2299,N_24907,N_24564);
or UO_2300 (O_2300,N_24498,N_24797);
nand UO_2301 (O_2301,N_24262,N_24739);
nand UO_2302 (O_2302,N_24506,N_24546);
nand UO_2303 (O_2303,N_24291,N_24786);
or UO_2304 (O_2304,N_24445,N_24540);
nand UO_2305 (O_2305,N_24363,N_24658);
nand UO_2306 (O_2306,N_24150,N_24610);
or UO_2307 (O_2307,N_24706,N_24626);
xnor UO_2308 (O_2308,N_24689,N_24330);
xor UO_2309 (O_2309,N_24990,N_24738);
nand UO_2310 (O_2310,N_24028,N_24736);
xnor UO_2311 (O_2311,N_24603,N_24388);
nand UO_2312 (O_2312,N_24935,N_24887);
and UO_2313 (O_2313,N_24707,N_24448);
nor UO_2314 (O_2314,N_24426,N_24711);
and UO_2315 (O_2315,N_24016,N_24342);
or UO_2316 (O_2316,N_24693,N_24274);
or UO_2317 (O_2317,N_24500,N_24784);
or UO_2318 (O_2318,N_24940,N_24069);
and UO_2319 (O_2319,N_24978,N_24501);
and UO_2320 (O_2320,N_24507,N_24546);
nor UO_2321 (O_2321,N_24125,N_24482);
nand UO_2322 (O_2322,N_24656,N_24342);
or UO_2323 (O_2323,N_24266,N_24613);
or UO_2324 (O_2324,N_24872,N_24929);
xor UO_2325 (O_2325,N_24833,N_24013);
xnor UO_2326 (O_2326,N_24821,N_24235);
xor UO_2327 (O_2327,N_24347,N_24430);
nor UO_2328 (O_2328,N_24546,N_24416);
nor UO_2329 (O_2329,N_24598,N_24290);
xnor UO_2330 (O_2330,N_24196,N_24896);
nand UO_2331 (O_2331,N_24320,N_24154);
and UO_2332 (O_2332,N_24717,N_24204);
and UO_2333 (O_2333,N_24097,N_24876);
nand UO_2334 (O_2334,N_24489,N_24259);
xor UO_2335 (O_2335,N_24580,N_24765);
or UO_2336 (O_2336,N_24863,N_24321);
xnor UO_2337 (O_2337,N_24468,N_24350);
nor UO_2338 (O_2338,N_24936,N_24775);
and UO_2339 (O_2339,N_24891,N_24979);
nand UO_2340 (O_2340,N_24908,N_24508);
or UO_2341 (O_2341,N_24948,N_24304);
xnor UO_2342 (O_2342,N_24651,N_24184);
xor UO_2343 (O_2343,N_24468,N_24659);
nor UO_2344 (O_2344,N_24915,N_24443);
xnor UO_2345 (O_2345,N_24273,N_24901);
nor UO_2346 (O_2346,N_24283,N_24360);
nor UO_2347 (O_2347,N_24476,N_24737);
nand UO_2348 (O_2348,N_24486,N_24963);
nor UO_2349 (O_2349,N_24157,N_24267);
nand UO_2350 (O_2350,N_24334,N_24121);
and UO_2351 (O_2351,N_24774,N_24359);
xnor UO_2352 (O_2352,N_24828,N_24222);
nor UO_2353 (O_2353,N_24887,N_24410);
or UO_2354 (O_2354,N_24635,N_24214);
xor UO_2355 (O_2355,N_24561,N_24784);
or UO_2356 (O_2356,N_24382,N_24497);
xor UO_2357 (O_2357,N_24581,N_24197);
xor UO_2358 (O_2358,N_24781,N_24760);
and UO_2359 (O_2359,N_24311,N_24397);
and UO_2360 (O_2360,N_24601,N_24110);
nor UO_2361 (O_2361,N_24378,N_24405);
or UO_2362 (O_2362,N_24037,N_24161);
nand UO_2363 (O_2363,N_24439,N_24400);
and UO_2364 (O_2364,N_24286,N_24480);
or UO_2365 (O_2365,N_24156,N_24790);
xor UO_2366 (O_2366,N_24727,N_24734);
nor UO_2367 (O_2367,N_24916,N_24662);
nor UO_2368 (O_2368,N_24703,N_24232);
nor UO_2369 (O_2369,N_24282,N_24367);
xnor UO_2370 (O_2370,N_24553,N_24044);
xnor UO_2371 (O_2371,N_24622,N_24904);
nor UO_2372 (O_2372,N_24521,N_24385);
or UO_2373 (O_2373,N_24876,N_24332);
nor UO_2374 (O_2374,N_24052,N_24274);
nor UO_2375 (O_2375,N_24830,N_24870);
and UO_2376 (O_2376,N_24337,N_24385);
or UO_2377 (O_2377,N_24378,N_24551);
or UO_2378 (O_2378,N_24912,N_24386);
and UO_2379 (O_2379,N_24730,N_24710);
and UO_2380 (O_2380,N_24206,N_24726);
nand UO_2381 (O_2381,N_24847,N_24482);
nor UO_2382 (O_2382,N_24404,N_24999);
or UO_2383 (O_2383,N_24108,N_24279);
nand UO_2384 (O_2384,N_24934,N_24365);
nand UO_2385 (O_2385,N_24348,N_24560);
nand UO_2386 (O_2386,N_24571,N_24109);
xnor UO_2387 (O_2387,N_24438,N_24561);
nand UO_2388 (O_2388,N_24977,N_24177);
xnor UO_2389 (O_2389,N_24725,N_24410);
nor UO_2390 (O_2390,N_24592,N_24043);
or UO_2391 (O_2391,N_24836,N_24889);
nor UO_2392 (O_2392,N_24129,N_24917);
nor UO_2393 (O_2393,N_24807,N_24252);
nand UO_2394 (O_2394,N_24629,N_24489);
and UO_2395 (O_2395,N_24736,N_24014);
nand UO_2396 (O_2396,N_24557,N_24670);
nand UO_2397 (O_2397,N_24016,N_24118);
nor UO_2398 (O_2398,N_24184,N_24165);
xor UO_2399 (O_2399,N_24213,N_24255);
nand UO_2400 (O_2400,N_24223,N_24728);
and UO_2401 (O_2401,N_24241,N_24175);
nand UO_2402 (O_2402,N_24469,N_24921);
or UO_2403 (O_2403,N_24846,N_24095);
nor UO_2404 (O_2404,N_24667,N_24509);
or UO_2405 (O_2405,N_24212,N_24628);
nor UO_2406 (O_2406,N_24004,N_24017);
nand UO_2407 (O_2407,N_24596,N_24030);
and UO_2408 (O_2408,N_24875,N_24408);
nor UO_2409 (O_2409,N_24131,N_24986);
xnor UO_2410 (O_2410,N_24075,N_24876);
nand UO_2411 (O_2411,N_24158,N_24585);
or UO_2412 (O_2412,N_24144,N_24395);
or UO_2413 (O_2413,N_24716,N_24973);
xor UO_2414 (O_2414,N_24656,N_24910);
xnor UO_2415 (O_2415,N_24260,N_24705);
or UO_2416 (O_2416,N_24520,N_24902);
xor UO_2417 (O_2417,N_24833,N_24288);
xor UO_2418 (O_2418,N_24300,N_24983);
xor UO_2419 (O_2419,N_24715,N_24954);
nand UO_2420 (O_2420,N_24319,N_24387);
and UO_2421 (O_2421,N_24114,N_24620);
or UO_2422 (O_2422,N_24409,N_24545);
xor UO_2423 (O_2423,N_24539,N_24852);
or UO_2424 (O_2424,N_24364,N_24575);
and UO_2425 (O_2425,N_24557,N_24650);
and UO_2426 (O_2426,N_24143,N_24171);
nor UO_2427 (O_2427,N_24100,N_24496);
nor UO_2428 (O_2428,N_24335,N_24992);
nand UO_2429 (O_2429,N_24533,N_24550);
xnor UO_2430 (O_2430,N_24553,N_24426);
nor UO_2431 (O_2431,N_24025,N_24017);
xor UO_2432 (O_2432,N_24882,N_24326);
xor UO_2433 (O_2433,N_24934,N_24813);
and UO_2434 (O_2434,N_24383,N_24969);
or UO_2435 (O_2435,N_24040,N_24467);
nand UO_2436 (O_2436,N_24520,N_24104);
or UO_2437 (O_2437,N_24153,N_24135);
xor UO_2438 (O_2438,N_24718,N_24704);
nor UO_2439 (O_2439,N_24563,N_24330);
nor UO_2440 (O_2440,N_24650,N_24635);
xnor UO_2441 (O_2441,N_24109,N_24278);
nor UO_2442 (O_2442,N_24590,N_24568);
and UO_2443 (O_2443,N_24575,N_24311);
nand UO_2444 (O_2444,N_24429,N_24860);
xnor UO_2445 (O_2445,N_24661,N_24438);
and UO_2446 (O_2446,N_24006,N_24193);
xor UO_2447 (O_2447,N_24702,N_24823);
and UO_2448 (O_2448,N_24545,N_24390);
or UO_2449 (O_2449,N_24442,N_24042);
or UO_2450 (O_2450,N_24688,N_24115);
xnor UO_2451 (O_2451,N_24773,N_24684);
nor UO_2452 (O_2452,N_24716,N_24875);
and UO_2453 (O_2453,N_24958,N_24966);
or UO_2454 (O_2454,N_24429,N_24534);
or UO_2455 (O_2455,N_24619,N_24688);
or UO_2456 (O_2456,N_24440,N_24481);
nand UO_2457 (O_2457,N_24704,N_24605);
or UO_2458 (O_2458,N_24435,N_24213);
nand UO_2459 (O_2459,N_24904,N_24619);
xnor UO_2460 (O_2460,N_24911,N_24690);
or UO_2461 (O_2461,N_24862,N_24381);
nand UO_2462 (O_2462,N_24045,N_24421);
and UO_2463 (O_2463,N_24357,N_24682);
nand UO_2464 (O_2464,N_24434,N_24247);
or UO_2465 (O_2465,N_24588,N_24678);
and UO_2466 (O_2466,N_24931,N_24528);
nand UO_2467 (O_2467,N_24026,N_24503);
or UO_2468 (O_2468,N_24238,N_24399);
and UO_2469 (O_2469,N_24742,N_24725);
or UO_2470 (O_2470,N_24980,N_24055);
xnor UO_2471 (O_2471,N_24715,N_24312);
nor UO_2472 (O_2472,N_24512,N_24686);
nand UO_2473 (O_2473,N_24463,N_24698);
and UO_2474 (O_2474,N_24270,N_24578);
nand UO_2475 (O_2475,N_24666,N_24059);
nor UO_2476 (O_2476,N_24187,N_24730);
or UO_2477 (O_2477,N_24271,N_24069);
or UO_2478 (O_2478,N_24986,N_24932);
nor UO_2479 (O_2479,N_24631,N_24467);
and UO_2480 (O_2480,N_24436,N_24122);
or UO_2481 (O_2481,N_24889,N_24532);
or UO_2482 (O_2482,N_24459,N_24940);
or UO_2483 (O_2483,N_24015,N_24365);
nand UO_2484 (O_2484,N_24987,N_24373);
and UO_2485 (O_2485,N_24121,N_24135);
nor UO_2486 (O_2486,N_24412,N_24444);
xnor UO_2487 (O_2487,N_24625,N_24754);
nor UO_2488 (O_2488,N_24118,N_24780);
xnor UO_2489 (O_2489,N_24918,N_24186);
and UO_2490 (O_2490,N_24287,N_24111);
nand UO_2491 (O_2491,N_24123,N_24873);
and UO_2492 (O_2492,N_24702,N_24320);
xnor UO_2493 (O_2493,N_24438,N_24845);
or UO_2494 (O_2494,N_24120,N_24308);
nand UO_2495 (O_2495,N_24478,N_24110);
xnor UO_2496 (O_2496,N_24189,N_24846);
xnor UO_2497 (O_2497,N_24890,N_24300);
nand UO_2498 (O_2498,N_24293,N_24721);
and UO_2499 (O_2499,N_24889,N_24132);
or UO_2500 (O_2500,N_24326,N_24029);
nand UO_2501 (O_2501,N_24040,N_24645);
nand UO_2502 (O_2502,N_24794,N_24660);
nand UO_2503 (O_2503,N_24306,N_24002);
and UO_2504 (O_2504,N_24006,N_24410);
or UO_2505 (O_2505,N_24430,N_24696);
or UO_2506 (O_2506,N_24849,N_24453);
xor UO_2507 (O_2507,N_24867,N_24499);
xor UO_2508 (O_2508,N_24999,N_24989);
xor UO_2509 (O_2509,N_24220,N_24425);
xnor UO_2510 (O_2510,N_24612,N_24413);
and UO_2511 (O_2511,N_24559,N_24762);
or UO_2512 (O_2512,N_24765,N_24606);
nor UO_2513 (O_2513,N_24275,N_24323);
or UO_2514 (O_2514,N_24826,N_24774);
nand UO_2515 (O_2515,N_24724,N_24410);
xnor UO_2516 (O_2516,N_24257,N_24082);
nor UO_2517 (O_2517,N_24145,N_24987);
and UO_2518 (O_2518,N_24532,N_24020);
or UO_2519 (O_2519,N_24187,N_24620);
nand UO_2520 (O_2520,N_24437,N_24466);
xnor UO_2521 (O_2521,N_24499,N_24330);
or UO_2522 (O_2522,N_24982,N_24180);
or UO_2523 (O_2523,N_24246,N_24494);
and UO_2524 (O_2524,N_24814,N_24296);
or UO_2525 (O_2525,N_24784,N_24713);
or UO_2526 (O_2526,N_24461,N_24450);
or UO_2527 (O_2527,N_24740,N_24723);
nand UO_2528 (O_2528,N_24291,N_24226);
nor UO_2529 (O_2529,N_24028,N_24392);
nand UO_2530 (O_2530,N_24202,N_24954);
xor UO_2531 (O_2531,N_24311,N_24619);
nand UO_2532 (O_2532,N_24455,N_24697);
nor UO_2533 (O_2533,N_24128,N_24443);
or UO_2534 (O_2534,N_24408,N_24353);
nand UO_2535 (O_2535,N_24271,N_24038);
nand UO_2536 (O_2536,N_24559,N_24091);
and UO_2537 (O_2537,N_24580,N_24013);
xnor UO_2538 (O_2538,N_24672,N_24208);
nand UO_2539 (O_2539,N_24632,N_24008);
nor UO_2540 (O_2540,N_24635,N_24952);
xor UO_2541 (O_2541,N_24046,N_24356);
nor UO_2542 (O_2542,N_24195,N_24991);
and UO_2543 (O_2543,N_24564,N_24365);
nand UO_2544 (O_2544,N_24139,N_24809);
xnor UO_2545 (O_2545,N_24450,N_24688);
and UO_2546 (O_2546,N_24818,N_24057);
nand UO_2547 (O_2547,N_24464,N_24737);
nor UO_2548 (O_2548,N_24863,N_24473);
xor UO_2549 (O_2549,N_24526,N_24744);
and UO_2550 (O_2550,N_24097,N_24752);
and UO_2551 (O_2551,N_24907,N_24751);
nor UO_2552 (O_2552,N_24736,N_24911);
and UO_2553 (O_2553,N_24712,N_24811);
or UO_2554 (O_2554,N_24571,N_24917);
nand UO_2555 (O_2555,N_24166,N_24669);
or UO_2556 (O_2556,N_24823,N_24852);
nor UO_2557 (O_2557,N_24130,N_24796);
xor UO_2558 (O_2558,N_24263,N_24133);
and UO_2559 (O_2559,N_24907,N_24909);
and UO_2560 (O_2560,N_24276,N_24256);
or UO_2561 (O_2561,N_24174,N_24579);
nor UO_2562 (O_2562,N_24693,N_24900);
or UO_2563 (O_2563,N_24263,N_24452);
xnor UO_2564 (O_2564,N_24667,N_24669);
xnor UO_2565 (O_2565,N_24867,N_24826);
nor UO_2566 (O_2566,N_24866,N_24277);
or UO_2567 (O_2567,N_24143,N_24580);
nand UO_2568 (O_2568,N_24727,N_24986);
and UO_2569 (O_2569,N_24896,N_24751);
xnor UO_2570 (O_2570,N_24968,N_24481);
or UO_2571 (O_2571,N_24217,N_24636);
xor UO_2572 (O_2572,N_24183,N_24752);
nand UO_2573 (O_2573,N_24220,N_24555);
nor UO_2574 (O_2574,N_24998,N_24689);
nor UO_2575 (O_2575,N_24118,N_24524);
and UO_2576 (O_2576,N_24134,N_24624);
nor UO_2577 (O_2577,N_24209,N_24929);
and UO_2578 (O_2578,N_24537,N_24048);
or UO_2579 (O_2579,N_24945,N_24650);
or UO_2580 (O_2580,N_24277,N_24170);
nor UO_2581 (O_2581,N_24722,N_24215);
xnor UO_2582 (O_2582,N_24502,N_24978);
nor UO_2583 (O_2583,N_24803,N_24995);
and UO_2584 (O_2584,N_24235,N_24448);
and UO_2585 (O_2585,N_24386,N_24817);
or UO_2586 (O_2586,N_24663,N_24731);
and UO_2587 (O_2587,N_24216,N_24025);
nor UO_2588 (O_2588,N_24889,N_24472);
and UO_2589 (O_2589,N_24037,N_24617);
nor UO_2590 (O_2590,N_24631,N_24177);
nand UO_2591 (O_2591,N_24918,N_24914);
and UO_2592 (O_2592,N_24179,N_24486);
and UO_2593 (O_2593,N_24562,N_24150);
or UO_2594 (O_2594,N_24959,N_24866);
or UO_2595 (O_2595,N_24607,N_24810);
nor UO_2596 (O_2596,N_24899,N_24710);
nand UO_2597 (O_2597,N_24188,N_24837);
nand UO_2598 (O_2598,N_24233,N_24443);
and UO_2599 (O_2599,N_24941,N_24975);
nand UO_2600 (O_2600,N_24451,N_24904);
or UO_2601 (O_2601,N_24057,N_24429);
and UO_2602 (O_2602,N_24173,N_24934);
or UO_2603 (O_2603,N_24093,N_24660);
nor UO_2604 (O_2604,N_24838,N_24884);
nand UO_2605 (O_2605,N_24270,N_24187);
and UO_2606 (O_2606,N_24494,N_24828);
nand UO_2607 (O_2607,N_24643,N_24842);
xor UO_2608 (O_2608,N_24796,N_24777);
nor UO_2609 (O_2609,N_24235,N_24404);
xor UO_2610 (O_2610,N_24756,N_24314);
or UO_2611 (O_2611,N_24402,N_24997);
xor UO_2612 (O_2612,N_24473,N_24105);
nor UO_2613 (O_2613,N_24832,N_24769);
nand UO_2614 (O_2614,N_24055,N_24373);
xnor UO_2615 (O_2615,N_24840,N_24454);
or UO_2616 (O_2616,N_24690,N_24729);
xor UO_2617 (O_2617,N_24648,N_24644);
nand UO_2618 (O_2618,N_24304,N_24385);
nand UO_2619 (O_2619,N_24035,N_24004);
nand UO_2620 (O_2620,N_24222,N_24917);
or UO_2621 (O_2621,N_24510,N_24503);
nand UO_2622 (O_2622,N_24199,N_24546);
and UO_2623 (O_2623,N_24310,N_24926);
and UO_2624 (O_2624,N_24795,N_24764);
nor UO_2625 (O_2625,N_24455,N_24955);
nand UO_2626 (O_2626,N_24697,N_24122);
nand UO_2627 (O_2627,N_24190,N_24358);
and UO_2628 (O_2628,N_24913,N_24672);
nand UO_2629 (O_2629,N_24583,N_24022);
or UO_2630 (O_2630,N_24390,N_24774);
or UO_2631 (O_2631,N_24706,N_24612);
nor UO_2632 (O_2632,N_24285,N_24455);
or UO_2633 (O_2633,N_24899,N_24068);
or UO_2634 (O_2634,N_24566,N_24174);
nand UO_2635 (O_2635,N_24948,N_24723);
or UO_2636 (O_2636,N_24325,N_24874);
and UO_2637 (O_2637,N_24388,N_24962);
nor UO_2638 (O_2638,N_24517,N_24616);
or UO_2639 (O_2639,N_24192,N_24560);
or UO_2640 (O_2640,N_24958,N_24372);
nor UO_2641 (O_2641,N_24635,N_24414);
and UO_2642 (O_2642,N_24005,N_24874);
and UO_2643 (O_2643,N_24309,N_24762);
xnor UO_2644 (O_2644,N_24728,N_24824);
nor UO_2645 (O_2645,N_24694,N_24518);
nor UO_2646 (O_2646,N_24201,N_24949);
nor UO_2647 (O_2647,N_24891,N_24887);
nor UO_2648 (O_2648,N_24578,N_24402);
nor UO_2649 (O_2649,N_24350,N_24209);
nor UO_2650 (O_2650,N_24837,N_24362);
xor UO_2651 (O_2651,N_24018,N_24630);
nor UO_2652 (O_2652,N_24238,N_24482);
nor UO_2653 (O_2653,N_24222,N_24397);
or UO_2654 (O_2654,N_24679,N_24278);
nand UO_2655 (O_2655,N_24859,N_24630);
and UO_2656 (O_2656,N_24095,N_24775);
xor UO_2657 (O_2657,N_24543,N_24035);
or UO_2658 (O_2658,N_24184,N_24825);
xor UO_2659 (O_2659,N_24333,N_24346);
nor UO_2660 (O_2660,N_24671,N_24809);
nor UO_2661 (O_2661,N_24322,N_24567);
xor UO_2662 (O_2662,N_24591,N_24326);
nor UO_2663 (O_2663,N_24697,N_24260);
xor UO_2664 (O_2664,N_24087,N_24244);
nor UO_2665 (O_2665,N_24333,N_24788);
nor UO_2666 (O_2666,N_24369,N_24065);
nor UO_2667 (O_2667,N_24221,N_24575);
and UO_2668 (O_2668,N_24775,N_24614);
or UO_2669 (O_2669,N_24352,N_24984);
nand UO_2670 (O_2670,N_24211,N_24730);
xnor UO_2671 (O_2671,N_24119,N_24657);
nor UO_2672 (O_2672,N_24800,N_24681);
or UO_2673 (O_2673,N_24979,N_24727);
nor UO_2674 (O_2674,N_24077,N_24488);
xor UO_2675 (O_2675,N_24452,N_24588);
nand UO_2676 (O_2676,N_24449,N_24876);
nand UO_2677 (O_2677,N_24133,N_24191);
and UO_2678 (O_2678,N_24743,N_24471);
nand UO_2679 (O_2679,N_24550,N_24313);
nand UO_2680 (O_2680,N_24862,N_24115);
xnor UO_2681 (O_2681,N_24961,N_24452);
xor UO_2682 (O_2682,N_24999,N_24442);
nor UO_2683 (O_2683,N_24014,N_24041);
xor UO_2684 (O_2684,N_24348,N_24715);
nand UO_2685 (O_2685,N_24588,N_24857);
or UO_2686 (O_2686,N_24946,N_24533);
nor UO_2687 (O_2687,N_24437,N_24602);
nor UO_2688 (O_2688,N_24577,N_24560);
and UO_2689 (O_2689,N_24310,N_24400);
and UO_2690 (O_2690,N_24730,N_24764);
nand UO_2691 (O_2691,N_24657,N_24168);
nand UO_2692 (O_2692,N_24448,N_24953);
nand UO_2693 (O_2693,N_24317,N_24810);
nand UO_2694 (O_2694,N_24685,N_24734);
nand UO_2695 (O_2695,N_24194,N_24478);
nor UO_2696 (O_2696,N_24049,N_24912);
and UO_2697 (O_2697,N_24026,N_24374);
nor UO_2698 (O_2698,N_24413,N_24223);
and UO_2699 (O_2699,N_24498,N_24916);
nor UO_2700 (O_2700,N_24157,N_24107);
xor UO_2701 (O_2701,N_24499,N_24740);
nand UO_2702 (O_2702,N_24811,N_24211);
nor UO_2703 (O_2703,N_24969,N_24415);
xor UO_2704 (O_2704,N_24296,N_24369);
nor UO_2705 (O_2705,N_24927,N_24776);
xnor UO_2706 (O_2706,N_24582,N_24670);
and UO_2707 (O_2707,N_24193,N_24069);
xor UO_2708 (O_2708,N_24582,N_24563);
or UO_2709 (O_2709,N_24309,N_24556);
nand UO_2710 (O_2710,N_24058,N_24215);
and UO_2711 (O_2711,N_24259,N_24296);
and UO_2712 (O_2712,N_24607,N_24110);
xnor UO_2713 (O_2713,N_24923,N_24967);
or UO_2714 (O_2714,N_24028,N_24512);
nor UO_2715 (O_2715,N_24581,N_24623);
and UO_2716 (O_2716,N_24808,N_24887);
nor UO_2717 (O_2717,N_24430,N_24461);
xor UO_2718 (O_2718,N_24226,N_24129);
or UO_2719 (O_2719,N_24615,N_24980);
and UO_2720 (O_2720,N_24219,N_24117);
nand UO_2721 (O_2721,N_24799,N_24168);
or UO_2722 (O_2722,N_24194,N_24970);
nand UO_2723 (O_2723,N_24903,N_24601);
nand UO_2724 (O_2724,N_24567,N_24041);
nand UO_2725 (O_2725,N_24873,N_24903);
xor UO_2726 (O_2726,N_24760,N_24765);
or UO_2727 (O_2727,N_24689,N_24784);
xnor UO_2728 (O_2728,N_24609,N_24443);
or UO_2729 (O_2729,N_24645,N_24801);
or UO_2730 (O_2730,N_24208,N_24586);
nor UO_2731 (O_2731,N_24600,N_24450);
or UO_2732 (O_2732,N_24179,N_24372);
nor UO_2733 (O_2733,N_24051,N_24743);
and UO_2734 (O_2734,N_24248,N_24200);
and UO_2735 (O_2735,N_24638,N_24930);
and UO_2736 (O_2736,N_24723,N_24731);
and UO_2737 (O_2737,N_24745,N_24479);
xnor UO_2738 (O_2738,N_24715,N_24287);
or UO_2739 (O_2739,N_24251,N_24511);
nand UO_2740 (O_2740,N_24225,N_24336);
xnor UO_2741 (O_2741,N_24267,N_24547);
and UO_2742 (O_2742,N_24155,N_24737);
xor UO_2743 (O_2743,N_24372,N_24209);
nor UO_2744 (O_2744,N_24731,N_24372);
nand UO_2745 (O_2745,N_24808,N_24832);
and UO_2746 (O_2746,N_24485,N_24921);
xnor UO_2747 (O_2747,N_24692,N_24663);
and UO_2748 (O_2748,N_24498,N_24165);
nand UO_2749 (O_2749,N_24075,N_24632);
nor UO_2750 (O_2750,N_24362,N_24853);
and UO_2751 (O_2751,N_24888,N_24260);
nand UO_2752 (O_2752,N_24185,N_24955);
or UO_2753 (O_2753,N_24895,N_24446);
nor UO_2754 (O_2754,N_24838,N_24675);
nand UO_2755 (O_2755,N_24079,N_24743);
and UO_2756 (O_2756,N_24883,N_24865);
nand UO_2757 (O_2757,N_24219,N_24299);
and UO_2758 (O_2758,N_24457,N_24427);
and UO_2759 (O_2759,N_24401,N_24645);
nand UO_2760 (O_2760,N_24219,N_24368);
and UO_2761 (O_2761,N_24845,N_24059);
xor UO_2762 (O_2762,N_24104,N_24389);
nand UO_2763 (O_2763,N_24967,N_24410);
xor UO_2764 (O_2764,N_24003,N_24883);
and UO_2765 (O_2765,N_24048,N_24361);
or UO_2766 (O_2766,N_24505,N_24812);
or UO_2767 (O_2767,N_24595,N_24706);
or UO_2768 (O_2768,N_24075,N_24028);
or UO_2769 (O_2769,N_24143,N_24651);
or UO_2770 (O_2770,N_24902,N_24722);
or UO_2771 (O_2771,N_24223,N_24873);
nand UO_2772 (O_2772,N_24125,N_24352);
nand UO_2773 (O_2773,N_24559,N_24173);
nand UO_2774 (O_2774,N_24123,N_24424);
xor UO_2775 (O_2775,N_24477,N_24103);
or UO_2776 (O_2776,N_24188,N_24339);
or UO_2777 (O_2777,N_24843,N_24643);
and UO_2778 (O_2778,N_24213,N_24425);
nor UO_2779 (O_2779,N_24993,N_24906);
nand UO_2780 (O_2780,N_24765,N_24068);
or UO_2781 (O_2781,N_24109,N_24602);
and UO_2782 (O_2782,N_24176,N_24698);
nor UO_2783 (O_2783,N_24944,N_24964);
and UO_2784 (O_2784,N_24510,N_24733);
or UO_2785 (O_2785,N_24481,N_24186);
or UO_2786 (O_2786,N_24596,N_24634);
nand UO_2787 (O_2787,N_24982,N_24953);
or UO_2788 (O_2788,N_24900,N_24053);
or UO_2789 (O_2789,N_24935,N_24903);
nor UO_2790 (O_2790,N_24988,N_24885);
and UO_2791 (O_2791,N_24955,N_24458);
xnor UO_2792 (O_2792,N_24738,N_24967);
and UO_2793 (O_2793,N_24877,N_24727);
xor UO_2794 (O_2794,N_24842,N_24109);
xor UO_2795 (O_2795,N_24325,N_24279);
or UO_2796 (O_2796,N_24382,N_24208);
and UO_2797 (O_2797,N_24231,N_24893);
nor UO_2798 (O_2798,N_24039,N_24294);
and UO_2799 (O_2799,N_24478,N_24857);
xnor UO_2800 (O_2800,N_24317,N_24288);
and UO_2801 (O_2801,N_24666,N_24904);
or UO_2802 (O_2802,N_24378,N_24125);
xor UO_2803 (O_2803,N_24664,N_24776);
xor UO_2804 (O_2804,N_24968,N_24302);
nor UO_2805 (O_2805,N_24910,N_24070);
or UO_2806 (O_2806,N_24601,N_24753);
or UO_2807 (O_2807,N_24950,N_24613);
or UO_2808 (O_2808,N_24271,N_24334);
nor UO_2809 (O_2809,N_24444,N_24165);
nor UO_2810 (O_2810,N_24905,N_24928);
nor UO_2811 (O_2811,N_24484,N_24449);
nor UO_2812 (O_2812,N_24436,N_24526);
and UO_2813 (O_2813,N_24284,N_24055);
xnor UO_2814 (O_2814,N_24989,N_24564);
nand UO_2815 (O_2815,N_24298,N_24386);
xor UO_2816 (O_2816,N_24571,N_24993);
xor UO_2817 (O_2817,N_24343,N_24759);
and UO_2818 (O_2818,N_24245,N_24585);
nand UO_2819 (O_2819,N_24935,N_24825);
nand UO_2820 (O_2820,N_24197,N_24280);
xor UO_2821 (O_2821,N_24256,N_24778);
nand UO_2822 (O_2822,N_24597,N_24039);
xor UO_2823 (O_2823,N_24314,N_24583);
or UO_2824 (O_2824,N_24798,N_24363);
and UO_2825 (O_2825,N_24076,N_24750);
xor UO_2826 (O_2826,N_24011,N_24095);
nor UO_2827 (O_2827,N_24628,N_24990);
nor UO_2828 (O_2828,N_24568,N_24451);
nor UO_2829 (O_2829,N_24748,N_24879);
nand UO_2830 (O_2830,N_24469,N_24626);
nor UO_2831 (O_2831,N_24617,N_24525);
or UO_2832 (O_2832,N_24010,N_24006);
and UO_2833 (O_2833,N_24297,N_24816);
and UO_2834 (O_2834,N_24479,N_24721);
and UO_2835 (O_2835,N_24317,N_24474);
nand UO_2836 (O_2836,N_24119,N_24804);
and UO_2837 (O_2837,N_24523,N_24193);
nand UO_2838 (O_2838,N_24457,N_24643);
or UO_2839 (O_2839,N_24124,N_24121);
nor UO_2840 (O_2840,N_24103,N_24889);
xor UO_2841 (O_2841,N_24047,N_24642);
and UO_2842 (O_2842,N_24025,N_24922);
and UO_2843 (O_2843,N_24971,N_24491);
nand UO_2844 (O_2844,N_24316,N_24536);
nor UO_2845 (O_2845,N_24639,N_24800);
and UO_2846 (O_2846,N_24034,N_24793);
nand UO_2847 (O_2847,N_24217,N_24787);
xnor UO_2848 (O_2848,N_24813,N_24608);
nor UO_2849 (O_2849,N_24177,N_24108);
nor UO_2850 (O_2850,N_24915,N_24343);
or UO_2851 (O_2851,N_24346,N_24141);
nor UO_2852 (O_2852,N_24581,N_24692);
nand UO_2853 (O_2853,N_24975,N_24164);
nor UO_2854 (O_2854,N_24676,N_24881);
xor UO_2855 (O_2855,N_24447,N_24017);
or UO_2856 (O_2856,N_24808,N_24534);
and UO_2857 (O_2857,N_24853,N_24543);
xor UO_2858 (O_2858,N_24954,N_24028);
and UO_2859 (O_2859,N_24335,N_24589);
nand UO_2860 (O_2860,N_24197,N_24029);
and UO_2861 (O_2861,N_24374,N_24358);
and UO_2862 (O_2862,N_24814,N_24592);
nand UO_2863 (O_2863,N_24472,N_24786);
or UO_2864 (O_2864,N_24172,N_24292);
and UO_2865 (O_2865,N_24835,N_24908);
xnor UO_2866 (O_2866,N_24533,N_24220);
xor UO_2867 (O_2867,N_24587,N_24535);
and UO_2868 (O_2868,N_24357,N_24624);
or UO_2869 (O_2869,N_24465,N_24763);
nand UO_2870 (O_2870,N_24517,N_24234);
or UO_2871 (O_2871,N_24572,N_24733);
nor UO_2872 (O_2872,N_24109,N_24343);
xnor UO_2873 (O_2873,N_24619,N_24567);
xnor UO_2874 (O_2874,N_24948,N_24413);
and UO_2875 (O_2875,N_24951,N_24655);
nor UO_2876 (O_2876,N_24666,N_24871);
or UO_2877 (O_2877,N_24448,N_24851);
nor UO_2878 (O_2878,N_24144,N_24691);
nand UO_2879 (O_2879,N_24637,N_24632);
xor UO_2880 (O_2880,N_24708,N_24277);
nand UO_2881 (O_2881,N_24337,N_24340);
nand UO_2882 (O_2882,N_24434,N_24394);
nand UO_2883 (O_2883,N_24931,N_24658);
xnor UO_2884 (O_2884,N_24400,N_24266);
nor UO_2885 (O_2885,N_24761,N_24177);
nor UO_2886 (O_2886,N_24777,N_24695);
nor UO_2887 (O_2887,N_24930,N_24553);
xor UO_2888 (O_2888,N_24203,N_24534);
nor UO_2889 (O_2889,N_24953,N_24849);
nand UO_2890 (O_2890,N_24721,N_24569);
nor UO_2891 (O_2891,N_24655,N_24138);
xor UO_2892 (O_2892,N_24463,N_24876);
xor UO_2893 (O_2893,N_24356,N_24580);
xnor UO_2894 (O_2894,N_24989,N_24610);
nor UO_2895 (O_2895,N_24553,N_24914);
or UO_2896 (O_2896,N_24991,N_24911);
and UO_2897 (O_2897,N_24178,N_24879);
and UO_2898 (O_2898,N_24359,N_24033);
and UO_2899 (O_2899,N_24463,N_24509);
and UO_2900 (O_2900,N_24767,N_24681);
and UO_2901 (O_2901,N_24391,N_24087);
xnor UO_2902 (O_2902,N_24311,N_24494);
nor UO_2903 (O_2903,N_24089,N_24468);
and UO_2904 (O_2904,N_24862,N_24002);
or UO_2905 (O_2905,N_24117,N_24047);
nor UO_2906 (O_2906,N_24787,N_24369);
and UO_2907 (O_2907,N_24620,N_24322);
nand UO_2908 (O_2908,N_24715,N_24898);
xor UO_2909 (O_2909,N_24303,N_24449);
nor UO_2910 (O_2910,N_24035,N_24531);
and UO_2911 (O_2911,N_24696,N_24819);
nor UO_2912 (O_2912,N_24251,N_24325);
and UO_2913 (O_2913,N_24431,N_24848);
nor UO_2914 (O_2914,N_24580,N_24117);
xnor UO_2915 (O_2915,N_24160,N_24077);
nor UO_2916 (O_2916,N_24801,N_24943);
or UO_2917 (O_2917,N_24107,N_24296);
or UO_2918 (O_2918,N_24881,N_24234);
and UO_2919 (O_2919,N_24927,N_24183);
nand UO_2920 (O_2920,N_24181,N_24997);
xnor UO_2921 (O_2921,N_24108,N_24067);
or UO_2922 (O_2922,N_24354,N_24928);
or UO_2923 (O_2923,N_24754,N_24683);
nand UO_2924 (O_2924,N_24361,N_24245);
nand UO_2925 (O_2925,N_24686,N_24552);
and UO_2926 (O_2926,N_24326,N_24628);
and UO_2927 (O_2927,N_24555,N_24623);
or UO_2928 (O_2928,N_24217,N_24979);
and UO_2929 (O_2929,N_24925,N_24706);
or UO_2930 (O_2930,N_24131,N_24759);
xnor UO_2931 (O_2931,N_24195,N_24361);
nor UO_2932 (O_2932,N_24386,N_24301);
xor UO_2933 (O_2933,N_24338,N_24229);
nor UO_2934 (O_2934,N_24797,N_24472);
nor UO_2935 (O_2935,N_24985,N_24823);
or UO_2936 (O_2936,N_24317,N_24664);
nor UO_2937 (O_2937,N_24247,N_24537);
nor UO_2938 (O_2938,N_24379,N_24094);
or UO_2939 (O_2939,N_24906,N_24871);
nand UO_2940 (O_2940,N_24469,N_24289);
xor UO_2941 (O_2941,N_24615,N_24177);
or UO_2942 (O_2942,N_24544,N_24276);
and UO_2943 (O_2943,N_24004,N_24408);
nand UO_2944 (O_2944,N_24982,N_24295);
or UO_2945 (O_2945,N_24396,N_24673);
xor UO_2946 (O_2946,N_24191,N_24025);
nor UO_2947 (O_2947,N_24792,N_24129);
nor UO_2948 (O_2948,N_24237,N_24638);
nand UO_2949 (O_2949,N_24474,N_24090);
nor UO_2950 (O_2950,N_24909,N_24008);
xnor UO_2951 (O_2951,N_24045,N_24883);
nand UO_2952 (O_2952,N_24038,N_24236);
nand UO_2953 (O_2953,N_24992,N_24357);
or UO_2954 (O_2954,N_24289,N_24705);
nand UO_2955 (O_2955,N_24448,N_24467);
or UO_2956 (O_2956,N_24414,N_24392);
nor UO_2957 (O_2957,N_24274,N_24112);
xor UO_2958 (O_2958,N_24064,N_24742);
and UO_2959 (O_2959,N_24283,N_24164);
nor UO_2960 (O_2960,N_24703,N_24635);
and UO_2961 (O_2961,N_24741,N_24978);
xor UO_2962 (O_2962,N_24124,N_24588);
nand UO_2963 (O_2963,N_24534,N_24773);
nor UO_2964 (O_2964,N_24541,N_24692);
or UO_2965 (O_2965,N_24921,N_24935);
xor UO_2966 (O_2966,N_24574,N_24167);
nand UO_2967 (O_2967,N_24663,N_24275);
and UO_2968 (O_2968,N_24095,N_24718);
and UO_2969 (O_2969,N_24491,N_24095);
nor UO_2970 (O_2970,N_24896,N_24219);
nand UO_2971 (O_2971,N_24493,N_24011);
nor UO_2972 (O_2972,N_24660,N_24055);
nor UO_2973 (O_2973,N_24638,N_24321);
and UO_2974 (O_2974,N_24948,N_24818);
nand UO_2975 (O_2975,N_24261,N_24040);
xnor UO_2976 (O_2976,N_24118,N_24130);
nand UO_2977 (O_2977,N_24934,N_24034);
or UO_2978 (O_2978,N_24309,N_24013);
xor UO_2979 (O_2979,N_24817,N_24428);
nor UO_2980 (O_2980,N_24566,N_24874);
nand UO_2981 (O_2981,N_24715,N_24017);
nand UO_2982 (O_2982,N_24258,N_24265);
or UO_2983 (O_2983,N_24188,N_24297);
xnor UO_2984 (O_2984,N_24828,N_24462);
nand UO_2985 (O_2985,N_24200,N_24589);
xor UO_2986 (O_2986,N_24783,N_24195);
or UO_2987 (O_2987,N_24932,N_24212);
and UO_2988 (O_2988,N_24705,N_24094);
and UO_2989 (O_2989,N_24478,N_24032);
xnor UO_2990 (O_2990,N_24972,N_24822);
and UO_2991 (O_2991,N_24321,N_24298);
nor UO_2992 (O_2992,N_24352,N_24195);
and UO_2993 (O_2993,N_24853,N_24985);
and UO_2994 (O_2994,N_24742,N_24363);
nand UO_2995 (O_2995,N_24345,N_24578);
or UO_2996 (O_2996,N_24053,N_24717);
nor UO_2997 (O_2997,N_24862,N_24653);
nor UO_2998 (O_2998,N_24993,N_24817);
or UO_2999 (O_2999,N_24175,N_24765);
endmodule