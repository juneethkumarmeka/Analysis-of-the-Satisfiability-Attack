module basic_750_5000_1000_2_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2503,N_2504,N_2505,N_2506,N_2507,N_2511,N_2512,N_2513,N_2514,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2526,N_2528,N_2529,N_2530,N_2531,N_2532,N_2534,N_2535,N_2537,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2550,N_2552,N_2553,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2564,N_2565,N_2566,N_2567,N_2568,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2577,N_2578,N_2579,N_2580,N_2581,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2603,N_2604,N_2606,N_2607,N_2608,N_2609,N_2612,N_2613,N_2614,N_2616,N_2617,N_2618,N_2619,N_2620,N_2622,N_2623,N_2624,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2654,N_2655,N_2656,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2665,N_2666,N_2667,N_2668,N_2670,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2688,N_2690,N_2692,N_2694,N_2695,N_2696,N_2697,N_2699,N_2701,N_2702,N_2703,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2715,N_2717,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2757,N_2759,N_2760,N_2761,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2770,N_2771,N_2772,N_2774,N_2776,N_2777,N_2778,N_2780,N_2781,N_2782,N_2783,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2792,N_2793,N_2796,N_2797,N_2798,N_2799,N_2800,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2818,N_2820,N_2822,N_2823,N_2824,N_2826,N_2827,N_2828,N_2829,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2839,N_2840,N_2841,N_2842,N_2843,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2858,N_2859,N_2860,N_2862,N_2863,N_2864,N_2866,N_2867,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2890,N_2891,N_2893,N_2894,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2906,N_2908,N_2910,N_2911,N_2913,N_2914,N_2915,N_2918,N_2919,N_2920,N_2922,N_2923,N_2924,N_2926,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2949,N_2950,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2963,N_2964,N_2965,N_2967,N_2968,N_2969,N_2971,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2997,N_2999,N_3000,N_3002,N_3004,N_3006,N_3007,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3020,N_3021,N_3022,N_3023,N_3024,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3037,N_3038,N_3039,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3087,N_3088,N_3089,N_3090,N_3091,N_3093,N_3095,N_3097,N_3098,N_3099,N_3100,N_3101,N_3103,N_3104,N_3108,N_3109,N_3110,N_3112,N_3113,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3140,N_3141,N_3142,N_3143,N_3144,N_3146,N_3147,N_3148,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3171,N_3172,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3204,N_3205,N_3206,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3216,N_3217,N_3219,N_3220,N_3221,N_3222,N_3224,N_3226,N_3227,N_3228,N_3229,N_3231,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3253,N_3254,N_3256,N_3257,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3268,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3291,N_3292,N_3293,N_3294,N_3295,N_3297,N_3299,N_3300,N_3301,N_3303,N_3304,N_3306,N_3307,N_3308,N_3309,N_3311,N_3312,N_3314,N_3316,N_3317,N_3319,N_3320,N_3321,N_3323,N_3324,N_3326,N_3330,N_3332,N_3333,N_3334,N_3335,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3345,N_3346,N_3348,N_3349,N_3350,N_3353,N_3354,N_3356,N_3357,N_3358,N_3361,N_3362,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3374,N_3375,N_3377,N_3378,N_3379,N_3380,N_3382,N_3383,N_3384,N_3385,N_3387,N_3389,N_3390,N_3391,N_3392,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3403,N_3404,N_3405,N_3406,N_3407,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3436,N_3437,N_3438,N_3439,N_3441,N_3443,N_3444,N_3445,N_3446,N_3448,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3503,N_3505,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3515,N_3517,N_3519,N_3520,N_3521,N_3524,N_3525,N_3526,N_3527,N_3529,N_3531,N_3532,N_3533,N_3535,N_3536,N_3537,N_3538,N_3540,N_3541,N_3542,N_3543,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3570,N_3571,N_3572,N_3574,N_3575,N_3576,N_3577,N_3578,N_3580,N_3582,N_3583,N_3584,N_3586,N_3587,N_3588,N_3590,N_3591,N_3592,N_3593,N_3594,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3606,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3645,N_3646,N_3647,N_3648,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3666,N_3667,N_3668,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3679,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3689,N_3690,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3705,N_3707,N_3708,N_3710,N_3711,N_3712,N_3713,N_3714,N_3716,N_3718,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3728,N_3729,N_3730,N_3731,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3742,N_3743,N_3744,N_3745,N_3746,N_3748,N_3749,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3760,N_3761,N_3762,N_3765,N_3767,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3778,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3788,N_3789,N_3791,N_3792,N_3794,N_3795,N_3796,N_3797,N_3801,N_3802,N_3803,N_3804,N_3805,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3814,N_3815,N_3816,N_3817,N_3819,N_3820,N_3821,N_3822,N_3823,N_3825,N_3826,N_3827,N_3830,N_3831,N_3834,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3849,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3868,N_3871,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3884,N_3885,N_3886,N_3887,N_3888,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3899,N_3900,N_3901,N_3902,N_3904,N_3905,N_3906,N_3908,N_3909,N_3910,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3920,N_3921,N_3922,N_3923,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3938,N_3939,N_3940,N_3941,N_3942,N_3944,N_3945,N_3946,N_3947,N_3949,N_3950,N_3951,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3960,N_3961,N_3963,N_3965,N_3966,N_3967,N_3968,N_3971,N_3972,N_3975,N_3977,N_3978,N_3979,N_3980,N_3981,N_3984,N_3985,N_3987,N_3988,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_4001,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4061,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4080,N_4083,N_4086,N_4088,N_4089,N_4090,N_4091,N_4092,N_4096,N_4097,N_4098,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4117,N_4118,N_4119,N_4120,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4131,N_4132,N_4133,N_4135,N_4136,N_4139,N_4140,N_4142,N_4144,N_4145,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4155,N_4157,N_4158,N_4161,N_4162,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4182,N_4184,N_4185,N_4187,N_4188,N_4190,N_4191,N_4192,N_4193,N_4194,N_4197,N_4198,N_4199,N_4200,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4262,N_4263,N_4264,N_4265,N_4266,N_4268,N_4269,N_4270,N_4271,N_4273,N_4274,N_4275,N_4276,N_4278,N_4279,N_4280,N_4282,N_4284,N_4285,N_4286,N_4288,N_4289,N_4290,N_4291,N_4293,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4306,N_4307,N_4308,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4321,N_4323,N_4325,N_4326,N_4328,N_4329,N_4330,N_4331,N_4333,N_4334,N_4335,N_4336,N_4338,N_4339,N_4340,N_4343,N_4347,N_4348,N_4349,N_4351,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4361,N_4362,N_4363,N_4364,N_4365,N_4367,N_4368,N_4369,N_4372,N_4373,N_4375,N_4377,N_4378,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4412,N_4413,N_4414,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4425,N_4426,N_4427,N_4428,N_4429,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4456,N_4457,N_4458,N_4459,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4483,N_4484,N_4485,N_4486,N_4487,N_4489,N_4490,N_4491,N_4492,N_4493,N_4495,N_4496,N_4498,N_4499,N_4500,N_4502,N_4503,N_4505,N_4507,N_4508,N_4510,N_4513,N_4515,N_4517,N_4518,N_4519,N_4520,N_4522,N_4523,N_4524,N_4525,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4570,N_4572,N_4573,N_4574,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4584,N_4585,N_4586,N_4587,N_4589,N_4590,N_4593,N_4596,N_4597,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4608,N_4609,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4629,N_4632,N_4633,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4665,N_4666,N_4667,N_4668,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4679,N_4680,N_4681,N_4684,N_4685,N_4686,N_4688,N_4689,N_4690,N_4691,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4701,N_4703,N_4705,N_4706,N_4707,N_4708,N_4709,N_4711,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4721,N_4722,N_4723,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4756,N_4758,N_4759,N_4760,N_4761,N_4762,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4785,N_4787,N_4788,N_4789,N_4791,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4823,N_4824,N_4827,N_4828,N_4829,N_4830,N_4833,N_4834,N_4835,N_4836,N_4839,N_4840,N_4841,N_4843,N_4844,N_4845,N_4846,N_4848,N_4850,N_4851,N_4852,N_4853,N_4855,N_4856,N_4857,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4866,N_4867,N_4868,N_4870,N_4871,N_4872,N_4874,N_4875,N_4876,N_4877,N_4878,N_4880,N_4881,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4890,N_4891,N_4892,N_4894,N_4896,N_4898,N_4899,N_4900,N_4902,N_4903,N_4905,N_4906,N_4907,N_4909,N_4910,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4939,N_4940,N_4942,N_4943,N_4944,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4967,N_4968,N_4970,N_4972,N_4973,N_4975,N_4976,N_4980,N_4982,N_4983,N_4984,N_4987,N_4988,N_4989,N_4990,N_4992,N_4993,N_4994,N_4995,N_4996,N_4998,N_4999;
or U0 (N_0,In_346,In_538);
and U1 (N_1,In_411,In_22);
or U2 (N_2,In_200,In_603);
and U3 (N_3,In_686,In_67);
nor U4 (N_4,In_627,In_334);
and U5 (N_5,In_460,In_720);
and U6 (N_6,In_501,In_746);
nor U7 (N_7,In_278,In_144);
or U8 (N_8,In_10,In_436);
and U9 (N_9,In_288,In_254);
nor U10 (N_10,In_240,In_407);
nand U11 (N_11,In_111,In_551);
nand U12 (N_12,In_170,In_96);
nand U13 (N_13,In_54,In_262);
and U14 (N_14,In_721,In_675);
nand U15 (N_15,In_374,In_238);
nor U16 (N_16,In_12,In_119);
nor U17 (N_17,In_402,In_21);
nand U18 (N_18,In_671,In_504);
nand U19 (N_19,In_483,In_745);
or U20 (N_20,In_716,In_13);
nor U21 (N_21,In_398,In_228);
nor U22 (N_22,In_148,In_279);
nand U23 (N_23,In_340,In_133);
or U24 (N_24,In_500,In_71);
and U25 (N_25,In_48,In_49);
nor U26 (N_26,In_308,In_134);
or U27 (N_27,In_364,In_492);
nand U28 (N_28,In_257,In_25);
and U29 (N_29,In_422,In_469);
nand U30 (N_30,In_92,In_568);
and U31 (N_31,In_673,In_314);
and U32 (N_32,In_418,In_56);
nor U33 (N_33,In_624,In_209);
nand U34 (N_34,In_327,In_302);
nor U35 (N_35,In_408,In_130);
and U36 (N_36,In_516,In_517);
nand U37 (N_37,In_737,In_511);
and U38 (N_38,In_616,In_692);
nand U39 (N_39,In_174,In_585);
nand U40 (N_40,In_309,In_345);
or U41 (N_41,In_728,In_747);
nor U42 (N_42,In_506,In_732);
or U43 (N_43,In_566,In_105);
or U44 (N_44,In_444,In_385);
or U45 (N_45,In_175,In_1);
or U46 (N_46,In_318,In_575);
or U47 (N_47,In_199,In_196);
nor U48 (N_48,In_290,In_547);
or U49 (N_49,In_740,In_331);
or U50 (N_50,In_699,In_635);
and U51 (N_51,In_555,In_68);
xor U52 (N_52,In_378,In_696);
or U53 (N_53,In_285,In_493);
nor U54 (N_54,In_706,In_355);
and U55 (N_55,In_125,In_61);
or U56 (N_56,In_214,In_729);
or U57 (N_57,In_232,In_390);
and U58 (N_58,In_410,In_412);
or U59 (N_59,In_625,In_584);
nor U60 (N_60,In_578,In_190);
nand U61 (N_61,In_74,In_252);
or U62 (N_62,In_428,In_362);
or U63 (N_63,In_221,In_234);
nand U64 (N_64,In_678,In_642);
or U65 (N_65,In_265,In_649);
nand U66 (N_66,In_354,In_167);
nor U67 (N_67,In_156,In_27);
nor U68 (N_68,In_51,In_689);
nor U69 (N_69,In_574,In_672);
and U70 (N_70,In_179,In_690);
or U71 (N_71,In_187,In_205);
nor U72 (N_72,In_631,In_427);
nor U73 (N_73,In_136,In_352);
nand U74 (N_74,In_650,In_58);
nor U75 (N_75,In_186,In_475);
nor U76 (N_76,In_425,In_465);
or U77 (N_77,In_90,In_739);
nand U78 (N_78,In_694,In_734);
nand U79 (N_79,In_305,In_363);
or U80 (N_80,In_225,In_332);
nand U81 (N_81,In_736,In_23);
or U82 (N_82,In_315,In_297);
or U83 (N_83,In_473,In_623);
nor U84 (N_84,In_260,In_135);
or U85 (N_85,In_264,In_556);
nand U86 (N_86,In_645,In_705);
nor U87 (N_87,In_541,In_487);
and U88 (N_88,In_558,In_122);
nor U89 (N_89,In_20,In_535);
nand U90 (N_90,In_89,In_204);
or U91 (N_91,In_521,In_701);
nand U92 (N_92,In_409,In_477);
or U93 (N_93,In_66,In_165);
nand U94 (N_94,In_415,In_19);
nor U95 (N_95,In_271,In_69);
or U96 (N_96,In_294,In_459);
nor U97 (N_97,In_661,In_283);
nor U98 (N_98,In_383,In_490);
nand U99 (N_99,In_185,In_7);
and U100 (N_100,In_582,In_321);
and U101 (N_101,In_524,In_162);
or U102 (N_102,In_651,In_78);
nand U103 (N_103,In_46,In_31);
xnor U104 (N_104,In_680,In_674);
and U105 (N_105,In_550,In_534);
or U106 (N_106,In_79,In_152);
or U107 (N_107,In_608,In_195);
nand U108 (N_108,In_607,In_405);
nand U109 (N_109,In_344,In_273);
and U110 (N_110,In_284,In_268);
or U111 (N_111,In_660,In_348);
or U112 (N_112,In_280,In_276);
nor U113 (N_113,In_508,In_60);
nor U114 (N_114,In_634,In_420);
or U115 (N_115,In_569,In_256);
nand U116 (N_116,In_206,In_394);
or U117 (N_117,In_494,In_65);
and U118 (N_118,In_289,In_724);
nand U119 (N_119,In_733,In_57);
xor U120 (N_120,In_401,In_178);
xnor U121 (N_121,In_502,In_188);
nor U122 (N_122,In_522,In_684);
or U123 (N_123,In_472,In_639);
and U124 (N_124,In_24,In_382);
xor U125 (N_125,In_208,In_147);
or U126 (N_126,In_29,In_338);
nand U127 (N_127,In_589,In_527);
and U128 (N_128,In_41,In_384);
or U129 (N_129,In_266,In_143);
or U130 (N_130,In_386,In_37);
nand U131 (N_131,In_326,In_5);
and U132 (N_132,In_261,In_463);
or U133 (N_133,In_579,In_180);
nand U134 (N_134,In_498,In_738);
and U135 (N_135,In_381,In_154);
or U136 (N_136,In_59,In_670);
and U137 (N_137,In_668,In_72);
nand U138 (N_138,In_351,In_718);
xnor U139 (N_139,In_219,In_104);
and U140 (N_140,In_621,In_210);
nor U141 (N_141,In_269,In_536);
and U142 (N_142,In_543,In_388);
or U143 (N_143,In_115,In_513);
nand U144 (N_144,In_400,In_447);
nor U145 (N_145,In_212,In_18);
xor U146 (N_146,In_38,In_549);
nor U147 (N_147,In_368,In_662);
and U148 (N_148,In_141,In_140);
and U149 (N_149,In_499,In_617);
xor U150 (N_150,In_138,In_395);
nor U151 (N_151,In_11,In_638);
nor U152 (N_152,In_528,In_697);
nor U153 (N_153,In_433,In_613);
xnor U154 (N_154,In_466,In_570);
or U155 (N_155,In_202,In_726);
xnor U156 (N_156,In_274,In_588);
nand U157 (N_157,In_600,In_544);
xnor U158 (N_158,In_198,In_430);
nor U159 (N_159,In_479,In_343);
nand U160 (N_160,In_328,In_80);
and U161 (N_161,In_424,In_110);
nand U162 (N_162,In_630,In_158);
and U163 (N_163,In_137,In_665);
nand U164 (N_164,In_667,In_453);
and U165 (N_165,In_310,In_723);
or U166 (N_166,In_648,In_376);
and U167 (N_167,In_486,In_223);
nand U168 (N_168,In_192,In_215);
nor U169 (N_169,In_677,In_583);
nand U170 (N_170,In_127,In_275);
and U171 (N_171,In_611,In_529);
and U172 (N_172,In_519,In_231);
or U173 (N_173,In_207,In_380);
xor U174 (N_174,In_34,In_282);
or U175 (N_175,In_299,In_197);
nor U176 (N_176,In_698,In_748);
nand U177 (N_177,In_581,In_357);
and U178 (N_178,In_693,In_461);
nor U179 (N_179,In_391,In_614);
nor U180 (N_180,In_358,In_171);
and U181 (N_181,In_485,In_303);
or U182 (N_182,In_471,In_622);
nand U183 (N_183,In_683,In_572);
and U184 (N_184,In_731,In_30);
xnor U185 (N_185,In_604,In_476);
or U186 (N_186,In_416,In_478);
or U187 (N_187,In_539,In_191);
or U188 (N_188,In_177,In_116);
or U189 (N_189,In_591,In_619);
or U190 (N_190,In_244,In_17);
and U191 (N_191,In_176,In_403);
and U192 (N_192,In_55,In_586);
nor U193 (N_193,In_373,In_250);
or U194 (N_194,In_40,In_301);
nor U195 (N_195,In_560,In_628);
or U196 (N_196,In_15,In_632);
or U197 (N_197,In_329,In_421);
nor U198 (N_198,In_107,In_270);
nor U199 (N_199,In_230,In_546);
and U200 (N_200,In_82,In_322);
and U201 (N_201,In_666,In_711);
or U202 (N_202,In_319,In_335);
nand U203 (N_203,In_452,In_263);
nor U204 (N_204,In_679,In_458);
nor U205 (N_205,In_552,In_169);
nor U206 (N_206,In_446,In_236);
nand U207 (N_207,In_599,In_742);
or U208 (N_208,In_341,In_474);
and U209 (N_209,In_641,In_510);
or U210 (N_210,In_372,In_296);
and U211 (N_211,In_682,In_640);
nor U212 (N_212,In_99,In_160);
nor U213 (N_213,In_128,In_593);
nor U214 (N_214,In_35,In_377);
nand U215 (N_215,In_168,In_150);
and U216 (N_216,In_562,In_157);
and U217 (N_217,In_676,In_153);
nand U218 (N_218,In_43,In_533);
and U219 (N_219,In_507,In_126);
nand U220 (N_220,In_488,In_653);
nand U221 (N_221,In_610,In_658);
nand U222 (N_222,In_577,In_468);
nor U223 (N_223,In_730,In_243);
and U224 (N_224,In_311,In_565);
or U225 (N_225,In_183,In_129);
or U226 (N_226,In_464,In_235);
nand U227 (N_227,In_323,In_531);
or U228 (N_228,In_456,In_505);
nor U229 (N_229,In_28,In_307);
and U230 (N_230,In_455,In_744);
and U231 (N_231,In_443,In_434);
and U232 (N_232,In_325,In_44);
nor U233 (N_233,In_218,In_497);
and U234 (N_234,In_489,In_451);
nand U235 (N_235,In_573,In_559);
and U236 (N_236,In_248,In_664);
nand U237 (N_237,In_304,In_596);
or U238 (N_238,In_467,In_655);
nand U239 (N_239,In_159,In_606);
or U240 (N_240,In_749,In_438);
or U241 (N_241,In_389,In_164);
nand U242 (N_242,In_100,In_480);
xor U243 (N_243,In_712,In_93);
and U244 (N_244,In_495,In_114);
nand U245 (N_245,In_542,In_435);
or U246 (N_246,In_6,In_298);
and U247 (N_247,In_42,In_633);
nor U248 (N_248,In_367,In_347);
nor U249 (N_249,In_448,In_342);
nand U250 (N_250,In_330,In_520);
nor U251 (N_251,In_609,In_417);
nor U252 (N_252,In_484,In_124);
nand U253 (N_253,In_636,In_226);
or U254 (N_254,In_91,In_481);
or U255 (N_255,In_85,In_349);
nor U256 (N_256,In_602,In_258);
nor U257 (N_257,In_76,In_594);
nor U258 (N_258,In_439,In_312);
nand U259 (N_259,In_47,In_687);
or U260 (N_260,In_454,In_605);
xor U261 (N_261,In_652,In_702);
nor U262 (N_262,In_576,In_654);
and U263 (N_263,In_442,In_317);
nand U264 (N_264,In_426,In_84);
and U265 (N_265,In_445,In_36);
or U266 (N_266,In_216,In_53);
nor U267 (N_267,In_695,In_580);
nand U268 (N_268,In_399,In_688);
nand U269 (N_269,In_371,In_103);
nor U270 (N_270,In_437,In_518);
and U271 (N_271,In_450,In_87);
or U272 (N_272,In_704,In_503);
or U273 (N_273,In_45,In_626);
or U274 (N_274,In_429,In_73);
and U275 (N_275,In_194,In_714);
or U276 (N_276,In_548,In_201);
and U277 (N_277,In_155,In_8);
nor U278 (N_278,In_470,In_710);
nor U279 (N_279,In_392,In_142);
and U280 (N_280,In_404,In_166);
nor U281 (N_281,In_64,In_118);
xor U282 (N_282,In_722,In_184);
nand U283 (N_283,In_253,In_112);
and U284 (N_284,In_557,In_77);
and U285 (N_285,In_9,In_245);
or U286 (N_286,In_540,In_239);
nor U287 (N_287,In_163,In_300);
and U288 (N_288,In_644,In_211);
nand U289 (N_289,In_643,In_669);
and U290 (N_290,In_16,In_735);
or U291 (N_291,In_63,In_587);
nand U292 (N_292,In_172,In_715);
and U293 (N_293,In_379,In_365);
or U294 (N_294,In_2,In_316);
nand U295 (N_295,In_95,In_14);
nand U296 (N_296,In_32,In_241);
nand U297 (N_297,In_512,In_646);
nand U298 (N_298,In_393,In_595);
and U299 (N_299,In_707,In_217);
or U300 (N_300,In_597,In_4);
and U301 (N_301,In_491,In_62);
nand U302 (N_302,In_33,In_656);
nor U303 (N_303,In_413,In_281);
or U304 (N_304,In_295,In_532);
and U305 (N_305,In_590,In_182);
and U306 (N_306,In_0,In_359);
and U307 (N_307,In_743,In_369);
and U308 (N_308,In_242,In_131);
or U309 (N_309,In_109,In_75);
nand U310 (N_310,In_313,In_292);
nand U311 (N_311,In_237,In_106);
and U312 (N_312,In_691,In_336);
nand U313 (N_313,In_681,In_139);
and U314 (N_314,In_108,In_146);
nand U315 (N_315,In_286,In_523);
nor U316 (N_316,In_3,In_181);
or U317 (N_317,In_50,In_515);
nor U318 (N_318,In_375,In_618);
nor U319 (N_319,In_440,In_366);
and U320 (N_320,In_509,In_123);
nand U321 (N_321,In_397,In_102);
nor U322 (N_322,In_685,In_419);
nand U323 (N_323,In_350,In_339);
or U324 (N_324,In_637,In_620);
or U325 (N_325,In_26,In_612);
or U326 (N_326,In_259,In_423);
nor U327 (N_327,In_229,In_189);
nand U328 (N_328,In_414,In_370);
or U329 (N_329,In_81,In_249);
or U330 (N_330,In_709,In_277);
or U331 (N_331,In_121,In_615);
nor U332 (N_332,In_396,In_554);
nand U333 (N_333,In_233,In_117);
nor U334 (N_334,In_657,In_406);
or U335 (N_335,In_324,In_120);
and U336 (N_336,In_39,In_545);
or U337 (N_337,In_203,In_88);
or U338 (N_338,In_741,In_251);
nor U339 (N_339,In_224,In_561);
nand U340 (N_340,In_52,In_291);
xor U341 (N_341,In_213,In_601);
nand U342 (N_342,In_659,In_449);
or U343 (N_343,In_113,In_227);
nor U344 (N_344,In_94,In_629);
nand U345 (N_345,In_86,In_432);
nor U346 (N_346,In_525,In_145);
and U347 (N_347,In_306,In_173);
or U348 (N_348,In_703,In_387);
and U349 (N_349,In_567,In_287);
and U350 (N_350,In_530,In_149);
or U351 (N_351,In_132,In_222);
nand U352 (N_352,In_663,In_272);
and U353 (N_353,In_293,In_647);
and U354 (N_354,In_247,In_514);
or U355 (N_355,In_267,In_246);
nor U356 (N_356,In_151,In_337);
and U357 (N_357,In_431,In_725);
nor U358 (N_358,In_161,In_563);
xnor U359 (N_359,In_361,In_441);
or U360 (N_360,In_193,In_571);
or U361 (N_361,In_462,In_70);
nand U362 (N_362,In_255,In_598);
and U363 (N_363,In_320,In_98);
or U364 (N_364,In_97,In_564);
nor U365 (N_365,In_360,In_496);
and U366 (N_366,In_457,In_719);
and U367 (N_367,In_537,In_708);
and U368 (N_368,In_717,In_101);
nand U369 (N_369,In_713,In_353);
or U370 (N_370,In_356,In_727);
or U371 (N_371,In_220,In_83);
and U372 (N_372,In_526,In_700);
nand U373 (N_373,In_482,In_553);
and U374 (N_374,In_333,In_592);
nor U375 (N_375,In_667,In_57);
or U376 (N_376,In_715,In_601);
nor U377 (N_377,In_211,In_468);
and U378 (N_378,In_628,In_575);
nand U379 (N_379,In_18,In_644);
nand U380 (N_380,In_105,In_292);
and U381 (N_381,In_338,In_509);
nor U382 (N_382,In_436,In_158);
and U383 (N_383,In_186,In_579);
nor U384 (N_384,In_709,In_121);
and U385 (N_385,In_79,In_469);
nor U386 (N_386,In_624,In_120);
nand U387 (N_387,In_377,In_265);
and U388 (N_388,In_508,In_494);
nor U389 (N_389,In_289,In_211);
or U390 (N_390,In_114,In_669);
nor U391 (N_391,In_741,In_733);
nor U392 (N_392,In_316,In_430);
nand U393 (N_393,In_440,In_363);
nor U394 (N_394,In_613,In_587);
nor U395 (N_395,In_481,In_163);
and U396 (N_396,In_256,In_655);
and U397 (N_397,In_626,In_128);
or U398 (N_398,In_110,In_676);
or U399 (N_399,In_575,In_21);
nor U400 (N_400,In_549,In_70);
nor U401 (N_401,In_592,In_718);
or U402 (N_402,In_92,In_598);
nand U403 (N_403,In_740,In_546);
nor U404 (N_404,In_288,In_26);
and U405 (N_405,In_351,In_467);
or U406 (N_406,In_170,In_40);
and U407 (N_407,In_359,In_315);
and U408 (N_408,In_587,In_74);
nor U409 (N_409,In_247,In_36);
and U410 (N_410,In_356,In_245);
and U411 (N_411,In_436,In_525);
nor U412 (N_412,In_365,In_465);
nor U413 (N_413,In_15,In_77);
or U414 (N_414,In_693,In_714);
nand U415 (N_415,In_681,In_477);
nand U416 (N_416,In_16,In_602);
nor U417 (N_417,In_326,In_746);
or U418 (N_418,In_514,In_398);
and U419 (N_419,In_286,In_310);
nor U420 (N_420,In_211,In_467);
or U421 (N_421,In_301,In_468);
or U422 (N_422,In_596,In_269);
nor U423 (N_423,In_682,In_97);
xnor U424 (N_424,In_573,In_367);
xnor U425 (N_425,In_239,In_686);
or U426 (N_426,In_634,In_560);
nor U427 (N_427,In_566,In_378);
and U428 (N_428,In_440,In_376);
and U429 (N_429,In_65,In_531);
and U430 (N_430,In_148,In_694);
and U431 (N_431,In_90,In_490);
nor U432 (N_432,In_70,In_546);
xnor U433 (N_433,In_197,In_255);
nand U434 (N_434,In_150,In_82);
and U435 (N_435,In_242,In_573);
nand U436 (N_436,In_305,In_472);
or U437 (N_437,In_404,In_251);
or U438 (N_438,In_62,In_53);
nor U439 (N_439,In_272,In_25);
or U440 (N_440,In_388,In_277);
and U441 (N_441,In_576,In_53);
and U442 (N_442,In_525,In_486);
nand U443 (N_443,In_266,In_547);
nand U444 (N_444,In_393,In_310);
and U445 (N_445,In_380,In_690);
nand U446 (N_446,In_253,In_665);
and U447 (N_447,In_423,In_530);
nor U448 (N_448,In_341,In_330);
and U449 (N_449,In_127,In_391);
nand U450 (N_450,In_506,In_428);
nor U451 (N_451,In_32,In_104);
nor U452 (N_452,In_318,In_179);
nand U453 (N_453,In_695,In_445);
or U454 (N_454,In_21,In_364);
and U455 (N_455,In_239,In_743);
or U456 (N_456,In_80,In_239);
nor U457 (N_457,In_685,In_516);
and U458 (N_458,In_222,In_282);
or U459 (N_459,In_590,In_199);
and U460 (N_460,In_467,In_13);
or U461 (N_461,In_560,In_350);
or U462 (N_462,In_378,In_510);
and U463 (N_463,In_494,In_362);
and U464 (N_464,In_176,In_211);
nor U465 (N_465,In_431,In_620);
and U466 (N_466,In_342,In_336);
nor U467 (N_467,In_613,In_328);
nand U468 (N_468,In_505,In_497);
or U469 (N_469,In_686,In_623);
and U470 (N_470,In_162,In_708);
nor U471 (N_471,In_484,In_305);
or U472 (N_472,In_557,In_710);
nand U473 (N_473,In_137,In_535);
nor U474 (N_474,In_278,In_69);
nand U475 (N_475,In_540,In_464);
nor U476 (N_476,In_518,In_20);
nor U477 (N_477,In_515,In_686);
or U478 (N_478,In_688,In_530);
and U479 (N_479,In_278,In_1);
and U480 (N_480,In_627,In_282);
nor U481 (N_481,In_107,In_157);
or U482 (N_482,In_487,In_174);
nand U483 (N_483,In_263,In_41);
and U484 (N_484,In_379,In_422);
and U485 (N_485,In_709,In_268);
nand U486 (N_486,In_363,In_554);
nand U487 (N_487,In_266,In_259);
nor U488 (N_488,In_62,In_604);
and U489 (N_489,In_600,In_42);
nand U490 (N_490,In_275,In_227);
or U491 (N_491,In_110,In_445);
nor U492 (N_492,In_560,In_404);
and U493 (N_493,In_173,In_482);
nor U494 (N_494,In_73,In_563);
and U495 (N_495,In_615,In_427);
or U496 (N_496,In_319,In_736);
nor U497 (N_497,In_578,In_650);
and U498 (N_498,In_339,In_630);
nor U499 (N_499,In_691,In_377);
nor U500 (N_500,In_213,In_707);
and U501 (N_501,In_606,In_329);
or U502 (N_502,In_208,In_5);
or U503 (N_503,In_142,In_695);
or U504 (N_504,In_97,In_40);
nand U505 (N_505,In_163,In_155);
nor U506 (N_506,In_477,In_351);
and U507 (N_507,In_549,In_445);
or U508 (N_508,In_39,In_644);
nand U509 (N_509,In_547,In_137);
or U510 (N_510,In_104,In_210);
and U511 (N_511,In_129,In_421);
and U512 (N_512,In_331,In_82);
nor U513 (N_513,In_459,In_119);
and U514 (N_514,In_415,In_613);
nand U515 (N_515,In_594,In_545);
or U516 (N_516,In_81,In_176);
and U517 (N_517,In_623,In_721);
nand U518 (N_518,In_600,In_449);
nand U519 (N_519,In_497,In_236);
nand U520 (N_520,In_253,In_370);
and U521 (N_521,In_473,In_615);
nor U522 (N_522,In_722,In_58);
nor U523 (N_523,In_263,In_369);
nand U524 (N_524,In_531,In_686);
nor U525 (N_525,In_283,In_717);
or U526 (N_526,In_100,In_593);
or U527 (N_527,In_473,In_175);
or U528 (N_528,In_711,In_718);
nor U529 (N_529,In_140,In_210);
or U530 (N_530,In_411,In_637);
nor U531 (N_531,In_533,In_52);
and U532 (N_532,In_232,In_524);
nand U533 (N_533,In_103,In_514);
and U534 (N_534,In_508,In_305);
or U535 (N_535,In_561,In_325);
or U536 (N_536,In_158,In_423);
or U537 (N_537,In_289,In_216);
and U538 (N_538,In_138,In_467);
nand U539 (N_539,In_318,In_344);
nand U540 (N_540,In_608,In_419);
and U541 (N_541,In_398,In_436);
or U542 (N_542,In_355,In_218);
nor U543 (N_543,In_390,In_60);
nand U544 (N_544,In_536,In_430);
and U545 (N_545,In_23,In_33);
or U546 (N_546,In_703,In_338);
and U547 (N_547,In_512,In_143);
and U548 (N_548,In_600,In_327);
or U549 (N_549,In_718,In_168);
nor U550 (N_550,In_422,In_462);
and U551 (N_551,In_533,In_506);
or U552 (N_552,In_255,In_701);
nand U553 (N_553,In_445,In_442);
nand U554 (N_554,In_399,In_230);
or U555 (N_555,In_59,In_56);
and U556 (N_556,In_508,In_27);
or U557 (N_557,In_264,In_114);
nand U558 (N_558,In_4,In_235);
or U559 (N_559,In_458,In_421);
nor U560 (N_560,In_217,In_698);
xnor U561 (N_561,In_273,In_696);
or U562 (N_562,In_465,In_726);
or U563 (N_563,In_412,In_223);
nor U564 (N_564,In_507,In_138);
and U565 (N_565,In_554,In_725);
and U566 (N_566,In_238,In_619);
xor U567 (N_567,In_543,In_76);
nand U568 (N_568,In_524,In_194);
nand U569 (N_569,In_709,In_678);
nor U570 (N_570,In_53,In_141);
and U571 (N_571,In_577,In_256);
and U572 (N_572,In_65,In_122);
and U573 (N_573,In_451,In_343);
and U574 (N_574,In_678,In_686);
and U575 (N_575,In_336,In_411);
nand U576 (N_576,In_455,In_454);
or U577 (N_577,In_242,In_727);
xor U578 (N_578,In_216,In_183);
or U579 (N_579,In_684,In_664);
or U580 (N_580,In_616,In_351);
nor U581 (N_581,In_320,In_66);
nor U582 (N_582,In_51,In_561);
and U583 (N_583,In_545,In_423);
or U584 (N_584,In_140,In_177);
nor U585 (N_585,In_360,In_268);
nand U586 (N_586,In_671,In_383);
nand U587 (N_587,In_513,In_480);
or U588 (N_588,In_149,In_264);
nor U589 (N_589,In_681,In_514);
and U590 (N_590,In_415,In_434);
nor U591 (N_591,In_357,In_346);
and U592 (N_592,In_610,In_228);
nor U593 (N_593,In_649,In_298);
and U594 (N_594,In_622,In_112);
and U595 (N_595,In_293,In_81);
and U596 (N_596,In_373,In_451);
and U597 (N_597,In_539,In_44);
or U598 (N_598,In_393,In_489);
nor U599 (N_599,In_465,In_479);
or U600 (N_600,In_138,In_50);
xnor U601 (N_601,In_730,In_384);
nand U602 (N_602,In_43,In_329);
and U603 (N_603,In_220,In_666);
and U604 (N_604,In_278,In_385);
nor U605 (N_605,In_541,In_338);
and U606 (N_606,In_534,In_394);
or U607 (N_607,In_194,In_473);
or U608 (N_608,In_223,In_334);
nand U609 (N_609,In_387,In_561);
or U610 (N_610,In_597,In_648);
and U611 (N_611,In_201,In_16);
and U612 (N_612,In_297,In_350);
nor U613 (N_613,In_287,In_506);
nand U614 (N_614,In_749,In_375);
and U615 (N_615,In_61,In_414);
nand U616 (N_616,In_327,In_52);
nor U617 (N_617,In_227,In_450);
nor U618 (N_618,In_92,In_384);
and U619 (N_619,In_675,In_221);
nor U620 (N_620,In_21,In_211);
or U621 (N_621,In_254,In_389);
nor U622 (N_622,In_576,In_572);
or U623 (N_623,In_297,In_419);
and U624 (N_624,In_443,In_255);
and U625 (N_625,In_183,In_109);
xnor U626 (N_626,In_157,In_193);
or U627 (N_627,In_60,In_79);
nor U628 (N_628,In_3,In_225);
nand U629 (N_629,In_389,In_535);
nand U630 (N_630,In_509,In_70);
nor U631 (N_631,In_599,In_61);
and U632 (N_632,In_255,In_397);
nand U633 (N_633,In_249,In_571);
nor U634 (N_634,In_373,In_73);
nand U635 (N_635,In_317,In_666);
nor U636 (N_636,In_42,In_738);
nor U637 (N_637,In_195,In_69);
and U638 (N_638,In_74,In_621);
or U639 (N_639,In_404,In_402);
and U640 (N_640,In_696,In_408);
nor U641 (N_641,In_633,In_333);
nand U642 (N_642,In_724,In_708);
nor U643 (N_643,In_590,In_286);
or U644 (N_644,In_439,In_247);
nor U645 (N_645,In_503,In_558);
and U646 (N_646,In_329,In_218);
or U647 (N_647,In_112,In_744);
or U648 (N_648,In_39,In_641);
or U649 (N_649,In_149,In_200);
nor U650 (N_650,In_506,In_36);
and U651 (N_651,In_1,In_622);
or U652 (N_652,In_491,In_449);
or U653 (N_653,In_165,In_422);
nand U654 (N_654,In_107,In_196);
and U655 (N_655,In_400,In_340);
nand U656 (N_656,In_120,In_735);
nor U657 (N_657,In_464,In_0);
nor U658 (N_658,In_374,In_541);
nor U659 (N_659,In_733,In_430);
nor U660 (N_660,In_4,In_51);
or U661 (N_661,In_136,In_369);
xor U662 (N_662,In_74,In_168);
xnor U663 (N_663,In_423,In_745);
nand U664 (N_664,In_201,In_369);
nor U665 (N_665,In_694,In_591);
xnor U666 (N_666,In_235,In_383);
or U667 (N_667,In_705,In_629);
nand U668 (N_668,In_94,In_585);
nand U669 (N_669,In_215,In_442);
nor U670 (N_670,In_552,In_621);
nand U671 (N_671,In_572,In_660);
or U672 (N_672,In_309,In_372);
nand U673 (N_673,In_57,In_444);
or U674 (N_674,In_373,In_139);
and U675 (N_675,In_492,In_148);
nand U676 (N_676,In_402,In_582);
and U677 (N_677,In_123,In_413);
nand U678 (N_678,In_276,In_139);
or U679 (N_679,In_483,In_559);
xnor U680 (N_680,In_257,In_150);
nand U681 (N_681,In_640,In_126);
or U682 (N_682,In_184,In_671);
nor U683 (N_683,In_542,In_23);
nor U684 (N_684,In_252,In_250);
xnor U685 (N_685,In_586,In_704);
nor U686 (N_686,In_24,In_445);
and U687 (N_687,In_102,In_431);
nand U688 (N_688,In_71,In_597);
nor U689 (N_689,In_610,In_376);
or U690 (N_690,In_168,In_586);
nor U691 (N_691,In_101,In_325);
nor U692 (N_692,In_342,In_739);
and U693 (N_693,In_97,In_649);
nand U694 (N_694,In_727,In_422);
and U695 (N_695,In_26,In_335);
and U696 (N_696,In_59,In_107);
or U697 (N_697,In_116,In_647);
xor U698 (N_698,In_322,In_652);
and U699 (N_699,In_35,In_220);
nor U700 (N_700,In_204,In_685);
nand U701 (N_701,In_645,In_67);
or U702 (N_702,In_675,In_107);
or U703 (N_703,In_195,In_544);
and U704 (N_704,In_550,In_294);
and U705 (N_705,In_312,In_86);
nor U706 (N_706,In_378,In_38);
and U707 (N_707,In_700,In_132);
and U708 (N_708,In_32,In_459);
and U709 (N_709,In_190,In_410);
nand U710 (N_710,In_681,In_491);
or U711 (N_711,In_702,In_409);
nor U712 (N_712,In_2,In_156);
nor U713 (N_713,In_380,In_652);
or U714 (N_714,In_618,In_257);
or U715 (N_715,In_498,In_504);
nor U716 (N_716,In_680,In_501);
nor U717 (N_717,In_84,In_526);
and U718 (N_718,In_90,In_374);
and U719 (N_719,In_417,In_201);
or U720 (N_720,In_287,In_491);
and U721 (N_721,In_615,In_88);
nand U722 (N_722,In_649,In_611);
nor U723 (N_723,In_224,In_661);
or U724 (N_724,In_467,In_698);
and U725 (N_725,In_186,In_104);
or U726 (N_726,In_706,In_418);
nand U727 (N_727,In_739,In_568);
or U728 (N_728,In_559,In_157);
and U729 (N_729,In_669,In_745);
or U730 (N_730,In_396,In_395);
nand U731 (N_731,In_449,In_516);
nor U732 (N_732,In_613,In_607);
nand U733 (N_733,In_217,In_378);
and U734 (N_734,In_515,In_185);
nor U735 (N_735,In_288,In_340);
and U736 (N_736,In_633,In_168);
and U737 (N_737,In_579,In_630);
or U738 (N_738,In_421,In_37);
nand U739 (N_739,In_70,In_280);
and U740 (N_740,In_484,In_684);
nor U741 (N_741,In_617,In_610);
nor U742 (N_742,In_720,In_17);
and U743 (N_743,In_393,In_311);
nor U744 (N_744,In_535,In_560);
nand U745 (N_745,In_618,In_498);
and U746 (N_746,In_568,In_588);
xor U747 (N_747,In_262,In_424);
nand U748 (N_748,In_596,In_40);
and U749 (N_749,In_584,In_259);
and U750 (N_750,In_109,In_219);
and U751 (N_751,In_631,In_340);
or U752 (N_752,In_670,In_77);
nand U753 (N_753,In_91,In_56);
xnor U754 (N_754,In_598,In_317);
nand U755 (N_755,In_532,In_259);
or U756 (N_756,In_527,In_58);
and U757 (N_757,In_684,In_351);
nand U758 (N_758,In_367,In_64);
and U759 (N_759,In_89,In_436);
nand U760 (N_760,In_639,In_341);
nand U761 (N_761,In_36,In_404);
or U762 (N_762,In_120,In_599);
and U763 (N_763,In_630,In_230);
or U764 (N_764,In_258,In_346);
or U765 (N_765,In_722,In_386);
nand U766 (N_766,In_392,In_40);
nor U767 (N_767,In_131,In_352);
nand U768 (N_768,In_702,In_631);
nand U769 (N_769,In_167,In_61);
and U770 (N_770,In_632,In_82);
nor U771 (N_771,In_376,In_122);
and U772 (N_772,In_15,In_112);
nor U773 (N_773,In_269,In_185);
nand U774 (N_774,In_60,In_274);
nor U775 (N_775,In_420,In_319);
nor U776 (N_776,In_689,In_306);
nor U777 (N_777,In_55,In_385);
nand U778 (N_778,In_250,In_444);
nand U779 (N_779,In_434,In_564);
and U780 (N_780,In_715,In_304);
or U781 (N_781,In_189,In_719);
nand U782 (N_782,In_736,In_440);
nand U783 (N_783,In_36,In_150);
nor U784 (N_784,In_81,In_252);
and U785 (N_785,In_244,In_664);
nor U786 (N_786,In_565,In_339);
xnor U787 (N_787,In_651,In_428);
nor U788 (N_788,In_143,In_431);
and U789 (N_789,In_512,In_626);
nand U790 (N_790,In_472,In_46);
or U791 (N_791,In_529,In_235);
or U792 (N_792,In_119,In_723);
nor U793 (N_793,In_225,In_731);
and U794 (N_794,In_51,In_542);
nor U795 (N_795,In_617,In_336);
nor U796 (N_796,In_244,In_438);
nor U797 (N_797,In_275,In_104);
or U798 (N_798,In_712,In_172);
nand U799 (N_799,In_598,In_578);
nand U800 (N_800,In_506,In_100);
nand U801 (N_801,In_244,In_594);
nor U802 (N_802,In_275,In_612);
and U803 (N_803,In_537,In_682);
and U804 (N_804,In_486,In_207);
nor U805 (N_805,In_98,In_458);
nand U806 (N_806,In_499,In_51);
or U807 (N_807,In_610,In_708);
and U808 (N_808,In_719,In_81);
nor U809 (N_809,In_64,In_127);
and U810 (N_810,In_601,In_177);
and U811 (N_811,In_467,In_542);
nand U812 (N_812,In_714,In_169);
and U813 (N_813,In_405,In_411);
nand U814 (N_814,In_96,In_556);
and U815 (N_815,In_8,In_633);
and U816 (N_816,In_315,In_166);
nand U817 (N_817,In_205,In_171);
nand U818 (N_818,In_65,In_613);
nand U819 (N_819,In_132,In_414);
nand U820 (N_820,In_614,In_675);
or U821 (N_821,In_57,In_490);
xnor U822 (N_822,In_656,In_584);
or U823 (N_823,In_163,In_661);
and U824 (N_824,In_433,In_586);
nand U825 (N_825,In_465,In_393);
or U826 (N_826,In_569,In_663);
nand U827 (N_827,In_251,In_374);
or U828 (N_828,In_510,In_17);
or U829 (N_829,In_29,In_640);
xor U830 (N_830,In_521,In_431);
and U831 (N_831,In_683,In_600);
nor U832 (N_832,In_235,In_179);
nand U833 (N_833,In_388,In_668);
or U834 (N_834,In_572,In_658);
nand U835 (N_835,In_308,In_180);
or U836 (N_836,In_139,In_5);
and U837 (N_837,In_314,In_65);
nand U838 (N_838,In_290,In_322);
or U839 (N_839,In_240,In_393);
nor U840 (N_840,In_422,In_381);
xor U841 (N_841,In_498,In_413);
or U842 (N_842,In_477,In_174);
nor U843 (N_843,In_169,In_596);
nor U844 (N_844,In_479,In_94);
or U845 (N_845,In_124,In_143);
and U846 (N_846,In_258,In_351);
nand U847 (N_847,In_687,In_133);
xor U848 (N_848,In_175,In_600);
or U849 (N_849,In_532,In_192);
nor U850 (N_850,In_717,In_110);
nand U851 (N_851,In_670,In_745);
and U852 (N_852,In_713,In_594);
nand U853 (N_853,In_639,In_278);
and U854 (N_854,In_496,In_455);
nor U855 (N_855,In_30,In_165);
and U856 (N_856,In_381,In_353);
and U857 (N_857,In_194,In_553);
and U858 (N_858,In_426,In_63);
and U859 (N_859,In_387,In_736);
nand U860 (N_860,In_264,In_10);
nor U861 (N_861,In_209,In_671);
nor U862 (N_862,In_214,In_88);
nor U863 (N_863,In_466,In_391);
and U864 (N_864,In_469,In_305);
nor U865 (N_865,In_5,In_28);
nand U866 (N_866,In_353,In_23);
nand U867 (N_867,In_65,In_587);
nand U868 (N_868,In_44,In_699);
or U869 (N_869,In_264,In_210);
or U870 (N_870,In_633,In_283);
nand U871 (N_871,In_641,In_246);
and U872 (N_872,In_690,In_136);
or U873 (N_873,In_573,In_515);
nor U874 (N_874,In_54,In_454);
or U875 (N_875,In_463,In_89);
and U876 (N_876,In_535,In_333);
and U877 (N_877,In_479,In_679);
or U878 (N_878,In_73,In_538);
or U879 (N_879,In_217,In_229);
or U880 (N_880,In_373,In_749);
and U881 (N_881,In_123,In_55);
nor U882 (N_882,In_554,In_549);
or U883 (N_883,In_273,In_92);
nor U884 (N_884,In_664,In_82);
or U885 (N_885,In_211,In_663);
or U886 (N_886,In_325,In_608);
nand U887 (N_887,In_389,In_450);
or U888 (N_888,In_235,In_729);
nor U889 (N_889,In_212,In_314);
nand U890 (N_890,In_691,In_546);
or U891 (N_891,In_392,In_228);
and U892 (N_892,In_34,In_403);
xnor U893 (N_893,In_231,In_482);
or U894 (N_894,In_451,In_483);
or U895 (N_895,In_387,In_157);
and U896 (N_896,In_286,In_528);
nand U897 (N_897,In_594,In_231);
or U898 (N_898,In_287,In_565);
or U899 (N_899,In_549,In_485);
and U900 (N_900,In_559,In_104);
nor U901 (N_901,In_520,In_689);
nand U902 (N_902,In_314,In_429);
nor U903 (N_903,In_127,In_452);
nand U904 (N_904,In_466,In_293);
nor U905 (N_905,In_371,In_176);
or U906 (N_906,In_287,In_60);
nand U907 (N_907,In_496,In_270);
or U908 (N_908,In_118,In_633);
or U909 (N_909,In_188,In_312);
nor U910 (N_910,In_681,In_557);
and U911 (N_911,In_564,In_75);
and U912 (N_912,In_50,In_364);
or U913 (N_913,In_487,In_464);
and U914 (N_914,In_285,In_388);
nand U915 (N_915,In_254,In_704);
or U916 (N_916,In_734,In_212);
nand U917 (N_917,In_195,In_82);
and U918 (N_918,In_137,In_13);
nor U919 (N_919,In_456,In_438);
xor U920 (N_920,In_613,In_600);
or U921 (N_921,In_416,In_709);
nand U922 (N_922,In_736,In_733);
or U923 (N_923,In_580,In_490);
or U924 (N_924,In_638,In_684);
or U925 (N_925,In_86,In_208);
or U926 (N_926,In_227,In_239);
or U927 (N_927,In_180,In_209);
or U928 (N_928,In_655,In_112);
nor U929 (N_929,In_747,In_446);
xor U930 (N_930,In_489,In_669);
and U931 (N_931,In_138,In_695);
nor U932 (N_932,In_450,In_686);
or U933 (N_933,In_513,In_354);
and U934 (N_934,In_102,In_61);
and U935 (N_935,In_726,In_370);
or U936 (N_936,In_94,In_348);
nor U937 (N_937,In_307,In_365);
and U938 (N_938,In_306,In_292);
and U939 (N_939,In_358,In_727);
nor U940 (N_940,In_337,In_289);
and U941 (N_941,In_589,In_124);
nor U942 (N_942,In_457,In_381);
and U943 (N_943,In_547,In_434);
nor U944 (N_944,In_624,In_144);
or U945 (N_945,In_31,In_508);
and U946 (N_946,In_20,In_566);
or U947 (N_947,In_328,In_747);
or U948 (N_948,In_268,In_468);
nor U949 (N_949,In_19,In_690);
nor U950 (N_950,In_414,In_153);
nand U951 (N_951,In_410,In_687);
and U952 (N_952,In_649,In_128);
and U953 (N_953,In_448,In_462);
nor U954 (N_954,In_36,In_626);
nor U955 (N_955,In_648,In_15);
nand U956 (N_956,In_339,In_718);
or U957 (N_957,In_334,In_160);
and U958 (N_958,In_414,In_463);
or U959 (N_959,In_0,In_146);
nand U960 (N_960,In_474,In_243);
nand U961 (N_961,In_360,In_673);
nor U962 (N_962,In_48,In_540);
or U963 (N_963,In_52,In_647);
nor U964 (N_964,In_252,In_595);
and U965 (N_965,In_441,In_287);
nor U966 (N_966,In_77,In_571);
and U967 (N_967,In_556,In_745);
or U968 (N_968,In_380,In_85);
nand U969 (N_969,In_365,In_687);
nand U970 (N_970,In_734,In_364);
nand U971 (N_971,In_370,In_142);
nor U972 (N_972,In_169,In_520);
nor U973 (N_973,In_239,In_648);
nor U974 (N_974,In_29,In_402);
or U975 (N_975,In_323,In_717);
or U976 (N_976,In_77,In_691);
xor U977 (N_977,In_16,In_693);
nor U978 (N_978,In_545,In_132);
and U979 (N_979,In_692,In_305);
nor U980 (N_980,In_610,In_727);
nand U981 (N_981,In_62,In_530);
nor U982 (N_982,In_103,In_253);
and U983 (N_983,In_35,In_30);
and U984 (N_984,In_557,In_421);
xnor U985 (N_985,In_526,In_620);
nor U986 (N_986,In_233,In_209);
nor U987 (N_987,In_141,In_696);
nor U988 (N_988,In_507,In_535);
nand U989 (N_989,In_611,In_19);
nor U990 (N_990,In_364,In_30);
or U991 (N_991,In_301,In_19);
and U992 (N_992,In_34,In_581);
and U993 (N_993,In_140,In_125);
nand U994 (N_994,In_377,In_234);
nand U995 (N_995,In_173,In_448);
nand U996 (N_996,In_575,In_162);
nand U997 (N_997,In_717,In_315);
and U998 (N_998,In_8,In_574);
and U999 (N_999,In_343,In_38);
and U1000 (N_1000,In_614,In_59);
and U1001 (N_1001,In_539,In_76);
and U1002 (N_1002,In_344,In_742);
nand U1003 (N_1003,In_240,In_684);
or U1004 (N_1004,In_126,In_345);
nor U1005 (N_1005,In_20,In_288);
nand U1006 (N_1006,In_28,In_299);
nor U1007 (N_1007,In_734,In_549);
or U1008 (N_1008,In_393,In_578);
nand U1009 (N_1009,In_747,In_248);
nand U1010 (N_1010,In_668,In_647);
nor U1011 (N_1011,In_391,In_534);
nand U1012 (N_1012,In_76,In_84);
or U1013 (N_1013,In_347,In_49);
nor U1014 (N_1014,In_658,In_194);
or U1015 (N_1015,In_163,In_472);
nor U1016 (N_1016,In_684,In_569);
nand U1017 (N_1017,In_21,In_521);
or U1018 (N_1018,In_241,In_606);
nand U1019 (N_1019,In_169,In_715);
nand U1020 (N_1020,In_253,In_613);
and U1021 (N_1021,In_633,In_676);
or U1022 (N_1022,In_38,In_144);
nand U1023 (N_1023,In_353,In_481);
nor U1024 (N_1024,In_14,In_590);
xnor U1025 (N_1025,In_200,In_706);
and U1026 (N_1026,In_173,In_463);
or U1027 (N_1027,In_12,In_587);
nand U1028 (N_1028,In_276,In_13);
nor U1029 (N_1029,In_586,In_699);
nand U1030 (N_1030,In_130,In_140);
nand U1031 (N_1031,In_474,In_186);
or U1032 (N_1032,In_446,In_157);
and U1033 (N_1033,In_182,In_237);
nand U1034 (N_1034,In_633,In_432);
or U1035 (N_1035,In_631,In_194);
nor U1036 (N_1036,In_727,In_68);
nand U1037 (N_1037,In_553,In_542);
and U1038 (N_1038,In_301,In_152);
nand U1039 (N_1039,In_711,In_708);
or U1040 (N_1040,In_669,In_375);
and U1041 (N_1041,In_186,In_545);
nand U1042 (N_1042,In_73,In_331);
nand U1043 (N_1043,In_370,In_176);
and U1044 (N_1044,In_482,In_709);
nor U1045 (N_1045,In_40,In_258);
nand U1046 (N_1046,In_135,In_680);
nor U1047 (N_1047,In_692,In_176);
nor U1048 (N_1048,In_699,In_562);
nand U1049 (N_1049,In_613,In_512);
or U1050 (N_1050,In_480,In_423);
or U1051 (N_1051,In_307,In_739);
or U1052 (N_1052,In_641,In_55);
nand U1053 (N_1053,In_655,In_356);
nor U1054 (N_1054,In_76,In_566);
nor U1055 (N_1055,In_633,In_288);
or U1056 (N_1056,In_666,In_246);
and U1057 (N_1057,In_197,In_495);
or U1058 (N_1058,In_360,In_653);
nand U1059 (N_1059,In_141,In_286);
nor U1060 (N_1060,In_234,In_123);
or U1061 (N_1061,In_457,In_484);
xor U1062 (N_1062,In_89,In_741);
or U1063 (N_1063,In_634,In_677);
nor U1064 (N_1064,In_161,In_68);
and U1065 (N_1065,In_451,In_79);
xor U1066 (N_1066,In_619,In_375);
nor U1067 (N_1067,In_632,In_641);
nand U1068 (N_1068,In_623,In_466);
nand U1069 (N_1069,In_737,In_126);
and U1070 (N_1070,In_685,In_3);
nor U1071 (N_1071,In_59,In_579);
nand U1072 (N_1072,In_659,In_183);
nor U1073 (N_1073,In_314,In_351);
nor U1074 (N_1074,In_613,In_374);
nand U1075 (N_1075,In_269,In_635);
nor U1076 (N_1076,In_97,In_273);
and U1077 (N_1077,In_88,In_116);
nor U1078 (N_1078,In_576,In_419);
and U1079 (N_1079,In_9,In_140);
and U1080 (N_1080,In_625,In_653);
nor U1081 (N_1081,In_403,In_549);
or U1082 (N_1082,In_700,In_442);
nand U1083 (N_1083,In_747,In_475);
and U1084 (N_1084,In_547,In_213);
nor U1085 (N_1085,In_431,In_515);
or U1086 (N_1086,In_747,In_504);
nor U1087 (N_1087,In_142,In_522);
nand U1088 (N_1088,In_158,In_290);
or U1089 (N_1089,In_27,In_414);
nor U1090 (N_1090,In_133,In_523);
xor U1091 (N_1091,In_199,In_581);
nand U1092 (N_1092,In_543,In_586);
and U1093 (N_1093,In_15,In_640);
and U1094 (N_1094,In_500,In_749);
and U1095 (N_1095,In_358,In_735);
or U1096 (N_1096,In_696,In_418);
nand U1097 (N_1097,In_572,In_634);
nand U1098 (N_1098,In_70,In_481);
nor U1099 (N_1099,In_3,In_737);
and U1100 (N_1100,In_736,In_49);
and U1101 (N_1101,In_658,In_127);
nor U1102 (N_1102,In_312,In_277);
nand U1103 (N_1103,In_714,In_48);
or U1104 (N_1104,In_492,In_559);
nand U1105 (N_1105,In_97,In_598);
or U1106 (N_1106,In_192,In_4);
nor U1107 (N_1107,In_321,In_707);
nand U1108 (N_1108,In_669,In_41);
nand U1109 (N_1109,In_267,In_285);
nand U1110 (N_1110,In_269,In_121);
or U1111 (N_1111,In_576,In_656);
and U1112 (N_1112,In_206,In_749);
and U1113 (N_1113,In_452,In_714);
nor U1114 (N_1114,In_40,In_498);
nor U1115 (N_1115,In_683,In_21);
and U1116 (N_1116,In_696,In_217);
nor U1117 (N_1117,In_307,In_717);
and U1118 (N_1118,In_377,In_646);
or U1119 (N_1119,In_255,In_626);
or U1120 (N_1120,In_641,In_178);
nand U1121 (N_1121,In_589,In_126);
and U1122 (N_1122,In_33,In_48);
and U1123 (N_1123,In_646,In_77);
or U1124 (N_1124,In_39,In_236);
nor U1125 (N_1125,In_422,In_359);
or U1126 (N_1126,In_564,In_625);
and U1127 (N_1127,In_371,In_308);
and U1128 (N_1128,In_584,In_331);
nor U1129 (N_1129,In_182,In_93);
nand U1130 (N_1130,In_618,In_379);
and U1131 (N_1131,In_136,In_517);
and U1132 (N_1132,In_346,In_498);
nor U1133 (N_1133,In_214,In_296);
or U1134 (N_1134,In_199,In_372);
or U1135 (N_1135,In_698,In_606);
nand U1136 (N_1136,In_193,In_725);
nand U1137 (N_1137,In_661,In_516);
nor U1138 (N_1138,In_585,In_270);
xor U1139 (N_1139,In_557,In_673);
xnor U1140 (N_1140,In_600,In_72);
and U1141 (N_1141,In_716,In_737);
nand U1142 (N_1142,In_634,In_409);
or U1143 (N_1143,In_640,In_616);
nand U1144 (N_1144,In_84,In_91);
and U1145 (N_1145,In_648,In_47);
nor U1146 (N_1146,In_695,In_602);
nor U1147 (N_1147,In_233,In_409);
nand U1148 (N_1148,In_45,In_578);
and U1149 (N_1149,In_460,In_69);
or U1150 (N_1150,In_279,In_306);
nand U1151 (N_1151,In_460,In_445);
and U1152 (N_1152,In_67,In_123);
or U1153 (N_1153,In_468,In_145);
nand U1154 (N_1154,In_731,In_15);
nor U1155 (N_1155,In_493,In_567);
nand U1156 (N_1156,In_514,In_454);
and U1157 (N_1157,In_226,In_30);
nand U1158 (N_1158,In_13,In_735);
nand U1159 (N_1159,In_42,In_320);
or U1160 (N_1160,In_562,In_110);
nor U1161 (N_1161,In_264,In_532);
or U1162 (N_1162,In_235,In_26);
and U1163 (N_1163,In_456,In_332);
nand U1164 (N_1164,In_414,In_198);
or U1165 (N_1165,In_164,In_360);
nand U1166 (N_1166,In_136,In_36);
nand U1167 (N_1167,In_465,In_472);
or U1168 (N_1168,In_307,In_483);
and U1169 (N_1169,In_703,In_573);
and U1170 (N_1170,In_532,In_299);
and U1171 (N_1171,In_187,In_95);
or U1172 (N_1172,In_720,In_15);
xnor U1173 (N_1173,In_310,In_375);
nor U1174 (N_1174,In_130,In_514);
nand U1175 (N_1175,In_709,In_704);
nor U1176 (N_1176,In_131,In_113);
nor U1177 (N_1177,In_27,In_314);
nor U1178 (N_1178,In_223,In_296);
nor U1179 (N_1179,In_613,In_486);
or U1180 (N_1180,In_182,In_121);
nand U1181 (N_1181,In_593,In_574);
nand U1182 (N_1182,In_483,In_419);
nand U1183 (N_1183,In_401,In_353);
nor U1184 (N_1184,In_62,In_609);
nand U1185 (N_1185,In_602,In_75);
nand U1186 (N_1186,In_131,In_356);
nand U1187 (N_1187,In_77,In_436);
or U1188 (N_1188,In_405,In_109);
xnor U1189 (N_1189,In_84,In_172);
and U1190 (N_1190,In_588,In_138);
nor U1191 (N_1191,In_333,In_573);
nor U1192 (N_1192,In_293,In_205);
or U1193 (N_1193,In_635,In_328);
and U1194 (N_1194,In_647,In_400);
nor U1195 (N_1195,In_736,In_478);
or U1196 (N_1196,In_293,In_200);
nor U1197 (N_1197,In_423,In_475);
nand U1198 (N_1198,In_210,In_341);
nor U1199 (N_1199,In_15,In_555);
nor U1200 (N_1200,In_643,In_655);
nor U1201 (N_1201,In_440,In_208);
and U1202 (N_1202,In_330,In_736);
and U1203 (N_1203,In_624,In_161);
xor U1204 (N_1204,In_352,In_446);
or U1205 (N_1205,In_278,In_42);
nand U1206 (N_1206,In_386,In_556);
or U1207 (N_1207,In_602,In_261);
and U1208 (N_1208,In_616,In_233);
and U1209 (N_1209,In_412,In_219);
or U1210 (N_1210,In_85,In_318);
nand U1211 (N_1211,In_701,In_47);
nand U1212 (N_1212,In_24,In_135);
nand U1213 (N_1213,In_232,In_188);
nor U1214 (N_1214,In_580,In_70);
and U1215 (N_1215,In_533,In_324);
or U1216 (N_1216,In_543,In_637);
nor U1217 (N_1217,In_709,In_312);
nand U1218 (N_1218,In_359,In_33);
and U1219 (N_1219,In_82,In_299);
and U1220 (N_1220,In_412,In_51);
nand U1221 (N_1221,In_391,In_265);
or U1222 (N_1222,In_185,In_261);
nand U1223 (N_1223,In_587,In_56);
xor U1224 (N_1224,In_685,In_282);
nand U1225 (N_1225,In_536,In_558);
xnor U1226 (N_1226,In_700,In_643);
or U1227 (N_1227,In_121,In_136);
nor U1228 (N_1228,In_352,In_508);
or U1229 (N_1229,In_181,In_506);
nor U1230 (N_1230,In_739,In_53);
and U1231 (N_1231,In_691,In_102);
nand U1232 (N_1232,In_631,In_721);
nor U1233 (N_1233,In_399,In_574);
or U1234 (N_1234,In_28,In_496);
or U1235 (N_1235,In_67,In_712);
nor U1236 (N_1236,In_258,In_39);
nor U1237 (N_1237,In_583,In_211);
and U1238 (N_1238,In_143,In_487);
or U1239 (N_1239,In_230,In_451);
nand U1240 (N_1240,In_55,In_435);
and U1241 (N_1241,In_422,In_442);
xor U1242 (N_1242,In_455,In_478);
or U1243 (N_1243,In_523,In_328);
nand U1244 (N_1244,In_221,In_24);
or U1245 (N_1245,In_408,In_182);
and U1246 (N_1246,In_520,In_501);
nor U1247 (N_1247,In_691,In_50);
nor U1248 (N_1248,In_149,In_159);
nand U1249 (N_1249,In_607,In_197);
or U1250 (N_1250,In_515,In_733);
and U1251 (N_1251,In_680,In_261);
or U1252 (N_1252,In_403,In_634);
nor U1253 (N_1253,In_660,In_620);
and U1254 (N_1254,In_703,In_599);
and U1255 (N_1255,In_619,In_1);
nand U1256 (N_1256,In_389,In_732);
or U1257 (N_1257,In_295,In_107);
nand U1258 (N_1258,In_686,In_194);
or U1259 (N_1259,In_65,In_588);
nand U1260 (N_1260,In_280,In_345);
or U1261 (N_1261,In_624,In_580);
nand U1262 (N_1262,In_493,In_10);
or U1263 (N_1263,In_417,In_169);
or U1264 (N_1264,In_428,In_370);
xnor U1265 (N_1265,In_735,In_394);
and U1266 (N_1266,In_501,In_742);
nor U1267 (N_1267,In_380,In_269);
and U1268 (N_1268,In_514,In_563);
and U1269 (N_1269,In_246,In_418);
and U1270 (N_1270,In_420,In_583);
or U1271 (N_1271,In_45,In_511);
xnor U1272 (N_1272,In_370,In_290);
and U1273 (N_1273,In_73,In_730);
or U1274 (N_1274,In_206,In_595);
or U1275 (N_1275,In_50,In_170);
or U1276 (N_1276,In_227,In_507);
nand U1277 (N_1277,In_297,In_525);
nor U1278 (N_1278,In_377,In_383);
and U1279 (N_1279,In_454,In_81);
nand U1280 (N_1280,In_472,In_487);
and U1281 (N_1281,In_237,In_170);
or U1282 (N_1282,In_586,In_414);
or U1283 (N_1283,In_554,In_87);
and U1284 (N_1284,In_356,In_109);
nor U1285 (N_1285,In_712,In_199);
and U1286 (N_1286,In_51,In_299);
or U1287 (N_1287,In_137,In_493);
nand U1288 (N_1288,In_75,In_627);
nor U1289 (N_1289,In_208,In_311);
and U1290 (N_1290,In_723,In_223);
or U1291 (N_1291,In_307,In_747);
nor U1292 (N_1292,In_743,In_373);
or U1293 (N_1293,In_645,In_232);
and U1294 (N_1294,In_67,In_419);
or U1295 (N_1295,In_473,In_606);
nand U1296 (N_1296,In_484,In_574);
or U1297 (N_1297,In_179,In_282);
nor U1298 (N_1298,In_537,In_476);
nor U1299 (N_1299,In_710,In_247);
nand U1300 (N_1300,In_450,In_73);
nor U1301 (N_1301,In_248,In_433);
and U1302 (N_1302,In_534,In_587);
nand U1303 (N_1303,In_447,In_322);
nand U1304 (N_1304,In_453,In_149);
nand U1305 (N_1305,In_692,In_371);
nand U1306 (N_1306,In_335,In_292);
and U1307 (N_1307,In_100,In_520);
nand U1308 (N_1308,In_99,In_414);
and U1309 (N_1309,In_173,In_376);
nand U1310 (N_1310,In_78,In_522);
or U1311 (N_1311,In_30,In_461);
nand U1312 (N_1312,In_55,In_463);
or U1313 (N_1313,In_107,In_588);
and U1314 (N_1314,In_585,In_692);
and U1315 (N_1315,In_586,In_489);
nor U1316 (N_1316,In_360,In_643);
nand U1317 (N_1317,In_45,In_37);
nor U1318 (N_1318,In_384,In_581);
nand U1319 (N_1319,In_391,In_85);
and U1320 (N_1320,In_165,In_256);
or U1321 (N_1321,In_25,In_351);
nor U1322 (N_1322,In_335,In_506);
or U1323 (N_1323,In_347,In_530);
nor U1324 (N_1324,In_618,In_258);
nand U1325 (N_1325,In_486,In_98);
nor U1326 (N_1326,In_267,In_474);
and U1327 (N_1327,In_692,In_737);
nor U1328 (N_1328,In_43,In_420);
nor U1329 (N_1329,In_172,In_697);
and U1330 (N_1330,In_650,In_653);
nor U1331 (N_1331,In_620,In_52);
nor U1332 (N_1332,In_402,In_279);
nor U1333 (N_1333,In_689,In_323);
and U1334 (N_1334,In_338,In_57);
xnor U1335 (N_1335,In_232,In_364);
or U1336 (N_1336,In_5,In_698);
and U1337 (N_1337,In_129,In_605);
and U1338 (N_1338,In_312,In_201);
and U1339 (N_1339,In_74,In_425);
or U1340 (N_1340,In_260,In_97);
nor U1341 (N_1341,In_83,In_392);
nand U1342 (N_1342,In_574,In_407);
nor U1343 (N_1343,In_69,In_463);
or U1344 (N_1344,In_224,In_236);
nand U1345 (N_1345,In_348,In_391);
nor U1346 (N_1346,In_652,In_363);
nor U1347 (N_1347,In_238,In_146);
nor U1348 (N_1348,In_749,In_668);
and U1349 (N_1349,In_315,In_6);
nor U1350 (N_1350,In_63,In_422);
and U1351 (N_1351,In_356,In_283);
nand U1352 (N_1352,In_122,In_668);
nor U1353 (N_1353,In_89,In_240);
and U1354 (N_1354,In_325,In_109);
or U1355 (N_1355,In_415,In_42);
and U1356 (N_1356,In_257,In_152);
nand U1357 (N_1357,In_470,In_321);
nand U1358 (N_1358,In_92,In_697);
nand U1359 (N_1359,In_0,In_614);
or U1360 (N_1360,In_640,In_524);
or U1361 (N_1361,In_487,In_61);
nand U1362 (N_1362,In_56,In_262);
nand U1363 (N_1363,In_234,In_533);
or U1364 (N_1364,In_453,In_66);
or U1365 (N_1365,In_595,In_277);
and U1366 (N_1366,In_421,In_2);
nand U1367 (N_1367,In_417,In_576);
nand U1368 (N_1368,In_149,In_569);
nand U1369 (N_1369,In_151,In_156);
nor U1370 (N_1370,In_526,In_210);
or U1371 (N_1371,In_578,In_194);
nor U1372 (N_1372,In_329,In_666);
nand U1373 (N_1373,In_86,In_285);
and U1374 (N_1374,In_749,In_652);
and U1375 (N_1375,In_28,In_699);
or U1376 (N_1376,In_206,In_167);
and U1377 (N_1377,In_429,In_742);
nand U1378 (N_1378,In_27,In_709);
nand U1379 (N_1379,In_260,In_104);
nand U1380 (N_1380,In_602,In_444);
or U1381 (N_1381,In_706,In_126);
nor U1382 (N_1382,In_444,In_541);
nand U1383 (N_1383,In_579,In_190);
and U1384 (N_1384,In_701,In_395);
or U1385 (N_1385,In_124,In_54);
nand U1386 (N_1386,In_690,In_38);
nand U1387 (N_1387,In_721,In_737);
and U1388 (N_1388,In_279,In_545);
and U1389 (N_1389,In_402,In_362);
nand U1390 (N_1390,In_461,In_543);
nor U1391 (N_1391,In_708,In_668);
and U1392 (N_1392,In_311,In_517);
nor U1393 (N_1393,In_5,In_262);
nor U1394 (N_1394,In_50,In_743);
nor U1395 (N_1395,In_176,In_109);
nor U1396 (N_1396,In_355,In_276);
nor U1397 (N_1397,In_488,In_651);
and U1398 (N_1398,In_457,In_380);
nand U1399 (N_1399,In_708,In_733);
or U1400 (N_1400,In_535,In_444);
nand U1401 (N_1401,In_602,In_243);
or U1402 (N_1402,In_423,In_42);
and U1403 (N_1403,In_60,In_678);
or U1404 (N_1404,In_544,In_135);
and U1405 (N_1405,In_487,In_141);
or U1406 (N_1406,In_214,In_667);
nand U1407 (N_1407,In_295,In_132);
and U1408 (N_1408,In_720,In_711);
and U1409 (N_1409,In_21,In_662);
or U1410 (N_1410,In_258,In_714);
and U1411 (N_1411,In_390,In_307);
or U1412 (N_1412,In_496,In_404);
xor U1413 (N_1413,In_209,In_447);
nor U1414 (N_1414,In_515,In_167);
and U1415 (N_1415,In_220,In_85);
nor U1416 (N_1416,In_80,In_552);
and U1417 (N_1417,In_608,In_516);
nor U1418 (N_1418,In_692,In_88);
and U1419 (N_1419,In_727,In_421);
and U1420 (N_1420,In_344,In_268);
nand U1421 (N_1421,In_714,In_190);
xor U1422 (N_1422,In_711,In_609);
nor U1423 (N_1423,In_295,In_245);
nand U1424 (N_1424,In_321,In_643);
nand U1425 (N_1425,In_99,In_229);
nor U1426 (N_1426,In_65,In_329);
nor U1427 (N_1427,In_67,In_287);
and U1428 (N_1428,In_267,In_137);
and U1429 (N_1429,In_323,In_574);
nor U1430 (N_1430,In_13,In_296);
nor U1431 (N_1431,In_586,In_369);
nor U1432 (N_1432,In_638,In_704);
or U1433 (N_1433,In_487,In_200);
nand U1434 (N_1434,In_244,In_315);
nand U1435 (N_1435,In_580,In_136);
and U1436 (N_1436,In_725,In_407);
nor U1437 (N_1437,In_334,In_225);
or U1438 (N_1438,In_40,In_440);
nand U1439 (N_1439,In_720,In_26);
and U1440 (N_1440,In_112,In_251);
nand U1441 (N_1441,In_377,In_469);
or U1442 (N_1442,In_234,In_115);
and U1443 (N_1443,In_136,In_93);
and U1444 (N_1444,In_208,In_512);
nor U1445 (N_1445,In_467,In_694);
nand U1446 (N_1446,In_325,In_304);
and U1447 (N_1447,In_696,In_281);
nand U1448 (N_1448,In_266,In_699);
and U1449 (N_1449,In_543,In_523);
or U1450 (N_1450,In_610,In_649);
or U1451 (N_1451,In_724,In_393);
or U1452 (N_1452,In_391,In_735);
nor U1453 (N_1453,In_279,In_285);
nand U1454 (N_1454,In_430,In_413);
nand U1455 (N_1455,In_704,In_93);
and U1456 (N_1456,In_430,In_253);
or U1457 (N_1457,In_269,In_230);
nand U1458 (N_1458,In_4,In_363);
and U1459 (N_1459,In_513,In_123);
and U1460 (N_1460,In_302,In_342);
nand U1461 (N_1461,In_689,In_110);
or U1462 (N_1462,In_53,In_36);
or U1463 (N_1463,In_439,In_398);
xor U1464 (N_1464,In_508,In_57);
and U1465 (N_1465,In_443,In_292);
nor U1466 (N_1466,In_32,In_337);
and U1467 (N_1467,In_662,In_730);
nor U1468 (N_1468,In_61,In_479);
or U1469 (N_1469,In_48,In_203);
nand U1470 (N_1470,In_698,In_638);
nor U1471 (N_1471,In_363,In_5);
nand U1472 (N_1472,In_390,In_497);
and U1473 (N_1473,In_688,In_312);
nand U1474 (N_1474,In_111,In_614);
or U1475 (N_1475,In_315,In_383);
nor U1476 (N_1476,In_417,In_489);
or U1477 (N_1477,In_727,In_8);
or U1478 (N_1478,In_519,In_262);
nor U1479 (N_1479,In_674,In_150);
and U1480 (N_1480,In_63,In_538);
and U1481 (N_1481,In_692,In_323);
nor U1482 (N_1482,In_420,In_246);
or U1483 (N_1483,In_262,In_223);
and U1484 (N_1484,In_251,In_53);
nand U1485 (N_1485,In_222,In_331);
nand U1486 (N_1486,In_2,In_63);
or U1487 (N_1487,In_260,In_627);
nand U1488 (N_1488,In_657,In_714);
and U1489 (N_1489,In_395,In_588);
nor U1490 (N_1490,In_64,In_682);
nor U1491 (N_1491,In_375,In_534);
nand U1492 (N_1492,In_360,In_670);
nor U1493 (N_1493,In_158,In_380);
and U1494 (N_1494,In_725,In_261);
and U1495 (N_1495,In_722,In_129);
nand U1496 (N_1496,In_489,In_253);
or U1497 (N_1497,In_300,In_110);
or U1498 (N_1498,In_720,In_291);
and U1499 (N_1499,In_348,In_525);
nor U1500 (N_1500,In_228,In_493);
nand U1501 (N_1501,In_718,In_608);
or U1502 (N_1502,In_653,In_329);
nor U1503 (N_1503,In_527,In_436);
or U1504 (N_1504,In_91,In_590);
and U1505 (N_1505,In_686,In_369);
or U1506 (N_1506,In_168,In_596);
nand U1507 (N_1507,In_682,In_129);
nor U1508 (N_1508,In_390,In_370);
and U1509 (N_1509,In_521,In_425);
nor U1510 (N_1510,In_170,In_141);
or U1511 (N_1511,In_481,In_172);
or U1512 (N_1512,In_714,In_583);
or U1513 (N_1513,In_673,In_408);
and U1514 (N_1514,In_627,In_484);
nand U1515 (N_1515,In_742,In_246);
and U1516 (N_1516,In_554,In_142);
or U1517 (N_1517,In_450,In_193);
and U1518 (N_1518,In_391,In_424);
nand U1519 (N_1519,In_257,In_619);
and U1520 (N_1520,In_454,In_4);
and U1521 (N_1521,In_695,In_624);
nand U1522 (N_1522,In_497,In_363);
nor U1523 (N_1523,In_176,In_588);
nand U1524 (N_1524,In_718,In_433);
and U1525 (N_1525,In_577,In_731);
or U1526 (N_1526,In_378,In_447);
or U1527 (N_1527,In_224,In_597);
nor U1528 (N_1528,In_648,In_737);
and U1529 (N_1529,In_21,In_406);
nor U1530 (N_1530,In_415,In_406);
and U1531 (N_1531,In_272,In_55);
or U1532 (N_1532,In_506,In_633);
and U1533 (N_1533,In_267,In_652);
nand U1534 (N_1534,In_449,In_374);
or U1535 (N_1535,In_342,In_558);
or U1536 (N_1536,In_248,In_693);
and U1537 (N_1537,In_41,In_710);
and U1538 (N_1538,In_85,In_725);
nand U1539 (N_1539,In_218,In_610);
nor U1540 (N_1540,In_279,In_308);
nand U1541 (N_1541,In_157,In_733);
nor U1542 (N_1542,In_338,In_97);
nand U1543 (N_1543,In_519,In_465);
nor U1544 (N_1544,In_716,In_651);
or U1545 (N_1545,In_702,In_705);
and U1546 (N_1546,In_90,In_465);
nand U1547 (N_1547,In_553,In_243);
and U1548 (N_1548,In_342,In_401);
and U1549 (N_1549,In_79,In_392);
or U1550 (N_1550,In_401,In_51);
or U1551 (N_1551,In_157,In_362);
nand U1552 (N_1552,In_403,In_42);
xor U1553 (N_1553,In_619,In_610);
nand U1554 (N_1554,In_399,In_296);
or U1555 (N_1555,In_532,In_370);
nand U1556 (N_1556,In_404,In_491);
xnor U1557 (N_1557,In_372,In_612);
nor U1558 (N_1558,In_195,In_613);
nor U1559 (N_1559,In_410,In_629);
nor U1560 (N_1560,In_7,In_622);
and U1561 (N_1561,In_131,In_586);
or U1562 (N_1562,In_362,In_523);
or U1563 (N_1563,In_389,In_623);
and U1564 (N_1564,In_578,In_239);
and U1565 (N_1565,In_465,In_222);
nand U1566 (N_1566,In_305,In_588);
nor U1567 (N_1567,In_506,In_625);
nor U1568 (N_1568,In_525,In_400);
nand U1569 (N_1569,In_133,In_275);
nand U1570 (N_1570,In_74,In_481);
and U1571 (N_1571,In_306,In_102);
and U1572 (N_1572,In_695,In_746);
nor U1573 (N_1573,In_654,In_214);
nor U1574 (N_1574,In_6,In_645);
and U1575 (N_1575,In_78,In_475);
or U1576 (N_1576,In_472,In_741);
nand U1577 (N_1577,In_331,In_514);
and U1578 (N_1578,In_58,In_430);
nand U1579 (N_1579,In_648,In_700);
and U1580 (N_1580,In_436,In_533);
nand U1581 (N_1581,In_460,In_131);
and U1582 (N_1582,In_37,In_731);
nor U1583 (N_1583,In_493,In_151);
nand U1584 (N_1584,In_323,In_28);
or U1585 (N_1585,In_661,In_162);
nor U1586 (N_1586,In_336,In_354);
nor U1587 (N_1587,In_340,In_18);
and U1588 (N_1588,In_632,In_539);
nand U1589 (N_1589,In_733,In_680);
and U1590 (N_1590,In_165,In_134);
nand U1591 (N_1591,In_732,In_261);
nor U1592 (N_1592,In_164,In_278);
and U1593 (N_1593,In_689,In_678);
and U1594 (N_1594,In_398,In_410);
nand U1595 (N_1595,In_681,In_192);
and U1596 (N_1596,In_118,In_614);
and U1597 (N_1597,In_40,In_308);
nand U1598 (N_1598,In_591,In_92);
nand U1599 (N_1599,In_150,In_263);
or U1600 (N_1600,In_478,In_453);
and U1601 (N_1601,In_449,In_686);
and U1602 (N_1602,In_72,In_507);
xnor U1603 (N_1603,In_133,In_309);
nand U1604 (N_1604,In_349,In_509);
nor U1605 (N_1605,In_526,In_714);
and U1606 (N_1606,In_714,In_644);
nand U1607 (N_1607,In_131,In_621);
and U1608 (N_1608,In_445,In_645);
nand U1609 (N_1609,In_449,In_588);
and U1610 (N_1610,In_735,In_280);
nand U1611 (N_1611,In_45,In_728);
nor U1612 (N_1612,In_2,In_529);
and U1613 (N_1613,In_684,In_503);
nor U1614 (N_1614,In_604,In_48);
and U1615 (N_1615,In_224,In_623);
or U1616 (N_1616,In_45,In_43);
nand U1617 (N_1617,In_186,In_109);
and U1618 (N_1618,In_460,In_71);
nor U1619 (N_1619,In_82,In_672);
nor U1620 (N_1620,In_383,In_65);
nor U1621 (N_1621,In_395,In_452);
nor U1622 (N_1622,In_139,In_414);
or U1623 (N_1623,In_333,In_625);
and U1624 (N_1624,In_684,In_458);
and U1625 (N_1625,In_84,In_393);
nand U1626 (N_1626,In_259,In_613);
or U1627 (N_1627,In_664,In_382);
and U1628 (N_1628,In_610,In_549);
and U1629 (N_1629,In_11,In_625);
xnor U1630 (N_1630,In_91,In_213);
and U1631 (N_1631,In_184,In_418);
nand U1632 (N_1632,In_522,In_513);
and U1633 (N_1633,In_322,In_260);
nand U1634 (N_1634,In_344,In_203);
xor U1635 (N_1635,In_404,In_689);
nor U1636 (N_1636,In_660,In_183);
or U1637 (N_1637,In_690,In_516);
nand U1638 (N_1638,In_350,In_679);
xnor U1639 (N_1639,In_515,In_232);
or U1640 (N_1640,In_448,In_550);
nand U1641 (N_1641,In_363,In_407);
nor U1642 (N_1642,In_407,In_215);
nor U1643 (N_1643,In_12,In_343);
nor U1644 (N_1644,In_415,In_51);
and U1645 (N_1645,In_740,In_498);
and U1646 (N_1646,In_153,In_640);
nand U1647 (N_1647,In_227,In_184);
nand U1648 (N_1648,In_201,In_448);
nor U1649 (N_1649,In_653,In_408);
nor U1650 (N_1650,In_507,In_488);
nand U1651 (N_1651,In_38,In_250);
nand U1652 (N_1652,In_180,In_556);
and U1653 (N_1653,In_427,In_363);
nor U1654 (N_1654,In_435,In_516);
nor U1655 (N_1655,In_180,In_740);
nor U1656 (N_1656,In_105,In_98);
nor U1657 (N_1657,In_197,In_445);
nand U1658 (N_1658,In_26,In_508);
or U1659 (N_1659,In_454,In_329);
and U1660 (N_1660,In_361,In_55);
nand U1661 (N_1661,In_680,In_3);
or U1662 (N_1662,In_673,In_315);
and U1663 (N_1663,In_360,In_427);
xor U1664 (N_1664,In_603,In_511);
or U1665 (N_1665,In_256,In_714);
nor U1666 (N_1666,In_717,In_695);
nor U1667 (N_1667,In_664,In_319);
nor U1668 (N_1668,In_399,In_106);
and U1669 (N_1669,In_364,In_584);
nand U1670 (N_1670,In_710,In_743);
and U1671 (N_1671,In_458,In_136);
and U1672 (N_1672,In_477,In_250);
or U1673 (N_1673,In_14,In_565);
nor U1674 (N_1674,In_86,In_110);
nand U1675 (N_1675,In_730,In_748);
and U1676 (N_1676,In_447,In_398);
nor U1677 (N_1677,In_23,In_304);
and U1678 (N_1678,In_348,In_285);
nand U1679 (N_1679,In_157,In_255);
nand U1680 (N_1680,In_342,In_55);
or U1681 (N_1681,In_470,In_729);
and U1682 (N_1682,In_618,In_529);
or U1683 (N_1683,In_377,In_174);
or U1684 (N_1684,In_370,In_166);
nand U1685 (N_1685,In_266,In_349);
nor U1686 (N_1686,In_709,In_301);
and U1687 (N_1687,In_151,In_230);
nand U1688 (N_1688,In_367,In_570);
nand U1689 (N_1689,In_494,In_168);
nor U1690 (N_1690,In_168,In_357);
nand U1691 (N_1691,In_252,In_79);
xnor U1692 (N_1692,In_682,In_647);
or U1693 (N_1693,In_102,In_329);
nand U1694 (N_1694,In_474,In_623);
or U1695 (N_1695,In_81,In_342);
nand U1696 (N_1696,In_140,In_665);
and U1697 (N_1697,In_690,In_44);
or U1698 (N_1698,In_619,In_203);
nor U1699 (N_1699,In_224,In_218);
nand U1700 (N_1700,In_443,In_345);
or U1701 (N_1701,In_80,In_396);
nor U1702 (N_1702,In_137,In_53);
nor U1703 (N_1703,In_76,In_628);
or U1704 (N_1704,In_706,In_0);
or U1705 (N_1705,In_732,In_184);
or U1706 (N_1706,In_505,In_665);
nor U1707 (N_1707,In_577,In_333);
or U1708 (N_1708,In_214,In_497);
nand U1709 (N_1709,In_200,In_57);
nor U1710 (N_1710,In_641,In_693);
nor U1711 (N_1711,In_547,In_360);
or U1712 (N_1712,In_570,In_220);
nand U1713 (N_1713,In_230,In_652);
or U1714 (N_1714,In_236,In_659);
or U1715 (N_1715,In_114,In_496);
or U1716 (N_1716,In_235,In_55);
xor U1717 (N_1717,In_566,In_27);
nor U1718 (N_1718,In_576,In_335);
nand U1719 (N_1719,In_478,In_204);
or U1720 (N_1720,In_535,In_362);
and U1721 (N_1721,In_706,In_137);
or U1722 (N_1722,In_4,In_209);
nor U1723 (N_1723,In_588,In_199);
nand U1724 (N_1724,In_156,In_628);
or U1725 (N_1725,In_657,In_44);
nor U1726 (N_1726,In_325,In_31);
nand U1727 (N_1727,In_438,In_90);
or U1728 (N_1728,In_403,In_397);
nor U1729 (N_1729,In_610,In_273);
or U1730 (N_1730,In_719,In_571);
nor U1731 (N_1731,In_291,In_543);
or U1732 (N_1732,In_479,In_730);
nor U1733 (N_1733,In_634,In_426);
or U1734 (N_1734,In_390,In_372);
and U1735 (N_1735,In_205,In_652);
and U1736 (N_1736,In_404,In_645);
nand U1737 (N_1737,In_740,In_637);
nand U1738 (N_1738,In_435,In_329);
nand U1739 (N_1739,In_485,In_244);
and U1740 (N_1740,In_408,In_194);
nor U1741 (N_1741,In_719,In_327);
and U1742 (N_1742,In_637,In_43);
nor U1743 (N_1743,In_259,In_188);
nor U1744 (N_1744,In_259,In_595);
nor U1745 (N_1745,In_569,In_84);
and U1746 (N_1746,In_394,In_393);
nand U1747 (N_1747,In_104,In_232);
nand U1748 (N_1748,In_347,In_273);
and U1749 (N_1749,In_706,In_741);
or U1750 (N_1750,In_161,In_653);
and U1751 (N_1751,In_377,In_299);
and U1752 (N_1752,In_310,In_617);
and U1753 (N_1753,In_194,In_705);
or U1754 (N_1754,In_599,In_509);
or U1755 (N_1755,In_70,In_141);
and U1756 (N_1756,In_83,In_692);
and U1757 (N_1757,In_650,In_599);
and U1758 (N_1758,In_387,In_35);
nor U1759 (N_1759,In_204,In_153);
nand U1760 (N_1760,In_462,In_545);
or U1761 (N_1761,In_37,In_715);
nor U1762 (N_1762,In_221,In_749);
xnor U1763 (N_1763,In_640,In_569);
or U1764 (N_1764,In_538,In_235);
nor U1765 (N_1765,In_560,In_647);
nor U1766 (N_1766,In_233,In_380);
or U1767 (N_1767,In_680,In_670);
nor U1768 (N_1768,In_746,In_105);
and U1769 (N_1769,In_237,In_435);
and U1770 (N_1770,In_714,In_31);
xor U1771 (N_1771,In_352,In_346);
nor U1772 (N_1772,In_154,In_610);
and U1773 (N_1773,In_733,In_375);
nor U1774 (N_1774,In_486,In_255);
nor U1775 (N_1775,In_18,In_176);
nor U1776 (N_1776,In_324,In_402);
nand U1777 (N_1777,In_235,In_63);
or U1778 (N_1778,In_18,In_547);
nand U1779 (N_1779,In_443,In_254);
or U1780 (N_1780,In_28,In_145);
and U1781 (N_1781,In_118,In_23);
or U1782 (N_1782,In_392,In_666);
nor U1783 (N_1783,In_281,In_444);
nand U1784 (N_1784,In_15,In_425);
or U1785 (N_1785,In_267,In_468);
and U1786 (N_1786,In_82,In_396);
nand U1787 (N_1787,In_235,In_540);
nand U1788 (N_1788,In_432,In_648);
and U1789 (N_1789,In_116,In_654);
or U1790 (N_1790,In_229,In_16);
and U1791 (N_1791,In_576,In_133);
or U1792 (N_1792,In_308,In_665);
nand U1793 (N_1793,In_658,In_376);
nand U1794 (N_1794,In_697,In_348);
nand U1795 (N_1795,In_614,In_492);
nor U1796 (N_1796,In_317,In_489);
or U1797 (N_1797,In_535,In_40);
nor U1798 (N_1798,In_337,In_55);
nand U1799 (N_1799,In_740,In_56);
or U1800 (N_1800,In_549,In_544);
or U1801 (N_1801,In_156,In_637);
and U1802 (N_1802,In_508,In_572);
nand U1803 (N_1803,In_399,In_466);
nand U1804 (N_1804,In_431,In_610);
nor U1805 (N_1805,In_669,In_134);
nand U1806 (N_1806,In_95,In_461);
and U1807 (N_1807,In_143,In_715);
nand U1808 (N_1808,In_525,In_119);
and U1809 (N_1809,In_439,In_318);
nor U1810 (N_1810,In_206,In_506);
and U1811 (N_1811,In_546,In_430);
or U1812 (N_1812,In_745,In_118);
nor U1813 (N_1813,In_671,In_405);
nand U1814 (N_1814,In_335,In_5);
nand U1815 (N_1815,In_6,In_196);
nor U1816 (N_1816,In_158,In_429);
or U1817 (N_1817,In_251,In_91);
or U1818 (N_1818,In_436,In_617);
nand U1819 (N_1819,In_550,In_598);
nor U1820 (N_1820,In_479,In_439);
nand U1821 (N_1821,In_741,In_537);
and U1822 (N_1822,In_248,In_274);
nor U1823 (N_1823,In_552,In_58);
or U1824 (N_1824,In_181,In_172);
xnor U1825 (N_1825,In_528,In_153);
nand U1826 (N_1826,In_521,In_476);
nor U1827 (N_1827,In_340,In_679);
nand U1828 (N_1828,In_487,In_396);
nor U1829 (N_1829,In_502,In_351);
nor U1830 (N_1830,In_461,In_665);
xnor U1831 (N_1831,In_710,In_547);
nor U1832 (N_1832,In_305,In_157);
or U1833 (N_1833,In_516,In_703);
and U1834 (N_1834,In_640,In_741);
nand U1835 (N_1835,In_746,In_288);
nand U1836 (N_1836,In_492,In_32);
and U1837 (N_1837,In_715,In_277);
and U1838 (N_1838,In_201,In_403);
nand U1839 (N_1839,In_440,In_317);
or U1840 (N_1840,In_168,In_446);
nor U1841 (N_1841,In_48,In_311);
nor U1842 (N_1842,In_1,In_334);
or U1843 (N_1843,In_189,In_134);
and U1844 (N_1844,In_361,In_121);
or U1845 (N_1845,In_255,In_146);
nor U1846 (N_1846,In_264,In_409);
and U1847 (N_1847,In_40,In_64);
nor U1848 (N_1848,In_357,In_579);
nor U1849 (N_1849,In_512,In_730);
nand U1850 (N_1850,In_449,In_417);
and U1851 (N_1851,In_650,In_160);
or U1852 (N_1852,In_267,In_648);
nor U1853 (N_1853,In_596,In_607);
xor U1854 (N_1854,In_321,In_383);
nand U1855 (N_1855,In_407,In_709);
and U1856 (N_1856,In_361,In_651);
or U1857 (N_1857,In_101,In_301);
or U1858 (N_1858,In_113,In_412);
nand U1859 (N_1859,In_407,In_224);
nor U1860 (N_1860,In_459,In_587);
nand U1861 (N_1861,In_404,In_469);
or U1862 (N_1862,In_729,In_332);
nor U1863 (N_1863,In_255,In_69);
xor U1864 (N_1864,In_250,In_230);
and U1865 (N_1865,In_173,In_502);
nor U1866 (N_1866,In_246,In_127);
or U1867 (N_1867,In_461,In_141);
nor U1868 (N_1868,In_605,In_372);
nand U1869 (N_1869,In_97,In_220);
nor U1870 (N_1870,In_472,In_516);
nor U1871 (N_1871,In_722,In_660);
nor U1872 (N_1872,In_55,In_20);
nand U1873 (N_1873,In_337,In_537);
or U1874 (N_1874,In_208,In_505);
nor U1875 (N_1875,In_658,In_594);
nor U1876 (N_1876,In_375,In_42);
or U1877 (N_1877,In_634,In_109);
nand U1878 (N_1878,In_220,In_528);
and U1879 (N_1879,In_693,In_593);
or U1880 (N_1880,In_206,In_593);
nor U1881 (N_1881,In_274,In_661);
nor U1882 (N_1882,In_184,In_278);
nor U1883 (N_1883,In_487,In_208);
or U1884 (N_1884,In_587,In_105);
nor U1885 (N_1885,In_207,In_65);
nand U1886 (N_1886,In_643,In_377);
nand U1887 (N_1887,In_392,In_340);
nor U1888 (N_1888,In_457,In_535);
and U1889 (N_1889,In_65,In_594);
nand U1890 (N_1890,In_454,In_675);
nand U1891 (N_1891,In_457,In_408);
nand U1892 (N_1892,In_54,In_706);
nor U1893 (N_1893,In_537,In_231);
nand U1894 (N_1894,In_637,In_74);
and U1895 (N_1895,In_464,In_201);
nor U1896 (N_1896,In_695,In_590);
or U1897 (N_1897,In_692,In_610);
nand U1898 (N_1898,In_190,In_541);
and U1899 (N_1899,In_577,In_63);
xor U1900 (N_1900,In_214,In_427);
and U1901 (N_1901,In_464,In_379);
and U1902 (N_1902,In_2,In_171);
or U1903 (N_1903,In_187,In_476);
or U1904 (N_1904,In_228,In_535);
nor U1905 (N_1905,In_434,In_45);
and U1906 (N_1906,In_511,In_558);
or U1907 (N_1907,In_200,In_248);
or U1908 (N_1908,In_598,In_326);
and U1909 (N_1909,In_537,In_735);
nor U1910 (N_1910,In_545,In_741);
or U1911 (N_1911,In_42,In_448);
and U1912 (N_1912,In_144,In_257);
and U1913 (N_1913,In_261,In_147);
or U1914 (N_1914,In_439,In_1);
and U1915 (N_1915,In_645,In_462);
nor U1916 (N_1916,In_698,In_485);
and U1917 (N_1917,In_23,In_573);
nand U1918 (N_1918,In_629,In_748);
or U1919 (N_1919,In_267,In_122);
and U1920 (N_1920,In_747,In_606);
nand U1921 (N_1921,In_320,In_53);
nor U1922 (N_1922,In_52,In_459);
and U1923 (N_1923,In_264,In_12);
nand U1924 (N_1924,In_25,In_450);
nand U1925 (N_1925,In_535,In_281);
nand U1926 (N_1926,In_508,In_25);
and U1927 (N_1927,In_263,In_682);
nand U1928 (N_1928,In_691,In_80);
nand U1929 (N_1929,In_697,In_323);
nand U1930 (N_1930,In_475,In_73);
and U1931 (N_1931,In_578,In_352);
nor U1932 (N_1932,In_497,In_366);
or U1933 (N_1933,In_334,In_683);
or U1934 (N_1934,In_60,In_489);
nor U1935 (N_1935,In_476,In_0);
or U1936 (N_1936,In_478,In_644);
nand U1937 (N_1937,In_404,In_99);
nand U1938 (N_1938,In_579,In_744);
nor U1939 (N_1939,In_514,In_165);
or U1940 (N_1940,In_483,In_195);
xnor U1941 (N_1941,In_550,In_289);
or U1942 (N_1942,In_38,In_272);
nand U1943 (N_1943,In_569,In_545);
nor U1944 (N_1944,In_263,In_459);
nor U1945 (N_1945,In_640,In_748);
or U1946 (N_1946,In_405,In_385);
and U1947 (N_1947,In_101,In_74);
and U1948 (N_1948,In_575,In_109);
and U1949 (N_1949,In_74,In_444);
and U1950 (N_1950,In_133,In_455);
nor U1951 (N_1951,In_92,In_134);
and U1952 (N_1952,In_486,In_441);
nand U1953 (N_1953,In_504,In_302);
nor U1954 (N_1954,In_74,In_735);
nor U1955 (N_1955,In_232,In_541);
nor U1956 (N_1956,In_283,In_297);
nand U1957 (N_1957,In_289,In_685);
or U1958 (N_1958,In_650,In_195);
xor U1959 (N_1959,In_183,In_712);
and U1960 (N_1960,In_246,In_373);
and U1961 (N_1961,In_476,In_634);
nand U1962 (N_1962,In_123,In_321);
nand U1963 (N_1963,In_567,In_32);
nand U1964 (N_1964,In_497,In_288);
or U1965 (N_1965,In_141,In_634);
nand U1966 (N_1966,In_458,In_711);
nor U1967 (N_1967,In_202,In_386);
and U1968 (N_1968,In_327,In_680);
and U1969 (N_1969,In_460,In_627);
and U1970 (N_1970,In_600,In_113);
and U1971 (N_1971,In_602,In_667);
and U1972 (N_1972,In_712,In_397);
or U1973 (N_1973,In_514,In_403);
nand U1974 (N_1974,In_117,In_106);
or U1975 (N_1975,In_213,In_598);
nor U1976 (N_1976,In_219,In_225);
and U1977 (N_1977,In_722,In_424);
nand U1978 (N_1978,In_625,In_670);
and U1979 (N_1979,In_674,In_342);
or U1980 (N_1980,In_581,In_421);
nand U1981 (N_1981,In_413,In_691);
nand U1982 (N_1982,In_48,In_211);
nand U1983 (N_1983,In_219,In_527);
or U1984 (N_1984,In_29,In_647);
nand U1985 (N_1985,In_406,In_0);
nand U1986 (N_1986,In_680,In_693);
nor U1987 (N_1987,In_31,In_449);
or U1988 (N_1988,In_722,In_29);
and U1989 (N_1989,In_214,In_685);
nand U1990 (N_1990,In_444,In_314);
nor U1991 (N_1991,In_555,In_25);
nand U1992 (N_1992,In_217,In_79);
and U1993 (N_1993,In_611,In_422);
nand U1994 (N_1994,In_191,In_592);
nor U1995 (N_1995,In_84,In_429);
nand U1996 (N_1996,In_411,In_224);
nor U1997 (N_1997,In_646,In_379);
or U1998 (N_1998,In_508,In_328);
or U1999 (N_1999,In_686,In_656);
nor U2000 (N_2000,In_182,In_72);
and U2001 (N_2001,In_672,In_36);
nand U2002 (N_2002,In_146,In_239);
nor U2003 (N_2003,In_483,In_579);
and U2004 (N_2004,In_555,In_398);
nor U2005 (N_2005,In_691,In_696);
and U2006 (N_2006,In_443,In_458);
or U2007 (N_2007,In_519,In_97);
or U2008 (N_2008,In_535,In_264);
xnor U2009 (N_2009,In_345,In_736);
nand U2010 (N_2010,In_83,In_341);
and U2011 (N_2011,In_744,In_67);
and U2012 (N_2012,In_11,In_582);
nand U2013 (N_2013,In_280,In_62);
nor U2014 (N_2014,In_245,In_666);
or U2015 (N_2015,In_99,In_555);
or U2016 (N_2016,In_644,In_548);
nand U2017 (N_2017,In_419,In_100);
or U2018 (N_2018,In_41,In_521);
nand U2019 (N_2019,In_159,In_482);
or U2020 (N_2020,In_611,In_497);
nand U2021 (N_2021,In_178,In_381);
and U2022 (N_2022,In_518,In_444);
xor U2023 (N_2023,In_175,In_144);
nand U2024 (N_2024,In_286,In_544);
nor U2025 (N_2025,In_688,In_615);
and U2026 (N_2026,In_18,In_693);
or U2027 (N_2027,In_359,In_686);
nand U2028 (N_2028,In_733,In_4);
nor U2029 (N_2029,In_30,In_445);
or U2030 (N_2030,In_497,In_491);
and U2031 (N_2031,In_447,In_649);
or U2032 (N_2032,In_550,In_240);
or U2033 (N_2033,In_454,In_404);
or U2034 (N_2034,In_243,In_420);
nor U2035 (N_2035,In_548,In_83);
nor U2036 (N_2036,In_331,In_90);
nor U2037 (N_2037,In_200,In_380);
nand U2038 (N_2038,In_313,In_140);
nand U2039 (N_2039,In_360,In_266);
or U2040 (N_2040,In_248,In_553);
nand U2041 (N_2041,In_481,In_258);
nor U2042 (N_2042,In_307,In_92);
and U2043 (N_2043,In_402,In_702);
or U2044 (N_2044,In_390,In_492);
and U2045 (N_2045,In_161,In_381);
and U2046 (N_2046,In_23,In_321);
and U2047 (N_2047,In_728,In_340);
or U2048 (N_2048,In_636,In_447);
or U2049 (N_2049,In_412,In_523);
nand U2050 (N_2050,In_699,In_232);
nor U2051 (N_2051,In_237,In_105);
nand U2052 (N_2052,In_391,In_173);
or U2053 (N_2053,In_553,In_177);
nand U2054 (N_2054,In_681,In_489);
and U2055 (N_2055,In_741,In_462);
or U2056 (N_2056,In_629,In_167);
and U2057 (N_2057,In_259,In_433);
or U2058 (N_2058,In_322,In_450);
or U2059 (N_2059,In_172,In_505);
or U2060 (N_2060,In_170,In_82);
nor U2061 (N_2061,In_109,In_301);
nand U2062 (N_2062,In_176,In_667);
or U2063 (N_2063,In_536,In_126);
and U2064 (N_2064,In_309,In_494);
nor U2065 (N_2065,In_103,In_703);
and U2066 (N_2066,In_356,In_468);
or U2067 (N_2067,In_410,In_577);
or U2068 (N_2068,In_479,In_747);
nand U2069 (N_2069,In_67,In_669);
nor U2070 (N_2070,In_236,In_239);
and U2071 (N_2071,In_385,In_665);
or U2072 (N_2072,In_397,In_270);
or U2073 (N_2073,In_654,In_525);
or U2074 (N_2074,In_356,In_401);
or U2075 (N_2075,In_3,In_128);
nand U2076 (N_2076,In_28,In_353);
nand U2077 (N_2077,In_113,In_628);
nand U2078 (N_2078,In_391,In_590);
nor U2079 (N_2079,In_605,In_432);
nor U2080 (N_2080,In_408,In_724);
or U2081 (N_2081,In_287,In_362);
or U2082 (N_2082,In_324,In_623);
xnor U2083 (N_2083,In_601,In_174);
nand U2084 (N_2084,In_254,In_61);
or U2085 (N_2085,In_637,In_361);
nor U2086 (N_2086,In_499,In_91);
or U2087 (N_2087,In_352,In_574);
nand U2088 (N_2088,In_198,In_447);
nor U2089 (N_2089,In_329,In_417);
nor U2090 (N_2090,In_44,In_163);
nand U2091 (N_2091,In_178,In_583);
nor U2092 (N_2092,In_149,In_284);
xnor U2093 (N_2093,In_193,In_136);
or U2094 (N_2094,In_598,In_183);
and U2095 (N_2095,In_77,In_297);
nor U2096 (N_2096,In_213,In_732);
nor U2097 (N_2097,In_351,In_385);
and U2098 (N_2098,In_619,In_437);
or U2099 (N_2099,In_730,In_260);
or U2100 (N_2100,In_360,In_335);
nor U2101 (N_2101,In_57,In_683);
or U2102 (N_2102,In_111,In_262);
or U2103 (N_2103,In_706,In_651);
nand U2104 (N_2104,In_238,In_391);
and U2105 (N_2105,In_507,In_743);
and U2106 (N_2106,In_742,In_121);
or U2107 (N_2107,In_615,In_479);
or U2108 (N_2108,In_367,In_102);
nand U2109 (N_2109,In_480,In_344);
nor U2110 (N_2110,In_644,In_402);
nor U2111 (N_2111,In_717,In_21);
nor U2112 (N_2112,In_239,In_422);
or U2113 (N_2113,In_722,In_535);
nand U2114 (N_2114,In_351,In_584);
and U2115 (N_2115,In_103,In_585);
nand U2116 (N_2116,In_332,In_276);
and U2117 (N_2117,In_409,In_263);
nand U2118 (N_2118,In_667,In_647);
or U2119 (N_2119,In_646,In_636);
nand U2120 (N_2120,In_549,In_679);
nor U2121 (N_2121,In_27,In_538);
nor U2122 (N_2122,In_724,In_334);
nor U2123 (N_2123,In_571,In_12);
or U2124 (N_2124,In_587,In_88);
nor U2125 (N_2125,In_417,In_79);
nor U2126 (N_2126,In_519,In_556);
nand U2127 (N_2127,In_60,In_443);
nand U2128 (N_2128,In_92,In_691);
nor U2129 (N_2129,In_129,In_107);
nand U2130 (N_2130,In_536,In_741);
or U2131 (N_2131,In_492,In_63);
nand U2132 (N_2132,In_666,In_578);
and U2133 (N_2133,In_128,In_669);
or U2134 (N_2134,In_291,In_87);
and U2135 (N_2135,In_268,In_449);
nor U2136 (N_2136,In_173,In_413);
nand U2137 (N_2137,In_296,In_211);
nor U2138 (N_2138,In_87,In_269);
and U2139 (N_2139,In_27,In_698);
nand U2140 (N_2140,In_233,In_567);
nor U2141 (N_2141,In_304,In_9);
and U2142 (N_2142,In_151,In_711);
or U2143 (N_2143,In_276,In_716);
nor U2144 (N_2144,In_242,In_170);
or U2145 (N_2145,In_219,In_213);
nor U2146 (N_2146,In_365,In_84);
nand U2147 (N_2147,In_524,In_605);
xnor U2148 (N_2148,In_36,In_688);
nor U2149 (N_2149,In_429,In_687);
nand U2150 (N_2150,In_51,In_445);
nor U2151 (N_2151,In_212,In_447);
and U2152 (N_2152,In_601,In_729);
and U2153 (N_2153,In_18,In_110);
xnor U2154 (N_2154,In_567,In_242);
nor U2155 (N_2155,In_357,In_521);
nor U2156 (N_2156,In_560,In_722);
nor U2157 (N_2157,In_320,In_567);
and U2158 (N_2158,In_154,In_393);
nand U2159 (N_2159,In_517,In_495);
nand U2160 (N_2160,In_560,In_83);
nand U2161 (N_2161,In_490,In_113);
nor U2162 (N_2162,In_678,In_305);
nor U2163 (N_2163,In_713,In_362);
xor U2164 (N_2164,In_705,In_155);
nand U2165 (N_2165,In_369,In_565);
nor U2166 (N_2166,In_231,In_151);
and U2167 (N_2167,In_697,In_502);
or U2168 (N_2168,In_355,In_528);
nand U2169 (N_2169,In_444,In_305);
or U2170 (N_2170,In_435,In_425);
nand U2171 (N_2171,In_104,In_399);
and U2172 (N_2172,In_88,In_181);
and U2173 (N_2173,In_398,In_644);
nand U2174 (N_2174,In_592,In_703);
nor U2175 (N_2175,In_360,In_176);
nor U2176 (N_2176,In_473,In_343);
nand U2177 (N_2177,In_112,In_495);
nor U2178 (N_2178,In_388,In_238);
and U2179 (N_2179,In_238,In_659);
or U2180 (N_2180,In_125,In_183);
or U2181 (N_2181,In_687,In_142);
nor U2182 (N_2182,In_342,In_477);
and U2183 (N_2183,In_482,In_536);
or U2184 (N_2184,In_294,In_657);
nand U2185 (N_2185,In_376,In_215);
nor U2186 (N_2186,In_727,In_342);
nand U2187 (N_2187,In_390,In_653);
and U2188 (N_2188,In_674,In_507);
or U2189 (N_2189,In_114,In_359);
or U2190 (N_2190,In_666,In_698);
nor U2191 (N_2191,In_426,In_249);
and U2192 (N_2192,In_671,In_94);
nor U2193 (N_2193,In_301,In_159);
or U2194 (N_2194,In_532,In_24);
or U2195 (N_2195,In_701,In_381);
or U2196 (N_2196,In_9,In_670);
nand U2197 (N_2197,In_10,In_156);
and U2198 (N_2198,In_555,In_625);
and U2199 (N_2199,In_107,In_92);
or U2200 (N_2200,In_488,In_88);
or U2201 (N_2201,In_348,In_134);
nand U2202 (N_2202,In_472,In_244);
nor U2203 (N_2203,In_468,In_15);
nand U2204 (N_2204,In_359,In_696);
nand U2205 (N_2205,In_231,In_396);
nand U2206 (N_2206,In_144,In_212);
nor U2207 (N_2207,In_321,In_402);
or U2208 (N_2208,In_154,In_15);
or U2209 (N_2209,In_603,In_241);
and U2210 (N_2210,In_396,In_623);
nor U2211 (N_2211,In_94,In_597);
xor U2212 (N_2212,In_230,In_324);
or U2213 (N_2213,In_736,In_645);
or U2214 (N_2214,In_352,In_176);
or U2215 (N_2215,In_434,In_77);
and U2216 (N_2216,In_362,In_62);
or U2217 (N_2217,In_276,In_90);
and U2218 (N_2218,In_661,In_258);
nand U2219 (N_2219,In_279,In_544);
and U2220 (N_2220,In_649,In_555);
nand U2221 (N_2221,In_402,In_101);
nor U2222 (N_2222,In_354,In_246);
nor U2223 (N_2223,In_94,In_236);
nand U2224 (N_2224,In_442,In_328);
nor U2225 (N_2225,In_125,In_651);
and U2226 (N_2226,In_418,In_367);
and U2227 (N_2227,In_549,In_623);
or U2228 (N_2228,In_104,In_267);
nor U2229 (N_2229,In_730,In_77);
xnor U2230 (N_2230,In_368,In_350);
nand U2231 (N_2231,In_129,In_178);
nor U2232 (N_2232,In_140,In_562);
nor U2233 (N_2233,In_508,In_515);
nand U2234 (N_2234,In_79,In_663);
and U2235 (N_2235,In_193,In_76);
and U2236 (N_2236,In_162,In_715);
nor U2237 (N_2237,In_402,In_198);
or U2238 (N_2238,In_567,In_296);
and U2239 (N_2239,In_576,In_336);
or U2240 (N_2240,In_724,In_145);
or U2241 (N_2241,In_491,In_182);
nor U2242 (N_2242,In_79,In_402);
nor U2243 (N_2243,In_189,In_76);
or U2244 (N_2244,In_228,In_722);
and U2245 (N_2245,In_68,In_273);
and U2246 (N_2246,In_216,In_667);
nor U2247 (N_2247,In_720,In_127);
or U2248 (N_2248,In_410,In_460);
nor U2249 (N_2249,In_70,In_738);
nor U2250 (N_2250,In_369,In_341);
and U2251 (N_2251,In_275,In_305);
and U2252 (N_2252,In_525,In_500);
nor U2253 (N_2253,In_142,In_238);
or U2254 (N_2254,In_157,In_223);
or U2255 (N_2255,In_484,In_94);
nand U2256 (N_2256,In_124,In_63);
nor U2257 (N_2257,In_430,In_575);
nor U2258 (N_2258,In_522,In_749);
nor U2259 (N_2259,In_317,In_158);
or U2260 (N_2260,In_607,In_373);
and U2261 (N_2261,In_84,In_54);
or U2262 (N_2262,In_239,In_187);
and U2263 (N_2263,In_556,In_620);
nor U2264 (N_2264,In_402,In_459);
and U2265 (N_2265,In_277,In_351);
nand U2266 (N_2266,In_436,In_532);
nor U2267 (N_2267,In_52,In_193);
or U2268 (N_2268,In_452,In_38);
or U2269 (N_2269,In_446,In_535);
or U2270 (N_2270,In_731,In_530);
nand U2271 (N_2271,In_119,In_496);
and U2272 (N_2272,In_392,In_445);
nor U2273 (N_2273,In_477,In_225);
nand U2274 (N_2274,In_347,In_487);
nand U2275 (N_2275,In_420,In_306);
and U2276 (N_2276,In_656,In_328);
nor U2277 (N_2277,In_292,In_444);
and U2278 (N_2278,In_718,In_299);
or U2279 (N_2279,In_695,In_167);
or U2280 (N_2280,In_632,In_106);
and U2281 (N_2281,In_68,In_640);
or U2282 (N_2282,In_566,In_197);
and U2283 (N_2283,In_296,In_665);
and U2284 (N_2284,In_149,In_544);
or U2285 (N_2285,In_675,In_45);
nand U2286 (N_2286,In_38,In_456);
nor U2287 (N_2287,In_88,In_396);
or U2288 (N_2288,In_312,In_164);
nor U2289 (N_2289,In_163,In_679);
nand U2290 (N_2290,In_578,In_585);
nand U2291 (N_2291,In_251,In_142);
or U2292 (N_2292,In_721,In_492);
nor U2293 (N_2293,In_162,In_431);
or U2294 (N_2294,In_536,In_101);
nand U2295 (N_2295,In_57,In_336);
and U2296 (N_2296,In_519,In_135);
and U2297 (N_2297,In_449,In_376);
or U2298 (N_2298,In_92,In_93);
and U2299 (N_2299,In_461,In_746);
nand U2300 (N_2300,In_704,In_300);
nand U2301 (N_2301,In_395,In_311);
or U2302 (N_2302,In_726,In_188);
and U2303 (N_2303,In_271,In_349);
nand U2304 (N_2304,In_703,In_72);
nand U2305 (N_2305,In_345,In_740);
and U2306 (N_2306,In_382,In_17);
or U2307 (N_2307,In_313,In_555);
nor U2308 (N_2308,In_146,In_486);
and U2309 (N_2309,In_107,In_119);
or U2310 (N_2310,In_52,In_671);
and U2311 (N_2311,In_115,In_328);
nand U2312 (N_2312,In_543,In_735);
and U2313 (N_2313,In_7,In_598);
or U2314 (N_2314,In_338,In_71);
and U2315 (N_2315,In_729,In_507);
nand U2316 (N_2316,In_677,In_448);
nor U2317 (N_2317,In_471,In_129);
and U2318 (N_2318,In_708,In_592);
nand U2319 (N_2319,In_1,In_2);
nor U2320 (N_2320,In_65,In_130);
nor U2321 (N_2321,In_45,In_451);
xnor U2322 (N_2322,In_367,In_466);
nand U2323 (N_2323,In_218,In_477);
nor U2324 (N_2324,In_351,In_243);
nand U2325 (N_2325,In_637,In_301);
and U2326 (N_2326,In_481,In_748);
or U2327 (N_2327,In_558,In_688);
or U2328 (N_2328,In_128,In_158);
or U2329 (N_2329,In_427,In_18);
and U2330 (N_2330,In_587,In_1);
and U2331 (N_2331,In_636,In_29);
and U2332 (N_2332,In_256,In_622);
and U2333 (N_2333,In_496,In_263);
or U2334 (N_2334,In_676,In_570);
or U2335 (N_2335,In_103,In_241);
nor U2336 (N_2336,In_389,In_653);
nor U2337 (N_2337,In_220,In_633);
and U2338 (N_2338,In_34,In_627);
and U2339 (N_2339,In_89,In_558);
and U2340 (N_2340,In_241,In_348);
and U2341 (N_2341,In_628,In_272);
or U2342 (N_2342,In_550,In_345);
and U2343 (N_2343,In_729,In_234);
nor U2344 (N_2344,In_349,In_141);
nand U2345 (N_2345,In_268,In_299);
and U2346 (N_2346,In_341,In_453);
nand U2347 (N_2347,In_452,In_454);
nor U2348 (N_2348,In_416,In_37);
nand U2349 (N_2349,In_560,In_103);
nor U2350 (N_2350,In_64,In_422);
or U2351 (N_2351,In_262,In_576);
nor U2352 (N_2352,In_176,In_380);
nor U2353 (N_2353,In_671,In_358);
nor U2354 (N_2354,In_492,In_269);
nand U2355 (N_2355,In_240,In_42);
nand U2356 (N_2356,In_162,In_262);
nor U2357 (N_2357,In_302,In_314);
and U2358 (N_2358,In_565,In_264);
nand U2359 (N_2359,In_317,In_296);
nand U2360 (N_2360,In_475,In_672);
and U2361 (N_2361,In_702,In_196);
or U2362 (N_2362,In_128,In_256);
and U2363 (N_2363,In_595,In_138);
nor U2364 (N_2364,In_684,In_109);
and U2365 (N_2365,In_386,In_169);
nor U2366 (N_2366,In_672,In_332);
nor U2367 (N_2367,In_198,In_91);
or U2368 (N_2368,In_192,In_394);
or U2369 (N_2369,In_735,In_672);
nand U2370 (N_2370,In_108,In_335);
nand U2371 (N_2371,In_237,In_181);
nand U2372 (N_2372,In_13,In_234);
or U2373 (N_2373,In_641,In_659);
or U2374 (N_2374,In_559,In_663);
nor U2375 (N_2375,In_65,In_698);
or U2376 (N_2376,In_247,In_240);
or U2377 (N_2377,In_164,In_711);
nor U2378 (N_2378,In_78,In_430);
nand U2379 (N_2379,In_106,In_364);
nand U2380 (N_2380,In_448,In_96);
nand U2381 (N_2381,In_531,In_405);
or U2382 (N_2382,In_170,In_277);
or U2383 (N_2383,In_568,In_663);
and U2384 (N_2384,In_450,In_560);
nor U2385 (N_2385,In_704,In_645);
or U2386 (N_2386,In_123,In_569);
nor U2387 (N_2387,In_24,In_631);
xnor U2388 (N_2388,In_529,In_506);
and U2389 (N_2389,In_404,In_51);
nand U2390 (N_2390,In_208,In_201);
and U2391 (N_2391,In_251,In_272);
and U2392 (N_2392,In_120,In_91);
or U2393 (N_2393,In_32,In_368);
nand U2394 (N_2394,In_703,In_339);
nor U2395 (N_2395,In_1,In_476);
and U2396 (N_2396,In_6,In_691);
nor U2397 (N_2397,In_576,In_257);
xor U2398 (N_2398,In_426,In_477);
xnor U2399 (N_2399,In_101,In_542);
nand U2400 (N_2400,In_673,In_270);
nand U2401 (N_2401,In_329,In_229);
xnor U2402 (N_2402,In_541,In_392);
nand U2403 (N_2403,In_310,In_270);
and U2404 (N_2404,In_272,In_319);
and U2405 (N_2405,In_707,In_161);
nand U2406 (N_2406,In_383,In_320);
nor U2407 (N_2407,In_302,In_163);
nand U2408 (N_2408,In_621,In_542);
and U2409 (N_2409,In_428,In_736);
and U2410 (N_2410,In_59,In_279);
nand U2411 (N_2411,In_507,In_443);
and U2412 (N_2412,In_541,In_137);
or U2413 (N_2413,In_586,In_274);
and U2414 (N_2414,In_322,In_315);
nor U2415 (N_2415,In_182,In_640);
nor U2416 (N_2416,In_164,In_558);
nor U2417 (N_2417,In_506,In_277);
or U2418 (N_2418,In_180,In_602);
nand U2419 (N_2419,In_201,In_407);
and U2420 (N_2420,In_546,In_163);
nand U2421 (N_2421,In_238,In_104);
and U2422 (N_2422,In_384,In_366);
and U2423 (N_2423,In_333,In_150);
nor U2424 (N_2424,In_103,In_741);
nor U2425 (N_2425,In_174,In_218);
nor U2426 (N_2426,In_617,In_461);
nor U2427 (N_2427,In_546,In_700);
and U2428 (N_2428,In_398,In_298);
or U2429 (N_2429,In_337,In_602);
nand U2430 (N_2430,In_303,In_218);
nor U2431 (N_2431,In_154,In_688);
nor U2432 (N_2432,In_315,In_606);
nor U2433 (N_2433,In_259,In_449);
nor U2434 (N_2434,In_221,In_194);
nand U2435 (N_2435,In_465,In_614);
nand U2436 (N_2436,In_311,In_476);
nor U2437 (N_2437,In_535,In_555);
and U2438 (N_2438,In_486,In_74);
and U2439 (N_2439,In_286,In_237);
xnor U2440 (N_2440,In_595,In_402);
and U2441 (N_2441,In_433,In_169);
nor U2442 (N_2442,In_520,In_242);
nor U2443 (N_2443,In_734,In_271);
nand U2444 (N_2444,In_98,In_73);
or U2445 (N_2445,In_621,In_441);
or U2446 (N_2446,In_532,In_165);
and U2447 (N_2447,In_504,In_633);
nand U2448 (N_2448,In_285,In_522);
or U2449 (N_2449,In_575,In_724);
or U2450 (N_2450,In_251,In_58);
and U2451 (N_2451,In_60,In_194);
and U2452 (N_2452,In_203,In_260);
and U2453 (N_2453,In_413,In_484);
and U2454 (N_2454,In_443,In_483);
nand U2455 (N_2455,In_82,In_485);
nor U2456 (N_2456,In_400,In_306);
nor U2457 (N_2457,In_255,In_710);
nand U2458 (N_2458,In_532,In_413);
or U2459 (N_2459,In_324,In_443);
and U2460 (N_2460,In_371,In_301);
or U2461 (N_2461,In_264,In_337);
nand U2462 (N_2462,In_22,In_745);
nor U2463 (N_2463,In_200,In_267);
and U2464 (N_2464,In_196,In_393);
and U2465 (N_2465,In_203,In_207);
and U2466 (N_2466,In_574,In_536);
and U2467 (N_2467,In_213,In_460);
or U2468 (N_2468,In_162,In_697);
and U2469 (N_2469,In_381,In_724);
and U2470 (N_2470,In_612,In_206);
or U2471 (N_2471,In_635,In_662);
nand U2472 (N_2472,In_209,In_507);
and U2473 (N_2473,In_712,In_421);
nor U2474 (N_2474,In_541,In_248);
or U2475 (N_2475,In_593,In_363);
nand U2476 (N_2476,In_447,In_1);
nor U2477 (N_2477,In_286,In_404);
or U2478 (N_2478,In_328,In_36);
nor U2479 (N_2479,In_662,In_472);
and U2480 (N_2480,In_99,In_429);
or U2481 (N_2481,In_206,In_448);
and U2482 (N_2482,In_736,In_459);
and U2483 (N_2483,In_389,In_228);
and U2484 (N_2484,In_84,In_472);
nor U2485 (N_2485,In_41,In_169);
nor U2486 (N_2486,In_668,In_398);
or U2487 (N_2487,In_404,In_10);
and U2488 (N_2488,In_81,In_632);
or U2489 (N_2489,In_156,In_585);
nand U2490 (N_2490,In_529,In_66);
and U2491 (N_2491,In_587,In_256);
nand U2492 (N_2492,In_41,In_469);
nand U2493 (N_2493,In_97,In_572);
or U2494 (N_2494,In_437,In_429);
nor U2495 (N_2495,In_581,In_185);
and U2496 (N_2496,In_97,In_93);
nor U2497 (N_2497,In_212,In_506);
and U2498 (N_2498,In_339,In_618);
and U2499 (N_2499,In_355,In_191);
nand U2500 (N_2500,N_1583,N_2058);
and U2501 (N_2501,N_1603,N_499);
nand U2502 (N_2502,N_424,N_1270);
and U2503 (N_2503,N_1610,N_1456);
nand U2504 (N_2504,N_482,N_1068);
and U2505 (N_2505,N_626,N_1189);
or U2506 (N_2506,N_561,N_1835);
and U2507 (N_2507,N_584,N_743);
and U2508 (N_2508,N_2062,N_104);
nor U2509 (N_2509,N_2098,N_2313);
nor U2510 (N_2510,N_2239,N_659);
nand U2511 (N_2511,N_2064,N_1787);
or U2512 (N_2512,N_2006,N_1634);
nand U2513 (N_2513,N_420,N_2179);
and U2514 (N_2514,N_1544,N_2379);
nor U2515 (N_2515,N_2213,N_1993);
nor U2516 (N_2516,N_399,N_284);
and U2517 (N_2517,N_1744,N_2207);
nand U2518 (N_2518,N_877,N_277);
nand U2519 (N_2519,N_968,N_994);
nor U2520 (N_2520,N_1662,N_899);
nand U2521 (N_2521,N_1171,N_814);
nand U2522 (N_2522,N_171,N_1065);
nand U2523 (N_2523,N_1460,N_2496);
and U2524 (N_2524,N_738,N_2381);
xnor U2525 (N_2525,N_956,N_1176);
nor U2526 (N_2526,N_1138,N_106);
and U2527 (N_2527,N_1037,N_886);
xor U2528 (N_2528,N_2145,N_2216);
or U2529 (N_2529,N_176,N_250);
or U2530 (N_2530,N_68,N_2320);
nand U2531 (N_2531,N_1987,N_359);
or U2532 (N_2532,N_1367,N_1087);
nor U2533 (N_2533,N_1584,N_2197);
nand U2534 (N_2534,N_85,N_1889);
and U2535 (N_2535,N_2488,N_1243);
nor U2536 (N_2536,N_564,N_1130);
and U2537 (N_2537,N_1311,N_1006);
and U2538 (N_2538,N_973,N_531);
or U2539 (N_2539,N_1939,N_2270);
nand U2540 (N_2540,N_412,N_251);
and U2541 (N_2541,N_1286,N_1640);
or U2542 (N_2542,N_1979,N_2417);
nor U2543 (N_2543,N_1907,N_1041);
nor U2544 (N_2544,N_475,N_1962);
xor U2545 (N_2545,N_2302,N_1101);
and U2546 (N_2546,N_1660,N_1415);
nor U2547 (N_2547,N_2383,N_1362);
and U2548 (N_2548,N_1129,N_282);
nand U2549 (N_2549,N_1970,N_808);
and U2550 (N_2550,N_901,N_1025);
and U2551 (N_2551,N_711,N_1615);
nand U2552 (N_2552,N_1066,N_1566);
and U2553 (N_2553,N_1693,N_850);
and U2554 (N_2554,N_800,N_918);
or U2555 (N_2555,N_644,N_1128);
xnor U2556 (N_2556,N_893,N_461);
or U2557 (N_2557,N_386,N_1153);
or U2558 (N_2558,N_989,N_2156);
or U2559 (N_2559,N_241,N_1964);
and U2560 (N_2560,N_322,N_2415);
or U2561 (N_2561,N_2273,N_1611);
nor U2562 (N_2562,N_366,N_89);
nand U2563 (N_2563,N_1416,N_462);
nor U2564 (N_2564,N_2146,N_74);
nor U2565 (N_2565,N_343,N_970);
or U2566 (N_2566,N_1118,N_33);
and U2567 (N_2567,N_2253,N_831);
and U2568 (N_2568,N_1972,N_380);
nand U2569 (N_2569,N_78,N_1912);
and U2570 (N_2570,N_656,N_1717);
nor U2571 (N_2571,N_141,N_2209);
nor U2572 (N_2572,N_10,N_596);
or U2573 (N_2573,N_1304,N_1440);
or U2574 (N_2574,N_1312,N_1960);
nand U2575 (N_2575,N_1856,N_15);
xnor U2576 (N_2576,N_330,N_1436);
nor U2577 (N_2577,N_560,N_1223);
or U2578 (N_2578,N_164,N_221);
or U2579 (N_2579,N_2188,N_1982);
nor U2580 (N_2580,N_629,N_375);
or U2581 (N_2581,N_1809,N_1511);
or U2582 (N_2582,N_1620,N_1317);
or U2583 (N_2583,N_1748,N_1371);
nor U2584 (N_2584,N_1350,N_707);
nor U2585 (N_2585,N_356,N_1886);
or U2586 (N_2586,N_946,N_1810);
or U2587 (N_2587,N_126,N_1871);
nand U2588 (N_2588,N_1276,N_2404);
and U2589 (N_2589,N_2217,N_2106);
nand U2590 (N_2590,N_722,N_2051);
or U2591 (N_2591,N_640,N_1327);
and U2592 (N_2592,N_333,N_1149);
nor U2593 (N_2593,N_1109,N_2314);
nor U2594 (N_2594,N_1758,N_37);
or U2595 (N_2595,N_919,N_2305);
and U2596 (N_2596,N_812,N_134);
nand U2597 (N_2597,N_1769,N_194);
or U2598 (N_2598,N_617,N_1648);
or U2599 (N_2599,N_609,N_641);
nor U2600 (N_2600,N_2203,N_2167);
nand U2601 (N_2601,N_1530,N_2200);
and U2602 (N_2602,N_813,N_950);
and U2603 (N_2603,N_1088,N_1876);
or U2604 (N_2604,N_486,N_2294);
nor U2605 (N_2605,N_1731,N_572);
nand U2606 (N_2606,N_27,N_1576);
and U2607 (N_2607,N_2353,N_1759);
and U2608 (N_2608,N_1201,N_1913);
nand U2609 (N_2609,N_2390,N_1490);
nand U2610 (N_2610,N_2159,N_2067);
or U2611 (N_2611,N_295,N_763);
nand U2612 (N_2612,N_1542,N_487);
nor U2613 (N_2613,N_70,N_2070);
and U2614 (N_2614,N_2412,N_771);
nand U2615 (N_2615,N_205,N_5);
nand U2616 (N_2616,N_1600,N_1637);
or U2617 (N_2617,N_2277,N_1442);
nand U2618 (N_2618,N_1794,N_1654);
or U2619 (N_2619,N_464,N_1638);
nor U2620 (N_2620,N_480,N_1707);
nand U2621 (N_2621,N_1710,N_987);
nor U2622 (N_2622,N_2164,N_1392);
nand U2623 (N_2623,N_1,N_1523);
nand U2624 (N_2624,N_1299,N_577);
and U2625 (N_2625,N_1822,N_2123);
nor U2626 (N_2626,N_2369,N_1963);
nand U2627 (N_2627,N_2367,N_1625);
or U2628 (N_2628,N_1277,N_2074);
and U2629 (N_2629,N_667,N_1154);
and U2630 (N_2630,N_1612,N_600);
xnor U2631 (N_2631,N_1696,N_972);
nor U2632 (N_2632,N_892,N_8);
nand U2633 (N_2633,N_118,N_2225);
and U2634 (N_2634,N_95,N_1784);
nand U2635 (N_2635,N_1080,N_309);
or U2636 (N_2636,N_1084,N_1102);
nand U2637 (N_2637,N_9,N_1040);
or U2638 (N_2638,N_344,N_2174);
nor U2639 (N_2639,N_1909,N_730);
nand U2640 (N_2640,N_1191,N_844);
nor U2641 (N_2641,N_2433,N_1679);
nand U2642 (N_2642,N_780,N_422);
or U2643 (N_2643,N_1018,N_1527);
and U2644 (N_2644,N_231,N_222);
nand U2645 (N_2645,N_1984,N_1157);
nor U2646 (N_2646,N_138,N_1977);
nand U2647 (N_2647,N_910,N_1297);
nor U2648 (N_2648,N_2312,N_2068);
or U2649 (N_2649,N_1994,N_2427);
nor U2650 (N_2650,N_80,N_2300);
and U2651 (N_2651,N_1023,N_1681);
nand U2652 (N_2652,N_1198,N_1165);
or U2653 (N_2653,N_1205,N_2389);
nand U2654 (N_2654,N_155,N_1287);
nand U2655 (N_2655,N_1757,N_1378);
and U2656 (N_2656,N_902,N_975);
and U2657 (N_2657,N_492,N_1838);
or U2658 (N_2658,N_1282,N_56);
or U2659 (N_2659,N_1407,N_71);
and U2660 (N_2660,N_2194,N_455);
and U2661 (N_2661,N_540,N_862);
nor U2662 (N_2662,N_201,N_1894);
or U2663 (N_2663,N_174,N_2482);
and U2664 (N_2664,N_308,N_2298);
or U2665 (N_2665,N_606,N_2227);
nor U2666 (N_2666,N_2185,N_206);
and U2667 (N_2667,N_2032,N_669);
and U2668 (N_2668,N_558,N_1001);
and U2669 (N_2669,N_2272,N_2116);
and U2670 (N_2670,N_1800,N_1581);
nor U2671 (N_2671,N_2103,N_127);
and U2672 (N_2672,N_1035,N_1055);
and U2673 (N_2673,N_2307,N_1699);
and U2674 (N_2674,N_782,N_2316);
nand U2675 (N_2675,N_1903,N_2475);
or U2676 (N_2676,N_934,N_2398);
and U2677 (N_2677,N_587,N_2303);
or U2678 (N_2678,N_2291,N_2025);
nor U2679 (N_2679,N_2285,N_220);
and U2680 (N_2680,N_675,N_2345);
nor U2681 (N_2681,N_1403,N_1691);
nand U2682 (N_2682,N_636,N_2063);
nand U2683 (N_2683,N_1418,N_1202);
or U2684 (N_2684,N_2301,N_1275);
nand U2685 (N_2685,N_650,N_2124);
nor U2686 (N_2686,N_1424,N_1390);
nand U2687 (N_2687,N_2454,N_1877);
or U2688 (N_2688,N_1158,N_974);
and U2689 (N_2689,N_395,N_1649);
and U2690 (N_2690,N_2204,N_2241);
or U2691 (N_2691,N_1308,N_1496);
and U2692 (N_2692,N_1597,N_988);
nor U2693 (N_2693,N_215,N_755);
nor U2694 (N_2694,N_2045,N_815);
xnor U2695 (N_2695,N_1150,N_554);
and U2696 (N_2696,N_1184,N_1578);
or U2697 (N_2697,N_1229,N_1830);
and U2698 (N_2698,N_2077,N_903);
and U2699 (N_2699,N_1135,N_1756);
or U2700 (N_2700,N_130,N_2340);
and U2701 (N_2701,N_1177,N_1688);
xor U2702 (N_2702,N_1193,N_754);
or U2703 (N_2703,N_326,N_105);
or U2704 (N_2704,N_776,N_2292);
nand U2705 (N_2705,N_52,N_668);
and U2706 (N_2706,N_1968,N_2112);
and U2707 (N_2707,N_821,N_1535);
nand U2708 (N_2708,N_1412,N_2118);
and U2709 (N_2709,N_474,N_225);
and U2710 (N_2710,N_2085,N_188);
or U2711 (N_2711,N_2350,N_1561);
nor U2712 (N_2712,N_746,N_2288);
nor U2713 (N_2713,N_865,N_279);
nor U2714 (N_2714,N_2341,N_436);
nor U2715 (N_2715,N_2261,N_240);
nand U2716 (N_2716,N_2015,N_116);
or U2717 (N_2717,N_1241,N_278);
xnor U2718 (N_2718,N_2009,N_1899);
nor U2719 (N_2719,N_643,N_2342);
nor U2720 (N_2720,N_751,N_2022);
or U2721 (N_2721,N_1338,N_817);
nor U2722 (N_2722,N_2053,N_1030);
or U2723 (N_2723,N_1861,N_411);
or U2724 (N_2724,N_2352,N_55);
or U2725 (N_2725,N_242,N_2128);
or U2726 (N_2726,N_2095,N_2311);
and U2727 (N_2727,N_556,N_550);
nor U2728 (N_2728,N_2040,N_598);
or U2729 (N_2729,N_1017,N_1958);
or U2730 (N_2730,N_539,N_1720);
and U2731 (N_2731,N_819,N_2306);
nor U2732 (N_2732,N_1828,N_1268);
nor U2733 (N_2733,N_3,N_1341);
nor U2734 (N_2734,N_1079,N_1140);
nor U2735 (N_2735,N_2446,N_1665);
xor U2736 (N_2736,N_1428,N_1827);
and U2737 (N_2737,N_2013,N_161);
and U2738 (N_2738,N_1917,N_36);
nor U2739 (N_2739,N_1602,N_1770);
xnor U2740 (N_2740,N_1879,N_545);
nand U2741 (N_2741,N_1112,N_793);
nor U2742 (N_2742,N_2109,N_1022);
or U2743 (N_2743,N_926,N_38);
nor U2744 (N_2744,N_2406,N_1747);
nor U2745 (N_2745,N_81,N_1186);
and U2746 (N_2746,N_704,N_1959);
and U2747 (N_2747,N_158,N_719);
and U2748 (N_2748,N_849,N_619);
or U2749 (N_2749,N_2104,N_1237);
nor U2750 (N_2750,N_1045,N_2376);
nand U2751 (N_2751,N_1740,N_2466);
nor U2752 (N_2752,N_1499,N_752);
nor U2753 (N_2753,N_506,N_964);
and U2754 (N_2754,N_1393,N_2430);
and U2755 (N_2755,N_2082,N_1855);
and U2756 (N_2756,N_1567,N_1595);
nand U2757 (N_2757,N_1501,N_1207);
or U2758 (N_2758,N_1726,N_1589);
and U2759 (N_2759,N_288,N_652);
or U2760 (N_2760,N_1441,N_228);
nand U2761 (N_2761,N_2418,N_1547);
nand U2762 (N_2762,N_1840,N_2337);
nor U2763 (N_2763,N_287,N_1950);
nor U2764 (N_2764,N_845,N_1627);
or U2765 (N_2765,N_913,N_1108);
or U2766 (N_2766,N_1953,N_1414);
nand U2767 (N_2767,N_1656,N_616);
and U2768 (N_2768,N_2455,N_1905);
or U2769 (N_2769,N_1990,N_2157);
nor U2770 (N_2770,N_1888,N_941);
or U2771 (N_2771,N_2464,N_804);
and U2772 (N_2772,N_173,N_646);
and U2773 (N_2773,N_936,N_1537);
nor U2774 (N_2774,N_2171,N_1492);
or U2775 (N_2775,N_456,N_1026);
nor U2776 (N_2776,N_23,N_1347);
or U2777 (N_2777,N_198,N_214);
nand U2778 (N_2778,N_2132,N_1771);
or U2779 (N_2779,N_1812,N_2033);
nand U2780 (N_2780,N_1459,N_2208);
nand U2781 (N_2781,N_681,N_1995);
and U2782 (N_2782,N_1512,N_1447);
nand U2783 (N_2783,N_604,N_150);
nor U2784 (N_2784,N_1185,N_907);
or U2785 (N_2785,N_2142,N_1943);
nor U2786 (N_2786,N_61,N_2467);
or U2787 (N_2787,N_1116,N_2319);
nor U2788 (N_2788,N_637,N_2396);
nor U2789 (N_2789,N_129,N_196);
nor U2790 (N_2790,N_1676,N_2138);
and U2791 (N_2791,N_1251,N_671);
and U2792 (N_2792,N_1113,N_1009);
nor U2793 (N_2793,N_1947,N_1446);
or U2794 (N_2794,N_2444,N_2190);
xnor U2795 (N_2795,N_1435,N_1819);
nand U2796 (N_2796,N_180,N_700);
and U2797 (N_2797,N_642,N_417);
nand U2798 (N_2798,N_334,N_2287);
and U2799 (N_2799,N_1254,N_2290);
nor U2800 (N_2800,N_425,N_649);
nand U2801 (N_2801,N_483,N_1144);
nand U2802 (N_2802,N_1075,N_938);
or U2803 (N_2803,N_909,N_1238);
nand U2804 (N_2804,N_2166,N_680);
nor U2805 (N_2805,N_2386,N_513);
nand U2806 (N_2806,N_2091,N_774);
nor U2807 (N_2807,N_837,N_1348);
or U2808 (N_2808,N_175,N_234);
and U2809 (N_2809,N_1283,N_2178);
and U2810 (N_2810,N_271,N_696);
nand U2811 (N_2811,N_299,N_1120);
or U2812 (N_2812,N_4,N_592);
or U2813 (N_2813,N_608,N_371);
xnor U2814 (N_2814,N_354,N_53);
nor U2815 (N_2815,N_1701,N_1127);
nor U2816 (N_2816,N_1301,N_2248);
nor U2817 (N_2817,N_1450,N_576);
or U2818 (N_2818,N_98,N_2003);
or U2819 (N_2819,N_2193,N_2493);
nand U2820 (N_2820,N_1932,N_661);
or U2821 (N_2821,N_131,N_1639);
nand U2822 (N_2822,N_102,N_1767);
or U2823 (N_2823,N_1675,N_2094);
and U2824 (N_2824,N_123,N_984);
and U2825 (N_2825,N_2212,N_863);
nand U2826 (N_2826,N_409,N_1846);
nand U2827 (N_2827,N_703,N_699);
nand U2828 (N_2828,N_432,N_589);
or U2829 (N_2829,N_2245,N_2251);
nand U2830 (N_2830,N_2452,N_34);
or U2831 (N_2831,N_1636,N_1024);
nand U2832 (N_2832,N_1302,N_1300);
and U2833 (N_2833,N_1487,N_1292);
nand U2834 (N_2834,N_1839,N_790);
nand U2835 (N_2835,N_1672,N_1339);
nand U2836 (N_2836,N_695,N_1797);
nand U2837 (N_2837,N_1021,N_1773);
and U2838 (N_2838,N_147,N_1356);
and U2839 (N_2839,N_810,N_1044);
nor U2840 (N_2840,N_958,N_122);
nor U2841 (N_2841,N_20,N_2497);
nand U2842 (N_2842,N_2061,N_2000);
or U2843 (N_2843,N_69,N_1653);
or U2844 (N_2844,N_1346,N_648);
or U2845 (N_2845,N_146,N_144);
or U2846 (N_2846,N_1577,N_532);
and U2847 (N_2847,N_772,N_2122);
xnor U2848 (N_2848,N_1867,N_256);
nor U2849 (N_2849,N_2355,N_178);
nand U2850 (N_2850,N_534,N_2384);
nor U2851 (N_2851,N_1337,N_355);
nand U2852 (N_2852,N_2411,N_2492);
nand U2853 (N_2853,N_1100,N_1221);
or U2854 (N_2854,N_1494,N_2036);
and U2855 (N_2855,N_133,N_18);
or U2856 (N_2856,N_383,N_184);
and U2857 (N_2857,N_306,N_2479);
nor U2858 (N_2858,N_93,N_663);
and U2859 (N_2859,N_0,N_1569);
and U2860 (N_2860,N_2478,N_2465);
and U2861 (N_2861,N_947,N_1253);
or U2862 (N_2862,N_1107,N_99);
nor U2863 (N_2863,N_1461,N_779);
nor U2864 (N_2864,N_1399,N_581);
nor U2865 (N_2865,N_313,N_718);
or U2866 (N_2866,N_578,N_585);
and U2867 (N_2867,N_361,N_1764);
and U2868 (N_2868,N_49,N_1126);
nor U2869 (N_2869,N_923,N_1209);
or U2870 (N_2870,N_1574,N_1694);
or U2871 (N_2871,N_1357,N_1965);
nand U2872 (N_2872,N_1141,N_2175);
nor U2873 (N_2873,N_1005,N_1563);
nand U2874 (N_2874,N_2257,N_630);
or U2875 (N_2875,N_2325,N_832);
nor U2876 (N_2876,N_84,N_2005);
or U2877 (N_2877,N_1851,N_635);
and U2878 (N_2878,N_1365,N_1658);
nand U2879 (N_2879,N_2323,N_2419);
or U2880 (N_2880,N_1735,N_1434);
or U2881 (N_2881,N_823,N_603);
nor U2882 (N_2882,N_767,N_182);
nand U2883 (N_2883,N_1247,N_2247);
and U2884 (N_2884,N_1884,N_1902);
and U2885 (N_2885,N_1272,N_633);
nor U2886 (N_2886,N_13,N_1881);
nor U2887 (N_2887,N_2065,N_1775);
or U2888 (N_2888,N_549,N_1857);
or U2889 (N_2889,N_1410,N_245);
or U2890 (N_2890,N_2049,N_1908);
and U2891 (N_2891,N_1073,N_413);
and U2892 (N_2892,N_582,N_1433);
and U2893 (N_2893,N_1874,N_1183);
or U2894 (N_2894,N_1944,N_517);
nand U2895 (N_2895,N_1796,N_1230);
or U2896 (N_2896,N_43,N_931);
nor U2897 (N_2897,N_112,N_1147);
or U2898 (N_2898,N_1821,N_1674);
nand U2899 (N_2899,N_1956,N_1466);
nor U2900 (N_2900,N_338,N_2357);
nand U2901 (N_2901,N_686,N_79);
nand U2902 (N_2902,N_398,N_1265);
and U2903 (N_2903,N_153,N_567);
or U2904 (N_2904,N_871,N_280);
nand U2905 (N_2905,N_732,N_441);
or U2906 (N_2906,N_423,N_791);
nor U2907 (N_2907,N_219,N_1043);
nand U2908 (N_2908,N_1246,N_889);
or U2909 (N_2909,N_2391,N_1047);
nand U2910 (N_2910,N_2490,N_202);
or U2911 (N_2911,N_1697,N_429);
nand U2912 (N_2912,N_2279,N_1159);
nand U2913 (N_2913,N_1279,N_83);
nand U2914 (N_2914,N_94,N_347);
nand U2915 (N_2915,N_2133,N_2180);
nor U2916 (N_2916,N_1449,N_446);
and U2917 (N_2917,N_2232,N_1741);
nor U2918 (N_2918,N_1380,N_2387);
and U2919 (N_2919,N_364,N_1829);
and U2920 (N_2920,N_2289,N_2250);
nor U2921 (N_2921,N_1751,N_1869);
and U2922 (N_2922,N_1476,N_1472);
xor U2923 (N_2923,N_544,N_1755);
nand U2924 (N_2924,N_613,N_741);
nor U2925 (N_2925,N_1271,N_1700);
or U2926 (N_2926,N_2026,N_1844);
nor U2927 (N_2927,N_1248,N_1863);
nor U2928 (N_2928,N_828,N_166);
nor U2929 (N_2929,N_1772,N_875);
nand U2930 (N_2930,N_1682,N_860);
nor U2931 (N_2931,N_2362,N_634);
nor U2932 (N_2932,N_67,N_211);
and U2933 (N_2933,N_1992,N_895);
nand U2934 (N_2934,N_1724,N_1920);
and U2935 (N_2935,N_58,N_1099);
xnor U2936 (N_2936,N_639,N_691);
nand U2937 (N_2937,N_1922,N_1659);
nor U2938 (N_2938,N_345,N_627);
or U2939 (N_2939,N_2101,N_2089);
or U2940 (N_2940,N_1580,N_1722);
nand U2941 (N_2941,N_2263,N_1196);
nor U2942 (N_2942,N_445,N_1208);
nor U2943 (N_2943,N_1910,N_1485);
nand U2944 (N_2944,N_798,N_533);
or U2945 (N_2945,N_368,N_1663);
nand U2946 (N_2946,N_2086,N_1454);
or U2947 (N_2947,N_1285,N_2436);
or U2948 (N_2948,N_382,N_318);
nand U2949 (N_2949,N_583,N_1211);
nand U2950 (N_2950,N_1139,N_2059);
nand U2951 (N_2951,N_861,N_208);
or U2952 (N_2952,N_128,N_880);
or U2953 (N_2953,N_809,N_512);
nand U2954 (N_2954,N_1808,N_933);
or U2955 (N_2955,N_1556,N_1323);
or U2956 (N_2956,N_1242,N_1936);
or U2957 (N_2957,N_2234,N_2283);
or U2958 (N_2958,N_1632,N_204);
nor U2959 (N_2959,N_2218,N_2470);
or U2960 (N_2960,N_1590,N_1618);
nand U2961 (N_2961,N_2335,N_1227);
nor U2962 (N_2962,N_1121,N_1942);
and U2963 (N_2963,N_1924,N_1083);
nor U2964 (N_2964,N_320,N_607);
or U2965 (N_2965,N_2428,N_1579);
nand U2966 (N_2966,N_2468,N_297);
and U2967 (N_2967,N_193,N_1295);
nor U2968 (N_2968,N_1318,N_357);
and U2969 (N_2969,N_2471,N_1749);
nand U2970 (N_2970,N_479,N_160);
nand U2971 (N_2971,N_54,N_1174);
or U2972 (N_2972,N_2210,N_1374);
and U2973 (N_2973,N_2299,N_1303);
nand U2974 (N_2974,N_1536,N_2226);
nand U2975 (N_2975,N_1564,N_744);
nand U2976 (N_2976,N_2407,N_2240);
nor U2977 (N_2977,N_319,N_1714);
nand U2978 (N_2978,N_2282,N_981);
and U2979 (N_2979,N_2141,N_1517);
or U2980 (N_2980,N_1010,N_2451);
nand U2981 (N_2981,N_1225,N_1409);
nor U2982 (N_2982,N_290,N_507);
nor U2983 (N_2983,N_185,N_283);
nor U2984 (N_2984,N_1506,N_1885);
nand U2985 (N_2985,N_1622,N_296);
nand U2986 (N_2986,N_237,N_30);
nor U2987 (N_2987,N_806,N_1952);
or U2988 (N_2988,N_294,N_1353);
nand U2989 (N_2989,N_1900,N_927);
or U2990 (N_2990,N_784,N_145);
nor U2991 (N_2991,N_2429,N_2198);
nor U2992 (N_2992,N_1873,N_65);
nor U2993 (N_2993,N_706,N_2149);
nor U2994 (N_2994,N_2181,N_1172);
and U2995 (N_2995,N_514,N_135);
nor U2996 (N_2996,N_2016,N_2229);
nor U2997 (N_2997,N_1235,N_731);
nand U2998 (N_2998,N_1534,N_217);
and U2999 (N_2999,N_235,N_932);
nor U3000 (N_3000,N_1491,N_2486);
nand U3001 (N_3001,N_1182,N_28);
nand U3002 (N_3002,N_316,N_467);
nor U3003 (N_3003,N_358,N_911);
nor U3004 (N_3004,N_495,N_1507);
nand U3005 (N_3005,N_762,N_2459);
and U3006 (N_3006,N_439,N_121);
xnor U3007 (N_3007,N_723,N_1451);
nor U3008 (N_3008,N_1645,N_1685);
and U3009 (N_3009,N_472,N_1175);
nand U3010 (N_3010,N_216,N_304);
nand U3011 (N_3011,N_1252,N_266);
nand U3012 (N_3012,N_262,N_1131);
or U3013 (N_3013,N_1188,N_2333);
and U3014 (N_3014,N_1854,N_2246);
nor U3015 (N_3015,N_1818,N_773);
nor U3016 (N_3016,N_82,N_1841);
nand U3017 (N_3017,N_1815,N_573);
nor U3018 (N_3018,N_737,N_1666);
and U3019 (N_3019,N_1897,N_310);
nand U3020 (N_3020,N_969,N_855);
or U3021 (N_3021,N_1760,N_142);
or U3022 (N_3022,N_342,N_381);
nor U3023 (N_3023,N_2228,N_1684);
and U3024 (N_3024,N_2110,N_500);
or U3025 (N_3025,N_1915,N_745);
and U3026 (N_3026,N_264,N_300);
nor U3027 (N_3027,N_1761,N_1289);
xnor U3028 (N_3028,N_2060,N_1480);
and U3029 (N_3029,N_2476,N_1661);
or U3030 (N_3030,N_418,N_1245);
or U3031 (N_3031,N_1678,N_1505);
or U3032 (N_3032,N_1199,N_716);
nor U3033 (N_3033,N_733,N_1599);
xnor U3034 (N_3034,N_1309,N_2400);
nor U3035 (N_3035,N_2155,N_103);
and U3036 (N_3036,N_586,N_1053);
nor U3037 (N_3037,N_1557,N_2432);
or U3038 (N_3038,N_2150,N_2019);
nand U3039 (N_3039,N_360,N_1048);
and U3040 (N_3040,N_1504,N_2462);
and U3041 (N_3041,N_469,N_1224);
nand U3042 (N_3042,N_735,N_2154);
nor U3043 (N_3043,N_2498,N_655);
or U3044 (N_3044,N_945,N_1373);
nand U3045 (N_3045,N_2403,N_1051);
and U3046 (N_3046,N_739,N_484);
or U3047 (N_3047,N_298,N_1551);
or U3048 (N_3048,N_2011,N_1477);
nand U3049 (N_3049,N_244,N_100);
nand U3050 (N_3050,N_2349,N_2365);
and U3051 (N_3051,N_503,N_1190);
nand U3052 (N_3052,N_1866,N_1419);
nor U3053 (N_3053,N_961,N_758);
or U3054 (N_3054,N_327,N_460);
nor U3055 (N_3055,N_1164,N_2423);
nor U3056 (N_3056,N_1671,N_2329);
or U3057 (N_3057,N_2017,N_1807);
or U3058 (N_3058,N_2205,N_720);
or U3059 (N_3059,N_2107,N_1096);
and U3060 (N_3060,N_1345,N_682);
or U3061 (N_3061,N_2230,N_1732);
nand U3062 (N_3062,N_2258,N_232);
or U3063 (N_3063,N_891,N_1008);
and U3064 (N_3064,N_2281,N_541);
nand U3065 (N_3065,N_1291,N_1432);
or U3066 (N_3066,N_1788,N_497);
nand U3067 (N_3067,N_1488,N_2259);
nand U3068 (N_3068,N_468,N_1898);
and U3069 (N_3069,N_1954,N_66);
nor U3070 (N_3070,N_897,N_1985);
nor U3071 (N_3071,N_400,N_1883);
nand U3072 (N_3072,N_2297,N_260);
or U3073 (N_3073,N_2371,N_157);
and U3074 (N_3074,N_210,N_1422);
and U3075 (N_3075,N_614,N_1290);
or U3076 (N_3076,N_203,N_1368);
nand U3077 (N_3077,N_369,N_1039);
or U3078 (N_3078,N_593,N_1896);
and U3079 (N_3079,N_1988,N_2012);
or U3080 (N_3080,N_29,N_238);
nand U3081 (N_3081,N_548,N_992);
nor U3082 (N_3082,N_1533,N_1930);
nor U3083 (N_3083,N_951,N_843);
or U3084 (N_3084,N_187,N_611);
nand U3085 (N_3085,N_579,N_942);
or U3086 (N_3086,N_2438,N_2426);
nand U3087 (N_3087,N_2183,N_397);
nor U3088 (N_3088,N_959,N_1475);
nor U3089 (N_3089,N_485,N_2158);
nor U3090 (N_3090,N_2047,N_1617);
or U3091 (N_3091,N_2394,N_1020);
or U3092 (N_3092,N_1389,N_96);
and U3093 (N_3093,N_374,N_2043);
nand U3094 (N_3094,N_267,N_1064);
nor U3095 (N_3095,N_998,N_708);
or U3096 (N_3096,N_459,N_1514);
and U3097 (N_3097,N_1594,N_1552);
nand U3098 (N_3098,N_2274,N_1532);
and U3099 (N_3099,N_736,N_935);
nand U3100 (N_3100,N_1354,N_1683);
or U3101 (N_3101,N_2322,N_165);
or U3102 (N_3102,N_2126,N_1893);
and U3103 (N_3103,N_978,N_726);
nand U3104 (N_3104,N_1971,N_2363);
and U3105 (N_3105,N_683,N_713);
or U3106 (N_3106,N_2372,N_1923);
and U3107 (N_3107,N_1782,N_796);
or U3108 (N_3108,N_1626,N_647);
nor U3109 (N_3109,N_1421,N_1833);
nor U3110 (N_3110,N_307,N_908);
nor U3111 (N_3111,N_410,N_1444);
and U3112 (N_3112,N_529,N_999);
or U3113 (N_3113,N_528,N_1934);
nor U3114 (N_3114,N_601,N_602);
and U3115 (N_3115,N_516,N_1473);
or U3116 (N_3116,N_876,N_2148);
and U3117 (N_3117,N_1195,N_768);
nor U3118 (N_3118,N_431,N_1882);
nor U3119 (N_3119,N_1019,N_1555);
or U3120 (N_3120,N_2020,N_824);
nor U3121 (N_3121,N_520,N_1134);
or U3122 (N_3122,N_470,N_1336);
or U3123 (N_3123,N_834,N_1515);
or U3124 (N_3124,N_742,N_1789);
nor U3125 (N_3125,N_1034,N_2121);
and U3126 (N_3126,N_2420,N_1834);
nand U3127 (N_3127,N_77,N_115);
nor U3128 (N_3128,N_303,N_1408);
nand U3129 (N_3129,N_1904,N_624);
xnor U3130 (N_3130,N_392,N_1716);
nand U3131 (N_3131,N_189,N_505);
and U3132 (N_3132,N_1862,N_1545);
nor U3133 (N_3133,N_1728,N_2334);
and U3134 (N_3134,N_826,N_1465);
or U3135 (N_3135,N_1091,N_664);
nor U3136 (N_3136,N_2176,N_335);
nand U3137 (N_3137,N_1591,N_465);
or U3138 (N_3138,N_1669,N_243);
and U3139 (N_3139,N_408,N_177);
or U3140 (N_3140,N_1550,N_688);
or U3141 (N_3141,N_1911,N_2);
nor U3142 (N_3142,N_2206,N_524);
nand U3143 (N_3143,N_1852,N_1957);
or U3144 (N_3144,N_1624,N_181);
or U3145 (N_3145,N_47,N_426);
nor U3146 (N_3146,N_1249,N_1817);
nor U3147 (N_3147,N_1146,N_1032);
or U3148 (N_3148,N_1482,N_2081);
and U3149 (N_3149,N_1273,N_565);
nor U3150 (N_3150,N_2048,N_1430);
or U3151 (N_3151,N_2055,N_90);
nand U3152 (N_3152,N_783,N_230);
nand U3153 (N_3153,N_255,N_2494);
or U3154 (N_3154,N_363,N_1321);
or U3155 (N_3155,N_949,N_523);
or U3156 (N_3156,N_1847,N_904);
and U3157 (N_3157,N_2080,N_818);
or U3158 (N_3158,N_677,N_2160);
or U3159 (N_3159,N_2318,N_1217);
nand U3160 (N_3160,N_1587,N_591);
nor U3161 (N_3161,N_1402,N_2268);
xnor U3162 (N_3162,N_1895,N_1396);
nand U3163 (N_3163,N_957,N_2260);
or U3164 (N_3164,N_1056,N_57);
or U3165 (N_3165,N_1776,N_1631);
or U3166 (N_3166,N_894,N_2172);
nor U3167 (N_3167,N_1837,N_1156);
nor U3168 (N_3168,N_2457,N_906);
and U3169 (N_3169,N_2131,N_1742);
and U3170 (N_3170,N_1986,N_454);
or U3171 (N_3171,N_1085,N_2021);
xnor U3172 (N_3172,N_599,N_2254);
nand U3173 (N_3173,N_88,N_2029);
and U3174 (N_3174,N_1180,N_1293);
and U3175 (N_3175,N_1133,N_2382);
nand U3176 (N_3176,N_254,N_404);
or U3177 (N_3177,N_662,N_1468);
or U3178 (N_3178,N_2317,N_2071);
or U3179 (N_3179,N_2023,N_1431);
or U3180 (N_3180,N_2249,N_433);
and U3181 (N_3181,N_233,N_2356);
nor U3182 (N_3182,N_888,N_525);
or U3183 (N_3183,N_898,N_665);
and U3184 (N_3184,N_727,N_1937);
or U3185 (N_3185,N_2007,N_1042);
nand U3186 (N_3186,N_170,N_421);
and U3187 (N_3187,N_1360,N_1049);
and U3188 (N_3188,N_325,N_2324);
and U3189 (N_3189,N_19,N_976);
and U3190 (N_3190,N_1929,N_1668);
nor U3191 (N_3191,N_1878,N_881);
or U3192 (N_3192,N_1935,N_1945);
nand U3193 (N_3193,N_1234,N_2066);
or U3194 (N_3194,N_1750,N_515);
nand U3195 (N_3195,N_1453,N_687);
nand U3196 (N_3196,N_728,N_990);
or U3197 (N_3197,N_1799,N_2222);
nand U3198 (N_3198,N_1723,N_2186);
or U3199 (N_3199,N_2439,N_2402);
nand U3200 (N_3200,N_1388,N_997);
and U3201 (N_3201,N_62,N_2408);
or U3202 (N_3202,N_983,N_2368);
and U3203 (N_3203,N_802,N_884);
nor U3204 (N_3204,N_494,N_848);
nand U3205 (N_3205,N_2087,N_842);
nand U3206 (N_3206,N_678,N_2264);
nand U3207 (N_3207,N_1027,N_1256);
nand U3208 (N_3208,N_2373,N_1200);
and U3209 (N_3209,N_263,N_167);
and U3210 (N_3210,N_265,N_2125);
nor U3211 (N_3211,N_1058,N_1093);
and U3212 (N_3212,N_466,N_1340);
nor U3213 (N_3213,N_2244,N_977);
and U3214 (N_3214,N_1664,N_1016);
nand U3215 (N_3215,N_2293,N_775);
nand U3216 (N_3216,N_1330,N_1733);
and U3217 (N_3217,N_2030,N_807);
or U3218 (N_3218,N_1014,N_1377);
nand U3219 (N_3219,N_1652,N_86);
and U3220 (N_3220,N_1715,N_1015);
and U3221 (N_3221,N_2269,N_305);
and U3222 (N_3222,N_2393,N_163);
nor U3223 (N_3223,N_471,N_236);
or U3224 (N_3224,N_1738,N_1978);
and U3225 (N_3225,N_2395,N_1206);
or U3226 (N_3226,N_2143,N_1470);
and U3227 (N_3227,N_542,N_1495);
nor U3228 (N_3228,N_1106,N_1647);
nand U3229 (N_3229,N_1062,N_1592);
or U3230 (N_3230,N_555,N_154);
and U3231 (N_3231,N_463,N_1702);
nor U3232 (N_3232,N_1921,N_882);
nand U3233 (N_3233,N_1887,N_1801);
and U3234 (N_3234,N_2364,N_858);
nand U3235 (N_3235,N_1437,N_1739);
or U3236 (N_3236,N_1160,N_2296);
or U3237 (N_3237,N_1711,N_1215);
nand U3238 (N_3238,N_489,N_2484);
nor U3239 (N_3239,N_148,N_218);
nand U3240 (N_3240,N_490,N_1692);
nor U3241 (N_3241,N_2388,N_2010);
nand U3242 (N_3242,N_476,N_1305);
nand U3243 (N_3243,N_427,N_948);
and U3244 (N_3244,N_393,N_632);
nor U3245 (N_3245,N_1145,N_124);
nand U3246 (N_3246,N_449,N_757);
and U3247 (N_3247,N_536,N_1226);
nand U3248 (N_3248,N_1778,N_1097);
or U3249 (N_3249,N_2092,N_1281);
and U3250 (N_3250,N_1541,N_2182);
nand U3251 (N_3251,N_618,N_190);
nand U3252 (N_3252,N_1549,N_1858);
nand U3253 (N_3253,N_689,N_1294);
or U3254 (N_3254,N_2196,N_1498);
nand U3255 (N_3255,N_405,N_2130);
or U3256 (N_3256,N_2461,N_651);
or U3257 (N_3257,N_797,N_753);
nor U3258 (N_3258,N_2078,N_654);
nand U3259 (N_3259,N_2344,N_340);
or U3260 (N_3260,N_137,N_281);
nor U3261 (N_3261,N_1439,N_1452);
xnor U3262 (N_3262,N_292,N_1072);
and U3263 (N_3263,N_183,N_1076);
nor U3264 (N_3264,N_2278,N_623);
or U3265 (N_3265,N_1614,N_2027);
nor U3266 (N_3266,N_291,N_1998);
and U3267 (N_3267,N_2147,N_1479);
xnor U3268 (N_3268,N_75,N_92);
or U3269 (N_3269,N_1050,N_444);
nor U3270 (N_3270,N_2079,N_1497);
or U3271 (N_3271,N_1162,N_2448);
or U3272 (N_3272,N_1785,N_1060);
nand U3273 (N_3273,N_21,N_1793);
or U3274 (N_3274,N_712,N_841);
nor U3275 (N_3275,N_152,N_1832);
or U3276 (N_3276,N_715,N_352);
nor U3277 (N_3277,N_1457,N_1232);
and U3278 (N_3278,N_2108,N_1351);
nand U3279 (N_3279,N_801,N_1680);
or U3280 (N_3280,N_660,N_1705);
nor U3281 (N_3281,N_329,N_453);
nand U3282 (N_3282,N_605,N_631);
and U3283 (N_3283,N_1280,N_1335);
and U3284 (N_3284,N_1142,N_769);
nand U3285 (N_3285,N_778,N_7);
nor U3286 (N_3286,N_1948,N_458);
and U3287 (N_3287,N_2487,N_1725);
nor U3288 (N_3288,N_868,N_1999);
nand U3289 (N_3289,N_2453,N_1036);
or U3290 (N_3290,N_995,N_1927);
and U3291 (N_3291,N_1464,N_353);
nor U3292 (N_3292,N_1513,N_1598);
or U3293 (N_3293,N_1605,N_546);
and U3294 (N_3294,N_1489,N_491);
xnor U3295 (N_3295,N_2309,N_498);
or U3296 (N_3296,N_14,N_1836);
and U3297 (N_3297,N_172,N_2339);
nor U3298 (N_3298,N_980,N_2201);
and U3299 (N_3299,N_1386,N_2119);
nand U3300 (N_3300,N_1752,N_521);
and U3301 (N_3301,N_1804,N_1445);
or U3302 (N_3302,N_963,N_2491);
nor U3303 (N_3303,N_2267,N_274);
and U3304 (N_3304,N_1926,N_559);
nor U3305 (N_3305,N_2024,N_42);
or U3306 (N_3306,N_996,N_317);
nand U3307 (N_3307,N_2437,N_1059);
nor U3308 (N_3308,N_1967,N_1805);
or U3309 (N_3309,N_725,N_1002);
nand U3310 (N_3310,N_846,N_1111);
or U3311 (N_3311,N_1730,N_419);
and U3312 (N_3312,N_117,N_32);
nor U3313 (N_3313,N_1067,N_2332);
nor U3314 (N_3314,N_1802,N_272);
and U3315 (N_3315,N_873,N_562);
nand U3316 (N_3316,N_1503,N_1559);
nand U3317 (N_3317,N_451,N_1928);
and U3318 (N_3318,N_2202,N_199);
nor U3319 (N_3319,N_2327,N_1628);
nand U3320 (N_3320,N_1267,N_1554);
and U3321 (N_3321,N_2449,N_1548);
nand U3322 (N_3322,N_1791,N_87);
nand U3323 (N_3323,N_1650,N_1167);
and U3324 (N_3324,N_2271,N_1262);
and U3325 (N_3325,N_1078,N_63);
or U3326 (N_3326,N_2331,N_1997);
nand U3327 (N_3327,N_1359,N_1427);
or U3328 (N_3328,N_2134,N_827);
nand U3329 (N_3329,N_2105,N_853);
or U3330 (N_3330,N_1086,N_416);
or U3331 (N_3331,N_870,N_2414);
and U3332 (N_3332,N_389,N_162);
nand U3333 (N_3333,N_1307,N_1651);
or U3334 (N_3334,N_1187,N_1766);
nand U3335 (N_3335,N_1991,N_547);
nand U3336 (N_3336,N_612,N_1375);
nand U3337 (N_3337,N_2315,N_246);
nor U3338 (N_3338,N_1210,N_1125);
nand U3339 (N_3339,N_685,N_1163);
nor U3340 (N_3340,N_1098,N_213);
or U3341 (N_3341,N_1092,N_2195);
nand U3342 (N_3342,N_1105,N_2187);
nor U3343 (N_3343,N_1783,N_1329);
nor U3344 (N_3344,N_1868,N_1219);
nand U3345 (N_3345,N_2284,N_1762);
nand U3346 (N_3346,N_2485,N_1864);
or U3347 (N_3347,N_2135,N_921);
nor U3348 (N_3348,N_2235,N_349);
and U3349 (N_3349,N_674,N_2237);
nor U3350 (N_3350,N_1931,N_76);
and U3351 (N_3351,N_1763,N_854);
nand U3352 (N_3352,N_1316,N_1471);
nor U3353 (N_3353,N_2004,N_535);
and U3354 (N_3354,N_835,N_2044);
nor U3355 (N_3355,N_885,N_1786);
or U3356 (N_3356,N_955,N_1604);
nand U3357 (N_3357,N_1568,N_557);
and U3358 (N_3358,N_943,N_1181);
or U3359 (N_3359,N_1914,N_16);
or U3360 (N_3360,N_851,N_1850);
and U3361 (N_3361,N_1395,N_1781);
and U3362 (N_3362,N_452,N_1601);
or U3363 (N_3363,N_729,N_143);
nand U3364 (N_3364,N_1729,N_1397);
and U3365 (N_3365,N_1173,N_2275);
nor U3366 (N_3366,N_341,N_259);
and U3367 (N_3367,N_1746,N_777);
nand U3368 (N_3368,N_496,N_740);
or U3369 (N_3369,N_1284,N_2401);
or U3370 (N_3370,N_2266,N_1298);
or U3371 (N_3371,N_917,N_403);
xnor U3372 (N_3372,N_1481,N_1609);
nand U3373 (N_3373,N_2469,N_1826);
or U3374 (N_3374,N_805,N_538);
and U3375 (N_3375,N_2286,N_2495);
nor U3376 (N_3376,N_1644,N_1077);
nor U3377 (N_3377,N_478,N_2221);
nor U3378 (N_3378,N_2321,N_64);
or U3379 (N_3379,N_714,N_110);
or U3380 (N_3380,N_1906,N_2140);
nand U3381 (N_3381,N_367,N_830);
nor U3382 (N_3382,N_622,N_518);
nor U3383 (N_3383,N_286,N_396);
nor U3384 (N_3384,N_1519,N_2370);
and U3385 (N_3385,N_1820,N_816);
or U3386 (N_3386,N_2168,N_2425);
nand U3387 (N_3387,N_377,N_2392);
nand U3388 (N_3388,N_900,N_1366);
and U3389 (N_3389,N_1596,N_1860);
or U3390 (N_3390,N_2001,N_1222);
or U3391 (N_3391,N_1754,N_721);
nand U3392 (N_3392,N_569,N_1673);
nand U3393 (N_3393,N_887,N_1629);
and U3394 (N_3394,N_1104,N_1795);
nor U3395 (N_3395,N_1220,N_73);
and U3396 (N_3396,N_1961,N_1462);
or U3397 (N_3397,N_1765,N_925);
and U3398 (N_3398,N_2328,N_1657);
and U3399 (N_3399,N_151,N_1119);
or U3400 (N_3400,N_179,N_119);
or U3401 (N_3401,N_2358,N_328);
nand U3402 (N_3402,N_1777,N_552);
nand U3403 (N_3403,N_795,N_508);
nor U3404 (N_3404,N_384,N_1274);
nand U3405 (N_3405,N_1115,N_1244);
and U3406 (N_3406,N_962,N_1737);
or U3407 (N_3407,N_270,N_1538);
or U3408 (N_3408,N_2280,N_45);
or U3409 (N_3409,N_350,N_22);
and U3410 (N_3410,N_1721,N_2440);
nor U3411 (N_3411,N_24,N_109);
nand U3412 (N_3412,N_1520,N_1500);
nor U3413 (N_3413,N_1266,N_1089);
nor U3414 (N_3414,N_1606,N_1233);
nand U3415 (N_3415,N_1417,N_2360);
nand U3416 (N_3416,N_1709,N_1973);
and U3417 (N_3417,N_2093,N_615);
nand U3418 (N_3418,N_2256,N_1204);
nand U3419 (N_3419,N_2170,N_59);
nand U3420 (N_3420,N_1753,N_373);
nand U3421 (N_3421,N_2069,N_679);
nor U3422 (N_3422,N_820,N_944);
nand U3423 (N_3423,N_1814,N_694);
or U3424 (N_3424,N_2114,N_1980);
nor U3425 (N_3425,N_510,N_2262);
and U3426 (N_3426,N_1012,N_1052);
nor U3427 (N_3427,N_226,N_1094);
and U3428 (N_3428,N_676,N_1239);
nor U3429 (N_3429,N_1352,N_1843);
nor U3430 (N_3430,N_597,N_2238);
and U3431 (N_3431,N_765,N_1469);
xor U3432 (N_3432,N_41,N_1194);
nand U3433 (N_3433,N_1613,N_2380);
nor U3434 (N_3434,N_1969,N_966);
or U3435 (N_3435,N_1803,N_1543);
nand U3436 (N_3436,N_1261,N_434);
nor U3437 (N_3437,N_372,N_1891);
or U3438 (N_3438,N_437,N_1708);
or U3439 (N_3439,N_1000,N_2199);
or U3440 (N_3440,N_1736,N_2137);
and U3441 (N_3441,N_1727,N_1212);
or U3442 (N_3442,N_2443,N_847);
nand U3443 (N_3443,N_1508,N_108);
nor U3444 (N_3444,N_2374,N_610);
or U3445 (N_3445,N_72,N_139);
and U3446 (N_3446,N_1288,N_428);
or U3447 (N_3447,N_12,N_2102);
or U3448 (N_3448,N_1455,N_2456);
nor U3449 (N_3449,N_2162,N_2090);
nand U3450 (N_3450,N_1326,N_401);
nand U3451 (N_3451,N_125,N_209);
nor U3452 (N_3452,N_551,N_836);
or U3453 (N_3453,N_1486,N_1546);
nand U3454 (N_3454,N_684,N_40);
nand U3455 (N_3455,N_2083,N_339);
or U3456 (N_3456,N_1933,N_2073);
nand U3457 (N_3457,N_46,N_930);
and U3458 (N_3458,N_566,N_749);
or U3459 (N_3459,N_6,N_1571);
or U3460 (N_3460,N_2224,N_1522);
or U3461 (N_3461,N_362,N_1429);
xnor U3462 (N_3462,N_1405,N_833);
or U3463 (N_3463,N_993,N_2480);
nor U3464 (N_3464,N_1213,N_1955);
nor U3465 (N_3465,N_1892,N_1007);
or U3466 (N_3466,N_44,N_1168);
xor U3467 (N_3467,N_939,N_2097);
and U3468 (N_3468,N_1319,N_2233);
nand U3469 (N_3469,N_670,N_1358);
or U3470 (N_3470,N_111,N_1901);
and U3471 (N_3471,N_1949,N_1703);
and U3472 (N_3472,N_406,N_879);
nand U3473 (N_3473,N_1484,N_1192);
or U3474 (N_3474,N_302,N_869);
and U3475 (N_3475,N_2214,N_756);
or U3476 (N_3476,N_1690,N_1103);
and U3477 (N_3477,N_2310,N_365);
xor U3478 (N_3478,N_673,N_575);
and U3479 (N_3479,N_1540,N_526);
nor U3480 (N_3480,N_872,N_435);
or U3481 (N_3481,N_35,N_1379);
nand U3482 (N_3482,N_2192,N_1057);
nor U3483 (N_3483,N_301,N_1667);
nor U3484 (N_3484,N_114,N_1214);
and U3485 (N_3485,N_390,N_2377);
or U3486 (N_3486,N_2115,N_1918);
nor U3487 (N_3487,N_2375,N_764);
and U3488 (N_3488,N_156,N_1525);
nand U3489 (N_3489,N_1779,N_457);
nor U3490 (N_3490,N_2338,N_2050);
or U3491 (N_3491,N_1334,N_1774);
nor U3492 (N_3492,N_1258,N_1925);
nor U3493 (N_3493,N_1570,N_1231);
or U3494 (N_3494,N_1197,N_1361);
nand U3495 (N_3495,N_2031,N_2265);
xor U3496 (N_3496,N_692,N_2242);
nor U3497 (N_3497,N_1394,N_1478);
or U3498 (N_3498,N_1263,N_1938);
nand U3499 (N_3499,N_2474,N_2295);
nor U3500 (N_3500,N_1013,N_2359);
and U3501 (N_3501,N_1257,N_1400);
and U3502 (N_3502,N_840,N_1033);
nand U3503 (N_3503,N_1148,N_1996);
nor U3504 (N_3504,N_1588,N_1313);
nor U3505 (N_3505,N_2144,N_212);
nor U3506 (N_3506,N_1706,N_838);
or U3507 (N_3507,N_653,N_672);
or U3508 (N_3508,N_1641,N_1054);
and U3509 (N_3509,N_1349,N_481);
and U3510 (N_3510,N_2460,N_60);
and U3511 (N_3511,N_1919,N_2354);
and U3512 (N_3512,N_1376,N_1179);
or U3513 (N_3513,N_1816,N_323);
or U3514 (N_3514,N_1236,N_1081);
or U3515 (N_3515,N_883,N_442);
or U3516 (N_3516,N_1420,N_971);
and U3517 (N_3517,N_1619,N_2385);
nand U3518 (N_3518,N_2037,N_2421);
or U3519 (N_3519,N_1404,N_2191);
or U3520 (N_3520,N_803,N_2431);
or U3521 (N_3521,N_2445,N_1114);
or U3522 (N_3522,N_1011,N_312);
or U3523 (N_3523,N_2378,N_248);
nor U3524 (N_3524,N_488,N_2219);
or U3525 (N_3525,N_2076,N_985);
or U3526 (N_3526,N_1798,N_1363);
nor U3527 (N_3527,N_1516,N_2450);
or U3528 (N_3528,N_2481,N_920);
and U3529 (N_3529,N_169,N_223);
and U3530 (N_3530,N_388,N_822);
nor U3531 (N_3531,N_1768,N_315);
nand U3532 (N_3532,N_1524,N_2211);
or U3533 (N_3533,N_1178,N_2038);
nand U3534 (N_3534,N_207,N_1734);
and U3535 (N_3535,N_588,N_1218);
nor U3536 (N_3536,N_2189,N_1974);
nand U3537 (N_3537,N_799,N_2041);
nand U3538 (N_3538,N_1046,N_1074);
or U3539 (N_3539,N_1687,N_200);
and U3540 (N_3540,N_781,N_1166);
nor U3541 (N_3541,N_1712,N_811);
nor U3542 (N_3542,N_1123,N_568);
nand U3543 (N_3543,N_1413,N_1502);
or U3544 (N_3544,N_1719,N_1170);
xor U3545 (N_3545,N_385,N_1332);
nand U3546 (N_3546,N_937,N_1813);
nor U3547 (N_3547,N_2057,N_1743);
and U3548 (N_3548,N_1872,N_1704);
nand U3549 (N_3549,N_2117,N_1845);
or U3550 (N_3550,N_859,N_2348);
and U3551 (N_3551,N_1865,N_1940);
and U3552 (N_3552,N_2463,N_1848);
and U3553 (N_3553,N_2347,N_2088);
nor U3554 (N_3554,N_257,N_1790);
and U3555 (N_3555,N_1510,N_1322);
nand U3556 (N_3556,N_39,N_1582);
or U3557 (N_3557,N_391,N_1063);
or U3558 (N_3558,N_1981,N_1824);
xor U3559 (N_3559,N_132,N_1565);
and U3560 (N_3560,N_1369,N_590);
xor U3561 (N_3561,N_1151,N_2099);
nor U3562 (N_3562,N_1575,N_1643);
or U3563 (N_3563,N_1355,N_1364);
and U3564 (N_3564,N_890,N_1324);
or U3565 (N_3565,N_760,N_1136);
nor U3566 (N_3566,N_1635,N_1387);
xor U3567 (N_3567,N_594,N_289);
nor U3568 (N_3568,N_2215,N_878);
and U3569 (N_3569,N_159,N_2236);
nor U3570 (N_3570,N_440,N_285);
or U3571 (N_3571,N_2424,N_625);
nand U3572 (N_3572,N_750,N_1342);
or U3573 (N_3573,N_1203,N_1382);
nor U3574 (N_3574,N_1966,N_1391);
nor U3575 (N_3575,N_1260,N_852);
or U3576 (N_3576,N_370,N_1825);
or U3577 (N_3577,N_759,N_1521);
nand U3578 (N_3578,N_1946,N_952);
nand U3579 (N_3579,N_101,N_2252);
nor U3580 (N_3580,N_1381,N_2096);
or U3581 (N_3581,N_864,N_2304);
or U3582 (N_3582,N_1448,N_1069);
xor U3583 (N_3583,N_2153,N_1344);
nand U3584 (N_3584,N_638,N_2405);
nand U3585 (N_3585,N_224,N_1398);
and U3586 (N_3586,N_249,N_1003);
and U3587 (N_3587,N_1328,N_2447);
and U3588 (N_3588,N_1689,N_2008);
or U3589 (N_3589,N_247,N_1122);
or U3590 (N_3590,N_1240,N_2326);
xor U3591 (N_3591,N_839,N_563);
nor U3592 (N_3592,N_25,N_1458);
nor U3593 (N_3593,N_1941,N_91);
and U3594 (N_3594,N_2161,N_1383);
or U3595 (N_3595,N_1539,N_1558);
nand U3596 (N_3596,N_789,N_2223);
and U3597 (N_3597,N_31,N_1983);
nand U3598 (N_3598,N_527,N_1695);
nand U3599 (N_3599,N_448,N_1038);
nand U3600 (N_3600,N_570,N_268);
nand U3601 (N_3601,N_331,N_2035);
or U3602 (N_3602,N_2120,N_402);
nand U3603 (N_3603,N_1621,N_1633);
or U3604 (N_3604,N_1333,N_414);
or U3605 (N_3605,N_2472,N_915);
and U3606 (N_3606,N_2255,N_1372);
xor U3607 (N_3607,N_2416,N_1745);
or U3608 (N_3608,N_387,N_168);
and U3609 (N_3609,N_1916,N_2100);
nand U3610 (N_3610,N_928,N_574);
nor U3611 (N_3611,N_261,N_120);
nor U3612 (N_3612,N_2002,N_1853);
nor U3613 (N_3613,N_2084,N_321);
or U3614 (N_3614,N_1880,N_1384);
or U3615 (N_3615,N_2056,N_2136);
nor U3616 (N_3616,N_1070,N_407);
xnor U3617 (N_3617,N_967,N_378);
nor U3618 (N_3618,N_734,N_1296);
or U3619 (N_3619,N_924,N_698);
and U3620 (N_3620,N_1028,N_502);
nor U3621 (N_3621,N_1875,N_825);
and U3622 (N_3622,N_1411,N_991);
nor U3623 (N_3623,N_717,N_1493);
and U3624 (N_3624,N_2361,N_253);
nand U3625 (N_3625,N_276,N_1529);
nand U3626 (N_3626,N_960,N_351);
and U3627 (N_3627,N_511,N_1483);
nor U3628 (N_3628,N_874,N_2308);
or U3629 (N_3629,N_17,N_658);
or U3630 (N_3630,N_2046,N_191);
and U3631 (N_3631,N_929,N_1975);
nor U3632 (N_3632,N_1823,N_794);
or U3633 (N_3633,N_1137,N_97);
and U3634 (N_3634,N_2243,N_275);
and U3635 (N_3635,N_621,N_1646);
or U3636 (N_3636,N_553,N_693);
or U3637 (N_3637,N_443,N_2169);
and U3638 (N_3638,N_2410,N_11);
nand U3639 (N_3639,N_690,N_1370);
and U3640 (N_3640,N_1004,N_293);
and U3641 (N_3641,N_195,N_2173);
or U3642 (N_3642,N_113,N_1169);
and U3643 (N_3643,N_438,N_1811);
nand U3644 (N_3644,N_979,N_2052);
or U3645 (N_3645,N_2139,N_258);
nor U3646 (N_3646,N_229,N_269);
nor U3647 (N_3647,N_2499,N_954);
or U3648 (N_3648,N_1031,N_1315);
nor U3649 (N_3649,N_1976,N_530);
nand U3650 (N_3650,N_1806,N_311);
nand U3651 (N_3651,N_48,N_1325);
nand U3652 (N_3652,N_620,N_1117);
nor U3653 (N_3653,N_1870,N_376);
nand U3654 (N_3654,N_986,N_571);
and U3655 (N_3655,N_916,N_1718);
or U3656 (N_3656,N_2075,N_982);
nand U3657 (N_3657,N_787,N_2163);
nor U3658 (N_3658,N_1474,N_829);
or U3659 (N_3659,N_1630,N_2028);
nor U3660 (N_3660,N_2366,N_522);
nor U3661 (N_3661,N_2177,N_1831);
nand U3662 (N_3662,N_2014,N_2111);
nor U3663 (N_3663,N_1677,N_2165);
and U3664 (N_3664,N_1278,N_192);
nor U3665 (N_3665,N_394,N_1526);
or U3666 (N_3666,N_450,N_186);
nand U3667 (N_3667,N_2397,N_1528);
and U3668 (N_3668,N_2220,N_1842);
nand U3669 (N_3669,N_2489,N_1849);
nand U3670 (N_3670,N_2442,N_1314);
nand U3671 (N_3671,N_2127,N_1426);
nand U3672 (N_3672,N_2477,N_2473);
xor U3673 (N_3673,N_595,N_766);
nor U3674 (N_3674,N_2034,N_1531);
nor U3675 (N_3675,N_697,N_314);
nand U3676 (N_3676,N_519,N_628);
nor U3677 (N_3677,N_2343,N_1608);
or U3678 (N_3678,N_1713,N_149);
or U3679 (N_3679,N_1642,N_940);
nand U3680 (N_3680,N_1518,N_2409);
nor U3681 (N_3681,N_1890,N_1585);
and U3682 (N_3682,N_761,N_788);
nand U3683 (N_3683,N_1155,N_866);
nor U3684 (N_3684,N_702,N_1792);
nor U3685 (N_3685,N_136,N_477);
or U3686 (N_3686,N_792,N_580);
and U3687 (N_3687,N_1623,N_504);
or U3688 (N_3688,N_1443,N_2113);
and U3689 (N_3689,N_337,N_447);
or U3690 (N_3690,N_867,N_701);
or U3691 (N_3691,N_107,N_2330);
or U3692 (N_3692,N_415,N_332);
and U3693 (N_3693,N_953,N_2422);
nor U3694 (N_3694,N_666,N_273);
and U3695 (N_3695,N_709,N_324);
and U3696 (N_3696,N_2346,N_1320);
and U3697 (N_3697,N_239,N_197);
nand U3698 (N_3698,N_1780,N_1463);
and U3699 (N_3699,N_914,N_1686);
or U3700 (N_3700,N_786,N_1616);
nand U3701 (N_3701,N_2399,N_922);
or U3702 (N_3702,N_1509,N_657);
or U3703 (N_3703,N_493,N_1401);
nand U3704 (N_3704,N_2336,N_1423);
and U3705 (N_3705,N_2458,N_856);
nor U3706 (N_3706,N_748,N_2413);
nor U3707 (N_3707,N_1670,N_501);
and U3708 (N_3708,N_1425,N_2072);
nor U3709 (N_3709,N_1255,N_1082);
or U3710 (N_3710,N_1560,N_2018);
or U3711 (N_3711,N_965,N_1607);
and U3712 (N_3712,N_1061,N_51);
and U3713 (N_3713,N_1438,N_140);
or U3714 (N_3714,N_2441,N_705);
nand U3715 (N_3715,N_1228,N_50);
and U3716 (N_3716,N_905,N_1259);
nor U3717 (N_3717,N_1859,N_537);
and U3718 (N_3718,N_1989,N_346);
or U3719 (N_3719,N_1143,N_1310);
nor U3720 (N_3720,N_1586,N_1562);
nand U3721 (N_3721,N_1593,N_1152);
and U3722 (N_3722,N_1110,N_1951);
or U3723 (N_3723,N_1161,N_2039);
nand U3724 (N_3724,N_473,N_1029);
nor U3725 (N_3725,N_2435,N_2434);
or U3726 (N_3726,N_747,N_2276);
nand U3727 (N_3727,N_379,N_1572);
or U3728 (N_3728,N_509,N_430);
nor U3729 (N_3729,N_2351,N_1655);
and U3730 (N_3730,N_1698,N_1553);
or U3731 (N_3731,N_1406,N_336);
and U3732 (N_3732,N_710,N_1124);
nand U3733 (N_3733,N_1132,N_2151);
and U3734 (N_3734,N_252,N_1269);
or U3735 (N_3735,N_857,N_1250);
and U3736 (N_3736,N_1343,N_2483);
nand U3737 (N_3737,N_227,N_1095);
and U3738 (N_3738,N_26,N_896);
nor U3739 (N_3739,N_724,N_543);
or U3740 (N_3740,N_1306,N_1264);
nand U3741 (N_3741,N_2042,N_645);
or U3742 (N_3742,N_2231,N_348);
nor U3743 (N_3743,N_785,N_1331);
or U3744 (N_3744,N_1385,N_1090);
or U3745 (N_3745,N_1467,N_2184);
xor U3746 (N_3746,N_1573,N_1216);
and U3747 (N_3747,N_2152,N_912);
nand U3748 (N_3748,N_770,N_1071);
or U3749 (N_3749,N_2129,N_2054);
nor U3750 (N_3750,N_718,N_600);
nor U3751 (N_3751,N_424,N_323);
nor U3752 (N_3752,N_129,N_707);
nor U3753 (N_3753,N_2276,N_2216);
nor U3754 (N_3754,N_735,N_418);
nand U3755 (N_3755,N_923,N_358);
or U3756 (N_3756,N_2395,N_1790);
nand U3757 (N_3757,N_422,N_1760);
nor U3758 (N_3758,N_1129,N_2166);
and U3759 (N_3759,N_959,N_686);
and U3760 (N_3760,N_664,N_485);
nor U3761 (N_3761,N_50,N_1601);
and U3762 (N_3762,N_540,N_2448);
or U3763 (N_3763,N_933,N_2243);
or U3764 (N_3764,N_2124,N_2349);
and U3765 (N_3765,N_1664,N_1428);
nor U3766 (N_3766,N_1678,N_2289);
and U3767 (N_3767,N_1351,N_2275);
nand U3768 (N_3768,N_2354,N_1728);
nor U3769 (N_3769,N_1379,N_1478);
and U3770 (N_3770,N_1807,N_595);
and U3771 (N_3771,N_1277,N_19);
xnor U3772 (N_3772,N_601,N_334);
and U3773 (N_3773,N_1831,N_946);
and U3774 (N_3774,N_909,N_2385);
or U3775 (N_3775,N_1608,N_423);
nand U3776 (N_3776,N_1284,N_2219);
nand U3777 (N_3777,N_582,N_1205);
nand U3778 (N_3778,N_1399,N_814);
or U3779 (N_3779,N_1784,N_2488);
nand U3780 (N_3780,N_973,N_2406);
nor U3781 (N_3781,N_1171,N_847);
and U3782 (N_3782,N_828,N_265);
or U3783 (N_3783,N_793,N_1401);
or U3784 (N_3784,N_1897,N_28);
and U3785 (N_3785,N_1648,N_267);
or U3786 (N_3786,N_1790,N_1167);
nor U3787 (N_3787,N_1889,N_904);
or U3788 (N_3788,N_333,N_2317);
xnor U3789 (N_3789,N_1074,N_98);
or U3790 (N_3790,N_430,N_566);
or U3791 (N_3791,N_1341,N_1193);
nor U3792 (N_3792,N_322,N_1632);
nor U3793 (N_3793,N_1794,N_2491);
and U3794 (N_3794,N_1830,N_1349);
or U3795 (N_3795,N_679,N_1709);
nand U3796 (N_3796,N_97,N_1471);
or U3797 (N_3797,N_2220,N_2412);
nand U3798 (N_3798,N_663,N_161);
and U3799 (N_3799,N_1107,N_409);
or U3800 (N_3800,N_150,N_122);
nand U3801 (N_3801,N_100,N_420);
nor U3802 (N_3802,N_557,N_2065);
nand U3803 (N_3803,N_839,N_1279);
nor U3804 (N_3804,N_1806,N_2120);
and U3805 (N_3805,N_814,N_800);
nor U3806 (N_3806,N_1480,N_212);
and U3807 (N_3807,N_1206,N_1755);
or U3808 (N_3808,N_2455,N_8);
or U3809 (N_3809,N_10,N_180);
and U3810 (N_3810,N_1404,N_283);
and U3811 (N_3811,N_2235,N_2176);
nand U3812 (N_3812,N_1173,N_1178);
nor U3813 (N_3813,N_1921,N_586);
nand U3814 (N_3814,N_307,N_777);
and U3815 (N_3815,N_1848,N_2422);
nor U3816 (N_3816,N_1622,N_11);
nand U3817 (N_3817,N_2366,N_350);
nor U3818 (N_3818,N_330,N_1270);
or U3819 (N_3819,N_606,N_1088);
and U3820 (N_3820,N_2104,N_598);
nor U3821 (N_3821,N_1461,N_2054);
or U3822 (N_3822,N_355,N_983);
and U3823 (N_3823,N_1407,N_1296);
and U3824 (N_3824,N_1200,N_805);
nand U3825 (N_3825,N_357,N_755);
or U3826 (N_3826,N_2102,N_190);
or U3827 (N_3827,N_1781,N_1349);
nand U3828 (N_3828,N_1353,N_579);
xor U3829 (N_3829,N_865,N_1068);
nor U3830 (N_3830,N_2123,N_666);
nor U3831 (N_3831,N_2239,N_1316);
and U3832 (N_3832,N_1705,N_2098);
and U3833 (N_3833,N_1580,N_1691);
nor U3834 (N_3834,N_726,N_1254);
nand U3835 (N_3835,N_190,N_204);
and U3836 (N_3836,N_1598,N_33);
nor U3837 (N_3837,N_1665,N_2006);
nand U3838 (N_3838,N_1680,N_520);
or U3839 (N_3839,N_1562,N_2209);
and U3840 (N_3840,N_214,N_2302);
or U3841 (N_3841,N_196,N_1533);
or U3842 (N_3842,N_719,N_93);
and U3843 (N_3843,N_2053,N_1704);
or U3844 (N_3844,N_782,N_85);
and U3845 (N_3845,N_2264,N_1600);
or U3846 (N_3846,N_257,N_539);
or U3847 (N_3847,N_1409,N_1924);
nand U3848 (N_3848,N_1401,N_697);
or U3849 (N_3849,N_1876,N_802);
nand U3850 (N_3850,N_359,N_1597);
nand U3851 (N_3851,N_285,N_1449);
and U3852 (N_3852,N_1798,N_2214);
or U3853 (N_3853,N_1140,N_1605);
or U3854 (N_3854,N_1728,N_1900);
or U3855 (N_3855,N_1863,N_453);
or U3856 (N_3856,N_855,N_1943);
and U3857 (N_3857,N_2307,N_2456);
nand U3858 (N_3858,N_105,N_2289);
nor U3859 (N_3859,N_2295,N_562);
and U3860 (N_3860,N_1100,N_393);
xnor U3861 (N_3861,N_1123,N_2372);
nor U3862 (N_3862,N_512,N_1319);
or U3863 (N_3863,N_474,N_552);
and U3864 (N_3864,N_1585,N_48);
and U3865 (N_3865,N_596,N_840);
or U3866 (N_3866,N_466,N_1523);
nor U3867 (N_3867,N_2493,N_514);
and U3868 (N_3868,N_2156,N_87);
and U3869 (N_3869,N_39,N_1937);
nand U3870 (N_3870,N_2319,N_1915);
or U3871 (N_3871,N_348,N_664);
and U3872 (N_3872,N_38,N_1435);
nor U3873 (N_3873,N_117,N_866);
and U3874 (N_3874,N_1060,N_2219);
nor U3875 (N_3875,N_1529,N_2402);
and U3876 (N_3876,N_1906,N_287);
or U3877 (N_3877,N_1955,N_2436);
and U3878 (N_3878,N_1127,N_1872);
nand U3879 (N_3879,N_433,N_683);
nor U3880 (N_3880,N_1781,N_343);
and U3881 (N_3881,N_295,N_1388);
xor U3882 (N_3882,N_813,N_880);
nand U3883 (N_3883,N_875,N_570);
or U3884 (N_3884,N_2334,N_568);
nor U3885 (N_3885,N_2376,N_738);
and U3886 (N_3886,N_1062,N_846);
nor U3887 (N_3887,N_550,N_365);
or U3888 (N_3888,N_2460,N_1454);
and U3889 (N_3889,N_1495,N_24);
nand U3890 (N_3890,N_1386,N_579);
or U3891 (N_3891,N_1205,N_1780);
nand U3892 (N_3892,N_1492,N_1931);
or U3893 (N_3893,N_2021,N_2438);
and U3894 (N_3894,N_1145,N_1641);
and U3895 (N_3895,N_354,N_1347);
nand U3896 (N_3896,N_2267,N_90);
nand U3897 (N_3897,N_1676,N_34);
nand U3898 (N_3898,N_417,N_1632);
nor U3899 (N_3899,N_1731,N_99);
nand U3900 (N_3900,N_562,N_1745);
nand U3901 (N_3901,N_110,N_230);
or U3902 (N_3902,N_1016,N_925);
nor U3903 (N_3903,N_1490,N_819);
and U3904 (N_3904,N_140,N_151);
and U3905 (N_3905,N_2283,N_476);
or U3906 (N_3906,N_2306,N_606);
and U3907 (N_3907,N_1964,N_1746);
nor U3908 (N_3908,N_552,N_110);
and U3909 (N_3909,N_886,N_1914);
nand U3910 (N_3910,N_107,N_2328);
and U3911 (N_3911,N_1246,N_171);
or U3912 (N_3912,N_606,N_1922);
nor U3913 (N_3913,N_192,N_1685);
and U3914 (N_3914,N_796,N_1094);
nor U3915 (N_3915,N_635,N_1188);
nor U3916 (N_3916,N_178,N_1027);
nand U3917 (N_3917,N_1753,N_195);
nor U3918 (N_3918,N_2349,N_798);
or U3919 (N_3919,N_619,N_1808);
and U3920 (N_3920,N_1214,N_277);
nor U3921 (N_3921,N_1880,N_2362);
nor U3922 (N_3922,N_1752,N_996);
nand U3923 (N_3923,N_1946,N_1774);
or U3924 (N_3924,N_2205,N_931);
and U3925 (N_3925,N_1436,N_1692);
nor U3926 (N_3926,N_2391,N_348);
nor U3927 (N_3927,N_201,N_560);
nand U3928 (N_3928,N_728,N_2155);
nand U3929 (N_3929,N_321,N_1916);
and U3930 (N_3930,N_446,N_1401);
nand U3931 (N_3931,N_789,N_1260);
and U3932 (N_3932,N_399,N_1211);
nor U3933 (N_3933,N_2090,N_1470);
and U3934 (N_3934,N_2497,N_155);
or U3935 (N_3935,N_2467,N_232);
or U3936 (N_3936,N_1824,N_1909);
xnor U3937 (N_3937,N_1909,N_540);
nand U3938 (N_3938,N_403,N_123);
nand U3939 (N_3939,N_1276,N_1799);
and U3940 (N_3940,N_1020,N_141);
nand U3941 (N_3941,N_1637,N_2174);
nor U3942 (N_3942,N_269,N_309);
nand U3943 (N_3943,N_2141,N_475);
nor U3944 (N_3944,N_1492,N_1422);
nand U3945 (N_3945,N_1800,N_1975);
nand U3946 (N_3946,N_379,N_981);
or U3947 (N_3947,N_277,N_1249);
or U3948 (N_3948,N_467,N_232);
nor U3949 (N_3949,N_1119,N_751);
xnor U3950 (N_3950,N_785,N_1357);
nand U3951 (N_3951,N_1131,N_2351);
nand U3952 (N_3952,N_2138,N_261);
nand U3953 (N_3953,N_202,N_1466);
and U3954 (N_3954,N_1953,N_1960);
and U3955 (N_3955,N_859,N_1614);
or U3956 (N_3956,N_1366,N_2103);
nor U3957 (N_3957,N_1121,N_1842);
and U3958 (N_3958,N_116,N_2299);
and U3959 (N_3959,N_2294,N_1849);
or U3960 (N_3960,N_1900,N_49);
nor U3961 (N_3961,N_2347,N_470);
and U3962 (N_3962,N_449,N_1694);
or U3963 (N_3963,N_1967,N_1309);
and U3964 (N_3964,N_2353,N_2308);
or U3965 (N_3965,N_437,N_1168);
and U3966 (N_3966,N_1693,N_2400);
or U3967 (N_3967,N_1545,N_353);
or U3968 (N_3968,N_1136,N_175);
nor U3969 (N_3969,N_1125,N_1751);
or U3970 (N_3970,N_272,N_1014);
and U3971 (N_3971,N_1601,N_415);
nor U3972 (N_3972,N_2355,N_841);
and U3973 (N_3973,N_1303,N_868);
or U3974 (N_3974,N_1095,N_1908);
nand U3975 (N_3975,N_1068,N_66);
or U3976 (N_3976,N_219,N_2486);
nor U3977 (N_3977,N_196,N_641);
and U3978 (N_3978,N_2462,N_1160);
and U3979 (N_3979,N_312,N_2413);
or U3980 (N_3980,N_651,N_1535);
or U3981 (N_3981,N_1420,N_342);
or U3982 (N_3982,N_701,N_2120);
and U3983 (N_3983,N_263,N_1842);
nor U3984 (N_3984,N_117,N_368);
nor U3985 (N_3985,N_1068,N_706);
nor U3986 (N_3986,N_1179,N_673);
nor U3987 (N_3987,N_2229,N_80);
or U3988 (N_3988,N_1276,N_1280);
or U3989 (N_3989,N_1135,N_1450);
nand U3990 (N_3990,N_1762,N_1052);
and U3991 (N_3991,N_443,N_1959);
or U3992 (N_3992,N_781,N_2280);
nor U3993 (N_3993,N_1303,N_1569);
nand U3994 (N_3994,N_1533,N_812);
or U3995 (N_3995,N_485,N_490);
nand U3996 (N_3996,N_95,N_1712);
or U3997 (N_3997,N_1358,N_2401);
or U3998 (N_3998,N_1316,N_2450);
or U3999 (N_3999,N_84,N_1214);
nor U4000 (N_4000,N_2241,N_259);
or U4001 (N_4001,N_938,N_596);
nand U4002 (N_4002,N_2177,N_477);
and U4003 (N_4003,N_1401,N_2271);
or U4004 (N_4004,N_2105,N_1920);
or U4005 (N_4005,N_1366,N_2171);
nand U4006 (N_4006,N_549,N_885);
nand U4007 (N_4007,N_724,N_871);
and U4008 (N_4008,N_1922,N_1340);
nand U4009 (N_4009,N_368,N_2209);
nand U4010 (N_4010,N_1682,N_2211);
or U4011 (N_4011,N_1142,N_1947);
and U4012 (N_4012,N_1487,N_2162);
nor U4013 (N_4013,N_2394,N_1723);
nor U4014 (N_4014,N_1237,N_1235);
xor U4015 (N_4015,N_1414,N_1667);
or U4016 (N_4016,N_847,N_1725);
nand U4017 (N_4017,N_2246,N_1555);
and U4018 (N_4018,N_828,N_443);
or U4019 (N_4019,N_1129,N_1197);
and U4020 (N_4020,N_910,N_1461);
nor U4021 (N_4021,N_2450,N_1547);
or U4022 (N_4022,N_1775,N_1451);
and U4023 (N_4023,N_2003,N_1997);
and U4024 (N_4024,N_1616,N_2466);
and U4025 (N_4025,N_1177,N_2353);
nand U4026 (N_4026,N_1860,N_454);
nor U4027 (N_4027,N_495,N_897);
nand U4028 (N_4028,N_52,N_854);
and U4029 (N_4029,N_887,N_2262);
and U4030 (N_4030,N_197,N_1979);
and U4031 (N_4031,N_2393,N_1751);
and U4032 (N_4032,N_750,N_638);
and U4033 (N_4033,N_1228,N_1857);
nand U4034 (N_4034,N_856,N_2289);
nor U4035 (N_4035,N_858,N_1261);
nand U4036 (N_4036,N_1957,N_2012);
or U4037 (N_4037,N_753,N_1119);
nor U4038 (N_4038,N_1422,N_2442);
and U4039 (N_4039,N_2226,N_49);
or U4040 (N_4040,N_132,N_84);
nor U4041 (N_4041,N_550,N_1927);
nand U4042 (N_4042,N_703,N_1950);
nand U4043 (N_4043,N_1796,N_1961);
or U4044 (N_4044,N_2040,N_2187);
and U4045 (N_4045,N_242,N_1163);
nand U4046 (N_4046,N_2112,N_1969);
and U4047 (N_4047,N_622,N_75);
nor U4048 (N_4048,N_1894,N_796);
and U4049 (N_4049,N_1963,N_2486);
or U4050 (N_4050,N_1400,N_539);
nand U4051 (N_4051,N_1702,N_777);
and U4052 (N_4052,N_1656,N_682);
nor U4053 (N_4053,N_2108,N_1948);
nand U4054 (N_4054,N_1211,N_601);
and U4055 (N_4055,N_2183,N_218);
or U4056 (N_4056,N_1128,N_826);
or U4057 (N_4057,N_1608,N_574);
nor U4058 (N_4058,N_1158,N_143);
or U4059 (N_4059,N_1798,N_2229);
nand U4060 (N_4060,N_2469,N_570);
nor U4061 (N_4061,N_380,N_2230);
or U4062 (N_4062,N_62,N_1719);
nand U4063 (N_4063,N_1103,N_1711);
nor U4064 (N_4064,N_2359,N_1569);
nor U4065 (N_4065,N_2158,N_630);
and U4066 (N_4066,N_4,N_524);
or U4067 (N_4067,N_348,N_1546);
or U4068 (N_4068,N_1422,N_1811);
nor U4069 (N_4069,N_54,N_1180);
and U4070 (N_4070,N_641,N_1208);
nor U4071 (N_4071,N_1534,N_2247);
or U4072 (N_4072,N_339,N_1061);
nor U4073 (N_4073,N_1820,N_369);
and U4074 (N_4074,N_2360,N_1066);
and U4075 (N_4075,N_1056,N_477);
or U4076 (N_4076,N_151,N_891);
nor U4077 (N_4077,N_1491,N_818);
nor U4078 (N_4078,N_2149,N_363);
nand U4079 (N_4079,N_2362,N_1465);
nor U4080 (N_4080,N_1066,N_83);
and U4081 (N_4081,N_2052,N_1502);
nor U4082 (N_4082,N_1941,N_137);
and U4083 (N_4083,N_1197,N_2079);
nor U4084 (N_4084,N_1091,N_2040);
or U4085 (N_4085,N_1609,N_1410);
nor U4086 (N_4086,N_1147,N_158);
nor U4087 (N_4087,N_2194,N_2411);
and U4088 (N_4088,N_2076,N_1404);
or U4089 (N_4089,N_1198,N_525);
and U4090 (N_4090,N_1959,N_1968);
and U4091 (N_4091,N_1414,N_172);
and U4092 (N_4092,N_929,N_78);
nand U4093 (N_4093,N_1097,N_62);
or U4094 (N_4094,N_454,N_5);
nor U4095 (N_4095,N_1945,N_1912);
nand U4096 (N_4096,N_1393,N_774);
and U4097 (N_4097,N_2285,N_542);
nand U4098 (N_4098,N_708,N_374);
and U4099 (N_4099,N_1449,N_345);
nand U4100 (N_4100,N_1762,N_547);
nor U4101 (N_4101,N_442,N_237);
nor U4102 (N_4102,N_602,N_1621);
nor U4103 (N_4103,N_1738,N_1037);
and U4104 (N_4104,N_2013,N_1408);
and U4105 (N_4105,N_1491,N_745);
and U4106 (N_4106,N_2069,N_46);
or U4107 (N_4107,N_1622,N_2484);
and U4108 (N_4108,N_784,N_822);
or U4109 (N_4109,N_917,N_51);
or U4110 (N_4110,N_606,N_736);
nor U4111 (N_4111,N_1569,N_2337);
or U4112 (N_4112,N_263,N_446);
or U4113 (N_4113,N_1094,N_2102);
nand U4114 (N_4114,N_1388,N_1182);
nand U4115 (N_4115,N_242,N_1509);
and U4116 (N_4116,N_164,N_394);
and U4117 (N_4117,N_2140,N_631);
nor U4118 (N_4118,N_2300,N_1876);
nand U4119 (N_4119,N_215,N_1960);
or U4120 (N_4120,N_2222,N_2310);
and U4121 (N_4121,N_622,N_2251);
xnor U4122 (N_4122,N_149,N_874);
or U4123 (N_4123,N_304,N_1213);
nand U4124 (N_4124,N_1672,N_54);
and U4125 (N_4125,N_1110,N_1042);
and U4126 (N_4126,N_1637,N_945);
or U4127 (N_4127,N_1696,N_599);
and U4128 (N_4128,N_500,N_1661);
nand U4129 (N_4129,N_1054,N_1052);
nand U4130 (N_4130,N_843,N_1434);
or U4131 (N_4131,N_2316,N_48);
nor U4132 (N_4132,N_1803,N_529);
and U4133 (N_4133,N_1319,N_525);
nor U4134 (N_4134,N_2391,N_938);
nor U4135 (N_4135,N_184,N_1325);
nand U4136 (N_4136,N_1954,N_1065);
or U4137 (N_4137,N_761,N_954);
nand U4138 (N_4138,N_2070,N_916);
nand U4139 (N_4139,N_618,N_2417);
nand U4140 (N_4140,N_1339,N_1817);
nand U4141 (N_4141,N_919,N_2358);
nor U4142 (N_4142,N_2306,N_1195);
nand U4143 (N_4143,N_292,N_1429);
nor U4144 (N_4144,N_749,N_1184);
or U4145 (N_4145,N_1786,N_823);
nand U4146 (N_4146,N_891,N_1991);
and U4147 (N_4147,N_936,N_2233);
nor U4148 (N_4148,N_1770,N_1905);
nand U4149 (N_4149,N_1573,N_724);
or U4150 (N_4150,N_2057,N_1246);
or U4151 (N_4151,N_2254,N_1159);
nand U4152 (N_4152,N_1021,N_656);
or U4153 (N_4153,N_567,N_708);
nor U4154 (N_4154,N_61,N_929);
nor U4155 (N_4155,N_2046,N_1931);
nor U4156 (N_4156,N_2473,N_1147);
nor U4157 (N_4157,N_1504,N_1982);
nand U4158 (N_4158,N_1383,N_887);
or U4159 (N_4159,N_2133,N_564);
and U4160 (N_4160,N_1836,N_122);
or U4161 (N_4161,N_267,N_1085);
or U4162 (N_4162,N_2095,N_1767);
nand U4163 (N_4163,N_156,N_568);
and U4164 (N_4164,N_1203,N_1217);
nor U4165 (N_4165,N_2060,N_1033);
nand U4166 (N_4166,N_994,N_915);
nand U4167 (N_4167,N_1605,N_637);
xor U4168 (N_4168,N_1854,N_1389);
nor U4169 (N_4169,N_1413,N_1511);
and U4170 (N_4170,N_634,N_865);
nor U4171 (N_4171,N_964,N_1150);
or U4172 (N_4172,N_1988,N_1341);
and U4173 (N_4173,N_278,N_1202);
or U4174 (N_4174,N_1303,N_997);
or U4175 (N_4175,N_2443,N_775);
nand U4176 (N_4176,N_2172,N_1586);
nor U4177 (N_4177,N_2249,N_2309);
and U4178 (N_4178,N_2253,N_1518);
or U4179 (N_4179,N_1610,N_1729);
and U4180 (N_4180,N_1845,N_869);
and U4181 (N_4181,N_1552,N_1938);
nand U4182 (N_4182,N_998,N_2222);
nand U4183 (N_4183,N_354,N_733);
and U4184 (N_4184,N_2068,N_1515);
and U4185 (N_4185,N_1944,N_2063);
nor U4186 (N_4186,N_876,N_1537);
or U4187 (N_4187,N_1546,N_1109);
nor U4188 (N_4188,N_2137,N_313);
or U4189 (N_4189,N_1859,N_561);
and U4190 (N_4190,N_1406,N_786);
nand U4191 (N_4191,N_1580,N_1050);
and U4192 (N_4192,N_1018,N_1757);
nor U4193 (N_4193,N_1649,N_232);
nand U4194 (N_4194,N_835,N_1229);
xor U4195 (N_4195,N_1406,N_317);
or U4196 (N_4196,N_502,N_394);
or U4197 (N_4197,N_199,N_2019);
or U4198 (N_4198,N_291,N_149);
or U4199 (N_4199,N_56,N_242);
and U4200 (N_4200,N_425,N_1034);
xor U4201 (N_4201,N_472,N_1910);
nor U4202 (N_4202,N_19,N_773);
nand U4203 (N_4203,N_816,N_288);
or U4204 (N_4204,N_1619,N_1920);
and U4205 (N_4205,N_576,N_212);
xnor U4206 (N_4206,N_550,N_2371);
and U4207 (N_4207,N_1967,N_2311);
or U4208 (N_4208,N_264,N_1489);
nor U4209 (N_4209,N_1267,N_677);
or U4210 (N_4210,N_2280,N_103);
nor U4211 (N_4211,N_812,N_136);
nand U4212 (N_4212,N_774,N_2222);
nor U4213 (N_4213,N_2265,N_763);
nor U4214 (N_4214,N_470,N_2201);
nor U4215 (N_4215,N_674,N_651);
or U4216 (N_4216,N_1038,N_95);
or U4217 (N_4217,N_1230,N_81);
or U4218 (N_4218,N_1019,N_1151);
and U4219 (N_4219,N_1237,N_901);
and U4220 (N_4220,N_1408,N_526);
or U4221 (N_4221,N_793,N_1619);
and U4222 (N_4222,N_1119,N_2254);
and U4223 (N_4223,N_2360,N_1025);
nand U4224 (N_4224,N_1543,N_1797);
nand U4225 (N_4225,N_1052,N_622);
nor U4226 (N_4226,N_2338,N_685);
or U4227 (N_4227,N_2251,N_1221);
or U4228 (N_4228,N_1954,N_1171);
or U4229 (N_4229,N_590,N_1104);
or U4230 (N_4230,N_1342,N_857);
and U4231 (N_4231,N_6,N_2413);
or U4232 (N_4232,N_1348,N_399);
and U4233 (N_4233,N_1622,N_2326);
or U4234 (N_4234,N_2268,N_1677);
or U4235 (N_4235,N_2082,N_125);
or U4236 (N_4236,N_737,N_1374);
and U4237 (N_4237,N_131,N_956);
nand U4238 (N_4238,N_2299,N_449);
or U4239 (N_4239,N_998,N_6);
nand U4240 (N_4240,N_1173,N_243);
nor U4241 (N_4241,N_1700,N_516);
and U4242 (N_4242,N_1467,N_1631);
and U4243 (N_4243,N_1424,N_741);
xnor U4244 (N_4244,N_251,N_1211);
or U4245 (N_4245,N_1196,N_2369);
or U4246 (N_4246,N_701,N_2354);
and U4247 (N_4247,N_915,N_916);
or U4248 (N_4248,N_615,N_945);
and U4249 (N_4249,N_1606,N_1376);
or U4250 (N_4250,N_307,N_2063);
nand U4251 (N_4251,N_852,N_2281);
and U4252 (N_4252,N_326,N_44);
nand U4253 (N_4253,N_1124,N_2183);
and U4254 (N_4254,N_621,N_2024);
and U4255 (N_4255,N_763,N_953);
xnor U4256 (N_4256,N_151,N_754);
and U4257 (N_4257,N_1245,N_71);
or U4258 (N_4258,N_2335,N_1964);
or U4259 (N_4259,N_1148,N_1324);
and U4260 (N_4260,N_1185,N_2240);
nor U4261 (N_4261,N_1285,N_2278);
and U4262 (N_4262,N_272,N_2130);
and U4263 (N_4263,N_1195,N_2331);
and U4264 (N_4264,N_1098,N_1384);
nand U4265 (N_4265,N_533,N_809);
and U4266 (N_4266,N_1170,N_2181);
nand U4267 (N_4267,N_252,N_1148);
nor U4268 (N_4268,N_2401,N_2209);
and U4269 (N_4269,N_713,N_2150);
or U4270 (N_4270,N_1140,N_754);
and U4271 (N_4271,N_510,N_838);
xor U4272 (N_4272,N_2448,N_1586);
or U4273 (N_4273,N_1181,N_1304);
nor U4274 (N_4274,N_2482,N_2265);
and U4275 (N_4275,N_347,N_109);
nor U4276 (N_4276,N_2218,N_2249);
and U4277 (N_4277,N_399,N_552);
or U4278 (N_4278,N_1718,N_589);
and U4279 (N_4279,N_2301,N_495);
and U4280 (N_4280,N_1600,N_1880);
and U4281 (N_4281,N_1034,N_1549);
nor U4282 (N_4282,N_2155,N_1052);
or U4283 (N_4283,N_96,N_265);
or U4284 (N_4284,N_1256,N_366);
nor U4285 (N_4285,N_469,N_1113);
xor U4286 (N_4286,N_1355,N_1353);
or U4287 (N_4287,N_503,N_2015);
nor U4288 (N_4288,N_137,N_1927);
nand U4289 (N_4289,N_2198,N_135);
or U4290 (N_4290,N_1844,N_271);
nor U4291 (N_4291,N_1333,N_811);
nor U4292 (N_4292,N_585,N_464);
or U4293 (N_4293,N_1037,N_814);
and U4294 (N_4294,N_458,N_521);
and U4295 (N_4295,N_2074,N_149);
nor U4296 (N_4296,N_319,N_1058);
nor U4297 (N_4297,N_1117,N_1518);
nand U4298 (N_4298,N_1918,N_2496);
and U4299 (N_4299,N_1564,N_444);
nor U4300 (N_4300,N_103,N_1416);
and U4301 (N_4301,N_1409,N_18);
and U4302 (N_4302,N_1503,N_1803);
nor U4303 (N_4303,N_232,N_1130);
nor U4304 (N_4304,N_2351,N_1550);
nor U4305 (N_4305,N_1217,N_246);
nand U4306 (N_4306,N_1971,N_283);
nor U4307 (N_4307,N_1040,N_1331);
xor U4308 (N_4308,N_1674,N_1147);
or U4309 (N_4309,N_1890,N_767);
or U4310 (N_4310,N_2027,N_372);
and U4311 (N_4311,N_1046,N_1181);
or U4312 (N_4312,N_329,N_1851);
nand U4313 (N_4313,N_1770,N_1147);
nand U4314 (N_4314,N_362,N_492);
or U4315 (N_4315,N_1959,N_1908);
nand U4316 (N_4316,N_1449,N_247);
or U4317 (N_4317,N_269,N_201);
or U4318 (N_4318,N_82,N_1018);
or U4319 (N_4319,N_1688,N_2098);
or U4320 (N_4320,N_245,N_1467);
and U4321 (N_4321,N_964,N_1173);
or U4322 (N_4322,N_1932,N_314);
and U4323 (N_4323,N_1857,N_786);
or U4324 (N_4324,N_1412,N_886);
and U4325 (N_4325,N_195,N_501);
nand U4326 (N_4326,N_341,N_656);
and U4327 (N_4327,N_1555,N_1250);
nand U4328 (N_4328,N_843,N_1076);
xor U4329 (N_4329,N_1897,N_1449);
or U4330 (N_4330,N_986,N_1381);
or U4331 (N_4331,N_623,N_289);
or U4332 (N_4332,N_751,N_62);
xnor U4333 (N_4333,N_458,N_1667);
nor U4334 (N_4334,N_599,N_1394);
or U4335 (N_4335,N_512,N_2080);
or U4336 (N_4336,N_513,N_1161);
nand U4337 (N_4337,N_1574,N_918);
and U4338 (N_4338,N_1428,N_2334);
or U4339 (N_4339,N_2341,N_2261);
or U4340 (N_4340,N_1812,N_791);
nor U4341 (N_4341,N_1798,N_1259);
nor U4342 (N_4342,N_1988,N_199);
and U4343 (N_4343,N_2188,N_1524);
or U4344 (N_4344,N_250,N_997);
or U4345 (N_4345,N_1921,N_2185);
nor U4346 (N_4346,N_2357,N_2182);
or U4347 (N_4347,N_1543,N_833);
and U4348 (N_4348,N_1357,N_2052);
nor U4349 (N_4349,N_331,N_322);
or U4350 (N_4350,N_2044,N_244);
and U4351 (N_4351,N_145,N_2059);
and U4352 (N_4352,N_1781,N_254);
nor U4353 (N_4353,N_1141,N_1859);
nand U4354 (N_4354,N_2262,N_1035);
nor U4355 (N_4355,N_345,N_2397);
nand U4356 (N_4356,N_2007,N_799);
nand U4357 (N_4357,N_2221,N_716);
or U4358 (N_4358,N_916,N_696);
nor U4359 (N_4359,N_30,N_809);
or U4360 (N_4360,N_2435,N_1357);
or U4361 (N_4361,N_239,N_2001);
nand U4362 (N_4362,N_120,N_2342);
nand U4363 (N_4363,N_926,N_1976);
or U4364 (N_4364,N_552,N_71);
nand U4365 (N_4365,N_2472,N_1859);
nor U4366 (N_4366,N_145,N_691);
nor U4367 (N_4367,N_773,N_910);
and U4368 (N_4368,N_781,N_1706);
nor U4369 (N_4369,N_2384,N_675);
and U4370 (N_4370,N_745,N_1508);
and U4371 (N_4371,N_98,N_797);
nand U4372 (N_4372,N_2483,N_458);
and U4373 (N_4373,N_521,N_1363);
nand U4374 (N_4374,N_42,N_825);
nand U4375 (N_4375,N_363,N_1133);
or U4376 (N_4376,N_2365,N_1639);
and U4377 (N_4377,N_971,N_1655);
and U4378 (N_4378,N_1618,N_2443);
nor U4379 (N_4379,N_2054,N_816);
or U4380 (N_4380,N_163,N_1261);
nand U4381 (N_4381,N_129,N_1731);
and U4382 (N_4382,N_1951,N_537);
and U4383 (N_4383,N_631,N_571);
nand U4384 (N_4384,N_731,N_1182);
nand U4385 (N_4385,N_1504,N_436);
nand U4386 (N_4386,N_76,N_735);
or U4387 (N_4387,N_180,N_2171);
and U4388 (N_4388,N_1251,N_1840);
and U4389 (N_4389,N_747,N_1169);
and U4390 (N_4390,N_551,N_562);
or U4391 (N_4391,N_1863,N_1709);
nand U4392 (N_4392,N_1515,N_1329);
nor U4393 (N_4393,N_652,N_586);
nand U4394 (N_4394,N_2482,N_2341);
or U4395 (N_4395,N_542,N_832);
nor U4396 (N_4396,N_893,N_1451);
or U4397 (N_4397,N_1799,N_862);
or U4398 (N_4398,N_1112,N_937);
or U4399 (N_4399,N_261,N_1440);
or U4400 (N_4400,N_1749,N_2243);
nor U4401 (N_4401,N_300,N_215);
xnor U4402 (N_4402,N_137,N_1486);
and U4403 (N_4403,N_1581,N_987);
and U4404 (N_4404,N_1438,N_1503);
nor U4405 (N_4405,N_923,N_1479);
and U4406 (N_4406,N_1445,N_1654);
nand U4407 (N_4407,N_2109,N_658);
nor U4408 (N_4408,N_109,N_251);
or U4409 (N_4409,N_2236,N_1635);
nand U4410 (N_4410,N_1279,N_204);
nand U4411 (N_4411,N_574,N_911);
and U4412 (N_4412,N_745,N_1343);
nor U4413 (N_4413,N_1491,N_546);
and U4414 (N_4414,N_2370,N_492);
nand U4415 (N_4415,N_2351,N_1054);
nor U4416 (N_4416,N_2463,N_63);
and U4417 (N_4417,N_1491,N_2270);
nor U4418 (N_4418,N_2497,N_2440);
nor U4419 (N_4419,N_1175,N_159);
nor U4420 (N_4420,N_908,N_696);
or U4421 (N_4421,N_961,N_118);
and U4422 (N_4422,N_2047,N_1513);
or U4423 (N_4423,N_2049,N_453);
and U4424 (N_4424,N_1733,N_2145);
nor U4425 (N_4425,N_1142,N_186);
nor U4426 (N_4426,N_1527,N_319);
nand U4427 (N_4427,N_1608,N_1946);
nand U4428 (N_4428,N_1620,N_1910);
nand U4429 (N_4429,N_2070,N_296);
and U4430 (N_4430,N_426,N_975);
or U4431 (N_4431,N_220,N_2330);
nand U4432 (N_4432,N_456,N_821);
and U4433 (N_4433,N_314,N_671);
and U4434 (N_4434,N_2321,N_2006);
nand U4435 (N_4435,N_1956,N_2159);
nor U4436 (N_4436,N_1722,N_405);
nor U4437 (N_4437,N_1897,N_903);
nor U4438 (N_4438,N_83,N_2090);
nand U4439 (N_4439,N_872,N_1284);
or U4440 (N_4440,N_1207,N_1546);
or U4441 (N_4441,N_739,N_843);
xnor U4442 (N_4442,N_1718,N_124);
nor U4443 (N_4443,N_825,N_1113);
and U4444 (N_4444,N_1894,N_490);
nor U4445 (N_4445,N_1166,N_1023);
or U4446 (N_4446,N_1217,N_238);
nand U4447 (N_4447,N_1413,N_8);
or U4448 (N_4448,N_110,N_2137);
xnor U4449 (N_4449,N_1581,N_839);
nor U4450 (N_4450,N_1080,N_53);
nor U4451 (N_4451,N_1566,N_772);
or U4452 (N_4452,N_1917,N_2411);
and U4453 (N_4453,N_1765,N_777);
and U4454 (N_4454,N_298,N_663);
and U4455 (N_4455,N_685,N_182);
or U4456 (N_4456,N_1493,N_728);
or U4457 (N_4457,N_767,N_1372);
or U4458 (N_4458,N_2261,N_2052);
nand U4459 (N_4459,N_2220,N_2403);
nor U4460 (N_4460,N_1948,N_590);
or U4461 (N_4461,N_656,N_826);
xnor U4462 (N_4462,N_1774,N_78);
or U4463 (N_4463,N_281,N_1049);
or U4464 (N_4464,N_411,N_1493);
and U4465 (N_4465,N_2022,N_925);
nand U4466 (N_4466,N_1434,N_1305);
nor U4467 (N_4467,N_689,N_1076);
nand U4468 (N_4468,N_197,N_2209);
nor U4469 (N_4469,N_241,N_1273);
nor U4470 (N_4470,N_195,N_1191);
nand U4471 (N_4471,N_1652,N_1912);
nand U4472 (N_4472,N_1371,N_1017);
nand U4473 (N_4473,N_747,N_500);
and U4474 (N_4474,N_369,N_1013);
nand U4475 (N_4475,N_1533,N_2100);
nand U4476 (N_4476,N_1927,N_1432);
nor U4477 (N_4477,N_2220,N_1353);
nor U4478 (N_4478,N_1532,N_139);
and U4479 (N_4479,N_1387,N_1205);
or U4480 (N_4480,N_647,N_379);
or U4481 (N_4481,N_154,N_290);
or U4482 (N_4482,N_2475,N_1899);
nand U4483 (N_4483,N_2039,N_1001);
and U4484 (N_4484,N_337,N_1494);
and U4485 (N_4485,N_1219,N_819);
or U4486 (N_4486,N_995,N_1036);
or U4487 (N_4487,N_2256,N_445);
nor U4488 (N_4488,N_1942,N_527);
nor U4489 (N_4489,N_963,N_997);
nand U4490 (N_4490,N_1928,N_1755);
nand U4491 (N_4491,N_1721,N_139);
or U4492 (N_4492,N_2343,N_1098);
and U4493 (N_4493,N_322,N_1939);
nand U4494 (N_4494,N_2204,N_410);
nor U4495 (N_4495,N_2198,N_1404);
nor U4496 (N_4496,N_2384,N_908);
and U4497 (N_4497,N_924,N_410);
nor U4498 (N_4498,N_2080,N_656);
nand U4499 (N_4499,N_1092,N_215);
nor U4500 (N_4500,N_1946,N_124);
nor U4501 (N_4501,N_349,N_1553);
and U4502 (N_4502,N_9,N_568);
nand U4503 (N_4503,N_1049,N_554);
nand U4504 (N_4504,N_1003,N_1295);
and U4505 (N_4505,N_1567,N_1830);
nand U4506 (N_4506,N_484,N_1829);
or U4507 (N_4507,N_1865,N_742);
or U4508 (N_4508,N_2066,N_2361);
nor U4509 (N_4509,N_2272,N_253);
nor U4510 (N_4510,N_906,N_928);
nor U4511 (N_4511,N_578,N_446);
and U4512 (N_4512,N_159,N_982);
and U4513 (N_4513,N_2064,N_296);
nor U4514 (N_4514,N_1868,N_1800);
or U4515 (N_4515,N_932,N_37);
nand U4516 (N_4516,N_1238,N_2051);
and U4517 (N_4517,N_1604,N_1835);
and U4518 (N_4518,N_495,N_564);
or U4519 (N_4519,N_376,N_2342);
and U4520 (N_4520,N_1372,N_726);
and U4521 (N_4521,N_1188,N_300);
or U4522 (N_4522,N_1052,N_4);
or U4523 (N_4523,N_2349,N_1387);
and U4524 (N_4524,N_618,N_1364);
and U4525 (N_4525,N_1062,N_2140);
and U4526 (N_4526,N_621,N_2108);
nor U4527 (N_4527,N_2376,N_504);
nor U4528 (N_4528,N_1544,N_1730);
and U4529 (N_4529,N_1358,N_2353);
and U4530 (N_4530,N_1024,N_1765);
and U4531 (N_4531,N_945,N_1704);
nor U4532 (N_4532,N_1057,N_198);
or U4533 (N_4533,N_668,N_566);
nand U4534 (N_4534,N_298,N_1827);
and U4535 (N_4535,N_1361,N_1812);
nor U4536 (N_4536,N_1388,N_1595);
nor U4537 (N_4537,N_164,N_1548);
and U4538 (N_4538,N_941,N_654);
or U4539 (N_4539,N_1990,N_2464);
nor U4540 (N_4540,N_353,N_643);
nand U4541 (N_4541,N_710,N_886);
nand U4542 (N_4542,N_1785,N_63);
or U4543 (N_4543,N_2186,N_124);
nor U4544 (N_4544,N_137,N_1306);
and U4545 (N_4545,N_2019,N_66);
nand U4546 (N_4546,N_1072,N_2255);
nor U4547 (N_4547,N_242,N_1475);
or U4548 (N_4548,N_1331,N_2463);
nor U4549 (N_4549,N_1320,N_2255);
and U4550 (N_4550,N_1325,N_344);
nor U4551 (N_4551,N_541,N_1789);
nor U4552 (N_4552,N_1141,N_1889);
or U4553 (N_4553,N_301,N_2244);
nor U4554 (N_4554,N_283,N_311);
or U4555 (N_4555,N_96,N_1740);
nor U4556 (N_4556,N_791,N_2413);
nand U4557 (N_4557,N_904,N_2312);
or U4558 (N_4558,N_1595,N_1177);
or U4559 (N_4559,N_1144,N_2013);
nand U4560 (N_4560,N_1633,N_177);
nor U4561 (N_4561,N_1620,N_727);
or U4562 (N_4562,N_929,N_661);
nand U4563 (N_4563,N_1869,N_493);
nor U4564 (N_4564,N_27,N_75);
nor U4565 (N_4565,N_2180,N_2444);
and U4566 (N_4566,N_1146,N_647);
nand U4567 (N_4567,N_2382,N_65);
or U4568 (N_4568,N_1060,N_1419);
or U4569 (N_4569,N_672,N_1624);
and U4570 (N_4570,N_1643,N_1119);
or U4571 (N_4571,N_1969,N_1009);
nor U4572 (N_4572,N_1281,N_377);
and U4573 (N_4573,N_86,N_1625);
or U4574 (N_4574,N_73,N_808);
nor U4575 (N_4575,N_508,N_666);
or U4576 (N_4576,N_1035,N_164);
or U4577 (N_4577,N_2199,N_1984);
nand U4578 (N_4578,N_613,N_1549);
nand U4579 (N_4579,N_575,N_705);
nor U4580 (N_4580,N_1412,N_179);
and U4581 (N_4581,N_2493,N_347);
nor U4582 (N_4582,N_286,N_714);
nor U4583 (N_4583,N_2349,N_2170);
nand U4584 (N_4584,N_1417,N_1763);
and U4585 (N_4585,N_870,N_1539);
and U4586 (N_4586,N_1304,N_2336);
nand U4587 (N_4587,N_2197,N_1444);
nor U4588 (N_4588,N_872,N_2031);
nor U4589 (N_4589,N_2381,N_1032);
nand U4590 (N_4590,N_944,N_1670);
or U4591 (N_4591,N_1794,N_1960);
nand U4592 (N_4592,N_1816,N_525);
or U4593 (N_4593,N_351,N_1530);
and U4594 (N_4594,N_1520,N_2061);
or U4595 (N_4595,N_650,N_474);
and U4596 (N_4596,N_2315,N_1732);
or U4597 (N_4597,N_148,N_391);
and U4598 (N_4598,N_1572,N_1388);
and U4599 (N_4599,N_395,N_591);
or U4600 (N_4600,N_296,N_615);
xor U4601 (N_4601,N_1906,N_1024);
and U4602 (N_4602,N_462,N_2462);
nand U4603 (N_4603,N_2206,N_1379);
xor U4604 (N_4604,N_1713,N_1375);
or U4605 (N_4605,N_555,N_2352);
nand U4606 (N_4606,N_2304,N_1145);
and U4607 (N_4607,N_1277,N_2480);
or U4608 (N_4608,N_1991,N_1689);
or U4609 (N_4609,N_1513,N_293);
nor U4610 (N_4610,N_122,N_1384);
and U4611 (N_4611,N_47,N_975);
or U4612 (N_4612,N_490,N_1211);
nor U4613 (N_4613,N_1567,N_489);
nor U4614 (N_4614,N_738,N_1397);
nor U4615 (N_4615,N_434,N_607);
and U4616 (N_4616,N_2236,N_2029);
nor U4617 (N_4617,N_1917,N_1062);
nand U4618 (N_4618,N_1779,N_2356);
xor U4619 (N_4619,N_776,N_1244);
nand U4620 (N_4620,N_932,N_459);
nand U4621 (N_4621,N_1349,N_2455);
nand U4622 (N_4622,N_2036,N_468);
and U4623 (N_4623,N_1874,N_1831);
or U4624 (N_4624,N_2277,N_699);
and U4625 (N_4625,N_1976,N_1208);
nand U4626 (N_4626,N_2041,N_274);
nor U4627 (N_4627,N_789,N_864);
and U4628 (N_4628,N_1920,N_1271);
or U4629 (N_4629,N_522,N_1085);
nand U4630 (N_4630,N_768,N_1782);
nand U4631 (N_4631,N_2044,N_291);
nor U4632 (N_4632,N_713,N_917);
nand U4633 (N_4633,N_556,N_1670);
nor U4634 (N_4634,N_397,N_491);
and U4635 (N_4635,N_836,N_1221);
or U4636 (N_4636,N_1763,N_2434);
or U4637 (N_4637,N_602,N_1206);
nand U4638 (N_4638,N_986,N_1287);
and U4639 (N_4639,N_31,N_830);
nor U4640 (N_4640,N_1016,N_1561);
nor U4641 (N_4641,N_2168,N_325);
nand U4642 (N_4642,N_1397,N_104);
nand U4643 (N_4643,N_61,N_132);
nor U4644 (N_4644,N_340,N_283);
or U4645 (N_4645,N_641,N_2363);
nor U4646 (N_4646,N_858,N_1068);
nand U4647 (N_4647,N_1364,N_1154);
and U4648 (N_4648,N_2286,N_2271);
nand U4649 (N_4649,N_2348,N_731);
nand U4650 (N_4650,N_1737,N_738);
and U4651 (N_4651,N_2488,N_466);
or U4652 (N_4652,N_1266,N_508);
nand U4653 (N_4653,N_2497,N_103);
nor U4654 (N_4654,N_81,N_198);
xnor U4655 (N_4655,N_2209,N_1142);
nand U4656 (N_4656,N_1717,N_1027);
nand U4657 (N_4657,N_1323,N_1705);
nand U4658 (N_4658,N_1175,N_1722);
and U4659 (N_4659,N_1595,N_2167);
nor U4660 (N_4660,N_487,N_1411);
nor U4661 (N_4661,N_2297,N_1997);
and U4662 (N_4662,N_1155,N_386);
nor U4663 (N_4663,N_2099,N_787);
nand U4664 (N_4664,N_200,N_1988);
nor U4665 (N_4665,N_803,N_110);
nand U4666 (N_4666,N_111,N_452);
or U4667 (N_4667,N_2194,N_52);
nor U4668 (N_4668,N_2180,N_126);
and U4669 (N_4669,N_2335,N_363);
nor U4670 (N_4670,N_1448,N_1303);
nand U4671 (N_4671,N_621,N_2159);
nand U4672 (N_4672,N_126,N_976);
nand U4673 (N_4673,N_42,N_894);
or U4674 (N_4674,N_2423,N_1486);
and U4675 (N_4675,N_1739,N_888);
nand U4676 (N_4676,N_73,N_1);
nand U4677 (N_4677,N_1328,N_1385);
and U4678 (N_4678,N_2159,N_1868);
nor U4679 (N_4679,N_1225,N_2339);
or U4680 (N_4680,N_1327,N_59);
and U4681 (N_4681,N_1259,N_2069);
or U4682 (N_4682,N_403,N_1362);
nand U4683 (N_4683,N_955,N_825);
nand U4684 (N_4684,N_2205,N_241);
nand U4685 (N_4685,N_557,N_2331);
nor U4686 (N_4686,N_797,N_1899);
nand U4687 (N_4687,N_502,N_297);
nor U4688 (N_4688,N_1590,N_2207);
nor U4689 (N_4689,N_681,N_1134);
nand U4690 (N_4690,N_1877,N_1065);
nor U4691 (N_4691,N_1803,N_896);
nand U4692 (N_4692,N_1636,N_1010);
nand U4693 (N_4693,N_1247,N_835);
and U4694 (N_4694,N_7,N_2023);
or U4695 (N_4695,N_490,N_2311);
or U4696 (N_4696,N_1610,N_1863);
and U4697 (N_4697,N_2368,N_441);
or U4698 (N_4698,N_1158,N_1287);
and U4699 (N_4699,N_2444,N_421);
and U4700 (N_4700,N_2190,N_1548);
or U4701 (N_4701,N_2228,N_551);
or U4702 (N_4702,N_639,N_2159);
xnor U4703 (N_4703,N_2164,N_825);
nor U4704 (N_4704,N_681,N_1385);
nor U4705 (N_4705,N_2447,N_1652);
or U4706 (N_4706,N_1646,N_1774);
and U4707 (N_4707,N_1897,N_969);
nor U4708 (N_4708,N_2306,N_1352);
and U4709 (N_4709,N_786,N_643);
nor U4710 (N_4710,N_2493,N_1223);
nand U4711 (N_4711,N_354,N_757);
and U4712 (N_4712,N_1719,N_636);
and U4713 (N_4713,N_2457,N_1995);
nor U4714 (N_4714,N_2470,N_381);
and U4715 (N_4715,N_1301,N_657);
nand U4716 (N_4716,N_394,N_1770);
nor U4717 (N_4717,N_2097,N_969);
and U4718 (N_4718,N_1500,N_337);
and U4719 (N_4719,N_1809,N_9);
xor U4720 (N_4720,N_7,N_1277);
and U4721 (N_4721,N_1808,N_1611);
and U4722 (N_4722,N_1052,N_894);
and U4723 (N_4723,N_343,N_1449);
or U4724 (N_4724,N_332,N_78);
nor U4725 (N_4725,N_1392,N_502);
nor U4726 (N_4726,N_2084,N_495);
or U4727 (N_4727,N_253,N_1969);
nand U4728 (N_4728,N_645,N_1617);
or U4729 (N_4729,N_1421,N_223);
or U4730 (N_4730,N_792,N_1171);
nor U4731 (N_4731,N_2109,N_2367);
xor U4732 (N_4732,N_792,N_369);
xnor U4733 (N_4733,N_149,N_48);
nor U4734 (N_4734,N_262,N_2441);
or U4735 (N_4735,N_2314,N_1451);
or U4736 (N_4736,N_1604,N_645);
and U4737 (N_4737,N_766,N_2351);
nor U4738 (N_4738,N_1451,N_1115);
xor U4739 (N_4739,N_251,N_591);
or U4740 (N_4740,N_1293,N_2464);
or U4741 (N_4741,N_440,N_239);
nor U4742 (N_4742,N_1684,N_1577);
nand U4743 (N_4743,N_1862,N_1236);
and U4744 (N_4744,N_1706,N_1475);
nor U4745 (N_4745,N_1603,N_409);
and U4746 (N_4746,N_2301,N_1581);
nand U4747 (N_4747,N_755,N_717);
or U4748 (N_4748,N_2053,N_1199);
nand U4749 (N_4749,N_1015,N_1403);
and U4750 (N_4750,N_2198,N_2425);
or U4751 (N_4751,N_861,N_803);
nor U4752 (N_4752,N_456,N_1795);
nand U4753 (N_4753,N_1097,N_687);
nand U4754 (N_4754,N_2414,N_1183);
nand U4755 (N_4755,N_1107,N_1931);
nor U4756 (N_4756,N_976,N_1227);
and U4757 (N_4757,N_583,N_1758);
or U4758 (N_4758,N_344,N_457);
or U4759 (N_4759,N_1562,N_2154);
nor U4760 (N_4760,N_542,N_1960);
or U4761 (N_4761,N_806,N_2294);
nor U4762 (N_4762,N_2130,N_380);
or U4763 (N_4763,N_278,N_2013);
nor U4764 (N_4764,N_1890,N_950);
and U4765 (N_4765,N_532,N_1697);
nand U4766 (N_4766,N_1135,N_808);
nor U4767 (N_4767,N_1253,N_432);
nand U4768 (N_4768,N_271,N_1232);
and U4769 (N_4769,N_1425,N_40);
nor U4770 (N_4770,N_1857,N_2359);
nor U4771 (N_4771,N_2470,N_2298);
and U4772 (N_4772,N_966,N_1330);
or U4773 (N_4773,N_396,N_748);
nand U4774 (N_4774,N_97,N_891);
nor U4775 (N_4775,N_653,N_1106);
and U4776 (N_4776,N_2124,N_507);
or U4777 (N_4777,N_1501,N_2221);
or U4778 (N_4778,N_144,N_34);
nor U4779 (N_4779,N_2215,N_6);
nand U4780 (N_4780,N_1615,N_942);
or U4781 (N_4781,N_1920,N_1578);
and U4782 (N_4782,N_2334,N_2039);
nand U4783 (N_4783,N_1010,N_2113);
nand U4784 (N_4784,N_1287,N_637);
nand U4785 (N_4785,N_1633,N_1663);
nor U4786 (N_4786,N_167,N_1831);
or U4787 (N_4787,N_1431,N_1374);
or U4788 (N_4788,N_1259,N_1074);
nor U4789 (N_4789,N_1647,N_2261);
nor U4790 (N_4790,N_2446,N_1621);
nand U4791 (N_4791,N_2263,N_576);
nand U4792 (N_4792,N_433,N_1717);
or U4793 (N_4793,N_1121,N_1623);
and U4794 (N_4794,N_1272,N_1023);
nor U4795 (N_4795,N_925,N_1239);
nand U4796 (N_4796,N_1121,N_718);
or U4797 (N_4797,N_16,N_737);
or U4798 (N_4798,N_518,N_641);
nand U4799 (N_4799,N_1951,N_2047);
nor U4800 (N_4800,N_691,N_2100);
or U4801 (N_4801,N_1204,N_2341);
or U4802 (N_4802,N_2045,N_1071);
nor U4803 (N_4803,N_282,N_2485);
nor U4804 (N_4804,N_1297,N_1580);
nor U4805 (N_4805,N_1567,N_163);
nand U4806 (N_4806,N_124,N_1238);
nor U4807 (N_4807,N_2147,N_1455);
nand U4808 (N_4808,N_869,N_1581);
nor U4809 (N_4809,N_1777,N_2413);
xor U4810 (N_4810,N_757,N_2225);
or U4811 (N_4811,N_1915,N_564);
nand U4812 (N_4812,N_811,N_687);
and U4813 (N_4813,N_1782,N_793);
xor U4814 (N_4814,N_1636,N_718);
nand U4815 (N_4815,N_966,N_282);
nand U4816 (N_4816,N_1653,N_243);
or U4817 (N_4817,N_490,N_279);
and U4818 (N_4818,N_1462,N_990);
nand U4819 (N_4819,N_1966,N_1089);
xnor U4820 (N_4820,N_1738,N_749);
or U4821 (N_4821,N_1535,N_1550);
or U4822 (N_4822,N_1798,N_451);
and U4823 (N_4823,N_1620,N_1608);
and U4824 (N_4824,N_1447,N_986);
and U4825 (N_4825,N_31,N_1881);
or U4826 (N_4826,N_287,N_196);
and U4827 (N_4827,N_1580,N_976);
nand U4828 (N_4828,N_881,N_1872);
or U4829 (N_4829,N_1256,N_2136);
or U4830 (N_4830,N_1640,N_734);
or U4831 (N_4831,N_2081,N_2037);
nor U4832 (N_4832,N_894,N_2066);
nand U4833 (N_4833,N_660,N_136);
nand U4834 (N_4834,N_719,N_635);
and U4835 (N_4835,N_2497,N_2371);
nor U4836 (N_4836,N_1823,N_2378);
nor U4837 (N_4837,N_2288,N_810);
and U4838 (N_4838,N_1934,N_685);
or U4839 (N_4839,N_1348,N_2026);
nand U4840 (N_4840,N_1489,N_923);
nor U4841 (N_4841,N_1738,N_1584);
and U4842 (N_4842,N_846,N_2379);
nand U4843 (N_4843,N_1153,N_520);
or U4844 (N_4844,N_1002,N_555);
or U4845 (N_4845,N_1042,N_2321);
nand U4846 (N_4846,N_2398,N_1506);
nand U4847 (N_4847,N_1734,N_2003);
nor U4848 (N_4848,N_2188,N_470);
nor U4849 (N_4849,N_1571,N_1681);
nor U4850 (N_4850,N_1240,N_2398);
nor U4851 (N_4851,N_1807,N_249);
and U4852 (N_4852,N_633,N_290);
and U4853 (N_4853,N_2379,N_2124);
nand U4854 (N_4854,N_1122,N_1085);
or U4855 (N_4855,N_2433,N_700);
and U4856 (N_4856,N_1804,N_742);
nand U4857 (N_4857,N_1043,N_851);
xnor U4858 (N_4858,N_1500,N_63);
nor U4859 (N_4859,N_272,N_1659);
nor U4860 (N_4860,N_2145,N_1990);
and U4861 (N_4861,N_867,N_1428);
and U4862 (N_4862,N_1158,N_2301);
nand U4863 (N_4863,N_1205,N_870);
or U4864 (N_4864,N_1382,N_2279);
nand U4865 (N_4865,N_1671,N_2078);
nand U4866 (N_4866,N_283,N_940);
or U4867 (N_4867,N_2173,N_2441);
nand U4868 (N_4868,N_1585,N_2212);
nand U4869 (N_4869,N_321,N_1707);
nor U4870 (N_4870,N_1801,N_407);
and U4871 (N_4871,N_946,N_1397);
or U4872 (N_4872,N_1169,N_1717);
nand U4873 (N_4873,N_1986,N_1003);
nand U4874 (N_4874,N_1385,N_1977);
nand U4875 (N_4875,N_2285,N_1936);
nand U4876 (N_4876,N_1163,N_788);
nand U4877 (N_4877,N_1674,N_1768);
and U4878 (N_4878,N_1525,N_2258);
nand U4879 (N_4879,N_2430,N_51);
nor U4880 (N_4880,N_1108,N_245);
and U4881 (N_4881,N_1575,N_532);
xor U4882 (N_4882,N_117,N_2284);
nor U4883 (N_4883,N_2297,N_2345);
and U4884 (N_4884,N_653,N_804);
nor U4885 (N_4885,N_197,N_1183);
nand U4886 (N_4886,N_1210,N_280);
nand U4887 (N_4887,N_874,N_974);
and U4888 (N_4888,N_1310,N_2172);
and U4889 (N_4889,N_2309,N_1373);
nand U4890 (N_4890,N_1506,N_135);
nor U4891 (N_4891,N_922,N_1505);
nand U4892 (N_4892,N_1971,N_242);
xnor U4893 (N_4893,N_1672,N_35);
nand U4894 (N_4894,N_1092,N_2451);
nand U4895 (N_4895,N_163,N_1409);
and U4896 (N_4896,N_1131,N_219);
nor U4897 (N_4897,N_1070,N_1661);
nand U4898 (N_4898,N_1129,N_2408);
nand U4899 (N_4899,N_1925,N_739);
nor U4900 (N_4900,N_1274,N_1167);
xor U4901 (N_4901,N_1585,N_1210);
and U4902 (N_4902,N_1120,N_123);
nand U4903 (N_4903,N_2194,N_2293);
nand U4904 (N_4904,N_900,N_256);
and U4905 (N_4905,N_1306,N_1217);
and U4906 (N_4906,N_642,N_343);
nand U4907 (N_4907,N_2076,N_2158);
nand U4908 (N_4908,N_1950,N_2464);
nor U4909 (N_4909,N_2391,N_1991);
nand U4910 (N_4910,N_1429,N_684);
or U4911 (N_4911,N_2066,N_786);
nor U4912 (N_4912,N_980,N_1643);
and U4913 (N_4913,N_672,N_2250);
or U4914 (N_4914,N_833,N_61);
nor U4915 (N_4915,N_596,N_41);
and U4916 (N_4916,N_787,N_212);
or U4917 (N_4917,N_286,N_161);
and U4918 (N_4918,N_1251,N_1849);
or U4919 (N_4919,N_1894,N_1995);
or U4920 (N_4920,N_1554,N_2356);
or U4921 (N_4921,N_167,N_1460);
nand U4922 (N_4922,N_789,N_513);
or U4923 (N_4923,N_2170,N_1566);
and U4924 (N_4924,N_2453,N_2040);
nor U4925 (N_4925,N_828,N_2436);
nor U4926 (N_4926,N_1125,N_1426);
or U4927 (N_4927,N_989,N_1006);
nor U4928 (N_4928,N_98,N_929);
nand U4929 (N_4929,N_1519,N_722);
and U4930 (N_4930,N_1759,N_371);
nand U4931 (N_4931,N_1587,N_2442);
and U4932 (N_4932,N_1593,N_1781);
nor U4933 (N_4933,N_597,N_1230);
nor U4934 (N_4934,N_190,N_1500);
nor U4935 (N_4935,N_933,N_1084);
nor U4936 (N_4936,N_1464,N_2397);
nand U4937 (N_4937,N_1912,N_538);
xnor U4938 (N_4938,N_1312,N_1062);
nor U4939 (N_4939,N_890,N_729);
and U4940 (N_4940,N_2036,N_1818);
xnor U4941 (N_4941,N_2032,N_1260);
nor U4942 (N_4942,N_803,N_136);
and U4943 (N_4943,N_2212,N_236);
or U4944 (N_4944,N_1685,N_897);
xnor U4945 (N_4945,N_2452,N_578);
nand U4946 (N_4946,N_730,N_2162);
xor U4947 (N_4947,N_1808,N_335);
nand U4948 (N_4948,N_1104,N_152);
and U4949 (N_4949,N_1200,N_2049);
nand U4950 (N_4950,N_1591,N_1285);
or U4951 (N_4951,N_2467,N_2438);
or U4952 (N_4952,N_355,N_1179);
and U4953 (N_4953,N_1649,N_366);
and U4954 (N_4954,N_1990,N_1168);
or U4955 (N_4955,N_632,N_1108);
nor U4956 (N_4956,N_1855,N_1942);
or U4957 (N_4957,N_1930,N_939);
nor U4958 (N_4958,N_1432,N_2021);
xor U4959 (N_4959,N_65,N_724);
or U4960 (N_4960,N_309,N_502);
nor U4961 (N_4961,N_1063,N_271);
and U4962 (N_4962,N_1816,N_1544);
and U4963 (N_4963,N_1593,N_788);
nor U4964 (N_4964,N_2005,N_1322);
nand U4965 (N_4965,N_572,N_721);
nand U4966 (N_4966,N_1961,N_1791);
nor U4967 (N_4967,N_1948,N_711);
and U4968 (N_4968,N_1931,N_684);
and U4969 (N_4969,N_729,N_1860);
nor U4970 (N_4970,N_42,N_2143);
nor U4971 (N_4971,N_581,N_70);
and U4972 (N_4972,N_362,N_1466);
nor U4973 (N_4973,N_1667,N_2241);
nor U4974 (N_4974,N_761,N_2078);
nor U4975 (N_4975,N_1123,N_1983);
and U4976 (N_4976,N_2491,N_1447);
and U4977 (N_4977,N_1755,N_1944);
nand U4978 (N_4978,N_2329,N_2116);
nand U4979 (N_4979,N_1862,N_1308);
or U4980 (N_4980,N_2142,N_1365);
or U4981 (N_4981,N_1286,N_1000);
nor U4982 (N_4982,N_1203,N_753);
or U4983 (N_4983,N_1257,N_1951);
nand U4984 (N_4984,N_2182,N_1478);
nor U4985 (N_4985,N_931,N_1872);
nor U4986 (N_4986,N_1208,N_1416);
nor U4987 (N_4987,N_439,N_2060);
nor U4988 (N_4988,N_814,N_517);
nor U4989 (N_4989,N_1632,N_242);
nand U4990 (N_4990,N_801,N_626);
nand U4991 (N_4991,N_1140,N_166);
and U4992 (N_4992,N_1526,N_1645);
and U4993 (N_4993,N_1166,N_628);
nor U4994 (N_4994,N_2471,N_231);
nand U4995 (N_4995,N_1339,N_2169);
nor U4996 (N_4996,N_1111,N_1147);
and U4997 (N_4997,N_869,N_984);
nor U4998 (N_4998,N_1761,N_161);
and U4999 (N_4999,N_1892,N_1757);
nor UO_0 (O_0,N_2900,N_4373);
and UO_1 (O_1,N_4714,N_4868);
nand UO_2 (O_2,N_4399,N_4336);
nor UO_3 (O_3,N_3289,N_4733);
or UO_4 (O_4,N_4993,N_2613);
and UO_5 (O_5,N_4756,N_2644);
nor UO_6 (O_6,N_3404,N_4067);
xor UO_7 (O_7,N_4329,N_2749);
and UO_8 (O_8,N_3217,N_4128);
nand UO_9 (O_9,N_3583,N_3666);
and UO_10 (O_10,N_3905,N_4213);
nand UO_11 (O_11,N_3819,N_3391);
nand UO_12 (O_12,N_4553,N_3985);
and UO_13 (O_13,N_3875,N_3262);
nor UO_14 (O_14,N_4012,N_4279);
and UO_15 (O_15,N_2884,N_3711);
and UO_16 (O_16,N_3786,N_4654);
or UO_17 (O_17,N_4058,N_4609);
nor UO_18 (O_18,N_3453,N_4843);
nand UO_19 (O_19,N_4441,N_2634);
nor UO_20 (O_20,N_2748,N_4800);
or UO_21 (O_21,N_3109,N_3226);
nand UO_22 (O_22,N_4080,N_4754);
or UO_23 (O_23,N_4225,N_2759);
nand UO_24 (O_24,N_4813,N_4939);
or UO_25 (O_25,N_2877,N_2592);
and UO_26 (O_26,N_3771,N_3265);
or UO_27 (O_27,N_3316,N_3270);
nor UO_28 (O_28,N_2807,N_2934);
nand UO_29 (O_29,N_3834,N_2876);
nor UO_30 (O_30,N_4902,N_2706);
nand UO_31 (O_31,N_2908,N_3157);
nand UO_32 (O_32,N_2781,N_4871);
and UO_33 (O_33,N_3148,N_3564);
nand UO_34 (O_34,N_2730,N_2688);
or UO_35 (O_35,N_4896,N_2945);
nor UO_36 (O_36,N_3358,N_2572);
nand UO_37 (O_37,N_4912,N_4405);
and UO_38 (O_38,N_3737,N_3444);
nand UO_39 (O_39,N_4590,N_3049);
and UO_40 (O_40,N_2674,N_3701);
or UO_41 (O_41,N_2528,N_2826);
nand UO_42 (O_42,N_3321,N_3868);
nand UO_43 (O_43,N_3946,N_4883);
or UO_44 (O_44,N_3736,N_4585);
or UO_45 (O_45,N_4735,N_3707);
or UO_46 (O_46,N_3757,N_3740);
and UO_47 (O_47,N_4353,N_4219);
and UO_48 (O_48,N_4243,N_4625);
or UO_49 (O_49,N_4451,N_3896);
nand UO_50 (O_50,N_2673,N_3231);
xnor UO_51 (O_51,N_3703,N_3547);
nor UO_52 (O_52,N_4476,N_4852);
and UO_53 (O_53,N_3980,N_4214);
nor UO_54 (O_54,N_3184,N_4527);
nor UO_55 (O_55,N_4918,N_4270);
and UO_56 (O_56,N_4034,N_4659);
nand UO_57 (O_57,N_2696,N_3100);
nor UO_58 (O_58,N_4528,N_3987);
nor UO_59 (O_59,N_2635,N_3853);
and UO_60 (O_60,N_3253,N_4321);
xor UO_61 (O_61,N_2935,N_4386);
or UO_62 (O_62,N_4537,N_4300);
or UO_63 (O_63,N_3977,N_3445);
or UO_64 (O_64,N_2516,N_4523);
nand UO_65 (O_65,N_4866,N_4463);
or UO_66 (O_66,N_4030,N_4139);
and UO_67 (O_67,N_3017,N_3811);
nor UO_68 (O_68,N_2547,N_4247);
or UO_69 (O_69,N_4589,N_2656);
nor UO_70 (O_70,N_2741,N_3197);
and UO_71 (O_71,N_3576,N_4905);
or UO_72 (O_72,N_4355,N_4357);
nor UO_73 (O_73,N_4119,N_4125);
or UO_74 (O_74,N_4185,N_3561);
nand UO_75 (O_75,N_4269,N_4846);
or UO_76 (O_76,N_4926,N_2624);
nand UO_77 (O_77,N_4556,N_2926);
nor UO_78 (O_78,N_2731,N_4809);
or UO_79 (O_79,N_4639,N_3609);
nand UO_80 (O_80,N_3125,N_3050);
nor UO_81 (O_81,N_4972,N_2575);
nor UO_82 (O_82,N_2586,N_3146);
nand UO_83 (O_83,N_4005,N_3879);
nand UO_84 (O_84,N_4362,N_3407);
nand UO_85 (O_85,N_3187,N_2999);
and UO_86 (O_86,N_2782,N_4383);
nor UO_87 (O_87,N_3618,N_3721);
and UO_88 (O_88,N_3130,N_3694);
nor UO_89 (O_89,N_3411,N_3744);
or UO_90 (O_90,N_2660,N_3511);
and UO_91 (O_91,N_2898,N_3929);
nand UO_92 (O_92,N_2710,N_2846);
nand UO_93 (O_93,N_2973,N_4178);
and UO_94 (O_94,N_2974,N_4326);
nand UO_95 (O_95,N_4867,N_4235);
or UO_96 (O_96,N_4412,N_3945);
nand UO_97 (O_97,N_4211,N_4472);
nand UO_98 (O_98,N_4608,N_4807);
nor UO_99 (O_99,N_3873,N_4471);
or UO_100 (O_100,N_4611,N_3472);
nand UO_101 (O_101,N_4486,N_4909);
nor UO_102 (O_102,N_2518,N_4387);
nand UO_103 (O_103,N_2943,N_4439);
or UO_104 (O_104,N_4285,N_2896);
or UO_105 (O_105,N_3981,N_3635);
or UO_106 (O_106,N_4182,N_4690);
nand UO_107 (O_107,N_3256,N_3091);
nor UO_108 (O_108,N_4582,N_4970);
or UO_109 (O_109,N_4064,N_2694);
or UO_110 (O_110,N_4817,N_4330);
nand UO_111 (O_111,N_3916,N_3084);
nor UO_112 (O_112,N_3405,N_3780);
nor UO_113 (O_113,N_3788,N_4890);
nor UO_114 (O_114,N_4769,N_3622);
nand UO_115 (O_115,N_4892,N_3314);
and UO_116 (O_116,N_2672,N_4007);
nand UO_117 (O_117,N_3881,N_3884);
or UO_118 (O_118,N_4835,N_4586);
and UO_119 (O_119,N_3326,N_4098);
or UO_120 (O_120,N_3438,N_4742);
nand UO_121 (O_121,N_3816,N_3068);
nor UO_122 (O_122,N_3079,N_4886);
nor UO_123 (O_123,N_3441,N_4951);
and UO_124 (O_124,N_2836,N_4145);
or UO_125 (O_125,N_2562,N_4340);
xor UO_126 (O_126,N_4660,N_3186);
nand UO_127 (O_127,N_3007,N_2760);
nand UO_128 (O_128,N_3216,N_4249);
or UO_129 (O_129,N_4447,N_4377);
and UO_130 (O_130,N_4133,N_3515);
nor UO_131 (O_131,N_2500,N_2663);
or UO_132 (O_132,N_4502,N_4927);
or UO_133 (O_133,N_3675,N_4400);
or UO_134 (O_134,N_2863,N_3593);
and UO_135 (O_135,N_4793,N_4144);
nand UO_136 (O_136,N_3335,N_4730);
and UO_137 (O_137,N_4522,N_3702);
nand UO_138 (O_138,N_2918,N_3473);
or UO_139 (O_139,N_4587,N_4333);
nand UO_140 (O_140,N_4117,N_4574);
nor UO_141 (O_141,N_4808,N_2705);
or UO_142 (O_142,N_2995,N_2537);
and UO_143 (O_143,N_3141,N_4198);
and UO_144 (O_144,N_4767,N_4859);
or UO_145 (O_145,N_3241,N_3574);
nand UO_146 (O_146,N_4711,N_3596);
and UO_147 (O_147,N_4567,N_2632);
and UO_148 (O_148,N_4738,N_4017);
nand UO_149 (O_149,N_4202,N_3199);
nor UO_150 (O_150,N_2997,N_4490);
nand UO_151 (O_151,N_3083,N_3932);
and UO_152 (O_152,N_3159,N_4581);
nand UO_153 (O_153,N_4789,N_2699);
or UO_154 (O_154,N_4372,N_4311);
nor UO_155 (O_155,N_3074,N_3155);
nor UO_156 (O_156,N_3949,N_3133);
nor UO_157 (O_157,N_4860,N_2579);
nand UO_158 (O_158,N_4445,N_3023);
nand UO_159 (O_159,N_4264,N_3295);
or UO_160 (O_160,N_2893,N_3910);
nor UO_161 (O_161,N_3591,N_3636);
xor UO_162 (O_162,N_3261,N_4422);
nand UO_163 (O_163,N_3206,N_4550);
or UO_164 (O_164,N_4426,N_3380);
nor UO_165 (O_165,N_4815,N_3024);
nor UO_166 (O_166,N_3132,N_4656);
or UO_167 (O_167,N_3641,N_4197);
nor UO_168 (O_168,N_3501,N_3679);
nor UO_169 (O_169,N_3052,N_3088);
nand UO_170 (O_170,N_3282,N_2789);
and UO_171 (O_171,N_4487,N_3496);
or UO_172 (O_172,N_4915,N_4788);
nor UO_173 (O_173,N_3893,N_4772);
nand UO_174 (O_174,N_4618,N_2690);
nand UO_175 (O_175,N_3890,N_4452);
and UO_176 (O_176,N_3423,N_2859);
and UO_177 (O_177,N_3698,N_3204);
nor UO_178 (O_178,N_4498,N_2866);
and UO_179 (O_179,N_3708,N_2890);
nor UO_180 (O_180,N_4407,N_3785);
and UO_181 (O_181,N_4232,N_4059);
nand UO_182 (O_182,N_3099,N_4947);
nor UO_183 (O_183,N_2954,N_2991);
or UO_184 (O_184,N_2507,N_4127);
nand UO_185 (O_185,N_4072,N_4170);
nor UO_186 (O_186,N_2722,N_4919);
and UO_187 (O_187,N_2679,N_2670);
nor UO_188 (O_188,N_4237,N_4599);
nand UO_189 (O_189,N_2858,N_3251);
nand UO_190 (O_190,N_3730,N_4676);
xnor UO_191 (O_191,N_4680,N_3193);
and UO_192 (O_192,N_2897,N_3723);
or UO_193 (O_193,N_4958,N_2941);
nand UO_194 (O_194,N_3044,N_3754);
and UO_195 (O_195,N_4877,N_3880);
and UO_196 (O_196,N_3720,N_4126);
or UO_197 (O_197,N_3604,N_3934);
and UO_198 (O_198,N_4520,N_4713);
nor UO_199 (O_199,N_3430,N_3060);
or UO_200 (O_200,N_3761,N_2543);
or UO_201 (O_201,N_4338,N_3654);
or UO_202 (O_202,N_3554,N_3953);
or UO_203 (O_203,N_3236,N_4983);
nor UO_204 (O_204,N_2922,N_3891);
and UO_205 (O_205,N_3914,N_4762);
and UO_206 (O_206,N_4151,N_2649);
nand UO_207 (O_207,N_3668,N_2546);
or UO_208 (O_208,N_4819,N_3551);
nor UO_209 (O_209,N_4612,N_2702);
and UO_210 (O_210,N_2519,N_3975);
and UO_211 (O_211,N_4217,N_3971);
nor UO_212 (O_212,N_2755,N_4318);
and UO_213 (O_213,N_2733,N_3863);
and UO_214 (O_214,N_3057,N_4510);
nor UO_215 (O_215,N_2595,N_3960);
nand UO_216 (O_216,N_3436,N_4949);
nor UO_217 (O_217,N_4263,N_3613);
and UO_218 (O_218,N_2622,N_3926);
nor UO_219 (O_219,N_3004,N_4777);
or UO_220 (O_220,N_3807,N_4177);
nor UO_221 (O_221,N_3051,N_3724);
nor UO_222 (O_222,N_4105,N_4932);
and UO_223 (O_223,N_3876,N_3810);
nand UO_224 (O_224,N_3421,N_4507);
nor UO_225 (O_225,N_2530,N_2556);
or UO_226 (O_226,N_3546,N_3093);
or UO_227 (O_227,N_4922,N_4050);
or UO_228 (O_228,N_3240,N_4066);
nand UO_229 (O_229,N_4316,N_3428);
nor UO_230 (O_230,N_3112,N_2647);
nor UO_231 (O_231,N_2697,N_4291);
or UO_232 (O_232,N_3965,N_2923);
or UO_233 (O_233,N_3794,N_3073);
xnor UO_234 (O_234,N_4814,N_3429);
nand UO_235 (O_235,N_4031,N_3513);
nor UO_236 (O_236,N_4552,N_2963);
and UO_237 (O_237,N_4614,N_4049);
nand UO_238 (O_238,N_4544,N_4748);
nor UO_239 (O_239,N_3979,N_3734);
or UO_240 (O_240,N_3791,N_2937);
nor UO_241 (O_241,N_4440,N_3471);
nand UO_242 (O_242,N_4651,N_4454);
nor UO_243 (O_243,N_3566,N_2899);
xor UO_244 (O_244,N_3568,N_3415);
nand UO_245 (O_245,N_4899,N_2541);
and UO_246 (O_246,N_3221,N_4543);
nand UO_247 (O_247,N_4004,N_3018);
nand UO_248 (O_248,N_3454,N_2577);
or UO_249 (O_249,N_3032,N_2578);
and UO_250 (O_250,N_4434,N_4334);
nand UO_251 (O_251,N_4572,N_4238);
nand UO_252 (O_252,N_2982,N_3395);
and UO_253 (O_253,N_2902,N_4262);
nor UO_254 (O_254,N_4500,N_4484);
nor UO_255 (O_255,N_4752,N_3409);
nand UO_256 (O_256,N_2983,N_3128);
nor UO_257 (O_257,N_2667,N_4071);
or UO_258 (O_258,N_3469,N_4429);
nand UO_259 (O_259,N_3812,N_4057);
and UO_260 (O_260,N_3722,N_2992);
nor UO_261 (O_261,N_4204,N_3189);
xnor UO_262 (O_262,N_2910,N_4406);
and UO_263 (O_263,N_4534,N_4018);
nand UO_264 (O_264,N_4136,N_3277);
nor UO_265 (O_265,N_4694,N_4104);
nor UO_266 (O_266,N_3663,N_2676);
nand UO_267 (O_267,N_3346,N_3555);
and UO_268 (O_268,N_4044,N_4479);
or UO_269 (O_269,N_3307,N_3567);
or UO_270 (O_270,N_4090,N_3375);
nor UO_271 (O_271,N_3684,N_2831);
nor UO_272 (O_272,N_3944,N_3648);
and UO_273 (O_273,N_4940,N_4880);
nand UO_274 (O_274,N_3103,N_3237);
and UO_275 (O_275,N_3718,N_4698);
or UO_276 (O_276,N_3478,N_4111);
nor UO_277 (O_277,N_3739,N_3419);
and UO_278 (O_278,N_4875,N_2581);
or UO_279 (O_279,N_4175,N_4816);
nand UO_280 (O_280,N_4266,N_2639);
and UO_281 (O_281,N_3802,N_4041);
xnor UO_282 (O_282,N_4759,N_4753);
nand UO_283 (O_283,N_4848,N_2885);
nand UO_284 (O_284,N_3144,N_3293);
or UO_285 (O_285,N_2604,N_4519);
or UO_286 (O_286,N_3278,N_3385);
and UO_287 (O_287,N_4914,N_2854);
nor UO_288 (O_288,N_4741,N_2571);
nor UO_289 (O_289,N_2681,N_3765);
and UO_290 (O_290,N_3260,N_3210);
nand UO_291 (O_291,N_4118,N_4395);
nand UO_292 (O_292,N_4073,N_3394);
and UO_293 (O_293,N_4369,N_4083);
nand UO_294 (O_294,N_2531,N_3667);
or UO_295 (O_295,N_2612,N_4620);
nand UO_296 (O_296,N_3940,N_4290);
nand UO_297 (O_297,N_3175,N_3520);
or UO_298 (O_298,N_4339,N_3466);
or UO_299 (O_299,N_3121,N_4470);
xnor UO_300 (O_300,N_4900,N_4718);
or UO_301 (O_301,N_2596,N_4576);
or UO_302 (O_302,N_2813,N_3682);
or UO_303 (O_303,N_3259,N_4558);
and UO_304 (O_304,N_3545,N_2906);
nor UO_305 (O_305,N_3176,N_4420);
nor UO_306 (O_306,N_3039,N_4349);
nand UO_307 (O_307,N_3458,N_3340);
nand UO_308 (O_308,N_4980,N_3066);
and UO_309 (O_309,N_3951,N_4776);
and UO_310 (O_310,N_2609,N_4088);
and UO_311 (O_311,N_4293,N_3901);
nor UO_312 (O_312,N_3416,N_3499);
and UO_313 (O_313,N_4649,N_4076);
or UO_314 (O_314,N_4679,N_3205);
and UO_315 (O_315,N_4910,N_2734);
nand UO_316 (O_316,N_2805,N_4925);
or UO_317 (O_317,N_4008,N_3238);
nand UO_318 (O_318,N_4990,N_4248);
nand UO_319 (O_319,N_2882,N_2641);
and UO_320 (O_320,N_3597,N_2559);
or UO_321 (O_321,N_4035,N_3201);
or UO_322 (O_322,N_3572,N_4695);
nor UO_323 (O_323,N_2847,N_3550);
nor UO_324 (O_324,N_2665,N_3578);
nand UO_325 (O_325,N_4906,N_2603);
or UO_326 (O_326,N_4568,N_2685);
nor UO_327 (O_327,N_3291,N_4674);
or UO_328 (O_328,N_3378,N_3163);
or UO_329 (O_329,N_2545,N_3081);
or UO_330 (O_330,N_3072,N_4207);
nor UO_331 (O_331,N_2732,N_3733);
or UO_332 (O_332,N_2631,N_3921);
or UO_333 (O_333,N_2852,N_3273);
and UO_334 (O_334,N_3892,N_4228);
nand UO_335 (O_335,N_2812,N_4021);
nand UO_336 (O_336,N_4302,N_4023);
and UO_337 (O_337,N_3772,N_2867);
and UO_338 (O_338,N_3517,N_4257);
or UO_339 (O_339,N_4856,N_4106);
and UO_340 (O_340,N_4428,N_3271);
nand UO_341 (O_341,N_4070,N_4390);
nor UO_342 (O_342,N_4554,N_3131);
and UO_343 (O_343,N_4536,N_4288);
nand UO_344 (O_344,N_3285,N_3016);
or UO_345 (O_345,N_3065,N_4295);
and UO_346 (O_346,N_2560,N_3500);
and UO_347 (O_347,N_3955,N_3681);
nand UO_348 (O_348,N_2557,N_4312);
nor UO_349 (O_349,N_3653,N_4965);
nor UO_350 (O_350,N_4715,N_2588);
nor UO_351 (O_351,N_3821,N_3913);
or UO_352 (O_352,N_2662,N_4220);
and UO_353 (O_353,N_4954,N_4758);
or UO_354 (O_354,N_3098,N_2591);
or UO_355 (O_355,N_4414,N_3882);
nor UO_356 (O_356,N_3571,N_4162);
and UO_357 (O_357,N_2753,N_3180);
and UO_358 (O_358,N_4193,N_3686);
nand UO_359 (O_359,N_4529,N_2980);
xnor UO_360 (O_360,N_2558,N_4466);
nand UO_361 (O_361,N_2853,N_4408);
and UO_362 (O_362,N_2872,N_2953);
nor UO_363 (O_363,N_3457,N_4063);
or UO_364 (O_364,N_2529,N_4839);
and UO_365 (O_365,N_4449,N_3958);
or UO_366 (O_366,N_3283,N_3448);
nand UO_367 (O_367,N_4596,N_4169);
and UO_368 (O_368,N_4891,N_3961);
nand UO_369 (O_369,N_3587,N_2677);
nand UO_370 (O_370,N_4184,N_3580);
and UO_371 (O_371,N_2593,N_4666);
nor UO_372 (O_372,N_2565,N_4770);
and UO_373 (O_373,N_4524,N_3645);
or UO_374 (O_374,N_3915,N_4124);
nand UO_375 (O_375,N_3337,N_3610);
nor UO_376 (O_376,N_3954,N_2648);
and UO_377 (O_377,N_4465,N_2790);
nor UO_378 (O_378,N_3598,N_4040);
and UO_379 (O_379,N_3617,N_4354);
nor UO_380 (O_380,N_4650,N_4483);
nor UO_381 (O_381,N_3713,N_3117);
nand UO_382 (O_382,N_3652,N_4917);
and UO_383 (O_383,N_4240,N_2608);
or UO_384 (O_384,N_3775,N_4564);
nor UO_385 (O_385,N_4097,N_3067);
nor UO_386 (O_386,N_4029,N_2640);
and UO_387 (O_387,N_2520,N_3918);
nor UO_388 (O_388,N_3728,N_2598);
or UO_389 (O_389,N_4233,N_2633);
and UO_390 (O_390,N_3410,N_4280);
and UO_391 (O_391,N_4468,N_3615);
or UO_392 (O_392,N_3185,N_3994);
nand UO_393 (O_393,N_4367,N_3966);
or UO_394 (O_394,N_3877,N_2600);
or UO_395 (O_395,N_3590,N_4560);
and UO_396 (O_396,N_4881,N_3178);
nand UO_397 (O_397,N_3705,N_4950);
nand UO_398 (O_398,N_2797,N_4047);
nand UO_399 (O_399,N_4706,N_2567);
nand UO_400 (O_400,N_3214,N_3753);
nand UO_401 (O_401,N_2940,N_3862);
nand UO_402 (O_402,N_4619,N_3297);
nor UO_403 (O_403,N_4768,N_3383);
nor UO_404 (O_404,N_3027,N_3181);
nand UO_405 (O_405,N_3420,N_3026);
and UO_406 (O_406,N_2879,N_3227);
nand UO_407 (O_407,N_4398,N_3938);
nor UO_408 (O_408,N_4026,N_3699);
and UO_409 (O_409,N_3059,N_2810);
nor UO_410 (O_410,N_4923,N_4684);
and UO_411 (O_411,N_2947,N_3855);
or UO_412 (O_412,N_4056,N_2564);
nor UO_413 (O_413,N_4164,N_3367);
nor UO_414 (O_414,N_2566,N_4132);
and UO_415 (O_415,N_4389,N_2944);
and UO_416 (O_416,N_4165,N_4485);
nand UO_417 (O_417,N_2580,N_2764);
or UO_418 (O_418,N_3817,N_4190);
and UO_419 (O_419,N_3127,N_3563);
nor UO_420 (O_420,N_2659,N_4999);
and UO_421 (O_421,N_3743,N_4976);
or UO_422 (O_422,N_4039,N_3446);
and UO_423 (O_423,N_2961,N_4131);
nor UO_424 (O_424,N_3333,N_3245);
and UO_425 (O_425,N_3984,N_3219);
and UO_426 (O_426,N_3532,N_3138);
nand UO_427 (O_427,N_4323,N_3840);
or UO_428 (O_428,N_4024,N_2772);
nand UO_429 (O_429,N_4982,N_2534);
nand UO_430 (O_430,N_2642,N_4584);
and UO_431 (O_431,N_4045,N_2505);
nor UO_432 (O_432,N_4559,N_2763);
and UO_433 (O_433,N_2783,N_4862);
and UO_434 (O_434,N_4351,N_2855);
nor UO_435 (O_435,N_2501,N_4729);
nand UO_436 (O_436,N_3778,N_4149);
or UO_437 (O_437,N_2637,N_2978);
nor UO_438 (O_438,N_3726,N_2971);
nand UO_439 (O_439,N_4179,N_4531);
nand UO_440 (O_440,N_3368,N_4653);
or UO_441 (O_441,N_4301,N_4123);
and UO_442 (O_442,N_4419,N_4824);
nand UO_443 (O_443,N_2620,N_2803);
nand UO_444 (O_444,N_4037,N_3776);
and UO_445 (O_445,N_3838,N_4703);
nor UO_446 (O_446,N_4600,N_2800);
nor UO_447 (O_447,N_4436,N_2870);
and UO_448 (O_448,N_3745,N_4423);
or UO_449 (O_449,N_4987,N_2939);
or UO_450 (O_450,N_3406,N_3630);
and UO_451 (O_451,N_2862,N_4109);
and UO_452 (O_452,N_4089,N_4348);
or UO_453 (O_453,N_3303,N_2989);
or UO_454 (O_454,N_4404,N_3519);
nor UO_455 (O_455,N_4462,N_3382);
or UO_456 (O_456,N_4110,N_2771);
nand UO_457 (O_457,N_2747,N_2832);
nor UO_458 (O_458,N_4798,N_3494);
and UO_459 (O_459,N_3126,N_2841);
nor UO_460 (O_460,N_3047,N_3996);
nand UO_461 (O_461,N_3600,N_2616);
nand UO_462 (O_462,N_3090,N_3431);
and UO_463 (O_463,N_3789,N_2960);
nor UO_464 (O_464,N_3837,N_4646);
nand UO_465 (O_465,N_3043,N_3165);
and UO_466 (O_466,N_4697,N_3113);
nand UO_467 (O_467,N_3467,N_3055);
nor UO_468 (O_468,N_2720,N_4624);
xnor UO_469 (O_469,N_4314,N_2684);
nand UO_470 (O_470,N_4781,N_2550);
and UO_471 (O_471,N_3010,N_4744);
or UO_472 (O_472,N_2745,N_4884);
or UO_473 (O_473,N_3276,N_4731);
nand UO_474 (O_474,N_4061,N_3755);
and UO_475 (O_475,N_3006,N_3491);
nand UO_476 (O_476,N_3797,N_4092);
and UO_477 (O_477,N_3925,N_4096);
nor UO_478 (O_478,N_2652,N_2904);
nor UO_479 (O_479,N_3056,N_4944);
nand UO_480 (O_480,N_3859,N_3234);
nand UO_481 (O_481,N_3069,N_3443);
or UO_482 (O_482,N_4384,N_2845);
nand UO_483 (O_483,N_4378,N_3371);
and UO_484 (O_484,N_3168,N_3485);
or UO_485 (O_485,N_3941,N_4019);
and UO_486 (O_486,N_3468,N_4913);
nand UO_487 (O_487,N_2668,N_2606);
and UO_488 (O_488,N_2919,N_3486);
or UO_489 (O_489,N_4229,N_3369);
nand UO_490 (O_490,N_3582,N_4491);
or UO_491 (O_491,N_4226,N_3871);
or UO_492 (O_492,N_3783,N_4864);
nor UO_493 (O_493,N_3095,N_3338);
nor UO_494 (O_494,N_4172,N_4167);
nand UO_495 (O_495,N_3830,N_3748);
xor UO_496 (O_496,N_3841,N_3957);
and UO_497 (O_497,N_4274,N_4791);
nand UO_498 (O_498,N_4747,N_4048);
and UO_499 (O_499,N_3076,N_4885);
nand UO_500 (O_500,N_3606,N_3455);
xor UO_501 (O_501,N_3858,N_4086);
nand UO_502 (O_502,N_4432,N_3620);
nor UO_503 (O_503,N_4481,N_3320);
nand UO_504 (O_504,N_4736,N_4402);
and UO_505 (O_505,N_4806,N_3809);
and UO_506 (O_506,N_3235,N_3200);
nand UO_507 (O_507,N_4025,N_2726);
and UO_508 (O_508,N_2975,N_3451);
and UO_509 (O_509,N_3601,N_2820);
nor UO_510 (O_510,N_4299,N_3599);
or UO_511 (O_511,N_4566,N_4227);
and UO_512 (O_512,N_3939,N_4577);
nand UO_513 (O_513,N_2988,N_4397);
or UO_514 (O_514,N_4532,N_3147);
nor UO_515 (O_515,N_3612,N_3061);
and UO_516 (O_516,N_4540,N_2617);
xnor UO_517 (O_517,N_3403,N_3505);
and UO_518 (O_518,N_3104,N_4681);
or UO_519 (O_519,N_2587,N_3250);
nand UO_520 (O_520,N_2822,N_3120);
and UO_521 (O_521,N_4701,N_3509);
nor UO_522 (O_522,N_4805,N_4187);
or UO_523 (O_523,N_4606,N_2686);
nor UO_524 (O_524,N_4003,N_2654);
nor UO_525 (O_525,N_4006,N_4894);
nor UO_526 (O_526,N_3424,N_3693);
nand UO_527 (O_527,N_2682,N_2522);
or UO_528 (O_528,N_4916,N_3264);
and UO_529 (O_529,N_4746,N_3878);
or UO_530 (O_530,N_4459,N_4036);
or UO_531 (O_531,N_3012,N_3845);
or UO_532 (O_532,N_2875,N_4750);
or UO_533 (O_533,N_4464,N_2860);
nor UO_534 (O_534,N_3341,N_4331);
nor UO_535 (O_535,N_3030,N_3650);
or UO_536 (O_536,N_4723,N_3412);
nand UO_537 (O_537,N_3548,N_4020);
or UO_538 (O_538,N_3209,N_3479);
nor UO_539 (O_539,N_4928,N_4166);
nand UO_540 (O_540,N_3498,N_4513);
or UO_541 (O_541,N_3427,N_4936);
nor UO_542 (O_542,N_4276,N_4903);
and UO_543 (O_543,N_4212,N_4103);
nand UO_544 (O_544,N_3631,N_2986);
and UO_545 (O_545,N_3602,N_4218);
xnor UO_546 (O_546,N_4953,N_2707);
nand UO_547 (O_547,N_4783,N_4765);
and UO_548 (O_548,N_3792,N_3171);
and UO_549 (O_549,N_3639,N_4091);
nor UO_550 (O_550,N_4642,N_4861);
or UO_551 (O_551,N_3632,N_3844);
or UO_552 (O_552,N_3621,N_4810);
nor UO_553 (O_553,N_2661,N_3167);
or UO_554 (O_554,N_4959,N_4284);
or UO_555 (O_555,N_3220,N_3134);
or UO_556 (O_556,N_4766,N_4563);
and UO_557 (O_557,N_2651,N_3142);
nor UO_558 (O_558,N_4787,N_3452);
nand UO_559 (O_559,N_2931,N_2767);
xnor UO_560 (O_560,N_3366,N_3527);
nor UO_561 (O_561,N_2938,N_4113);
xnor UO_562 (O_562,N_3784,N_3137);
and UO_563 (O_563,N_4937,N_2990);
or UO_564 (O_564,N_3174,N_3249);
nand UO_565 (O_565,N_4493,N_4231);
nand UO_566 (O_566,N_2643,N_2936);
nand UO_567 (O_567,N_3396,N_4492);
nor UO_568 (O_568,N_4597,N_3274);
nand UO_569 (O_569,N_2514,N_2757);
or UO_570 (O_570,N_4998,N_3474);
nand UO_571 (O_571,N_4009,N_3425);
nand UO_572 (O_572,N_2542,N_4641);
nand UO_573 (O_573,N_3738,N_2787);
and UO_574 (O_574,N_3674,N_3480);
nand UO_575 (O_575,N_4273,N_3450);
xnor UO_576 (O_576,N_2880,N_2738);
and UO_577 (O_577,N_3046,N_3160);
nand UO_578 (O_578,N_2804,N_4975);
nor UO_579 (O_579,N_4836,N_3968);
and UO_580 (O_580,N_3002,N_3646);
nand UO_581 (O_581,N_3284,N_4647);
nor UO_582 (O_582,N_3592,N_3731);
nor UO_583 (O_583,N_3244,N_3909);
or UO_584 (O_584,N_3456,N_3263);
and UO_585 (O_585,N_2928,N_3541);
xor UO_586 (O_586,N_4392,N_4289);
and UO_587 (O_587,N_3339,N_3689);
nor UO_588 (O_588,N_3194,N_3332);
or UO_589 (O_589,N_2808,N_2658);
nand UO_590 (O_590,N_4194,N_3370);
nor UO_591 (O_591,N_3584,N_4851);
nand UO_592 (O_592,N_2555,N_2964);
and UO_593 (O_593,N_2843,N_4627);
and UO_594 (O_594,N_4246,N_3865);
or UO_595 (O_595,N_4033,N_2766);
nand UO_596 (O_596,N_2628,N_2746);
or UO_597 (O_597,N_4356,N_4538);
nor UO_598 (O_598,N_2619,N_3773);
and UO_599 (O_599,N_3933,N_4192);
xor UO_600 (O_600,N_2815,N_3922);
nor UO_601 (O_601,N_4632,N_3000);
or UO_602 (O_602,N_2725,N_3161);
or UO_603 (O_603,N_2574,N_4394);
and UO_604 (O_604,N_3993,N_3508);
nor UO_605 (O_605,N_2589,N_3714);
and UO_606 (O_606,N_3033,N_2967);
or UO_607 (O_607,N_4850,N_4253);
nor UO_608 (O_608,N_3956,N_4359);
xor UO_609 (O_609,N_3856,N_4841);
nand UO_610 (O_610,N_3037,N_3661);
or UO_611 (O_611,N_4996,N_3796);
and UO_612 (O_612,N_4241,N_4603);
or UO_613 (O_613,N_3135,N_4545);
nand UO_614 (O_614,N_3512,N_2743);
nor UO_615 (O_615,N_4709,N_4409);
nor UO_616 (O_616,N_4475,N_4271);
nor UO_617 (O_617,N_3687,N_3577);
and UO_618 (O_618,N_3062,N_4995);
or UO_619 (O_619,N_3224,N_2709);
nand UO_620 (O_620,N_4173,N_3317);
or UO_621 (O_621,N_2946,N_4046);
nor UO_622 (O_622,N_4548,N_4203);
nor UO_623 (O_623,N_4988,N_4623);
nand UO_624 (O_624,N_4478,N_2915);
or UO_625 (O_625,N_3475,N_3696);
or UO_626 (O_626,N_3762,N_2834);
or UO_627 (O_627,N_4561,N_3553);
and UO_628 (O_628,N_4751,N_2942);
or UO_629 (O_629,N_3348,N_3746);
and UO_630 (O_630,N_3963,N_2785);
and UO_631 (O_631,N_2513,N_3857);
and UO_632 (O_632,N_4107,N_3233);
and UO_633 (O_633,N_4551,N_3034);
nor UO_634 (O_634,N_4503,N_4863);
or UO_635 (O_635,N_2985,N_4508);
and UO_636 (O_636,N_4557,N_2675);
or UO_637 (O_637,N_3272,N_2788);
nand UO_638 (O_638,N_3823,N_2993);
and UO_639 (O_639,N_4474,N_2930);
or UO_640 (O_640,N_4032,N_4967);
xnor UO_641 (O_641,N_2511,N_4208);
and UO_642 (O_642,N_4148,N_3154);
nor UO_643 (O_643,N_2828,N_3437);
or UO_644 (O_644,N_3070,N_4437);
or UO_645 (O_645,N_3015,N_3439);
nand UO_646 (O_646,N_2768,N_2765);
or UO_647 (O_647,N_4306,N_2761);
and UO_648 (O_648,N_2903,N_2887);
nor UO_649 (O_649,N_3729,N_3392);
or UO_650 (O_650,N_4616,N_2977);
and UO_651 (O_651,N_4446,N_4638);
nor UO_652 (O_652,N_2869,N_4604);
or UO_653 (O_653,N_3673,N_4014);
nor UO_654 (O_654,N_2840,N_4968);
nand UO_655 (O_655,N_3183,N_2950);
or UO_656 (O_656,N_3350,N_3038);
nand UO_657 (O_657,N_3695,N_3470);
nor UO_658 (O_658,N_2729,N_4308);
and UO_659 (O_659,N_3414,N_4921);
nand UO_660 (O_660,N_4870,N_4633);
nand UO_661 (O_661,N_4686,N_3942);
nand UO_662 (O_662,N_3334,N_4418);
or UO_663 (O_663,N_4542,N_4027);
and UO_664 (O_664,N_4942,N_3533);
nor UO_665 (O_665,N_3182,N_4275);
or UO_666 (O_666,N_3831,N_3920);
and UO_667 (O_667,N_3384,N_2750);
or UO_668 (O_668,N_2535,N_4898);
nor UO_669 (O_669,N_4844,N_3657);
nand UO_670 (O_670,N_2721,N_3935);
and UO_671 (O_671,N_4458,N_4347);
and UO_672 (O_672,N_4011,N_3995);
and UO_673 (O_673,N_3895,N_3054);
nand UO_674 (O_674,N_4931,N_3904);
nor UO_675 (O_675,N_4438,N_3637);
nor UO_676 (O_676,N_4602,N_2965);
nor UO_677 (O_677,N_3751,N_4533);
nor UO_678 (O_678,N_3166,N_3153);
or UO_679 (O_679,N_4413,N_3053);
or UO_680 (O_680,N_4114,N_4685);
and UO_681 (O_681,N_3361,N_3526);
nor UO_682 (O_682,N_3638,N_3886);
or UO_683 (O_683,N_4210,N_3634);
and UO_684 (O_684,N_3725,N_4645);
and UO_685 (O_685,N_4401,N_3849);
or UO_686 (O_686,N_3805,N_3124);
and UO_687 (O_687,N_2680,N_4622);
or UO_688 (O_688,N_4343,N_3188);
or UO_689 (O_689,N_2864,N_2933);
nor UO_690 (O_690,N_2856,N_3864);
or UO_691 (O_691,N_4042,N_4161);
or UO_692 (O_692,N_2532,N_3575);
and UO_693 (O_693,N_3110,N_3774);
nor UO_694 (O_694,N_2792,N_4963);
nand UO_695 (O_695,N_3286,N_3462);
nor UO_696 (O_696,N_3839,N_4457);
or UO_697 (O_697,N_4727,N_2703);
or UO_698 (O_698,N_4448,N_3874);
nand UO_699 (O_699,N_2568,N_2913);
or UO_700 (O_700,N_3354,N_3662);
nor UO_701 (O_701,N_4078,N_3432);
or UO_702 (O_702,N_3389,N_2957);
nor UO_703 (O_703,N_3507,N_4887);
and UO_704 (O_704,N_2655,N_2824);
or UO_705 (O_705,N_4827,N_4637);
nor UO_706 (O_706,N_3815,N_2894);
xor UO_707 (O_707,N_3353,N_3021);
or UO_708 (O_708,N_4473,N_3042);
nand UO_709 (O_709,N_4176,N_4297);
nor UO_710 (O_710,N_4075,N_4802);
and UO_711 (O_711,N_4601,N_3490);
and UO_712 (O_712,N_2958,N_3118);
and UO_713 (O_713,N_4251,N_2976);
nor UO_714 (O_714,N_2968,N_4693);
nor UO_715 (O_715,N_3825,N_4224);
nand UO_716 (O_716,N_4317,N_3268);
nand UO_717 (O_717,N_3531,N_4853);
or UO_718 (O_718,N_2994,N_3543);
nand UO_719 (O_719,N_4876,N_3097);
or UO_720 (O_720,N_3628,N_4665);
and UO_721 (O_721,N_3770,N_2544);
or UO_722 (O_722,N_3082,N_3521);
nand UO_723 (O_723,N_3179,N_4661);
nand UO_724 (O_724,N_3659,N_4244);
nor UO_725 (O_725,N_4872,N_3319);
nand UO_726 (O_726,N_2523,N_3362);
and UO_727 (O_727,N_3247,N_4525);
or UO_728 (O_728,N_4874,N_4153);
or UO_729 (O_729,N_2776,N_3211);
nor UO_730 (O_730,N_2517,N_2929);
and UO_731 (O_731,N_3022,N_3801);
and UO_732 (O_732,N_2552,N_3246);
or UO_733 (O_733,N_3676,N_4252);
nor UO_734 (O_734,N_4992,N_3542);
nand UO_735 (O_735,N_2736,N_4668);
nor UO_736 (O_736,N_4823,N_2585);
nand UO_737 (O_737,N_2818,N_4068);
nand UO_738 (O_738,N_4477,N_3860);
nor UO_739 (O_739,N_4150,N_3324);
nand UO_740 (O_740,N_3014,N_4652);
or UO_741 (O_741,N_4450,N_2878);
or UO_742 (O_742,N_4530,N_4135);
or UO_743 (O_743,N_2901,N_2959);
nand UO_744 (O_744,N_3417,N_3312);
nand UO_745 (O_745,N_3923,N_4617);
or UO_746 (O_746,N_3642,N_3013);
nand UO_747 (O_747,N_3767,N_3029);
and UO_748 (O_748,N_2786,N_2780);
nand UO_749 (O_749,N_4794,N_4268);
or UO_750 (O_750,N_4811,N_3752);
nor UO_751 (O_751,N_4778,N_4382);
and UO_752 (O_752,N_4515,N_4427);
or UO_753 (O_753,N_4122,N_2539);
or UO_754 (O_754,N_4740,N_3356);
nor UO_755 (O_755,N_3536,N_3677);
or UO_756 (O_756,N_3558,N_2524);
nand UO_757 (O_757,N_2842,N_4570);
and UO_758 (O_758,N_2891,N_3894);
or UO_759 (O_759,N_4761,N_4829);
or UO_760 (O_760,N_3198,N_2793);
nor UO_761 (O_761,N_4368,N_3357);
and UO_762 (O_762,N_4315,N_4380);
or UO_763 (O_763,N_2506,N_4174);
or UO_764 (O_764,N_3594,N_3433);
and UO_765 (O_765,N_3465,N_3978);
nand UO_766 (O_766,N_4716,N_3342);
nor UO_767 (O_767,N_4705,N_3483);
and UO_768 (O_768,N_2952,N_4857);
xnor UO_769 (O_769,N_4728,N_2512);
or UO_770 (O_770,N_3660,N_4845);
nand UO_771 (O_771,N_4726,N_3190);
nand UO_772 (O_772,N_4734,N_4820);
xnor UO_773 (O_773,N_3899,N_3345);
and UO_774 (O_774,N_4381,N_4797);
and UO_775 (O_775,N_4102,N_2849);
and UO_776 (O_776,N_3769,N_4689);
or UO_777 (O_777,N_4155,N_4688);
nand UO_778 (O_778,N_2583,N_4365);
or UO_779 (O_779,N_4010,N_4675);
or UO_780 (O_780,N_2540,N_3257);
nor UO_781 (O_781,N_3900,N_2692);
or UO_782 (O_782,N_3931,N_3742);
nor UO_783 (O_783,N_4774,N_2723);
or UO_784 (O_784,N_2503,N_4888);
and UO_785 (O_785,N_4721,N_4549);
nand UO_786 (O_786,N_4546,N_3058);
nor UO_787 (O_787,N_3808,N_4722);
and UO_788 (O_788,N_4496,N_4022);
and UO_789 (O_789,N_3967,N_4779);
nor UO_790 (O_790,N_4957,N_3795);
or UO_791 (O_791,N_3588,N_2932);
nand UO_792 (O_792,N_4948,N_2981);
and UO_793 (O_793,N_2701,N_3390);
and UO_794 (O_794,N_4640,N_4101);
nand UO_795 (O_795,N_4635,N_3524);
or UO_796 (O_796,N_3492,N_2739);
or UO_797 (O_797,N_2802,N_4431);
nor UO_798 (O_798,N_3804,N_4952);
or UO_799 (O_799,N_2754,N_4929);
nor UO_800 (O_800,N_3998,N_3623);
or UO_801 (O_801,N_4388,N_4001);
nand UO_802 (O_802,N_4760,N_4456);
nor UO_803 (O_803,N_4051,N_3299);
and UO_804 (O_804,N_2623,N_3075);
nor UO_805 (O_805,N_2969,N_3484);
nor UO_806 (O_806,N_3413,N_4840);
or UO_807 (O_807,N_4828,N_3685);
and UO_808 (O_808,N_3009,N_4286);
and UO_809 (O_809,N_4821,N_3888);
nor UO_810 (O_810,N_3902,N_4555);
or UO_811 (O_811,N_3242,N_4956);
nor UO_812 (O_812,N_4296,N_3537);
nor UO_813 (O_813,N_4112,N_3172);
and UO_814 (O_814,N_4256,N_4499);
or UO_815 (O_815,N_4396,N_3992);
nor UO_816 (O_816,N_3169,N_2715);
nor UO_817 (O_817,N_4313,N_3683);
nor UO_818 (O_818,N_4489,N_4605);
nor UO_819 (O_819,N_4209,N_4303);
nor UO_820 (O_820,N_3349,N_4421);
nand UO_821 (O_821,N_2650,N_4245);
or UO_822 (O_822,N_4573,N_4518);
nand UO_823 (O_823,N_2599,N_2751);
nor UO_824 (O_824,N_3664,N_4541);
nor UO_825 (O_825,N_4655,N_4964);
and UO_826 (O_826,N_3288,N_3028);
nand UO_827 (O_827,N_4505,N_4168);
or UO_828 (O_828,N_2740,N_2886);
nor UO_829 (O_829,N_3861,N_4708);
or UO_830 (O_830,N_2924,N_3077);
or UO_831 (O_831,N_4038,N_4644);
and UO_832 (O_832,N_4028,N_2752);
nand UO_833 (O_833,N_3301,N_3822);
or UO_834 (O_834,N_4696,N_4662);
nor UO_835 (O_835,N_3177,N_3482);
or UO_836 (O_836,N_3309,N_2799);
and UO_837 (O_837,N_4785,N_3690);
nor UO_838 (O_838,N_3866,N_4361);
nand UO_839 (O_839,N_2778,N_2774);
nor UO_840 (O_840,N_3712,N_3426);
and UO_841 (O_841,N_4278,N_2521);
and UO_842 (O_842,N_2570,N_3158);
nand UO_843 (O_843,N_2920,N_4565);
and UO_844 (O_844,N_2735,N_2829);
nand UO_845 (O_845,N_3078,N_3464);
or UO_846 (O_846,N_2573,N_2851);
nand UO_847 (O_847,N_4771,N_3885);
or UO_848 (O_848,N_4158,N_3108);
nand UO_849 (O_849,N_4410,N_4310);
nor UO_850 (O_850,N_4115,N_3330);
or UO_851 (O_851,N_3195,N_2956);
nor UO_852 (O_852,N_3846,N_3854);
nand UO_853 (O_853,N_4636,N_4935);
nor UO_854 (O_854,N_3372,N_4223);
or UO_855 (O_855,N_4960,N_3281);
nand UO_856 (O_856,N_4615,N_3827);
nand UO_857 (O_857,N_3308,N_4142);
nor UO_858 (O_858,N_2683,N_4480);
nor UO_859 (O_859,N_3140,N_4725);
and UO_860 (O_860,N_4580,N_2724);
and UO_861 (O_861,N_4773,N_4658);
and UO_862 (O_862,N_2850,N_3710);
and UO_863 (O_863,N_3525,N_3031);
and UO_864 (O_864,N_3624,N_3990);
nand UO_865 (O_865,N_4495,N_4234);
or UO_866 (O_866,N_4328,N_4055);
or UO_867 (O_867,N_4930,N_4717);
nand UO_868 (O_868,N_3045,N_2618);
xnor UO_869 (O_869,N_4200,N_4943);
or UO_870 (O_870,N_4962,N_3287);
nand UO_871 (O_871,N_4855,N_3756);
nor UO_872 (O_872,N_4745,N_3565);
or UO_873 (O_873,N_3930,N_4629);
nand UO_874 (O_874,N_3749,N_4385);
and UO_875 (O_875,N_3820,N_3972);
or UO_876 (O_876,N_3988,N_3212);
nand UO_877 (O_877,N_3847,N_4298);
and UO_878 (O_878,N_3115,N_3379);
or UO_879 (O_879,N_2811,N_3089);
or UO_880 (O_880,N_4934,N_2814);
nand UO_881 (O_881,N_2614,N_3143);
nand UO_882 (O_882,N_4672,N_4782);
nand UO_883 (O_883,N_3672,N_3556);
nand UO_884 (O_884,N_2744,N_3228);
nor UO_885 (O_885,N_3897,N_3540);
and UO_886 (O_886,N_4265,N_4834);
nand UO_887 (O_887,N_3196,N_3586);
and UO_888 (O_888,N_4907,N_2871);
nor UO_889 (O_889,N_4707,N_2984);
nor UO_890 (O_890,N_4621,N_2949);
and UO_891 (O_891,N_3222,N_3611);
and UO_892 (O_892,N_3156,N_3658);
nand UO_893 (O_893,N_4236,N_3048);
nand UO_894 (O_894,N_3311,N_3020);
nor UO_895 (O_895,N_4335,N_4364);
or UO_896 (O_896,N_3487,N_3493);
nor UO_897 (O_897,N_3254,N_3323);
nand UO_898 (O_898,N_2708,N_4043);
and UO_899 (O_899,N_3560,N_4626);
or UO_900 (O_900,N_3782,N_4282);
or UO_901 (O_901,N_2881,N_2835);
or UO_902 (O_902,N_3917,N_4054);
or UO_903 (O_903,N_3164,N_3947);
or UO_904 (O_904,N_2526,N_2911);
or UO_905 (O_905,N_4796,N_3459);
and UO_906 (O_906,N_4065,N_3616);
nor UO_907 (O_907,N_3626,N_3399);
xor UO_908 (O_908,N_3603,N_3129);
nor UO_909 (O_909,N_2883,N_4363);
nand UO_910 (O_910,N_3481,N_4562);
nor UO_911 (O_911,N_4994,N_4391);
nor UO_912 (O_912,N_4157,N_4242);
or UO_913 (O_913,N_3398,N_4547);
nor UO_914 (O_914,N_3397,N_3387);
nand UO_915 (O_915,N_4239,N_4254);
or UO_916 (O_916,N_2727,N_3928);
nor UO_917 (O_917,N_3119,N_2590);
and UO_918 (O_918,N_3400,N_3529);
or UO_919 (O_919,N_3085,N_3041);
or UO_920 (O_920,N_3758,N_3997);
or UO_921 (O_921,N_3300,N_3950);
or UO_922 (O_922,N_2823,N_4453);
or UO_923 (O_923,N_3570,N_4191);
and UO_924 (O_924,N_4663,N_3306);
and UO_925 (O_925,N_3735,N_3843);
nor UO_926 (O_926,N_3814,N_4795);
nor UO_927 (O_927,N_4578,N_2627);
nand UO_928 (O_928,N_4878,N_3080);
and UO_929 (O_929,N_4780,N_4425);
or UO_930 (O_930,N_4961,N_2597);
nor UO_931 (O_931,N_4325,N_3700);
or UO_932 (O_932,N_3489,N_3852);
nor UO_933 (O_933,N_2914,N_4152);
or UO_934 (O_934,N_3418,N_4469);
nor UO_935 (O_935,N_4764,N_2666);
and UO_936 (O_936,N_2636,N_3552);
nor UO_937 (O_937,N_2561,N_4222);
nand UO_938 (O_938,N_4691,N_4435);
or UO_939 (O_939,N_4989,N_3535);
or UO_940 (O_940,N_2638,N_4517);
and UO_941 (O_941,N_3136,N_3803);
and UO_942 (O_942,N_3401,N_4804);
nor UO_943 (O_943,N_2695,N_4206);
and UO_944 (O_944,N_4984,N_2833);
or UO_945 (O_945,N_3087,N_2717);
nand UO_946 (O_946,N_3627,N_3614);
nor UO_947 (O_947,N_3549,N_4920);
or UO_948 (O_948,N_3294,N_2584);
nor UO_949 (O_949,N_4433,N_4830);
nand UO_950 (O_950,N_3619,N_4403);
nand UO_951 (O_951,N_3640,N_3280);
nor UO_952 (O_952,N_3647,N_4924);
nand UO_953 (O_953,N_2987,N_4013);
and UO_954 (O_954,N_3826,N_4739);
nand UO_955 (O_955,N_4100,N_4230);
xnor UO_956 (O_956,N_3760,N_3651);
or UO_957 (O_957,N_3497,N_3559);
or UO_958 (O_958,N_4593,N_4732);
nand UO_959 (O_959,N_3304,N_3510);
nand UO_960 (O_960,N_3633,N_4648);
nor UO_961 (O_961,N_4799,N_4221);
nor UO_962 (O_962,N_2874,N_3538);
or UO_963 (O_963,N_4307,N_4973);
nand UO_964 (O_964,N_3011,N_2777);
or UO_965 (O_965,N_4467,N_4358);
xnor UO_966 (O_966,N_3629,N_2796);
nand UO_967 (O_967,N_2607,N_3275);
nor UO_968 (O_968,N_4667,N_3377);
nand UO_969 (O_969,N_4539,N_3557);
nand UO_970 (O_970,N_4375,N_2798);
nor UO_971 (O_971,N_4579,N_3927);
or UO_972 (O_972,N_4120,N_3716);
or UO_973 (O_973,N_2646,N_3906);
nor UO_974 (O_974,N_3035,N_3116);
nand UO_975 (O_975,N_2848,N_3697);
nor UO_976 (O_976,N_3460,N_4749);
nor UO_977 (O_977,N_3991,N_4933);
xnor UO_978 (O_978,N_4077,N_4613);
or UO_979 (O_979,N_2873,N_3463);
or UO_980 (O_980,N_2955,N_2827);
xor UO_981 (O_981,N_3842,N_3248);
or UO_982 (O_982,N_4743,N_4319);
nand UO_983 (O_983,N_3229,N_4673);
or UO_984 (O_984,N_3279,N_4074);
nor UO_985 (O_985,N_3781,N_3655);
and UO_986 (O_986,N_4801,N_4015);
or UO_987 (O_987,N_2770,N_4188);
or UO_988 (O_988,N_3374,N_4140);
nand UO_989 (O_989,N_4199,N_3503);
or UO_990 (O_990,N_3213,N_4833);
nor UO_991 (O_991,N_3656,N_4171);
nor UO_992 (O_992,N_3122,N_4255);
or UO_993 (O_993,N_2806,N_3908);
and UO_994 (O_994,N_2742,N_2629);
and UO_995 (O_995,N_2504,N_3292);
nor UO_996 (O_996,N_4205,N_3101);
and UO_997 (O_997,N_2553,N_4671);
nor UO_998 (O_998,N_2839,N_3887);
nand UO_999 (O_999,N_3243,N_4818);
endmodule