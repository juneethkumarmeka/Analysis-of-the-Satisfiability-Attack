module basic_1500_15000_2000_30_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_714,In_851);
nor U1 (N_1,In_428,In_566);
nand U2 (N_2,In_875,In_1071);
nor U3 (N_3,In_1229,In_585);
nor U4 (N_4,In_409,In_391);
nor U5 (N_5,In_582,In_1116);
nand U6 (N_6,In_93,In_55);
xnor U7 (N_7,In_1240,In_273);
nand U8 (N_8,In_716,In_833);
or U9 (N_9,In_1061,In_850);
or U10 (N_10,In_81,In_183);
nand U11 (N_11,In_1107,In_415);
and U12 (N_12,In_304,In_408);
xor U13 (N_13,In_583,In_620);
nor U14 (N_14,In_1227,In_1131);
nor U15 (N_15,In_102,In_1425);
and U16 (N_16,In_1224,In_1378);
and U17 (N_17,In_1267,In_1339);
and U18 (N_18,In_219,In_98);
xor U19 (N_19,In_788,In_1041);
nand U20 (N_20,In_691,In_883);
and U21 (N_21,In_1482,In_766);
nor U22 (N_22,In_310,In_212);
nand U23 (N_23,In_62,In_393);
and U24 (N_24,In_128,In_1443);
nand U25 (N_25,In_1178,In_39);
nand U26 (N_26,In_892,In_992);
nand U27 (N_27,In_363,In_198);
or U28 (N_28,In_1458,In_831);
and U29 (N_29,In_278,In_915);
xnor U30 (N_30,In_1044,In_1266);
nor U31 (N_31,In_160,In_323);
or U32 (N_32,In_483,In_1419);
or U33 (N_33,In_1036,In_552);
nand U34 (N_34,In_621,In_759);
xnor U35 (N_35,In_295,In_1140);
and U36 (N_36,In_1464,In_1136);
nor U37 (N_37,In_610,In_333);
xor U38 (N_38,In_424,In_594);
nand U39 (N_39,In_392,In_1189);
xor U40 (N_40,In_1194,In_107);
or U41 (N_41,In_784,In_549);
or U42 (N_42,In_988,In_254);
xor U43 (N_43,In_1334,In_403);
nand U44 (N_44,In_1110,In_478);
nor U45 (N_45,In_730,In_361);
and U46 (N_46,In_1070,In_913);
nand U47 (N_47,In_624,In_601);
and U48 (N_48,In_445,In_1310);
xnor U49 (N_49,In_1397,In_457);
xnor U50 (N_50,In_922,In_1206);
and U51 (N_51,In_68,In_1420);
nand U52 (N_52,In_359,In_365);
nor U53 (N_53,In_516,In_786);
nand U54 (N_54,In_665,In_397);
nand U55 (N_55,In_1368,In_1328);
nor U56 (N_56,In_31,In_433);
and U57 (N_57,In_1440,In_332);
nor U58 (N_58,In_614,In_802);
nand U59 (N_59,In_1415,In_1470);
and U60 (N_60,In_945,In_900);
nand U61 (N_61,In_1492,In_448);
and U62 (N_62,In_487,In_794);
nand U63 (N_63,In_490,In_570);
nor U64 (N_64,In_751,In_1104);
or U65 (N_65,In_899,In_640);
and U66 (N_66,In_1066,In_280);
nor U67 (N_67,In_949,In_436);
nor U68 (N_68,In_808,In_1283);
and U69 (N_69,In_1427,In_1150);
or U70 (N_70,In_1387,In_776);
nand U71 (N_71,In_952,In_1209);
xnor U72 (N_72,In_151,In_1028);
nor U73 (N_73,In_511,In_739);
xnor U74 (N_74,In_769,In_320);
nor U75 (N_75,In_752,In_971);
nor U76 (N_76,In_1467,In_241);
nor U77 (N_77,In_858,In_548);
or U78 (N_78,In_1393,In_1217);
xor U79 (N_79,In_1327,In_1202);
nor U80 (N_80,In_401,In_543);
nor U81 (N_81,In_667,In_700);
or U82 (N_82,In_1157,In_1304);
and U83 (N_83,In_171,In_1210);
nand U84 (N_84,In_461,In_947);
nor U85 (N_85,In_1193,In_874);
nor U86 (N_86,In_16,In_658);
and U87 (N_87,In_429,In_1456);
nand U88 (N_88,In_663,In_630);
or U89 (N_89,In_1170,In_978);
and U90 (N_90,In_1333,In_1353);
nor U91 (N_91,In_1048,In_1023);
nor U92 (N_92,In_905,In_300);
nor U93 (N_93,In_1450,In_4);
and U94 (N_94,In_1300,In_674);
or U95 (N_95,In_565,In_426);
and U96 (N_96,In_1392,In_243);
nor U97 (N_97,In_637,In_354);
nor U98 (N_98,In_239,In_1388);
xnor U99 (N_99,In_1377,In_1349);
xnor U100 (N_100,In_884,In_912);
or U101 (N_101,In_189,In_909);
nor U102 (N_102,In_1001,In_513);
xnor U103 (N_103,In_290,In_1342);
or U104 (N_104,In_449,In_411);
nor U105 (N_105,In_1158,In_1487);
and U106 (N_106,In_812,In_147);
or U107 (N_107,In_1265,In_593);
or U108 (N_108,In_231,In_1400);
xnor U109 (N_109,In_315,In_626);
nor U110 (N_110,In_1499,In_1276);
or U111 (N_111,In_417,In_58);
nor U112 (N_112,In_169,In_1137);
nor U113 (N_113,In_1059,In_272);
nand U114 (N_114,In_676,In_326);
and U115 (N_115,In_113,In_244);
xnor U116 (N_116,In_595,In_775);
nor U117 (N_117,In_1361,In_1360);
xnor U118 (N_118,In_1476,In_617);
nand U119 (N_119,In_870,In_576);
xnor U120 (N_120,In_1416,In_591);
nor U121 (N_121,In_723,In_1332);
and U122 (N_122,In_15,In_534);
nand U123 (N_123,In_250,In_18);
or U124 (N_124,In_1187,In_1122);
nor U125 (N_125,In_754,In_935);
and U126 (N_126,In_203,In_696);
or U127 (N_127,In_480,In_246);
xor U128 (N_128,In_69,In_685);
nor U129 (N_129,In_941,In_901);
or U130 (N_130,In_832,In_844);
or U131 (N_131,In_1463,In_281);
nand U132 (N_132,In_218,In_496);
nor U133 (N_133,In_1246,In_687);
nor U134 (N_134,In_1340,In_101);
and U135 (N_135,In_825,In_140);
nor U136 (N_136,In_347,In_1376);
and U137 (N_137,In_997,In_704);
nor U138 (N_138,In_934,In_73);
xnor U139 (N_139,In_167,In_589);
nand U140 (N_140,In_36,In_849);
or U141 (N_141,In_1371,In_761);
or U142 (N_142,In_406,In_951);
nor U143 (N_143,In_384,In_387);
or U144 (N_144,In_131,In_1016);
or U145 (N_145,In_1115,In_264);
nor U146 (N_146,In_651,In_762);
or U147 (N_147,In_1106,In_1483);
and U148 (N_148,In_823,In_758);
nand U149 (N_149,In_450,In_828);
or U150 (N_150,In_360,In_504);
or U151 (N_151,In_1290,In_659);
or U152 (N_152,In_917,In_514);
or U153 (N_153,In_1111,In_643);
and U154 (N_154,In_1186,In_71);
nor U155 (N_155,In_1411,In_771);
nand U156 (N_156,In_877,In_74);
nor U157 (N_157,In_503,In_763);
nor U158 (N_158,In_438,In_59);
xnor U159 (N_159,In_571,In_983);
nand U160 (N_160,In_261,In_30);
and U161 (N_161,In_33,In_1173);
nor U162 (N_162,In_404,In_1469);
or U163 (N_163,In_1155,In_1451);
and U164 (N_164,In_914,In_115);
and U165 (N_165,In_328,In_508);
nor U166 (N_166,In_108,In_1135);
xnor U167 (N_167,In_1083,In_135);
or U168 (N_168,In_600,In_611);
nand U169 (N_169,In_327,In_451);
nand U170 (N_170,In_1241,In_801);
nor U171 (N_171,In_1214,In_1268);
nand U172 (N_172,In_72,In_459);
nor U173 (N_173,In_265,In_342);
nor U174 (N_174,In_588,In_757);
nand U175 (N_175,In_827,In_956);
nor U176 (N_176,In_475,In_398);
and U177 (N_177,In_1293,In_1091);
xor U178 (N_178,In_960,In_777);
or U179 (N_179,In_190,In_148);
nor U180 (N_180,In_1174,In_930);
and U181 (N_181,In_492,In_1203);
nor U182 (N_182,In_1336,In_842);
nor U183 (N_183,In_778,In_744);
or U184 (N_184,In_535,In_252);
nor U185 (N_185,In_61,In_857);
nand U186 (N_186,In_1441,In_701);
nor U187 (N_187,In_351,In_839);
and U188 (N_188,In_998,In_214);
or U189 (N_189,In_352,In_1384);
nand U190 (N_190,In_1382,In_888);
or U191 (N_191,In_486,In_1424);
and U192 (N_192,In_928,In_863);
xor U193 (N_193,In_1218,In_105);
or U194 (N_194,In_1271,In_312);
nor U195 (N_195,In_834,In_454);
and U196 (N_196,In_50,In_27);
or U197 (N_197,In_1148,In_690);
nor U198 (N_198,In_1294,In_1068);
nand U199 (N_199,In_597,In_45);
nor U200 (N_200,In_926,In_470);
or U201 (N_201,In_558,In_89);
and U202 (N_202,In_1395,In_334);
or U203 (N_203,In_519,In_258);
nor U204 (N_204,In_100,In_1261);
nand U205 (N_205,In_1191,In_309);
xnor U206 (N_206,In_793,In_505);
and U207 (N_207,In_481,In_1330);
nand U208 (N_208,In_1277,In_1162);
and U209 (N_209,In_178,In_143);
xor U210 (N_210,In_321,In_1413);
nor U211 (N_211,In_1027,In_837);
and U212 (N_212,In_852,In_1303);
nor U213 (N_213,In_179,In_544);
nor U214 (N_214,In_1414,In_256);
and U215 (N_215,In_860,In_1350);
nand U216 (N_216,In_1329,In_554);
nor U217 (N_217,In_134,In_586);
and U218 (N_218,In_336,In_1259);
and U219 (N_219,In_790,In_880);
or U220 (N_220,In_208,In_1233);
nand U221 (N_221,In_1043,In_974);
and U222 (N_222,In_712,In_1171);
or U223 (N_223,In_52,In_871);
xnor U224 (N_224,In_639,In_152);
and U225 (N_225,In_371,In_1172);
nor U226 (N_226,In_234,In_1374);
nor U227 (N_227,In_902,In_670);
and U228 (N_228,In_965,In_1211);
or U229 (N_229,In_64,In_1185);
and U230 (N_230,In_1347,In_1236);
nor U231 (N_231,In_906,In_703);
xor U232 (N_232,In_1264,In_1497);
or U233 (N_233,In_1437,In_943);
and U234 (N_234,In_638,In_785);
and U235 (N_235,In_24,In_405);
and U236 (N_236,In_1154,In_804);
and U237 (N_237,In_287,In_1076);
xor U238 (N_238,In_201,In_694);
nor U239 (N_239,In_476,In_528);
or U240 (N_240,In_623,In_1129);
and U241 (N_241,In_897,In_1100);
nor U242 (N_242,In_237,In_1359);
nand U243 (N_243,In_137,In_255);
nand U244 (N_244,In_629,In_145);
and U245 (N_245,In_726,In_43);
and U246 (N_246,In_742,In_1121);
nor U247 (N_247,In_1285,In_668);
or U248 (N_248,In_161,In_299);
xor U249 (N_249,In_242,In_257);
xor U250 (N_250,In_976,In_331);
or U251 (N_251,In_887,In_753);
or U252 (N_252,In_38,In_42);
and U253 (N_253,In_118,In_641);
and U254 (N_254,In_939,In_881);
and U255 (N_255,In_644,In_866);
nand U256 (N_256,In_1288,In_603);
nand U257 (N_257,In_921,In_0);
and U258 (N_258,In_1495,In_1417);
and U259 (N_259,In_645,In_423);
nand U260 (N_260,In_488,In_609);
nor U261 (N_261,In_764,In_1431);
nor U262 (N_262,In_1069,In_655);
nand U263 (N_263,In_2,In_132);
nor U264 (N_264,In_185,In_985);
nor U265 (N_265,In_957,In_1446);
xnor U266 (N_266,In_1055,In_263);
nand U267 (N_267,In_1379,In_1095);
or U268 (N_268,In_1452,In_418);
or U269 (N_269,In_181,In_836);
nor U270 (N_270,In_604,In_702);
nand U271 (N_271,In_7,In_509);
and U272 (N_272,In_1181,In_865);
nor U273 (N_273,In_1337,In_968);
or U274 (N_274,In_862,In_732);
nand U275 (N_275,In_379,In_1144);
nor U276 (N_276,In_302,In_170);
and U277 (N_277,In_907,In_821);
or U278 (N_278,In_740,In_373);
or U279 (N_279,In_292,In_568);
or U280 (N_280,In_471,In_933);
xor U281 (N_281,In_104,In_106);
and U282 (N_282,In_1089,In_119);
or U283 (N_283,In_1093,In_1404);
nand U284 (N_284,In_1024,In_1295);
nor U285 (N_285,In_746,In_9);
nor U286 (N_286,In_592,In_1109);
nor U287 (N_287,In_350,In_590);
nor U288 (N_288,In_17,In_1366);
xor U289 (N_289,In_410,In_807);
and U290 (N_290,In_826,In_1117);
nor U291 (N_291,In_1432,In_247);
xor U292 (N_292,In_288,In_618);
nand U293 (N_293,In_26,In_1345);
nand U294 (N_294,In_484,In_1183);
and U295 (N_295,In_796,In_14);
and U296 (N_296,In_745,In_979);
or U297 (N_297,In_1130,In_669);
or U298 (N_298,In_1145,In_1381);
and U299 (N_299,In_1344,In_1049);
and U300 (N_300,In_349,In_1280);
nand U301 (N_301,In_79,In_1372);
nand U302 (N_302,In_1273,In_467);
nor U303 (N_303,In_1084,In_1412);
nand U304 (N_304,In_846,In_193);
xnor U305 (N_305,In_1447,In_1286);
nor U306 (N_306,In_1270,In_556);
or U307 (N_307,In_818,In_1282);
or U308 (N_308,In_579,In_307);
nand U309 (N_309,In_267,In_378);
or U310 (N_310,In_550,In_1401);
and U311 (N_311,In_1245,In_1255);
and U312 (N_312,In_961,In_814);
xnor U313 (N_313,In_491,In_1406);
nor U314 (N_314,In_274,In_525);
or U315 (N_315,In_1468,In_5);
nand U316 (N_316,In_962,In_366);
nor U317 (N_317,In_569,In_19);
nand U318 (N_318,In_416,In_1159);
and U319 (N_319,In_799,In_130);
nand U320 (N_320,In_707,In_1430);
nand U321 (N_321,In_749,In_783);
nand U322 (N_322,In_1077,In_35);
and U323 (N_323,In_1320,In_547);
nand U324 (N_324,In_1008,In_657);
or U325 (N_325,In_787,In_518);
or U326 (N_326,In_1099,In_217);
xnor U327 (N_327,In_682,In_1355);
nor U328 (N_328,In_308,In_28);
xor U329 (N_329,In_599,In_1363);
xor U330 (N_330,In_995,In_1453);
nand U331 (N_331,In_446,In_1152);
nand U332 (N_332,In_1298,In_1038);
nand U333 (N_333,In_103,In_1369);
or U334 (N_334,In_822,In_722);
and U335 (N_335,In_878,In_678);
or U336 (N_336,In_176,In_82);
and U337 (N_337,In_681,In_204);
and U338 (N_338,In_1498,In_395);
nand U339 (N_339,In_437,In_838);
xnor U340 (N_340,In_1247,In_1146);
nor U341 (N_341,In_602,In_810);
or U342 (N_342,In_1449,In_1221);
or U343 (N_343,In_559,In_233);
and U344 (N_344,In_444,In_699);
or U345 (N_345,In_577,In_1421);
nand U346 (N_346,In_537,In_898);
nand U347 (N_347,In_1390,In_1139);
xnor U348 (N_348,In_1092,In_129);
nand U349 (N_349,In_944,In_647);
and U350 (N_350,In_1317,In_1260);
nor U351 (N_351,In_1087,In_389);
or U352 (N_352,In_1465,In_277);
nor U353 (N_353,In_348,In_159);
nor U354 (N_354,In_1346,In_153);
nor U355 (N_355,In_524,In_688);
xor U356 (N_356,In_982,In_249);
and U357 (N_357,In_1205,In_1274);
nor U358 (N_358,In_847,In_861);
and U359 (N_359,In_114,In_374);
or U360 (N_360,In_1,In_1079);
and U361 (N_361,In_206,In_421);
or U362 (N_362,In_996,In_990);
and U363 (N_363,In_1284,In_209);
or U364 (N_364,In_911,In_635);
or U365 (N_365,In_236,In_708);
and U366 (N_366,In_680,In_419);
nor U367 (N_367,In_973,In_1272);
or U368 (N_368,In_684,In_29);
or U369 (N_369,In_458,In_541);
nand U370 (N_370,In_561,In_1105);
nand U371 (N_371,In_196,In_222);
nor U372 (N_372,In_1471,In_710);
or U373 (N_373,In_1075,In_743);
and U374 (N_374,In_574,In_37);
or U375 (N_375,In_824,In_622);
xnor U376 (N_376,In_380,In_1364);
and U377 (N_377,In_948,In_507);
or U378 (N_378,In_1046,In_869);
or U379 (N_379,In_1118,In_1020);
nand U380 (N_380,In_1223,In_1423);
nor U381 (N_381,In_344,In_356);
or U382 (N_382,In_1034,In_1324);
xnor U383 (N_383,In_1056,In_755);
nor U384 (N_384,In_133,In_619);
xnor U385 (N_385,In_506,In_1114);
or U386 (N_386,In_1220,In_970);
nand U387 (N_387,In_671,In_1047);
and U388 (N_388,In_184,In_362);
xnor U389 (N_389,In_1479,In_177);
and U390 (N_390,In_1442,In_1254);
or U391 (N_391,In_813,In_538);
nor U392 (N_392,In_1019,In_1493);
nor U393 (N_393,In_1169,In_469);
or U394 (N_394,In_527,In_339);
nor U395 (N_395,In_1488,In_894);
or U396 (N_396,In_1014,In_390);
or U397 (N_397,In_1323,In_522);
nand U398 (N_398,In_285,In_1040);
and U399 (N_399,In_1239,In_197);
nor U400 (N_400,In_845,In_573);
and U401 (N_401,In_1072,In_141);
and U402 (N_402,In_294,In_1439);
nand U403 (N_403,In_737,In_738);
or U404 (N_404,In_1007,In_400);
and U405 (N_405,In_422,In_495);
nand U406 (N_406,In_1200,In_425);
xnor U407 (N_407,In_1216,In_372);
nor U408 (N_408,In_1062,In_924);
and U409 (N_409,In_654,In_1184);
and U410 (N_410,In_596,In_1120);
and U411 (N_411,In_253,In_1316);
nand U412 (N_412,In_1005,In_925);
xor U413 (N_413,In_993,In_489);
nand U414 (N_414,In_1491,In_1331);
nand U415 (N_415,In_259,In_741);
and U416 (N_416,In_1409,In_367);
and U417 (N_417,In_747,In_1052);
xor U418 (N_418,In_8,In_187);
and U419 (N_419,In_1167,In_412);
and U420 (N_420,In_346,In_1480);
nor U421 (N_421,In_864,In_512);
and U422 (N_422,In_1385,In_1029);
and U423 (N_423,In_432,In_493);
nor U424 (N_424,In_715,In_632);
or U425 (N_425,In_1164,In_22);
xnor U426 (N_426,In_608,In_1269);
or U427 (N_427,In_482,In_13);
nand U428 (N_428,In_1188,In_648);
nand U429 (N_429,In_464,In_1011);
nand U430 (N_430,In_1179,In_1238);
nand U431 (N_431,In_1230,In_268);
and U432 (N_432,In_1315,In_317);
xnor U433 (N_433,In_567,In_1134);
and U434 (N_434,In_182,In_683);
and U435 (N_435,In_724,In_1396);
or U436 (N_436,In_1389,In_442);
or U437 (N_437,In_1006,In_805);
nor U438 (N_438,In_245,In_1244);
nor U439 (N_439,In_498,In_439);
xor U440 (N_440,In_86,In_499);
and U441 (N_441,In_6,In_555);
and U442 (N_442,In_1082,In_1094);
nand U443 (N_443,In_664,In_1318);
nor U444 (N_444,In_291,In_1090);
or U445 (N_445,In_918,In_936);
and U446 (N_446,In_1484,In_606);
nand U447 (N_447,In_735,In_1481);
nor U448 (N_448,In_109,In_774);
and U449 (N_449,In_841,In_867);
nor U450 (N_450,In_1213,In_1243);
nor U451 (N_451,In_1128,In_329);
or U452 (N_452,In_44,In_235);
nor U453 (N_453,In_843,In_1305);
or U454 (N_454,In_1362,In_848);
nand U455 (N_455,In_338,In_1461);
nor U456 (N_456,In_1462,In_1042);
nor U457 (N_457,In_205,In_238);
or U458 (N_458,In_1457,In_817);
nand U459 (N_459,In_275,In_456);
and U460 (N_460,In_840,In_1478);
or U461 (N_461,In_165,In_697);
or U462 (N_462,In_1035,In_337);
or U463 (N_463,In_23,In_1031);
nor U464 (N_464,In_500,In_1250);
nor U465 (N_465,In_815,In_1065);
or U466 (N_466,In_1289,In_560);
and U467 (N_467,In_90,In_795);
or U468 (N_468,In_904,In_10);
nand U469 (N_469,In_210,In_46);
nand U470 (N_470,In_502,In_276);
and U471 (N_471,In_314,In_1141);
nand U472 (N_472,In_903,In_1474);
nand U473 (N_473,In_1226,In_293);
or U474 (N_474,In_1103,In_660);
and U475 (N_475,In_67,In_455);
or U476 (N_476,In_1428,In_497);
and U477 (N_477,In_859,In_199);
or U478 (N_478,In_953,In_124);
and U479 (N_479,In_138,In_616);
or U480 (N_480,In_1215,In_123);
and U481 (N_481,In_311,In_1367);
and U482 (N_482,In_1190,In_40);
nand U483 (N_483,In_1033,In_959);
nand U484 (N_484,In_927,In_111);
nor U485 (N_485,In_76,In_646);
xor U486 (N_486,In_972,In_1196);
and U487 (N_487,In_1127,In_25);
and U488 (N_488,In_937,In_240);
nor U489 (N_489,In_1078,In_1138);
nor U490 (N_490,In_1192,In_48);
or U491 (N_491,In_895,In_650);
or U492 (N_492,In_780,In_431);
and U493 (N_493,In_1301,In_1197);
xnor U494 (N_494,In_958,In_158);
nand U495 (N_495,In_226,In_144);
or U496 (N_496,In_121,In_1161);
and U497 (N_497,In_180,In_501);
nor U498 (N_498,In_531,In_946);
xnor U499 (N_499,In_453,In_1195);
and U500 (N_500,In_1113,In_386);
nor U501 (N_501,In_1370,In_540);
and U502 (N_502,In_353,In_835);
nand U503 (N_503,In_1199,N_416);
nand U504 (N_504,In_1352,In_1380);
or U505 (N_505,In_675,N_257);
nand U506 (N_506,In_381,In_673);
nor U507 (N_507,N_57,N_383);
or U508 (N_508,N_42,N_166);
or U509 (N_509,In_270,In_720);
or U510 (N_510,N_445,In_1263);
nor U511 (N_511,N_79,In_57);
nor U512 (N_512,N_335,N_275);
nand U513 (N_513,N_248,N_112);
and U514 (N_514,N_281,In_1088);
or U515 (N_515,N_88,In_394);
or U516 (N_516,In_1287,N_124);
nand U517 (N_517,In_873,In_553);
and U518 (N_518,N_482,N_480);
or U519 (N_519,N_341,In_283);
xor U520 (N_520,N_56,N_110);
or U521 (N_521,N_152,N_286);
or U522 (N_522,In_466,N_435);
or U523 (N_523,N_154,N_153);
nand U524 (N_524,In_91,N_486);
and U525 (N_525,In_1234,N_121);
nor U526 (N_526,N_179,N_247);
nor U527 (N_527,In_83,N_293);
nor U528 (N_528,In_1151,N_54);
nor U529 (N_529,In_1278,In_1383);
and U530 (N_530,In_262,N_374);
and U531 (N_531,In_441,N_89);
or U532 (N_532,In_1039,N_401);
or U533 (N_533,N_447,N_317);
xnor U534 (N_534,N_464,In_584);
xor U535 (N_535,In_191,N_109);
nor U536 (N_536,In_440,In_142);
or U537 (N_537,N_135,In_811);
nor U538 (N_538,N_332,In_709);
or U539 (N_539,N_351,N_60);
nor U540 (N_540,In_931,N_246);
nor U541 (N_541,N_323,N_45);
nand U542 (N_542,In_1426,In_791);
and U543 (N_543,N_240,N_303);
and U544 (N_544,N_188,N_59);
and U545 (N_545,In_886,In_1489);
or U546 (N_546,N_236,In_1455);
nor U547 (N_547,In_613,N_47);
nor U548 (N_548,N_470,N_251);
nand U549 (N_549,In_1050,N_143);
xor U550 (N_550,In_1351,In_929);
and U551 (N_551,N_51,N_245);
nand U552 (N_552,In_224,N_333);
nand U553 (N_553,N_499,In_164);
nor U554 (N_554,In_731,In_230);
and U555 (N_555,N_487,N_216);
nand U556 (N_556,N_127,N_313);
and U557 (N_557,In_202,In_1321);
nor U558 (N_558,N_363,N_226);
nor U559 (N_559,In_967,N_162);
nand U560 (N_560,In_662,In_1208);
xnor U561 (N_561,N_64,In_1433);
or U562 (N_562,N_425,N_271);
and U563 (N_563,N_442,In_1054);
nand U564 (N_564,In_383,N_25);
or U565 (N_565,N_171,N_481);
or U566 (N_566,N_96,In_1309);
or U567 (N_567,N_410,N_324);
and U568 (N_568,N_209,In_1472);
nand U569 (N_569,In_54,In_760);
nand U570 (N_570,In_297,In_211);
nor U571 (N_571,N_190,In_462);
nor U572 (N_572,In_542,N_299);
nand U573 (N_573,N_229,In_1257);
xor U574 (N_574,N_104,N_373);
and U575 (N_575,N_189,In_1022);
nor U576 (N_576,In_162,In_335);
nor U577 (N_577,In_1133,In_910);
and U578 (N_578,N_268,In_885);
nand U579 (N_579,N_367,N_419);
or U580 (N_580,In_581,N_231);
and U581 (N_581,N_202,N_39);
nor U582 (N_582,In_1073,In_194);
nand U583 (N_583,In_789,In_175);
nand U584 (N_584,In_572,N_457);
xnor U585 (N_585,N_241,In_955);
or U586 (N_586,In_987,N_78);
nand U587 (N_587,N_87,In_521);
nand U588 (N_588,N_289,N_441);
nor U589 (N_589,N_267,N_430);
nand U590 (N_590,In_1444,In_1126);
nand U591 (N_591,In_896,In_303);
nor U592 (N_592,In_1163,In_1102);
and U593 (N_593,N_455,N_163);
nand U594 (N_594,In_1053,In_1002);
and U595 (N_595,In_1375,In_345);
and U596 (N_596,In_563,In_994);
or U597 (N_597,In_318,In_56);
and U598 (N_598,N_312,In_92);
and U599 (N_599,In_631,N_46);
or U600 (N_600,N_6,In_1057);
nand U601 (N_601,In_260,In_78);
and U602 (N_602,In_1232,In_963);
nand U603 (N_603,In_376,N_309);
or U604 (N_604,N_398,In_174);
and U605 (N_605,In_340,N_95);
and U606 (N_606,In_1299,In_1182);
nor U607 (N_607,In_472,N_352);
nor U608 (N_608,In_1410,In_652);
or U609 (N_609,N_205,N_68);
nand U610 (N_610,In_473,In_1281);
and U611 (N_611,In_51,N_195);
nand U612 (N_612,In_942,In_1262);
nand U613 (N_613,N_469,In_364);
and U614 (N_614,N_26,N_33);
and U615 (N_615,N_250,N_227);
nand U616 (N_616,In_923,In_1296);
or U617 (N_617,N_219,N_478);
and U618 (N_618,N_73,In_341);
or U619 (N_619,N_28,In_698);
nand U620 (N_620,In_649,N_149);
and U621 (N_621,N_284,In_729);
and U622 (N_622,N_402,N_167);
xnor U623 (N_623,In_872,N_392);
or U624 (N_624,In_1132,In_156);
or U625 (N_625,In_578,In_279);
nand U626 (N_626,N_197,In_494);
xnor U627 (N_627,N_370,N_156);
or U628 (N_628,N_242,In_725);
or U629 (N_629,N_111,N_473);
nor U630 (N_630,N_123,N_360);
and U631 (N_631,N_41,In_986);
and U632 (N_632,N_278,N_22);
nand U633 (N_633,N_142,N_67);
or U634 (N_634,In_319,In_1123);
xnor U635 (N_635,N_307,In_402);
nor U636 (N_636,In_32,N_66);
xor U637 (N_637,N_12,In_85);
nor U638 (N_638,In_34,N_400);
nor U639 (N_639,In_284,N_159);
nor U640 (N_640,In_188,In_1060);
and U641 (N_641,In_797,In_479);
and U642 (N_642,In_1494,N_338);
xnor U643 (N_643,N_431,N_220);
nor U644 (N_644,In_1386,In_313);
nand U645 (N_645,In_413,N_65);
nand U646 (N_646,In_248,N_40);
or U647 (N_647,In_53,N_43);
or U648 (N_648,N_349,N_155);
nor U649 (N_649,In_1147,N_388);
nor U650 (N_650,In_1175,N_255);
nor U651 (N_651,N_35,N_412);
nand U652 (N_652,N_18,N_382);
or U653 (N_653,N_193,N_343);
or U654 (N_654,N_378,In_615);
or U655 (N_655,In_661,N_477);
nand U656 (N_656,In_1045,N_20);
xnor U657 (N_657,In_65,In_1422);
xor U658 (N_658,In_1017,In_1198);
or U659 (N_659,In_1004,N_458);
nand U660 (N_660,In_1242,In_1252);
and U661 (N_661,In_330,In_692);
nand U662 (N_662,N_376,In_186);
nor U663 (N_663,N_1,N_172);
or U664 (N_664,In_536,N_235);
nand U665 (N_665,In_207,In_803);
nor U666 (N_666,N_224,N_23);
xnor U667 (N_667,N_350,N_183);
or U668 (N_668,N_479,In_225);
xnor U669 (N_669,N_223,In_1064);
and U670 (N_670,N_315,In_1436);
and U671 (N_671,N_140,In_435);
nand U672 (N_672,N_75,N_21);
nand U673 (N_673,In_1222,N_347);
and U674 (N_674,In_1097,In_298);
or U675 (N_675,In_125,In_964);
and U676 (N_676,In_88,N_280);
nand U677 (N_677,N_192,In_1357);
nand U678 (N_678,In_1026,In_1166);
and U679 (N_679,In_1438,In_1063);
or U680 (N_680,N_102,N_474);
or U681 (N_681,In_1405,In_1085);
nand U682 (N_682,In_520,In_430);
and U683 (N_683,In_1338,In_122);
and U684 (N_684,In_155,In_1398);
nand U685 (N_685,N_186,In_1000);
or U686 (N_686,N_308,In_1399);
nand U687 (N_687,In_414,In_1275);
and U688 (N_688,N_443,In_1365);
or U689 (N_689,N_476,N_471);
and U690 (N_690,In_1475,N_37);
nand U691 (N_691,In_721,In_636);
nor U692 (N_692,N_133,In_1403);
or U693 (N_693,N_85,In_1249);
and U694 (N_694,N_494,N_175);
and U695 (N_695,N_314,N_161);
or U696 (N_696,In_713,N_379);
or U697 (N_697,In_60,In_213);
nor U698 (N_698,In_666,N_92);
nand U699 (N_699,N_488,In_447);
nor U700 (N_700,N_173,In_1319);
nor U701 (N_701,N_8,N_258);
and U702 (N_702,In_605,N_94);
and U703 (N_703,N_264,In_221);
nand U704 (N_704,In_1153,In_301);
and U705 (N_705,In_999,N_483);
or U706 (N_706,In_728,In_358);
nand U707 (N_707,In_551,N_145);
nand U708 (N_708,N_237,In_733);
xor U709 (N_709,N_141,N_105);
or U710 (N_710,In_316,In_1256);
nor U711 (N_711,In_434,In_1302);
and U712 (N_712,In_216,N_261);
nand U713 (N_713,In_768,N_125);
xnor U714 (N_714,N_468,N_32);
and U715 (N_715,In_1394,In_168);
and U716 (N_716,N_326,N_201);
or U717 (N_717,In_1248,N_475);
or U718 (N_718,In_1490,N_428);
or U719 (N_719,In_1165,N_148);
nor U720 (N_720,N_128,N_492);
nor U721 (N_721,N_437,N_342);
nand U722 (N_722,In_546,In_868);
nor U723 (N_723,In_1225,N_331);
or U724 (N_724,In_463,N_69);
or U725 (N_725,N_348,In_1253);
nor U726 (N_726,In_325,N_218);
xnor U727 (N_727,In_679,In_950);
nor U728 (N_728,In_460,In_628);
or U729 (N_729,In_1292,N_456);
nor U730 (N_730,N_199,In_1448);
or U731 (N_731,In_1032,In_529);
xnor U732 (N_732,N_265,In_1018);
and U733 (N_733,In_1402,N_221);
or U734 (N_734,In_587,N_361);
xor U735 (N_735,In_1343,In_653);
and U736 (N_736,N_157,In_1108);
or U737 (N_737,In_695,In_117);
nand U738 (N_738,N_176,In_474);
nor U739 (N_739,N_337,N_31);
nand U740 (N_740,N_48,In_1015);
and U741 (N_741,In_557,N_10);
nor U742 (N_742,In_1021,In_70);
or U743 (N_743,N_296,N_164);
nand U744 (N_744,In_1312,N_485);
nor U745 (N_745,In_809,N_346);
xnor U746 (N_746,In_677,N_44);
nor U747 (N_747,N_119,In_1391);
or U748 (N_748,N_198,N_321);
nand U749 (N_749,In_1201,In_966);
nor U750 (N_750,In_782,N_403);
or U751 (N_751,In_127,In_1435);
nor U752 (N_752,In_1168,N_362);
and U753 (N_753,N_459,In_286);
nor U754 (N_754,N_182,In_1354);
and U755 (N_755,N_397,N_83);
nand U756 (N_756,In_633,N_290);
nand U757 (N_757,N_463,In_1418);
nand U758 (N_758,In_919,In_539);
nand U759 (N_759,N_387,N_353);
or U760 (N_760,N_34,N_239);
nor U761 (N_761,In_1156,N_49);
and U762 (N_762,In_1496,N_233);
or U763 (N_763,In_21,In_1485);
and U764 (N_764,In_220,In_792);
nor U765 (N_765,In_781,N_263);
or U766 (N_766,N_160,In_120);
nor U767 (N_767,In_932,N_300);
xor U768 (N_768,N_270,In_1341);
nand U769 (N_769,In_136,N_30);
nor U770 (N_770,N_191,In_269);
nand U771 (N_771,N_204,N_11);
and U772 (N_772,N_62,In_916);
xor U773 (N_773,N_151,N_404);
nor U774 (N_774,In_1325,In_893);
and U775 (N_775,In_1080,N_100);
and U776 (N_776,N_215,N_0);
or U777 (N_777,N_15,N_413);
nor U778 (N_778,N_150,N_139);
nand U779 (N_779,N_276,N_391);
nand U780 (N_780,N_107,In_271);
and U781 (N_781,In_95,N_394);
and U782 (N_782,N_116,In_830);
xor U783 (N_783,N_336,N_279);
nand U784 (N_784,N_210,N_439);
or U785 (N_785,In_940,In_452);
xor U786 (N_786,In_1279,In_1306);
xor U787 (N_787,In_1149,N_364);
nor U788 (N_788,In_580,N_345);
and U789 (N_789,N_212,In_756);
nor U790 (N_790,In_1012,N_327);
nand U791 (N_791,In_1180,N_385);
and U792 (N_792,N_408,In_195);
and U793 (N_793,N_436,N_446);
xor U794 (N_794,N_243,In_533);
and U795 (N_795,In_399,In_266);
nor U796 (N_796,In_232,In_607);
nand U797 (N_797,N_266,N_415);
nor U798 (N_798,N_424,N_63);
and U799 (N_799,In_355,In_882);
or U800 (N_800,In_1030,N_355);
and U801 (N_801,N_365,N_302);
or U802 (N_802,In_1466,N_228);
and U803 (N_803,N_287,N_70);
nand U804 (N_804,N_136,In_375);
and U805 (N_805,N_366,N_433);
nor U806 (N_806,In_1434,In_172);
nand U807 (N_807,N_106,N_414);
or U808 (N_808,In_146,N_249);
xor U809 (N_809,In_343,In_289);
or U810 (N_810,In_150,N_187);
or U811 (N_811,In_1212,In_154);
or U812 (N_812,In_736,N_418);
nor U813 (N_813,N_294,N_3);
xnor U814 (N_814,N_304,N_399);
xnor U815 (N_815,In_969,N_438);
or U816 (N_816,N_498,In_1112);
and U817 (N_817,In_642,N_449);
nor U818 (N_818,N_291,In_523);
nor U819 (N_819,In_1251,In_532);
nand U820 (N_820,In_718,N_207);
or U821 (N_821,In_1311,N_80);
or U822 (N_822,In_1096,N_217);
nand U823 (N_823,N_377,N_375);
nor U824 (N_824,N_423,In_94);
nor U825 (N_825,N_452,In_96);
nor U826 (N_826,N_465,N_101);
nand U827 (N_827,N_138,In_820);
nand U828 (N_828,In_526,In_477);
nor U829 (N_829,N_434,In_1373);
or U830 (N_830,N_126,In_1160);
nor U831 (N_831,N_200,N_320);
or U832 (N_832,In_99,In_750);
xnor U833 (N_833,N_7,In_1086);
nand U834 (N_834,In_1010,N_84);
and U835 (N_835,In_706,N_82);
nor U836 (N_836,N_211,In_854);
and U837 (N_837,N_17,In_1308);
or U838 (N_838,In_192,In_984);
or U839 (N_839,N_24,N_120);
xnor U840 (N_840,In_686,In_1025);
nor U841 (N_841,N_395,N_472);
xor U842 (N_842,In_306,In_980);
nand U843 (N_843,In_420,In_1231);
nand U844 (N_844,In_1460,N_311);
or U845 (N_845,N_467,In_1408);
or U846 (N_846,N_253,In_3);
nand U847 (N_847,N_356,In_1258);
nor U848 (N_848,N_232,In_1009);
and U849 (N_849,In_829,In_1291);
nor U850 (N_850,In_672,N_390);
and U851 (N_851,N_178,N_386);
and U852 (N_852,In_634,N_177);
nand U853 (N_853,In_20,N_393);
and U854 (N_854,N_260,In_296);
and U855 (N_855,In_116,N_493);
and U856 (N_856,N_357,In_1037);
or U857 (N_857,N_371,N_180);
nor U858 (N_858,N_273,In_856);
or U859 (N_859,In_1297,In_1407);
nor U860 (N_860,In_368,N_234);
xor U861 (N_861,N_14,N_460);
nor U862 (N_862,In_173,In_77);
or U863 (N_863,N_117,N_339);
xnor U864 (N_864,N_427,In_1124);
nor U865 (N_865,In_377,In_806);
or U866 (N_866,N_497,In_1013);
or U867 (N_867,In_819,In_1326);
and U868 (N_868,In_1356,N_318);
and U869 (N_869,In_625,In_388);
or U870 (N_870,In_1429,N_194);
nand U871 (N_871,N_448,N_491);
xnor U872 (N_872,N_86,N_196);
nor U873 (N_873,In_530,In_765);
nand U874 (N_874,N_55,N_292);
nand U875 (N_875,N_131,N_19);
or U876 (N_876,In_517,In_1477);
xor U877 (N_877,N_462,N_130);
nor U878 (N_878,N_359,In_1486);
or U879 (N_879,In_989,In_215);
and U880 (N_880,In_656,N_169);
or U881 (N_881,N_214,N_36);
or U882 (N_882,N_340,In_954);
and U883 (N_883,In_223,In_427);
nor U884 (N_884,N_283,In_1207);
or U885 (N_885,In_1067,In_1142);
or U886 (N_886,N_108,N_181);
and U887 (N_887,N_13,In_1119);
nor U888 (N_888,In_12,N_432);
or U889 (N_889,In_1098,N_238);
nand U890 (N_890,N_310,In_1228);
and U891 (N_891,In_800,N_396);
nand U892 (N_892,N_454,In_562);
nand U893 (N_893,In_1051,N_38);
nand U894 (N_894,N_76,In_1473);
nand U895 (N_895,In_734,In_97);
nor U896 (N_896,In_1003,N_453);
xnor U897 (N_897,In_991,N_417);
or U898 (N_898,N_222,In_689);
and U899 (N_899,In_891,N_58);
and U900 (N_900,N_206,In_981);
or U901 (N_901,N_113,In_227);
nand U902 (N_902,In_228,N_134);
xnor U903 (N_903,N_262,In_49);
and U904 (N_904,In_748,N_225);
or U905 (N_905,In_282,In_1313);
or U906 (N_906,In_382,N_496);
or U907 (N_907,N_184,N_203);
and U908 (N_908,In_47,In_1143);
xnor U909 (N_909,N_165,In_719);
and U910 (N_910,N_252,In_798);
nand U911 (N_911,In_767,In_575);
nor U912 (N_912,N_298,N_484);
nand U913 (N_913,In_515,N_407);
nand U914 (N_914,In_772,In_975);
nand U915 (N_915,N_354,N_269);
nor U916 (N_916,N_288,In_163);
and U917 (N_917,N_490,N_322);
or U918 (N_918,In_396,N_384);
nand U919 (N_919,In_773,N_144);
xor U920 (N_920,In_1445,N_50);
and U921 (N_921,N_90,In_1237);
and U922 (N_922,N_495,In_166);
or U923 (N_923,N_132,In_564);
nor U924 (N_924,N_5,N_440);
nand U925 (N_925,N_461,In_1204);
or U926 (N_926,In_126,In_465);
and U927 (N_927,N_295,N_115);
nor U928 (N_928,In_855,N_168);
xnor U929 (N_929,N_137,In_853);
or U930 (N_930,N_213,N_369);
nor U931 (N_931,N_185,In_1314);
or U932 (N_932,N_426,In_139);
or U933 (N_933,N_358,In_385);
nor U934 (N_934,In_305,N_380);
nand U935 (N_935,In_41,N_429);
xor U936 (N_936,In_627,In_80);
nor U937 (N_937,In_1219,N_421);
nor U938 (N_938,In_1235,N_329);
and U939 (N_939,In_876,N_305);
or U940 (N_940,In_200,N_98);
nor U941 (N_941,N_301,N_256);
or U942 (N_942,N_53,N_319);
nand U943 (N_943,N_277,N_328);
or U944 (N_944,In_1101,In_816);
nand U945 (N_945,In_63,In_87);
nor U946 (N_946,In_149,N_450);
and U947 (N_947,N_230,N_72);
xnor U948 (N_948,In_727,In_370);
and U949 (N_949,In_545,N_451);
nand U950 (N_950,N_334,N_444);
xor U951 (N_951,In_1058,N_97);
xnor U952 (N_952,In_879,In_1074);
nor U953 (N_953,N_285,In_11);
or U954 (N_954,N_297,In_84);
and U955 (N_955,In_110,N_420);
nor U956 (N_956,N_406,In_322);
nor U957 (N_957,N_174,In_938);
nor U958 (N_958,N_2,N_147);
nor U959 (N_959,In_369,In_711);
nor U960 (N_960,N_306,In_324);
nor U961 (N_961,N_272,N_4);
or U962 (N_962,N_259,In_66);
nor U963 (N_963,In_1081,In_407);
nand U964 (N_964,N_103,In_357);
xnor U965 (N_965,N_244,N_389);
nand U966 (N_966,N_381,N_146);
nand U967 (N_967,N_122,N_409);
and U968 (N_968,N_9,In_889);
xnor U969 (N_969,N_325,In_598);
nor U970 (N_970,N_422,N_158);
xor U971 (N_971,N_254,In_717);
or U972 (N_972,N_74,In_1459);
nand U973 (N_973,In_1348,N_368);
nand U974 (N_974,In_693,N_61);
or U975 (N_975,In_1177,In_890);
nor U976 (N_976,N_129,N_372);
nand U977 (N_977,In_251,In_1176);
or U978 (N_978,N_405,In_443);
and U979 (N_979,N_466,In_1322);
or U980 (N_980,N_27,N_170);
or U981 (N_981,In_468,In_908);
nand U982 (N_982,N_93,In_920);
and U983 (N_983,In_705,In_485);
and U984 (N_984,N_16,In_612);
or U985 (N_985,In_112,N_91);
xor U986 (N_986,N_330,In_157);
nand U987 (N_987,N_411,In_1307);
and U988 (N_988,In_779,In_1454);
nor U989 (N_989,N_99,N_114);
nand U990 (N_990,N_274,In_75);
and U991 (N_991,In_1125,N_489);
nor U992 (N_992,N_77,N_29);
xor U993 (N_993,In_510,In_977);
and U994 (N_994,N_118,N_316);
nor U995 (N_995,N_282,N_71);
nand U996 (N_996,In_1358,In_1335);
nand U997 (N_997,In_229,N_208);
and U998 (N_998,In_770,N_344);
or U999 (N_999,N_52,N_81);
or U1000 (N_1000,N_508,N_869);
nor U1001 (N_1001,N_976,N_915);
or U1002 (N_1002,N_536,N_700);
and U1003 (N_1003,N_801,N_964);
and U1004 (N_1004,N_583,N_658);
or U1005 (N_1005,N_659,N_704);
nand U1006 (N_1006,N_682,N_766);
nand U1007 (N_1007,N_809,N_894);
nand U1008 (N_1008,N_714,N_965);
xor U1009 (N_1009,N_823,N_604);
or U1010 (N_1010,N_875,N_743);
and U1011 (N_1011,N_722,N_789);
xnor U1012 (N_1012,N_500,N_834);
or U1013 (N_1013,N_958,N_685);
nor U1014 (N_1014,N_668,N_721);
or U1015 (N_1015,N_888,N_776);
or U1016 (N_1016,N_567,N_832);
and U1017 (N_1017,N_913,N_863);
nor U1018 (N_1018,N_858,N_650);
and U1019 (N_1019,N_754,N_527);
and U1020 (N_1020,N_708,N_826);
nand U1021 (N_1021,N_727,N_608);
nor U1022 (N_1022,N_720,N_988);
nor U1023 (N_1023,N_734,N_916);
and U1024 (N_1024,N_849,N_639);
xor U1025 (N_1025,N_865,N_502);
xnor U1026 (N_1026,N_590,N_617);
nor U1027 (N_1027,N_748,N_752);
nor U1028 (N_1028,N_575,N_841);
and U1029 (N_1029,N_963,N_648);
and U1030 (N_1030,N_615,N_821);
and U1031 (N_1031,N_605,N_645);
nand U1032 (N_1032,N_936,N_808);
nor U1033 (N_1033,N_922,N_635);
nor U1034 (N_1034,N_982,N_678);
or U1035 (N_1035,N_599,N_642);
and U1036 (N_1036,N_800,N_825);
nor U1037 (N_1037,N_530,N_879);
and U1038 (N_1038,N_581,N_920);
nor U1039 (N_1039,N_926,N_775);
and U1040 (N_1040,N_514,N_791);
or U1041 (N_1041,N_562,N_880);
nand U1042 (N_1042,N_819,N_525);
nor U1043 (N_1043,N_790,N_519);
nand U1044 (N_1044,N_881,N_620);
xnor U1045 (N_1045,N_522,N_701);
xor U1046 (N_1046,N_598,N_890);
or U1047 (N_1047,N_961,N_884);
or U1048 (N_1048,N_625,N_867);
nor U1049 (N_1049,N_957,N_626);
or U1050 (N_1050,N_883,N_864);
xor U1051 (N_1051,N_795,N_836);
nor U1052 (N_1052,N_991,N_877);
nand U1053 (N_1053,N_702,N_686);
nor U1054 (N_1054,N_785,N_955);
xnor U1055 (N_1055,N_802,N_588);
and U1056 (N_1056,N_859,N_874);
or U1057 (N_1057,N_813,N_528);
or U1058 (N_1058,N_811,N_644);
and U1059 (N_1059,N_649,N_968);
nand U1060 (N_1060,N_699,N_548);
nor U1061 (N_1061,N_878,N_917);
and U1062 (N_1062,N_866,N_844);
and U1063 (N_1063,N_543,N_824);
nand U1064 (N_1064,N_990,N_895);
nor U1065 (N_1065,N_940,N_549);
nor U1066 (N_1066,N_524,N_749);
and U1067 (N_1067,N_898,N_511);
and U1068 (N_1068,N_691,N_715);
and U1069 (N_1069,N_983,N_818);
or U1070 (N_1070,N_560,N_728);
or U1071 (N_1071,N_788,N_593);
nand U1072 (N_1072,N_725,N_817);
nand U1073 (N_1073,N_710,N_535);
or U1074 (N_1074,N_646,N_756);
nor U1075 (N_1075,N_633,N_746);
nor U1076 (N_1076,N_774,N_778);
or U1077 (N_1077,N_794,N_768);
nand U1078 (N_1078,N_741,N_882);
xnor U1079 (N_1079,N_661,N_896);
nand U1080 (N_1080,N_671,N_759);
or U1081 (N_1081,N_757,N_815);
or U1082 (N_1082,N_838,N_529);
nor U1083 (N_1083,N_840,N_871);
nor U1084 (N_1084,N_510,N_600);
or U1085 (N_1085,N_925,N_724);
nor U1086 (N_1086,N_951,N_876);
or U1087 (N_1087,N_665,N_541);
or U1088 (N_1088,N_980,N_960);
and U1089 (N_1089,N_807,N_566);
xor U1090 (N_1090,N_651,N_814);
nor U1091 (N_1091,N_780,N_868);
and U1092 (N_1092,N_504,N_911);
and U1093 (N_1093,N_934,N_655);
nor U1094 (N_1094,N_923,N_718);
nor U1095 (N_1095,N_556,N_733);
or U1096 (N_1096,N_565,N_989);
xnor U1097 (N_1097,N_779,N_770);
nor U1098 (N_1098,N_924,N_979);
or U1099 (N_1099,N_705,N_892);
nand U1100 (N_1100,N_767,N_506);
nand U1101 (N_1101,N_576,N_953);
nand U1102 (N_1102,N_555,N_601);
and U1103 (N_1103,N_579,N_580);
and U1104 (N_1104,N_613,N_551);
nand U1105 (N_1105,N_603,N_930);
or U1106 (N_1106,N_696,N_634);
nor U1107 (N_1107,N_783,N_845);
nor U1108 (N_1108,N_638,N_706);
and U1109 (N_1109,N_798,N_839);
nand U1110 (N_1110,N_792,N_739);
and U1111 (N_1111,N_669,N_578);
nor U1112 (N_1112,N_908,N_829);
or U1113 (N_1113,N_697,N_899);
nand U1114 (N_1114,N_550,N_750);
nand U1115 (N_1115,N_657,N_545);
nand U1116 (N_1116,N_861,N_939);
nor U1117 (N_1117,N_676,N_558);
or U1118 (N_1118,N_698,N_969);
nor U1119 (N_1119,N_931,N_542);
nand U1120 (N_1120,N_501,N_656);
nand U1121 (N_1121,N_966,N_831);
and U1122 (N_1122,N_744,N_606);
or U1123 (N_1123,N_629,N_816);
or U1124 (N_1124,N_632,N_610);
xor U1125 (N_1125,N_544,N_731);
nand U1126 (N_1126,N_607,N_828);
xor U1127 (N_1127,N_797,N_897);
and U1128 (N_1128,N_573,N_730);
and U1129 (N_1129,N_747,N_726);
or U1130 (N_1130,N_666,N_860);
xnor U1131 (N_1131,N_689,N_855);
and U1132 (N_1132,N_850,N_589);
and U1133 (N_1133,N_932,N_793);
xor U1134 (N_1134,N_561,N_812);
and U1135 (N_1135,N_919,N_518);
xnor U1136 (N_1136,N_942,N_630);
nand U1137 (N_1137,N_810,N_695);
or U1138 (N_1138,N_787,N_835);
nor U1139 (N_1139,N_672,N_538);
xnor U1140 (N_1140,N_893,N_950);
nand U1141 (N_1141,N_554,N_712);
or U1142 (N_1142,N_609,N_948);
nor U1143 (N_1143,N_777,N_856);
nor U1144 (N_1144,N_675,N_563);
nor U1145 (N_1145,N_660,N_827);
nor U1146 (N_1146,N_516,N_684);
xor U1147 (N_1147,N_941,N_967);
nand U1148 (N_1148,N_843,N_833);
nand U1149 (N_1149,N_614,N_738);
nor U1150 (N_1150,N_673,N_984);
nor U1151 (N_1151,N_690,N_719);
or U1152 (N_1152,N_803,N_570);
or U1153 (N_1153,N_621,N_667);
and U1154 (N_1154,N_526,N_582);
xnor U1155 (N_1155,N_933,N_680);
and U1156 (N_1156,N_995,N_531);
or U1157 (N_1157,N_901,N_758);
xor U1158 (N_1158,N_569,N_938);
nor U1159 (N_1159,N_977,N_972);
nor U1160 (N_1160,N_799,N_641);
nor U1161 (N_1161,N_574,N_905);
nand U1162 (N_1162,N_717,N_513);
and U1163 (N_1163,N_643,N_568);
nor U1164 (N_1164,N_996,N_847);
nand U1165 (N_1165,N_796,N_918);
nor U1166 (N_1166,N_854,N_520);
nor U1167 (N_1167,N_975,N_970);
nand U1168 (N_1168,N_993,N_611);
or U1169 (N_1169,N_912,N_753);
or U1170 (N_1170,N_822,N_851);
or U1171 (N_1171,N_585,N_902);
and U1172 (N_1172,N_534,N_755);
or U1173 (N_1173,N_540,N_857);
nor U1174 (N_1174,N_713,N_886);
nand U1175 (N_1175,N_740,N_662);
and U1176 (N_1176,N_547,N_559);
or U1177 (N_1177,N_679,N_505);
nor U1178 (N_1178,N_956,N_592);
and U1179 (N_1179,N_557,N_729);
nor U1180 (N_1180,N_806,N_987);
and U1181 (N_1181,N_962,N_946);
nor U1182 (N_1182,N_670,N_910);
nor U1183 (N_1183,N_891,N_521);
nand U1184 (N_1184,N_586,N_602);
nor U1185 (N_1185,N_654,N_677);
nor U1186 (N_1186,N_782,N_873);
and U1187 (N_1187,N_949,N_596);
and U1188 (N_1188,N_769,N_994);
nor U1189 (N_1189,N_591,N_723);
xnor U1190 (N_1190,N_537,N_647);
and U1191 (N_1191,N_587,N_954);
nor U1192 (N_1192,N_546,N_903);
xnor U1193 (N_1193,N_564,N_862);
nor U1194 (N_1194,N_532,N_999);
nor U1195 (N_1195,N_929,N_636);
and U1196 (N_1196,N_853,N_765);
or U1197 (N_1197,N_889,N_703);
or U1198 (N_1198,N_577,N_640);
and U1199 (N_1199,N_732,N_927);
or U1200 (N_1200,N_503,N_928);
nor U1201 (N_1201,N_664,N_781);
xor U1202 (N_1202,N_515,N_687);
and U1203 (N_1203,N_618,N_992);
nand U1204 (N_1204,N_997,N_947);
and U1205 (N_1205,N_552,N_623);
nor U1206 (N_1206,N_681,N_761);
nor U1207 (N_1207,N_907,N_909);
nand U1208 (N_1208,N_597,N_805);
nand U1209 (N_1209,N_595,N_986);
nor U1210 (N_1210,N_981,N_572);
and U1211 (N_1211,N_935,N_716);
or U1212 (N_1212,N_784,N_904);
and U1213 (N_1213,N_745,N_653);
xnor U1214 (N_1214,N_804,N_945);
and U1215 (N_1215,N_523,N_846);
and U1216 (N_1216,N_943,N_921);
nand U1217 (N_1217,N_944,N_533);
nor U1218 (N_1218,N_772,N_906);
and U1219 (N_1219,N_622,N_693);
or U1220 (N_1220,N_735,N_707);
nor U1221 (N_1221,N_627,N_571);
nor U1222 (N_1222,N_631,N_594);
and U1223 (N_1223,N_842,N_692);
nand U1224 (N_1224,N_694,N_517);
or U1225 (N_1225,N_914,N_762);
nand U1226 (N_1226,N_848,N_837);
or U1227 (N_1227,N_773,N_820);
and U1228 (N_1228,N_637,N_683);
or U1229 (N_1229,N_998,N_539);
xor U1230 (N_1230,N_764,N_612);
and U1231 (N_1231,N_652,N_786);
nand U1232 (N_1232,N_830,N_674);
and U1233 (N_1233,N_736,N_509);
and U1234 (N_1234,N_985,N_512);
nor U1235 (N_1235,N_971,N_663);
nor U1236 (N_1236,N_885,N_619);
xnor U1237 (N_1237,N_959,N_771);
nor U1238 (N_1238,N_711,N_584);
xnor U1239 (N_1239,N_887,N_507);
xnor U1240 (N_1240,N_978,N_973);
nand U1241 (N_1241,N_751,N_709);
or U1242 (N_1242,N_974,N_760);
nor U1243 (N_1243,N_553,N_688);
and U1244 (N_1244,N_737,N_870);
xnor U1245 (N_1245,N_624,N_872);
or U1246 (N_1246,N_852,N_763);
nor U1247 (N_1247,N_742,N_937);
nor U1248 (N_1248,N_628,N_616);
xnor U1249 (N_1249,N_952,N_900);
xnor U1250 (N_1250,N_753,N_585);
or U1251 (N_1251,N_831,N_834);
nand U1252 (N_1252,N_787,N_514);
nor U1253 (N_1253,N_877,N_636);
nand U1254 (N_1254,N_623,N_705);
or U1255 (N_1255,N_884,N_752);
xnor U1256 (N_1256,N_706,N_935);
and U1257 (N_1257,N_640,N_850);
and U1258 (N_1258,N_774,N_720);
nor U1259 (N_1259,N_556,N_804);
and U1260 (N_1260,N_747,N_770);
and U1261 (N_1261,N_595,N_972);
nor U1262 (N_1262,N_834,N_826);
or U1263 (N_1263,N_504,N_891);
nor U1264 (N_1264,N_618,N_942);
xnor U1265 (N_1265,N_898,N_831);
and U1266 (N_1266,N_590,N_585);
nand U1267 (N_1267,N_707,N_792);
or U1268 (N_1268,N_758,N_635);
and U1269 (N_1269,N_834,N_630);
xor U1270 (N_1270,N_695,N_868);
or U1271 (N_1271,N_513,N_905);
xor U1272 (N_1272,N_682,N_726);
nor U1273 (N_1273,N_560,N_720);
nand U1274 (N_1274,N_617,N_518);
or U1275 (N_1275,N_649,N_905);
nor U1276 (N_1276,N_954,N_730);
and U1277 (N_1277,N_950,N_861);
nor U1278 (N_1278,N_826,N_552);
and U1279 (N_1279,N_599,N_832);
nor U1280 (N_1280,N_812,N_614);
nand U1281 (N_1281,N_686,N_976);
and U1282 (N_1282,N_756,N_949);
nor U1283 (N_1283,N_979,N_542);
nor U1284 (N_1284,N_733,N_805);
nand U1285 (N_1285,N_744,N_845);
nand U1286 (N_1286,N_723,N_651);
and U1287 (N_1287,N_716,N_968);
nand U1288 (N_1288,N_679,N_782);
and U1289 (N_1289,N_929,N_610);
nor U1290 (N_1290,N_939,N_830);
and U1291 (N_1291,N_834,N_668);
or U1292 (N_1292,N_904,N_645);
xor U1293 (N_1293,N_508,N_532);
or U1294 (N_1294,N_546,N_690);
nor U1295 (N_1295,N_694,N_810);
nor U1296 (N_1296,N_805,N_537);
nor U1297 (N_1297,N_667,N_734);
nand U1298 (N_1298,N_750,N_717);
nor U1299 (N_1299,N_994,N_525);
nand U1300 (N_1300,N_714,N_554);
and U1301 (N_1301,N_821,N_755);
and U1302 (N_1302,N_506,N_993);
nor U1303 (N_1303,N_645,N_734);
or U1304 (N_1304,N_777,N_853);
or U1305 (N_1305,N_760,N_766);
and U1306 (N_1306,N_889,N_549);
and U1307 (N_1307,N_765,N_681);
xor U1308 (N_1308,N_696,N_654);
or U1309 (N_1309,N_923,N_588);
or U1310 (N_1310,N_769,N_837);
nor U1311 (N_1311,N_602,N_622);
nand U1312 (N_1312,N_999,N_893);
nor U1313 (N_1313,N_627,N_881);
xor U1314 (N_1314,N_542,N_575);
nor U1315 (N_1315,N_816,N_676);
nand U1316 (N_1316,N_968,N_622);
or U1317 (N_1317,N_603,N_650);
xor U1318 (N_1318,N_888,N_893);
and U1319 (N_1319,N_694,N_944);
or U1320 (N_1320,N_918,N_976);
nand U1321 (N_1321,N_981,N_646);
nor U1322 (N_1322,N_856,N_942);
nand U1323 (N_1323,N_679,N_924);
and U1324 (N_1324,N_893,N_800);
and U1325 (N_1325,N_997,N_866);
nand U1326 (N_1326,N_981,N_782);
or U1327 (N_1327,N_995,N_820);
nor U1328 (N_1328,N_938,N_680);
or U1329 (N_1329,N_675,N_550);
and U1330 (N_1330,N_593,N_847);
nor U1331 (N_1331,N_989,N_768);
nor U1332 (N_1332,N_559,N_631);
or U1333 (N_1333,N_923,N_806);
nand U1334 (N_1334,N_596,N_930);
and U1335 (N_1335,N_978,N_511);
and U1336 (N_1336,N_731,N_804);
nand U1337 (N_1337,N_740,N_630);
or U1338 (N_1338,N_569,N_675);
and U1339 (N_1339,N_794,N_971);
or U1340 (N_1340,N_553,N_921);
or U1341 (N_1341,N_800,N_753);
nand U1342 (N_1342,N_705,N_884);
nand U1343 (N_1343,N_605,N_603);
and U1344 (N_1344,N_900,N_760);
or U1345 (N_1345,N_733,N_892);
nand U1346 (N_1346,N_910,N_646);
xor U1347 (N_1347,N_874,N_832);
nand U1348 (N_1348,N_533,N_901);
nor U1349 (N_1349,N_556,N_828);
nand U1350 (N_1350,N_877,N_674);
and U1351 (N_1351,N_702,N_538);
and U1352 (N_1352,N_772,N_764);
and U1353 (N_1353,N_984,N_876);
nor U1354 (N_1354,N_655,N_622);
or U1355 (N_1355,N_632,N_582);
nand U1356 (N_1356,N_805,N_758);
nor U1357 (N_1357,N_665,N_670);
nand U1358 (N_1358,N_846,N_985);
or U1359 (N_1359,N_809,N_524);
or U1360 (N_1360,N_843,N_576);
xor U1361 (N_1361,N_881,N_709);
and U1362 (N_1362,N_552,N_739);
xnor U1363 (N_1363,N_581,N_976);
nand U1364 (N_1364,N_616,N_552);
or U1365 (N_1365,N_833,N_693);
nand U1366 (N_1366,N_510,N_643);
nand U1367 (N_1367,N_991,N_810);
nand U1368 (N_1368,N_728,N_798);
nor U1369 (N_1369,N_672,N_704);
or U1370 (N_1370,N_771,N_547);
and U1371 (N_1371,N_914,N_792);
nand U1372 (N_1372,N_670,N_552);
nor U1373 (N_1373,N_589,N_981);
or U1374 (N_1374,N_775,N_789);
nor U1375 (N_1375,N_730,N_634);
and U1376 (N_1376,N_899,N_676);
or U1377 (N_1377,N_872,N_826);
nor U1378 (N_1378,N_839,N_620);
and U1379 (N_1379,N_713,N_653);
nand U1380 (N_1380,N_650,N_894);
and U1381 (N_1381,N_891,N_797);
or U1382 (N_1382,N_751,N_797);
xor U1383 (N_1383,N_532,N_513);
and U1384 (N_1384,N_849,N_747);
nand U1385 (N_1385,N_557,N_967);
xnor U1386 (N_1386,N_626,N_947);
nor U1387 (N_1387,N_670,N_694);
or U1388 (N_1388,N_740,N_530);
nand U1389 (N_1389,N_723,N_676);
nor U1390 (N_1390,N_941,N_916);
and U1391 (N_1391,N_672,N_562);
and U1392 (N_1392,N_584,N_936);
nand U1393 (N_1393,N_704,N_793);
nor U1394 (N_1394,N_965,N_854);
or U1395 (N_1395,N_908,N_598);
nand U1396 (N_1396,N_772,N_733);
or U1397 (N_1397,N_635,N_750);
or U1398 (N_1398,N_521,N_515);
nor U1399 (N_1399,N_746,N_535);
and U1400 (N_1400,N_608,N_775);
and U1401 (N_1401,N_546,N_952);
nor U1402 (N_1402,N_985,N_607);
or U1403 (N_1403,N_984,N_764);
or U1404 (N_1404,N_648,N_707);
and U1405 (N_1405,N_680,N_757);
nor U1406 (N_1406,N_559,N_757);
and U1407 (N_1407,N_639,N_566);
and U1408 (N_1408,N_936,N_925);
nor U1409 (N_1409,N_932,N_882);
and U1410 (N_1410,N_925,N_921);
and U1411 (N_1411,N_620,N_547);
nand U1412 (N_1412,N_615,N_588);
and U1413 (N_1413,N_528,N_506);
nand U1414 (N_1414,N_810,N_520);
nor U1415 (N_1415,N_740,N_889);
nor U1416 (N_1416,N_688,N_884);
and U1417 (N_1417,N_628,N_970);
nor U1418 (N_1418,N_520,N_554);
or U1419 (N_1419,N_689,N_655);
nor U1420 (N_1420,N_990,N_998);
nor U1421 (N_1421,N_953,N_883);
or U1422 (N_1422,N_520,N_883);
and U1423 (N_1423,N_761,N_523);
nand U1424 (N_1424,N_684,N_503);
nor U1425 (N_1425,N_838,N_759);
nor U1426 (N_1426,N_662,N_913);
and U1427 (N_1427,N_555,N_854);
or U1428 (N_1428,N_841,N_572);
and U1429 (N_1429,N_658,N_684);
nand U1430 (N_1430,N_987,N_796);
or U1431 (N_1431,N_586,N_706);
nand U1432 (N_1432,N_588,N_782);
nand U1433 (N_1433,N_904,N_746);
nor U1434 (N_1434,N_690,N_687);
xnor U1435 (N_1435,N_992,N_503);
and U1436 (N_1436,N_958,N_909);
nand U1437 (N_1437,N_981,N_884);
and U1438 (N_1438,N_922,N_879);
or U1439 (N_1439,N_584,N_681);
or U1440 (N_1440,N_828,N_775);
xnor U1441 (N_1441,N_893,N_990);
xnor U1442 (N_1442,N_815,N_554);
and U1443 (N_1443,N_673,N_736);
and U1444 (N_1444,N_950,N_786);
or U1445 (N_1445,N_582,N_927);
nand U1446 (N_1446,N_827,N_826);
nand U1447 (N_1447,N_745,N_970);
or U1448 (N_1448,N_991,N_608);
xor U1449 (N_1449,N_659,N_747);
and U1450 (N_1450,N_880,N_635);
and U1451 (N_1451,N_713,N_686);
and U1452 (N_1452,N_849,N_841);
nand U1453 (N_1453,N_552,N_856);
and U1454 (N_1454,N_722,N_646);
nand U1455 (N_1455,N_658,N_548);
and U1456 (N_1456,N_961,N_829);
nor U1457 (N_1457,N_554,N_587);
xnor U1458 (N_1458,N_732,N_999);
nor U1459 (N_1459,N_847,N_987);
nand U1460 (N_1460,N_714,N_641);
or U1461 (N_1461,N_541,N_505);
nor U1462 (N_1462,N_588,N_771);
nand U1463 (N_1463,N_540,N_611);
nand U1464 (N_1464,N_576,N_638);
nor U1465 (N_1465,N_727,N_594);
nor U1466 (N_1466,N_751,N_838);
nand U1467 (N_1467,N_524,N_811);
nor U1468 (N_1468,N_695,N_646);
nor U1469 (N_1469,N_542,N_620);
or U1470 (N_1470,N_950,N_737);
or U1471 (N_1471,N_710,N_775);
and U1472 (N_1472,N_706,N_750);
or U1473 (N_1473,N_989,N_987);
nand U1474 (N_1474,N_889,N_714);
and U1475 (N_1475,N_689,N_814);
xnor U1476 (N_1476,N_711,N_563);
nor U1477 (N_1477,N_951,N_927);
nor U1478 (N_1478,N_765,N_555);
nor U1479 (N_1479,N_977,N_721);
nand U1480 (N_1480,N_975,N_604);
xor U1481 (N_1481,N_956,N_770);
nor U1482 (N_1482,N_849,N_921);
xnor U1483 (N_1483,N_770,N_825);
nand U1484 (N_1484,N_920,N_592);
and U1485 (N_1485,N_675,N_866);
xor U1486 (N_1486,N_702,N_841);
and U1487 (N_1487,N_777,N_504);
xor U1488 (N_1488,N_782,N_612);
nor U1489 (N_1489,N_841,N_637);
nand U1490 (N_1490,N_994,N_964);
nand U1491 (N_1491,N_581,N_808);
and U1492 (N_1492,N_924,N_822);
nor U1493 (N_1493,N_710,N_556);
and U1494 (N_1494,N_817,N_606);
and U1495 (N_1495,N_588,N_847);
nor U1496 (N_1496,N_639,N_622);
or U1497 (N_1497,N_659,N_878);
nand U1498 (N_1498,N_960,N_528);
and U1499 (N_1499,N_716,N_863);
nor U1500 (N_1500,N_1376,N_1365);
and U1501 (N_1501,N_1048,N_1317);
nor U1502 (N_1502,N_1435,N_1203);
nand U1503 (N_1503,N_1320,N_1343);
nor U1504 (N_1504,N_1225,N_1424);
and U1505 (N_1505,N_1447,N_1255);
xor U1506 (N_1506,N_1165,N_1257);
nand U1507 (N_1507,N_1064,N_1101);
nor U1508 (N_1508,N_1332,N_1175);
and U1509 (N_1509,N_1252,N_1199);
and U1510 (N_1510,N_1303,N_1398);
nor U1511 (N_1511,N_1227,N_1336);
or U1512 (N_1512,N_1053,N_1393);
and U1513 (N_1513,N_1406,N_1243);
and U1514 (N_1514,N_1049,N_1330);
xnor U1515 (N_1515,N_1129,N_1143);
and U1516 (N_1516,N_1479,N_1246);
or U1517 (N_1517,N_1400,N_1170);
nor U1518 (N_1518,N_1464,N_1296);
and U1519 (N_1519,N_1042,N_1200);
or U1520 (N_1520,N_1459,N_1073);
nand U1521 (N_1521,N_1329,N_1472);
nand U1522 (N_1522,N_1190,N_1024);
or U1523 (N_1523,N_1371,N_1453);
nand U1524 (N_1524,N_1160,N_1044);
nand U1525 (N_1525,N_1364,N_1440);
nor U1526 (N_1526,N_1331,N_1071);
or U1527 (N_1527,N_1055,N_1110);
nor U1528 (N_1528,N_1058,N_1282);
nor U1529 (N_1529,N_1210,N_1146);
nor U1530 (N_1530,N_1347,N_1293);
nand U1531 (N_1531,N_1063,N_1346);
nor U1532 (N_1532,N_1433,N_1120);
nor U1533 (N_1533,N_1272,N_1294);
nand U1534 (N_1534,N_1168,N_1208);
or U1535 (N_1535,N_1380,N_1095);
and U1536 (N_1536,N_1133,N_1216);
nor U1537 (N_1537,N_1370,N_1138);
and U1538 (N_1538,N_1496,N_1494);
xor U1539 (N_1539,N_1311,N_1434);
nand U1540 (N_1540,N_1491,N_1323);
nor U1541 (N_1541,N_1070,N_1167);
nand U1542 (N_1542,N_1213,N_1467);
nand U1543 (N_1543,N_1345,N_1201);
or U1544 (N_1544,N_1418,N_1035);
and U1545 (N_1545,N_1209,N_1454);
nor U1546 (N_1546,N_1244,N_1162);
nand U1547 (N_1547,N_1436,N_1391);
and U1548 (N_1548,N_1384,N_1461);
and U1549 (N_1549,N_1358,N_1124);
xnor U1550 (N_1550,N_1137,N_1083);
and U1551 (N_1551,N_1261,N_1313);
nand U1552 (N_1552,N_1100,N_1022);
nand U1553 (N_1553,N_1362,N_1423);
nand U1554 (N_1554,N_1181,N_1113);
nor U1555 (N_1555,N_1369,N_1250);
or U1556 (N_1556,N_1289,N_1020);
nand U1557 (N_1557,N_1169,N_1401);
nor U1558 (N_1558,N_1003,N_1005);
or U1559 (N_1559,N_1059,N_1354);
or U1560 (N_1560,N_1164,N_1262);
nand U1561 (N_1561,N_1037,N_1182);
and U1562 (N_1562,N_1316,N_1019);
and U1563 (N_1563,N_1488,N_1002);
and U1564 (N_1564,N_1414,N_1215);
or U1565 (N_1565,N_1153,N_1135);
nor U1566 (N_1566,N_1178,N_1279);
xnor U1567 (N_1567,N_1211,N_1089);
or U1568 (N_1568,N_1076,N_1228);
xnor U1569 (N_1569,N_1388,N_1273);
nor U1570 (N_1570,N_1079,N_1399);
nand U1571 (N_1571,N_1307,N_1416);
nand U1572 (N_1572,N_1412,N_1457);
nor U1573 (N_1573,N_1127,N_1402);
nand U1574 (N_1574,N_1297,N_1087);
xor U1575 (N_1575,N_1150,N_1237);
nor U1576 (N_1576,N_1102,N_1154);
or U1577 (N_1577,N_1134,N_1045);
nor U1578 (N_1578,N_1098,N_1016);
and U1579 (N_1579,N_1093,N_1309);
nor U1580 (N_1580,N_1470,N_1231);
and U1581 (N_1581,N_1158,N_1027);
and U1582 (N_1582,N_1342,N_1419);
and U1583 (N_1583,N_1367,N_1455);
or U1584 (N_1584,N_1431,N_1439);
or U1585 (N_1585,N_1305,N_1015);
nor U1586 (N_1586,N_1196,N_1310);
nor U1587 (N_1587,N_1374,N_1094);
or U1588 (N_1588,N_1258,N_1214);
nor U1589 (N_1589,N_1006,N_1166);
nand U1590 (N_1590,N_1148,N_1284);
nor U1591 (N_1591,N_1333,N_1013);
nor U1592 (N_1592,N_1359,N_1281);
nand U1593 (N_1593,N_1119,N_1446);
or U1594 (N_1594,N_1217,N_1179);
or U1595 (N_1595,N_1482,N_1242);
nor U1596 (N_1596,N_1408,N_1264);
or U1597 (N_1597,N_1476,N_1449);
nand U1598 (N_1598,N_1223,N_1066);
or U1599 (N_1599,N_1067,N_1263);
nand U1600 (N_1600,N_1394,N_1009);
xor U1601 (N_1601,N_1497,N_1247);
nand U1602 (N_1602,N_1368,N_1465);
or U1603 (N_1603,N_1385,N_1381);
nand U1604 (N_1604,N_1256,N_1484);
nor U1605 (N_1605,N_1032,N_1108);
nor U1606 (N_1606,N_1474,N_1004);
or U1607 (N_1607,N_1239,N_1437);
xnor U1608 (N_1608,N_1144,N_1448);
or U1609 (N_1609,N_1241,N_1157);
nand U1610 (N_1610,N_1292,N_1460);
or U1611 (N_1611,N_1428,N_1269);
nor U1612 (N_1612,N_1340,N_1417);
nor U1613 (N_1613,N_1018,N_1413);
nand U1614 (N_1614,N_1145,N_1373);
or U1615 (N_1615,N_1286,N_1421);
and U1616 (N_1616,N_1238,N_1017);
nor U1617 (N_1617,N_1014,N_1130);
and U1618 (N_1618,N_1151,N_1056);
xor U1619 (N_1619,N_1462,N_1205);
nor U1620 (N_1620,N_1051,N_1366);
nand U1621 (N_1621,N_1288,N_1147);
nor U1622 (N_1622,N_1312,N_1357);
nand U1623 (N_1623,N_1389,N_1031);
and U1624 (N_1624,N_1084,N_1029);
nor U1625 (N_1625,N_1236,N_1010);
or U1626 (N_1626,N_1001,N_1325);
nand U1627 (N_1627,N_1041,N_1403);
nor U1628 (N_1628,N_1287,N_1328);
and U1629 (N_1629,N_1277,N_1422);
and U1630 (N_1630,N_1081,N_1266);
nor U1631 (N_1631,N_1226,N_1099);
nand U1632 (N_1632,N_1473,N_1061);
or U1633 (N_1633,N_1283,N_1046);
or U1634 (N_1634,N_1280,N_1379);
and U1635 (N_1635,N_1234,N_1180);
nor U1636 (N_1636,N_1382,N_1298);
nor U1637 (N_1637,N_1337,N_1097);
nor U1638 (N_1638,N_1060,N_1030);
or U1639 (N_1639,N_1039,N_1232);
nor U1640 (N_1640,N_1353,N_1132);
nand U1641 (N_1641,N_1189,N_1350);
xnor U1642 (N_1642,N_1360,N_1410);
nor U1643 (N_1643,N_1278,N_1253);
nand U1644 (N_1644,N_1112,N_1349);
nor U1645 (N_1645,N_1352,N_1334);
nand U1646 (N_1646,N_1355,N_1427);
xnor U1647 (N_1647,N_1128,N_1052);
and U1648 (N_1648,N_1174,N_1008);
nor U1649 (N_1649,N_1485,N_1483);
and U1650 (N_1650,N_1198,N_1319);
xor U1651 (N_1651,N_1078,N_1088);
and U1652 (N_1652,N_1033,N_1220);
nor U1653 (N_1653,N_1351,N_1072);
nor U1654 (N_1654,N_1490,N_1458);
and U1655 (N_1655,N_1300,N_1304);
or U1656 (N_1656,N_1397,N_1314);
nor U1657 (N_1657,N_1411,N_1092);
and U1658 (N_1658,N_1259,N_1091);
and U1659 (N_1659,N_1426,N_1396);
and U1660 (N_1660,N_1390,N_1121);
nor U1661 (N_1661,N_1085,N_1106);
and U1662 (N_1662,N_1194,N_1173);
nand U1663 (N_1663,N_1021,N_1131);
nand U1664 (N_1664,N_1191,N_1152);
nor U1665 (N_1665,N_1090,N_1140);
nand U1666 (N_1666,N_1276,N_1224);
nand U1667 (N_1667,N_1268,N_1271);
or U1668 (N_1668,N_1486,N_1267);
and U1669 (N_1669,N_1341,N_1075);
or U1670 (N_1670,N_1062,N_1193);
nand U1671 (N_1671,N_1235,N_1065);
or U1672 (N_1672,N_1468,N_1222);
and U1673 (N_1673,N_1372,N_1429);
or U1674 (N_1674,N_1012,N_1007);
nor U1675 (N_1675,N_1477,N_1043);
nor U1676 (N_1676,N_1103,N_1326);
or U1677 (N_1677,N_1197,N_1432);
or U1678 (N_1678,N_1047,N_1176);
or U1679 (N_1679,N_1469,N_1318);
nand U1680 (N_1680,N_1383,N_1187);
xnor U1681 (N_1681,N_1363,N_1080);
xor U1682 (N_1682,N_1077,N_1425);
and U1683 (N_1683,N_1212,N_1274);
xnor U1684 (N_1684,N_1285,N_1492);
and U1685 (N_1685,N_1348,N_1438);
and U1686 (N_1686,N_1171,N_1322);
and U1687 (N_1687,N_1295,N_1495);
or U1688 (N_1688,N_1395,N_1245);
or U1689 (N_1689,N_1186,N_1475);
nand U1690 (N_1690,N_1386,N_1034);
and U1691 (N_1691,N_1221,N_1463);
and U1692 (N_1692,N_1117,N_1415);
or U1693 (N_1693,N_1159,N_1392);
nor U1694 (N_1694,N_1270,N_1344);
nand U1695 (N_1695,N_1096,N_1183);
nor U1696 (N_1696,N_1115,N_1229);
xor U1697 (N_1697,N_1338,N_1142);
nand U1698 (N_1698,N_1141,N_1233);
nand U1699 (N_1699,N_1188,N_1441);
xnor U1700 (N_1700,N_1161,N_1387);
and U1701 (N_1701,N_1306,N_1456);
and U1702 (N_1702,N_1251,N_1026);
and U1703 (N_1703,N_1038,N_1123);
nor U1704 (N_1704,N_1445,N_1156);
nor U1705 (N_1705,N_1054,N_1487);
nand U1706 (N_1706,N_1324,N_1050);
nor U1707 (N_1707,N_1471,N_1248);
and U1708 (N_1708,N_1025,N_1126);
nand U1709 (N_1709,N_1116,N_1155);
nor U1710 (N_1710,N_1105,N_1011);
nor U1711 (N_1711,N_1184,N_1265);
and U1712 (N_1712,N_1204,N_1260);
or U1713 (N_1713,N_1122,N_1202);
nand U1714 (N_1714,N_1040,N_1420);
xor U1715 (N_1715,N_1498,N_1430);
xor U1716 (N_1716,N_1407,N_1206);
nor U1717 (N_1717,N_1109,N_1139);
and U1718 (N_1718,N_1450,N_1082);
and U1719 (N_1719,N_1442,N_1111);
nor U1720 (N_1720,N_1361,N_1335);
and U1721 (N_1721,N_1028,N_1192);
nor U1722 (N_1722,N_1023,N_1356);
and U1723 (N_1723,N_1339,N_1321);
and U1724 (N_1724,N_1219,N_1290);
xnor U1725 (N_1725,N_1404,N_1493);
or U1726 (N_1726,N_1409,N_1302);
nand U1727 (N_1727,N_1378,N_1249);
nor U1728 (N_1728,N_1185,N_1195);
and U1729 (N_1729,N_1375,N_1086);
nand U1730 (N_1730,N_1114,N_1481);
xnor U1731 (N_1731,N_1136,N_1478);
or U1732 (N_1732,N_1069,N_1068);
nand U1733 (N_1733,N_1036,N_1149);
and U1734 (N_1734,N_1489,N_1377);
nand U1735 (N_1735,N_1172,N_1451);
nand U1736 (N_1736,N_1308,N_1466);
nor U1737 (N_1737,N_1275,N_1444);
nor U1738 (N_1738,N_1207,N_1074);
or U1739 (N_1739,N_1315,N_1163);
nor U1740 (N_1740,N_1177,N_1301);
or U1741 (N_1741,N_1107,N_1405);
xnor U1742 (N_1742,N_1057,N_1104);
xor U1743 (N_1743,N_1218,N_1291);
xor U1744 (N_1744,N_1240,N_1125);
nand U1745 (N_1745,N_1443,N_1299);
or U1746 (N_1746,N_1480,N_1118);
nor U1747 (N_1747,N_1254,N_1000);
nand U1748 (N_1748,N_1230,N_1499);
and U1749 (N_1749,N_1452,N_1327);
nor U1750 (N_1750,N_1200,N_1049);
and U1751 (N_1751,N_1447,N_1221);
nor U1752 (N_1752,N_1172,N_1082);
xor U1753 (N_1753,N_1072,N_1049);
and U1754 (N_1754,N_1377,N_1234);
nor U1755 (N_1755,N_1124,N_1417);
and U1756 (N_1756,N_1270,N_1457);
or U1757 (N_1757,N_1236,N_1020);
or U1758 (N_1758,N_1224,N_1320);
and U1759 (N_1759,N_1036,N_1366);
nand U1760 (N_1760,N_1361,N_1190);
or U1761 (N_1761,N_1456,N_1191);
nand U1762 (N_1762,N_1194,N_1232);
and U1763 (N_1763,N_1279,N_1157);
and U1764 (N_1764,N_1457,N_1092);
and U1765 (N_1765,N_1389,N_1220);
and U1766 (N_1766,N_1137,N_1400);
nand U1767 (N_1767,N_1053,N_1084);
and U1768 (N_1768,N_1054,N_1474);
nor U1769 (N_1769,N_1094,N_1288);
nand U1770 (N_1770,N_1159,N_1226);
and U1771 (N_1771,N_1450,N_1290);
or U1772 (N_1772,N_1372,N_1463);
nor U1773 (N_1773,N_1441,N_1156);
nor U1774 (N_1774,N_1245,N_1253);
or U1775 (N_1775,N_1444,N_1372);
nor U1776 (N_1776,N_1472,N_1181);
nand U1777 (N_1777,N_1219,N_1047);
xnor U1778 (N_1778,N_1359,N_1415);
nor U1779 (N_1779,N_1032,N_1196);
xor U1780 (N_1780,N_1496,N_1073);
xnor U1781 (N_1781,N_1316,N_1148);
or U1782 (N_1782,N_1283,N_1112);
or U1783 (N_1783,N_1480,N_1422);
and U1784 (N_1784,N_1242,N_1279);
nand U1785 (N_1785,N_1027,N_1048);
nor U1786 (N_1786,N_1328,N_1254);
or U1787 (N_1787,N_1035,N_1264);
nand U1788 (N_1788,N_1180,N_1226);
and U1789 (N_1789,N_1450,N_1042);
nor U1790 (N_1790,N_1428,N_1330);
nand U1791 (N_1791,N_1126,N_1184);
xor U1792 (N_1792,N_1433,N_1225);
nand U1793 (N_1793,N_1421,N_1019);
nor U1794 (N_1794,N_1381,N_1354);
or U1795 (N_1795,N_1016,N_1469);
and U1796 (N_1796,N_1453,N_1129);
and U1797 (N_1797,N_1396,N_1383);
xnor U1798 (N_1798,N_1039,N_1027);
or U1799 (N_1799,N_1429,N_1027);
or U1800 (N_1800,N_1052,N_1163);
nand U1801 (N_1801,N_1471,N_1469);
or U1802 (N_1802,N_1339,N_1088);
and U1803 (N_1803,N_1209,N_1468);
and U1804 (N_1804,N_1406,N_1423);
nor U1805 (N_1805,N_1240,N_1295);
nand U1806 (N_1806,N_1425,N_1177);
nand U1807 (N_1807,N_1144,N_1174);
and U1808 (N_1808,N_1309,N_1005);
nor U1809 (N_1809,N_1080,N_1219);
nor U1810 (N_1810,N_1306,N_1322);
or U1811 (N_1811,N_1394,N_1279);
or U1812 (N_1812,N_1445,N_1253);
or U1813 (N_1813,N_1286,N_1397);
and U1814 (N_1814,N_1403,N_1498);
nor U1815 (N_1815,N_1120,N_1390);
and U1816 (N_1816,N_1277,N_1197);
or U1817 (N_1817,N_1103,N_1428);
and U1818 (N_1818,N_1399,N_1498);
nand U1819 (N_1819,N_1137,N_1495);
xnor U1820 (N_1820,N_1068,N_1201);
nand U1821 (N_1821,N_1496,N_1139);
nand U1822 (N_1822,N_1280,N_1397);
and U1823 (N_1823,N_1240,N_1458);
xor U1824 (N_1824,N_1059,N_1010);
or U1825 (N_1825,N_1247,N_1428);
nor U1826 (N_1826,N_1125,N_1365);
and U1827 (N_1827,N_1086,N_1232);
nor U1828 (N_1828,N_1142,N_1042);
and U1829 (N_1829,N_1456,N_1089);
nand U1830 (N_1830,N_1004,N_1109);
nor U1831 (N_1831,N_1115,N_1059);
and U1832 (N_1832,N_1070,N_1201);
or U1833 (N_1833,N_1380,N_1201);
nand U1834 (N_1834,N_1182,N_1121);
or U1835 (N_1835,N_1459,N_1313);
and U1836 (N_1836,N_1264,N_1050);
or U1837 (N_1837,N_1118,N_1368);
nor U1838 (N_1838,N_1429,N_1031);
nor U1839 (N_1839,N_1378,N_1401);
and U1840 (N_1840,N_1110,N_1024);
and U1841 (N_1841,N_1251,N_1440);
nand U1842 (N_1842,N_1422,N_1316);
xnor U1843 (N_1843,N_1357,N_1164);
and U1844 (N_1844,N_1238,N_1495);
nand U1845 (N_1845,N_1444,N_1083);
nor U1846 (N_1846,N_1318,N_1060);
or U1847 (N_1847,N_1019,N_1494);
nor U1848 (N_1848,N_1214,N_1431);
nand U1849 (N_1849,N_1073,N_1343);
or U1850 (N_1850,N_1159,N_1345);
or U1851 (N_1851,N_1181,N_1358);
nand U1852 (N_1852,N_1122,N_1091);
or U1853 (N_1853,N_1157,N_1284);
and U1854 (N_1854,N_1175,N_1302);
nor U1855 (N_1855,N_1302,N_1083);
nand U1856 (N_1856,N_1459,N_1053);
and U1857 (N_1857,N_1347,N_1117);
nand U1858 (N_1858,N_1232,N_1373);
or U1859 (N_1859,N_1456,N_1235);
or U1860 (N_1860,N_1370,N_1262);
or U1861 (N_1861,N_1447,N_1000);
nor U1862 (N_1862,N_1366,N_1237);
nor U1863 (N_1863,N_1059,N_1382);
nor U1864 (N_1864,N_1141,N_1098);
and U1865 (N_1865,N_1122,N_1268);
or U1866 (N_1866,N_1159,N_1026);
and U1867 (N_1867,N_1070,N_1120);
or U1868 (N_1868,N_1002,N_1192);
or U1869 (N_1869,N_1014,N_1196);
nand U1870 (N_1870,N_1337,N_1154);
nand U1871 (N_1871,N_1197,N_1101);
and U1872 (N_1872,N_1182,N_1375);
and U1873 (N_1873,N_1202,N_1406);
nor U1874 (N_1874,N_1386,N_1006);
nor U1875 (N_1875,N_1162,N_1212);
or U1876 (N_1876,N_1045,N_1005);
nand U1877 (N_1877,N_1348,N_1384);
nand U1878 (N_1878,N_1471,N_1080);
nor U1879 (N_1879,N_1123,N_1048);
nand U1880 (N_1880,N_1216,N_1459);
nand U1881 (N_1881,N_1327,N_1238);
or U1882 (N_1882,N_1171,N_1497);
nand U1883 (N_1883,N_1335,N_1302);
nand U1884 (N_1884,N_1198,N_1168);
nand U1885 (N_1885,N_1212,N_1456);
and U1886 (N_1886,N_1168,N_1179);
nand U1887 (N_1887,N_1153,N_1431);
nand U1888 (N_1888,N_1365,N_1308);
nor U1889 (N_1889,N_1320,N_1466);
nand U1890 (N_1890,N_1105,N_1080);
nor U1891 (N_1891,N_1307,N_1363);
xor U1892 (N_1892,N_1036,N_1164);
nor U1893 (N_1893,N_1160,N_1398);
and U1894 (N_1894,N_1157,N_1360);
and U1895 (N_1895,N_1310,N_1104);
nand U1896 (N_1896,N_1380,N_1291);
nor U1897 (N_1897,N_1261,N_1371);
and U1898 (N_1898,N_1194,N_1258);
nand U1899 (N_1899,N_1303,N_1377);
xor U1900 (N_1900,N_1422,N_1392);
nor U1901 (N_1901,N_1127,N_1102);
nand U1902 (N_1902,N_1176,N_1125);
nor U1903 (N_1903,N_1230,N_1317);
and U1904 (N_1904,N_1166,N_1454);
nor U1905 (N_1905,N_1482,N_1132);
nand U1906 (N_1906,N_1469,N_1295);
and U1907 (N_1907,N_1129,N_1447);
or U1908 (N_1908,N_1287,N_1285);
xor U1909 (N_1909,N_1176,N_1038);
xor U1910 (N_1910,N_1235,N_1239);
and U1911 (N_1911,N_1469,N_1365);
and U1912 (N_1912,N_1142,N_1476);
nor U1913 (N_1913,N_1181,N_1084);
nand U1914 (N_1914,N_1253,N_1459);
or U1915 (N_1915,N_1304,N_1274);
and U1916 (N_1916,N_1240,N_1362);
or U1917 (N_1917,N_1288,N_1133);
and U1918 (N_1918,N_1286,N_1237);
and U1919 (N_1919,N_1390,N_1426);
nand U1920 (N_1920,N_1071,N_1201);
nand U1921 (N_1921,N_1011,N_1098);
or U1922 (N_1922,N_1433,N_1488);
nor U1923 (N_1923,N_1075,N_1020);
xnor U1924 (N_1924,N_1416,N_1294);
nor U1925 (N_1925,N_1173,N_1147);
and U1926 (N_1926,N_1373,N_1070);
nor U1927 (N_1927,N_1026,N_1229);
nand U1928 (N_1928,N_1063,N_1321);
nor U1929 (N_1929,N_1066,N_1327);
nor U1930 (N_1930,N_1463,N_1423);
or U1931 (N_1931,N_1396,N_1074);
nand U1932 (N_1932,N_1128,N_1235);
nand U1933 (N_1933,N_1040,N_1352);
xnor U1934 (N_1934,N_1076,N_1022);
and U1935 (N_1935,N_1491,N_1179);
nor U1936 (N_1936,N_1257,N_1357);
nand U1937 (N_1937,N_1418,N_1047);
nand U1938 (N_1938,N_1033,N_1317);
xnor U1939 (N_1939,N_1448,N_1010);
nor U1940 (N_1940,N_1434,N_1484);
nor U1941 (N_1941,N_1260,N_1201);
nand U1942 (N_1942,N_1086,N_1038);
nor U1943 (N_1943,N_1285,N_1134);
or U1944 (N_1944,N_1249,N_1459);
or U1945 (N_1945,N_1002,N_1070);
nand U1946 (N_1946,N_1070,N_1006);
and U1947 (N_1947,N_1022,N_1063);
and U1948 (N_1948,N_1041,N_1420);
nor U1949 (N_1949,N_1260,N_1332);
or U1950 (N_1950,N_1463,N_1269);
nand U1951 (N_1951,N_1119,N_1262);
or U1952 (N_1952,N_1313,N_1052);
nand U1953 (N_1953,N_1310,N_1345);
and U1954 (N_1954,N_1268,N_1446);
and U1955 (N_1955,N_1343,N_1120);
and U1956 (N_1956,N_1326,N_1115);
xnor U1957 (N_1957,N_1196,N_1103);
or U1958 (N_1958,N_1211,N_1435);
or U1959 (N_1959,N_1361,N_1152);
nand U1960 (N_1960,N_1221,N_1444);
xnor U1961 (N_1961,N_1218,N_1066);
nand U1962 (N_1962,N_1261,N_1005);
xnor U1963 (N_1963,N_1096,N_1254);
nand U1964 (N_1964,N_1099,N_1371);
nand U1965 (N_1965,N_1325,N_1383);
nand U1966 (N_1966,N_1301,N_1058);
and U1967 (N_1967,N_1267,N_1413);
xnor U1968 (N_1968,N_1489,N_1315);
nor U1969 (N_1969,N_1496,N_1174);
nor U1970 (N_1970,N_1403,N_1341);
or U1971 (N_1971,N_1028,N_1460);
nor U1972 (N_1972,N_1080,N_1305);
nor U1973 (N_1973,N_1240,N_1449);
nor U1974 (N_1974,N_1111,N_1254);
or U1975 (N_1975,N_1164,N_1483);
xor U1976 (N_1976,N_1264,N_1387);
xnor U1977 (N_1977,N_1387,N_1422);
nand U1978 (N_1978,N_1051,N_1142);
and U1979 (N_1979,N_1355,N_1253);
nand U1980 (N_1980,N_1435,N_1065);
xor U1981 (N_1981,N_1177,N_1075);
and U1982 (N_1982,N_1073,N_1267);
nand U1983 (N_1983,N_1322,N_1173);
or U1984 (N_1984,N_1484,N_1495);
nor U1985 (N_1985,N_1271,N_1425);
or U1986 (N_1986,N_1133,N_1426);
and U1987 (N_1987,N_1225,N_1407);
nor U1988 (N_1988,N_1066,N_1183);
xnor U1989 (N_1989,N_1125,N_1154);
or U1990 (N_1990,N_1200,N_1448);
and U1991 (N_1991,N_1448,N_1373);
nor U1992 (N_1992,N_1285,N_1345);
and U1993 (N_1993,N_1192,N_1152);
and U1994 (N_1994,N_1080,N_1496);
and U1995 (N_1995,N_1278,N_1072);
nand U1996 (N_1996,N_1007,N_1140);
or U1997 (N_1997,N_1398,N_1497);
or U1998 (N_1998,N_1339,N_1276);
and U1999 (N_1999,N_1398,N_1093);
nand U2000 (N_2000,N_1583,N_1812);
nor U2001 (N_2001,N_1937,N_1848);
xor U2002 (N_2002,N_1602,N_1729);
nand U2003 (N_2003,N_1934,N_1961);
nand U2004 (N_2004,N_1738,N_1927);
or U2005 (N_2005,N_1733,N_1632);
nand U2006 (N_2006,N_1702,N_1629);
nand U2007 (N_2007,N_1554,N_1687);
and U2008 (N_2008,N_1813,N_1655);
nor U2009 (N_2009,N_1557,N_1933);
xnor U2010 (N_2010,N_1590,N_1775);
nand U2011 (N_2011,N_1841,N_1668);
nor U2012 (N_2012,N_1845,N_1849);
and U2013 (N_2013,N_1788,N_1571);
nor U2014 (N_2014,N_1858,N_1640);
nand U2015 (N_2015,N_1534,N_1781);
nand U2016 (N_2016,N_1824,N_1711);
or U2017 (N_2017,N_1965,N_1521);
xor U2018 (N_2018,N_1890,N_1635);
nor U2019 (N_2019,N_1701,N_1610);
nor U2020 (N_2020,N_1783,N_1770);
nor U2021 (N_2021,N_1815,N_1984);
nor U2022 (N_2022,N_1892,N_1740);
or U2023 (N_2023,N_1794,N_1593);
nor U2024 (N_2024,N_1985,N_1952);
and U2025 (N_2025,N_1761,N_1680);
xnor U2026 (N_2026,N_1630,N_1878);
or U2027 (N_2027,N_1966,N_1540);
and U2028 (N_2028,N_1539,N_1808);
nor U2029 (N_2029,N_1888,N_1889);
nand U2030 (N_2030,N_1504,N_1564);
and U2031 (N_2031,N_1737,N_1930);
and U2032 (N_2032,N_1720,N_1672);
and U2033 (N_2033,N_1653,N_1774);
and U2034 (N_2034,N_1975,N_1697);
nand U2035 (N_2035,N_1957,N_1713);
nand U2036 (N_2036,N_1634,N_1716);
or U2037 (N_2037,N_1580,N_1923);
nand U2038 (N_2038,N_1605,N_1698);
nand U2039 (N_2039,N_1928,N_1636);
nand U2040 (N_2040,N_1842,N_1659);
nor U2041 (N_2041,N_1859,N_1932);
and U2042 (N_2042,N_1675,N_1512);
or U2043 (N_2043,N_1947,N_1862);
xnor U2044 (N_2044,N_1663,N_1976);
or U2045 (N_2045,N_1501,N_1851);
and U2046 (N_2046,N_1739,N_1596);
nand U2047 (N_2047,N_1613,N_1936);
xnor U2048 (N_2048,N_1891,N_1728);
nor U2049 (N_2049,N_1818,N_1826);
nand U2050 (N_2050,N_1520,N_1718);
nor U2051 (N_2051,N_1692,N_1550);
nor U2052 (N_2052,N_1765,N_1832);
and U2053 (N_2053,N_1552,N_1569);
nor U2054 (N_2054,N_1676,N_1920);
nand U2055 (N_2055,N_1866,N_1855);
nor U2056 (N_2056,N_1657,N_1879);
nor U2057 (N_2057,N_1639,N_1938);
or U2058 (N_2058,N_1853,N_1750);
xor U2059 (N_2059,N_1523,N_1964);
or U2060 (N_2060,N_1903,N_1731);
or U2061 (N_2061,N_1695,N_1780);
xor U2062 (N_2062,N_1846,N_1727);
nor U2063 (N_2063,N_1665,N_1861);
xnor U2064 (N_2064,N_1648,N_1752);
nand U2065 (N_2065,N_1751,N_1766);
or U2066 (N_2066,N_1584,N_1837);
xor U2067 (N_2067,N_1784,N_1873);
and U2068 (N_2068,N_1608,N_1791);
nand U2069 (N_2069,N_1627,N_1746);
nor U2070 (N_2070,N_1979,N_1913);
or U2071 (N_2071,N_1943,N_1662);
nor U2072 (N_2072,N_1759,N_1717);
and U2073 (N_2073,N_1881,N_1545);
and U2074 (N_2074,N_1789,N_1960);
or U2075 (N_2075,N_1650,N_1631);
or U2076 (N_2076,N_1696,N_1921);
nand U2077 (N_2077,N_1978,N_1754);
nand U2078 (N_2078,N_1962,N_1516);
nor U2079 (N_2079,N_1642,N_1579);
nor U2080 (N_2080,N_1967,N_1758);
nand U2081 (N_2081,N_1707,N_1505);
and U2082 (N_2082,N_1940,N_1556);
and U2083 (N_2083,N_1773,N_1949);
and U2084 (N_2084,N_1973,N_1799);
nor U2085 (N_2085,N_1693,N_1527);
nand U2086 (N_2086,N_1797,N_1690);
nor U2087 (N_2087,N_1798,N_1868);
and U2088 (N_2088,N_1651,N_1756);
or U2089 (N_2089,N_1852,N_1532);
xor U2090 (N_2090,N_1743,N_1922);
nor U2091 (N_2091,N_1500,N_1721);
or U2092 (N_2092,N_1628,N_1897);
or U2093 (N_2093,N_1969,N_1679);
and U2094 (N_2094,N_1768,N_1677);
xor U2095 (N_2095,N_1656,N_1912);
nor U2096 (N_2096,N_1772,N_1604);
and U2097 (N_2097,N_1914,N_1518);
nand U2098 (N_2098,N_1997,N_1594);
and U2099 (N_2099,N_1524,N_1620);
nor U2100 (N_2100,N_1804,N_1712);
xnor U2101 (N_2101,N_1586,N_1622);
xor U2102 (N_2102,N_1592,N_1953);
nand U2103 (N_2103,N_1652,N_1819);
and U2104 (N_2104,N_1685,N_1863);
xor U2105 (N_2105,N_1730,N_1507);
and U2106 (N_2106,N_1896,N_1814);
and U2107 (N_2107,N_1694,N_1745);
and U2108 (N_2108,N_1736,N_1755);
xnor U2109 (N_2109,N_1753,N_1546);
or U2110 (N_2110,N_1547,N_1836);
nor U2111 (N_2111,N_1939,N_1839);
nand U2112 (N_2112,N_1795,N_1587);
nor U2113 (N_2113,N_1776,N_1537);
or U2114 (N_2114,N_1591,N_1983);
nor U2115 (N_2115,N_1667,N_1887);
or U2116 (N_2116,N_1948,N_1699);
nand U2117 (N_2117,N_1559,N_1802);
nand U2118 (N_2118,N_1638,N_1958);
nand U2119 (N_2119,N_1840,N_1529);
nand U2120 (N_2120,N_1519,N_1528);
or U2121 (N_2121,N_1654,N_1769);
nor U2122 (N_2122,N_1830,N_1792);
nand U2123 (N_2123,N_1671,N_1658);
nand U2124 (N_2124,N_1793,N_1709);
nand U2125 (N_2125,N_1637,N_1807);
nand U2126 (N_2126,N_1597,N_1993);
nor U2127 (N_2127,N_1601,N_1760);
nor U2128 (N_2128,N_1549,N_1996);
nor U2129 (N_2129,N_1644,N_1786);
and U2130 (N_2130,N_1778,N_1649);
nand U2131 (N_2131,N_1562,N_1906);
or U2132 (N_2132,N_1777,N_1573);
nor U2133 (N_2133,N_1909,N_1929);
nand U2134 (N_2134,N_1991,N_1683);
nand U2135 (N_2135,N_1763,N_1918);
xor U2136 (N_2136,N_1551,N_1682);
or U2137 (N_2137,N_1609,N_1911);
and U2138 (N_2138,N_1618,N_1522);
nand U2139 (N_2139,N_1904,N_1955);
nor U2140 (N_2140,N_1847,N_1850);
or U2141 (N_2141,N_1616,N_1843);
or U2142 (N_2142,N_1502,N_1875);
nor U2143 (N_2143,N_1872,N_1577);
and U2144 (N_2144,N_1894,N_1645);
nor U2145 (N_2145,N_1531,N_1735);
nor U2146 (N_2146,N_1764,N_1732);
and U2147 (N_2147,N_1741,N_1691);
nor U2148 (N_2148,N_1612,N_1542);
and U2149 (N_2149,N_1902,N_1581);
nor U2150 (N_2150,N_1661,N_1869);
nand U2151 (N_2151,N_1595,N_1538);
or U2152 (N_2152,N_1660,N_1822);
or U2153 (N_2153,N_1633,N_1681);
xor U2154 (N_2154,N_1901,N_1876);
nand U2155 (N_2155,N_1974,N_1941);
or U2156 (N_2156,N_1615,N_1995);
nor U2157 (N_2157,N_1684,N_1576);
and U2158 (N_2158,N_1990,N_1611);
nor U2159 (N_2159,N_1907,N_1513);
xor U2160 (N_2160,N_1899,N_1705);
nand U2161 (N_2161,N_1543,N_1726);
and U2162 (N_2162,N_1544,N_1910);
nand U2163 (N_2163,N_1871,N_1561);
or U2164 (N_2164,N_1885,N_1915);
nor U2165 (N_2165,N_1510,N_1771);
xnor U2166 (N_2166,N_1567,N_1865);
nand U2167 (N_2167,N_1833,N_1674);
or U2168 (N_2168,N_1686,N_1509);
nand U2169 (N_2169,N_1508,N_1882);
nand U2170 (N_2170,N_1560,N_1511);
or U2171 (N_2171,N_1688,N_1607);
nand U2172 (N_2172,N_1796,N_1575);
or U2173 (N_2173,N_1817,N_1874);
and U2174 (N_2174,N_1809,N_1748);
and U2175 (N_2175,N_1989,N_1762);
and U2176 (N_2176,N_1998,N_1582);
or U2177 (N_2177,N_1719,N_1884);
and U2178 (N_2178,N_1898,N_1744);
and U2179 (N_2179,N_1747,N_1810);
or U2180 (N_2180,N_1787,N_1666);
nand U2181 (N_2181,N_1572,N_1599);
nor U2182 (N_2182,N_1536,N_1782);
nor U2183 (N_2183,N_1623,N_1956);
and U2184 (N_2184,N_1968,N_1805);
or U2185 (N_2185,N_1844,N_1980);
or U2186 (N_2186,N_1823,N_1916);
nor U2187 (N_2187,N_1563,N_1785);
nor U2188 (N_2188,N_1829,N_1603);
nand U2189 (N_2189,N_1647,N_1908);
nor U2190 (N_2190,N_1870,N_1566);
nor U2191 (N_2191,N_1806,N_1749);
or U2192 (N_2192,N_1886,N_1570);
or U2193 (N_2193,N_1954,N_1625);
or U2194 (N_2194,N_1641,N_1919);
and U2195 (N_2195,N_1811,N_1526);
xnor U2196 (N_2196,N_1700,N_1517);
nor U2197 (N_2197,N_1803,N_1626);
nor U2198 (N_2198,N_1689,N_1959);
and U2199 (N_2199,N_1558,N_1568);
nor U2200 (N_2200,N_1506,N_1801);
xnor U2201 (N_2201,N_1742,N_1779);
or U2202 (N_2202,N_1703,N_1827);
or U2203 (N_2203,N_1854,N_1893);
nand U2204 (N_2204,N_1946,N_1828);
xor U2205 (N_2205,N_1515,N_1883);
and U2206 (N_2206,N_1838,N_1800);
and U2207 (N_2207,N_1617,N_1944);
nor U2208 (N_2208,N_1723,N_1619);
or U2209 (N_2209,N_1820,N_1734);
nand U2210 (N_2210,N_1670,N_1895);
nand U2211 (N_2211,N_1917,N_1541);
nand U2212 (N_2212,N_1673,N_1621);
nand U2213 (N_2213,N_1514,N_1790);
and U2214 (N_2214,N_1880,N_1646);
and U2215 (N_2215,N_1834,N_1994);
or U2216 (N_2216,N_1935,N_1643);
or U2217 (N_2217,N_1600,N_1715);
nor U2218 (N_2218,N_1767,N_1982);
and U2219 (N_2219,N_1664,N_1835);
and U2220 (N_2220,N_1963,N_1971);
or U2221 (N_2221,N_1905,N_1624);
nor U2222 (N_2222,N_1924,N_1831);
nand U2223 (N_2223,N_1588,N_1706);
nor U2224 (N_2224,N_1669,N_1951);
xnor U2225 (N_2225,N_1606,N_1589);
nor U2226 (N_2226,N_1999,N_1992);
xnor U2227 (N_2227,N_1942,N_1598);
nand U2228 (N_2228,N_1574,N_1704);
and U2229 (N_2229,N_1821,N_1578);
or U2230 (N_2230,N_1926,N_1988);
or U2231 (N_2231,N_1555,N_1825);
xor U2232 (N_2232,N_1931,N_1972);
nand U2233 (N_2233,N_1864,N_1678);
xnor U2234 (N_2234,N_1981,N_1977);
nor U2235 (N_2235,N_1710,N_1535);
and U2236 (N_2236,N_1925,N_1708);
and U2237 (N_2237,N_1987,N_1860);
nand U2238 (N_2238,N_1970,N_1986);
nor U2239 (N_2239,N_1877,N_1553);
nor U2240 (N_2240,N_1548,N_1867);
nand U2241 (N_2241,N_1530,N_1722);
and U2242 (N_2242,N_1525,N_1950);
and U2243 (N_2243,N_1533,N_1816);
or U2244 (N_2244,N_1900,N_1724);
nor U2245 (N_2245,N_1725,N_1945);
nand U2246 (N_2246,N_1565,N_1856);
or U2247 (N_2247,N_1857,N_1614);
nor U2248 (N_2248,N_1503,N_1585);
nor U2249 (N_2249,N_1714,N_1757);
and U2250 (N_2250,N_1510,N_1754);
nand U2251 (N_2251,N_1750,N_1882);
and U2252 (N_2252,N_1784,N_1705);
or U2253 (N_2253,N_1840,N_1660);
and U2254 (N_2254,N_1933,N_1651);
nand U2255 (N_2255,N_1580,N_1764);
or U2256 (N_2256,N_1720,N_1979);
and U2257 (N_2257,N_1560,N_1808);
or U2258 (N_2258,N_1854,N_1508);
and U2259 (N_2259,N_1946,N_1686);
or U2260 (N_2260,N_1959,N_1923);
nor U2261 (N_2261,N_1698,N_1941);
nand U2262 (N_2262,N_1809,N_1561);
and U2263 (N_2263,N_1529,N_1804);
and U2264 (N_2264,N_1662,N_1507);
or U2265 (N_2265,N_1593,N_1716);
nor U2266 (N_2266,N_1811,N_1897);
nor U2267 (N_2267,N_1900,N_1586);
nand U2268 (N_2268,N_1866,N_1967);
and U2269 (N_2269,N_1759,N_1734);
nor U2270 (N_2270,N_1739,N_1903);
nand U2271 (N_2271,N_1936,N_1535);
xnor U2272 (N_2272,N_1887,N_1506);
and U2273 (N_2273,N_1959,N_1756);
or U2274 (N_2274,N_1723,N_1841);
and U2275 (N_2275,N_1961,N_1896);
nor U2276 (N_2276,N_1974,N_1787);
nor U2277 (N_2277,N_1716,N_1515);
nor U2278 (N_2278,N_1922,N_1686);
or U2279 (N_2279,N_1810,N_1970);
or U2280 (N_2280,N_1892,N_1596);
or U2281 (N_2281,N_1806,N_1983);
and U2282 (N_2282,N_1863,N_1531);
nand U2283 (N_2283,N_1700,N_1649);
and U2284 (N_2284,N_1754,N_1823);
or U2285 (N_2285,N_1877,N_1952);
nand U2286 (N_2286,N_1882,N_1798);
and U2287 (N_2287,N_1954,N_1559);
or U2288 (N_2288,N_1632,N_1777);
xnor U2289 (N_2289,N_1994,N_1853);
nand U2290 (N_2290,N_1929,N_1518);
and U2291 (N_2291,N_1756,N_1518);
or U2292 (N_2292,N_1703,N_1734);
xor U2293 (N_2293,N_1979,N_1971);
and U2294 (N_2294,N_1533,N_1598);
nand U2295 (N_2295,N_1568,N_1817);
and U2296 (N_2296,N_1778,N_1764);
nor U2297 (N_2297,N_1869,N_1504);
nand U2298 (N_2298,N_1801,N_1748);
or U2299 (N_2299,N_1546,N_1639);
nor U2300 (N_2300,N_1884,N_1643);
and U2301 (N_2301,N_1928,N_1528);
nor U2302 (N_2302,N_1555,N_1912);
and U2303 (N_2303,N_1596,N_1803);
or U2304 (N_2304,N_1756,N_1957);
xnor U2305 (N_2305,N_1723,N_1708);
or U2306 (N_2306,N_1714,N_1742);
nand U2307 (N_2307,N_1833,N_1587);
and U2308 (N_2308,N_1565,N_1976);
nor U2309 (N_2309,N_1896,N_1760);
and U2310 (N_2310,N_1573,N_1627);
nor U2311 (N_2311,N_1514,N_1986);
xnor U2312 (N_2312,N_1521,N_1717);
or U2313 (N_2313,N_1539,N_1934);
or U2314 (N_2314,N_1703,N_1739);
or U2315 (N_2315,N_1976,N_1887);
and U2316 (N_2316,N_1900,N_1746);
nand U2317 (N_2317,N_1967,N_1566);
or U2318 (N_2318,N_1540,N_1826);
and U2319 (N_2319,N_1895,N_1896);
xnor U2320 (N_2320,N_1587,N_1630);
nand U2321 (N_2321,N_1672,N_1689);
and U2322 (N_2322,N_1750,N_1924);
or U2323 (N_2323,N_1767,N_1525);
nor U2324 (N_2324,N_1681,N_1760);
nand U2325 (N_2325,N_1690,N_1655);
nand U2326 (N_2326,N_1864,N_1846);
and U2327 (N_2327,N_1740,N_1858);
or U2328 (N_2328,N_1760,N_1572);
and U2329 (N_2329,N_1629,N_1822);
and U2330 (N_2330,N_1881,N_1920);
xnor U2331 (N_2331,N_1943,N_1843);
and U2332 (N_2332,N_1729,N_1798);
and U2333 (N_2333,N_1711,N_1538);
xnor U2334 (N_2334,N_1827,N_1837);
and U2335 (N_2335,N_1954,N_1787);
or U2336 (N_2336,N_1765,N_1667);
xnor U2337 (N_2337,N_1763,N_1863);
nand U2338 (N_2338,N_1952,N_1707);
nand U2339 (N_2339,N_1691,N_1752);
and U2340 (N_2340,N_1918,N_1743);
nand U2341 (N_2341,N_1613,N_1883);
and U2342 (N_2342,N_1894,N_1539);
nand U2343 (N_2343,N_1714,N_1940);
nor U2344 (N_2344,N_1930,N_1524);
nor U2345 (N_2345,N_1706,N_1978);
and U2346 (N_2346,N_1994,N_1902);
or U2347 (N_2347,N_1752,N_1878);
nand U2348 (N_2348,N_1992,N_1628);
and U2349 (N_2349,N_1836,N_1510);
or U2350 (N_2350,N_1922,N_1912);
or U2351 (N_2351,N_1595,N_1676);
nor U2352 (N_2352,N_1942,N_1790);
and U2353 (N_2353,N_1723,N_1964);
nor U2354 (N_2354,N_1613,N_1519);
nand U2355 (N_2355,N_1528,N_1759);
nand U2356 (N_2356,N_1617,N_1746);
nand U2357 (N_2357,N_1637,N_1828);
and U2358 (N_2358,N_1731,N_1778);
nand U2359 (N_2359,N_1612,N_1857);
nand U2360 (N_2360,N_1770,N_1645);
or U2361 (N_2361,N_1925,N_1886);
and U2362 (N_2362,N_1989,N_1689);
or U2363 (N_2363,N_1902,N_1701);
nand U2364 (N_2364,N_1929,N_1804);
xnor U2365 (N_2365,N_1576,N_1534);
and U2366 (N_2366,N_1583,N_1998);
and U2367 (N_2367,N_1734,N_1816);
and U2368 (N_2368,N_1783,N_1830);
nor U2369 (N_2369,N_1557,N_1966);
and U2370 (N_2370,N_1726,N_1643);
nor U2371 (N_2371,N_1865,N_1543);
and U2372 (N_2372,N_1722,N_1567);
nand U2373 (N_2373,N_1606,N_1626);
nand U2374 (N_2374,N_1670,N_1568);
or U2375 (N_2375,N_1739,N_1802);
nor U2376 (N_2376,N_1953,N_1920);
and U2377 (N_2377,N_1512,N_1822);
and U2378 (N_2378,N_1765,N_1986);
or U2379 (N_2379,N_1719,N_1564);
nand U2380 (N_2380,N_1594,N_1964);
xor U2381 (N_2381,N_1764,N_1879);
or U2382 (N_2382,N_1662,N_1925);
nor U2383 (N_2383,N_1726,N_1907);
nor U2384 (N_2384,N_1861,N_1783);
nor U2385 (N_2385,N_1667,N_1873);
nand U2386 (N_2386,N_1619,N_1932);
and U2387 (N_2387,N_1687,N_1638);
nor U2388 (N_2388,N_1759,N_1950);
or U2389 (N_2389,N_1763,N_1597);
nand U2390 (N_2390,N_1855,N_1858);
and U2391 (N_2391,N_1819,N_1687);
nor U2392 (N_2392,N_1506,N_1976);
nor U2393 (N_2393,N_1812,N_1669);
or U2394 (N_2394,N_1942,N_1503);
nor U2395 (N_2395,N_1637,N_1992);
nor U2396 (N_2396,N_1912,N_1810);
or U2397 (N_2397,N_1937,N_1906);
and U2398 (N_2398,N_1578,N_1702);
nand U2399 (N_2399,N_1685,N_1992);
nor U2400 (N_2400,N_1961,N_1531);
or U2401 (N_2401,N_1533,N_1806);
or U2402 (N_2402,N_1886,N_1500);
or U2403 (N_2403,N_1802,N_1754);
xor U2404 (N_2404,N_1689,N_1922);
xnor U2405 (N_2405,N_1752,N_1639);
and U2406 (N_2406,N_1609,N_1657);
nand U2407 (N_2407,N_1630,N_1891);
or U2408 (N_2408,N_1941,N_1891);
nor U2409 (N_2409,N_1942,N_1978);
nor U2410 (N_2410,N_1758,N_1962);
and U2411 (N_2411,N_1549,N_1535);
xnor U2412 (N_2412,N_1737,N_1665);
and U2413 (N_2413,N_1981,N_1582);
nand U2414 (N_2414,N_1821,N_1545);
nand U2415 (N_2415,N_1609,N_1827);
nor U2416 (N_2416,N_1895,N_1722);
nand U2417 (N_2417,N_1672,N_1515);
or U2418 (N_2418,N_1543,N_1546);
and U2419 (N_2419,N_1831,N_1565);
and U2420 (N_2420,N_1574,N_1874);
and U2421 (N_2421,N_1975,N_1625);
and U2422 (N_2422,N_1587,N_1505);
or U2423 (N_2423,N_1592,N_1686);
nand U2424 (N_2424,N_1809,N_1952);
xor U2425 (N_2425,N_1792,N_1834);
xor U2426 (N_2426,N_1559,N_1943);
and U2427 (N_2427,N_1915,N_1943);
and U2428 (N_2428,N_1565,N_1836);
nor U2429 (N_2429,N_1790,N_1537);
nor U2430 (N_2430,N_1854,N_1922);
or U2431 (N_2431,N_1825,N_1588);
nand U2432 (N_2432,N_1589,N_1920);
or U2433 (N_2433,N_1929,N_1989);
xnor U2434 (N_2434,N_1855,N_1807);
or U2435 (N_2435,N_1717,N_1708);
and U2436 (N_2436,N_1986,N_1791);
or U2437 (N_2437,N_1772,N_1992);
nor U2438 (N_2438,N_1647,N_1823);
nor U2439 (N_2439,N_1892,N_1641);
nor U2440 (N_2440,N_1746,N_1650);
nor U2441 (N_2441,N_1838,N_1978);
and U2442 (N_2442,N_1971,N_1840);
and U2443 (N_2443,N_1918,N_1606);
nor U2444 (N_2444,N_1646,N_1799);
nor U2445 (N_2445,N_1663,N_1515);
nor U2446 (N_2446,N_1510,N_1597);
nand U2447 (N_2447,N_1531,N_1733);
nor U2448 (N_2448,N_1995,N_1843);
and U2449 (N_2449,N_1811,N_1520);
nand U2450 (N_2450,N_1636,N_1904);
xor U2451 (N_2451,N_1738,N_1909);
or U2452 (N_2452,N_1533,N_1543);
nor U2453 (N_2453,N_1625,N_1881);
nor U2454 (N_2454,N_1773,N_1906);
and U2455 (N_2455,N_1806,N_1796);
nor U2456 (N_2456,N_1773,N_1663);
or U2457 (N_2457,N_1993,N_1536);
or U2458 (N_2458,N_1629,N_1808);
and U2459 (N_2459,N_1861,N_1920);
nand U2460 (N_2460,N_1559,N_1856);
nand U2461 (N_2461,N_1610,N_1695);
and U2462 (N_2462,N_1938,N_1740);
xor U2463 (N_2463,N_1522,N_1926);
nand U2464 (N_2464,N_1709,N_1528);
nand U2465 (N_2465,N_1862,N_1700);
xor U2466 (N_2466,N_1920,N_1600);
or U2467 (N_2467,N_1958,N_1676);
or U2468 (N_2468,N_1641,N_1682);
or U2469 (N_2469,N_1879,N_1902);
and U2470 (N_2470,N_1806,N_1693);
nand U2471 (N_2471,N_1875,N_1595);
or U2472 (N_2472,N_1699,N_1704);
and U2473 (N_2473,N_1569,N_1693);
nor U2474 (N_2474,N_1577,N_1888);
xor U2475 (N_2475,N_1988,N_1743);
or U2476 (N_2476,N_1618,N_1895);
or U2477 (N_2477,N_1866,N_1641);
nor U2478 (N_2478,N_1725,N_1957);
nand U2479 (N_2479,N_1596,N_1663);
and U2480 (N_2480,N_1896,N_1654);
nor U2481 (N_2481,N_1911,N_1516);
nor U2482 (N_2482,N_1585,N_1671);
xnor U2483 (N_2483,N_1565,N_1579);
nand U2484 (N_2484,N_1548,N_1683);
and U2485 (N_2485,N_1635,N_1540);
nor U2486 (N_2486,N_1669,N_1945);
nand U2487 (N_2487,N_1750,N_1629);
xnor U2488 (N_2488,N_1661,N_1984);
nand U2489 (N_2489,N_1931,N_1890);
nor U2490 (N_2490,N_1911,N_1779);
and U2491 (N_2491,N_1904,N_1512);
or U2492 (N_2492,N_1935,N_1705);
nand U2493 (N_2493,N_1949,N_1500);
and U2494 (N_2494,N_1987,N_1639);
and U2495 (N_2495,N_1518,N_1516);
nor U2496 (N_2496,N_1656,N_1658);
or U2497 (N_2497,N_1927,N_1737);
nand U2498 (N_2498,N_1650,N_1899);
and U2499 (N_2499,N_1520,N_1824);
xor U2500 (N_2500,N_2225,N_2217);
and U2501 (N_2501,N_2365,N_2362);
or U2502 (N_2502,N_2131,N_2441);
xnor U2503 (N_2503,N_2435,N_2292);
xor U2504 (N_2504,N_2282,N_2094);
nor U2505 (N_2505,N_2467,N_2159);
nor U2506 (N_2506,N_2246,N_2495);
nand U2507 (N_2507,N_2076,N_2029);
or U2508 (N_2508,N_2129,N_2251);
or U2509 (N_2509,N_2314,N_2095);
nor U2510 (N_2510,N_2455,N_2174);
nand U2511 (N_2511,N_2258,N_2078);
nand U2512 (N_2512,N_2419,N_2352);
nand U2513 (N_2513,N_2265,N_2142);
nor U2514 (N_2514,N_2428,N_2236);
and U2515 (N_2515,N_2433,N_2499);
or U2516 (N_2516,N_2297,N_2053);
nand U2517 (N_2517,N_2006,N_2107);
and U2518 (N_2518,N_2263,N_2026);
or U2519 (N_2519,N_2337,N_2137);
and U2520 (N_2520,N_2284,N_2481);
or U2521 (N_2521,N_2484,N_2064);
xnor U2522 (N_2522,N_2322,N_2100);
nor U2523 (N_2523,N_2390,N_2168);
or U2524 (N_2524,N_2332,N_2154);
and U2525 (N_2525,N_2418,N_2203);
nand U2526 (N_2526,N_2115,N_2187);
and U2527 (N_2527,N_2468,N_2404);
or U2528 (N_2528,N_2393,N_2194);
and U2529 (N_2529,N_2215,N_2123);
nand U2530 (N_2530,N_2234,N_2060);
xor U2531 (N_2531,N_2457,N_2066);
nand U2532 (N_2532,N_2102,N_2180);
or U2533 (N_2533,N_2077,N_2272);
and U2534 (N_2534,N_2268,N_2376);
nand U2535 (N_2535,N_2465,N_2036);
and U2536 (N_2536,N_2132,N_2039);
nor U2537 (N_2537,N_2092,N_2151);
nor U2538 (N_2538,N_2489,N_2114);
and U2539 (N_2539,N_2456,N_2400);
and U2540 (N_2540,N_2331,N_2323);
nor U2541 (N_2541,N_2289,N_2061);
nor U2542 (N_2542,N_2055,N_2235);
and U2543 (N_2543,N_2408,N_2392);
nor U2544 (N_2544,N_2196,N_2249);
nor U2545 (N_2545,N_2113,N_2188);
and U2546 (N_2546,N_2080,N_2072);
or U2547 (N_2547,N_2042,N_2295);
or U2548 (N_2548,N_2243,N_2030);
and U2549 (N_2549,N_2206,N_2473);
or U2550 (N_2550,N_2054,N_2377);
nor U2551 (N_2551,N_2202,N_2049);
or U2552 (N_2552,N_2069,N_2470);
nor U2553 (N_2553,N_2220,N_2333);
nor U2554 (N_2554,N_2436,N_2155);
nor U2555 (N_2555,N_2166,N_2124);
and U2556 (N_2556,N_2172,N_2306);
and U2557 (N_2557,N_2002,N_2296);
and U2558 (N_2558,N_2460,N_2007);
nand U2559 (N_2559,N_2287,N_2379);
nor U2560 (N_2560,N_2099,N_2093);
nor U2561 (N_2561,N_2381,N_2308);
or U2562 (N_2562,N_2126,N_2449);
xor U2563 (N_2563,N_2046,N_2452);
nand U2564 (N_2564,N_2320,N_2025);
nand U2565 (N_2565,N_2276,N_2480);
xor U2566 (N_2566,N_2299,N_2421);
nand U2567 (N_2567,N_2430,N_2406);
nor U2568 (N_2568,N_2440,N_2254);
or U2569 (N_2569,N_2367,N_2425);
and U2570 (N_2570,N_2471,N_2338);
nor U2571 (N_2571,N_2143,N_2157);
or U2572 (N_2572,N_2040,N_2253);
nand U2573 (N_2573,N_2027,N_2207);
nor U2574 (N_2574,N_2490,N_2056);
and U2575 (N_2575,N_2085,N_2405);
or U2576 (N_2576,N_2190,N_2363);
or U2577 (N_2577,N_2104,N_2271);
nor U2578 (N_2578,N_2375,N_2412);
nor U2579 (N_2579,N_2186,N_2402);
or U2580 (N_2580,N_2148,N_2205);
or U2581 (N_2581,N_2161,N_2339);
and U2582 (N_2582,N_2237,N_2310);
and U2583 (N_2583,N_2261,N_2313);
nor U2584 (N_2584,N_2398,N_2476);
or U2585 (N_2585,N_2149,N_2221);
and U2586 (N_2586,N_2138,N_2141);
and U2587 (N_2587,N_2275,N_2063);
nor U2588 (N_2588,N_2183,N_2201);
and U2589 (N_2589,N_2477,N_2073);
nor U2590 (N_2590,N_2209,N_2368);
or U2591 (N_2591,N_2252,N_2461);
or U2592 (N_2592,N_2448,N_2328);
and U2593 (N_2593,N_2110,N_2108);
and U2594 (N_2594,N_2396,N_2020);
nand U2595 (N_2595,N_2179,N_2475);
and U2596 (N_2596,N_2199,N_2173);
and U2597 (N_2597,N_2346,N_2387);
nand U2598 (N_2598,N_2413,N_2195);
nor U2599 (N_2599,N_2164,N_2324);
or U2600 (N_2600,N_2019,N_2382);
nor U2601 (N_2601,N_2079,N_2106);
or U2602 (N_2602,N_2302,N_2366);
xnor U2603 (N_2603,N_2045,N_2011);
nand U2604 (N_2604,N_2033,N_2169);
nand U2605 (N_2605,N_2062,N_2122);
nand U2606 (N_2606,N_2232,N_2226);
or U2607 (N_2607,N_2486,N_2058);
and U2608 (N_2608,N_2444,N_2277);
xor U2609 (N_2609,N_2311,N_2429);
nor U2610 (N_2610,N_2147,N_2176);
and U2611 (N_2611,N_2130,N_2270);
nor U2612 (N_2612,N_2008,N_2178);
xnor U2613 (N_2613,N_2315,N_2278);
nor U2614 (N_2614,N_2330,N_2358);
xor U2615 (N_2615,N_2407,N_2478);
nand U2616 (N_2616,N_2288,N_2443);
nor U2617 (N_2617,N_2422,N_2192);
and U2618 (N_2618,N_2083,N_2244);
nor U2619 (N_2619,N_2013,N_2394);
or U2620 (N_2620,N_2374,N_2482);
and U2621 (N_2621,N_2096,N_2032);
nor U2622 (N_2622,N_2321,N_2239);
or U2623 (N_2623,N_2351,N_2028);
and U2624 (N_2624,N_2373,N_2181);
nand U2625 (N_2625,N_2163,N_2015);
and U2626 (N_2626,N_2081,N_2487);
nor U2627 (N_2627,N_2498,N_2336);
and U2628 (N_2628,N_2070,N_2426);
and U2629 (N_2629,N_2128,N_2326);
nand U2630 (N_2630,N_2454,N_2485);
nand U2631 (N_2631,N_2453,N_2241);
and U2632 (N_2632,N_2293,N_2037);
nand U2633 (N_2633,N_2139,N_2091);
xnor U2634 (N_2634,N_2354,N_2193);
or U2635 (N_2635,N_2127,N_2259);
xnor U2636 (N_2636,N_2230,N_2052);
or U2637 (N_2637,N_2160,N_2103);
nor U2638 (N_2638,N_2000,N_2384);
or U2639 (N_2639,N_2197,N_2493);
or U2640 (N_2640,N_2135,N_2140);
or U2641 (N_2641,N_2458,N_2152);
nor U2642 (N_2642,N_2118,N_2432);
and U2643 (N_2643,N_2423,N_2101);
nor U2644 (N_2644,N_2090,N_2222);
and U2645 (N_2645,N_2247,N_2001);
nand U2646 (N_2646,N_2451,N_2316);
or U2647 (N_2647,N_2211,N_2109);
nor U2648 (N_2648,N_2041,N_2361);
nand U2649 (N_2649,N_2356,N_2388);
and U2650 (N_2650,N_2403,N_2309);
nor U2651 (N_2651,N_2009,N_2450);
and U2652 (N_2652,N_2372,N_2319);
nor U2653 (N_2653,N_2198,N_2410);
nand U2654 (N_2654,N_2117,N_2304);
and U2655 (N_2655,N_2255,N_2116);
and U2656 (N_2656,N_2047,N_2156);
or U2657 (N_2657,N_2350,N_2228);
nand U2658 (N_2658,N_2380,N_2213);
nand U2659 (N_2659,N_2262,N_2170);
or U2660 (N_2660,N_2158,N_2219);
nor U2661 (N_2661,N_2389,N_2134);
and U2662 (N_2662,N_2018,N_2105);
or U2663 (N_2663,N_2267,N_2023);
nand U2664 (N_2664,N_2245,N_2150);
and U2665 (N_2665,N_2329,N_2120);
nor U2666 (N_2666,N_2248,N_2301);
and U2667 (N_2667,N_2364,N_2399);
and U2668 (N_2668,N_2231,N_2048);
nor U2669 (N_2669,N_2347,N_2177);
and U2670 (N_2670,N_2401,N_2146);
nand U2671 (N_2671,N_2024,N_2153);
or U2672 (N_2672,N_2204,N_2307);
or U2673 (N_2673,N_2415,N_2281);
xor U2674 (N_2674,N_2012,N_2218);
nand U2675 (N_2675,N_2437,N_2464);
nor U2676 (N_2676,N_2459,N_2191);
and U2677 (N_2677,N_2463,N_2305);
xnor U2678 (N_2678,N_2411,N_2086);
nor U2679 (N_2679,N_2233,N_2466);
and U2680 (N_2680,N_2111,N_2447);
and U2681 (N_2681,N_2003,N_2479);
and U2682 (N_2682,N_2416,N_2355);
and U2683 (N_2683,N_2397,N_2185);
nor U2684 (N_2684,N_2483,N_2427);
and U2685 (N_2685,N_2335,N_2269);
nor U2686 (N_2686,N_2383,N_2439);
xor U2687 (N_2687,N_2385,N_2274);
or U2688 (N_2688,N_2214,N_2353);
or U2689 (N_2689,N_2189,N_2496);
nor U2690 (N_2690,N_2369,N_2256);
and U2691 (N_2691,N_2238,N_2260);
nand U2692 (N_2692,N_2184,N_2098);
xor U2693 (N_2693,N_2133,N_2162);
and U2694 (N_2694,N_2283,N_2016);
nand U2695 (N_2695,N_2395,N_2343);
nor U2696 (N_2696,N_2325,N_2165);
and U2697 (N_2697,N_2294,N_2212);
nand U2698 (N_2698,N_2065,N_2022);
and U2699 (N_2699,N_2462,N_2119);
and U2700 (N_2700,N_2059,N_2494);
xor U2701 (N_2701,N_2431,N_2434);
nor U2702 (N_2702,N_2031,N_2446);
nand U2703 (N_2703,N_2286,N_2112);
or U2704 (N_2704,N_2472,N_2442);
and U2705 (N_2705,N_2317,N_2175);
or U2706 (N_2706,N_2391,N_2171);
xor U2707 (N_2707,N_2264,N_2348);
xor U2708 (N_2708,N_2349,N_2144);
xnor U2709 (N_2709,N_2136,N_2227);
and U2710 (N_2710,N_2200,N_2327);
or U2711 (N_2711,N_2409,N_2334);
nor U2712 (N_2712,N_2474,N_2224);
xor U2713 (N_2713,N_2280,N_2082);
or U2714 (N_2714,N_2370,N_2378);
and U2715 (N_2715,N_2492,N_2341);
and U2716 (N_2716,N_2050,N_2125);
and U2717 (N_2717,N_2497,N_2257);
or U2718 (N_2718,N_2298,N_2071);
and U2719 (N_2719,N_2051,N_2145);
xnor U2720 (N_2720,N_2034,N_2291);
and U2721 (N_2721,N_2043,N_2121);
nand U2722 (N_2722,N_2074,N_2360);
nand U2723 (N_2723,N_2469,N_2182);
xor U2724 (N_2724,N_2216,N_2344);
or U2725 (N_2725,N_2240,N_2010);
and U2726 (N_2726,N_2057,N_2067);
nand U2727 (N_2727,N_2491,N_2250);
and U2728 (N_2728,N_2312,N_2273);
nand U2729 (N_2729,N_2229,N_2084);
or U2730 (N_2730,N_2285,N_2420);
xnor U2731 (N_2731,N_2424,N_2097);
xnor U2732 (N_2732,N_2021,N_2386);
xor U2733 (N_2733,N_2223,N_2068);
or U2734 (N_2734,N_2345,N_2303);
or U2735 (N_2735,N_2005,N_2445);
nand U2736 (N_2736,N_2087,N_2075);
nor U2737 (N_2737,N_2371,N_2014);
xnor U2738 (N_2738,N_2359,N_2279);
and U2739 (N_2739,N_2017,N_2290);
nand U2740 (N_2740,N_2438,N_2035);
xnor U2741 (N_2741,N_2242,N_2300);
or U2742 (N_2742,N_2044,N_2417);
or U2743 (N_2743,N_2167,N_2357);
xor U2744 (N_2744,N_2208,N_2342);
xor U2745 (N_2745,N_2004,N_2088);
and U2746 (N_2746,N_2210,N_2488);
and U2747 (N_2747,N_2089,N_2038);
and U2748 (N_2748,N_2340,N_2318);
nor U2749 (N_2749,N_2414,N_2266);
or U2750 (N_2750,N_2218,N_2185);
and U2751 (N_2751,N_2149,N_2344);
xor U2752 (N_2752,N_2313,N_2134);
and U2753 (N_2753,N_2163,N_2064);
nor U2754 (N_2754,N_2206,N_2492);
nor U2755 (N_2755,N_2366,N_2387);
nor U2756 (N_2756,N_2482,N_2137);
and U2757 (N_2757,N_2250,N_2067);
or U2758 (N_2758,N_2469,N_2419);
and U2759 (N_2759,N_2356,N_2024);
nor U2760 (N_2760,N_2497,N_2432);
nor U2761 (N_2761,N_2062,N_2143);
and U2762 (N_2762,N_2316,N_2386);
xnor U2763 (N_2763,N_2410,N_2420);
nor U2764 (N_2764,N_2148,N_2436);
xor U2765 (N_2765,N_2390,N_2019);
xnor U2766 (N_2766,N_2206,N_2104);
or U2767 (N_2767,N_2141,N_2336);
nand U2768 (N_2768,N_2083,N_2429);
or U2769 (N_2769,N_2343,N_2153);
and U2770 (N_2770,N_2190,N_2105);
or U2771 (N_2771,N_2233,N_2474);
or U2772 (N_2772,N_2302,N_2415);
and U2773 (N_2773,N_2191,N_2222);
xor U2774 (N_2774,N_2360,N_2034);
nand U2775 (N_2775,N_2075,N_2343);
xnor U2776 (N_2776,N_2001,N_2055);
and U2777 (N_2777,N_2025,N_2084);
or U2778 (N_2778,N_2438,N_2327);
or U2779 (N_2779,N_2198,N_2438);
xor U2780 (N_2780,N_2051,N_2485);
nand U2781 (N_2781,N_2044,N_2142);
nor U2782 (N_2782,N_2117,N_2146);
nand U2783 (N_2783,N_2130,N_2149);
xnor U2784 (N_2784,N_2164,N_2478);
or U2785 (N_2785,N_2039,N_2221);
and U2786 (N_2786,N_2411,N_2177);
nand U2787 (N_2787,N_2233,N_2281);
nand U2788 (N_2788,N_2097,N_2028);
nand U2789 (N_2789,N_2086,N_2360);
and U2790 (N_2790,N_2093,N_2367);
or U2791 (N_2791,N_2361,N_2105);
or U2792 (N_2792,N_2273,N_2180);
or U2793 (N_2793,N_2329,N_2109);
or U2794 (N_2794,N_2227,N_2470);
or U2795 (N_2795,N_2283,N_2407);
nand U2796 (N_2796,N_2175,N_2418);
or U2797 (N_2797,N_2026,N_2409);
nor U2798 (N_2798,N_2361,N_2320);
or U2799 (N_2799,N_2335,N_2097);
and U2800 (N_2800,N_2193,N_2110);
nand U2801 (N_2801,N_2155,N_2373);
nor U2802 (N_2802,N_2147,N_2327);
xnor U2803 (N_2803,N_2020,N_2328);
nand U2804 (N_2804,N_2340,N_2211);
or U2805 (N_2805,N_2332,N_2293);
and U2806 (N_2806,N_2253,N_2163);
nand U2807 (N_2807,N_2023,N_2107);
nor U2808 (N_2808,N_2031,N_2066);
nand U2809 (N_2809,N_2177,N_2434);
nor U2810 (N_2810,N_2383,N_2292);
or U2811 (N_2811,N_2310,N_2320);
nand U2812 (N_2812,N_2109,N_2186);
nand U2813 (N_2813,N_2293,N_2486);
nand U2814 (N_2814,N_2127,N_2278);
nand U2815 (N_2815,N_2028,N_2280);
nand U2816 (N_2816,N_2389,N_2333);
and U2817 (N_2817,N_2384,N_2092);
xor U2818 (N_2818,N_2451,N_2044);
or U2819 (N_2819,N_2192,N_2231);
or U2820 (N_2820,N_2102,N_2422);
and U2821 (N_2821,N_2236,N_2392);
xnor U2822 (N_2822,N_2278,N_2297);
or U2823 (N_2823,N_2428,N_2472);
nand U2824 (N_2824,N_2024,N_2125);
xnor U2825 (N_2825,N_2115,N_2338);
xnor U2826 (N_2826,N_2263,N_2039);
or U2827 (N_2827,N_2042,N_2029);
xnor U2828 (N_2828,N_2157,N_2206);
nor U2829 (N_2829,N_2308,N_2313);
nand U2830 (N_2830,N_2347,N_2324);
and U2831 (N_2831,N_2256,N_2099);
nor U2832 (N_2832,N_2497,N_2231);
nand U2833 (N_2833,N_2267,N_2394);
nand U2834 (N_2834,N_2138,N_2034);
or U2835 (N_2835,N_2389,N_2152);
nand U2836 (N_2836,N_2067,N_2025);
nand U2837 (N_2837,N_2193,N_2332);
nand U2838 (N_2838,N_2117,N_2481);
or U2839 (N_2839,N_2344,N_2146);
nor U2840 (N_2840,N_2438,N_2077);
or U2841 (N_2841,N_2130,N_2336);
xnor U2842 (N_2842,N_2241,N_2044);
and U2843 (N_2843,N_2461,N_2190);
and U2844 (N_2844,N_2016,N_2351);
and U2845 (N_2845,N_2357,N_2266);
nor U2846 (N_2846,N_2055,N_2461);
nor U2847 (N_2847,N_2347,N_2400);
nor U2848 (N_2848,N_2413,N_2142);
nand U2849 (N_2849,N_2094,N_2089);
or U2850 (N_2850,N_2496,N_2390);
and U2851 (N_2851,N_2144,N_2186);
nor U2852 (N_2852,N_2258,N_2123);
nand U2853 (N_2853,N_2439,N_2319);
xor U2854 (N_2854,N_2213,N_2410);
nor U2855 (N_2855,N_2053,N_2010);
and U2856 (N_2856,N_2138,N_2189);
nor U2857 (N_2857,N_2192,N_2218);
nor U2858 (N_2858,N_2147,N_2119);
and U2859 (N_2859,N_2330,N_2216);
xnor U2860 (N_2860,N_2408,N_2352);
and U2861 (N_2861,N_2025,N_2154);
xnor U2862 (N_2862,N_2288,N_2323);
and U2863 (N_2863,N_2163,N_2408);
and U2864 (N_2864,N_2334,N_2035);
nand U2865 (N_2865,N_2197,N_2186);
and U2866 (N_2866,N_2120,N_2029);
xor U2867 (N_2867,N_2384,N_2153);
or U2868 (N_2868,N_2442,N_2111);
xnor U2869 (N_2869,N_2009,N_2225);
and U2870 (N_2870,N_2420,N_2247);
and U2871 (N_2871,N_2082,N_2380);
nor U2872 (N_2872,N_2188,N_2467);
xnor U2873 (N_2873,N_2127,N_2250);
nor U2874 (N_2874,N_2092,N_2118);
and U2875 (N_2875,N_2167,N_2214);
and U2876 (N_2876,N_2056,N_2331);
nand U2877 (N_2877,N_2213,N_2220);
and U2878 (N_2878,N_2215,N_2446);
nor U2879 (N_2879,N_2415,N_2397);
or U2880 (N_2880,N_2153,N_2070);
nand U2881 (N_2881,N_2380,N_2498);
and U2882 (N_2882,N_2254,N_2323);
nor U2883 (N_2883,N_2488,N_2009);
nor U2884 (N_2884,N_2439,N_2179);
and U2885 (N_2885,N_2374,N_2444);
nand U2886 (N_2886,N_2140,N_2168);
nand U2887 (N_2887,N_2063,N_2144);
xor U2888 (N_2888,N_2297,N_2214);
or U2889 (N_2889,N_2122,N_2208);
and U2890 (N_2890,N_2351,N_2422);
xor U2891 (N_2891,N_2496,N_2354);
nor U2892 (N_2892,N_2442,N_2328);
nand U2893 (N_2893,N_2275,N_2084);
nor U2894 (N_2894,N_2066,N_2187);
nand U2895 (N_2895,N_2339,N_2235);
xnor U2896 (N_2896,N_2248,N_2015);
nor U2897 (N_2897,N_2475,N_2456);
or U2898 (N_2898,N_2173,N_2390);
xor U2899 (N_2899,N_2405,N_2038);
nor U2900 (N_2900,N_2013,N_2392);
or U2901 (N_2901,N_2321,N_2288);
nor U2902 (N_2902,N_2482,N_2268);
or U2903 (N_2903,N_2452,N_2443);
and U2904 (N_2904,N_2071,N_2093);
nand U2905 (N_2905,N_2184,N_2182);
xnor U2906 (N_2906,N_2093,N_2013);
nand U2907 (N_2907,N_2419,N_2493);
nand U2908 (N_2908,N_2136,N_2146);
or U2909 (N_2909,N_2484,N_2003);
and U2910 (N_2910,N_2262,N_2375);
or U2911 (N_2911,N_2385,N_2358);
or U2912 (N_2912,N_2192,N_2325);
nor U2913 (N_2913,N_2494,N_2372);
and U2914 (N_2914,N_2069,N_2209);
nand U2915 (N_2915,N_2072,N_2054);
or U2916 (N_2916,N_2468,N_2460);
nor U2917 (N_2917,N_2258,N_2044);
nand U2918 (N_2918,N_2351,N_2179);
nand U2919 (N_2919,N_2257,N_2448);
xor U2920 (N_2920,N_2141,N_2225);
or U2921 (N_2921,N_2089,N_2217);
or U2922 (N_2922,N_2315,N_2487);
and U2923 (N_2923,N_2100,N_2242);
or U2924 (N_2924,N_2080,N_2127);
or U2925 (N_2925,N_2354,N_2419);
or U2926 (N_2926,N_2445,N_2389);
nor U2927 (N_2927,N_2104,N_2098);
nand U2928 (N_2928,N_2460,N_2453);
nor U2929 (N_2929,N_2170,N_2451);
and U2930 (N_2930,N_2033,N_2097);
and U2931 (N_2931,N_2221,N_2202);
and U2932 (N_2932,N_2276,N_2201);
or U2933 (N_2933,N_2376,N_2154);
nor U2934 (N_2934,N_2118,N_2443);
nor U2935 (N_2935,N_2296,N_2325);
or U2936 (N_2936,N_2263,N_2021);
and U2937 (N_2937,N_2345,N_2482);
nand U2938 (N_2938,N_2430,N_2201);
or U2939 (N_2939,N_2012,N_2116);
nand U2940 (N_2940,N_2134,N_2402);
or U2941 (N_2941,N_2497,N_2453);
and U2942 (N_2942,N_2283,N_2124);
xnor U2943 (N_2943,N_2149,N_2010);
xnor U2944 (N_2944,N_2006,N_2314);
or U2945 (N_2945,N_2044,N_2435);
nor U2946 (N_2946,N_2266,N_2262);
nand U2947 (N_2947,N_2244,N_2405);
nor U2948 (N_2948,N_2234,N_2003);
or U2949 (N_2949,N_2265,N_2238);
or U2950 (N_2950,N_2105,N_2058);
xor U2951 (N_2951,N_2126,N_2313);
or U2952 (N_2952,N_2358,N_2333);
xor U2953 (N_2953,N_2211,N_2439);
and U2954 (N_2954,N_2165,N_2423);
and U2955 (N_2955,N_2361,N_2281);
nor U2956 (N_2956,N_2290,N_2457);
or U2957 (N_2957,N_2353,N_2037);
nor U2958 (N_2958,N_2255,N_2097);
nand U2959 (N_2959,N_2459,N_2290);
xnor U2960 (N_2960,N_2039,N_2169);
or U2961 (N_2961,N_2462,N_2281);
and U2962 (N_2962,N_2099,N_2049);
nand U2963 (N_2963,N_2223,N_2264);
or U2964 (N_2964,N_2392,N_2135);
or U2965 (N_2965,N_2466,N_2453);
or U2966 (N_2966,N_2186,N_2222);
nor U2967 (N_2967,N_2395,N_2263);
or U2968 (N_2968,N_2100,N_2354);
or U2969 (N_2969,N_2398,N_2081);
nor U2970 (N_2970,N_2272,N_2175);
nand U2971 (N_2971,N_2141,N_2169);
nor U2972 (N_2972,N_2045,N_2103);
nand U2973 (N_2973,N_2455,N_2358);
xor U2974 (N_2974,N_2435,N_2077);
and U2975 (N_2975,N_2436,N_2362);
xnor U2976 (N_2976,N_2442,N_2373);
or U2977 (N_2977,N_2425,N_2471);
nor U2978 (N_2978,N_2134,N_2046);
or U2979 (N_2979,N_2378,N_2130);
and U2980 (N_2980,N_2401,N_2069);
nand U2981 (N_2981,N_2472,N_2142);
and U2982 (N_2982,N_2481,N_2441);
and U2983 (N_2983,N_2142,N_2491);
and U2984 (N_2984,N_2036,N_2071);
and U2985 (N_2985,N_2157,N_2101);
and U2986 (N_2986,N_2409,N_2163);
and U2987 (N_2987,N_2425,N_2198);
or U2988 (N_2988,N_2249,N_2020);
and U2989 (N_2989,N_2034,N_2282);
and U2990 (N_2990,N_2265,N_2006);
or U2991 (N_2991,N_2265,N_2448);
nand U2992 (N_2992,N_2025,N_2272);
and U2993 (N_2993,N_2295,N_2014);
nor U2994 (N_2994,N_2075,N_2182);
and U2995 (N_2995,N_2231,N_2072);
and U2996 (N_2996,N_2420,N_2193);
and U2997 (N_2997,N_2498,N_2299);
xor U2998 (N_2998,N_2233,N_2212);
nand U2999 (N_2999,N_2104,N_2132);
and U3000 (N_3000,N_2893,N_2999);
nor U3001 (N_3001,N_2990,N_2816);
nor U3002 (N_3002,N_2536,N_2580);
or U3003 (N_3003,N_2672,N_2900);
nand U3004 (N_3004,N_2593,N_2813);
nand U3005 (N_3005,N_2909,N_2969);
nand U3006 (N_3006,N_2686,N_2815);
nand U3007 (N_3007,N_2948,N_2719);
or U3008 (N_3008,N_2917,N_2976);
nor U3009 (N_3009,N_2645,N_2992);
nor U3010 (N_3010,N_2818,N_2890);
xnor U3011 (N_3011,N_2944,N_2779);
or U3012 (N_3012,N_2766,N_2661);
nor U3013 (N_3013,N_2665,N_2675);
nor U3014 (N_3014,N_2799,N_2885);
nor U3015 (N_3015,N_2589,N_2736);
nor U3016 (N_3016,N_2571,N_2621);
xnor U3017 (N_3017,N_2983,N_2875);
and U3018 (N_3018,N_2648,N_2868);
nor U3019 (N_3019,N_2666,N_2787);
nand U3020 (N_3020,N_2817,N_2943);
and U3021 (N_3021,N_2535,N_2549);
nor U3022 (N_3022,N_2572,N_2634);
nor U3023 (N_3023,N_2507,N_2579);
and U3024 (N_3024,N_2761,N_2502);
and U3025 (N_3025,N_2737,N_2929);
xnor U3026 (N_3026,N_2640,N_2770);
and U3027 (N_3027,N_2691,N_2935);
nor U3028 (N_3028,N_2695,N_2716);
or U3029 (N_3029,N_2851,N_2807);
and U3030 (N_3030,N_2711,N_2925);
xnor U3031 (N_3031,N_2837,N_2653);
and U3032 (N_3032,N_2626,N_2870);
or U3033 (N_3033,N_2913,N_2866);
nor U3034 (N_3034,N_2606,N_2898);
or U3035 (N_3035,N_2590,N_2584);
xor U3036 (N_3036,N_2820,N_2783);
and U3037 (N_3037,N_2884,N_2897);
nor U3038 (N_3038,N_2708,N_2694);
nor U3039 (N_3039,N_2765,N_2906);
and U3040 (N_3040,N_2633,N_2703);
nand U3041 (N_3041,N_2771,N_2971);
nor U3042 (N_3042,N_2876,N_2618);
nand U3043 (N_3043,N_2947,N_2923);
or U3044 (N_3044,N_2528,N_2669);
xor U3045 (N_3045,N_2750,N_2790);
nand U3046 (N_3046,N_2822,N_2577);
and U3047 (N_3047,N_2836,N_2751);
and U3048 (N_3048,N_2553,N_2841);
and U3049 (N_3049,N_2855,N_2550);
and U3050 (N_3050,N_2699,N_2782);
nor U3051 (N_3051,N_2950,N_2762);
nand U3052 (N_3052,N_2594,N_2639);
and U3053 (N_3053,N_2683,N_2561);
or U3054 (N_3054,N_2786,N_2518);
nand U3055 (N_3055,N_2768,N_2792);
and U3056 (N_3056,N_2718,N_2916);
and U3057 (N_3057,N_2854,N_2838);
xor U3058 (N_3058,N_2834,N_2952);
or U3059 (N_3059,N_2982,N_2956);
nand U3060 (N_3060,N_2616,N_2509);
nand U3061 (N_3061,N_2702,N_2805);
nor U3062 (N_3062,N_2953,N_2714);
xnor U3063 (N_3063,N_2968,N_2674);
nand U3064 (N_3064,N_2595,N_2707);
nor U3065 (N_3065,N_2814,N_2505);
and U3066 (N_3066,N_2721,N_2617);
xor U3067 (N_3067,N_2588,N_2788);
nor U3068 (N_3068,N_2993,N_2551);
nand U3069 (N_3069,N_2903,N_2965);
nor U3070 (N_3070,N_2743,N_2628);
nand U3071 (N_3071,N_2659,N_2632);
nand U3072 (N_3072,N_2864,N_2717);
nor U3073 (N_3073,N_2696,N_2769);
and U3074 (N_3074,N_2775,N_2763);
or U3075 (N_3075,N_2915,N_2605);
or U3076 (N_3076,N_2733,N_2583);
and U3077 (N_3077,N_2684,N_2902);
nor U3078 (N_3078,N_2882,N_2501);
nand U3079 (N_3079,N_2731,N_2678);
nor U3080 (N_3080,N_2567,N_2725);
or U3081 (N_3081,N_2794,N_2531);
nor U3082 (N_3082,N_2773,N_2940);
or U3083 (N_3083,N_2552,N_2513);
or U3084 (N_3084,N_2701,N_2881);
and U3085 (N_3085,N_2798,N_2828);
or U3086 (N_3086,N_2564,N_2607);
xnor U3087 (N_3087,N_2514,N_2705);
nor U3088 (N_3088,N_2730,N_2521);
nand U3089 (N_3089,N_2647,N_2597);
nand U3090 (N_3090,N_2693,N_2789);
nor U3091 (N_3091,N_2918,N_2927);
and U3092 (N_3092,N_2544,N_2889);
and U3093 (N_3093,N_2877,N_2772);
nand U3094 (N_3094,N_2614,N_2734);
nor U3095 (N_3095,N_2748,N_2832);
and U3096 (N_3096,N_2957,N_2879);
and U3097 (N_3097,N_2986,N_2874);
nand U3098 (N_3098,N_2537,N_2596);
and U3099 (N_3099,N_2599,N_2939);
and U3100 (N_3100,N_2995,N_2987);
or U3101 (N_3101,N_2573,N_2526);
or U3102 (N_3102,N_2860,N_2586);
nor U3103 (N_3103,N_2955,N_2824);
or U3104 (N_3104,N_2777,N_2742);
nand U3105 (N_3105,N_2872,N_2997);
xnor U3106 (N_3106,N_2858,N_2920);
xor U3107 (N_3107,N_2755,N_2933);
nand U3108 (N_3108,N_2547,N_2942);
nand U3109 (N_3109,N_2585,N_2515);
nor U3110 (N_3110,N_2978,N_2891);
nand U3111 (N_3111,N_2587,N_2706);
nor U3112 (N_3112,N_2994,N_2778);
nor U3113 (N_3113,N_2859,N_2525);
nor U3114 (N_3114,N_2985,N_2801);
xnor U3115 (N_3115,N_2548,N_2687);
nand U3116 (N_3116,N_2975,N_2928);
nor U3117 (N_3117,N_2563,N_2895);
nor U3118 (N_3118,N_2979,N_2753);
nand U3119 (N_3119,N_2869,N_2738);
or U3120 (N_3120,N_2700,N_2519);
or U3121 (N_3121,N_2949,N_2689);
nor U3122 (N_3122,N_2578,N_2911);
and U3123 (N_3123,N_2624,N_2608);
nand U3124 (N_3124,N_2861,N_2932);
or U3125 (N_3125,N_2541,N_2892);
and U3126 (N_3126,N_2853,N_2631);
or U3127 (N_3127,N_2998,N_2727);
nand U3128 (N_3128,N_2615,N_2641);
nand U3129 (N_3129,N_2679,N_2862);
or U3130 (N_3130,N_2520,N_2803);
nor U3131 (N_3131,N_2811,N_2758);
xnor U3132 (N_3132,N_2936,N_2904);
nand U3133 (N_3133,N_2601,N_2697);
or U3134 (N_3134,N_2980,N_2937);
or U3135 (N_3135,N_2996,N_2619);
and U3136 (N_3136,N_2849,N_2649);
or U3137 (N_3137,N_2781,N_2873);
and U3138 (N_3138,N_2545,N_2517);
nand U3139 (N_3139,N_2611,N_2912);
nor U3140 (N_3140,N_2793,N_2625);
nor U3141 (N_3141,N_2991,N_2668);
xnor U3142 (N_3142,N_2559,N_2622);
nand U3143 (N_3143,N_2662,N_2774);
and U3144 (N_3144,N_2886,N_2646);
and U3145 (N_3145,N_2840,N_2746);
or U3146 (N_3146,N_2945,N_2581);
xnor U3147 (N_3147,N_2598,N_2565);
or U3148 (N_3148,N_2812,N_2575);
or U3149 (N_3149,N_2511,N_2627);
nor U3150 (N_3150,N_2557,N_2613);
nor U3151 (N_3151,N_2922,N_2726);
and U3152 (N_3152,N_2643,N_2780);
and U3153 (N_3153,N_2914,N_2764);
and U3154 (N_3154,N_2833,N_2845);
or U3155 (N_3155,N_2591,N_2776);
or U3156 (N_3156,N_2655,N_2685);
nor U3157 (N_3157,N_2800,N_2728);
or U3158 (N_3158,N_2852,N_2506);
or U3159 (N_3159,N_2558,N_2963);
nand U3160 (N_3160,N_2842,N_2974);
nor U3161 (N_3161,N_2908,N_2752);
nor U3162 (N_3162,N_2958,N_2620);
nor U3163 (N_3163,N_2523,N_2878);
or U3164 (N_3164,N_2988,N_2612);
nor U3165 (N_3165,N_2574,N_2830);
nand U3166 (N_3166,N_2809,N_2656);
and U3167 (N_3167,N_2880,N_2516);
nand U3168 (N_3168,N_2749,N_2568);
nand U3169 (N_3169,N_2522,N_2823);
nor U3170 (N_3170,N_2680,N_2871);
and U3171 (N_3171,N_2629,N_2977);
and U3172 (N_3172,N_2938,N_2715);
nor U3173 (N_3173,N_2538,N_2735);
nor U3174 (N_3174,N_2709,N_2970);
nand U3175 (N_3175,N_2887,N_2896);
or U3176 (N_3176,N_2796,N_2682);
and U3177 (N_3177,N_2543,N_2671);
and U3178 (N_3178,N_2961,N_2660);
nand U3179 (N_3179,N_2946,N_2821);
nand U3180 (N_3180,N_2905,N_2825);
or U3181 (N_3181,N_2797,N_2829);
nor U3182 (N_3182,N_2582,N_2767);
or U3183 (N_3183,N_2533,N_2635);
nor U3184 (N_3184,N_2981,N_2967);
nor U3185 (N_3185,N_2512,N_2973);
and U3186 (N_3186,N_2741,N_2754);
nor U3187 (N_3187,N_2642,N_2791);
or U3188 (N_3188,N_2802,N_2539);
and U3189 (N_3189,N_2542,N_2554);
nand U3190 (N_3190,N_2724,N_2835);
and U3191 (N_3191,N_2857,N_2592);
and U3192 (N_3192,N_2658,N_2951);
nand U3193 (N_3193,N_2710,N_2546);
and U3194 (N_3194,N_2560,N_2888);
nand U3195 (N_3195,N_2540,N_2704);
nor U3196 (N_3196,N_2910,N_2712);
nand U3197 (N_3197,N_2600,N_2610);
nor U3198 (N_3198,N_2722,N_2664);
nor U3199 (N_3199,N_2555,N_2739);
and U3200 (N_3200,N_2847,N_2637);
and U3201 (N_3201,N_2919,N_2907);
or U3202 (N_3202,N_2839,N_2785);
or U3203 (N_3203,N_2530,N_2819);
and U3204 (N_3204,N_2831,N_2894);
or U3205 (N_3205,N_2534,N_2856);
or U3206 (N_3206,N_2745,N_2865);
nand U3207 (N_3207,N_2690,N_2650);
nor U3208 (N_3208,N_2652,N_2759);
xnor U3209 (N_3209,N_2795,N_2934);
nor U3210 (N_3210,N_2504,N_2848);
and U3211 (N_3211,N_2972,N_2850);
nor U3212 (N_3212,N_2964,N_2732);
or U3213 (N_3213,N_2500,N_2954);
or U3214 (N_3214,N_2698,N_2931);
nor U3215 (N_3215,N_2930,N_2556);
and U3216 (N_3216,N_2744,N_2569);
or U3217 (N_3217,N_2503,N_2677);
or U3218 (N_3218,N_2688,N_2810);
or U3219 (N_3219,N_2959,N_2603);
or U3220 (N_3220,N_2576,N_2638);
or U3221 (N_3221,N_2989,N_2663);
nor U3222 (N_3222,N_2827,N_2508);
or U3223 (N_3223,N_2562,N_2676);
nand U3224 (N_3224,N_2670,N_2740);
nor U3225 (N_3225,N_2984,N_2604);
and U3226 (N_3226,N_2692,N_2899);
or U3227 (N_3227,N_2843,N_2926);
or U3228 (N_3228,N_2867,N_2651);
or U3229 (N_3229,N_2729,N_2527);
nand U3230 (N_3230,N_2673,N_2960);
nor U3231 (N_3231,N_2804,N_2756);
xnor U3232 (N_3232,N_2636,N_2570);
xor U3233 (N_3233,N_2623,N_2941);
nand U3234 (N_3234,N_2524,N_2808);
or U3235 (N_3235,N_2784,N_2962);
or U3236 (N_3236,N_2529,N_2644);
or U3237 (N_3237,N_2924,N_2806);
xnor U3238 (N_3238,N_2760,N_2901);
nor U3239 (N_3239,N_2846,N_2602);
xnor U3240 (N_3240,N_2966,N_2510);
nand U3241 (N_3241,N_2713,N_2609);
and U3242 (N_3242,N_2720,N_2667);
nor U3243 (N_3243,N_2681,N_2863);
nand U3244 (N_3244,N_2757,N_2723);
nand U3245 (N_3245,N_2532,N_2883);
nor U3246 (N_3246,N_2654,N_2657);
nor U3247 (N_3247,N_2921,N_2630);
or U3248 (N_3248,N_2844,N_2826);
nor U3249 (N_3249,N_2566,N_2747);
or U3250 (N_3250,N_2895,N_2634);
and U3251 (N_3251,N_2930,N_2717);
nor U3252 (N_3252,N_2704,N_2627);
nand U3253 (N_3253,N_2900,N_2994);
nand U3254 (N_3254,N_2877,N_2714);
nand U3255 (N_3255,N_2956,N_2960);
nand U3256 (N_3256,N_2666,N_2772);
or U3257 (N_3257,N_2742,N_2877);
nor U3258 (N_3258,N_2586,N_2542);
xor U3259 (N_3259,N_2552,N_2565);
and U3260 (N_3260,N_2801,N_2956);
nand U3261 (N_3261,N_2865,N_2628);
or U3262 (N_3262,N_2750,N_2947);
or U3263 (N_3263,N_2871,N_2715);
or U3264 (N_3264,N_2890,N_2569);
xnor U3265 (N_3265,N_2974,N_2985);
nand U3266 (N_3266,N_2883,N_2972);
or U3267 (N_3267,N_2962,N_2685);
nand U3268 (N_3268,N_2506,N_2574);
and U3269 (N_3269,N_2659,N_2826);
nand U3270 (N_3270,N_2739,N_2876);
and U3271 (N_3271,N_2799,N_2686);
or U3272 (N_3272,N_2666,N_2659);
nor U3273 (N_3273,N_2968,N_2860);
or U3274 (N_3274,N_2996,N_2872);
xor U3275 (N_3275,N_2953,N_2594);
and U3276 (N_3276,N_2748,N_2532);
or U3277 (N_3277,N_2678,N_2879);
nand U3278 (N_3278,N_2829,N_2672);
and U3279 (N_3279,N_2644,N_2980);
nand U3280 (N_3280,N_2646,N_2958);
nor U3281 (N_3281,N_2912,N_2680);
and U3282 (N_3282,N_2515,N_2790);
or U3283 (N_3283,N_2874,N_2588);
nand U3284 (N_3284,N_2669,N_2657);
xor U3285 (N_3285,N_2959,N_2534);
and U3286 (N_3286,N_2822,N_2681);
nand U3287 (N_3287,N_2668,N_2557);
or U3288 (N_3288,N_2760,N_2643);
nor U3289 (N_3289,N_2662,N_2715);
nand U3290 (N_3290,N_2585,N_2825);
nand U3291 (N_3291,N_2958,N_2863);
and U3292 (N_3292,N_2740,N_2843);
or U3293 (N_3293,N_2905,N_2833);
and U3294 (N_3294,N_2864,N_2528);
nor U3295 (N_3295,N_2942,N_2919);
nor U3296 (N_3296,N_2797,N_2803);
or U3297 (N_3297,N_2966,N_2762);
or U3298 (N_3298,N_2582,N_2855);
nor U3299 (N_3299,N_2948,N_2720);
nand U3300 (N_3300,N_2695,N_2544);
nor U3301 (N_3301,N_2671,N_2838);
nor U3302 (N_3302,N_2537,N_2514);
or U3303 (N_3303,N_2825,N_2847);
or U3304 (N_3304,N_2631,N_2849);
nor U3305 (N_3305,N_2601,N_2600);
xor U3306 (N_3306,N_2789,N_2632);
nor U3307 (N_3307,N_2518,N_2611);
nand U3308 (N_3308,N_2642,N_2560);
nor U3309 (N_3309,N_2646,N_2654);
xnor U3310 (N_3310,N_2726,N_2666);
nor U3311 (N_3311,N_2964,N_2707);
and U3312 (N_3312,N_2618,N_2842);
and U3313 (N_3313,N_2802,N_2590);
nor U3314 (N_3314,N_2642,N_2570);
and U3315 (N_3315,N_2621,N_2806);
xnor U3316 (N_3316,N_2766,N_2842);
or U3317 (N_3317,N_2944,N_2950);
nor U3318 (N_3318,N_2952,N_2687);
nand U3319 (N_3319,N_2762,N_2832);
nor U3320 (N_3320,N_2590,N_2930);
nor U3321 (N_3321,N_2981,N_2685);
nand U3322 (N_3322,N_2846,N_2792);
nor U3323 (N_3323,N_2817,N_2684);
xnor U3324 (N_3324,N_2657,N_2712);
and U3325 (N_3325,N_2774,N_2794);
or U3326 (N_3326,N_2553,N_2525);
nor U3327 (N_3327,N_2771,N_2527);
nand U3328 (N_3328,N_2948,N_2973);
and U3329 (N_3329,N_2760,N_2837);
xor U3330 (N_3330,N_2587,N_2564);
nor U3331 (N_3331,N_2709,N_2852);
and U3332 (N_3332,N_2928,N_2584);
or U3333 (N_3333,N_2770,N_2956);
nand U3334 (N_3334,N_2781,N_2943);
nand U3335 (N_3335,N_2588,N_2665);
nor U3336 (N_3336,N_2815,N_2852);
or U3337 (N_3337,N_2691,N_2839);
or U3338 (N_3338,N_2787,N_2973);
and U3339 (N_3339,N_2820,N_2865);
nor U3340 (N_3340,N_2593,N_2886);
nor U3341 (N_3341,N_2801,N_2605);
nand U3342 (N_3342,N_2642,N_2912);
and U3343 (N_3343,N_2845,N_2753);
or U3344 (N_3344,N_2672,N_2838);
or U3345 (N_3345,N_2588,N_2683);
and U3346 (N_3346,N_2593,N_2740);
xnor U3347 (N_3347,N_2769,N_2903);
and U3348 (N_3348,N_2552,N_2810);
nor U3349 (N_3349,N_2721,N_2787);
xnor U3350 (N_3350,N_2702,N_2724);
or U3351 (N_3351,N_2514,N_2993);
nor U3352 (N_3352,N_2751,N_2889);
or U3353 (N_3353,N_2593,N_2809);
or U3354 (N_3354,N_2915,N_2637);
nand U3355 (N_3355,N_2678,N_2598);
and U3356 (N_3356,N_2704,N_2932);
nand U3357 (N_3357,N_2690,N_2769);
or U3358 (N_3358,N_2804,N_2648);
nor U3359 (N_3359,N_2876,N_2833);
xnor U3360 (N_3360,N_2996,N_2961);
xnor U3361 (N_3361,N_2717,N_2596);
nand U3362 (N_3362,N_2892,N_2830);
nor U3363 (N_3363,N_2685,N_2946);
nand U3364 (N_3364,N_2763,N_2624);
nand U3365 (N_3365,N_2732,N_2790);
nor U3366 (N_3366,N_2649,N_2796);
and U3367 (N_3367,N_2859,N_2947);
and U3368 (N_3368,N_2601,N_2909);
nor U3369 (N_3369,N_2963,N_2510);
nor U3370 (N_3370,N_2861,N_2781);
nor U3371 (N_3371,N_2807,N_2542);
nor U3372 (N_3372,N_2989,N_2944);
or U3373 (N_3373,N_2939,N_2573);
nor U3374 (N_3374,N_2976,N_2968);
nand U3375 (N_3375,N_2720,N_2751);
xor U3376 (N_3376,N_2815,N_2991);
and U3377 (N_3377,N_2998,N_2828);
nand U3378 (N_3378,N_2668,N_2848);
nand U3379 (N_3379,N_2878,N_2566);
and U3380 (N_3380,N_2900,N_2823);
nand U3381 (N_3381,N_2851,N_2745);
or U3382 (N_3382,N_2771,N_2538);
nor U3383 (N_3383,N_2601,N_2703);
nor U3384 (N_3384,N_2900,N_2659);
or U3385 (N_3385,N_2936,N_2678);
nor U3386 (N_3386,N_2924,N_2752);
xnor U3387 (N_3387,N_2951,N_2526);
nand U3388 (N_3388,N_2928,N_2510);
nand U3389 (N_3389,N_2756,N_2572);
and U3390 (N_3390,N_2734,N_2689);
or U3391 (N_3391,N_2634,N_2651);
or U3392 (N_3392,N_2725,N_2664);
xnor U3393 (N_3393,N_2654,N_2990);
xnor U3394 (N_3394,N_2698,N_2864);
or U3395 (N_3395,N_2763,N_2647);
and U3396 (N_3396,N_2643,N_2983);
nand U3397 (N_3397,N_2866,N_2867);
or U3398 (N_3398,N_2825,N_2575);
nand U3399 (N_3399,N_2961,N_2882);
xor U3400 (N_3400,N_2727,N_2664);
and U3401 (N_3401,N_2644,N_2667);
nor U3402 (N_3402,N_2999,N_2770);
nor U3403 (N_3403,N_2538,N_2704);
or U3404 (N_3404,N_2792,N_2612);
or U3405 (N_3405,N_2809,N_2692);
or U3406 (N_3406,N_2616,N_2951);
and U3407 (N_3407,N_2691,N_2652);
nor U3408 (N_3408,N_2736,N_2742);
nand U3409 (N_3409,N_2967,N_2870);
and U3410 (N_3410,N_2566,N_2542);
nor U3411 (N_3411,N_2730,N_2751);
or U3412 (N_3412,N_2739,N_2764);
or U3413 (N_3413,N_2961,N_2593);
and U3414 (N_3414,N_2790,N_2583);
nor U3415 (N_3415,N_2993,N_2521);
or U3416 (N_3416,N_2812,N_2930);
nand U3417 (N_3417,N_2876,N_2714);
xor U3418 (N_3418,N_2675,N_2774);
and U3419 (N_3419,N_2532,N_2613);
nand U3420 (N_3420,N_2773,N_2959);
or U3421 (N_3421,N_2987,N_2949);
nand U3422 (N_3422,N_2639,N_2700);
and U3423 (N_3423,N_2809,N_2865);
and U3424 (N_3424,N_2682,N_2577);
xor U3425 (N_3425,N_2614,N_2994);
nor U3426 (N_3426,N_2548,N_2750);
nand U3427 (N_3427,N_2622,N_2605);
or U3428 (N_3428,N_2530,N_2772);
nand U3429 (N_3429,N_2811,N_2842);
or U3430 (N_3430,N_2939,N_2681);
nor U3431 (N_3431,N_2884,N_2676);
nor U3432 (N_3432,N_2983,N_2691);
and U3433 (N_3433,N_2829,N_2750);
or U3434 (N_3434,N_2676,N_2721);
xor U3435 (N_3435,N_2545,N_2504);
nand U3436 (N_3436,N_2986,N_2809);
nand U3437 (N_3437,N_2698,N_2724);
nand U3438 (N_3438,N_2630,N_2833);
and U3439 (N_3439,N_2500,N_2698);
or U3440 (N_3440,N_2708,N_2623);
xnor U3441 (N_3441,N_2961,N_2735);
nand U3442 (N_3442,N_2907,N_2671);
and U3443 (N_3443,N_2717,N_2987);
nor U3444 (N_3444,N_2577,N_2893);
nand U3445 (N_3445,N_2892,N_2548);
nor U3446 (N_3446,N_2961,N_2805);
and U3447 (N_3447,N_2790,N_2831);
or U3448 (N_3448,N_2601,N_2892);
and U3449 (N_3449,N_2966,N_2621);
and U3450 (N_3450,N_2855,N_2753);
and U3451 (N_3451,N_2529,N_2678);
nand U3452 (N_3452,N_2837,N_2934);
nand U3453 (N_3453,N_2770,N_2602);
and U3454 (N_3454,N_2559,N_2836);
or U3455 (N_3455,N_2601,N_2820);
or U3456 (N_3456,N_2544,N_2707);
xor U3457 (N_3457,N_2536,N_2517);
or U3458 (N_3458,N_2800,N_2810);
or U3459 (N_3459,N_2549,N_2798);
nor U3460 (N_3460,N_2595,N_2786);
nand U3461 (N_3461,N_2538,N_2893);
or U3462 (N_3462,N_2633,N_2721);
nor U3463 (N_3463,N_2945,N_2867);
nor U3464 (N_3464,N_2742,N_2806);
and U3465 (N_3465,N_2866,N_2798);
nor U3466 (N_3466,N_2666,N_2690);
nand U3467 (N_3467,N_2952,N_2705);
or U3468 (N_3468,N_2590,N_2938);
or U3469 (N_3469,N_2696,N_2832);
and U3470 (N_3470,N_2527,N_2573);
or U3471 (N_3471,N_2554,N_2630);
or U3472 (N_3472,N_2695,N_2901);
or U3473 (N_3473,N_2880,N_2917);
nand U3474 (N_3474,N_2928,N_2969);
nand U3475 (N_3475,N_2647,N_2922);
nor U3476 (N_3476,N_2758,N_2737);
nand U3477 (N_3477,N_2921,N_2688);
nand U3478 (N_3478,N_2908,N_2769);
nor U3479 (N_3479,N_2866,N_2733);
nor U3480 (N_3480,N_2872,N_2822);
nand U3481 (N_3481,N_2524,N_2915);
nand U3482 (N_3482,N_2821,N_2634);
nand U3483 (N_3483,N_2748,N_2860);
nor U3484 (N_3484,N_2926,N_2801);
nand U3485 (N_3485,N_2854,N_2940);
or U3486 (N_3486,N_2543,N_2616);
and U3487 (N_3487,N_2885,N_2662);
or U3488 (N_3488,N_2828,N_2624);
and U3489 (N_3489,N_2547,N_2855);
nand U3490 (N_3490,N_2620,N_2802);
nand U3491 (N_3491,N_2506,N_2933);
nor U3492 (N_3492,N_2734,N_2598);
nand U3493 (N_3493,N_2925,N_2670);
and U3494 (N_3494,N_2961,N_2953);
or U3495 (N_3495,N_2671,N_2899);
and U3496 (N_3496,N_2756,N_2639);
nand U3497 (N_3497,N_2883,N_2839);
and U3498 (N_3498,N_2759,N_2783);
nand U3499 (N_3499,N_2525,N_2939);
nand U3500 (N_3500,N_3245,N_3153);
nand U3501 (N_3501,N_3311,N_3075);
and U3502 (N_3502,N_3248,N_3031);
nor U3503 (N_3503,N_3186,N_3210);
or U3504 (N_3504,N_3390,N_3221);
xor U3505 (N_3505,N_3054,N_3293);
xor U3506 (N_3506,N_3430,N_3247);
xor U3507 (N_3507,N_3074,N_3070);
and U3508 (N_3508,N_3495,N_3159);
or U3509 (N_3509,N_3161,N_3331);
nand U3510 (N_3510,N_3276,N_3335);
or U3511 (N_3511,N_3488,N_3275);
xor U3512 (N_3512,N_3145,N_3058);
or U3513 (N_3513,N_3241,N_3137);
and U3514 (N_3514,N_3339,N_3396);
and U3515 (N_3515,N_3415,N_3484);
or U3516 (N_3516,N_3223,N_3472);
nor U3517 (N_3517,N_3359,N_3269);
nand U3518 (N_3518,N_3346,N_3177);
xor U3519 (N_3519,N_3330,N_3199);
or U3520 (N_3520,N_3315,N_3402);
nor U3521 (N_3521,N_3250,N_3085);
nor U3522 (N_3522,N_3071,N_3499);
nor U3523 (N_3523,N_3020,N_3427);
nand U3524 (N_3524,N_3291,N_3365);
and U3525 (N_3525,N_3312,N_3433);
nand U3526 (N_3526,N_3013,N_3176);
and U3527 (N_3527,N_3446,N_3483);
or U3528 (N_3528,N_3441,N_3323);
nor U3529 (N_3529,N_3404,N_3461);
nor U3530 (N_3530,N_3357,N_3094);
nand U3531 (N_3531,N_3324,N_3443);
nor U3532 (N_3532,N_3108,N_3478);
nor U3533 (N_3533,N_3208,N_3061);
and U3534 (N_3534,N_3367,N_3140);
or U3535 (N_3535,N_3188,N_3237);
and U3536 (N_3536,N_3406,N_3105);
nor U3537 (N_3537,N_3400,N_3109);
xor U3538 (N_3538,N_3340,N_3420);
xor U3539 (N_3539,N_3374,N_3416);
xnor U3540 (N_3540,N_3288,N_3240);
or U3541 (N_3541,N_3076,N_3278);
or U3542 (N_3542,N_3296,N_3120);
nor U3543 (N_3543,N_3325,N_3258);
xor U3544 (N_3544,N_3068,N_3086);
or U3545 (N_3545,N_3187,N_3169);
and U3546 (N_3546,N_3219,N_3381);
xor U3547 (N_3547,N_3313,N_3097);
nor U3548 (N_3548,N_3040,N_3473);
nand U3549 (N_3549,N_3211,N_3280);
xor U3550 (N_3550,N_3256,N_3066);
nand U3551 (N_3551,N_3289,N_3078);
nor U3552 (N_3552,N_3091,N_3203);
nor U3553 (N_3553,N_3053,N_3206);
or U3554 (N_3554,N_3236,N_3252);
nor U3555 (N_3555,N_3314,N_3398);
or U3556 (N_3556,N_3419,N_3093);
xor U3557 (N_3557,N_3361,N_3423);
xnor U3558 (N_3558,N_3224,N_3401);
nand U3559 (N_3559,N_3025,N_3360);
xor U3560 (N_3560,N_3294,N_3088);
nand U3561 (N_3561,N_3144,N_3142);
xor U3562 (N_3562,N_3307,N_3028);
nor U3563 (N_3563,N_3116,N_3050);
nor U3564 (N_3564,N_3281,N_3439);
nand U3565 (N_3565,N_3038,N_3336);
nor U3566 (N_3566,N_3225,N_3422);
and U3567 (N_3567,N_3164,N_3320);
and U3568 (N_3568,N_3175,N_3304);
and U3569 (N_3569,N_3363,N_3290);
and U3570 (N_3570,N_3214,N_3337);
and U3571 (N_3571,N_3309,N_3069);
nor U3572 (N_3572,N_3021,N_3003);
nand U3573 (N_3573,N_3101,N_3477);
nor U3574 (N_3574,N_3308,N_3274);
nor U3575 (N_3575,N_3270,N_3019);
and U3576 (N_3576,N_3128,N_3080);
nor U3577 (N_3577,N_3267,N_3466);
and U3578 (N_3578,N_3004,N_3012);
and U3579 (N_3579,N_3264,N_3182);
nand U3580 (N_3580,N_3067,N_3480);
xor U3581 (N_3581,N_3492,N_3371);
nor U3582 (N_3582,N_3233,N_3138);
or U3583 (N_3583,N_3130,N_3229);
and U3584 (N_3584,N_3372,N_3139);
nand U3585 (N_3585,N_3126,N_3190);
nand U3586 (N_3586,N_3005,N_3122);
and U3587 (N_3587,N_3351,N_3102);
nor U3588 (N_3588,N_3178,N_3165);
and U3589 (N_3589,N_3023,N_3462);
nor U3590 (N_3590,N_3016,N_3081);
nand U3591 (N_3591,N_3123,N_3077);
or U3592 (N_3592,N_3112,N_3437);
and U3593 (N_3593,N_3213,N_3015);
and U3594 (N_3594,N_3470,N_3448);
or U3595 (N_3595,N_3482,N_3300);
or U3596 (N_3596,N_3228,N_3118);
or U3597 (N_3597,N_3368,N_3306);
or U3598 (N_3598,N_3403,N_3060);
nor U3599 (N_3599,N_3163,N_3425);
and U3600 (N_3600,N_3471,N_3205);
or U3601 (N_3601,N_3172,N_3166);
nand U3602 (N_3602,N_3200,N_3295);
xor U3603 (N_3603,N_3405,N_3317);
and U3604 (N_3604,N_3469,N_3379);
nor U3605 (N_3605,N_3217,N_3260);
and U3606 (N_3606,N_3220,N_3171);
nand U3607 (N_3607,N_3111,N_3079);
nor U3608 (N_3608,N_3344,N_3442);
nand U3609 (N_3609,N_3431,N_3254);
and U3610 (N_3610,N_3132,N_3121);
or U3611 (N_3611,N_3271,N_3486);
and U3612 (N_3612,N_3418,N_3204);
nor U3613 (N_3613,N_3222,N_3387);
xor U3614 (N_3614,N_3485,N_3436);
nor U3615 (N_3615,N_3282,N_3487);
or U3616 (N_3616,N_3476,N_3407);
nor U3617 (N_3617,N_3460,N_3454);
nor U3618 (N_3618,N_3366,N_3251);
or U3619 (N_3619,N_3410,N_3388);
or U3620 (N_3620,N_3494,N_3035);
nand U3621 (N_3621,N_3029,N_3392);
and U3622 (N_3622,N_3207,N_3150);
nand U3623 (N_3623,N_3424,N_3393);
and U3624 (N_3624,N_3319,N_3095);
and U3625 (N_3625,N_3409,N_3239);
nand U3626 (N_3626,N_3292,N_3151);
xor U3627 (N_3627,N_3327,N_3244);
nor U3628 (N_3628,N_3378,N_3043);
xnor U3629 (N_3629,N_3168,N_3391);
nand U3630 (N_3630,N_3343,N_3198);
nor U3631 (N_3631,N_3302,N_3156);
and U3632 (N_3632,N_3183,N_3435);
or U3633 (N_3633,N_3475,N_3257);
or U3634 (N_3634,N_3285,N_3262);
or U3635 (N_3635,N_3273,N_3226);
and U3636 (N_3636,N_3113,N_3334);
or U3637 (N_3637,N_3106,N_3141);
xor U3638 (N_3638,N_3380,N_3065);
nor U3639 (N_3639,N_3179,N_3197);
and U3640 (N_3640,N_3232,N_3429);
and U3641 (N_3641,N_3303,N_3474);
and U3642 (N_3642,N_3155,N_3318);
nand U3643 (N_3643,N_3279,N_3459);
xor U3644 (N_3644,N_3463,N_3100);
nand U3645 (N_3645,N_3490,N_3215);
or U3646 (N_3646,N_3148,N_3457);
or U3647 (N_3647,N_3417,N_3234);
or U3648 (N_3648,N_3087,N_3310);
and U3649 (N_3649,N_3338,N_3468);
nand U3650 (N_3650,N_3026,N_3090);
or U3651 (N_3651,N_3052,N_3047);
and U3652 (N_3652,N_3453,N_3243);
nor U3653 (N_3653,N_3376,N_3249);
nor U3654 (N_3654,N_3063,N_3115);
nand U3655 (N_3655,N_3209,N_3147);
nor U3656 (N_3656,N_3125,N_3196);
nor U3657 (N_3657,N_3057,N_3297);
or U3658 (N_3658,N_3399,N_3193);
nor U3659 (N_3659,N_3456,N_3212);
nor U3660 (N_3660,N_3353,N_3041);
and U3661 (N_3661,N_3096,N_3014);
nand U3662 (N_3662,N_3479,N_3099);
and U3663 (N_3663,N_3298,N_3135);
or U3664 (N_3664,N_3369,N_3259);
nor U3665 (N_3665,N_3174,N_3497);
or U3666 (N_3666,N_3238,N_3027);
nand U3667 (N_3667,N_3467,N_3322);
xnor U3668 (N_3668,N_3286,N_3167);
and U3669 (N_3669,N_3024,N_3465);
nand U3670 (N_3670,N_3489,N_3354);
and U3671 (N_3671,N_3450,N_3265);
xor U3672 (N_3672,N_3133,N_3036);
nand U3673 (N_3673,N_3358,N_3434);
xor U3674 (N_3674,N_3355,N_3364);
nor U3675 (N_3675,N_3049,N_3373);
or U3676 (N_3676,N_3055,N_3333);
and U3677 (N_3677,N_3192,N_3328);
and U3678 (N_3678,N_3496,N_3356);
or U3679 (N_3679,N_3082,N_3493);
or U3680 (N_3680,N_3481,N_3136);
or U3681 (N_3681,N_3386,N_3129);
and U3682 (N_3682,N_3329,N_3152);
and U3683 (N_3683,N_3377,N_3117);
or U3684 (N_3684,N_3173,N_3498);
or U3685 (N_3685,N_3412,N_3154);
or U3686 (N_3686,N_3246,N_3455);
nand U3687 (N_3687,N_3134,N_3056);
or U3688 (N_3688,N_3006,N_3253);
nor U3689 (N_3689,N_3184,N_3255);
or U3690 (N_3690,N_3332,N_3449);
nand U3691 (N_3691,N_3157,N_3261);
nand U3692 (N_3692,N_3451,N_3440);
and U3693 (N_3693,N_3119,N_3149);
nor U3694 (N_3694,N_3321,N_3002);
nand U3695 (N_3695,N_3444,N_3202);
nor U3696 (N_3696,N_3131,N_3458);
and U3697 (N_3697,N_3413,N_3445);
or U3698 (N_3698,N_3326,N_3008);
and U3699 (N_3699,N_3411,N_3432);
nand U3700 (N_3700,N_3185,N_3037);
nor U3701 (N_3701,N_3143,N_3235);
nor U3702 (N_3702,N_3110,N_3084);
and U3703 (N_3703,N_3158,N_3341);
and U3704 (N_3704,N_3194,N_3051);
nand U3705 (N_3705,N_3370,N_3059);
nor U3706 (N_3706,N_3266,N_3064);
or U3707 (N_3707,N_3114,N_3042);
nor U3708 (N_3708,N_3438,N_3072);
nor U3709 (N_3709,N_3127,N_3218);
nand U3710 (N_3710,N_3414,N_3104);
or U3711 (N_3711,N_3352,N_3301);
nand U3712 (N_3712,N_3103,N_3464);
nor U3713 (N_3713,N_3045,N_3375);
or U3714 (N_3714,N_3385,N_3347);
xnor U3715 (N_3715,N_3010,N_3034);
and U3716 (N_3716,N_3170,N_3089);
nand U3717 (N_3717,N_3083,N_3046);
or U3718 (N_3718,N_3384,N_3287);
nor U3719 (N_3719,N_3011,N_3350);
nor U3720 (N_3720,N_3342,N_3033);
and U3721 (N_3721,N_3394,N_3382);
and U3722 (N_3722,N_3022,N_3428);
nor U3723 (N_3723,N_3272,N_3277);
nand U3724 (N_3724,N_3426,N_3421);
and U3725 (N_3725,N_3395,N_3268);
or U3726 (N_3726,N_3345,N_3007);
or U3727 (N_3727,N_3349,N_3397);
nand U3728 (N_3728,N_3009,N_3201);
nor U3729 (N_3729,N_3048,N_3231);
nor U3730 (N_3730,N_3124,N_3062);
and U3731 (N_3731,N_3098,N_3160);
or U3732 (N_3732,N_3018,N_3284);
nor U3733 (N_3733,N_3242,N_3146);
nor U3734 (N_3734,N_3039,N_3107);
nor U3735 (N_3735,N_3030,N_3180);
nor U3736 (N_3736,N_3283,N_3227);
and U3737 (N_3737,N_3017,N_3230);
xnor U3738 (N_3738,N_3299,N_3189);
or U3739 (N_3739,N_3044,N_3452);
xnor U3740 (N_3740,N_3162,N_3408);
and U3741 (N_3741,N_3305,N_3001);
and U3742 (N_3742,N_3181,N_3316);
nand U3743 (N_3743,N_3000,N_3195);
nor U3744 (N_3744,N_3348,N_3383);
nor U3745 (N_3745,N_3389,N_3491);
and U3746 (N_3746,N_3032,N_3092);
and U3747 (N_3747,N_3362,N_3191);
and U3748 (N_3748,N_3447,N_3073);
or U3749 (N_3749,N_3263,N_3216);
nand U3750 (N_3750,N_3050,N_3316);
or U3751 (N_3751,N_3496,N_3227);
and U3752 (N_3752,N_3354,N_3298);
xor U3753 (N_3753,N_3277,N_3424);
nand U3754 (N_3754,N_3008,N_3423);
xor U3755 (N_3755,N_3169,N_3295);
nand U3756 (N_3756,N_3107,N_3247);
and U3757 (N_3757,N_3278,N_3260);
or U3758 (N_3758,N_3009,N_3255);
xnor U3759 (N_3759,N_3480,N_3006);
or U3760 (N_3760,N_3320,N_3020);
nand U3761 (N_3761,N_3343,N_3334);
nor U3762 (N_3762,N_3109,N_3258);
or U3763 (N_3763,N_3327,N_3215);
or U3764 (N_3764,N_3066,N_3252);
and U3765 (N_3765,N_3477,N_3151);
or U3766 (N_3766,N_3438,N_3129);
nand U3767 (N_3767,N_3415,N_3155);
nand U3768 (N_3768,N_3102,N_3081);
or U3769 (N_3769,N_3096,N_3142);
or U3770 (N_3770,N_3495,N_3149);
xnor U3771 (N_3771,N_3199,N_3443);
nand U3772 (N_3772,N_3291,N_3457);
nand U3773 (N_3773,N_3191,N_3364);
nand U3774 (N_3774,N_3223,N_3424);
and U3775 (N_3775,N_3080,N_3162);
xor U3776 (N_3776,N_3362,N_3115);
and U3777 (N_3777,N_3310,N_3295);
nand U3778 (N_3778,N_3064,N_3315);
xnor U3779 (N_3779,N_3125,N_3386);
nor U3780 (N_3780,N_3423,N_3245);
and U3781 (N_3781,N_3200,N_3349);
or U3782 (N_3782,N_3438,N_3046);
and U3783 (N_3783,N_3392,N_3399);
nand U3784 (N_3784,N_3484,N_3260);
nor U3785 (N_3785,N_3098,N_3464);
nor U3786 (N_3786,N_3211,N_3024);
nor U3787 (N_3787,N_3211,N_3242);
nor U3788 (N_3788,N_3036,N_3258);
or U3789 (N_3789,N_3022,N_3134);
nand U3790 (N_3790,N_3084,N_3126);
xnor U3791 (N_3791,N_3115,N_3009);
and U3792 (N_3792,N_3338,N_3321);
or U3793 (N_3793,N_3417,N_3133);
xnor U3794 (N_3794,N_3081,N_3492);
and U3795 (N_3795,N_3454,N_3463);
nor U3796 (N_3796,N_3213,N_3203);
and U3797 (N_3797,N_3226,N_3415);
and U3798 (N_3798,N_3043,N_3262);
or U3799 (N_3799,N_3220,N_3230);
and U3800 (N_3800,N_3197,N_3079);
nand U3801 (N_3801,N_3137,N_3248);
or U3802 (N_3802,N_3440,N_3047);
xor U3803 (N_3803,N_3050,N_3417);
xnor U3804 (N_3804,N_3206,N_3434);
nor U3805 (N_3805,N_3002,N_3355);
nand U3806 (N_3806,N_3489,N_3408);
xnor U3807 (N_3807,N_3001,N_3137);
nor U3808 (N_3808,N_3015,N_3140);
and U3809 (N_3809,N_3393,N_3271);
xor U3810 (N_3810,N_3273,N_3473);
nand U3811 (N_3811,N_3249,N_3450);
nand U3812 (N_3812,N_3243,N_3122);
and U3813 (N_3813,N_3443,N_3362);
xor U3814 (N_3814,N_3052,N_3285);
xor U3815 (N_3815,N_3466,N_3442);
or U3816 (N_3816,N_3476,N_3196);
nand U3817 (N_3817,N_3207,N_3417);
or U3818 (N_3818,N_3258,N_3319);
or U3819 (N_3819,N_3419,N_3038);
and U3820 (N_3820,N_3214,N_3477);
and U3821 (N_3821,N_3016,N_3368);
nand U3822 (N_3822,N_3364,N_3395);
and U3823 (N_3823,N_3443,N_3448);
and U3824 (N_3824,N_3399,N_3294);
nand U3825 (N_3825,N_3024,N_3401);
nor U3826 (N_3826,N_3267,N_3310);
or U3827 (N_3827,N_3194,N_3443);
xor U3828 (N_3828,N_3032,N_3204);
and U3829 (N_3829,N_3152,N_3201);
nand U3830 (N_3830,N_3292,N_3340);
nor U3831 (N_3831,N_3311,N_3332);
or U3832 (N_3832,N_3066,N_3289);
and U3833 (N_3833,N_3271,N_3097);
and U3834 (N_3834,N_3286,N_3078);
or U3835 (N_3835,N_3001,N_3340);
nand U3836 (N_3836,N_3281,N_3136);
nor U3837 (N_3837,N_3356,N_3308);
nor U3838 (N_3838,N_3358,N_3124);
nand U3839 (N_3839,N_3200,N_3192);
or U3840 (N_3840,N_3027,N_3358);
or U3841 (N_3841,N_3420,N_3404);
or U3842 (N_3842,N_3206,N_3241);
nor U3843 (N_3843,N_3314,N_3278);
or U3844 (N_3844,N_3376,N_3090);
nor U3845 (N_3845,N_3049,N_3413);
or U3846 (N_3846,N_3225,N_3223);
or U3847 (N_3847,N_3484,N_3058);
or U3848 (N_3848,N_3315,N_3163);
or U3849 (N_3849,N_3405,N_3289);
nor U3850 (N_3850,N_3236,N_3253);
xnor U3851 (N_3851,N_3252,N_3489);
nand U3852 (N_3852,N_3079,N_3471);
and U3853 (N_3853,N_3270,N_3487);
nor U3854 (N_3854,N_3415,N_3162);
and U3855 (N_3855,N_3368,N_3121);
and U3856 (N_3856,N_3340,N_3110);
nor U3857 (N_3857,N_3411,N_3075);
nor U3858 (N_3858,N_3476,N_3054);
or U3859 (N_3859,N_3006,N_3136);
and U3860 (N_3860,N_3313,N_3471);
and U3861 (N_3861,N_3214,N_3368);
nand U3862 (N_3862,N_3032,N_3197);
nor U3863 (N_3863,N_3350,N_3320);
nand U3864 (N_3864,N_3079,N_3151);
nor U3865 (N_3865,N_3441,N_3269);
and U3866 (N_3866,N_3281,N_3485);
and U3867 (N_3867,N_3381,N_3448);
nor U3868 (N_3868,N_3049,N_3086);
nand U3869 (N_3869,N_3361,N_3225);
and U3870 (N_3870,N_3175,N_3339);
xor U3871 (N_3871,N_3303,N_3365);
and U3872 (N_3872,N_3200,N_3111);
nor U3873 (N_3873,N_3487,N_3164);
nand U3874 (N_3874,N_3061,N_3292);
or U3875 (N_3875,N_3356,N_3030);
nor U3876 (N_3876,N_3272,N_3120);
or U3877 (N_3877,N_3385,N_3205);
or U3878 (N_3878,N_3437,N_3303);
nand U3879 (N_3879,N_3213,N_3373);
nand U3880 (N_3880,N_3292,N_3455);
and U3881 (N_3881,N_3291,N_3339);
and U3882 (N_3882,N_3313,N_3300);
and U3883 (N_3883,N_3360,N_3386);
or U3884 (N_3884,N_3324,N_3059);
or U3885 (N_3885,N_3084,N_3273);
or U3886 (N_3886,N_3305,N_3384);
nand U3887 (N_3887,N_3212,N_3400);
and U3888 (N_3888,N_3115,N_3154);
or U3889 (N_3889,N_3443,N_3460);
nand U3890 (N_3890,N_3105,N_3292);
and U3891 (N_3891,N_3387,N_3382);
and U3892 (N_3892,N_3219,N_3169);
and U3893 (N_3893,N_3082,N_3004);
nor U3894 (N_3894,N_3109,N_3428);
and U3895 (N_3895,N_3202,N_3443);
nor U3896 (N_3896,N_3267,N_3181);
nand U3897 (N_3897,N_3060,N_3004);
and U3898 (N_3898,N_3075,N_3082);
nand U3899 (N_3899,N_3024,N_3041);
nor U3900 (N_3900,N_3277,N_3175);
and U3901 (N_3901,N_3090,N_3074);
nand U3902 (N_3902,N_3351,N_3064);
nor U3903 (N_3903,N_3265,N_3153);
nor U3904 (N_3904,N_3414,N_3112);
nand U3905 (N_3905,N_3456,N_3062);
or U3906 (N_3906,N_3040,N_3290);
nor U3907 (N_3907,N_3094,N_3428);
or U3908 (N_3908,N_3174,N_3492);
xor U3909 (N_3909,N_3201,N_3252);
and U3910 (N_3910,N_3376,N_3035);
or U3911 (N_3911,N_3051,N_3363);
nand U3912 (N_3912,N_3125,N_3476);
or U3913 (N_3913,N_3195,N_3073);
or U3914 (N_3914,N_3369,N_3458);
nor U3915 (N_3915,N_3039,N_3228);
nor U3916 (N_3916,N_3152,N_3205);
nand U3917 (N_3917,N_3489,N_3265);
nand U3918 (N_3918,N_3179,N_3435);
nand U3919 (N_3919,N_3152,N_3291);
and U3920 (N_3920,N_3104,N_3424);
or U3921 (N_3921,N_3418,N_3375);
nand U3922 (N_3922,N_3138,N_3156);
xnor U3923 (N_3923,N_3375,N_3306);
nand U3924 (N_3924,N_3176,N_3401);
nand U3925 (N_3925,N_3204,N_3037);
and U3926 (N_3926,N_3088,N_3168);
or U3927 (N_3927,N_3011,N_3009);
xnor U3928 (N_3928,N_3208,N_3036);
and U3929 (N_3929,N_3170,N_3384);
nand U3930 (N_3930,N_3106,N_3117);
nor U3931 (N_3931,N_3170,N_3035);
nand U3932 (N_3932,N_3058,N_3450);
nand U3933 (N_3933,N_3016,N_3206);
nand U3934 (N_3934,N_3008,N_3071);
or U3935 (N_3935,N_3446,N_3227);
xor U3936 (N_3936,N_3460,N_3306);
or U3937 (N_3937,N_3273,N_3179);
nor U3938 (N_3938,N_3421,N_3133);
nor U3939 (N_3939,N_3293,N_3136);
nor U3940 (N_3940,N_3263,N_3365);
nor U3941 (N_3941,N_3464,N_3248);
xnor U3942 (N_3942,N_3213,N_3100);
and U3943 (N_3943,N_3056,N_3361);
xor U3944 (N_3944,N_3186,N_3425);
or U3945 (N_3945,N_3033,N_3115);
and U3946 (N_3946,N_3435,N_3292);
or U3947 (N_3947,N_3190,N_3449);
nand U3948 (N_3948,N_3479,N_3471);
and U3949 (N_3949,N_3212,N_3463);
nor U3950 (N_3950,N_3122,N_3242);
nor U3951 (N_3951,N_3473,N_3055);
nor U3952 (N_3952,N_3487,N_3109);
or U3953 (N_3953,N_3331,N_3403);
nor U3954 (N_3954,N_3465,N_3316);
nand U3955 (N_3955,N_3484,N_3072);
and U3956 (N_3956,N_3029,N_3101);
nor U3957 (N_3957,N_3273,N_3241);
nand U3958 (N_3958,N_3135,N_3372);
and U3959 (N_3959,N_3391,N_3005);
nor U3960 (N_3960,N_3238,N_3036);
or U3961 (N_3961,N_3059,N_3169);
nand U3962 (N_3962,N_3338,N_3289);
nor U3963 (N_3963,N_3201,N_3042);
and U3964 (N_3964,N_3046,N_3335);
and U3965 (N_3965,N_3460,N_3010);
nor U3966 (N_3966,N_3101,N_3272);
nand U3967 (N_3967,N_3322,N_3125);
nand U3968 (N_3968,N_3266,N_3441);
nand U3969 (N_3969,N_3080,N_3220);
nor U3970 (N_3970,N_3354,N_3329);
and U3971 (N_3971,N_3275,N_3496);
nand U3972 (N_3972,N_3029,N_3428);
nor U3973 (N_3973,N_3463,N_3104);
nor U3974 (N_3974,N_3441,N_3348);
nor U3975 (N_3975,N_3242,N_3123);
nor U3976 (N_3976,N_3095,N_3326);
or U3977 (N_3977,N_3464,N_3019);
or U3978 (N_3978,N_3116,N_3386);
or U3979 (N_3979,N_3237,N_3160);
and U3980 (N_3980,N_3426,N_3497);
nor U3981 (N_3981,N_3271,N_3065);
or U3982 (N_3982,N_3349,N_3419);
nand U3983 (N_3983,N_3353,N_3059);
nand U3984 (N_3984,N_3171,N_3277);
nor U3985 (N_3985,N_3487,N_3001);
xor U3986 (N_3986,N_3090,N_3358);
nand U3987 (N_3987,N_3288,N_3379);
or U3988 (N_3988,N_3265,N_3448);
and U3989 (N_3989,N_3337,N_3052);
xor U3990 (N_3990,N_3167,N_3356);
nand U3991 (N_3991,N_3022,N_3147);
and U3992 (N_3992,N_3245,N_3159);
nand U3993 (N_3993,N_3267,N_3422);
nand U3994 (N_3994,N_3260,N_3368);
xnor U3995 (N_3995,N_3297,N_3088);
or U3996 (N_3996,N_3444,N_3438);
nand U3997 (N_3997,N_3439,N_3154);
nor U3998 (N_3998,N_3288,N_3220);
and U3999 (N_3999,N_3247,N_3362);
nand U4000 (N_4000,N_3572,N_3715);
nor U4001 (N_4001,N_3696,N_3523);
nand U4002 (N_4002,N_3993,N_3796);
nand U4003 (N_4003,N_3602,N_3971);
or U4004 (N_4004,N_3798,N_3877);
nand U4005 (N_4005,N_3812,N_3830);
xnor U4006 (N_4006,N_3789,N_3721);
and U4007 (N_4007,N_3799,N_3889);
xnor U4008 (N_4008,N_3778,N_3599);
and U4009 (N_4009,N_3703,N_3793);
nor U4010 (N_4010,N_3510,N_3831);
nor U4011 (N_4011,N_3724,N_3873);
nand U4012 (N_4012,N_3712,N_3671);
nor U4013 (N_4013,N_3591,N_3861);
and U4014 (N_4014,N_3905,N_3780);
xor U4015 (N_4015,N_3577,N_3891);
or U4016 (N_4016,N_3818,N_3823);
and U4017 (N_4017,N_3512,N_3767);
xor U4018 (N_4018,N_3554,N_3960);
nand U4019 (N_4019,N_3833,N_3965);
nand U4020 (N_4020,N_3963,N_3722);
and U4021 (N_4021,N_3999,N_3782);
or U4022 (N_4022,N_3566,N_3837);
or U4023 (N_4023,N_3855,N_3533);
or U4024 (N_4024,N_3895,N_3995);
nor U4025 (N_4025,N_3913,N_3632);
nor U4026 (N_4026,N_3879,N_3676);
xnor U4027 (N_4027,N_3740,N_3569);
nor U4028 (N_4028,N_3717,N_3675);
nand U4029 (N_4029,N_3530,N_3504);
xnor U4030 (N_4030,N_3841,N_3773);
nand U4031 (N_4031,N_3686,N_3662);
nand U4032 (N_4032,N_3856,N_3629);
and U4033 (N_4033,N_3628,N_3957);
and U4034 (N_4034,N_3862,N_3922);
nand U4035 (N_4035,N_3945,N_3790);
and U4036 (N_4036,N_3807,N_3754);
or U4037 (N_4037,N_3700,N_3802);
nor U4038 (N_4038,N_3911,N_3529);
xor U4039 (N_4039,N_3763,N_3613);
or U4040 (N_4040,N_3612,N_3786);
nor U4041 (N_4041,N_3770,N_3852);
xor U4042 (N_4042,N_3859,N_3977);
nand U4043 (N_4043,N_3906,N_3923);
and U4044 (N_4044,N_3944,N_3817);
and U4045 (N_4045,N_3570,N_3907);
and U4046 (N_4046,N_3926,N_3551);
nand U4047 (N_4047,N_3751,N_3701);
and U4048 (N_4048,N_3562,N_3985);
nand U4049 (N_4049,N_3594,N_3505);
nand U4050 (N_4050,N_3728,N_3667);
nand U4051 (N_4051,N_3956,N_3766);
xnor U4052 (N_4052,N_3947,N_3734);
nand U4053 (N_4053,N_3731,N_3981);
xnor U4054 (N_4054,N_3704,N_3994);
nand U4055 (N_4055,N_3986,N_3794);
or U4056 (N_4056,N_3730,N_3609);
nor U4057 (N_4057,N_3847,N_3652);
or U4058 (N_4058,N_3943,N_3908);
nor U4059 (N_4059,N_3635,N_3561);
nand U4060 (N_4060,N_3645,N_3500);
and U4061 (N_4061,N_3713,N_3509);
xor U4062 (N_4062,N_3982,N_3522);
or U4063 (N_4063,N_3863,N_3772);
nor U4064 (N_4064,N_3897,N_3586);
nand U4065 (N_4065,N_3804,N_3605);
nor U4066 (N_4066,N_3828,N_3540);
or U4067 (N_4067,N_3716,N_3653);
and U4068 (N_4068,N_3885,N_3867);
and U4069 (N_4069,N_3827,N_3611);
and U4070 (N_4070,N_3992,N_3596);
nand U4071 (N_4071,N_3840,N_3835);
and U4072 (N_4072,N_3702,N_3921);
nand U4073 (N_4073,N_3545,N_3816);
nand U4074 (N_4074,N_3669,N_3948);
and U4075 (N_4075,N_3688,N_3918);
nand U4076 (N_4076,N_3720,N_3881);
or U4077 (N_4077,N_3692,N_3845);
nand U4078 (N_4078,N_3511,N_3964);
nand U4079 (N_4079,N_3825,N_3544);
nor U4080 (N_4080,N_3539,N_3775);
or U4081 (N_4081,N_3822,N_3685);
xor U4082 (N_4082,N_3593,N_3501);
nor U4083 (N_4083,N_3542,N_3574);
and U4084 (N_4084,N_3746,N_3784);
and U4085 (N_4085,N_3541,N_3683);
nor U4086 (N_4086,N_3984,N_3508);
or U4087 (N_4087,N_3869,N_3709);
or U4088 (N_4088,N_3547,N_3564);
nor U4089 (N_4089,N_3699,N_3904);
nand U4090 (N_4090,N_3616,N_3990);
or U4091 (N_4091,N_3887,N_3914);
nor U4092 (N_4092,N_3806,N_3958);
nor U4093 (N_4093,N_3756,N_3664);
or U4094 (N_4094,N_3910,N_3502);
nand U4095 (N_4095,N_3872,N_3550);
or U4096 (N_4096,N_3689,N_3998);
and U4097 (N_4097,N_3567,N_3819);
or U4098 (N_4098,N_3896,N_3785);
nor U4099 (N_4099,N_3627,N_3748);
and U4100 (N_4100,N_3691,N_3900);
nor U4101 (N_4101,N_3928,N_3868);
nand U4102 (N_4102,N_3520,N_3656);
and U4103 (N_4103,N_3968,N_3880);
or U4104 (N_4104,N_3589,N_3949);
and U4105 (N_4105,N_3579,N_3739);
nand U4106 (N_4106,N_3864,N_3742);
nor U4107 (N_4107,N_3568,N_3648);
nor U4108 (N_4108,N_3610,N_3650);
and U4109 (N_4109,N_3838,N_3595);
or U4110 (N_4110,N_3848,N_3821);
nand U4111 (N_4111,N_3854,N_3665);
xnor U4112 (N_4112,N_3987,N_3902);
and U4113 (N_4113,N_3846,N_3557);
and U4114 (N_4114,N_3598,N_3558);
and U4115 (N_4115,N_3601,N_3776);
or U4116 (N_4116,N_3711,N_3800);
nand U4117 (N_4117,N_3658,N_3883);
and U4118 (N_4118,N_3563,N_3976);
nor U4119 (N_4119,N_3925,N_3916);
xor U4120 (N_4120,N_3513,N_3576);
nand U4121 (N_4121,N_3693,N_3970);
or U4122 (N_4122,N_3639,N_3638);
and U4123 (N_4123,N_3524,N_3866);
or U4124 (N_4124,N_3917,N_3655);
nor U4125 (N_4125,N_3608,N_3744);
or U4126 (N_4126,N_3663,N_3870);
and U4127 (N_4127,N_3884,N_3537);
or U4128 (N_4128,N_3587,N_3761);
or U4129 (N_4129,N_3829,N_3874);
and U4130 (N_4130,N_3849,N_3661);
and U4131 (N_4131,N_3506,N_3666);
or U4132 (N_4132,N_3839,N_3938);
or U4133 (N_4133,N_3826,N_3503);
nor U4134 (N_4134,N_3811,N_3953);
nor U4135 (N_4135,N_3860,N_3741);
nor U4136 (N_4136,N_3718,N_3725);
xnor U4137 (N_4137,N_3644,N_3969);
and U4138 (N_4138,N_3952,N_3955);
xor U4139 (N_4139,N_3525,N_3732);
or U4140 (N_4140,N_3603,N_3736);
nand U4141 (N_4141,N_3507,N_3706);
xor U4142 (N_4142,N_3912,N_3966);
or U4143 (N_4143,N_3585,N_3747);
or U4144 (N_4144,N_3946,N_3929);
nand U4145 (N_4145,N_3619,N_3961);
or U4146 (N_4146,N_3623,N_3707);
nand U4147 (N_4147,N_3774,N_3979);
or U4148 (N_4148,N_3634,N_3677);
xnor U4149 (N_4149,N_3705,N_3690);
nand U4150 (N_4150,N_3764,N_3901);
nand U4151 (N_4151,N_3927,N_3851);
nor U4152 (N_4152,N_3556,N_3548);
and U4153 (N_4153,N_3758,N_3626);
and U4154 (N_4154,N_3636,N_3824);
and U4155 (N_4155,N_3983,N_3573);
or U4156 (N_4156,N_3625,N_3515);
nand U4157 (N_4157,N_3934,N_3865);
nand U4158 (N_4158,N_3582,N_3850);
or U4159 (N_4159,N_3792,N_3719);
nor U4160 (N_4160,N_3814,N_3755);
nand U4161 (N_4161,N_3882,N_3890);
nor U4162 (N_4162,N_3803,N_3801);
nand U4163 (N_4163,N_3937,N_3678);
xor U4164 (N_4164,N_3622,N_3516);
nor U4165 (N_4165,N_3980,N_3941);
nor U4166 (N_4166,N_3942,N_3989);
nor U4167 (N_4167,N_3649,N_3588);
nand U4168 (N_4168,N_3538,N_3654);
and U4169 (N_4169,N_3931,N_3886);
and U4170 (N_4170,N_3519,N_3932);
or U4171 (N_4171,N_3749,N_3543);
nor U4172 (N_4172,N_3695,N_3876);
nand U4173 (N_4173,N_3991,N_3805);
and U4174 (N_4174,N_3681,N_3808);
and U4175 (N_4175,N_3777,N_3614);
nand U4176 (N_4176,N_3668,N_3621);
or U4177 (N_4177,N_3810,N_3682);
and U4178 (N_4178,N_3752,N_3973);
xnor U4179 (N_4179,N_3518,N_3624);
or U4180 (N_4180,N_3997,N_3618);
nand U4181 (N_4181,N_3679,N_3630);
xor U4182 (N_4182,N_3531,N_3844);
or U4183 (N_4183,N_3698,N_3714);
nand U4184 (N_4184,N_3894,N_3892);
xnor U4185 (N_4185,N_3580,N_3687);
nor U4186 (N_4186,N_3651,N_3735);
and U4187 (N_4187,N_3597,N_3898);
and U4188 (N_4188,N_3723,N_3590);
and U4189 (N_4189,N_3708,N_3517);
or U4190 (N_4190,N_3878,N_3673);
nand U4191 (N_4191,N_3527,N_3783);
or U4192 (N_4192,N_3647,N_3933);
or U4193 (N_4193,N_3578,N_3640);
nor U4194 (N_4194,N_3750,N_3972);
or U4195 (N_4195,N_3978,N_3920);
and U4196 (N_4196,N_3871,N_3974);
or U4197 (N_4197,N_3528,N_3710);
and U4198 (N_4198,N_3631,N_3820);
nor U4199 (N_4199,N_3738,N_3726);
or U4200 (N_4200,N_3779,N_3813);
or U4201 (N_4201,N_3620,N_3888);
and U4202 (N_4202,N_3549,N_3615);
nand U4203 (N_4203,N_3809,N_3743);
and U4204 (N_4204,N_3903,N_3657);
nor U4205 (N_4205,N_3836,N_3959);
or U4206 (N_4206,N_3858,N_3834);
nand U4207 (N_4207,N_3915,N_3534);
or U4208 (N_4208,N_3532,N_3521);
and U4209 (N_4209,N_3659,N_3733);
nor U4210 (N_4210,N_3924,N_3672);
or U4211 (N_4211,N_3787,N_3988);
nand U4212 (N_4212,N_3939,N_3617);
nand U4213 (N_4213,N_3514,N_3552);
nor U4214 (N_4214,N_3857,N_3769);
nor U4215 (N_4215,N_3757,N_3967);
and U4216 (N_4216,N_3697,N_3919);
or U4217 (N_4217,N_3553,N_3936);
and U4218 (N_4218,N_3575,N_3788);
nor U4219 (N_4219,N_3581,N_3600);
nor U4220 (N_4220,N_3940,N_3606);
or U4221 (N_4221,N_3555,N_3633);
nor U4222 (N_4222,N_3954,N_3660);
and U4223 (N_4223,N_3768,N_3760);
xor U4224 (N_4224,N_3584,N_3962);
nand U4225 (N_4225,N_3641,N_3674);
xnor U4226 (N_4226,N_3909,N_3727);
nand U4227 (N_4227,N_3996,N_3559);
or U4228 (N_4228,N_3607,N_3893);
or U4229 (N_4229,N_3729,N_3875);
xnor U4230 (N_4230,N_3791,N_3646);
nand U4231 (N_4231,N_3670,N_3771);
and U4232 (N_4232,N_3583,N_3842);
nor U4233 (N_4233,N_3604,N_3975);
xor U4234 (N_4234,N_3815,N_3951);
nand U4235 (N_4235,N_3930,N_3753);
and U4236 (N_4236,N_3592,N_3781);
and U4237 (N_4237,N_3853,N_3762);
and U4238 (N_4238,N_3680,N_3950);
nand U4239 (N_4239,N_3637,N_3759);
or U4240 (N_4240,N_3642,N_3745);
nor U4241 (N_4241,N_3935,N_3795);
and U4242 (N_4242,N_3797,N_3571);
and U4243 (N_4243,N_3899,N_3560);
and U4244 (N_4244,N_3832,N_3536);
nor U4245 (N_4245,N_3694,N_3535);
and U4246 (N_4246,N_3643,N_3843);
or U4247 (N_4247,N_3565,N_3765);
or U4248 (N_4248,N_3737,N_3684);
and U4249 (N_4249,N_3546,N_3526);
or U4250 (N_4250,N_3936,N_3858);
nand U4251 (N_4251,N_3916,N_3748);
nand U4252 (N_4252,N_3626,N_3789);
nand U4253 (N_4253,N_3832,N_3719);
nor U4254 (N_4254,N_3992,N_3719);
or U4255 (N_4255,N_3629,N_3571);
or U4256 (N_4256,N_3702,N_3510);
or U4257 (N_4257,N_3607,N_3939);
nand U4258 (N_4258,N_3616,N_3506);
nand U4259 (N_4259,N_3900,N_3798);
nor U4260 (N_4260,N_3688,N_3507);
nand U4261 (N_4261,N_3567,N_3838);
and U4262 (N_4262,N_3503,N_3878);
nand U4263 (N_4263,N_3942,N_3829);
nand U4264 (N_4264,N_3905,N_3742);
nor U4265 (N_4265,N_3670,N_3900);
nor U4266 (N_4266,N_3954,N_3605);
nor U4267 (N_4267,N_3883,N_3501);
xor U4268 (N_4268,N_3885,N_3833);
or U4269 (N_4269,N_3909,N_3640);
and U4270 (N_4270,N_3851,N_3670);
nand U4271 (N_4271,N_3828,N_3665);
nor U4272 (N_4272,N_3955,N_3946);
and U4273 (N_4273,N_3958,N_3551);
and U4274 (N_4274,N_3717,N_3839);
and U4275 (N_4275,N_3774,N_3687);
xnor U4276 (N_4276,N_3687,N_3890);
nand U4277 (N_4277,N_3690,N_3789);
xnor U4278 (N_4278,N_3825,N_3501);
and U4279 (N_4279,N_3518,N_3751);
and U4280 (N_4280,N_3625,N_3893);
nor U4281 (N_4281,N_3656,N_3785);
or U4282 (N_4282,N_3979,N_3816);
nor U4283 (N_4283,N_3972,N_3708);
nand U4284 (N_4284,N_3901,N_3576);
nor U4285 (N_4285,N_3810,N_3958);
nor U4286 (N_4286,N_3566,N_3741);
or U4287 (N_4287,N_3511,N_3896);
and U4288 (N_4288,N_3961,N_3523);
nand U4289 (N_4289,N_3996,N_3827);
and U4290 (N_4290,N_3858,N_3896);
and U4291 (N_4291,N_3532,N_3591);
and U4292 (N_4292,N_3550,N_3703);
or U4293 (N_4293,N_3845,N_3809);
nor U4294 (N_4294,N_3876,N_3905);
nor U4295 (N_4295,N_3632,N_3605);
and U4296 (N_4296,N_3519,N_3602);
nor U4297 (N_4297,N_3809,N_3744);
nor U4298 (N_4298,N_3929,N_3870);
and U4299 (N_4299,N_3975,N_3761);
or U4300 (N_4300,N_3508,N_3832);
and U4301 (N_4301,N_3657,N_3634);
nand U4302 (N_4302,N_3878,N_3725);
nand U4303 (N_4303,N_3837,N_3924);
or U4304 (N_4304,N_3545,N_3881);
nor U4305 (N_4305,N_3875,N_3893);
nand U4306 (N_4306,N_3709,N_3630);
or U4307 (N_4307,N_3746,N_3976);
nand U4308 (N_4308,N_3538,N_3804);
nand U4309 (N_4309,N_3541,N_3824);
nand U4310 (N_4310,N_3789,N_3817);
nand U4311 (N_4311,N_3557,N_3909);
and U4312 (N_4312,N_3536,N_3627);
nand U4313 (N_4313,N_3770,N_3519);
nor U4314 (N_4314,N_3649,N_3559);
or U4315 (N_4315,N_3549,N_3617);
nand U4316 (N_4316,N_3759,N_3714);
nand U4317 (N_4317,N_3586,N_3603);
or U4318 (N_4318,N_3730,N_3849);
or U4319 (N_4319,N_3567,N_3882);
or U4320 (N_4320,N_3963,N_3572);
nand U4321 (N_4321,N_3718,N_3607);
and U4322 (N_4322,N_3639,N_3727);
nor U4323 (N_4323,N_3609,N_3720);
and U4324 (N_4324,N_3563,N_3790);
and U4325 (N_4325,N_3754,N_3951);
and U4326 (N_4326,N_3643,N_3584);
and U4327 (N_4327,N_3841,N_3552);
nor U4328 (N_4328,N_3792,N_3838);
nor U4329 (N_4329,N_3613,N_3840);
xnor U4330 (N_4330,N_3912,N_3979);
nand U4331 (N_4331,N_3509,N_3576);
or U4332 (N_4332,N_3528,N_3561);
and U4333 (N_4333,N_3772,N_3614);
or U4334 (N_4334,N_3850,N_3641);
nand U4335 (N_4335,N_3663,N_3618);
nand U4336 (N_4336,N_3668,N_3955);
or U4337 (N_4337,N_3859,N_3520);
and U4338 (N_4338,N_3998,N_3715);
or U4339 (N_4339,N_3939,N_3754);
and U4340 (N_4340,N_3593,N_3802);
nand U4341 (N_4341,N_3973,N_3968);
or U4342 (N_4342,N_3972,N_3710);
or U4343 (N_4343,N_3692,N_3665);
nand U4344 (N_4344,N_3553,N_3598);
nand U4345 (N_4345,N_3649,N_3536);
and U4346 (N_4346,N_3696,N_3506);
nor U4347 (N_4347,N_3795,N_3503);
and U4348 (N_4348,N_3669,N_3553);
xor U4349 (N_4349,N_3637,N_3908);
and U4350 (N_4350,N_3859,N_3870);
nand U4351 (N_4351,N_3965,N_3871);
xor U4352 (N_4352,N_3808,N_3619);
and U4353 (N_4353,N_3964,N_3773);
or U4354 (N_4354,N_3660,N_3650);
and U4355 (N_4355,N_3864,N_3692);
nand U4356 (N_4356,N_3648,N_3949);
or U4357 (N_4357,N_3605,N_3653);
xor U4358 (N_4358,N_3815,N_3702);
and U4359 (N_4359,N_3866,N_3707);
nor U4360 (N_4360,N_3964,N_3998);
and U4361 (N_4361,N_3813,N_3733);
and U4362 (N_4362,N_3864,N_3632);
and U4363 (N_4363,N_3948,N_3586);
nand U4364 (N_4364,N_3773,N_3959);
and U4365 (N_4365,N_3894,N_3583);
and U4366 (N_4366,N_3819,N_3808);
nor U4367 (N_4367,N_3800,N_3995);
or U4368 (N_4368,N_3699,N_3749);
and U4369 (N_4369,N_3769,N_3773);
and U4370 (N_4370,N_3513,N_3526);
xor U4371 (N_4371,N_3578,N_3776);
and U4372 (N_4372,N_3588,N_3936);
and U4373 (N_4373,N_3918,N_3864);
nand U4374 (N_4374,N_3606,N_3693);
nor U4375 (N_4375,N_3709,N_3892);
nand U4376 (N_4376,N_3625,N_3635);
xnor U4377 (N_4377,N_3955,N_3940);
nor U4378 (N_4378,N_3913,N_3863);
nand U4379 (N_4379,N_3876,N_3626);
nand U4380 (N_4380,N_3523,N_3896);
nand U4381 (N_4381,N_3591,N_3781);
nand U4382 (N_4382,N_3578,N_3714);
nor U4383 (N_4383,N_3818,N_3588);
and U4384 (N_4384,N_3753,N_3932);
and U4385 (N_4385,N_3793,N_3971);
nor U4386 (N_4386,N_3694,N_3556);
nor U4387 (N_4387,N_3656,N_3776);
and U4388 (N_4388,N_3540,N_3562);
xnor U4389 (N_4389,N_3810,N_3908);
nor U4390 (N_4390,N_3771,N_3921);
or U4391 (N_4391,N_3591,N_3730);
nand U4392 (N_4392,N_3562,N_3753);
xor U4393 (N_4393,N_3865,N_3798);
nor U4394 (N_4394,N_3743,N_3547);
nor U4395 (N_4395,N_3825,N_3993);
and U4396 (N_4396,N_3973,N_3665);
nand U4397 (N_4397,N_3653,N_3954);
and U4398 (N_4398,N_3703,N_3875);
or U4399 (N_4399,N_3641,N_3604);
nor U4400 (N_4400,N_3707,N_3649);
nand U4401 (N_4401,N_3722,N_3645);
nor U4402 (N_4402,N_3983,N_3672);
and U4403 (N_4403,N_3511,N_3594);
or U4404 (N_4404,N_3682,N_3555);
xor U4405 (N_4405,N_3722,N_3913);
nand U4406 (N_4406,N_3789,N_3720);
nor U4407 (N_4407,N_3818,N_3920);
nand U4408 (N_4408,N_3959,N_3821);
nor U4409 (N_4409,N_3560,N_3611);
nand U4410 (N_4410,N_3500,N_3908);
nor U4411 (N_4411,N_3915,N_3807);
nor U4412 (N_4412,N_3515,N_3837);
nand U4413 (N_4413,N_3895,N_3835);
xnor U4414 (N_4414,N_3928,N_3552);
or U4415 (N_4415,N_3589,N_3506);
and U4416 (N_4416,N_3755,N_3592);
or U4417 (N_4417,N_3938,N_3523);
xnor U4418 (N_4418,N_3514,N_3767);
or U4419 (N_4419,N_3976,N_3609);
and U4420 (N_4420,N_3736,N_3888);
or U4421 (N_4421,N_3935,N_3709);
nor U4422 (N_4422,N_3702,N_3937);
nor U4423 (N_4423,N_3566,N_3638);
nand U4424 (N_4424,N_3837,N_3623);
nand U4425 (N_4425,N_3751,N_3883);
and U4426 (N_4426,N_3583,N_3777);
and U4427 (N_4427,N_3745,N_3681);
nor U4428 (N_4428,N_3894,N_3738);
nand U4429 (N_4429,N_3905,N_3680);
nor U4430 (N_4430,N_3596,N_3631);
nor U4431 (N_4431,N_3920,N_3604);
or U4432 (N_4432,N_3852,N_3627);
and U4433 (N_4433,N_3775,N_3885);
nand U4434 (N_4434,N_3615,N_3885);
and U4435 (N_4435,N_3500,N_3903);
nand U4436 (N_4436,N_3541,N_3991);
nor U4437 (N_4437,N_3512,N_3541);
and U4438 (N_4438,N_3992,N_3984);
nor U4439 (N_4439,N_3723,N_3703);
or U4440 (N_4440,N_3641,N_3687);
or U4441 (N_4441,N_3597,N_3648);
nor U4442 (N_4442,N_3867,N_3626);
xnor U4443 (N_4443,N_3966,N_3964);
xor U4444 (N_4444,N_3507,N_3793);
or U4445 (N_4445,N_3871,N_3841);
nor U4446 (N_4446,N_3591,N_3641);
nand U4447 (N_4447,N_3804,N_3544);
nor U4448 (N_4448,N_3613,N_3863);
or U4449 (N_4449,N_3669,N_3970);
nand U4450 (N_4450,N_3932,N_3611);
xor U4451 (N_4451,N_3522,N_3833);
nor U4452 (N_4452,N_3793,N_3919);
nand U4453 (N_4453,N_3787,N_3575);
xnor U4454 (N_4454,N_3914,N_3897);
and U4455 (N_4455,N_3748,N_3654);
nor U4456 (N_4456,N_3958,N_3878);
or U4457 (N_4457,N_3951,N_3592);
and U4458 (N_4458,N_3696,N_3848);
and U4459 (N_4459,N_3591,N_3550);
or U4460 (N_4460,N_3687,N_3809);
nor U4461 (N_4461,N_3582,N_3947);
or U4462 (N_4462,N_3999,N_3692);
nand U4463 (N_4463,N_3734,N_3980);
xnor U4464 (N_4464,N_3665,N_3708);
or U4465 (N_4465,N_3562,N_3589);
xor U4466 (N_4466,N_3718,N_3991);
xnor U4467 (N_4467,N_3810,N_3808);
nor U4468 (N_4468,N_3614,N_3662);
nand U4469 (N_4469,N_3953,N_3649);
nand U4470 (N_4470,N_3644,N_3722);
and U4471 (N_4471,N_3913,N_3697);
nand U4472 (N_4472,N_3801,N_3713);
nand U4473 (N_4473,N_3948,N_3817);
and U4474 (N_4474,N_3639,N_3965);
nor U4475 (N_4475,N_3904,N_3806);
or U4476 (N_4476,N_3609,N_3918);
nand U4477 (N_4477,N_3524,N_3716);
nor U4478 (N_4478,N_3945,N_3657);
xor U4479 (N_4479,N_3746,N_3850);
xor U4480 (N_4480,N_3885,N_3584);
nand U4481 (N_4481,N_3816,N_3865);
and U4482 (N_4482,N_3662,N_3602);
and U4483 (N_4483,N_3800,N_3716);
and U4484 (N_4484,N_3851,N_3502);
and U4485 (N_4485,N_3897,N_3908);
xnor U4486 (N_4486,N_3810,N_3815);
nor U4487 (N_4487,N_3762,N_3926);
or U4488 (N_4488,N_3969,N_3584);
and U4489 (N_4489,N_3863,N_3536);
nand U4490 (N_4490,N_3800,N_3734);
xnor U4491 (N_4491,N_3947,N_3517);
and U4492 (N_4492,N_3806,N_3675);
or U4493 (N_4493,N_3875,N_3836);
and U4494 (N_4494,N_3767,N_3947);
nand U4495 (N_4495,N_3618,N_3840);
nand U4496 (N_4496,N_3518,N_3682);
nor U4497 (N_4497,N_3855,N_3827);
nor U4498 (N_4498,N_3894,N_3631);
or U4499 (N_4499,N_3857,N_3638);
nor U4500 (N_4500,N_4048,N_4148);
nand U4501 (N_4501,N_4214,N_4140);
nand U4502 (N_4502,N_4345,N_4392);
xor U4503 (N_4503,N_4394,N_4313);
nor U4504 (N_4504,N_4248,N_4473);
or U4505 (N_4505,N_4360,N_4421);
nor U4506 (N_4506,N_4478,N_4070);
nor U4507 (N_4507,N_4013,N_4151);
nand U4508 (N_4508,N_4194,N_4146);
nor U4509 (N_4509,N_4073,N_4352);
or U4510 (N_4510,N_4293,N_4449);
and U4511 (N_4511,N_4155,N_4098);
xnor U4512 (N_4512,N_4351,N_4285);
and U4513 (N_4513,N_4016,N_4408);
nor U4514 (N_4514,N_4259,N_4290);
or U4515 (N_4515,N_4482,N_4172);
and U4516 (N_4516,N_4128,N_4284);
nor U4517 (N_4517,N_4252,N_4244);
nand U4518 (N_4518,N_4420,N_4493);
and U4519 (N_4519,N_4275,N_4471);
or U4520 (N_4520,N_4491,N_4231);
xnor U4521 (N_4521,N_4496,N_4350);
nor U4522 (N_4522,N_4370,N_4440);
nand U4523 (N_4523,N_4156,N_4029);
and U4524 (N_4524,N_4122,N_4355);
nand U4525 (N_4525,N_4267,N_4383);
nor U4526 (N_4526,N_4365,N_4183);
nor U4527 (N_4527,N_4340,N_4165);
or U4528 (N_4528,N_4095,N_4233);
nand U4529 (N_4529,N_4387,N_4154);
and U4530 (N_4530,N_4230,N_4141);
nor U4531 (N_4531,N_4067,N_4356);
or U4532 (N_4532,N_4081,N_4288);
and U4533 (N_4533,N_4018,N_4242);
and U4534 (N_4534,N_4386,N_4317);
nand U4535 (N_4535,N_4437,N_4008);
xnor U4536 (N_4536,N_4260,N_4077);
and U4537 (N_4537,N_4430,N_4120);
nor U4538 (N_4538,N_4298,N_4126);
and U4539 (N_4539,N_4379,N_4470);
or U4540 (N_4540,N_4041,N_4053);
nand U4541 (N_4541,N_4031,N_4039);
nor U4542 (N_4542,N_4448,N_4058);
nand U4543 (N_4543,N_4300,N_4338);
and U4544 (N_4544,N_4218,N_4316);
nand U4545 (N_4545,N_4223,N_4204);
nor U4546 (N_4546,N_4413,N_4017);
or U4547 (N_4547,N_4467,N_4357);
xor U4548 (N_4548,N_4004,N_4475);
or U4549 (N_4549,N_4221,N_4190);
or U4550 (N_4550,N_4498,N_4159);
or U4551 (N_4551,N_4212,N_4000);
nand U4552 (N_4552,N_4363,N_4377);
xor U4553 (N_4553,N_4436,N_4101);
and U4554 (N_4554,N_4118,N_4015);
xnor U4555 (N_4555,N_4035,N_4090);
or U4556 (N_4556,N_4005,N_4184);
and U4557 (N_4557,N_4001,N_4219);
or U4558 (N_4558,N_4033,N_4265);
or U4559 (N_4559,N_4270,N_4395);
or U4560 (N_4560,N_4235,N_4264);
nor U4561 (N_4561,N_4237,N_4331);
or U4562 (N_4562,N_4036,N_4393);
nand U4563 (N_4563,N_4157,N_4220);
and U4564 (N_4564,N_4411,N_4400);
nand U4565 (N_4565,N_4132,N_4086);
nand U4566 (N_4566,N_4339,N_4424);
nor U4567 (N_4567,N_4176,N_4245);
nor U4568 (N_4568,N_4150,N_4450);
or U4569 (N_4569,N_4243,N_4385);
nand U4570 (N_4570,N_4100,N_4107);
nor U4571 (N_4571,N_4232,N_4434);
nand U4572 (N_4572,N_4324,N_4181);
or U4573 (N_4573,N_4401,N_4366);
and U4574 (N_4574,N_4320,N_4404);
nand U4575 (N_4575,N_4346,N_4113);
or U4576 (N_4576,N_4145,N_4104);
nor U4577 (N_4577,N_4341,N_4037);
nand U4578 (N_4578,N_4326,N_4205);
and U4579 (N_4579,N_4251,N_4342);
nand U4580 (N_4580,N_4089,N_4144);
xnor U4581 (N_4581,N_4291,N_4179);
and U4582 (N_4582,N_4314,N_4359);
and U4583 (N_4583,N_4091,N_4410);
nand U4584 (N_4584,N_4207,N_4382);
nor U4585 (N_4585,N_4397,N_4225);
nor U4586 (N_4586,N_4097,N_4065);
or U4587 (N_4587,N_4398,N_4301);
or U4588 (N_4588,N_4047,N_4201);
and U4589 (N_4589,N_4289,N_4389);
nor U4590 (N_4590,N_4076,N_4419);
and U4591 (N_4591,N_4011,N_4453);
or U4592 (N_4592,N_4373,N_4049);
nand U4593 (N_4593,N_4136,N_4315);
and U4594 (N_4594,N_4364,N_4380);
xnor U4595 (N_4595,N_4173,N_4038);
and U4596 (N_4596,N_4280,N_4294);
nor U4597 (N_4597,N_4472,N_4337);
xnor U4598 (N_4598,N_4147,N_4149);
and U4599 (N_4599,N_4152,N_4188);
xnor U4600 (N_4600,N_4217,N_4202);
nand U4601 (N_4601,N_4481,N_4353);
nor U4602 (N_4602,N_4403,N_4269);
nor U4603 (N_4603,N_4348,N_4480);
and U4604 (N_4604,N_4461,N_4307);
nand U4605 (N_4605,N_4130,N_4323);
and U4606 (N_4606,N_4116,N_4296);
or U4607 (N_4607,N_4238,N_4465);
or U4608 (N_4608,N_4103,N_4322);
and U4609 (N_4609,N_4174,N_4131);
and U4610 (N_4610,N_4069,N_4175);
nor U4611 (N_4611,N_4329,N_4459);
nor U4612 (N_4612,N_4112,N_4192);
or U4613 (N_4613,N_4169,N_4247);
nor U4614 (N_4614,N_4186,N_4446);
or U4615 (N_4615,N_4416,N_4025);
nand U4616 (N_4616,N_4358,N_4388);
and U4617 (N_4617,N_4262,N_4479);
nand U4618 (N_4618,N_4161,N_4399);
or U4619 (N_4619,N_4158,N_4463);
xor U4620 (N_4620,N_4344,N_4312);
nand U4621 (N_4621,N_4209,N_4457);
nor U4622 (N_4622,N_4476,N_4071);
or U4623 (N_4623,N_4487,N_4052);
or U4624 (N_4624,N_4224,N_4096);
and U4625 (N_4625,N_4045,N_4414);
nand U4626 (N_4626,N_4253,N_4486);
and U4627 (N_4627,N_4299,N_4129);
or U4628 (N_4628,N_4378,N_4354);
nor U4629 (N_4629,N_4102,N_4455);
nand U4630 (N_4630,N_4497,N_4435);
nor U4631 (N_4631,N_4295,N_4425);
or U4632 (N_4632,N_4079,N_4330);
or U4633 (N_4633,N_4371,N_4203);
or U4634 (N_4634,N_4240,N_4372);
and U4635 (N_4635,N_4010,N_4111);
nor U4636 (N_4636,N_4124,N_4099);
nor U4637 (N_4637,N_4406,N_4305);
nor U4638 (N_4638,N_4271,N_4241);
nor U4639 (N_4639,N_4415,N_4279);
nand U4640 (N_4640,N_4072,N_4042);
nor U4641 (N_4641,N_4261,N_4115);
or U4642 (N_4642,N_4064,N_4046);
xor U4643 (N_4643,N_4133,N_4082);
nor U4644 (N_4644,N_4274,N_4108);
nor U4645 (N_4645,N_4423,N_4193);
and U4646 (N_4646,N_4304,N_4014);
and U4647 (N_4647,N_4164,N_4160);
and U4648 (N_4648,N_4277,N_4292);
or U4649 (N_4649,N_4327,N_4117);
nor U4650 (N_4650,N_4368,N_4211);
nor U4651 (N_4651,N_4198,N_4106);
and U4652 (N_4652,N_4075,N_4028);
nor U4653 (N_4653,N_4442,N_4443);
nor U4654 (N_4654,N_4138,N_4273);
or U4655 (N_4655,N_4412,N_4468);
or U4656 (N_4656,N_4228,N_4454);
nand U4657 (N_4657,N_4492,N_4407);
or U4658 (N_4658,N_4268,N_4068);
xnor U4659 (N_4659,N_4309,N_4061);
nor U4660 (N_4660,N_4375,N_4080);
xnor U4661 (N_4661,N_4325,N_4439);
nor U4662 (N_4662,N_4390,N_4137);
and U4663 (N_4663,N_4405,N_4417);
nand U4664 (N_4664,N_4216,N_4489);
or U4665 (N_4665,N_4032,N_4332);
or U4666 (N_4666,N_4063,N_4458);
nor U4667 (N_4667,N_4043,N_4362);
nor U4668 (N_4668,N_4376,N_4429);
nand U4669 (N_4669,N_4074,N_4433);
nand U4670 (N_4670,N_4227,N_4085);
or U4671 (N_4671,N_4059,N_4051);
and U4672 (N_4672,N_4428,N_4226);
nand U4673 (N_4673,N_4143,N_4034);
or U4674 (N_4674,N_4142,N_4056);
or U4675 (N_4675,N_4361,N_4206);
or U4676 (N_4676,N_4483,N_4427);
or U4677 (N_4677,N_4282,N_4177);
and U4678 (N_4678,N_4196,N_4283);
or U4679 (N_4679,N_4040,N_4087);
xnor U4680 (N_4680,N_4208,N_4084);
or U4681 (N_4681,N_4215,N_4418);
or U4682 (N_4682,N_4328,N_4441);
nand U4683 (N_4683,N_4066,N_4249);
nor U4684 (N_4684,N_4257,N_4006);
and U4685 (N_4685,N_4239,N_4024);
and U4686 (N_4686,N_4200,N_4134);
and U4687 (N_4687,N_4396,N_4374);
nor U4688 (N_4688,N_4431,N_4246);
xnor U4689 (N_4689,N_4027,N_4287);
nand U4690 (N_4690,N_4452,N_4191);
nor U4691 (N_4691,N_4474,N_4139);
or U4692 (N_4692,N_4255,N_4451);
nand U4693 (N_4693,N_4078,N_4162);
nand U4694 (N_4694,N_4092,N_4021);
and U4695 (N_4695,N_4445,N_4182);
nand U4696 (N_4696,N_4195,N_4499);
xnor U4697 (N_4697,N_4488,N_4409);
and U4698 (N_4698,N_4391,N_4153);
nand U4699 (N_4699,N_4187,N_4347);
and U4700 (N_4700,N_4254,N_4125);
nor U4701 (N_4701,N_4023,N_4229);
or U4702 (N_4702,N_4168,N_4306);
nand U4703 (N_4703,N_4171,N_4003);
xnor U4704 (N_4704,N_4180,N_4460);
or U4705 (N_4705,N_4197,N_4022);
nand U4706 (N_4706,N_4105,N_4222);
and U4707 (N_4707,N_4167,N_4127);
xor U4708 (N_4708,N_4057,N_4281);
xor U4709 (N_4709,N_4055,N_4485);
xor U4710 (N_4710,N_4333,N_4002);
and U4711 (N_4711,N_4121,N_4334);
nand U4712 (N_4712,N_4236,N_4319);
nor U4713 (N_4713,N_4189,N_4109);
nor U4714 (N_4714,N_4094,N_4349);
nand U4715 (N_4715,N_4213,N_4166);
nand U4716 (N_4716,N_4185,N_4447);
or U4717 (N_4717,N_4026,N_4178);
xnor U4718 (N_4718,N_4494,N_4456);
or U4719 (N_4719,N_4422,N_4367);
or U4720 (N_4720,N_4318,N_4343);
xor U4721 (N_4721,N_4266,N_4336);
nand U4722 (N_4722,N_4060,N_4114);
nor U4723 (N_4723,N_4335,N_4495);
xnor U4724 (N_4724,N_4163,N_4438);
nor U4725 (N_4725,N_4432,N_4369);
nor U4726 (N_4726,N_4250,N_4012);
nor U4727 (N_4727,N_4303,N_4278);
or U4728 (N_4728,N_4020,N_4466);
nor U4729 (N_4729,N_4384,N_4093);
or U4730 (N_4730,N_4110,N_4030);
nor U4731 (N_4731,N_4490,N_4135);
nor U4732 (N_4732,N_4381,N_4286);
nand U4733 (N_4733,N_4234,N_4302);
nor U4734 (N_4734,N_4019,N_4321);
and U4735 (N_4735,N_4007,N_4054);
xor U4736 (N_4736,N_4402,N_4123);
or U4737 (N_4737,N_4308,N_4050);
xnor U4738 (N_4738,N_4272,N_4083);
xnor U4739 (N_4739,N_4199,N_4464);
and U4740 (N_4740,N_4210,N_4119);
nor U4741 (N_4741,N_4062,N_4462);
and U4742 (N_4742,N_4258,N_4484);
nand U4743 (N_4743,N_4444,N_4297);
nand U4744 (N_4744,N_4256,N_4263);
and U4745 (N_4745,N_4310,N_4044);
nor U4746 (N_4746,N_4276,N_4170);
nand U4747 (N_4747,N_4477,N_4311);
or U4748 (N_4748,N_4469,N_4088);
and U4749 (N_4749,N_4426,N_4009);
or U4750 (N_4750,N_4498,N_4365);
or U4751 (N_4751,N_4182,N_4188);
and U4752 (N_4752,N_4468,N_4244);
nand U4753 (N_4753,N_4161,N_4216);
and U4754 (N_4754,N_4481,N_4162);
nand U4755 (N_4755,N_4007,N_4405);
or U4756 (N_4756,N_4047,N_4078);
xor U4757 (N_4757,N_4102,N_4376);
xnor U4758 (N_4758,N_4199,N_4010);
or U4759 (N_4759,N_4419,N_4455);
or U4760 (N_4760,N_4106,N_4072);
nor U4761 (N_4761,N_4064,N_4304);
or U4762 (N_4762,N_4304,N_4000);
and U4763 (N_4763,N_4065,N_4113);
nand U4764 (N_4764,N_4148,N_4096);
and U4765 (N_4765,N_4339,N_4241);
nand U4766 (N_4766,N_4449,N_4401);
nor U4767 (N_4767,N_4198,N_4111);
nor U4768 (N_4768,N_4324,N_4242);
nand U4769 (N_4769,N_4379,N_4154);
or U4770 (N_4770,N_4321,N_4026);
xor U4771 (N_4771,N_4192,N_4185);
nand U4772 (N_4772,N_4369,N_4230);
or U4773 (N_4773,N_4360,N_4150);
or U4774 (N_4774,N_4435,N_4175);
nor U4775 (N_4775,N_4070,N_4046);
nand U4776 (N_4776,N_4451,N_4209);
or U4777 (N_4777,N_4484,N_4363);
or U4778 (N_4778,N_4464,N_4339);
nor U4779 (N_4779,N_4341,N_4145);
or U4780 (N_4780,N_4328,N_4036);
and U4781 (N_4781,N_4005,N_4171);
nand U4782 (N_4782,N_4026,N_4171);
xor U4783 (N_4783,N_4023,N_4295);
nor U4784 (N_4784,N_4028,N_4045);
and U4785 (N_4785,N_4038,N_4246);
xnor U4786 (N_4786,N_4415,N_4106);
nand U4787 (N_4787,N_4282,N_4221);
and U4788 (N_4788,N_4217,N_4435);
and U4789 (N_4789,N_4203,N_4080);
and U4790 (N_4790,N_4404,N_4381);
and U4791 (N_4791,N_4339,N_4038);
nand U4792 (N_4792,N_4151,N_4102);
or U4793 (N_4793,N_4387,N_4315);
or U4794 (N_4794,N_4441,N_4266);
nor U4795 (N_4795,N_4424,N_4146);
or U4796 (N_4796,N_4083,N_4121);
xnor U4797 (N_4797,N_4466,N_4364);
nand U4798 (N_4798,N_4235,N_4056);
and U4799 (N_4799,N_4489,N_4034);
and U4800 (N_4800,N_4209,N_4387);
nand U4801 (N_4801,N_4410,N_4196);
xnor U4802 (N_4802,N_4025,N_4262);
and U4803 (N_4803,N_4061,N_4224);
or U4804 (N_4804,N_4266,N_4326);
nand U4805 (N_4805,N_4049,N_4164);
nor U4806 (N_4806,N_4447,N_4433);
or U4807 (N_4807,N_4097,N_4397);
or U4808 (N_4808,N_4345,N_4385);
nand U4809 (N_4809,N_4305,N_4317);
and U4810 (N_4810,N_4376,N_4049);
nand U4811 (N_4811,N_4475,N_4188);
nor U4812 (N_4812,N_4462,N_4008);
nor U4813 (N_4813,N_4462,N_4234);
nor U4814 (N_4814,N_4388,N_4080);
nand U4815 (N_4815,N_4311,N_4258);
nor U4816 (N_4816,N_4228,N_4313);
nor U4817 (N_4817,N_4496,N_4448);
or U4818 (N_4818,N_4130,N_4484);
and U4819 (N_4819,N_4382,N_4100);
xnor U4820 (N_4820,N_4181,N_4317);
nand U4821 (N_4821,N_4026,N_4080);
or U4822 (N_4822,N_4123,N_4378);
nor U4823 (N_4823,N_4425,N_4167);
and U4824 (N_4824,N_4414,N_4287);
and U4825 (N_4825,N_4270,N_4250);
nand U4826 (N_4826,N_4375,N_4461);
nand U4827 (N_4827,N_4426,N_4021);
nand U4828 (N_4828,N_4167,N_4280);
and U4829 (N_4829,N_4063,N_4125);
nand U4830 (N_4830,N_4114,N_4253);
nor U4831 (N_4831,N_4453,N_4115);
nand U4832 (N_4832,N_4440,N_4196);
or U4833 (N_4833,N_4051,N_4230);
and U4834 (N_4834,N_4222,N_4316);
and U4835 (N_4835,N_4342,N_4052);
nand U4836 (N_4836,N_4063,N_4427);
nor U4837 (N_4837,N_4340,N_4058);
nand U4838 (N_4838,N_4455,N_4325);
xor U4839 (N_4839,N_4187,N_4102);
nor U4840 (N_4840,N_4029,N_4354);
nand U4841 (N_4841,N_4380,N_4273);
and U4842 (N_4842,N_4153,N_4278);
or U4843 (N_4843,N_4395,N_4052);
nor U4844 (N_4844,N_4086,N_4325);
and U4845 (N_4845,N_4214,N_4204);
and U4846 (N_4846,N_4342,N_4362);
nor U4847 (N_4847,N_4430,N_4391);
nor U4848 (N_4848,N_4314,N_4021);
nand U4849 (N_4849,N_4123,N_4167);
nor U4850 (N_4850,N_4256,N_4305);
or U4851 (N_4851,N_4482,N_4248);
or U4852 (N_4852,N_4012,N_4226);
nand U4853 (N_4853,N_4155,N_4043);
nor U4854 (N_4854,N_4233,N_4213);
or U4855 (N_4855,N_4136,N_4214);
xnor U4856 (N_4856,N_4437,N_4050);
xor U4857 (N_4857,N_4355,N_4385);
or U4858 (N_4858,N_4193,N_4166);
xnor U4859 (N_4859,N_4325,N_4303);
and U4860 (N_4860,N_4425,N_4045);
nand U4861 (N_4861,N_4465,N_4468);
nand U4862 (N_4862,N_4023,N_4185);
nand U4863 (N_4863,N_4437,N_4156);
nand U4864 (N_4864,N_4288,N_4000);
nand U4865 (N_4865,N_4022,N_4337);
nor U4866 (N_4866,N_4414,N_4485);
nand U4867 (N_4867,N_4221,N_4187);
nand U4868 (N_4868,N_4464,N_4232);
or U4869 (N_4869,N_4176,N_4387);
nand U4870 (N_4870,N_4048,N_4168);
and U4871 (N_4871,N_4006,N_4437);
nand U4872 (N_4872,N_4423,N_4335);
nor U4873 (N_4873,N_4492,N_4190);
nand U4874 (N_4874,N_4065,N_4199);
or U4875 (N_4875,N_4338,N_4320);
or U4876 (N_4876,N_4329,N_4008);
nand U4877 (N_4877,N_4099,N_4366);
or U4878 (N_4878,N_4009,N_4215);
xnor U4879 (N_4879,N_4202,N_4084);
and U4880 (N_4880,N_4346,N_4175);
nor U4881 (N_4881,N_4183,N_4218);
or U4882 (N_4882,N_4290,N_4170);
xor U4883 (N_4883,N_4098,N_4456);
nor U4884 (N_4884,N_4326,N_4237);
nor U4885 (N_4885,N_4405,N_4002);
nand U4886 (N_4886,N_4246,N_4496);
and U4887 (N_4887,N_4006,N_4145);
or U4888 (N_4888,N_4002,N_4345);
or U4889 (N_4889,N_4411,N_4236);
nand U4890 (N_4890,N_4186,N_4001);
or U4891 (N_4891,N_4176,N_4131);
xnor U4892 (N_4892,N_4463,N_4476);
xnor U4893 (N_4893,N_4336,N_4153);
and U4894 (N_4894,N_4472,N_4075);
nand U4895 (N_4895,N_4075,N_4366);
nor U4896 (N_4896,N_4491,N_4465);
nand U4897 (N_4897,N_4210,N_4442);
xnor U4898 (N_4898,N_4334,N_4257);
nand U4899 (N_4899,N_4025,N_4067);
xnor U4900 (N_4900,N_4436,N_4304);
nor U4901 (N_4901,N_4025,N_4028);
nand U4902 (N_4902,N_4001,N_4180);
or U4903 (N_4903,N_4087,N_4445);
or U4904 (N_4904,N_4176,N_4449);
nand U4905 (N_4905,N_4399,N_4009);
or U4906 (N_4906,N_4310,N_4222);
nand U4907 (N_4907,N_4372,N_4237);
nand U4908 (N_4908,N_4194,N_4149);
nor U4909 (N_4909,N_4393,N_4141);
or U4910 (N_4910,N_4266,N_4309);
or U4911 (N_4911,N_4075,N_4142);
or U4912 (N_4912,N_4258,N_4337);
nor U4913 (N_4913,N_4492,N_4012);
or U4914 (N_4914,N_4330,N_4443);
nor U4915 (N_4915,N_4134,N_4480);
nand U4916 (N_4916,N_4130,N_4380);
xor U4917 (N_4917,N_4130,N_4240);
nor U4918 (N_4918,N_4331,N_4012);
nor U4919 (N_4919,N_4261,N_4429);
xor U4920 (N_4920,N_4271,N_4136);
or U4921 (N_4921,N_4040,N_4396);
xor U4922 (N_4922,N_4164,N_4440);
or U4923 (N_4923,N_4096,N_4073);
nand U4924 (N_4924,N_4289,N_4382);
xnor U4925 (N_4925,N_4428,N_4145);
or U4926 (N_4926,N_4356,N_4035);
and U4927 (N_4927,N_4494,N_4153);
or U4928 (N_4928,N_4299,N_4081);
or U4929 (N_4929,N_4275,N_4186);
or U4930 (N_4930,N_4210,N_4255);
and U4931 (N_4931,N_4014,N_4116);
nor U4932 (N_4932,N_4285,N_4450);
nand U4933 (N_4933,N_4051,N_4078);
and U4934 (N_4934,N_4440,N_4193);
and U4935 (N_4935,N_4074,N_4391);
or U4936 (N_4936,N_4038,N_4220);
nand U4937 (N_4937,N_4130,N_4175);
and U4938 (N_4938,N_4470,N_4120);
and U4939 (N_4939,N_4224,N_4484);
xnor U4940 (N_4940,N_4470,N_4038);
xor U4941 (N_4941,N_4201,N_4203);
or U4942 (N_4942,N_4202,N_4034);
nand U4943 (N_4943,N_4214,N_4032);
nand U4944 (N_4944,N_4145,N_4297);
nor U4945 (N_4945,N_4230,N_4346);
nor U4946 (N_4946,N_4251,N_4420);
or U4947 (N_4947,N_4280,N_4479);
and U4948 (N_4948,N_4248,N_4289);
or U4949 (N_4949,N_4444,N_4436);
nor U4950 (N_4950,N_4211,N_4099);
and U4951 (N_4951,N_4358,N_4313);
and U4952 (N_4952,N_4141,N_4104);
and U4953 (N_4953,N_4358,N_4258);
and U4954 (N_4954,N_4056,N_4083);
or U4955 (N_4955,N_4360,N_4030);
nand U4956 (N_4956,N_4394,N_4323);
nand U4957 (N_4957,N_4470,N_4481);
or U4958 (N_4958,N_4461,N_4211);
nor U4959 (N_4959,N_4298,N_4027);
nor U4960 (N_4960,N_4302,N_4205);
or U4961 (N_4961,N_4474,N_4271);
or U4962 (N_4962,N_4439,N_4458);
xnor U4963 (N_4963,N_4469,N_4391);
nor U4964 (N_4964,N_4290,N_4000);
nand U4965 (N_4965,N_4216,N_4201);
and U4966 (N_4966,N_4445,N_4346);
or U4967 (N_4967,N_4431,N_4170);
and U4968 (N_4968,N_4469,N_4195);
nand U4969 (N_4969,N_4467,N_4111);
and U4970 (N_4970,N_4484,N_4320);
and U4971 (N_4971,N_4176,N_4309);
nor U4972 (N_4972,N_4262,N_4460);
nor U4973 (N_4973,N_4424,N_4357);
nand U4974 (N_4974,N_4168,N_4004);
and U4975 (N_4975,N_4001,N_4422);
nor U4976 (N_4976,N_4298,N_4363);
xor U4977 (N_4977,N_4197,N_4331);
nand U4978 (N_4978,N_4119,N_4124);
nor U4979 (N_4979,N_4069,N_4343);
nand U4980 (N_4980,N_4366,N_4441);
nand U4981 (N_4981,N_4394,N_4023);
nor U4982 (N_4982,N_4383,N_4059);
or U4983 (N_4983,N_4354,N_4073);
and U4984 (N_4984,N_4244,N_4262);
nor U4985 (N_4985,N_4225,N_4074);
and U4986 (N_4986,N_4060,N_4077);
and U4987 (N_4987,N_4272,N_4200);
and U4988 (N_4988,N_4150,N_4036);
or U4989 (N_4989,N_4222,N_4296);
nand U4990 (N_4990,N_4244,N_4090);
and U4991 (N_4991,N_4480,N_4265);
nor U4992 (N_4992,N_4168,N_4060);
or U4993 (N_4993,N_4231,N_4235);
nand U4994 (N_4994,N_4177,N_4397);
nand U4995 (N_4995,N_4139,N_4479);
nand U4996 (N_4996,N_4298,N_4391);
and U4997 (N_4997,N_4015,N_4052);
and U4998 (N_4998,N_4355,N_4437);
and U4999 (N_4999,N_4349,N_4027);
and U5000 (N_5000,N_4721,N_4623);
and U5001 (N_5001,N_4634,N_4819);
nor U5002 (N_5002,N_4692,N_4504);
or U5003 (N_5003,N_4982,N_4562);
nand U5004 (N_5004,N_4963,N_4851);
nor U5005 (N_5005,N_4635,N_4994);
nand U5006 (N_5006,N_4974,N_4538);
or U5007 (N_5007,N_4732,N_4840);
and U5008 (N_5008,N_4603,N_4768);
nor U5009 (N_5009,N_4655,N_4886);
xor U5010 (N_5010,N_4565,N_4845);
or U5011 (N_5011,N_4854,N_4910);
or U5012 (N_5012,N_4563,N_4642);
xor U5013 (N_5013,N_4546,N_4570);
or U5014 (N_5014,N_4696,N_4700);
nor U5015 (N_5015,N_4584,N_4810);
and U5016 (N_5016,N_4615,N_4531);
and U5017 (N_5017,N_4956,N_4961);
and U5018 (N_5018,N_4764,N_4806);
nor U5019 (N_5019,N_4697,N_4580);
xnor U5020 (N_5020,N_4748,N_4751);
nand U5021 (N_5021,N_4761,N_4835);
or U5022 (N_5022,N_4646,N_4526);
or U5023 (N_5023,N_4632,N_4863);
nor U5024 (N_5024,N_4871,N_4979);
nand U5025 (N_5025,N_4657,N_4682);
and U5026 (N_5026,N_4596,N_4970);
nor U5027 (N_5027,N_4532,N_4985);
nor U5028 (N_5028,N_4541,N_4849);
and U5029 (N_5029,N_4966,N_4601);
nor U5030 (N_5030,N_4862,N_4540);
xor U5031 (N_5031,N_4534,N_4709);
nand U5032 (N_5032,N_4891,N_4805);
nor U5033 (N_5033,N_4576,N_4926);
or U5034 (N_5034,N_4904,N_4967);
nand U5035 (N_5035,N_4519,N_4788);
or U5036 (N_5036,N_4918,N_4989);
or U5037 (N_5037,N_4755,N_4848);
and U5038 (N_5038,N_4598,N_4801);
nor U5039 (N_5039,N_4738,N_4550);
nor U5040 (N_5040,N_4542,N_4671);
nand U5041 (N_5041,N_4830,N_4744);
or U5042 (N_5042,N_4885,N_4940);
or U5043 (N_5043,N_4828,N_4793);
nor U5044 (N_5044,N_4763,N_4503);
nand U5045 (N_5045,N_4826,N_4865);
and U5046 (N_5046,N_4633,N_4627);
nor U5047 (N_5047,N_4685,N_4586);
nor U5048 (N_5048,N_4521,N_4549);
nand U5049 (N_5049,N_4870,N_4831);
nor U5050 (N_5050,N_4752,N_4683);
nand U5051 (N_5051,N_4997,N_4593);
nor U5052 (N_5052,N_4869,N_4513);
nand U5053 (N_5053,N_4624,N_4606);
nor U5054 (N_5054,N_4759,N_4832);
nand U5055 (N_5055,N_4718,N_4781);
nand U5056 (N_5056,N_4780,N_4857);
or U5057 (N_5057,N_4592,N_4932);
nand U5058 (N_5058,N_4792,N_4686);
nor U5059 (N_5059,N_4935,N_4954);
nand U5060 (N_5060,N_4817,N_4929);
nor U5061 (N_5061,N_4607,N_4937);
nor U5062 (N_5062,N_4852,N_4548);
nand U5063 (N_5063,N_4841,N_4711);
and U5064 (N_5064,N_4557,N_4609);
nor U5065 (N_5065,N_4610,N_4585);
nand U5066 (N_5066,N_4903,N_4769);
or U5067 (N_5067,N_4799,N_4736);
nand U5068 (N_5068,N_4699,N_4790);
nand U5069 (N_5069,N_4838,N_4535);
or U5070 (N_5070,N_4500,N_4707);
or U5071 (N_5071,N_4859,N_4740);
and U5072 (N_5072,N_4803,N_4837);
nand U5073 (N_5073,N_4734,N_4706);
nand U5074 (N_5074,N_4704,N_4999);
nor U5075 (N_5075,N_4693,N_4753);
and U5076 (N_5076,N_4975,N_4778);
nand U5077 (N_5077,N_4833,N_4639);
nor U5078 (N_5078,N_4945,N_4847);
or U5079 (N_5079,N_4664,N_4583);
and U5080 (N_5080,N_4785,N_4716);
nor U5081 (N_5081,N_4813,N_4816);
nor U5082 (N_5082,N_4626,N_4992);
xor U5083 (N_5083,N_4516,N_4888);
or U5084 (N_5084,N_4743,N_4628);
or U5085 (N_5085,N_4856,N_4971);
xor U5086 (N_5086,N_4560,N_4529);
nor U5087 (N_5087,N_4976,N_4846);
nand U5088 (N_5088,N_4523,N_4795);
xor U5089 (N_5089,N_4774,N_4618);
nor U5090 (N_5090,N_4653,N_4784);
or U5091 (N_5091,N_4914,N_4578);
xnor U5092 (N_5092,N_4631,N_4812);
nor U5093 (N_5093,N_4575,N_4758);
nor U5094 (N_5094,N_4876,N_4714);
nor U5095 (N_5095,N_4561,N_4741);
and U5096 (N_5096,N_4919,N_4522);
xor U5097 (N_5097,N_4892,N_4551);
or U5098 (N_5098,N_4681,N_4501);
or U5099 (N_5099,N_4619,N_4860);
nor U5100 (N_5100,N_4511,N_4555);
and U5101 (N_5101,N_4737,N_4746);
nor U5102 (N_5102,N_4965,N_4957);
nor U5103 (N_5103,N_4951,N_4652);
nor U5104 (N_5104,N_4765,N_4977);
and U5105 (N_5105,N_4722,N_4739);
nor U5106 (N_5106,N_4648,N_4684);
nand U5107 (N_5107,N_4927,N_4938);
nor U5108 (N_5108,N_4878,N_4749);
nor U5109 (N_5109,N_4959,N_4622);
xnor U5110 (N_5110,N_4705,N_4934);
nand U5111 (N_5111,N_4782,N_4796);
and U5112 (N_5112,N_4571,N_4668);
nor U5113 (N_5113,N_4899,N_4507);
and U5114 (N_5114,N_4688,N_4595);
nor U5115 (N_5115,N_4559,N_4703);
and U5116 (N_5116,N_4553,N_4614);
nand U5117 (N_5117,N_4767,N_4656);
and U5118 (N_5118,N_4770,N_4822);
nor U5119 (N_5119,N_4530,N_4608);
nor U5120 (N_5120,N_4917,N_4829);
nand U5121 (N_5121,N_4920,N_4581);
and U5122 (N_5122,N_4930,N_4818);
nand U5123 (N_5123,N_4896,N_4771);
and U5124 (N_5124,N_4931,N_4775);
nor U5125 (N_5125,N_4510,N_4993);
or U5126 (N_5126,N_4922,N_4630);
or U5127 (N_5127,N_4777,N_4936);
or U5128 (N_5128,N_4766,N_4611);
or U5129 (N_5129,N_4990,N_4666);
and U5130 (N_5130,N_4544,N_4710);
or U5131 (N_5131,N_4789,N_4897);
nor U5132 (N_5132,N_4512,N_4539);
or U5133 (N_5133,N_4902,N_4713);
xor U5134 (N_5134,N_4514,N_4677);
and U5135 (N_5135,N_4582,N_4533);
or U5136 (N_5136,N_4811,N_4827);
and U5137 (N_5137,N_4773,N_4720);
nand U5138 (N_5138,N_4573,N_4679);
and U5139 (N_5139,N_4787,N_4660);
or U5140 (N_5140,N_4913,N_4879);
xnor U5141 (N_5141,N_4670,N_4823);
nand U5142 (N_5142,N_4698,N_4983);
nand U5143 (N_5143,N_4605,N_4745);
and U5144 (N_5144,N_4502,N_4760);
nand U5145 (N_5145,N_4733,N_4708);
nand U5146 (N_5146,N_4663,N_4800);
nand U5147 (N_5147,N_4853,N_4599);
and U5148 (N_5148,N_4928,N_4923);
and U5149 (N_5149,N_4579,N_4673);
and U5150 (N_5150,N_4941,N_4594);
nor U5151 (N_5151,N_4756,N_4536);
and U5152 (N_5152,N_4651,N_4667);
and U5153 (N_5153,N_4779,N_4636);
and U5154 (N_5154,N_4694,N_4855);
and U5155 (N_5155,N_4644,N_4729);
nand U5156 (N_5156,N_4702,N_4864);
or U5157 (N_5157,N_4872,N_4724);
or U5158 (N_5158,N_4844,N_4809);
nand U5159 (N_5159,N_4537,N_4730);
xor U5160 (N_5160,N_4695,N_4597);
or U5161 (N_5161,N_4960,N_4900);
nor U5162 (N_5162,N_4839,N_4527);
nand U5163 (N_5163,N_4807,N_4895);
or U5164 (N_5164,N_4717,N_4821);
xnor U5165 (N_5165,N_4661,N_4517);
nor U5166 (N_5166,N_4875,N_4973);
xor U5167 (N_5167,N_4617,N_4602);
and U5168 (N_5168,N_4691,N_4850);
nor U5169 (N_5169,N_4921,N_4726);
nor U5170 (N_5170,N_4794,N_4572);
nor U5171 (N_5171,N_4645,N_4890);
and U5172 (N_5172,N_4715,N_4658);
and U5173 (N_5173,N_4978,N_4647);
nand U5174 (N_5174,N_4884,N_4925);
xnor U5175 (N_5175,N_4915,N_4958);
or U5176 (N_5176,N_4554,N_4776);
nor U5177 (N_5177,N_4942,N_4727);
and U5178 (N_5178,N_4672,N_4988);
and U5179 (N_5179,N_4933,N_4556);
xor U5180 (N_5180,N_4867,N_4984);
or U5181 (N_5181,N_4909,N_4877);
nor U5182 (N_5182,N_4669,N_4612);
or U5183 (N_5183,N_4772,N_4754);
and U5184 (N_5184,N_4996,N_4986);
and U5185 (N_5185,N_4908,N_4783);
and U5186 (N_5186,N_4969,N_4883);
nor U5187 (N_5187,N_4898,N_4564);
nor U5188 (N_5188,N_4947,N_4750);
nand U5189 (N_5189,N_4843,N_4820);
and U5190 (N_5190,N_4747,N_4943);
or U5191 (N_5191,N_4620,N_4802);
and U5192 (N_5192,N_4874,N_4676);
xor U5193 (N_5193,N_4894,N_4650);
and U5194 (N_5194,N_4505,N_4728);
nor U5195 (N_5195,N_4723,N_4566);
and U5196 (N_5196,N_4604,N_4881);
and U5197 (N_5197,N_4991,N_4924);
or U5198 (N_5198,N_4613,N_4944);
and U5199 (N_5199,N_4952,N_4643);
nor U5200 (N_5200,N_4980,N_4689);
or U5201 (N_5201,N_4701,N_4757);
nand U5202 (N_5202,N_4680,N_4797);
nand U5203 (N_5203,N_4834,N_4804);
or U5204 (N_5204,N_4659,N_4880);
nand U5205 (N_5205,N_4654,N_4824);
nand U5206 (N_5206,N_4893,N_4520);
xor U5207 (N_5207,N_4836,N_4889);
nand U5208 (N_5208,N_4815,N_4616);
nand U5209 (N_5209,N_4907,N_4949);
or U5210 (N_5210,N_4825,N_4972);
nor U5211 (N_5211,N_4678,N_4662);
nand U5212 (N_5212,N_4868,N_4552);
xor U5213 (N_5213,N_4690,N_4725);
or U5214 (N_5214,N_4861,N_4791);
nor U5215 (N_5215,N_4912,N_4998);
nand U5216 (N_5216,N_4946,N_4916);
nor U5217 (N_5217,N_4950,N_4939);
or U5218 (N_5218,N_4528,N_4547);
and U5219 (N_5219,N_4962,N_4953);
nor U5220 (N_5220,N_4762,N_4808);
and U5221 (N_5221,N_4509,N_4687);
nor U5222 (N_5222,N_4590,N_4866);
nand U5223 (N_5223,N_4569,N_4524);
nor U5224 (N_5224,N_4731,N_4577);
and U5225 (N_5225,N_4882,N_4574);
nand U5226 (N_5226,N_4786,N_4887);
nand U5227 (N_5227,N_4518,N_4640);
and U5228 (N_5228,N_4814,N_4587);
or U5229 (N_5229,N_4911,N_4948);
or U5230 (N_5230,N_4742,N_4712);
and U5231 (N_5231,N_4600,N_4638);
or U5232 (N_5232,N_4649,N_4525);
nor U5233 (N_5233,N_4568,N_4591);
nand U5234 (N_5234,N_4567,N_4508);
nor U5235 (N_5235,N_4964,N_4545);
nand U5236 (N_5236,N_4629,N_4515);
nor U5237 (N_5237,N_4589,N_4858);
and U5238 (N_5238,N_4665,N_4543);
nor U5239 (N_5239,N_4674,N_4995);
and U5240 (N_5240,N_4621,N_4735);
xor U5241 (N_5241,N_4558,N_4641);
or U5242 (N_5242,N_4798,N_4675);
and U5243 (N_5243,N_4905,N_4842);
xor U5244 (N_5244,N_4901,N_4987);
or U5245 (N_5245,N_4906,N_4637);
xor U5246 (N_5246,N_4981,N_4625);
and U5247 (N_5247,N_4968,N_4588);
nor U5248 (N_5248,N_4719,N_4506);
nor U5249 (N_5249,N_4955,N_4873);
or U5250 (N_5250,N_4663,N_4886);
and U5251 (N_5251,N_4940,N_4868);
and U5252 (N_5252,N_4861,N_4980);
and U5253 (N_5253,N_4593,N_4578);
or U5254 (N_5254,N_4751,N_4699);
xnor U5255 (N_5255,N_4553,N_4788);
nor U5256 (N_5256,N_4754,N_4596);
nor U5257 (N_5257,N_4585,N_4760);
nor U5258 (N_5258,N_4506,N_4739);
nor U5259 (N_5259,N_4891,N_4821);
nor U5260 (N_5260,N_4908,N_4859);
nor U5261 (N_5261,N_4568,N_4801);
nand U5262 (N_5262,N_4879,N_4992);
nor U5263 (N_5263,N_4599,N_4586);
nand U5264 (N_5264,N_4986,N_4763);
nor U5265 (N_5265,N_4934,N_4571);
nand U5266 (N_5266,N_4555,N_4560);
nand U5267 (N_5267,N_4720,N_4824);
nand U5268 (N_5268,N_4587,N_4847);
nor U5269 (N_5269,N_4613,N_4982);
and U5270 (N_5270,N_4759,N_4865);
nor U5271 (N_5271,N_4826,N_4664);
and U5272 (N_5272,N_4605,N_4859);
or U5273 (N_5273,N_4518,N_4862);
nand U5274 (N_5274,N_4569,N_4790);
or U5275 (N_5275,N_4866,N_4843);
nor U5276 (N_5276,N_4931,N_4890);
nand U5277 (N_5277,N_4950,N_4959);
and U5278 (N_5278,N_4885,N_4553);
and U5279 (N_5279,N_4904,N_4618);
nand U5280 (N_5280,N_4542,N_4698);
and U5281 (N_5281,N_4797,N_4697);
or U5282 (N_5282,N_4616,N_4956);
and U5283 (N_5283,N_4732,N_4887);
and U5284 (N_5284,N_4839,N_4613);
nand U5285 (N_5285,N_4659,N_4504);
nand U5286 (N_5286,N_4702,N_4876);
or U5287 (N_5287,N_4710,N_4962);
and U5288 (N_5288,N_4974,N_4622);
nand U5289 (N_5289,N_4737,N_4992);
nand U5290 (N_5290,N_4855,N_4835);
nor U5291 (N_5291,N_4651,N_4567);
and U5292 (N_5292,N_4688,N_4826);
nand U5293 (N_5293,N_4906,N_4691);
and U5294 (N_5294,N_4943,N_4903);
nor U5295 (N_5295,N_4998,N_4803);
or U5296 (N_5296,N_4991,N_4997);
nor U5297 (N_5297,N_4568,N_4579);
nor U5298 (N_5298,N_4790,N_4879);
xor U5299 (N_5299,N_4802,N_4572);
or U5300 (N_5300,N_4706,N_4942);
or U5301 (N_5301,N_4857,N_4926);
xor U5302 (N_5302,N_4636,N_4912);
xnor U5303 (N_5303,N_4638,N_4567);
and U5304 (N_5304,N_4970,N_4928);
nor U5305 (N_5305,N_4948,N_4829);
nand U5306 (N_5306,N_4544,N_4879);
nor U5307 (N_5307,N_4777,N_4601);
nand U5308 (N_5308,N_4844,N_4597);
and U5309 (N_5309,N_4890,N_4936);
and U5310 (N_5310,N_4590,N_4896);
or U5311 (N_5311,N_4872,N_4538);
or U5312 (N_5312,N_4541,N_4566);
xnor U5313 (N_5313,N_4893,N_4798);
nor U5314 (N_5314,N_4715,N_4838);
and U5315 (N_5315,N_4605,N_4980);
nor U5316 (N_5316,N_4812,N_4950);
and U5317 (N_5317,N_4577,N_4882);
nand U5318 (N_5318,N_4990,N_4813);
and U5319 (N_5319,N_4848,N_4671);
nor U5320 (N_5320,N_4792,N_4616);
nand U5321 (N_5321,N_4723,N_4589);
and U5322 (N_5322,N_4725,N_4549);
nor U5323 (N_5323,N_4958,N_4854);
nand U5324 (N_5324,N_4898,N_4715);
and U5325 (N_5325,N_4819,N_4825);
nor U5326 (N_5326,N_4619,N_4725);
or U5327 (N_5327,N_4759,N_4981);
nor U5328 (N_5328,N_4840,N_4587);
and U5329 (N_5329,N_4831,N_4818);
nand U5330 (N_5330,N_4641,N_4889);
or U5331 (N_5331,N_4574,N_4512);
xor U5332 (N_5332,N_4653,N_4887);
or U5333 (N_5333,N_4998,N_4605);
nor U5334 (N_5334,N_4934,N_4585);
nor U5335 (N_5335,N_4893,N_4906);
nand U5336 (N_5336,N_4831,N_4672);
and U5337 (N_5337,N_4949,N_4975);
and U5338 (N_5338,N_4632,N_4776);
nor U5339 (N_5339,N_4885,N_4512);
nand U5340 (N_5340,N_4938,N_4926);
nor U5341 (N_5341,N_4828,N_4961);
nand U5342 (N_5342,N_4516,N_4929);
nand U5343 (N_5343,N_4565,N_4651);
nor U5344 (N_5344,N_4827,N_4828);
nor U5345 (N_5345,N_4782,N_4817);
nor U5346 (N_5346,N_4803,N_4750);
nand U5347 (N_5347,N_4985,N_4687);
xor U5348 (N_5348,N_4698,N_4604);
xnor U5349 (N_5349,N_4951,N_4995);
or U5350 (N_5350,N_4821,N_4990);
or U5351 (N_5351,N_4703,N_4983);
or U5352 (N_5352,N_4638,N_4625);
or U5353 (N_5353,N_4882,N_4841);
xor U5354 (N_5354,N_4595,N_4548);
nand U5355 (N_5355,N_4582,N_4936);
nor U5356 (N_5356,N_4772,N_4999);
and U5357 (N_5357,N_4835,N_4922);
xnor U5358 (N_5358,N_4968,N_4691);
nand U5359 (N_5359,N_4587,N_4904);
or U5360 (N_5360,N_4832,N_4712);
nand U5361 (N_5361,N_4756,N_4916);
or U5362 (N_5362,N_4681,N_4883);
or U5363 (N_5363,N_4536,N_4864);
or U5364 (N_5364,N_4644,N_4609);
nor U5365 (N_5365,N_4524,N_4697);
nor U5366 (N_5366,N_4667,N_4678);
nor U5367 (N_5367,N_4682,N_4568);
or U5368 (N_5368,N_4634,N_4728);
nor U5369 (N_5369,N_4904,N_4911);
and U5370 (N_5370,N_4844,N_4987);
or U5371 (N_5371,N_4831,N_4898);
nor U5372 (N_5372,N_4810,N_4676);
xor U5373 (N_5373,N_4722,N_4898);
nor U5374 (N_5374,N_4964,N_4585);
nor U5375 (N_5375,N_4913,N_4959);
and U5376 (N_5376,N_4666,N_4965);
nor U5377 (N_5377,N_4780,N_4885);
nor U5378 (N_5378,N_4752,N_4759);
nand U5379 (N_5379,N_4618,N_4521);
nand U5380 (N_5380,N_4956,N_4524);
xnor U5381 (N_5381,N_4993,N_4554);
or U5382 (N_5382,N_4661,N_4865);
nand U5383 (N_5383,N_4941,N_4920);
nor U5384 (N_5384,N_4795,N_4766);
or U5385 (N_5385,N_4563,N_4871);
nand U5386 (N_5386,N_4683,N_4597);
nand U5387 (N_5387,N_4726,N_4676);
nand U5388 (N_5388,N_4942,N_4729);
or U5389 (N_5389,N_4981,N_4956);
and U5390 (N_5390,N_4706,N_4928);
nand U5391 (N_5391,N_4547,N_4828);
and U5392 (N_5392,N_4843,N_4554);
nor U5393 (N_5393,N_4948,N_4735);
or U5394 (N_5394,N_4583,N_4610);
and U5395 (N_5395,N_4525,N_4680);
nor U5396 (N_5396,N_4778,N_4656);
or U5397 (N_5397,N_4806,N_4612);
and U5398 (N_5398,N_4595,N_4643);
nor U5399 (N_5399,N_4591,N_4662);
nand U5400 (N_5400,N_4549,N_4872);
and U5401 (N_5401,N_4821,N_4895);
nor U5402 (N_5402,N_4838,N_4764);
nand U5403 (N_5403,N_4637,N_4730);
or U5404 (N_5404,N_4765,N_4954);
xnor U5405 (N_5405,N_4801,N_4679);
xor U5406 (N_5406,N_4759,N_4605);
or U5407 (N_5407,N_4651,N_4623);
and U5408 (N_5408,N_4625,N_4668);
nor U5409 (N_5409,N_4821,N_4943);
xor U5410 (N_5410,N_4814,N_4797);
nand U5411 (N_5411,N_4598,N_4859);
and U5412 (N_5412,N_4816,N_4587);
nand U5413 (N_5413,N_4699,N_4862);
nand U5414 (N_5414,N_4793,N_4955);
or U5415 (N_5415,N_4768,N_4521);
and U5416 (N_5416,N_4590,N_4549);
nor U5417 (N_5417,N_4769,N_4927);
and U5418 (N_5418,N_4602,N_4823);
nand U5419 (N_5419,N_4840,N_4872);
nand U5420 (N_5420,N_4765,N_4623);
and U5421 (N_5421,N_4997,N_4988);
nor U5422 (N_5422,N_4648,N_4546);
or U5423 (N_5423,N_4625,N_4752);
nand U5424 (N_5424,N_4927,N_4976);
and U5425 (N_5425,N_4537,N_4784);
and U5426 (N_5426,N_4895,N_4871);
and U5427 (N_5427,N_4610,N_4801);
xor U5428 (N_5428,N_4537,N_4836);
xnor U5429 (N_5429,N_4641,N_4917);
nor U5430 (N_5430,N_4759,N_4895);
nor U5431 (N_5431,N_4858,N_4982);
nor U5432 (N_5432,N_4994,N_4849);
nor U5433 (N_5433,N_4599,N_4706);
and U5434 (N_5434,N_4635,N_4787);
and U5435 (N_5435,N_4758,N_4524);
and U5436 (N_5436,N_4661,N_4545);
nor U5437 (N_5437,N_4686,N_4659);
or U5438 (N_5438,N_4906,N_4681);
and U5439 (N_5439,N_4593,N_4876);
xnor U5440 (N_5440,N_4534,N_4904);
and U5441 (N_5441,N_4506,N_4523);
nor U5442 (N_5442,N_4508,N_4536);
xnor U5443 (N_5443,N_4905,N_4785);
nor U5444 (N_5444,N_4778,N_4676);
nand U5445 (N_5445,N_4806,N_4774);
nand U5446 (N_5446,N_4576,N_4985);
and U5447 (N_5447,N_4904,N_4993);
or U5448 (N_5448,N_4575,N_4688);
nor U5449 (N_5449,N_4782,N_4994);
nand U5450 (N_5450,N_4850,N_4705);
and U5451 (N_5451,N_4609,N_4752);
and U5452 (N_5452,N_4710,N_4524);
and U5453 (N_5453,N_4838,N_4798);
and U5454 (N_5454,N_4556,N_4989);
nor U5455 (N_5455,N_4816,N_4604);
and U5456 (N_5456,N_4841,N_4614);
and U5457 (N_5457,N_4688,N_4879);
and U5458 (N_5458,N_4711,N_4733);
nand U5459 (N_5459,N_4791,N_4859);
xor U5460 (N_5460,N_4922,N_4712);
and U5461 (N_5461,N_4976,N_4744);
nand U5462 (N_5462,N_4826,N_4996);
nor U5463 (N_5463,N_4742,N_4769);
or U5464 (N_5464,N_4829,N_4981);
or U5465 (N_5465,N_4771,N_4733);
nor U5466 (N_5466,N_4751,N_4589);
nand U5467 (N_5467,N_4793,N_4842);
and U5468 (N_5468,N_4942,N_4945);
or U5469 (N_5469,N_4972,N_4503);
nand U5470 (N_5470,N_4570,N_4537);
and U5471 (N_5471,N_4755,N_4909);
nor U5472 (N_5472,N_4632,N_4899);
or U5473 (N_5473,N_4874,N_4530);
nand U5474 (N_5474,N_4681,N_4656);
and U5475 (N_5475,N_4876,N_4952);
or U5476 (N_5476,N_4859,N_4557);
or U5477 (N_5477,N_4948,N_4860);
or U5478 (N_5478,N_4542,N_4875);
and U5479 (N_5479,N_4772,N_4811);
or U5480 (N_5480,N_4555,N_4650);
nand U5481 (N_5481,N_4526,N_4747);
xor U5482 (N_5482,N_4592,N_4991);
or U5483 (N_5483,N_4717,N_4901);
and U5484 (N_5484,N_4614,N_4655);
or U5485 (N_5485,N_4879,N_4536);
nor U5486 (N_5486,N_4521,N_4849);
and U5487 (N_5487,N_4877,N_4977);
or U5488 (N_5488,N_4579,N_4930);
nand U5489 (N_5489,N_4758,N_4766);
nand U5490 (N_5490,N_4864,N_4672);
nor U5491 (N_5491,N_4555,N_4770);
nor U5492 (N_5492,N_4739,N_4623);
nand U5493 (N_5493,N_4528,N_4741);
nor U5494 (N_5494,N_4629,N_4842);
nand U5495 (N_5495,N_4795,N_4539);
and U5496 (N_5496,N_4661,N_4508);
nor U5497 (N_5497,N_4898,N_4632);
nor U5498 (N_5498,N_4719,N_4994);
or U5499 (N_5499,N_4881,N_4728);
nand U5500 (N_5500,N_5241,N_5310);
or U5501 (N_5501,N_5442,N_5372);
or U5502 (N_5502,N_5279,N_5253);
nand U5503 (N_5503,N_5060,N_5357);
and U5504 (N_5504,N_5295,N_5132);
nor U5505 (N_5505,N_5321,N_5291);
xor U5506 (N_5506,N_5314,N_5477);
and U5507 (N_5507,N_5107,N_5037);
nand U5508 (N_5508,N_5334,N_5306);
and U5509 (N_5509,N_5034,N_5152);
xnor U5510 (N_5510,N_5359,N_5026);
or U5511 (N_5511,N_5033,N_5457);
xor U5512 (N_5512,N_5389,N_5488);
and U5513 (N_5513,N_5215,N_5064);
nor U5514 (N_5514,N_5169,N_5089);
or U5515 (N_5515,N_5467,N_5013);
xor U5516 (N_5516,N_5230,N_5146);
xnor U5517 (N_5517,N_5087,N_5054);
nand U5518 (N_5518,N_5300,N_5323);
xor U5519 (N_5519,N_5260,N_5237);
or U5520 (N_5520,N_5309,N_5434);
or U5521 (N_5521,N_5124,N_5205);
nand U5522 (N_5522,N_5119,N_5340);
nand U5523 (N_5523,N_5395,N_5282);
or U5524 (N_5524,N_5298,N_5272);
or U5525 (N_5525,N_5421,N_5185);
nor U5526 (N_5526,N_5112,N_5284);
nand U5527 (N_5527,N_5437,N_5096);
nor U5528 (N_5528,N_5375,N_5329);
and U5529 (N_5529,N_5407,N_5496);
and U5530 (N_5530,N_5181,N_5019);
or U5531 (N_5531,N_5045,N_5180);
or U5532 (N_5532,N_5247,N_5251);
or U5533 (N_5533,N_5402,N_5447);
xnor U5534 (N_5534,N_5242,N_5108);
and U5535 (N_5535,N_5497,N_5191);
nor U5536 (N_5536,N_5330,N_5418);
or U5537 (N_5537,N_5262,N_5393);
or U5538 (N_5538,N_5443,N_5209);
nor U5539 (N_5539,N_5490,N_5367);
or U5540 (N_5540,N_5120,N_5204);
nor U5541 (N_5541,N_5238,N_5322);
and U5542 (N_5542,N_5212,N_5479);
and U5543 (N_5543,N_5102,N_5485);
or U5544 (N_5544,N_5154,N_5118);
nand U5545 (N_5545,N_5266,N_5370);
xnor U5546 (N_5546,N_5377,N_5223);
nand U5547 (N_5547,N_5125,N_5428);
or U5548 (N_5548,N_5290,N_5148);
nand U5549 (N_5549,N_5369,N_5133);
and U5550 (N_5550,N_5127,N_5448);
xor U5551 (N_5551,N_5051,N_5287);
or U5552 (N_5552,N_5470,N_5097);
or U5553 (N_5553,N_5258,N_5243);
nor U5554 (N_5554,N_5214,N_5384);
and U5555 (N_5555,N_5140,N_5186);
or U5556 (N_5556,N_5208,N_5173);
nand U5557 (N_5557,N_5403,N_5203);
nand U5558 (N_5558,N_5065,N_5093);
or U5559 (N_5559,N_5368,N_5017);
or U5560 (N_5560,N_5195,N_5349);
nor U5561 (N_5561,N_5201,N_5299);
nor U5562 (N_5562,N_5240,N_5339);
or U5563 (N_5563,N_5158,N_5128);
nand U5564 (N_5564,N_5226,N_5441);
nor U5565 (N_5565,N_5382,N_5016);
and U5566 (N_5566,N_5345,N_5025);
or U5567 (N_5567,N_5378,N_5010);
nand U5568 (N_5568,N_5246,N_5333);
nor U5569 (N_5569,N_5233,N_5491);
nand U5570 (N_5570,N_5030,N_5465);
nand U5571 (N_5571,N_5385,N_5390);
or U5572 (N_5572,N_5342,N_5341);
or U5573 (N_5573,N_5250,N_5101);
and U5574 (N_5574,N_5256,N_5104);
or U5575 (N_5575,N_5244,N_5141);
nor U5576 (N_5576,N_5474,N_5024);
and U5577 (N_5577,N_5446,N_5379);
xnor U5578 (N_5578,N_5406,N_5399);
and U5579 (N_5579,N_5110,N_5380);
or U5580 (N_5580,N_5396,N_5464);
xnor U5581 (N_5581,N_5143,N_5175);
and U5582 (N_5582,N_5044,N_5021);
and U5583 (N_5583,N_5301,N_5014);
or U5584 (N_5584,N_5398,N_5009);
or U5585 (N_5585,N_5066,N_5072);
and U5586 (N_5586,N_5011,N_5095);
nand U5587 (N_5587,N_5248,N_5049);
nor U5588 (N_5588,N_5002,N_5289);
nor U5589 (N_5589,N_5028,N_5040);
or U5590 (N_5590,N_5471,N_5164);
and U5591 (N_5591,N_5417,N_5466);
nor U5592 (N_5592,N_5454,N_5356);
nor U5593 (N_5593,N_5171,N_5035);
nand U5594 (N_5594,N_5062,N_5346);
and U5595 (N_5595,N_5492,N_5217);
and U5596 (N_5596,N_5187,N_5387);
nand U5597 (N_5597,N_5271,N_5365);
or U5598 (N_5598,N_5015,N_5255);
nand U5599 (N_5599,N_5422,N_5235);
nor U5600 (N_5600,N_5332,N_5351);
nand U5601 (N_5601,N_5313,N_5225);
and U5602 (N_5602,N_5361,N_5023);
nor U5603 (N_5603,N_5106,N_5157);
and U5604 (N_5604,N_5394,N_5316);
and U5605 (N_5605,N_5177,N_5168);
nand U5606 (N_5606,N_5145,N_5219);
or U5607 (N_5607,N_5400,N_5027);
or U5608 (N_5608,N_5139,N_5222);
or U5609 (N_5609,N_5151,N_5355);
nand U5610 (N_5610,N_5381,N_5412);
and U5611 (N_5611,N_5468,N_5193);
or U5612 (N_5612,N_5461,N_5288);
and U5613 (N_5613,N_5259,N_5331);
nand U5614 (N_5614,N_5416,N_5000);
nand U5615 (N_5615,N_5162,N_5179);
nand U5616 (N_5616,N_5278,N_5047);
and U5617 (N_5617,N_5264,N_5493);
and U5618 (N_5618,N_5482,N_5254);
and U5619 (N_5619,N_5196,N_5307);
and U5620 (N_5620,N_5304,N_5336);
and U5621 (N_5621,N_5131,N_5392);
and U5622 (N_5622,N_5293,N_5232);
or U5623 (N_5623,N_5487,N_5194);
nor U5624 (N_5624,N_5170,N_5094);
nand U5625 (N_5625,N_5189,N_5480);
and U5626 (N_5626,N_5086,N_5001);
nand U5627 (N_5627,N_5135,N_5043);
and U5628 (N_5628,N_5354,N_5070);
nand U5629 (N_5629,N_5147,N_5167);
xor U5630 (N_5630,N_5294,N_5455);
and U5631 (N_5631,N_5489,N_5325);
nand U5632 (N_5632,N_5165,N_5042);
nand U5633 (N_5633,N_5268,N_5360);
or U5634 (N_5634,N_5456,N_5430);
nand U5635 (N_5635,N_5012,N_5075);
or U5636 (N_5636,N_5353,N_5426);
and U5637 (N_5637,N_5032,N_5252);
and U5638 (N_5638,N_5486,N_5444);
xor U5639 (N_5639,N_5363,N_5404);
and U5640 (N_5640,N_5200,N_5098);
and U5641 (N_5641,N_5211,N_5029);
and U5642 (N_5642,N_5216,N_5386);
nand U5643 (N_5643,N_5499,N_5156);
nor U5644 (N_5644,N_5319,N_5198);
and U5645 (N_5645,N_5144,N_5129);
nand U5646 (N_5646,N_5311,N_5275);
nor U5647 (N_5647,N_5458,N_5391);
nand U5648 (N_5648,N_5111,N_5324);
nor U5649 (N_5649,N_5183,N_5472);
or U5650 (N_5650,N_5058,N_5085);
nor U5651 (N_5651,N_5130,N_5149);
nor U5652 (N_5652,N_5338,N_5061);
and U5653 (N_5653,N_5199,N_5192);
or U5654 (N_5654,N_5285,N_5335);
or U5655 (N_5655,N_5231,N_5302);
and U5656 (N_5656,N_5092,N_5435);
and U5657 (N_5657,N_5292,N_5452);
nor U5658 (N_5658,N_5178,N_5445);
xnor U5659 (N_5659,N_5303,N_5245);
or U5660 (N_5660,N_5413,N_5305);
or U5661 (N_5661,N_5427,N_5174);
nand U5662 (N_5662,N_5206,N_5105);
nand U5663 (N_5663,N_5376,N_5041);
nand U5664 (N_5664,N_5383,N_5077);
nand U5665 (N_5665,N_5419,N_5048);
xor U5666 (N_5666,N_5213,N_5257);
or U5667 (N_5667,N_5004,N_5069);
nand U5668 (N_5668,N_5224,N_5283);
nand U5669 (N_5669,N_5270,N_5317);
or U5670 (N_5670,N_5082,N_5273);
nand U5671 (N_5671,N_5475,N_5197);
or U5672 (N_5672,N_5003,N_5005);
nand U5673 (N_5673,N_5440,N_5436);
and U5674 (N_5674,N_5153,N_5155);
and U5675 (N_5675,N_5308,N_5078);
nand U5676 (N_5676,N_5473,N_5320);
or U5677 (N_5677,N_5074,N_5439);
nand U5678 (N_5678,N_5059,N_5134);
nor U5679 (N_5679,N_5388,N_5022);
or U5680 (N_5680,N_5274,N_5207);
and U5681 (N_5681,N_5055,N_5121);
nor U5682 (N_5682,N_5073,N_5081);
nor U5683 (N_5683,N_5415,N_5343);
nor U5684 (N_5684,N_5462,N_5210);
nor U5685 (N_5685,N_5063,N_5056);
and U5686 (N_5686,N_5460,N_5176);
nor U5687 (N_5687,N_5008,N_5036);
and U5688 (N_5688,N_5449,N_5163);
nor U5689 (N_5689,N_5498,N_5067);
nor U5690 (N_5690,N_5166,N_5397);
nand U5691 (N_5691,N_5018,N_5431);
nand U5692 (N_5692,N_5184,N_5344);
xor U5693 (N_5693,N_5429,N_5068);
nor U5694 (N_5694,N_5052,N_5451);
nor U5695 (N_5695,N_5433,N_5090);
and U5696 (N_5696,N_5337,N_5265);
nor U5697 (N_5697,N_5432,N_5296);
nor U5698 (N_5698,N_5076,N_5160);
nor U5699 (N_5699,N_5236,N_5006);
and U5700 (N_5700,N_5116,N_5053);
or U5701 (N_5701,N_5234,N_5495);
xor U5702 (N_5702,N_5352,N_5050);
nand U5703 (N_5703,N_5039,N_5202);
xor U5704 (N_5704,N_5286,N_5228);
xor U5705 (N_5705,N_5142,N_5318);
nand U5706 (N_5706,N_5371,N_5281);
nand U5707 (N_5707,N_5373,N_5161);
nor U5708 (N_5708,N_5150,N_5221);
nor U5709 (N_5709,N_5159,N_5229);
nand U5710 (N_5710,N_5410,N_5326);
and U5711 (N_5711,N_5348,N_5020);
nand U5712 (N_5712,N_5476,N_5478);
nand U5713 (N_5713,N_5280,N_5083);
xnor U5714 (N_5714,N_5172,N_5038);
nor U5715 (N_5715,N_5057,N_5423);
or U5716 (N_5716,N_5113,N_5408);
and U5717 (N_5717,N_5084,N_5347);
and U5718 (N_5718,N_5100,N_5115);
nand U5719 (N_5719,N_5420,N_5414);
nor U5720 (N_5720,N_5091,N_5364);
and U5721 (N_5721,N_5276,N_5424);
and U5722 (N_5722,N_5182,N_5103);
or U5723 (N_5723,N_5297,N_5220);
and U5724 (N_5724,N_5249,N_5401);
or U5725 (N_5725,N_5328,N_5138);
nor U5726 (N_5726,N_5350,N_5079);
nor U5727 (N_5727,N_5405,N_5483);
and U5728 (N_5728,N_5453,N_5315);
and U5729 (N_5729,N_5463,N_5267);
or U5730 (N_5730,N_5218,N_5031);
or U5731 (N_5731,N_5190,N_5494);
nor U5732 (N_5732,N_5362,N_5277);
nor U5733 (N_5733,N_5137,N_5007);
or U5734 (N_5734,N_5358,N_5450);
xnor U5735 (N_5735,N_5046,N_5469);
nand U5736 (N_5736,N_5122,N_5136);
nor U5737 (N_5737,N_5374,N_5109);
or U5738 (N_5738,N_5438,N_5088);
and U5739 (N_5739,N_5188,N_5099);
nor U5740 (N_5740,N_5269,N_5080);
xor U5741 (N_5741,N_5123,N_5114);
nand U5742 (N_5742,N_5239,N_5126);
and U5743 (N_5743,N_5117,N_5227);
or U5744 (N_5744,N_5425,N_5261);
nor U5745 (N_5745,N_5409,N_5481);
and U5746 (N_5746,N_5263,N_5071);
and U5747 (N_5747,N_5484,N_5411);
nand U5748 (N_5748,N_5312,N_5327);
nand U5749 (N_5749,N_5459,N_5366);
nor U5750 (N_5750,N_5327,N_5020);
nand U5751 (N_5751,N_5298,N_5225);
nand U5752 (N_5752,N_5074,N_5199);
xnor U5753 (N_5753,N_5407,N_5223);
and U5754 (N_5754,N_5250,N_5352);
nor U5755 (N_5755,N_5371,N_5445);
or U5756 (N_5756,N_5138,N_5011);
nor U5757 (N_5757,N_5321,N_5289);
nor U5758 (N_5758,N_5158,N_5011);
and U5759 (N_5759,N_5101,N_5188);
nor U5760 (N_5760,N_5128,N_5029);
nor U5761 (N_5761,N_5126,N_5300);
and U5762 (N_5762,N_5444,N_5313);
nor U5763 (N_5763,N_5264,N_5183);
nor U5764 (N_5764,N_5012,N_5148);
nand U5765 (N_5765,N_5484,N_5455);
nand U5766 (N_5766,N_5403,N_5414);
and U5767 (N_5767,N_5410,N_5113);
or U5768 (N_5768,N_5134,N_5267);
nand U5769 (N_5769,N_5290,N_5489);
xor U5770 (N_5770,N_5322,N_5248);
or U5771 (N_5771,N_5251,N_5166);
nor U5772 (N_5772,N_5296,N_5365);
nand U5773 (N_5773,N_5035,N_5353);
nor U5774 (N_5774,N_5463,N_5417);
or U5775 (N_5775,N_5270,N_5045);
and U5776 (N_5776,N_5040,N_5170);
nor U5777 (N_5777,N_5487,N_5002);
nand U5778 (N_5778,N_5344,N_5012);
and U5779 (N_5779,N_5433,N_5155);
or U5780 (N_5780,N_5201,N_5337);
nor U5781 (N_5781,N_5247,N_5348);
nand U5782 (N_5782,N_5021,N_5323);
nor U5783 (N_5783,N_5422,N_5040);
or U5784 (N_5784,N_5029,N_5325);
nand U5785 (N_5785,N_5186,N_5118);
nor U5786 (N_5786,N_5067,N_5397);
and U5787 (N_5787,N_5367,N_5115);
and U5788 (N_5788,N_5428,N_5185);
or U5789 (N_5789,N_5398,N_5150);
nand U5790 (N_5790,N_5435,N_5451);
or U5791 (N_5791,N_5151,N_5118);
and U5792 (N_5792,N_5477,N_5312);
or U5793 (N_5793,N_5455,N_5099);
xnor U5794 (N_5794,N_5073,N_5372);
nor U5795 (N_5795,N_5129,N_5259);
and U5796 (N_5796,N_5254,N_5159);
nor U5797 (N_5797,N_5046,N_5271);
and U5798 (N_5798,N_5259,N_5207);
and U5799 (N_5799,N_5343,N_5272);
or U5800 (N_5800,N_5128,N_5386);
xnor U5801 (N_5801,N_5249,N_5030);
or U5802 (N_5802,N_5485,N_5198);
or U5803 (N_5803,N_5495,N_5418);
or U5804 (N_5804,N_5488,N_5022);
and U5805 (N_5805,N_5456,N_5197);
and U5806 (N_5806,N_5358,N_5047);
nand U5807 (N_5807,N_5345,N_5200);
nand U5808 (N_5808,N_5123,N_5277);
and U5809 (N_5809,N_5477,N_5078);
nor U5810 (N_5810,N_5359,N_5142);
nor U5811 (N_5811,N_5426,N_5458);
nor U5812 (N_5812,N_5410,N_5330);
and U5813 (N_5813,N_5051,N_5024);
xor U5814 (N_5814,N_5091,N_5142);
nor U5815 (N_5815,N_5264,N_5195);
and U5816 (N_5816,N_5052,N_5036);
xnor U5817 (N_5817,N_5446,N_5178);
or U5818 (N_5818,N_5270,N_5121);
and U5819 (N_5819,N_5151,N_5063);
nor U5820 (N_5820,N_5378,N_5250);
nand U5821 (N_5821,N_5198,N_5074);
nor U5822 (N_5822,N_5318,N_5134);
nand U5823 (N_5823,N_5428,N_5069);
nor U5824 (N_5824,N_5006,N_5130);
xnor U5825 (N_5825,N_5266,N_5401);
nand U5826 (N_5826,N_5269,N_5474);
or U5827 (N_5827,N_5009,N_5274);
or U5828 (N_5828,N_5417,N_5209);
nor U5829 (N_5829,N_5173,N_5321);
nand U5830 (N_5830,N_5476,N_5318);
and U5831 (N_5831,N_5036,N_5134);
and U5832 (N_5832,N_5320,N_5401);
and U5833 (N_5833,N_5020,N_5292);
or U5834 (N_5834,N_5014,N_5326);
nand U5835 (N_5835,N_5155,N_5034);
and U5836 (N_5836,N_5363,N_5390);
nor U5837 (N_5837,N_5238,N_5331);
or U5838 (N_5838,N_5098,N_5003);
or U5839 (N_5839,N_5259,N_5394);
and U5840 (N_5840,N_5005,N_5093);
nand U5841 (N_5841,N_5086,N_5272);
nand U5842 (N_5842,N_5105,N_5099);
and U5843 (N_5843,N_5354,N_5379);
or U5844 (N_5844,N_5294,N_5171);
or U5845 (N_5845,N_5263,N_5005);
nand U5846 (N_5846,N_5103,N_5210);
nor U5847 (N_5847,N_5262,N_5482);
or U5848 (N_5848,N_5303,N_5413);
nand U5849 (N_5849,N_5482,N_5090);
nand U5850 (N_5850,N_5336,N_5400);
nor U5851 (N_5851,N_5170,N_5293);
nor U5852 (N_5852,N_5449,N_5273);
or U5853 (N_5853,N_5006,N_5215);
nand U5854 (N_5854,N_5362,N_5152);
and U5855 (N_5855,N_5459,N_5208);
nand U5856 (N_5856,N_5354,N_5034);
nand U5857 (N_5857,N_5138,N_5400);
or U5858 (N_5858,N_5353,N_5472);
and U5859 (N_5859,N_5265,N_5374);
and U5860 (N_5860,N_5140,N_5358);
or U5861 (N_5861,N_5267,N_5218);
or U5862 (N_5862,N_5093,N_5155);
nor U5863 (N_5863,N_5009,N_5227);
nand U5864 (N_5864,N_5154,N_5012);
nor U5865 (N_5865,N_5460,N_5007);
nand U5866 (N_5866,N_5473,N_5151);
nor U5867 (N_5867,N_5229,N_5315);
nand U5868 (N_5868,N_5416,N_5087);
nand U5869 (N_5869,N_5046,N_5171);
and U5870 (N_5870,N_5107,N_5186);
nor U5871 (N_5871,N_5019,N_5221);
nand U5872 (N_5872,N_5106,N_5308);
nand U5873 (N_5873,N_5013,N_5115);
or U5874 (N_5874,N_5068,N_5302);
or U5875 (N_5875,N_5168,N_5459);
nand U5876 (N_5876,N_5476,N_5425);
nand U5877 (N_5877,N_5081,N_5150);
nor U5878 (N_5878,N_5040,N_5118);
nor U5879 (N_5879,N_5008,N_5428);
nand U5880 (N_5880,N_5095,N_5487);
or U5881 (N_5881,N_5049,N_5325);
nand U5882 (N_5882,N_5052,N_5265);
and U5883 (N_5883,N_5335,N_5365);
nor U5884 (N_5884,N_5114,N_5190);
and U5885 (N_5885,N_5473,N_5378);
or U5886 (N_5886,N_5243,N_5192);
xor U5887 (N_5887,N_5315,N_5465);
and U5888 (N_5888,N_5113,N_5434);
and U5889 (N_5889,N_5126,N_5067);
nand U5890 (N_5890,N_5344,N_5103);
and U5891 (N_5891,N_5405,N_5044);
nor U5892 (N_5892,N_5305,N_5491);
and U5893 (N_5893,N_5282,N_5001);
or U5894 (N_5894,N_5065,N_5416);
nand U5895 (N_5895,N_5202,N_5326);
or U5896 (N_5896,N_5371,N_5025);
and U5897 (N_5897,N_5415,N_5486);
and U5898 (N_5898,N_5097,N_5132);
nand U5899 (N_5899,N_5120,N_5250);
or U5900 (N_5900,N_5112,N_5116);
or U5901 (N_5901,N_5124,N_5033);
or U5902 (N_5902,N_5190,N_5391);
and U5903 (N_5903,N_5038,N_5407);
and U5904 (N_5904,N_5447,N_5249);
nor U5905 (N_5905,N_5446,N_5319);
or U5906 (N_5906,N_5282,N_5466);
or U5907 (N_5907,N_5200,N_5210);
and U5908 (N_5908,N_5258,N_5310);
or U5909 (N_5909,N_5206,N_5194);
nor U5910 (N_5910,N_5222,N_5210);
and U5911 (N_5911,N_5339,N_5297);
and U5912 (N_5912,N_5001,N_5456);
or U5913 (N_5913,N_5312,N_5030);
nand U5914 (N_5914,N_5319,N_5071);
and U5915 (N_5915,N_5272,N_5419);
nor U5916 (N_5916,N_5407,N_5071);
nor U5917 (N_5917,N_5076,N_5345);
and U5918 (N_5918,N_5286,N_5103);
or U5919 (N_5919,N_5149,N_5336);
or U5920 (N_5920,N_5445,N_5272);
nor U5921 (N_5921,N_5306,N_5127);
or U5922 (N_5922,N_5153,N_5349);
or U5923 (N_5923,N_5360,N_5092);
nand U5924 (N_5924,N_5140,N_5446);
and U5925 (N_5925,N_5122,N_5073);
nor U5926 (N_5926,N_5216,N_5334);
and U5927 (N_5927,N_5253,N_5290);
and U5928 (N_5928,N_5269,N_5484);
or U5929 (N_5929,N_5252,N_5137);
or U5930 (N_5930,N_5366,N_5018);
nand U5931 (N_5931,N_5491,N_5122);
or U5932 (N_5932,N_5248,N_5124);
or U5933 (N_5933,N_5056,N_5002);
or U5934 (N_5934,N_5249,N_5198);
or U5935 (N_5935,N_5070,N_5422);
and U5936 (N_5936,N_5122,N_5046);
nor U5937 (N_5937,N_5182,N_5269);
nor U5938 (N_5938,N_5359,N_5136);
nor U5939 (N_5939,N_5449,N_5490);
and U5940 (N_5940,N_5058,N_5128);
and U5941 (N_5941,N_5465,N_5039);
or U5942 (N_5942,N_5304,N_5171);
and U5943 (N_5943,N_5066,N_5412);
nor U5944 (N_5944,N_5290,N_5386);
nand U5945 (N_5945,N_5227,N_5150);
nor U5946 (N_5946,N_5159,N_5495);
nor U5947 (N_5947,N_5219,N_5261);
nor U5948 (N_5948,N_5070,N_5135);
nor U5949 (N_5949,N_5032,N_5343);
and U5950 (N_5950,N_5205,N_5043);
nor U5951 (N_5951,N_5343,N_5191);
or U5952 (N_5952,N_5164,N_5329);
and U5953 (N_5953,N_5311,N_5415);
and U5954 (N_5954,N_5483,N_5008);
nor U5955 (N_5955,N_5257,N_5072);
or U5956 (N_5956,N_5236,N_5072);
and U5957 (N_5957,N_5300,N_5008);
or U5958 (N_5958,N_5009,N_5100);
or U5959 (N_5959,N_5127,N_5212);
and U5960 (N_5960,N_5284,N_5121);
nor U5961 (N_5961,N_5481,N_5297);
nor U5962 (N_5962,N_5172,N_5424);
nor U5963 (N_5963,N_5007,N_5104);
and U5964 (N_5964,N_5196,N_5305);
and U5965 (N_5965,N_5131,N_5437);
xor U5966 (N_5966,N_5396,N_5380);
nand U5967 (N_5967,N_5419,N_5122);
nor U5968 (N_5968,N_5258,N_5459);
or U5969 (N_5969,N_5029,N_5262);
and U5970 (N_5970,N_5341,N_5495);
or U5971 (N_5971,N_5375,N_5372);
nand U5972 (N_5972,N_5282,N_5051);
nor U5973 (N_5973,N_5193,N_5195);
xor U5974 (N_5974,N_5298,N_5200);
or U5975 (N_5975,N_5104,N_5267);
and U5976 (N_5976,N_5354,N_5142);
or U5977 (N_5977,N_5245,N_5456);
nor U5978 (N_5978,N_5275,N_5239);
and U5979 (N_5979,N_5153,N_5251);
xor U5980 (N_5980,N_5448,N_5352);
and U5981 (N_5981,N_5355,N_5029);
and U5982 (N_5982,N_5012,N_5364);
nor U5983 (N_5983,N_5464,N_5483);
nand U5984 (N_5984,N_5238,N_5321);
nor U5985 (N_5985,N_5485,N_5271);
nand U5986 (N_5986,N_5475,N_5495);
or U5987 (N_5987,N_5371,N_5280);
nand U5988 (N_5988,N_5330,N_5411);
nand U5989 (N_5989,N_5385,N_5002);
and U5990 (N_5990,N_5199,N_5200);
nand U5991 (N_5991,N_5270,N_5063);
nand U5992 (N_5992,N_5369,N_5290);
nand U5993 (N_5993,N_5144,N_5289);
nor U5994 (N_5994,N_5352,N_5330);
nand U5995 (N_5995,N_5368,N_5097);
nor U5996 (N_5996,N_5021,N_5453);
xnor U5997 (N_5997,N_5266,N_5197);
nor U5998 (N_5998,N_5176,N_5224);
or U5999 (N_5999,N_5244,N_5229);
nand U6000 (N_6000,N_5668,N_5781);
and U6001 (N_6001,N_5586,N_5665);
or U6002 (N_6002,N_5900,N_5696);
nand U6003 (N_6003,N_5992,N_5980);
or U6004 (N_6004,N_5695,N_5858);
or U6005 (N_6005,N_5517,N_5930);
nand U6006 (N_6006,N_5567,N_5757);
or U6007 (N_6007,N_5521,N_5803);
xor U6008 (N_6008,N_5566,N_5963);
or U6009 (N_6009,N_5588,N_5537);
nor U6010 (N_6010,N_5699,N_5573);
xnor U6011 (N_6011,N_5706,N_5598);
nand U6012 (N_6012,N_5731,N_5880);
and U6013 (N_6013,N_5556,N_5984);
and U6014 (N_6014,N_5830,N_5794);
or U6015 (N_6015,N_5511,N_5810);
xor U6016 (N_6016,N_5946,N_5990);
and U6017 (N_6017,N_5952,N_5860);
nand U6018 (N_6018,N_5742,N_5605);
or U6019 (N_6019,N_5600,N_5898);
and U6020 (N_6020,N_5798,N_5863);
nand U6021 (N_6021,N_5532,N_5674);
nand U6022 (N_6022,N_5693,N_5680);
nor U6023 (N_6023,N_5604,N_5545);
nor U6024 (N_6024,N_5646,N_5761);
and U6025 (N_6025,N_5866,N_5628);
nand U6026 (N_6026,N_5637,N_5786);
xor U6027 (N_6027,N_5846,N_5844);
and U6028 (N_6028,N_5770,N_5893);
nor U6029 (N_6029,N_5635,N_5937);
nor U6030 (N_6030,N_5897,N_5750);
or U6031 (N_6031,N_5716,N_5998);
nand U6032 (N_6032,N_5621,N_5669);
nor U6033 (N_6033,N_5659,N_5953);
nor U6034 (N_6034,N_5778,N_5562);
nor U6035 (N_6035,N_5851,N_5585);
nor U6036 (N_6036,N_5554,N_5845);
or U6037 (N_6037,N_5656,N_5548);
xnor U6038 (N_6038,N_5741,N_5951);
nand U6039 (N_6039,N_5899,N_5597);
nand U6040 (N_6040,N_5964,N_5739);
nor U6041 (N_6041,N_5975,N_5772);
nand U6042 (N_6042,N_5785,N_5613);
nor U6043 (N_6043,N_5576,N_5634);
nand U6044 (N_6044,N_5994,N_5722);
nand U6045 (N_6045,N_5779,N_5692);
or U6046 (N_6046,N_5914,N_5957);
xnor U6047 (N_6047,N_5678,N_5821);
or U6048 (N_6048,N_5676,N_5728);
xor U6049 (N_6049,N_5662,N_5631);
nor U6050 (N_6050,N_5505,N_5666);
or U6051 (N_6051,N_5729,N_5753);
nand U6052 (N_6052,N_5891,N_5515);
nand U6053 (N_6053,N_5816,N_5721);
nand U6054 (N_6054,N_5825,N_5939);
and U6055 (N_6055,N_5620,N_5885);
or U6056 (N_6056,N_5758,N_5775);
xor U6057 (N_6057,N_5506,N_5861);
and U6058 (N_6058,N_5997,N_5657);
nand U6059 (N_6059,N_5911,N_5870);
or U6060 (N_6060,N_5852,N_5989);
and U6061 (N_6061,N_5912,N_5670);
or U6062 (N_6062,N_5767,N_5544);
nor U6063 (N_6063,N_5949,N_5811);
nand U6064 (N_6064,N_5967,N_5864);
nand U6065 (N_6065,N_5853,N_5787);
nor U6066 (N_6066,N_5649,N_5738);
nor U6067 (N_6067,N_5687,N_5812);
or U6068 (N_6068,N_5788,N_5549);
xnor U6069 (N_6069,N_5874,N_5538);
and U6070 (N_6070,N_5973,N_5632);
nor U6071 (N_6071,N_5726,N_5809);
nor U6072 (N_6072,N_5834,N_5942);
xor U6073 (N_6073,N_5815,N_5961);
nand U6074 (N_6074,N_5847,N_5901);
nor U6075 (N_6075,N_5652,N_5743);
nor U6076 (N_6076,N_5807,N_5614);
nand U6077 (N_6077,N_5882,N_5591);
xnor U6078 (N_6078,N_5854,N_5945);
and U6079 (N_6079,N_5983,N_5790);
nor U6080 (N_6080,N_5596,N_5641);
and U6081 (N_6081,N_5760,N_5651);
or U6082 (N_6082,N_5627,N_5580);
nand U6083 (N_6083,N_5615,N_5745);
nor U6084 (N_6084,N_5827,N_5644);
xor U6085 (N_6085,N_5601,N_5910);
nor U6086 (N_6086,N_5535,N_5671);
or U6087 (N_6087,N_5685,N_5660);
xor U6088 (N_6088,N_5648,N_5925);
xnor U6089 (N_6089,N_5971,N_5865);
nor U6090 (N_6090,N_5752,N_5623);
nand U6091 (N_6091,N_5813,N_5740);
and U6092 (N_6092,N_5697,N_5876);
or U6093 (N_6093,N_5565,N_5599);
nand U6094 (N_6094,N_5932,N_5579);
nand U6095 (N_6095,N_5985,N_5513);
and U6096 (N_6096,N_5675,N_5850);
or U6097 (N_6097,N_5658,N_5630);
and U6098 (N_6098,N_5751,N_5855);
nand U6099 (N_6099,N_5915,N_5818);
nand U6100 (N_6100,N_5645,N_5808);
or U6101 (N_6101,N_5875,N_5747);
xor U6102 (N_6102,N_5727,N_5711);
and U6103 (N_6103,N_5542,N_5619);
xnor U6104 (N_6104,N_5791,N_5749);
xnor U6105 (N_6105,N_5759,N_5793);
nor U6106 (N_6106,N_5768,N_5782);
nand U6107 (N_6107,N_5608,N_5958);
nand U6108 (N_6108,N_5895,N_5638);
nand U6109 (N_6109,N_5524,N_5650);
or U6110 (N_6110,N_5832,N_5969);
nand U6111 (N_6111,N_5633,N_5737);
or U6112 (N_6112,N_5709,N_5927);
and U6113 (N_6113,N_5718,N_5806);
or U6114 (N_6114,N_5654,N_5667);
or U6115 (N_6115,N_5530,N_5681);
nor U6116 (N_6116,N_5837,N_5878);
and U6117 (N_6117,N_5541,N_5869);
nor U6118 (N_6118,N_5777,N_5710);
or U6119 (N_6119,N_5966,N_5754);
nor U6120 (N_6120,N_5826,N_5841);
nand U6121 (N_6121,N_5636,N_5717);
and U6122 (N_6122,N_5501,N_5991);
or U6123 (N_6123,N_5823,N_5733);
xor U6124 (N_6124,N_5972,N_5609);
nor U6125 (N_6125,N_5887,N_5904);
and U6126 (N_6126,N_5574,N_5877);
nand U6127 (N_6127,N_5746,N_5606);
or U6128 (N_6128,N_5856,N_5756);
nor U6129 (N_6129,N_5928,N_5592);
nor U6130 (N_6130,N_5995,N_5610);
nand U6131 (N_6131,N_5618,N_5663);
or U6132 (N_6132,N_5974,N_5833);
nor U6133 (N_6133,N_5965,N_5577);
and U6134 (N_6134,N_5655,N_5944);
xnor U6135 (N_6135,N_5529,N_5929);
or U6136 (N_6136,N_5926,N_5546);
or U6137 (N_6137,N_5907,N_5642);
xnor U6138 (N_6138,N_5525,N_5744);
nand U6139 (N_6139,N_5800,N_5617);
nor U6140 (N_6140,N_5797,N_5734);
or U6141 (N_6141,N_5611,N_5873);
nor U6142 (N_6142,N_5802,N_5587);
xnor U6143 (N_6143,N_5672,N_5996);
nand U6144 (N_6144,N_5917,N_5702);
or U6145 (N_6145,N_5510,N_5715);
and U6146 (N_6146,N_5979,N_5552);
nand U6147 (N_6147,N_5842,N_5520);
or U6148 (N_6148,N_5884,N_5664);
or U6149 (N_6149,N_5694,N_5769);
nor U6150 (N_6150,N_5616,N_5819);
or U6151 (N_6151,N_5814,N_5590);
or U6152 (N_6152,N_5661,N_5922);
and U6153 (N_6153,N_5624,N_5647);
and U6154 (N_6154,N_5943,N_5843);
and U6155 (N_6155,N_5560,N_5575);
or U6156 (N_6156,N_5571,N_5730);
or U6157 (N_6157,N_5673,N_5539);
or U6158 (N_6158,N_5982,N_5999);
or U6159 (N_6159,N_5986,N_5547);
xor U6160 (N_6160,N_5602,N_5784);
nand U6161 (N_6161,N_5595,N_5504);
and U6162 (N_6162,N_5801,N_5507);
xnor U6163 (N_6163,N_5792,N_5516);
or U6164 (N_6164,N_5783,N_5955);
or U6165 (N_6165,N_5909,N_5931);
nand U6166 (N_6166,N_5522,N_5714);
or U6167 (N_6167,N_5581,N_5890);
and U6168 (N_6168,N_5677,N_5555);
nand U6169 (N_6169,N_5723,N_5805);
and U6170 (N_6170,N_5500,N_5684);
nor U6171 (N_6171,N_5748,N_5771);
or U6172 (N_6172,N_5840,N_5849);
nand U6173 (N_6173,N_5857,N_5872);
and U6174 (N_6174,N_5780,N_5795);
nor U6175 (N_6175,N_5977,N_5551);
xor U6176 (N_6176,N_5503,N_5941);
and U6177 (N_6177,N_5954,N_5643);
nand U6178 (N_6178,N_5838,N_5691);
or U6179 (N_6179,N_5701,N_5871);
and U6180 (N_6180,N_5527,N_5935);
xor U6181 (N_6181,N_5557,N_5987);
or U6182 (N_6182,N_5940,N_5594);
nand U6183 (N_6183,N_5707,N_5683);
or U6184 (N_6184,N_5584,N_5799);
nor U6185 (N_6185,N_5509,N_5950);
nor U6186 (N_6186,N_5564,N_5550);
nor U6187 (N_6187,N_5968,N_5703);
nor U6188 (N_6188,N_5578,N_5724);
nor U6189 (N_6189,N_5607,N_5916);
nand U6190 (N_6190,N_5888,N_5867);
xnor U6191 (N_6191,N_5906,N_5626);
nand U6192 (N_6192,N_5698,N_5713);
or U6193 (N_6193,N_5732,N_5923);
nand U6194 (N_6194,N_5705,N_5918);
xor U6195 (N_6195,N_5903,N_5755);
or U6196 (N_6196,N_5688,N_5981);
and U6197 (N_6197,N_5881,N_5708);
nand U6198 (N_6198,N_5921,N_5892);
and U6199 (N_6199,N_5774,N_5919);
or U6200 (N_6200,N_5603,N_5518);
xor U6201 (N_6201,N_5978,N_5736);
nand U6202 (N_6202,N_5540,N_5536);
nor U6203 (N_6203,N_5700,N_5976);
nor U6204 (N_6204,N_5924,N_5593);
and U6205 (N_6205,N_5913,N_5886);
and U6206 (N_6206,N_5612,N_5934);
or U6207 (N_6207,N_5835,N_5804);
nor U6208 (N_6208,N_5765,N_5558);
nand U6209 (N_6209,N_5773,N_5764);
and U6210 (N_6210,N_5948,N_5582);
nand U6211 (N_6211,N_5679,N_5938);
nand U6212 (N_6212,N_5817,N_5894);
nand U6213 (N_6213,N_5712,N_5762);
and U6214 (N_6214,N_5920,N_5640);
nor U6215 (N_6215,N_5993,N_5868);
and U6216 (N_6216,N_5639,N_5763);
nor U6217 (N_6217,N_5533,N_5570);
and U6218 (N_6218,N_5514,N_5563);
nor U6219 (N_6219,N_5796,N_5502);
xnor U6220 (N_6220,N_5589,N_5905);
or U6221 (N_6221,N_5789,N_5686);
nand U6222 (N_6222,N_5947,N_5959);
and U6223 (N_6223,N_5725,N_5508);
nand U6224 (N_6224,N_5690,N_5653);
or U6225 (N_6225,N_5528,N_5902);
or U6226 (N_6226,N_5682,N_5828);
and U6227 (N_6227,N_5862,N_5512);
nand U6228 (N_6228,N_5879,N_5526);
and U6229 (N_6229,N_5629,N_5908);
or U6230 (N_6230,N_5704,N_5572);
nor U6231 (N_6231,N_5776,N_5822);
nor U6232 (N_6232,N_5896,N_5583);
and U6233 (N_6233,N_5531,N_5622);
xnor U6234 (N_6234,N_5824,N_5689);
nor U6235 (N_6235,N_5720,N_5534);
and U6236 (N_6236,N_5519,N_5543);
or U6237 (N_6237,N_5956,N_5960);
nand U6238 (N_6238,N_5962,N_5848);
nand U6239 (N_6239,N_5936,N_5839);
nand U6240 (N_6240,N_5553,N_5568);
nand U6241 (N_6241,N_5829,N_5569);
nor U6242 (N_6242,N_5559,N_5988);
nor U6243 (N_6243,N_5970,N_5831);
xnor U6244 (N_6244,N_5719,N_5859);
nor U6245 (N_6245,N_5625,N_5883);
and U6246 (N_6246,N_5836,N_5889);
nand U6247 (N_6247,N_5820,N_5933);
xnor U6248 (N_6248,N_5766,N_5735);
nand U6249 (N_6249,N_5561,N_5523);
nor U6250 (N_6250,N_5750,N_5808);
nor U6251 (N_6251,N_5601,N_5923);
nand U6252 (N_6252,N_5852,N_5987);
and U6253 (N_6253,N_5510,N_5907);
or U6254 (N_6254,N_5530,N_5701);
nand U6255 (N_6255,N_5840,N_5903);
or U6256 (N_6256,N_5513,N_5959);
and U6257 (N_6257,N_5628,N_5586);
nand U6258 (N_6258,N_5795,N_5983);
and U6259 (N_6259,N_5600,N_5773);
nand U6260 (N_6260,N_5548,N_5752);
and U6261 (N_6261,N_5817,N_5992);
or U6262 (N_6262,N_5578,N_5849);
and U6263 (N_6263,N_5589,N_5706);
nand U6264 (N_6264,N_5898,N_5526);
or U6265 (N_6265,N_5636,N_5821);
and U6266 (N_6266,N_5620,N_5683);
xnor U6267 (N_6267,N_5989,N_5894);
nor U6268 (N_6268,N_5866,N_5602);
and U6269 (N_6269,N_5614,N_5849);
and U6270 (N_6270,N_5580,N_5959);
or U6271 (N_6271,N_5985,N_5625);
nor U6272 (N_6272,N_5845,N_5868);
xnor U6273 (N_6273,N_5793,N_5621);
or U6274 (N_6274,N_5558,N_5549);
xnor U6275 (N_6275,N_5837,N_5746);
and U6276 (N_6276,N_5828,N_5658);
or U6277 (N_6277,N_5704,N_5941);
and U6278 (N_6278,N_5626,N_5694);
nand U6279 (N_6279,N_5682,N_5970);
nor U6280 (N_6280,N_5690,N_5718);
xnor U6281 (N_6281,N_5799,N_5578);
nor U6282 (N_6282,N_5882,N_5727);
nand U6283 (N_6283,N_5656,N_5700);
and U6284 (N_6284,N_5779,N_5618);
or U6285 (N_6285,N_5583,N_5581);
and U6286 (N_6286,N_5551,N_5813);
xor U6287 (N_6287,N_5522,N_5631);
and U6288 (N_6288,N_5778,N_5815);
nand U6289 (N_6289,N_5749,N_5520);
xnor U6290 (N_6290,N_5808,N_5685);
nor U6291 (N_6291,N_5648,N_5581);
xnor U6292 (N_6292,N_5630,N_5786);
and U6293 (N_6293,N_5955,N_5694);
or U6294 (N_6294,N_5820,N_5740);
nand U6295 (N_6295,N_5654,N_5643);
xnor U6296 (N_6296,N_5957,N_5636);
xnor U6297 (N_6297,N_5505,N_5945);
and U6298 (N_6298,N_5701,N_5736);
nand U6299 (N_6299,N_5879,N_5820);
or U6300 (N_6300,N_5680,N_5822);
or U6301 (N_6301,N_5518,N_5912);
nor U6302 (N_6302,N_5923,N_5825);
or U6303 (N_6303,N_5592,N_5536);
nor U6304 (N_6304,N_5753,N_5868);
or U6305 (N_6305,N_5862,N_5875);
xor U6306 (N_6306,N_5559,N_5813);
xnor U6307 (N_6307,N_5784,N_5808);
nor U6308 (N_6308,N_5879,N_5833);
and U6309 (N_6309,N_5567,N_5874);
or U6310 (N_6310,N_5566,N_5567);
nor U6311 (N_6311,N_5909,N_5590);
or U6312 (N_6312,N_5633,N_5705);
xor U6313 (N_6313,N_5593,N_5868);
and U6314 (N_6314,N_5813,N_5527);
or U6315 (N_6315,N_5694,N_5964);
nor U6316 (N_6316,N_5673,N_5750);
or U6317 (N_6317,N_5948,N_5583);
xor U6318 (N_6318,N_5689,N_5712);
nand U6319 (N_6319,N_5972,N_5748);
and U6320 (N_6320,N_5619,N_5505);
or U6321 (N_6321,N_5727,N_5700);
xor U6322 (N_6322,N_5842,N_5951);
xor U6323 (N_6323,N_5805,N_5692);
and U6324 (N_6324,N_5682,N_5576);
xnor U6325 (N_6325,N_5943,N_5649);
nor U6326 (N_6326,N_5613,N_5621);
nand U6327 (N_6327,N_5733,N_5711);
or U6328 (N_6328,N_5570,N_5557);
and U6329 (N_6329,N_5964,N_5994);
xnor U6330 (N_6330,N_5681,N_5602);
and U6331 (N_6331,N_5900,N_5952);
and U6332 (N_6332,N_5581,N_5704);
or U6333 (N_6333,N_5879,N_5800);
nand U6334 (N_6334,N_5660,N_5898);
or U6335 (N_6335,N_5658,N_5536);
and U6336 (N_6336,N_5833,N_5661);
and U6337 (N_6337,N_5676,N_5556);
or U6338 (N_6338,N_5707,N_5825);
or U6339 (N_6339,N_5516,N_5971);
nor U6340 (N_6340,N_5683,N_5873);
nor U6341 (N_6341,N_5914,N_5524);
or U6342 (N_6342,N_5711,N_5776);
or U6343 (N_6343,N_5799,N_5546);
nor U6344 (N_6344,N_5532,N_5576);
and U6345 (N_6345,N_5727,N_5742);
nand U6346 (N_6346,N_5564,N_5972);
or U6347 (N_6347,N_5681,N_5850);
or U6348 (N_6348,N_5920,N_5746);
nand U6349 (N_6349,N_5717,N_5840);
xnor U6350 (N_6350,N_5547,N_5824);
nand U6351 (N_6351,N_5789,N_5897);
and U6352 (N_6352,N_5975,N_5831);
and U6353 (N_6353,N_5812,N_5755);
nand U6354 (N_6354,N_5550,N_5863);
or U6355 (N_6355,N_5681,N_5770);
or U6356 (N_6356,N_5524,N_5733);
nand U6357 (N_6357,N_5743,N_5842);
xnor U6358 (N_6358,N_5734,N_5807);
or U6359 (N_6359,N_5798,N_5956);
or U6360 (N_6360,N_5818,N_5806);
nand U6361 (N_6361,N_5564,N_5528);
xor U6362 (N_6362,N_5959,N_5830);
or U6363 (N_6363,N_5638,N_5949);
xnor U6364 (N_6364,N_5802,N_5761);
nand U6365 (N_6365,N_5523,N_5526);
or U6366 (N_6366,N_5827,N_5509);
nor U6367 (N_6367,N_5991,N_5515);
and U6368 (N_6368,N_5591,N_5708);
nand U6369 (N_6369,N_5505,N_5667);
xnor U6370 (N_6370,N_5798,N_5563);
and U6371 (N_6371,N_5637,N_5920);
nand U6372 (N_6372,N_5704,N_5641);
or U6373 (N_6373,N_5714,N_5603);
nor U6374 (N_6374,N_5674,N_5725);
or U6375 (N_6375,N_5961,N_5643);
nand U6376 (N_6376,N_5898,N_5668);
and U6377 (N_6377,N_5865,N_5585);
and U6378 (N_6378,N_5657,N_5870);
and U6379 (N_6379,N_5602,N_5837);
or U6380 (N_6380,N_5989,N_5982);
nor U6381 (N_6381,N_5710,N_5615);
nand U6382 (N_6382,N_5803,N_5597);
nand U6383 (N_6383,N_5937,N_5718);
or U6384 (N_6384,N_5896,N_5674);
or U6385 (N_6385,N_5627,N_5971);
xor U6386 (N_6386,N_5948,N_5594);
or U6387 (N_6387,N_5786,N_5937);
xor U6388 (N_6388,N_5557,N_5920);
nor U6389 (N_6389,N_5580,N_5736);
and U6390 (N_6390,N_5549,N_5825);
and U6391 (N_6391,N_5783,N_5868);
nand U6392 (N_6392,N_5595,N_5847);
nor U6393 (N_6393,N_5851,N_5533);
nor U6394 (N_6394,N_5738,N_5697);
nand U6395 (N_6395,N_5711,N_5628);
or U6396 (N_6396,N_5728,N_5952);
nand U6397 (N_6397,N_5909,N_5902);
xor U6398 (N_6398,N_5506,N_5865);
xor U6399 (N_6399,N_5547,N_5766);
nor U6400 (N_6400,N_5613,N_5807);
or U6401 (N_6401,N_5892,N_5667);
nand U6402 (N_6402,N_5733,N_5594);
or U6403 (N_6403,N_5502,N_5609);
nand U6404 (N_6404,N_5638,N_5793);
and U6405 (N_6405,N_5923,N_5983);
nor U6406 (N_6406,N_5723,N_5545);
nand U6407 (N_6407,N_5647,N_5552);
nand U6408 (N_6408,N_5880,N_5573);
nor U6409 (N_6409,N_5518,N_5827);
nand U6410 (N_6410,N_5735,N_5647);
or U6411 (N_6411,N_5593,N_5958);
or U6412 (N_6412,N_5942,N_5704);
nor U6413 (N_6413,N_5567,N_5630);
nor U6414 (N_6414,N_5725,N_5595);
nand U6415 (N_6415,N_5775,N_5517);
and U6416 (N_6416,N_5720,N_5744);
or U6417 (N_6417,N_5607,N_5748);
and U6418 (N_6418,N_5851,N_5951);
xnor U6419 (N_6419,N_5627,N_5818);
nand U6420 (N_6420,N_5981,N_5648);
nor U6421 (N_6421,N_5507,N_5855);
and U6422 (N_6422,N_5572,N_5679);
nor U6423 (N_6423,N_5660,N_5808);
or U6424 (N_6424,N_5605,N_5556);
xnor U6425 (N_6425,N_5797,N_5967);
nand U6426 (N_6426,N_5736,N_5713);
and U6427 (N_6427,N_5940,N_5702);
nand U6428 (N_6428,N_5935,N_5570);
or U6429 (N_6429,N_5600,N_5630);
xor U6430 (N_6430,N_5873,N_5561);
nor U6431 (N_6431,N_5918,N_5627);
or U6432 (N_6432,N_5690,N_5956);
nor U6433 (N_6433,N_5742,N_5713);
nor U6434 (N_6434,N_5758,N_5590);
nand U6435 (N_6435,N_5768,N_5861);
nor U6436 (N_6436,N_5537,N_5721);
nand U6437 (N_6437,N_5779,N_5811);
and U6438 (N_6438,N_5937,N_5989);
and U6439 (N_6439,N_5733,N_5559);
and U6440 (N_6440,N_5921,N_5821);
nand U6441 (N_6441,N_5935,N_5955);
or U6442 (N_6442,N_5913,N_5656);
or U6443 (N_6443,N_5693,N_5964);
nand U6444 (N_6444,N_5520,N_5745);
xnor U6445 (N_6445,N_5642,N_5761);
or U6446 (N_6446,N_5791,N_5658);
and U6447 (N_6447,N_5812,N_5789);
or U6448 (N_6448,N_5849,N_5655);
nor U6449 (N_6449,N_5778,N_5806);
nor U6450 (N_6450,N_5839,N_5626);
and U6451 (N_6451,N_5673,N_5800);
nand U6452 (N_6452,N_5715,N_5626);
xor U6453 (N_6453,N_5571,N_5754);
and U6454 (N_6454,N_5725,N_5623);
nor U6455 (N_6455,N_5721,N_5510);
nand U6456 (N_6456,N_5777,N_5994);
nor U6457 (N_6457,N_5665,N_5890);
or U6458 (N_6458,N_5519,N_5617);
and U6459 (N_6459,N_5555,N_5842);
and U6460 (N_6460,N_5707,N_5848);
nand U6461 (N_6461,N_5802,N_5502);
nor U6462 (N_6462,N_5586,N_5940);
nor U6463 (N_6463,N_5964,N_5779);
nand U6464 (N_6464,N_5803,N_5838);
nor U6465 (N_6465,N_5728,N_5855);
nand U6466 (N_6466,N_5734,N_5593);
nor U6467 (N_6467,N_5576,N_5522);
or U6468 (N_6468,N_5591,N_5843);
and U6469 (N_6469,N_5508,N_5794);
and U6470 (N_6470,N_5680,N_5607);
nor U6471 (N_6471,N_5997,N_5828);
nor U6472 (N_6472,N_5642,N_5729);
or U6473 (N_6473,N_5657,N_5635);
and U6474 (N_6474,N_5960,N_5515);
nand U6475 (N_6475,N_5851,N_5701);
nor U6476 (N_6476,N_5743,N_5828);
nand U6477 (N_6477,N_5898,N_5611);
or U6478 (N_6478,N_5994,N_5779);
or U6479 (N_6479,N_5800,N_5884);
and U6480 (N_6480,N_5750,N_5517);
nor U6481 (N_6481,N_5729,N_5885);
nand U6482 (N_6482,N_5617,N_5828);
xor U6483 (N_6483,N_5677,N_5646);
nor U6484 (N_6484,N_5821,N_5518);
or U6485 (N_6485,N_5768,N_5544);
nor U6486 (N_6486,N_5722,N_5599);
nand U6487 (N_6487,N_5679,N_5881);
or U6488 (N_6488,N_5630,N_5661);
nor U6489 (N_6489,N_5612,N_5710);
and U6490 (N_6490,N_5764,N_5518);
nor U6491 (N_6491,N_5849,N_5782);
nor U6492 (N_6492,N_5556,N_5567);
nand U6493 (N_6493,N_5870,N_5643);
nor U6494 (N_6494,N_5939,N_5624);
nand U6495 (N_6495,N_5657,N_5791);
nor U6496 (N_6496,N_5746,N_5614);
and U6497 (N_6497,N_5538,N_5980);
and U6498 (N_6498,N_5968,N_5825);
nand U6499 (N_6499,N_5505,N_5591);
nand U6500 (N_6500,N_6491,N_6145);
nand U6501 (N_6501,N_6488,N_6307);
nor U6502 (N_6502,N_6294,N_6258);
nand U6503 (N_6503,N_6462,N_6387);
and U6504 (N_6504,N_6003,N_6256);
or U6505 (N_6505,N_6227,N_6004);
or U6506 (N_6506,N_6395,N_6419);
or U6507 (N_6507,N_6349,N_6239);
or U6508 (N_6508,N_6441,N_6490);
xnor U6509 (N_6509,N_6305,N_6034);
xnor U6510 (N_6510,N_6027,N_6368);
and U6511 (N_6511,N_6377,N_6344);
and U6512 (N_6512,N_6206,N_6357);
or U6513 (N_6513,N_6224,N_6161);
nor U6514 (N_6514,N_6182,N_6235);
nand U6515 (N_6515,N_6121,N_6476);
nor U6516 (N_6516,N_6089,N_6383);
nor U6517 (N_6517,N_6229,N_6303);
and U6518 (N_6518,N_6168,N_6365);
or U6519 (N_6519,N_6468,N_6273);
nor U6520 (N_6520,N_6404,N_6405);
and U6521 (N_6521,N_6262,N_6088);
or U6522 (N_6522,N_6336,N_6246);
or U6523 (N_6523,N_6345,N_6274);
and U6524 (N_6524,N_6181,N_6080);
or U6525 (N_6525,N_6270,N_6021);
nor U6526 (N_6526,N_6077,N_6087);
nand U6527 (N_6527,N_6031,N_6352);
or U6528 (N_6528,N_6030,N_6110);
or U6529 (N_6529,N_6327,N_6390);
nor U6530 (N_6530,N_6183,N_6009);
xnor U6531 (N_6531,N_6407,N_6165);
nor U6532 (N_6532,N_6485,N_6230);
nor U6533 (N_6533,N_6221,N_6363);
nand U6534 (N_6534,N_6118,N_6494);
nand U6535 (N_6535,N_6474,N_6127);
or U6536 (N_6536,N_6310,N_6373);
nor U6537 (N_6537,N_6319,N_6228);
nand U6538 (N_6538,N_6320,N_6451);
and U6539 (N_6539,N_6125,N_6108);
nor U6540 (N_6540,N_6140,N_6210);
or U6541 (N_6541,N_6284,N_6251);
and U6542 (N_6542,N_6219,N_6142);
or U6543 (N_6543,N_6259,N_6151);
nand U6544 (N_6544,N_6185,N_6112);
nor U6545 (N_6545,N_6130,N_6323);
nand U6546 (N_6546,N_6155,N_6166);
or U6547 (N_6547,N_6209,N_6301);
nor U6548 (N_6548,N_6283,N_6374);
nor U6549 (N_6549,N_6314,N_6267);
and U6550 (N_6550,N_6146,N_6448);
nand U6551 (N_6551,N_6047,N_6137);
nor U6552 (N_6552,N_6300,N_6060);
or U6553 (N_6553,N_6065,N_6215);
nor U6554 (N_6554,N_6343,N_6340);
nor U6555 (N_6555,N_6296,N_6286);
or U6556 (N_6556,N_6147,N_6237);
nor U6557 (N_6557,N_6134,N_6200);
nor U6558 (N_6558,N_6226,N_6138);
nand U6559 (N_6559,N_6333,N_6434);
nor U6560 (N_6560,N_6175,N_6271);
nand U6561 (N_6561,N_6298,N_6417);
or U6562 (N_6562,N_6457,N_6002);
nor U6563 (N_6563,N_6094,N_6356);
and U6564 (N_6564,N_6443,N_6433);
nor U6565 (N_6565,N_6478,N_6119);
and U6566 (N_6566,N_6334,N_6008);
or U6567 (N_6567,N_6317,N_6430);
and U6568 (N_6568,N_6269,N_6242);
or U6569 (N_6569,N_6152,N_6326);
nor U6570 (N_6570,N_6391,N_6392);
xnor U6571 (N_6571,N_6055,N_6139);
xor U6572 (N_6572,N_6465,N_6136);
nor U6573 (N_6573,N_6149,N_6062);
and U6574 (N_6574,N_6007,N_6156);
and U6575 (N_6575,N_6299,N_6445);
nand U6576 (N_6576,N_6109,N_6222);
nor U6577 (N_6577,N_6176,N_6346);
xor U6578 (N_6578,N_6086,N_6179);
xor U6579 (N_6579,N_6042,N_6481);
or U6580 (N_6580,N_6464,N_6281);
or U6581 (N_6581,N_6420,N_6187);
or U6582 (N_6582,N_6066,N_6456);
nand U6583 (N_6583,N_6389,N_6359);
and U6584 (N_6584,N_6347,N_6120);
or U6585 (N_6585,N_6107,N_6201);
nand U6586 (N_6586,N_6382,N_6372);
nor U6587 (N_6587,N_6249,N_6331);
xnor U6588 (N_6588,N_6074,N_6339);
nand U6589 (N_6589,N_6102,N_6350);
nand U6590 (N_6590,N_6059,N_6297);
or U6591 (N_6591,N_6098,N_6467);
xnor U6592 (N_6592,N_6038,N_6067);
nor U6593 (N_6593,N_6208,N_6260);
or U6594 (N_6594,N_6424,N_6243);
nand U6595 (N_6595,N_6264,N_6045);
xor U6596 (N_6596,N_6411,N_6489);
nor U6597 (N_6597,N_6483,N_6452);
or U6598 (N_6598,N_6495,N_6068);
xor U6599 (N_6599,N_6380,N_6154);
nand U6600 (N_6600,N_6033,N_6036);
nand U6601 (N_6601,N_6435,N_6348);
or U6602 (N_6602,N_6289,N_6397);
or U6603 (N_6603,N_6124,N_6385);
nor U6604 (N_6604,N_6282,N_6414);
and U6605 (N_6605,N_6220,N_6313);
xnor U6606 (N_6606,N_6399,N_6085);
or U6607 (N_6607,N_6308,N_6095);
or U6608 (N_6608,N_6158,N_6439);
nand U6609 (N_6609,N_6263,N_6453);
nand U6610 (N_6610,N_6225,N_6254);
nor U6611 (N_6611,N_6255,N_6436);
or U6612 (N_6612,N_6113,N_6214);
nand U6613 (N_6613,N_6497,N_6160);
nor U6614 (N_6614,N_6261,N_6223);
nand U6615 (N_6615,N_6232,N_6437);
and U6616 (N_6616,N_6431,N_6213);
and U6617 (N_6617,N_6278,N_6005);
nor U6618 (N_6618,N_6234,N_6398);
nor U6619 (N_6619,N_6290,N_6469);
or U6620 (N_6620,N_6090,N_6167);
nor U6621 (N_6621,N_6370,N_6001);
xor U6622 (N_6622,N_6091,N_6361);
nor U6623 (N_6623,N_6403,N_6204);
nand U6624 (N_6624,N_6071,N_6479);
nor U6625 (N_6625,N_6024,N_6133);
or U6626 (N_6626,N_6114,N_6178);
nand U6627 (N_6627,N_6216,N_6432);
nor U6628 (N_6628,N_6444,N_6360);
nor U6629 (N_6629,N_6063,N_6366);
nand U6630 (N_6630,N_6293,N_6426);
nand U6631 (N_6631,N_6324,N_6455);
and U6632 (N_6632,N_6174,N_6078);
nor U6633 (N_6633,N_6014,N_6440);
and U6634 (N_6634,N_6409,N_6194);
or U6635 (N_6635,N_6484,N_6315);
or U6636 (N_6636,N_6381,N_6044);
and U6637 (N_6637,N_6266,N_6072);
or U6638 (N_6638,N_6459,N_6438);
nor U6639 (N_6639,N_6212,N_6265);
or U6640 (N_6640,N_6449,N_6203);
nor U6641 (N_6641,N_6351,N_6020);
or U6642 (N_6642,N_6141,N_6231);
or U6643 (N_6643,N_6442,N_6416);
nand U6644 (N_6644,N_6364,N_6247);
xor U6645 (N_6645,N_6458,N_6394);
nor U6646 (N_6646,N_6367,N_6472);
nor U6647 (N_6647,N_6000,N_6253);
nor U6648 (N_6648,N_6499,N_6032);
and U6649 (N_6649,N_6410,N_6454);
nor U6650 (N_6650,N_6013,N_6429);
xor U6651 (N_6651,N_6292,N_6084);
nand U6652 (N_6652,N_6016,N_6126);
and U6653 (N_6653,N_6169,N_6006);
nand U6654 (N_6654,N_6035,N_6309);
xor U6655 (N_6655,N_6241,N_6279);
and U6656 (N_6656,N_6048,N_6257);
nor U6657 (N_6657,N_6097,N_6069);
and U6658 (N_6658,N_6353,N_6143);
xnor U6659 (N_6659,N_6135,N_6362);
xnor U6660 (N_6660,N_6379,N_6199);
nand U6661 (N_6661,N_6358,N_6040);
nor U6662 (N_6662,N_6498,N_6422);
and U6663 (N_6663,N_6025,N_6192);
and U6664 (N_6664,N_6218,N_6184);
and U6665 (N_6665,N_6487,N_6460);
xor U6666 (N_6666,N_6415,N_6163);
or U6667 (N_6667,N_6012,N_6144);
nand U6668 (N_6668,N_6285,N_6295);
xor U6669 (N_6669,N_6196,N_6217);
and U6670 (N_6670,N_6116,N_6341);
or U6671 (N_6671,N_6191,N_6190);
xor U6672 (N_6672,N_6193,N_6401);
nor U6673 (N_6673,N_6207,N_6238);
nor U6674 (N_6674,N_6164,N_6486);
nand U6675 (N_6675,N_6475,N_6276);
nor U6676 (N_6676,N_6202,N_6096);
nor U6677 (N_6677,N_6450,N_6418);
or U6678 (N_6678,N_6287,N_6250);
nand U6679 (N_6679,N_6277,N_6412);
nand U6680 (N_6680,N_6354,N_6150);
or U6681 (N_6681,N_6342,N_6172);
or U6682 (N_6682,N_6131,N_6316);
or U6683 (N_6683,N_6393,N_6318);
nor U6684 (N_6684,N_6369,N_6322);
or U6685 (N_6685,N_6010,N_6471);
and U6686 (N_6686,N_6245,N_6105);
or U6687 (N_6687,N_6101,N_6043);
and U6688 (N_6688,N_6017,N_6321);
nand U6689 (N_6689,N_6054,N_6082);
and U6690 (N_6690,N_6400,N_6470);
and U6691 (N_6691,N_6328,N_6335);
nand U6692 (N_6692,N_6064,N_6236);
xnor U6693 (N_6693,N_6180,N_6244);
or U6694 (N_6694,N_6122,N_6029);
or U6695 (N_6695,N_6076,N_6157);
nor U6696 (N_6696,N_6325,N_6058);
nand U6697 (N_6697,N_6177,N_6466);
and U6698 (N_6698,N_6428,N_6473);
nand U6699 (N_6699,N_6026,N_6378);
xnor U6700 (N_6700,N_6492,N_6022);
or U6701 (N_6701,N_6148,N_6197);
and U6702 (N_6702,N_6018,N_6106);
and U6703 (N_6703,N_6446,N_6115);
nor U6704 (N_6704,N_6376,N_6195);
nor U6705 (N_6705,N_6050,N_6153);
xnor U6706 (N_6706,N_6388,N_6482);
and U6707 (N_6707,N_6103,N_6123);
nor U6708 (N_6708,N_6371,N_6070);
and U6709 (N_6709,N_6111,N_6100);
or U6710 (N_6710,N_6015,N_6051);
and U6711 (N_6711,N_6480,N_6011);
nor U6712 (N_6712,N_6198,N_6205);
nor U6713 (N_6713,N_6421,N_6425);
and U6714 (N_6714,N_6384,N_6132);
nor U6715 (N_6715,N_6280,N_6117);
nor U6716 (N_6716,N_6463,N_6046);
and U6717 (N_6717,N_6447,N_6311);
or U6718 (N_6718,N_6083,N_6355);
or U6719 (N_6719,N_6159,N_6337);
nor U6720 (N_6720,N_6306,N_6170);
nand U6721 (N_6721,N_6332,N_6252);
and U6722 (N_6722,N_6396,N_6081);
xor U6723 (N_6723,N_6268,N_6427);
or U6724 (N_6724,N_6288,N_6052);
nand U6725 (N_6725,N_6275,N_6240);
xor U6726 (N_6726,N_6248,N_6329);
and U6727 (N_6727,N_6056,N_6162);
nor U6728 (N_6728,N_6338,N_6019);
nor U6729 (N_6729,N_6493,N_6496);
nand U6730 (N_6730,N_6039,N_6189);
and U6731 (N_6731,N_6173,N_6171);
and U6732 (N_6732,N_6041,N_6188);
nor U6733 (N_6733,N_6211,N_6386);
xor U6734 (N_6734,N_6408,N_6304);
or U6735 (N_6735,N_6053,N_6128);
and U6736 (N_6736,N_6272,N_6302);
and U6737 (N_6737,N_6099,N_6092);
or U6738 (N_6738,N_6291,N_6406);
nand U6739 (N_6739,N_6461,N_6049);
or U6740 (N_6740,N_6330,N_6423);
nand U6741 (N_6741,N_6129,N_6186);
or U6742 (N_6742,N_6023,N_6477);
and U6743 (N_6743,N_6075,N_6073);
nand U6744 (N_6744,N_6413,N_6312);
nor U6745 (N_6745,N_6037,N_6104);
or U6746 (N_6746,N_6233,N_6402);
nor U6747 (N_6747,N_6028,N_6057);
xor U6748 (N_6748,N_6375,N_6093);
or U6749 (N_6749,N_6079,N_6061);
xor U6750 (N_6750,N_6053,N_6133);
xnor U6751 (N_6751,N_6012,N_6203);
xor U6752 (N_6752,N_6322,N_6012);
xnor U6753 (N_6753,N_6059,N_6129);
nor U6754 (N_6754,N_6382,N_6479);
and U6755 (N_6755,N_6321,N_6499);
and U6756 (N_6756,N_6081,N_6242);
nor U6757 (N_6757,N_6235,N_6200);
or U6758 (N_6758,N_6126,N_6376);
nand U6759 (N_6759,N_6002,N_6404);
nand U6760 (N_6760,N_6468,N_6229);
and U6761 (N_6761,N_6206,N_6461);
nor U6762 (N_6762,N_6125,N_6499);
nand U6763 (N_6763,N_6048,N_6413);
or U6764 (N_6764,N_6482,N_6400);
nand U6765 (N_6765,N_6021,N_6110);
nand U6766 (N_6766,N_6496,N_6156);
nand U6767 (N_6767,N_6148,N_6336);
or U6768 (N_6768,N_6189,N_6076);
or U6769 (N_6769,N_6182,N_6035);
nand U6770 (N_6770,N_6227,N_6020);
or U6771 (N_6771,N_6031,N_6213);
or U6772 (N_6772,N_6479,N_6030);
nand U6773 (N_6773,N_6098,N_6145);
nand U6774 (N_6774,N_6255,N_6470);
nor U6775 (N_6775,N_6255,N_6332);
nor U6776 (N_6776,N_6438,N_6312);
nor U6777 (N_6777,N_6201,N_6005);
nor U6778 (N_6778,N_6426,N_6016);
nand U6779 (N_6779,N_6281,N_6479);
and U6780 (N_6780,N_6127,N_6259);
or U6781 (N_6781,N_6492,N_6234);
and U6782 (N_6782,N_6153,N_6454);
or U6783 (N_6783,N_6115,N_6454);
nor U6784 (N_6784,N_6174,N_6429);
and U6785 (N_6785,N_6452,N_6478);
nor U6786 (N_6786,N_6088,N_6126);
nand U6787 (N_6787,N_6040,N_6299);
nand U6788 (N_6788,N_6019,N_6128);
nor U6789 (N_6789,N_6105,N_6303);
nor U6790 (N_6790,N_6168,N_6146);
and U6791 (N_6791,N_6060,N_6357);
and U6792 (N_6792,N_6264,N_6404);
nand U6793 (N_6793,N_6038,N_6259);
and U6794 (N_6794,N_6351,N_6320);
and U6795 (N_6795,N_6381,N_6012);
and U6796 (N_6796,N_6031,N_6141);
and U6797 (N_6797,N_6245,N_6058);
xnor U6798 (N_6798,N_6271,N_6453);
nand U6799 (N_6799,N_6457,N_6355);
nor U6800 (N_6800,N_6387,N_6147);
and U6801 (N_6801,N_6300,N_6315);
or U6802 (N_6802,N_6164,N_6062);
nand U6803 (N_6803,N_6121,N_6015);
nand U6804 (N_6804,N_6404,N_6115);
and U6805 (N_6805,N_6192,N_6064);
nand U6806 (N_6806,N_6201,N_6067);
and U6807 (N_6807,N_6080,N_6290);
nand U6808 (N_6808,N_6420,N_6467);
or U6809 (N_6809,N_6417,N_6120);
and U6810 (N_6810,N_6204,N_6299);
xnor U6811 (N_6811,N_6419,N_6256);
or U6812 (N_6812,N_6050,N_6074);
or U6813 (N_6813,N_6064,N_6462);
nand U6814 (N_6814,N_6040,N_6456);
nand U6815 (N_6815,N_6297,N_6002);
nand U6816 (N_6816,N_6402,N_6037);
xnor U6817 (N_6817,N_6137,N_6466);
xor U6818 (N_6818,N_6171,N_6061);
nor U6819 (N_6819,N_6049,N_6367);
nor U6820 (N_6820,N_6272,N_6064);
and U6821 (N_6821,N_6091,N_6429);
nand U6822 (N_6822,N_6154,N_6406);
nor U6823 (N_6823,N_6150,N_6210);
nor U6824 (N_6824,N_6381,N_6000);
nor U6825 (N_6825,N_6199,N_6186);
and U6826 (N_6826,N_6157,N_6441);
or U6827 (N_6827,N_6376,N_6377);
nor U6828 (N_6828,N_6231,N_6448);
and U6829 (N_6829,N_6334,N_6298);
nand U6830 (N_6830,N_6102,N_6097);
nand U6831 (N_6831,N_6470,N_6210);
nand U6832 (N_6832,N_6238,N_6099);
or U6833 (N_6833,N_6453,N_6018);
and U6834 (N_6834,N_6318,N_6084);
or U6835 (N_6835,N_6233,N_6337);
or U6836 (N_6836,N_6315,N_6347);
xnor U6837 (N_6837,N_6410,N_6382);
nand U6838 (N_6838,N_6124,N_6111);
nor U6839 (N_6839,N_6435,N_6308);
or U6840 (N_6840,N_6174,N_6478);
and U6841 (N_6841,N_6363,N_6052);
nor U6842 (N_6842,N_6451,N_6450);
and U6843 (N_6843,N_6069,N_6053);
xor U6844 (N_6844,N_6299,N_6237);
and U6845 (N_6845,N_6465,N_6376);
and U6846 (N_6846,N_6171,N_6332);
nor U6847 (N_6847,N_6441,N_6476);
nor U6848 (N_6848,N_6419,N_6044);
nand U6849 (N_6849,N_6307,N_6410);
xor U6850 (N_6850,N_6299,N_6375);
xnor U6851 (N_6851,N_6364,N_6385);
and U6852 (N_6852,N_6034,N_6362);
nor U6853 (N_6853,N_6286,N_6431);
and U6854 (N_6854,N_6205,N_6352);
and U6855 (N_6855,N_6095,N_6272);
nor U6856 (N_6856,N_6023,N_6156);
and U6857 (N_6857,N_6165,N_6036);
or U6858 (N_6858,N_6266,N_6162);
or U6859 (N_6859,N_6311,N_6380);
and U6860 (N_6860,N_6266,N_6387);
and U6861 (N_6861,N_6449,N_6263);
nor U6862 (N_6862,N_6274,N_6217);
and U6863 (N_6863,N_6208,N_6447);
nand U6864 (N_6864,N_6076,N_6316);
nor U6865 (N_6865,N_6172,N_6190);
and U6866 (N_6866,N_6181,N_6157);
or U6867 (N_6867,N_6158,N_6237);
xor U6868 (N_6868,N_6084,N_6487);
and U6869 (N_6869,N_6093,N_6371);
xor U6870 (N_6870,N_6394,N_6070);
and U6871 (N_6871,N_6275,N_6054);
or U6872 (N_6872,N_6271,N_6133);
and U6873 (N_6873,N_6270,N_6225);
nor U6874 (N_6874,N_6240,N_6257);
or U6875 (N_6875,N_6353,N_6435);
nor U6876 (N_6876,N_6447,N_6025);
or U6877 (N_6877,N_6421,N_6049);
nand U6878 (N_6878,N_6450,N_6117);
and U6879 (N_6879,N_6311,N_6373);
nand U6880 (N_6880,N_6196,N_6027);
and U6881 (N_6881,N_6255,N_6421);
nor U6882 (N_6882,N_6021,N_6312);
nand U6883 (N_6883,N_6082,N_6205);
nand U6884 (N_6884,N_6393,N_6054);
nand U6885 (N_6885,N_6321,N_6278);
nand U6886 (N_6886,N_6116,N_6273);
and U6887 (N_6887,N_6236,N_6051);
nor U6888 (N_6888,N_6474,N_6479);
xor U6889 (N_6889,N_6226,N_6112);
nor U6890 (N_6890,N_6416,N_6394);
and U6891 (N_6891,N_6199,N_6150);
nand U6892 (N_6892,N_6462,N_6235);
nor U6893 (N_6893,N_6338,N_6161);
nor U6894 (N_6894,N_6293,N_6049);
nor U6895 (N_6895,N_6439,N_6210);
or U6896 (N_6896,N_6469,N_6463);
xor U6897 (N_6897,N_6103,N_6357);
nor U6898 (N_6898,N_6288,N_6155);
nor U6899 (N_6899,N_6450,N_6266);
xnor U6900 (N_6900,N_6290,N_6101);
xor U6901 (N_6901,N_6070,N_6425);
xnor U6902 (N_6902,N_6242,N_6429);
xor U6903 (N_6903,N_6050,N_6465);
nand U6904 (N_6904,N_6133,N_6175);
xor U6905 (N_6905,N_6142,N_6452);
nand U6906 (N_6906,N_6497,N_6025);
nor U6907 (N_6907,N_6486,N_6124);
xnor U6908 (N_6908,N_6329,N_6019);
nor U6909 (N_6909,N_6135,N_6358);
nand U6910 (N_6910,N_6272,N_6286);
and U6911 (N_6911,N_6347,N_6061);
nor U6912 (N_6912,N_6129,N_6497);
xor U6913 (N_6913,N_6390,N_6097);
or U6914 (N_6914,N_6439,N_6049);
nand U6915 (N_6915,N_6081,N_6418);
nor U6916 (N_6916,N_6268,N_6462);
nor U6917 (N_6917,N_6213,N_6476);
nand U6918 (N_6918,N_6461,N_6400);
nand U6919 (N_6919,N_6139,N_6248);
nor U6920 (N_6920,N_6050,N_6228);
nor U6921 (N_6921,N_6032,N_6074);
nor U6922 (N_6922,N_6189,N_6085);
nand U6923 (N_6923,N_6313,N_6288);
and U6924 (N_6924,N_6327,N_6085);
and U6925 (N_6925,N_6315,N_6190);
nor U6926 (N_6926,N_6359,N_6115);
nor U6927 (N_6927,N_6497,N_6118);
or U6928 (N_6928,N_6177,N_6481);
and U6929 (N_6929,N_6075,N_6416);
xor U6930 (N_6930,N_6237,N_6396);
and U6931 (N_6931,N_6314,N_6435);
or U6932 (N_6932,N_6353,N_6261);
nand U6933 (N_6933,N_6051,N_6166);
nor U6934 (N_6934,N_6172,N_6494);
or U6935 (N_6935,N_6360,N_6232);
xnor U6936 (N_6936,N_6213,N_6148);
nor U6937 (N_6937,N_6482,N_6288);
nor U6938 (N_6938,N_6329,N_6026);
nor U6939 (N_6939,N_6064,N_6248);
nand U6940 (N_6940,N_6496,N_6235);
nor U6941 (N_6941,N_6259,N_6021);
or U6942 (N_6942,N_6286,N_6404);
and U6943 (N_6943,N_6247,N_6420);
nor U6944 (N_6944,N_6285,N_6031);
nand U6945 (N_6945,N_6385,N_6334);
or U6946 (N_6946,N_6133,N_6366);
or U6947 (N_6947,N_6109,N_6396);
nand U6948 (N_6948,N_6183,N_6276);
or U6949 (N_6949,N_6082,N_6496);
and U6950 (N_6950,N_6229,N_6239);
nor U6951 (N_6951,N_6176,N_6246);
and U6952 (N_6952,N_6490,N_6343);
nand U6953 (N_6953,N_6232,N_6016);
xnor U6954 (N_6954,N_6170,N_6202);
nor U6955 (N_6955,N_6144,N_6364);
nor U6956 (N_6956,N_6002,N_6369);
or U6957 (N_6957,N_6423,N_6027);
or U6958 (N_6958,N_6449,N_6247);
nor U6959 (N_6959,N_6297,N_6466);
or U6960 (N_6960,N_6101,N_6117);
and U6961 (N_6961,N_6002,N_6154);
or U6962 (N_6962,N_6104,N_6332);
nor U6963 (N_6963,N_6031,N_6405);
nor U6964 (N_6964,N_6288,N_6301);
nand U6965 (N_6965,N_6401,N_6366);
or U6966 (N_6966,N_6497,N_6361);
nor U6967 (N_6967,N_6163,N_6214);
and U6968 (N_6968,N_6499,N_6297);
and U6969 (N_6969,N_6380,N_6306);
and U6970 (N_6970,N_6305,N_6174);
nor U6971 (N_6971,N_6294,N_6076);
and U6972 (N_6972,N_6246,N_6052);
nor U6973 (N_6973,N_6118,N_6274);
nand U6974 (N_6974,N_6439,N_6368);
or U6975 (N_6975,N_6149,N_6079);
nor U6976 (N_6976,N_6289,N_6266);
xor U6977 (N_6977,N_6348,N_6445);
or U6978 (N_6978,N_6309,N_6296);
or U6979 (N_6979,N_6115,N_6274);
xnor U6980 (N_6980,N_6059,N_6409);
nor U6981 (N_6981,N_6291,N_6382);
nor U6982 (N_6982,N_6130,N_6471);
or U6983 (N_6983,N_6201,N_6291);
nand U6984 (N_6984,N_6388,N_6117);
or U6985 (N_6985,N_6313,N_6194);
and U6986 (N_6986,N_6371,N_6271);
or U6987 (N_6987,N_6324,N_6337);
or U6988 (N_6988,N_6022,N_6141);
xor U6989 (N_6989,N_6358,N_6000);
nand U6990 (N_6990,N_6313,N_6199);
or U6991 (N_6991,N_6312,N_6326);
or U6992 (N_6992,N_6189,N_6121);
nor U6993 (N_6993,N_6353,N_6213);
nand U6994 (N_6994,N_6337,N_6296);
nand U6995 (N_6995,N_6017,N_6081);
and U6996 (N_6996,N_6228,N_6271);
or U6997 (N_6997,N_6300,N_6214);
and U6998 (N_6998,N_6189,N_6277);
nand U6999 (N_6999,N_6092,N_6315);
nand U7000 (N_7000,N_6897,N_6594);
nor U7001 (N_7001,N_6538,N_6890);
or U7002 (N_7002,N_6543,N_6647);
nor U7003 (N_7003,N_6930,N_6631);
nor U7004 (N_7004,N_6925,N_6644);
nand U7005 (N_7005,N_6915,N_6593);
nor U7006 (N_7006,N_6696,N_6792);
nor U7007 (N_7007,N_6699,N_6733);
or U7008 (N_7008,N_6660,N_6682);
nor U7009 (N_7009,N_6749,N_6928);
nand U7010 (N_7010,N_6615,N_6746);
nand U7011 (N_7011,N_6941,N_6921);
xnor U7012 (N_7012,N_6542,N_6507);
and U7013 (N_7013,N_6949,N_6595);
or U7014 (N_7014,N_6689,N_6757);
or U7015 (N_7015,N_6790,N_6501);
nor U7016 (N_7016,N_6772,N_6681);
or U7017 (N_7017,N_6828,N_6807);
nor U7018 (N_7018,N_6835,N_6683);
nor U7019 (N_7019,N_6520,N_6996);
and U7020 (N_7020,N_6803,N_6658);
nor U7021 (N_7021,N_6611,N_6555);
nor U7022 (N_7022,N_6609,N_6731);
or U7023 (N_7023,N_6574,N_6766);
or U7024 (N_7024,N_6767,N_6533);
and U7025 (N_7025,N_6843,N_6840);
nand U7026 (N_7026,N_6550,N_6991);
nand U7027 (N_7027,N_6859,N_6986);
and U7028 (N_7028,N_6848,N_6794);
nand U7029 (N_7029,N_6971,N_6976);
and U7030 (N_7030,N_6561,N_6721);
or U7031 (N_7031,N_6628,N_6623);
or U7032 (N_7032,N_6619,N_6858);
nor U7033 (N_7033,N_6704,N_6761);
and U7034 (N_7034,N_6521,N_6978);
or U7035 (N_7035,N_6862,N_6977);
and U7036 (N_7036,N_6950,N_6529);
xnor U7037 (N_7037,N_6717,N_6518);
xnor U7038 (N_7038,N_6571,N_6936);
and U7039 (N_7039,N_6815,N_6750);
or U7040 (N_7040,N_6729,N_6566);
nand U7041 (N_7041,N_6888,N_6982);
and U7042 (N_7042,N_6500,N_6821);
or U7043 (N_7043,N_6741,N_6714);
or U7044 (N_7044,N_6706,N_6760);
nor U7045 (N_7045,N_6988,N_6612);
nor U7046 (N_7046,N_6908,N_6808);
nand U7047 (N_7047,N_6811,N_6953);
or U7048 (N_7048,N_6680,N_6563);
nand U7049 (N_7049,N_6919,N_6748);
nand U7050 (N_7050,N_6869,N_6942);
and U7051 (N_7051,N_6938,N_6514);
or U7052 (N_7052,N_6702,N_6802);
and U7053 (N_7053,N_6643,N_6670);
nand U7054 (N_7054,N_6512,N_6819);
nand U7055 (N_7055,N_6759,N_6810);
and U7056 (N_7056,N_6943,N_6678);
nor U7057 (N_7057,N_6684,N_6713);
or U7058 (N_7058,N_6637,N_6535);
and U7059 (N_7059,N_6944,N_6620);
nor U7060 (N_7060,N_6532,N_6645);
and U7061 (N_7061,N_6567,N_6534);
or U7062 (N_7062,N_6974,N_6562);
or U7063 (N_7063,N_6722,N_6753);
or U7064 (N_7064,N_6738,N_6509);
or U7065 (N_7065,N_6958,N_6674);
nand U7066 (N_7066,N_6822,N_6824);
and U7067 (N_7067,N_6607,N_6614);
nand U7068 (N_7068,N_6932,N_6565);
and U7069 (N_7069,N_6662,N_6723);
and U7070 (N_7070,N_6548,N_6876);
and U7071 (N_7071,N_6523,N_6906);
nor U7072 (N_7072,N_6575,N_6972);
nand U7073 (N_7073,N_6568,N_6719);
nor U7074 (N_7074,N_6804,N_6549);
and U7075 (N_7075,N_6724,N_6596);
nor U7076 (N_7076,N_6737,N_6629);
nand U7077 (N_7077,N_6646,N_6984);
and U7078 (N_7078,N_6918,N_6872);
and U7079 (N_7079,N_6875,N_6966);
and U7080 (N_7080,N_6933,N_6503);
and U7081 (N_7081,N_6911,N_6511);
nor U7082 (N_7082,N_6585,N_6954);
nor U7083 (N_7083,N_6831,N_6998);
xnor U7084 (N_7084,N_6960,N_6793);
nor U7085 (N_7085,N_6818,N_6798);
and U7086 (N_7086,N_6544,N_6912);
nand U7087 (N_7087,N_6904,N_6531);
nor U7088 (N_7088,N_6625,N_6913);
or U7089 (N_7089,N_6856,N_6539);
and U7090 (N_7090,N_6580,N_6554);
and U7091 (N_7091,N_6686,N_6700);
nor U7092 (N_7092,N_6636,N_6541);
xor U7093 (N_7093,N_6983,N_6718);
and U7094 (N_7094,N_6795,N_6981);
nand U7095 (N_7095,N_6837,N_6999);
nand U7096 (N_7096,N_6586,N_6886);
or U7097 (N_7097,N_6654,N_6652);
or U7098 (N_7098,N_6667,N_6854);
or U7099 (N_7099,N_6885,N_6616);
nor U7100 (N_7100,N_6598,N_6728);
nor U7101 (N_7101,N_6524,N_6774);
nand U7102 (N_7102,N_6602,N_6962);
or U7103 (N_7103,N_6841,N_6672);
nor U7104 (N_7104,N_6506,N_6877);
or U7105 (N_7105,N_6780,N_6707);
nand U7106 (N_7106,N_6703,N_6965);
nand U7107 (N_7107,N_6905,N_6832);
nor U7108 (N_7108,N_6902,N_6922);
nor U7109 (N_7109,N_6797,N_6517);
nand U7110 (N_7110,N_6515,N_6694);
and U7111 (N_7111,N_6909,N_6785);
nor U7112 (N_7112,N_6814,N_6677);
nor U7113 (N_7113,N_6838,N_6863);
and U7114 (N_7114,N_6676,N_6650);
nor U7115 (N_7115,N_6638,N_6924);
and U7116 (N_7116,N_6899,N_6553);
and U7117 (N_7117,N_6879,N_6603);
nor U7118 (N_7118,N_6964,N_6528);
nor U7119 (N_7119,N_6695,N_6659);
or U7120 (N_7120,N_6635,N_6881);
nor U7121 (N_7121,N_6587,N_6744);
or U7122 (N_7122,N_6675,N_6693);
xnor U7123 (N_7123,N_6970,N_6651);
nor U7124 (N_7124,N_6896,N_6963);
xor U7125 (N_7125,N_6923,N_6957);
and U7126 (N_7126,N_6784,N_6961);
nand U7127 (N_7127,N_6874,N_6851);
or U7128 (N_7128,N_6618,N_6861);
or U7129 (N_7129,N_6791,N_6648);
or U7130 (N_7130,N_6584,N_6882);
and U7131 (N_7131,N_6769,N_6685);
nand U7132 (N_7132,N_6871,N_6973);
and U7133 (N_7133,N_6864,N_6777);
or U7134 (N_7134,N_6985,N_6590);
nand U7135 (N_7135,N_6939,N_6935);
nand U7136 (N_7136,N_6513,N_6892);
nor U7137 (N_7137,N_6552,N_6855);
or U7138 (N_7138,N_6601,N_6758);
nor U7139 (N_7139,N_6556,N_6754);
or U7140 (N_7140,N_6765,N_6809);
nand U7141 (N_7141,N_6916,N_6947);
or U7142 (N_7142,N_6536,N_6557);
and U7143 (N_7143,N_6914,N_6632);
or U7144 (N_7144,N_6995,N_6679);
and U7145 (N_7145,N_6868,N_6505);
and U7146 (N_7146,N_6751,N_6917);
nand U7147 (N_7147,N_6829,N_6801);
nor U7148 (N_7148,N_6788,N_6573);
nand U7149 (N_7149,N_6716,N_6990);
xor U7150 (N_7150,N_6617,N_6727);
xnor U7151 (N_7151,N_6687,N_6697);
xnor U7152 (N_7152,N_6813,N_6730);
nand U7153 (N_7153,N_6641,N_6800);
nor U7154 (N_7154,N_6690,N_6903);
nand U7155 (N_7155,N_6889,N_6952);
or U7156 (N_7156,N_6987,N_6989);
nand U7157 (N_7157,N_6613,N_6663);
or U7158 (N_7158,N_6608,N_6867);
nand U7159 (N_7159,N_6664,N_6712);
and U7160 (N_7160,N_6673,N_6502);
and U7161 (N_7161,N_6900,N_6582);
and U7162 (N_7162,N_6599,N_6873);
nand U7163 (N_7163,N_6770,N_6993);
or U7164 (N_7164,N_6736,N_6768);
and U7165 (N_7165,N_6622,N_6526);
nor U7166 (N_7166,N_6830,N_6907);
and U7167 (N_7167,N_6893,N_6742);
nand U7168 (N_7168,N_6666,N_6934);
nand U7169 (N_7169,N_6711,N_6743);
and U7170 (N_7170,N_6715,N_6732);
nor U7171 (N_7171,N_6951,N_6853);
or U7172 (N_7172,N_6789,N_6865);
nand U7173 (N_7173,N_6570,N_6588);
nand U7174 (N_7174,N_6630,N_6852);
and U7175 (N_7175,N_6979,N_6895);
nor U7176 (N_7176,N_6519,N_6937);
nor U7177 (N_7177,N_6740,N_6649);
nor U7178 (N_7178,N_6583,N_6527);
or U7179 (N_7179,N_6734,N_6842);
or U7180 (N_7180,N_6726,N_6577);
nor U7181 (N_7181,N_6931,N_6833);
or U7182 (N_7182,N_6540,N_6787);
nor U7183 (N_7183,N_6834,N_6817);
and U7184 (N_7184,N_6870,N_6945);
nor U7185 (N_7185,N_6839,N_6516);
or U7186 (N_7186,N_6771,N_6551);
or U7187 (N_7187,N_6665,N_6569);
nor U7188 (N_7188,N_6655,N_6508);
nor U7189 (N_7189,N_6940,N_6735);
nor U7190 (N_7190,N_6698,N_6775);
nand U7191 (N_7191,N_6747,N_6847);
or U7192 (N_7192,N_6756,N_6806);
or U7193 (N_7193,N_6640,N_6600);
nor U7194 (N_7194,N_6816,N_6776);
nor U7195 (N_7195,N_6621,N_6688);
nand U7196 (N_7196,N_6796,N_6820);
and U7197 (N_7197,N_6762,N_6955);
nand U7198 (N_7198,N_6669,N_6605);
nor U7199 (N_7199,N_6642,N_6845);
nand U7200 (N_7200,N_6579,N_6967);
xnor U7201 (N_7201,N_6653,N_6671);
nand U7202 (N_7202,N_6846,N_6547);
xor U7203 (N_7203,N_6510,N_6720);
nand U7204 (N_7204,N_6825,N_6627);
and U7205 (N_7205,N_6606,N_6783);
and U7206 (N_7206,N_6812,N_6968);
nand U7207 (N_7207,N_6624,N_6849);
and U7208 (N_7208,N_6763,N_6564);
and U7209 (N_7209,N_6782,N_6626);
or U7210 (N_7210,N_6880,N_6927);
nor U7211 (N_7211,N_6826,N_6752);
nor U7212 (N_7212,N_6705,N_6764);
nor U7213 (N_7213,N_6891,N_6656);
nor U7214 (N_7214,N_6975,N_6725);
nand U7215 (N_7215,N_6572,N_6739);
nor U7216 (N_7216,N_6969,N_6589);
nand U7217 (N_7217,N_6633,N_6926);
nand U7218 (N_7218,N_6522,N_6545);
nor U7219 (N_7219,N_6910,N_6948);
and U7220 (N_7220,N_6558,N_6692);
or U7221 (N_7221,N_6592,N_6755);
nor U7222 (N_7222,N_6887,N_6581);
xnor U7223 (N_7223,N_6530,N_6884);
nor U7224 (N_7224,N_6778,N_6559);
xnor U7225 (N_7225,N_6560,N_6980);
or U7226 (N_7226,N_6597,N_6634);
and U7227 (N_7227,N_6857,N_6994);
or U7228 (N_7228,N_6850,N_6668);
nand U7229 (N_7229,N_6591,N_6946);
nand U7230 (N_7230,N_6959,N_6525);
nand U7231 (N_7231,N_6537,N_6691);
nor U7232 (N_7232,N_6860,N_6639);
nor U7233 (N_7233,N_6992,N_6844);
and U7234 (N_7234,N_6997,N_6701);
nor U7235 (N_7235,N_6929,N_6781);
or U7236 (N_7236,N_6898,N_6805);
or U7237 (N_7237,N_6657,N_6894);
and U7238 (N_7238,N_6827,N_6920);
or U7239 (N_7239,N_6956,N_6504);
and U7240 (N_7240,N_6786,N_6745);
nor U7241 (N_7241,N_6578,N_6883);
and U7242 (N_7242,N_6661,N_6878);
xor U7243 (N_7243,N_6708,N_6901);
nor U7244 (N_7244,N_6709,N_6823);
or U7245 (N_7245,N_6710,N_6576);
or U7246 (N_7246,N_6610,N_6546);
and U7247 (N_7247,N_6866,N_6604);
and U7248 (N_7248,N_6799,N_6836);
nand U7249 (N_7249,N_6773,N_6779);
or U7250 (N_7250,N_6567,N_6967);
nand U7251 (N_7251,N_6929,N_6628);
and U7252 (N_7252,N_6985,N_6816);
nand U7253 (N_7253,N_6547,N_6593);
nand U7254 (N_7254,N_6630,N_6824);
or U7255 (N_7255,N_6672,N_6502);
nand U7256 (N_7256,N_6639,N_6507);
or U7257 (N_7257,N_6672,N_6524);
nand U7258 (N_7258,N_6835,N_6855);
nor U7259 (N_7259,N_6519,N_6650);
or U7260 (N_7260,N_6797,N_6793);
nand U7261 (N_7261,N_6813,N_6995);
nand U7262 (N_7262,N_6534,N_6521);
and U7263 (N_7263,N_6737,N_6795);
or U7264 (N_7264,N_6793,N_6501);
nor U7265 (N_7265,N_6575,N_6733);
and U7266 (N_7266,N_6615,N_6776);
or U7267 (N_7267,N_6692,N_6502);
xnor U7268 (N_7268,N_6536,N_6970);
or U7269 (N_7269,N_6809,N_6797);
nor U7270 (N_7270,N_6963,N_6716);
and U7271 (N_7271,N_6537,N_6872);
xor U7272 (N_7272,N_6785,N_6817);
nand U7273 (N_7273,N_6512,N_6867);
nand U7274 (N_7274,N_6502,N_6600);
or U7275 (N_7275,N_6918,N_6928);
nor U7276 (N_7276,N_6535,N_6914);
nand U7277 (N_7277,N_6723,N_6650);
and U7278 (N_7278,N_6556,N_6702);
nor U7279 (N_7279,N_6692,N_6999);
nand U7280 (N_7280,N_6914,N_6833);
or U7281 (N_7281,N_6895,N_6694);
and U7282 (N_7282,N_6644,N_6626);
and U7283 (N_7283,N_6754,N_6928);
nor U7284 (N_7284,N_6911,N_6953);
or U7285 (N_7285,N_6782,N_6989);
nand U7286 (N_7286,N_6913,N_6684);
or U7287 (N_7287,N_6831,N_6809);
xor U7288 (N_7288,N_6678,N_6642);
or U7289 (N_7289,N_6991,N_6527);
or U7290 (N_7290,N_6539,N_6727);
xor U7291 (N_7291,N_6833,N_6589);
nand U7292 (N_7292,N_6938,N_6801);
nand U7293 (N_7293,N_6716,N_6701);
nor U7294 (N_7294,N_6689,N_6560);
and U7295 (N_7295,N_6966,N_6512);
or U7296 (N_7296,N_6836,N_6896);
nand U7297 (N_7297,N_6580,N_6969);
nor U7298 (N_7298,N_6607,N_6545);
nor U7299 (N_7299,N_6902,N_6545);
and U7300 (N_7300,N_6566,N_6646);
or U7301 (N_7301,N_6586,N_6558);
nor U7302 (N_7302,N_6798,N_6974);
nor U7303 (N_7303,N_6543,N_6561);
xor U7304 (N_7304,N_6764,N_6839);
nor U7305 (N_7305,N_6846,N_6706);
and U7306 (N_7306,N_6978,N_6667);
xnor U7307 (N_7307,N_6576,N_6786);
nor U7308 (N_7308,N_6563,N_6878);
or U7309 (N_7309,N_6946,N_6579);
and U7310 (N_7310,N_6790,N_6565);
nand U7311 (N_7311,N_6678,N_6965);
and U7312 (N_7312,N_6757,N_6627);
nand U7313 (N_7313,N_6875,N_6648);
nand U7314 (N_7314,N_6797,N_6834);
nand U7315 (N_7315,N_6969,N_6814);
nand U7316 (N_7316,N_6738,N_6532);
xnor U7317 (N_7317,N_6532,N_6865);
nand U7318 (N_7318,N_6784,N_6745);
nand U7319 (N_7319,N_6702,N_6886);
nor U7320 (N_7320,N_6932,N_6981);
nand U7321 (N_7321,N_6699,N_6650);
nand U7322 (N_7322,N_6572,N_6766);
and U7323 (N_7323,N_6856,N_6704);
nand U7324 (N_7324,N_6605,N_6743);
and U7325 (N_7325,N_6595,N_6509);
and U7326 (N_7326,N_6890,N_6717);
xnor U7327 (N_7327,N_6933,N_6684);
nand U7328 (N_7328,N_6568,N_6563);
nand U7329 (N_7329,N_6753,N_6802);
and U7330 (N_7330,N_6670,N_6669);
or U7331 (N_7331,N_6947,N_6888);
xnor U7332 (N_7332,N_6550,N_6990);
nand U7333 (N_7333,N_6563,N_6582);
or U7334 (N_7334,N_6642,N_6728);
nand U7335 (N_7335,N_6583,N_6552);
and U7336 (N_7336,N_6761,N_6686);
nand U7337 (N_7337,N_6696,N_6909);
nand U7338 (N_7338,N_6860,N_6924);
or U7339 (N_7339,N_6605,N_6747);
and U7340 (N_7340,N_6797,N_6534);
nor U7341 (N_7341,N_6519,N_6621);
and U7342 (N_7342,N_6841,N_6872);
nand U7343 (N_7343,N_6869,N_6812);
nand U7344 (N_7344,N_6820,N_6901);
xor U7345 (N_7345,N_6890,N_6938);
or U7346 (N_7346,N_6603,N_6549);
and U7347 (N_7347,N_6963,N_6600);
nand U7348 (N_7348,N_6555,N_6936);
or U7349 (N_7349,N_6702,N_6944);
and U7350 (N_7350,N_6616,N_6587);
nand U7351 (N_7351,N_6696,N_6852);
nand U7352 (N_7352,N_6906,N_6541);
and U7353 (N_7353,N_6895,N_6547);
and U7354 (N_7354,N_6752,N_6965);
or U7355 (N_7355,N_6859,N_6601);
or U7356 (N_7356,N_6777,N_6768);
and U7357 (N_7357,N_6931,N_6720);
and U7358 (N_7358,N_6615,N_6907);
xor U7359 (N_7359,N_6994,N_6595);
or U7360 (N_7360,N_6801,N_6685);
or U7361 (N_7361,N_6686,N_6685);
nor U7362 (N_7362,N_6623,N_6810);
nor U7363 (N_7363,N_6888,N_6804);
nand U7364 (N_7364,N_6555,N_6909);
nor U7365 (N_7365,N_6726,N_6825);
nand U7366 (N_7366,N_6773,N_6876);
nand U7367 (N_7367,N_6754,N_6640);
nand U7368 (N_7368,N_6558,N_6527);
nand U7369 (N_7369,N_6838,N_6801);
or U7370 (N_7370,N_6943,N_6879);
nand U7371 (N_7371,N_6874,N_6976);
nor U7372 (N_7372,N_6858,N_6790);
and U7373 (N_7373,N_6808,N_6738);
or U7374 (N_7374,N_6787,N_6882);
and U7375 (N_7375,N_6837,N_6806);
and U7376 (N_7376,N_6722,N_6607);
and U7377 (N_7377,N_6603,N_6555);
or U7378 (N_7378,N_6745,N_6876);
nand U7379 (N_7379,N_6722,N_6556);
and U7380 (N_7380,N_6540,N_6696);
xor U7381 (N_7381,N_6523,N_6971);
xnor U7382 (N_7382,N_6636,N_6941);
nand U7383 (N_7383,N_6818,N_6955);
nor U7384 (N_7384,N_6722,N_6529);
or U7385 (N_7385,N_6883,N_6701);
nor U7386 (N_7386,N_6505,N_6659);
or U7387 (N_7387,N_6882,N_6875);
and U7388 (N_7388,N_6696,N_6776);
nor U7389 (N_7389,N_6836,N_6888);
nor U7390 (N_7390,N_6782,N_6511);
and U7391 (N_7391,N_6876,N_6660);
or U7392 (N_7392,N_6569,N_6585);
or U7393 (N_7393,N_6761,N_6532);
nor U7394 (N_7394,N_6722,N_6614);
or U7395 (N_7395,N_6639,N_6765);
and U7396 (N_7396,N_6523,N_6658);
nor U7397 (N_7397,N_6629,N_6754);
or U7398 (N_7398,N_6580,N_6876);
and U7399 (N_7399,N_6988,N_6505);
nand U7400 (N_7400,N_6889,N_6713);
nor U7401 (N_7401,N_6978,N_6719);
nand U7402 (N_7402,N_6535,N_6544);
nand U7403 (N_7403,N_6556,N_6753);
and U7404 (N_7404,N_6822,N_6795);
nor U7405 (N_7405,N_6923,N_6609);
xnor U7406 (N_7406,N_6790,N_6875);
nor U7407 (N_7407,N_6902,N_6581);
nand U7408 (N_7408,N_6882,N_6895);
nand U7409 (N_7409,N_6770,N_6612);
and U7410 (N_7410,N_6742,N_6934);
nor U7411 (N_7411,N_6951,N_6781);
nor U7412 (N_7412,N_6849,N_6651);
nor U7413 (N_7413,N_6799,N_6846);
nor U7414 (N_7414,N_6892,N_6641);
xnor U7415 (N_7415,N_6500,N_6766);
or U7416 (N_7416,N_6889,N_6709);
nor U7417 (N_7417,N_6626,N_6746);
or U7418 (N_7418,N_6573,N_6946);
nor U7419 (N_7419,N_6903,N_6977);
nand U7420 (N_7420,N_6533,N_6773);
nor U7421 (N_7421,N_6819,N_6531);
nor U7422 (N_7422,N_6555,N_6544);
or U7423 (N_7423,N_6502,N_6955);
and U7424 (N_7424,N_6997,N_6922);
or U7425 (N_7425,N_6752,N_6775);
nand U7426 (N_7426,N_6627,N_6585);
or U7427 (N_7427,N_6591,N_6763);
xnor U7428 (N_7428,N_6931,N_6659);
and U7429 (N_7429,N_6766,N_6512);
nand U7430 (N_7430,N_6860,N_6833);
nand U7431 (N_7431,N_6960,N_6663);
or U7432 (N_7432,N_6769,N_6741);
or U7433 (N_7433,N_6652,N_6615);
and U7434 (N_7434,N_6530,N_6626);
nand U7435 (N_7435,N_6773,N_6515);
nor U7436 (N_7436,N_6562,N_6866);
and U7437 (N_7437,N_6608,N_6528);
or U7438 (N_7438,N_6945,N_6936);
or U7439 (N_7439,N_6937,N_6891);
nand U7440 (N_7440,N_6801,N_6724);
nand U7441 (N_7441,N_6921,N_6638);
or U7442 (N_7442,N_6733,N_6739);
and U7443 (N_7443,N_6949,N_6578);
or U7444 (N_7444,N_6551,N_6884);
xor U7445 (N_7445,N_6906,N_6767);
xnor U7446 (N_7446,N_6979,N_6609);
nor U7447 (N_7447,N_6897,N_6985);
or U7448 (N_7448,N_6962,N_6606);
nand U7449 (N_7449,N_6877,N_6754);
xor U7450 (N_7450,N_6729,N_6888);
nand U7451 (N_7451,N_6750,N_6837);
xnor U7452 (N_7452,N_6729,N_6591);
or U7453 (N_7453,N_6601,N_6541);
nor U7454 (N_7454,N_6809,N_6855);
or U7455 (N_7455,N_6643,N_6964);
nand U7456 (N_7456,N_6662,N_6793);
and U7457 (N_7457,N_6896,N_6887);
nor U7458 (N_7458,N_6520,N_6614);
nand U7459 (N_7459,N_6574,N_6500);
xnor U7460 (N_7460,N_6862,N_6832);
nor U7461 (N_7461,N_6711,N_6802);
nand U7462 (N_7462,N_6637,N_6520);
nor U7463 (N_7463,N_6742,N_6546);
or U7464 (N_7464,N_6942,N_6776);
and U7465 (N_7465,N_6590,N_6995);
nor U7466 (N_7466,N_6979,N_6698);
nor U7467 (N_7467,N_6625,N_6510);
nand U7468 (N_7468,N_6921,N_6728);
nand U7469 (N_7469,N_6877,N_6831);
nand U7470 (N_7470,N_6907,N_6714);
and U7471 (N_7471,N_6643,N_6865);
xnor U7472 (N_7472,N_6800,N_6659);
nand U7473 (N_7473,N_6828,N_6514);
nor U7474 (N_7474,N_6784,N_6552);
xnor U7475 (N_7475,N_6838,N_6793);
and U7476 (N_7476,N_6701,N_6934);
nand U7477 (N_7477,N_6537,N_6817);
or U7478 (N_7478,N_6964,N_6815);
nor U7479 (N_7479,N_6960,N_6686);
nand U7480 (N_7480,N_6820,N_6992);
and U7481 (N_7481,N_6768,N_6529);
nor U7482 (N_7482,N_6689,N_6692);
and U7483 (N_7483,N_6988,N_6881);
or U7484 (N_7484,N_6991,N_6776);
nor U7485 (N_7485,N_6934,N_6966);
nor U7486 (N_7486,N_6713,N_6542);
nor U7487 (N_7487,N_6677,N_6784);
nor U7488 (N_7488,N_6889,N_6971);
xor U7489 (N_7489,N_6578,N_6793);
and U7490 (N_7490,N_6619,N_6740);
nand U7491 (N_7491,N_6660,N_6805);
nand U7492 (N_7492,N_6545,N_6921);
nor U7493 (N_7493,N_6913,N_6545);
or U7494 (N_7494,N_6836,N_6636);
nand U7495 (N_7495,N_6985,N_6806);
xnor U7496 (N_7496,N_6837,N_6840);
nand U7497 (N_7497,N_6971,N_6773);
nand U7498 (N_7498,N_6792,N_6583);
and U7499 (N_7499,N_6732,N_6926);
nor U7500 (N_7500,N_7210,N_7004);
or U7501 (N_7501,N_7270,N_7146);
nor U7502 (N_7502,N_7472,N_7019);
nand U7503 (N_7503,N_7172,N_7195);
nor U7504 (N_7504,N_7257,N_7198);
nand U7505 (N_7505,N_7373,N_7462);
nand U7506 (N_7506,N_7309,N_7414);
xor U7507 (N_7507,N_7108,N_7178);
and U7508 (N_7508,N_7456,N_7349);
nor U7509 (N_7509,N_7293,N_7427);
and U7510 (N_7510,N_7048,N_7229);
or U7511 (N_7511,N_7356,N_7324);
nand U7512 (N_7512,N_7419,N_7377);
nand U7513 (N_7513,N_7221,N_7123);
nor U7514 (N_7514,N_7412,N_7245);
or U7515 (N_7515,N_7113,N_7128);
nand U7516 (N_7516,N_7188,N_7226);
nor U7517 (N_7517,N_7057,N_7460);
or U7518 (N_7518,N_7286,N_7050);
nand U7519 (N_7519,N_7042,N_7278);
nor U7520 (N_7520,N_7364,N_7209);
nand U7521 (N_7521,N_7211,N_7097);
nand U7522 (N_7522,N_7029,N_7081);
nor U7523 (N_7523,N_7134,N_7264);
nand U7524 (N_7524,N_7346,N_7441);
or U7525 (N_7525,N_7408,N_7492);
xnor U7526 (N_7526,N_7105,N_7085);
or U7527 (N_7527,N_7244,N_7459);
nand U7528 (N_7528,N_7475,N_7149);
nor U7529 (N_7529,N_7423,N_7145);
nand U7530 (N_7530,N_7398,N_7465);
or U7531 (N_7531,N_7409,N_7418);
and U7532 (N_7532,N_7480,N_7424);
xor U7533 (N_7533,N_7274,N_7322);
or U7534 (N_7534,N_7000,N_7199);
nand U7535 (N_7535,N_7137,N_7231);
nand U7536 (N_7536,N_7109,N_7086);
and U7537 (N_7537,N_7100,N_7069);
nor U7538 (N_7538,N_7115,N_7126);
xor U7539 (N_7539,N_7067,N_7101);
xnor U7540 (N_7540,N_7249,N_7442);
or U7541 (N_7541,N_7148,N_7341);
and U7542 (N_7542,N_7110,N_7489);
and U7543 (N_7543,N_7186,N_7432);
or U7544 (N_7544,N_7367,N_7215);
nor U7545 (N_7545,N_7045,N_7337);
and U7546 (N_7546,N_7080,N_7359);
and U7547 (N_7547,N_7079,N_7237);
nor U7548 (N_7548,N_7220,N_7205);
nand U7549 (N_7549,N_7248,N_7192);
and U7550 (N_7550,N_7203,N_7454);
nor U7551 (N_7551,N_7493,N_7151);
or U7552 (N_7552,N_7135,N_7162);
and U7553 (N_7553,N_7046,N_7160);
nand U7554 (N_7554,N_7425,N_7038);
xnor U7555 (N_7555,N_7259,N_7166);
and U7556 (N_7556,N_7252,N_7352);
nor U7557 (N_7557,N_7326,N_7066);
or U7558 (N_7558,N_7386,N_7173);
and U7559 (N_7559,N_7328,N_7007);
nand U7560 (N_7560,N_7315,N_7218);
or U7561 (N_7561,N_7474,N_7287);
and U7562 (N_7562,N_7167,N_7389);
nor U7563 (N_7563,N_7321,N_7091);
and U7564 (N_7564,N_7342,N_7375);
nand U7565 (N_7565,N_7329,N_7476);
xnor U7566 (N_7566,N_7376,N_7430);
or U7567 (N_7567,N_7217,N_7247);
nor U7568 (N_7568,N_7266,N_7301);
nand U7569 (N_7569,N_7457,N_7024);
nor U7570 (N_7570,N_7468,N_7020);
and U7571 (N_7571,N_7147,N_7494);
nor U7572 (N_7572,N_7275,N_7297);
and U7573 (N_7573,N_7250,N_7168);
or U7574 (N_7574,N_7305,N_7463);
or U7575 (N_7575,N_7095,N_7165);
xor U7576 (N_7576,N_7098,N_7345);
nand U7577 (N_7577,N_7005,N_7037);
nor U7578 (N_7578,N_7202,N_7455);
nand U7579 (N_7579,N_7406,N_7089);
nand U7580 (N_7580,N_7138,N_7204);
or U7581 (N_7581,N_7385,N_7490);
and U7582 (N_7582,N_7479,N_7331);
nor U7583 (N_7583,N_7272,N_7410);
or U7584 (N_7584,N_7399,N_7471);
and U7585 (N_7585,N_7319,N_7353);
and U7586 (N_7586,N_7267,N_7282);
and U7587 (N_7587,N_7285,N_7021);
and U7588 (N_7588,N_7082,N_7238);
and U7589 (N_7589,N_7429,N_7296);
or U7590 (N_7590,N_7200,N_7255);
and U7591 (N_7591,N_7362,N_7277);
nor U7592 (N_7592,N_7488,N_7180);
or U7593 (N_7593,N_7271,N_7347);
nor U7594 (N_7594,N_7018,N_7027);
nand U7595 (N_7595,N_7233,N_7336);
and U7596 (N_7596,N_7318,N_7054);
xnor U7597 (N_7597,N_7413,N_7022);
nand U7598 (N_7598,N_7496,N_7438);
nor U7599 (N_7599,N_7308,N_7119);
nand U7600 (N_7600,N_7458,N_7201);
or U7601 (N_7601,N_7451,N_7300);
nand U7602 (N_7602,N_7437,N_7295);
or U7603 (N_7603,N_7087,N_7360);
and U7604 (N_7604,N_7464,N_7302);
or U7605 (N_7605,N_7288,N_7372);
and U7606 (N_7606,N_7443,N_7461);
xnor U7607 (N_7607,N_7133,N_7394);
nand U7608 (N_7608,N_7339,N_7447);
xor U7609 (N_7609,N_7084,N_7121);
xor U7610 (N_7610,N_7403,N_7283);
xnor U7611 (N_7611,N_7235,N_7265);
nand U7612 (N_7612,N_7034,N_7120);
or U7613 (N_7613,N_7090,N_7156);
and U7614 (N_7614,N_7107,N_7382);
or U7615 (N_7615,N_7401,N_7491);
xnor U7616 (N_7616,N_7175,N_7263);
nand U7617 (N_7617,N_7106,N_7378);
or U7618 (N_7618,N_7068,N_7307);
and U7619 (N_7619,N_7365,N_7371);
nand U7620 (N_7620,N_7154,N_7348);
nor U7621 (N_7621,N_7466,N_7481);
xor U7622 (N_7622,N_7157,N_7290);
nor U7623 (N_7623,N_7239,N_7052);
nand U7624 (N_7624,N_7096,N_7150);
nor U7625 (N_7625,N_7473,N_7219);
and U7626 (N_7626,N_7258,N_7174);
and U7627 (N_7627,N_7152,N_7323);
nand U7628 (N_7628,N_7384,N_7040);
nor U7629 (N_7629,N_7312,N_7314);
nor U7630 (N_7630,N_7159,N_7072);
or U7631 (N_7631,N_7062,N_7189);
and U7632 (N_7632,N_7236,N_7182);
and U7633 (N_7633,N_7064,N_7453);
nand U7634 (N_7634,N_7390,N_7158);
or U7635 (N_7635,N_7338,N_7153);
and U7636 (N_7636,N_7125,N_7036);
nor U7637 (N_7637,N_7304,N_7484);
nand U7638 (N_7638,N_7388,N_7161);
and U7639 (N_7639,N_7313,N_7439);
and U7640 (N_7640,N_7495,N_7269);
nand U7641 (N_7641,N_7381,N_7142);
nand U7642 (N_7642,N_7369,N_7325);
xor U7643 (N_7643,N_7332,N_7032);
nand U7644 (N_7644,N_7224,N_7063);
nor U7645 (N_7645,N_7433,N_7363);
nand U7646 (N_7646,N_7370,N_7404);
nor U7647 (N_7647,N_7392,N_7051);
nand U7648 (N_7648,N_7444,N_7061);
nand U7649 (N_7649,N_7104,N_7099);
nor U7650 (N_7650,N_7289,N_7228);
or U7651 (N_7651,N_7074,N_7065);
and U7652 (N_7652,N_7094,N_7001);
and U7653 (N_7653,N_7102,N_7193);
nand U7654 (N_7654,N_7114,N_7380);
nor U7655 (N_7655,N_7088,N_7194);
or U7656 (N_7656,N_7317,N_7234);
xor U7657 (N_7657,N_7010,N_7334);
nor U7658 (N_7658,N_7243,N_7498);
nand U7659 (N_7659,N_7122,N_7103);
nor U7660 (N_7660,N_7207,N_7499);
nor U7661 (N_7661,N_7416,N_7185);
nand U7662 (N_7662,N_7124,N_7303);
or U7663 (N_7663,N_7187,N_7354);
nor U7664 (N_7664,N_7011,N_7246);
and U7665 (N_7665,N_7129,N_7469);
nand U7666 (N_7666,N_7139,N_7361);
nor U7667 (N_7667,N_7056,N_7387);
or U7668 (N_7668,N_7111,N_7177);
nor U7669 (N_7669,N_7391,N_7017);
and U7670 (N_7670,N_7344,N_7254);
and U7671 (N_7671,N_7031,N_7420);
nor U7672 (N_7672,N_7242,N_7232);
and U7673 (N_7673,N_7132,N_7033);
and U7674 (N_7674,N_7141,N_7327);
nor U7675 (N_7675,N_7415,N_7006);
and U7676 (N_7676,N_7191,N_7143);
or U7677 (N_7677,N_7030,N_7358);
or U7678 (N_7678,N_7333,N_7216);
nor U7679 (N_7679,N_7012,N_7059);
or U7680 (N_7680,N_7261,N_7196);
nand U7681 (N_7681,N_7130,N_7047);
nand U7682 (N_7682,N_7028,N_7155);
nor U7683 (N_7683,N_7251,N_7350);
nor U7684 (N_7684,N_7262,N_7470);
nor U7685 (N_7685,N_7169,N_7467);
nor U7686 (N_7686,N_7486,N_7240);
and U7687 (N_7687,N_7164,N_7482);
and U7688 (N_7688,N_7070,N_7009);
nand U7689 (N_7689,N_7446,N_7299);
nand U7690 (N_7690,N_7015,N_7411);
or U7691 (N_7691,N_7181,N_7292);
or U7692 (N_7692,N_7253,N_7112);
and U7693 (N_7693,N_7428,N_7276);
nor U7694 (N_7694,N_7140,N_7330);
nor U7695 (N_7695,N_7434,N_7163);
and U7696 (N_7696,N_7197,N_7093);
or U7697 (N_7697,N_7136,N_7092);
nand U7698 (N_7698,N_7402,N_7225);
and U7699 (N_7699,N_7208,N_7400);
nand U7700 (N_7700,N_7131,N_7223);
nor U7701 (N_7701,N_7343,N_7183);
or U7702 (N_7702,N_7417,N_7053);
and U7703 (N_7703,N_7144,N_7058);
nand U7704 (N_7704,N_7075,N_7260);
and U7705 (N_7705,N_7310,N_7436);
or U7706 (N_7706,N_7256,N_7077);
nand U7707 (N_7707,N_7013,N_7041);
xor U7708 (N_7708,N_7294,N_7025);
or U7709 (N_7709,N_7448,N_7268);
nand U7710 (N_7710,N_7379,N_7179);
nor U7711 (N_7711,N_7351,N_7452);
xnor U7712 (N_7712,N_7320,N_7213);
and U7713 (N_7713,N_7426,N_7335);
nand U7714 (N_7714,N_7355,N_7170);
or U7715 (N_7715,N_7171,N_7214);
xnor U7716 (N_7716,N_7071,N_7422);
nor U7717 (N_7717,N_7055,N_7060);
nand U7718 (N_7718,N_7176,N_7477);
nand U7719 (N_7719,N_7311,N_7184);
or U7720 (N_7720,N_7049,N_7076);
xnor U7721 (N_7721,N_7483,N_7222);
and U7722 (N_7722,N_7044,N_7279);
xor U7723 (N_7723,N_7073,N_7393);
nor U7724 (N_7724,N_7407,N_7421);
nand U7725 (N_7725,N_7306,N_7497);
nand U7726 (N_7726,N_7281,N_7241);
or U7727 (N_7727,N_7431,N_7396);
nor U7728 (N_7728,N_7449,N_7445);
or U7729 (N_7729,N_7039,N_7397);
or U7730 (N_7730,N_7118,N_7227);
nor U7731 (N_7731,N_7212,N_7035);
and U7732 (N_7732,N_7023,N_7273);
or U7733 (N_7733,N_7340,N_7002);
nand U7734 (N_7734,N_7230,N_7435);
nor U7735 (N_7735,N_7316,N_7206);
and U7736 (N_7736,N_7008,N_7078);
nand U7737 (N_7737,N_7357,N_7284);
or U7738 (N_7738,N_7083,N_7298);
nor U7739 (N_7739,N_7003,N_7127);
nor U7740 (N_7740,N_7014,N_7190);
and U7741 (N_7741,N_7374,N_7487);
nand U7742 (N_7742,N_7016,N_7405);
nand U7743 (N_7743,N_7291,N_7440);
nand U7744 (N_7744,N_7368,N_7383);
and U7745 (N_7745,N_7485,N_7026);
or U7746 (N_7746,N_7478,N_7395);
nand U7747 (N_7747,N_7366,N_7117);
nand U7748 (N_7748,N_7116,N_7043);
nor U7749 (N_7749,N_7280,N_7450);
nor U7750 (N_7750,N_7072,N_7013);
nand U7751 (N_7751,N_7378,N_7347);
nand U7752 (N_7752,N_7388,N_7333);
xnor U7753 (N_7753,N_7283,N_7275);
nor U7754 (N_7754,N_7464,N_7458);
nor U7755 (N_7755,N_7382,N_7082);
nor U7756 (N_7756,N_7168,N_7130);
and U7757 (N_7757,N_7077,N_7153);
nand U7758 (N_7758,N_7491,N_7191);
xor U7759 (N_7759,N_7199,N_7149);
nand U7760 (N_7760,N_7216,N_7278);
nor U7761 (N_7761,N_7223,N_7058);
nor U7762 (N_7762,N_7241,N_7215);
nor U7763 (N_7763,N_7378,N_7242);
and U7764 (N_7764,N_7482,N_7080);
nand U7765 (N_7765,N_7272,N_7296);
nor U7766 (N_7766,N_7127,N_7161);
nor U7767 (N_7767,N_7206,N_7395);
nor U7768 (N_7768,N_7238,N_7152);
or U7769 (N_7769,N_7491,N_7358);
nor U7770 (N_7770,N_7342,N_7417);
nor U7771 (N_7771,N_7075,N_7062);
nor U7772 (N_7772,N_7431,N_7311);
or U7773 (N_7773,N_7288,N_7219);
and U7774 (N_7774,N_7364,N_7066);
nand U7775 (N_7775,N_7332,N_7402);
or U7776 (N_7776,N_7025,N_7108);
or U7777 (N_7777,N_7104,N_7415);
nor U7778 (N_7778,N_7435,N_7033);
or U7779 (N_7779,N_7124,N_7101);
nor U7780 (N_7780,N_7372,N_7340);
or U7781 (N_7781,N_7489,N_7320);
nand U7782 (N_7782,N_7277,N_7121);
or U7783 (N_7783,N_7279,N_7408);
nand U7784 (N_7784,N_7467,N_7320);
xnor U7785 (N_7785,N_7332,N_7118);
nand U7786 (N_7786,N_7264,N_7060);
or U7787 (N_7787,N_7326,N_7483);
or U7788 (N_7788,N_7259,N_7491);
or U7789 (N_7789,N_7169,N_7293);
or U7790 (N_7790,N_7432,N_7463);
nor U7791 (N_7791,N_7441,N_7258);
and U7792 (N_7792,N_7227,N_7283);
nand U7793 (N_7793,N_7312,N_7221);
or U7794 (N_7794,N_7293,N_7323);
and U7795 (N_7795,N_7152,N_7268);
nor U7796 (N_7796,N_7223,N_7092);
nor U7797 (N_7797,N_7281,N_7104);
xor U7798 (N_7798,N_7239,N_7458);
or U7799 (N_7799,N_7393,N_7127);
or U7800 (N_7800,N_7006,N_7155);
and U7801 (N_7801,N_7352,N_7344);
nor U7802 (N_7802,N_7400,N_7385);
nand U7803 (N_7803,N_7325,N_7244);
nand U7804 (N_7804,N_7407,N_7147);
and U7805 (N_7805,N_7225,N_7461);
or U7806 (N_7806,N_7429,N_7367);
xor U7807 (N_7807,N_7320,N_7122);
xor U7808 (N_7808,N_7333,N_7320);
or U7809 (N_7809,N_7262,N_7146);
or U7810 (N_7810,N_7064,N_7335);
nor U7811 (N_7811,N_7008,N_7187);
nor U7812 (N_7812,N_7483,N_7452);
nand U7813 (N_7813,N_7063,N_7358);
nand U7814 (N_7814,N_7218,N_7221);
and U7815 (N_7815,N_7348,N_7211);
and U7816 (N_7816,N_7446,N_7236);
and U7817 (N_7817,N_7105,N_7297);
xor U7818 (N_7818,N_7020,N_7139);
and U7819 (N_7819,N_7256,N_7164);
and U7820 (N_7820,N_7374,N_7090);
and U7821 (N_7821,N_7306,N_7282);
xor U7822 (N_7822,N_7191,N_7407);
or U7823 (N_7823,N_7468,N_7082);
xnor U7824 (N_7824,N_7439,N_7153);
xnor U7825 (N_7825,N_7247,N_7193);
nand U7826 (N_7826,N_7289,N_7467);
or U7827 (N_7827,N_7449,N_7339);
xor U7828 (N_7828,N_7021,N_7417);
and U7829 (N_7829,N_7386,N_7107);
or U7830 (N_7830,N_7096,N_7165);
nor U7831 (N_7831,N_7301,N_7205);
xor U7832 (N_7832,N_7393,N_7241);
nand U7833 (N_7833,N_7012,N_7332);
or U7834 (N_7834,N_7136,N_7089);
or U7835 (N_7835,N_7443,N_7121);
nor U7836 (N_7836,N_7419,N_7349);
and U7837 (N_7837,N_7181,N_7467);
xnor U7838 (N_7838,N_7214,N_7318);
nand U7839 (N_7839,N_7081,N_7094);
and U7840 (N_7840,N_7297,N_7003);
nand U7841 (N_7841,N_7200,N_7244);
nor U7842 (N_7842,N_7453,N_7017);
and U7843 (N_7843,N_7186,N_7491);
nand U7844 (N_7844,N_7033,N_7248);
and U7845 (N_7845,N_7003,N_7047);
nor U7846 (N_7846,N_7065,N_7388);
and U7847 (N_7847,N_7348,N_7141);
and U7848 (N_7848,N_7340,N_7141);
nand U7849 (N_7849,N_7335,N_7429);
and U7850 (N_7850,N_7109,N_7164);
nor U7851 (N_7851,N_7334,N_7447);
xnor U7852 (N_7852,N_7117,N_7341);
xor U7853 (N_7853,N_7255,N_7141);
nand U7854 (N_7854,N_7067,N_7211);
nor U7855 (N_7855,N_7061,N_7424);
and U7856 (N_7856,N_7183,N_7118);
nand U7857 (N_7857,N_7012,N_7435);
and U7858 (N_7858,N_7172,N_7125);
or U7859 (N_7859,N_7141,N_7285);
xnor U7860 (N_7860,N_7209,N_7033);
nand U7861 (N_7861,N_7496,N_7071);
or U7862 (N_7862,N_7391,N_7243);
xor U7863 (N_7863,N_7458,N_7351);
and U7864 (N_7864,N_7487,N_7494);
nor U7865 (N_7865,N_7398,N_7162);
or U7866 (N_7866,N_7458,N_7317);
and U7867 (N_7867,N_7451,N_7329);
nor U7868 (N_7868,N_7331,N_7019);
nand U7869 (N_7869,N_7346,N_7017);
nand U7870 (N_7870,N_7189,N_7258);
or U7871 (N_7871,N_7179,N_7297);
and U7872 (N_7872,N_7061,N_7417);
xor U7873 (N_7873,N_7016,N_7346);
and U7874 (N_7874,N_7441,N_7084);
nor U7875 (N_7875,N_7318,N_7329);
and U7876 (N_7876,N_7393,N_7230);
and U7877 (N_7877,N_7207,N_7472);
or U7878 (N_7878,N_7378,N_7063);
nand U7879 (N_7879,N_7493,N_7406);
nor U7880 (N_7880,N_7368,N_7297);
or U7881 (N_7881,N_7076,N_7099);
nor U7882 (N_7882,N_7390,N_7089);
and U7883 (N_7883,N_7047,N_7198);
nor U7884 (N_7884,N_7382,N_7172);
and U7885 (N_7885,N_7329,N_7218);
or U7886 (N_7886,N_7307,N_7279);
nor U7887 (N_7887,N_7334,N_7481);
nand U7888 (N_7888,N_7294,N_7130);
or U7889 (N_7889,N_7029,N_7323);
and U7890 (N_7890,N_7095,N_7163);
nor U7891 (N_7891,N_7079,N_7094);
and U7892 (N_7892,N_7234,N_7111);
or U7893 (N_7893,N_7022,N_7124);
nand U7894 (N_7894,N_7107,N_7267);
or U7895 (N_7895,N_7373,N_7173);
nand U7896 (N_7896,N_7093,N_7277);
nand U7897 (N_7897,N_7096,N_7136);
nor U7898 (N_7898,N_7147,N_7393);
nand U7899 (N_7899,N_7275,N_7405);
nand U7900 (N_7900,N_7442,N_7069);
and U7901 (N_7901,N_7268,N_7312);
and U7902 (N_7902,N_7109,N_7328);
and U7903 (N_7903,N_7347,N_7050);
or U7904 (N_7904,N_7470,N_7236);
nor U7905 (N_7905,N_7179,N_7491);
nor U7906 (N_7906,N_7009,N_7160);
and U7907 (N_7907,N_7340,N_7251);
nor U7908 (N_7908,N_7256,N_7225);
nor U7909 (N_7909,N_7081,N_7238);
xor U7910 (N_7910,N_7143,N_7209);
nand U7911 (N_7911,N_7451,N_7453);
nor U7912 (N_7912,N_7437,N_7219);
or U7913 (N_7913,N_7311,N_7357);
nor U7914 (N_7914,N_7165,N_7394);
xor U7915 (N_7915,N_7068,N_7149);
nor U7916 (N_7916,N_7032,N_7360);
nand U7917 (N_7917,N_7486,N_7316);
nor U7918 (N_7918,N_7455,N_7402);
nor U7919 (N_7919,N_7327,N_7013);
or U7920 (N_7920,N_7440,N_7344);
or U7921 (N_7921,N_7006,N_7079);
nand U7922 (N_7922,N_7233,N_7087);
and U7923 (N_7923,N_7369,N_7105);
and U7924 (N_7924,N_7094,N_7060);
nand U7925 (N_7925,N_7038,N_7348);
nor U7926 (N_7926,N_7254,N_7071);
nor U7927 (N_7927,N_7201,N_7377);
nor U7928 (N_7928,N_7464,N_7359);
nor U7929 (N_7929,N_7459,N_7006);
nand U7930 (N_7930,N_7275,N_7471);
nand U7931 (N_7931,N_7382,N_7416);
nor U7932 (N_7932,N_7415,N_7280);
nand U7933 (N_7933,N_7037,N_7363);
nor U7934 (N_7934,N_7320,N_7137);
nor U7935 (N_7935,N_7120,N_7060);
or U7936 (N_7936,N_7083,N_7093);
nand U7937 (N_7937,N_7177,N_7268);
or U7938 (N_7938,N_7420,N_7098);
nand U7939 (N_7939,N_7013,N_7246);
and U7940 (N_7940,N_7280,N_7310);
nor U7941 (N_7941,N_7398,N_7325);
nor U7942 (N_7942,N_7238,N_7283);
nand U7943 (N_7943,N_7195,N_7193);
nand U7944 (N_7944,N_7269,N_7125);
or U7945 (N_7945,N_7045,N_7362);
nand U7946 (N_7946,N_7141,N_7428);
nor U7947 (N_7947,N_7384,N_7382);
nor U7948 (N_7948,N_7097,N_7010);
and U7949 (N_7949,N_7317,N_7161);
and U7950 (N_7950,N_7299,N_7144);
or U7951 (N_7951,N_7195,N_7019);
nor U7952 (N_7952,N_7164,N_7111);
nor U7953 (N_7953,N_7392,N_7461);
or U7954 (N_7954,N_7195,N_7054);
nand U7955 (N_7955,N_7093,N_7304);
nor U7956 (N_7956,N_7396,N_7344);
or U7957 (N_7957,N_7174,N_7014);
and U7958 (N_7958,N_7095,N_7459);
nor U7959 (N_7959,N_7196,N_7304);
nand U7960 (N_7960,N_7179,N_7004);
nor U7961 (N_7961,N_7159,N_7350);
and U7962 (N_7962,N_7355,N_7239);
or U7963 (N_7963,N_7238,N_7389);
or U7964 (N_7964,N_7119,N_7014);
and U7965 (N_7965,N_7282,N_7303);
nor U7966 (N_7966,N_7158,N_7073);
or U7967 (N_7967,N_7272,N_7404);
or U7968 (N_7968,N_7069,N_7119);
nor U7969 (N_7969,N_7325,N_7205);
and U7970 (N_7970,N_7339,N_7245);
and U7971 (N_7971,N_7337,N_7055);
or U7972 (N_7972,N_7381,N_7307);
xnor U7973 (N_7973,N_7420,N_7282);
or U7974 (N_7974,N_7161,N_7329);
nor U7975 (N_7975,N_7067,N_7386);
or U7976 (N_7976,N_7245,N_7273);
or U7977 (N_7977,N_7330,N_7359);
or U7978 (N_7978,N_7095,N_7061);
and U7979 (N_7979,N_7388,N_7384);
or U7980 (N_7980,N_7270,N_7373);
nand U7981 (N_7981,N_7119,N_7370);
and U7982 (N_7982,N_7041,N_7309);
and U7983 (N_7983,N_7130,N_7190);
and U7984 (N_7984,N_7131,N_7483);
nand U7985 (N_7985,N_7188,N_7273);
or U7986 (N_7986,N_7315,N_7456);
or U7987 (N_7987,N_7151,N_7139);
or U7988 (N_7988,N_7412,N_7067);
and U7989 (N_7989,N_7329,N_7242);
nor U7990 (N_7990,N_7419,N_7401);
or U7991 (N_7991,N_7291,N_7397);
nor U7992 (N_7992,N_7122,N_7330);
or U7993 (N_7993,N_7300,N_7475);
and U7994 (N_7994,N_7197,N_7212);
nor U7995 (N_7995,N_7218,N_7048);
nor U7996 (N_7996,N_7158,N_7178);
or U7997 (N_7997,N_7218,N_7033);
nand U7998 (N_7998,N_7213,N_7322);
or U7999 (N_7999,N_7252,N_7098);
and U8000 (N_8000,N_7996,N_7890);
or U8001 (N_8001,N_7663,N_7694);
nor U8002 (N_8002,N_7844,N_7531);
or U8003 (N_8003,N_7911,N_7571);
xnor U8004 (N_8004,N_7500,N_7568);
and U8005 (N_8005,N_7842,N_7725);
and U8006 (N_8006,N_7575,N_7516);
nand U8007 (N_8007,N_7888,N_7748);
or U8008 (N_8008,N_7608,N_7562);
nor U8009 (N_8009,N_7808,N_7975);
nor U8010 (N_8010,N_7533,N_7772);
xnor U8011 (N_8011,N_7632,N_7811);
or U8012 (N_8012,N_7731,N_7992);
nor U8013 (N_8013,N_7509,N_7827);
or U8014 (N_8014,N_7920,N_7918);
xor U8015 (N_8015,N_7603,N_7615);
or U8016 (N_8016,N_7702,N_7995);
nand U8017 (N_8017,N_7733,N_7578);
nand U8018 (N_8018,N_7592,N_7651);
and U8019 (N_8019,N_7938,N_7609);
nand U8020 (N_8020,N_7803,N_7939);
or U8021 (N_8021,N_7602,N_7908);
or U8022 (N_8022,N_7832,N_7659);
and U8023 (N_8023,N_7830,N_7940);
or U8024 (N_8024,N_7793,N_7744);
and U8025 (N_8025,N_7794,N_7859);
and U8026 (N_8026,N_7840,N_7504);
or U8027 (N_8027,N_7595,N_7957);
nand U8028 (N_8028,N_7955,N_7836);
and U8029 (N_8029,N_7580,N_7942);
nand U8030 (N_8030,N_7916,N_7593);
and U8031 (N_8031,N_7998,N_7610);
and U8032 (N_8032,N_7936,N_7770);
and U8033 (N_8033,N_7515,N_7687);
or U8034 (N_8034,N_7706,N_7508);
nor U8035 (N_8035,N_7849,N_7950);
and U8036 (N_8036,N_7743,N_7929);
nand U8037 (N_8037,N_7660,N_7596);
nand U8038 (N_8038,N_7644,N_7814);
nand U8039 (N_8039,N_7894,N_7551);
xor U8040 (N_8040,N_7789,N_7530);
or U8041 (N_8041,N_7764,N_7582);
or U8042 (N_8042,N_7798,N_7638);
or U8043 (N_8043,N_7716,N_7829);
and U8044 (N_8044,N_7962,N_7505);
and U8045 (N_8045,N_7944,N_7542);
and U8046 (N_8046,N_7721,N_7870);
and U8047 (N_8047,N_7834,N_7787);
nor U8048 (N_8048,N_7761,N_7853);
nand U8049 (N_8049,N_7757,N_7540);
nand U8050 (N_8050,N_7915,N_7614);
and U8051 (N_8051,N_7857,N_7963);
and U8052 (N_8052,N_7564,N_7601);
and U8053 (N_8053,N_7873,N_7735);
and U8054 (N_8054,N_7750,N_7521);
and U8055 (N_8055,N_7848,N_7876);
xnor U8056 (N_8056,N_7503,N_7692);
nor U8057 (N_8057,N_7906,N_7833);
nand U8058 (N_8058,N_7538,N_7847);
or U8059 (N_8059,N_7774,N_7947);
xor U8060 (N_8060,N_7980,N_7785);
or U8061 (N_8061,N_7924,N_7636);
or U8062 (N_8062,N_7835,N_7741);
and U8063 (N_8063,N_7749,N_7524);
nor U8064 (N_8064,N_7545,N_7559);
or U8065 (N_8065,N_7522,N_7755);
nand U8066 (N_8066,N_7856,N_7710);
nand U8067 (N_8067,N_7552,N_7622);
xor U8068 (N_8068,N_7588,N_7628);
nand U8069 (N_8069,N_7776,N_7838);
and U8070 (N_8070,N_7543,N_7520);
nand U8071 (N_8071,N_7556,N_7747);
nand U8072 (N_8072,N_7783,N_7535);
or U8073 (N_8073,N_7819,N_7567);
nand U8074 (N_8074,N_7788,N_7907);
and U8075 (N_8075,N_7587,N_7801);
or U8076 (N_8076,N_7901,N_7573);
and U8077 (N_8077,N_7983,N_7989);
nor U8078 (N_8078,N_7821,N_7717);
or U8079 (N_8079,N_7802,N_7946);
nand U8080 (N_8080,N_7700,N_7926);
xnor U8081 (N_8081,N_7919,N_7815);
nor U8082 (N_8082,N_7745,N_7536);
and U8083 (N_8083,N_7661,N_7928);
or U8084 (N_8084,N_7896,N_7686);
or U8085 (N_8085,N_7809,N_7646);
nor U8086 (N_8086,N_7952,N_7537);
or U8087 (N_8087,N_7519,N_7976);
and U8088 (N_8088,N_7855,N_7669);
nor U8089 (N_8089,N_7810,N_7956);
or U8090 (N_8090,N_7937,N_7675);
xnor U8091 (N_8091,N_7642,N_7941);
or U8092 (N_8092,N_7795,N_7804);
nand U8093 (N_8093,N_7607,N_7641);
xnor U8094 (N_8094,N_7704,N_7781);
nand U8095 (N_8095,N_7865,N_7586);
and U8096 (N_8096,N_7779,N_7875);
nor U8097 (N_8097,N_7862,N_7698);
nor U8098 (N_8098,N_7553,N_7742);
nand U8099 (N_8099,N_7726,N_7597);
or U8100 (N_8100,N_7913,N_7985);
xnor U8101 (N_8101,N_7673,N_7711);
or U8102 (N_8102,N_7885,N_7752);
nor U8103 (N_8103,N_7886,N_7969);
nor U8104 (N_8104,N_7696,N_7867);
nor U8105 (N_8105,N_7910,N_7773);
xnor U8106 (N_8106,N_7541,N_7624);
nand U8107 (N_8107,N_7997,N_7887);
nor U8108 (N_8108,N_7643,N_7902);
nor U8109 (N_8109,N_7714,N_7767);
nor U8110 (N_8110,N_7884,N_7507);
or U8111 (N_8111,N_7900,N_7999);
nand U8112 (N_8112,N_7868,N_7713);
and U8113 (N_8113,N_7612,N_7548);
and U8114 (N_8114,N_7839,N_7786);
nand U8115 (N_8115,N_7668,N_7925);
nand U8116 (N_8116,N_7554,N_7576);
and U8117 (N_8117,N_7816,N_7662);
nor U8118 (N_8118,N_7699,N_7558);
nand U8119 (N_8119,N_7871,N_7778);
or U8120 (N_8120,N_7591,N_7861);
and U8121 (N_8121,N_7828,N_7968);
nand U8122 (N_8122,N_7639,N_7528);
nand U8123 (N_8123,N_7506,N_7674);
xor U8124 (N_8124,N_7927,N_7967);
nor U8125 (N_8125,N_7518,N_7645);
nor U8126 (N_8126,N_7800,N_7818);
nor U8127 (N_8127,N_7600,N_7513);
or U8128 (N_8128,N_7824,N_7729);
and U8129 (N_8129,N_7945,N_7780);
nand U8130 (N_8130,N_7703,N_7977);
nand U8131 (N_8131,N_7647,N_7799);
and U8132 (N_8132,N_7547,N_7715);
nand U8133 (N_8133,N_7790,N_7720);
nor U8134 (N_8134,N_7617,N_7739);
nand U8135 (N_8135,N_7549,N_7579);
nand U8136 (N_8136,N_7690,N_7917);
nor U8137 (N_8137,N_7878,N_7589);
nor U8138 (N_8138,N_7680,N_7990);
or U8139 (N_8139,N_7685,N_7740);
nor U8140 (N_8140,N_7931,N_7572);
nor U8141 (N_8141,N_7759,N_7991);
nand U8142 (N_8142,N_7718,N_7972);
and U8143 (N_8143,N_7532,N_7523);
and U8144 (N_8144,N_7762,N_7891);
or U8145 (N_8145,N_7681,N_7728);
or U8146 (N_8146,N_7550,N_7649);
nand U8147 (N_8147,N_7866,N_7973);
or U8148 (N_8148,N_7514,N_7760);
nor U8149 (N_8149,N_7914,N_7805);
and U8150 (N_8150,N_7820,N_7796);
or U8151 (N_8151,N_7574,N_7974);
or U8152 (N_8152,N_7852,N_7619);
and U8153 (N_8153,N_7623,N_7934);
or U8154 (N_8154,N_7701,N_7527);
nor U8155 (N_8155,N_7670,N_7650);
and U8156 (N_8156,N_7843,N_7544);
or U8157 (N_8157,N_7583,N_7654);
nand U8158 (N_8158,N_7510,N_7889);
or U8159 (N_8159,N_7604,N_7961);
nand U8160 (N_8160,N_7869,N_7598);
xnor U8161 (N_8161,N_7970,N_7791);
or U8162 (N_8162,N_7708,N_7664);
and U8163 (N_8163,N_7775,N_7905);
nor U8164 (N_8164,N_7666,N_7611);
and U8165 (N_8165,N_7893,N_7812);
and U8166 (N_8166,N_7882,N_7599);
nand U8167 (N_8167,N_7695,N_7813);
or U8168 (N_8168,N_7935,N_7979);
nor U8169 (N_8169,N_7984,N_7502);
nor U8170 (N_8170,N_7863,N_7954);
or U8171 (N_8171,N_7620,N_7566);
or U8172 (N_8172,N_7782,N_7883);
or U8173 (N_8173,N_7555,N_7529);
nand U8174 (N_8174,N_7897,N_7831);
or U8175 (N_8175,N_7658,N_7964);
or U8176 (N_8176,N_7546,N_7960);
nand U8177 (N_8177,N_7948,N_7858);
nand U8178 (N_8178,N_7797,N_7943);
and U8179 (N_8179,N_7570,N_7584);
nor U8180 (N_8180,N_7665,N_7763);
nand U8181 (N_8181,N_7903,N_7605);
or U8182 (N_8182,N_7629,N_7616);
nand U8183 (N_8183,N_7724,N_7678);
nor U8184 (N_8184,N_7874,N_7734);
nor U8185 (N_8185,N_7994,N_7705);
and U8186 (N_8186,N_7534,N_7656);
and U8187 (N_8187,N_7892,N_7765);
and U8188 (N_8188,N_7951,N_7727);
or U8189 (N_8189,N_7958,N_7971);
nand U8190 (N_8190,N_7618,N_7606);
nand U8191 (N_8191,N_7630,N_7933);
nand U8192 (N_8192,N_7648,N_7879);
nor U8193 (N_8193,N_7806,N_7634);
nor U8194 (N_8194,N_7525,N_7921);
nor U8195 (N_8195,N_7557,N_7754);
and U8196 (N_8196,N_7904,N_7930);
and U8197 (N_8197,N_7766,N_7707);
nor U8198 (N_8198,N_7563,N_7684);
and U8199 (N_8199,N_7526,N_7657);
or U8200 (N_8200,N_7982,N_7736);
nand U8201 (N_8201,N_7966,N_7625);
nor U8202 (N_8202,N_7923,N_7898);
and U8203 (N_8203,N_7652,N_7682);
or U8204 (N_8204,N_7689,N_7993);
and U8205 (N_8205,N_7826,N_7746);
nor U8206 (N_8206,N_7922,N_7693);
or U8207 (N_8207,N_7565,N_7845);
nand U8208 (N_8208,N_7807,N_7577);
and U8209 (N_8209,N_7841,N_7676);
and U8210 (N_8210,N_7758,N_7895);
nand U8211 (N_8211,N_7719,N_7688);
or U8212 (N_8212,N_7512,N_7899);
nor U8213 (N_8213,N_7932,N_7986);
nand U8214 (N_8214,N_7511,N_7881);
and U8215 (N_8215,N_7822,N_7581);
and U8216 (N_8216,N_7539,N_7959);
and U8217 (N_8217,N_7709,N_7640);
xnor U8218 (N_8218,N_7594,N_7825);
nor U8219 (N_8219,N_7769,N_7756);
and U8220 (N_8220,N_7965,N_7712);
nand U8221 (N_8221,N_7880,N_7621);
or U8222 (N_8222,N_7730,N_7633);
nand U8223 (N_8223,N_7988,N_7851);
and U8224 (N_8224,N_7501,N_7846);
or U8225 (N_8225,N_7569,N_7912);
nor U8226 (N_8226,N_7854,N_7722);
nand U8227 (N_8227,N_7909,N_7823);
nand U8228 (N_8228,N_7683,N_7768);
nand U8229 (N_8229,N_7872,N_7561);
nand U8230 (N_8230,N_7723,N_7751);
nor U8231 (N_8231,N_7672,N_7978);
and U8232 (N_8232,N_7627,N_7817);
and U8233 (N_8233,N_7585,N_7635);
nor U8234 (N_8234,N_7691,N_7667);
xor U8235 (N_8235,N_7784,N_7949);
nor U8236 (N_8236,N_7953,N_7837);
nand U8237 (N_8237,N_7753,N_7677);
and U8238 (N_8238,N_7860,N_7737);
nand U8239 (N_8239,N_7792,N_7864);
nand U8240 (N_8240,N_7626,N_7877);
nand U8241 (N_8241,N_7613,N_7771);
or U8242 (N_8242,N_7631,N_7777);
xor U8243 (N_8243,N_7981,N_7590);
and U8244 (N_8244,N_7560,N_7679);
xnor U8245 (N_8245,N_7637,N_7987);
and U8246 (N_8246,N_7738,N_7671);
and U8247 (N_8247,N_7850,N_7517);
nor U8248 (N_8248,N_7655,N_7697);
xnor U8249 (N_8249,N_7653,N_7732);
and U8250 (N_8250,N_7838,N_7941);
nand U8251 (N_8251,N_7544,N_7948);
and U8252 (N_8252,N_7898,N_7973);
and U8253 (N_8253,N_7985,N_7931);
and U8254 (N_8254,N_7966,N_7793);
and U8255 (N_8255,N_7937,N_7534);
or U8256 (N_8256,N_7861,N_7763);
nor U8257 (N_8257,N_7892,N_7931);
or U8258 (N_8258,N_7763,N_7647);
nor U8259 (N_8259,N_7956,N_7925);
nor U8260 (N_8260,N_7507,N_7618);
and U8261 (N_8261,N_7679,N_7885);
and U8262 (N_8262,N_7540,N_7755);
xnor U8263 (N_8263,N_7569,N_7968);
or U8264 (N_8264,N_7859,N_7988);
xnor U8265 (N_8265,N_7710,N_7862);
xnor U8266 (N_8266,N_7825,N_7707);
nand U8267 (N_8267,N_7650,N_7869);
nor U8268 (N_8268,N_7724,N_7526);
nor U8269 (N_8269,N_7792,N_7962);
and U8270 (N_8270,N_7754,N_7999);
nor U8271 (N_8271,N_7727,N_7512);
nor U8272 (N_8272,N_7552,N_7584);
or U8273 (N_8273,N_7551,N_7956);
and U8274 (N_8274,N_7554,N_7716);
nor U8275 (N_8275,N_7774,N_7866);
and U8276 (N_8276,N_7573,N_7649);
or U8277 (N_8277,N_7937,N_7697);
nand U8278 (N_8278,N_7807,N_7536);
or U8279 (N_8279,N_7987,N_7902);
nand U8280 (N_8280,N_7848,N_7958);
nand U8281 (N_8281,N_7652,N_7813);
xor U8282 (N_8282,N_7684,N_7828);
nand U8283 (N_8283,N_7628,N_7637);
nor U8284 (N_8284,N_7811,N_7578);
nor U8285 (N_8285,N_7742,N_7758);
and U8286 (N_8286,N_7944,N_7707);
nand U8287 (N_8287,N_7693,N_7977);
and U8288 (N_8288,N_7823,N_7544);
or U8289 (N_8289,N_7889,N_7789);
and U8290 (N_8290,N_7991,N_7987);
or U8291 (N_8291,N_7536,N_7865);
nor U8292 (N_8292,N_7871,N_7500);
and U8293 (N_8293,N_7711,N_7693);
nand U8294 (N_8294,N_7505,N_7524);
and U8295 (N_8295,N_7862,N_7843);
and U8296 (N_8296,N_7552,N_7508);
nor U8297 (N_8297,N_7819,N_7980);
nor U8298 (N_8298,N_7919,N_7857);
nor U8299 (N_8299,N_7904,N_7554);
and U8300 (N_8300,N_7607,N_7848);
and U8301 (N_8301,N_7978,N_7856);
and U8302 (N_8302,N_7621,N_7568);
or U8303 (N_8303,N_7666,N_7711);
nor U8304 (N_8304,N_7991,N_7766);
xnor U8305 (N_8305,N_7626,N_7521);
or U8306 (N_8306,N_7872,N_7507);
or U8307 (N_8307,N_7576,N_7708);
and U8308 (N_8308,N_7784,N_7977);
or U8309 (N_8309,N_7593,N_7923);
xnor U8310 (N_8310,N_7995,N_7537);
nor U8311 (N_8311,N_7679,N_7810);
and U8312 (N_8312,N_7657,N_7522);
nand U8313 (N_8313,N_7739,N_7870);
nand U8314 (N_8314,N_7586,N_7779);
nand U8315 (N_8315,N_7599,N_7818);
nor U8316 (N_8316,N_7776,N_7976);
and U8317 (N_8317,N_7748,N_7924);
nand U8318 (N_8318,N_7508,N_7801);
nor U8319 (N_8319,N_7831,N_7787);
nor U8320 (N_8320,N_7805,N_7862);
or U8321 (N_8321,N_7586,N_7717);
or U8322 (N_8322,N_7946,N_7731);
nor U8323 (N_8323,N_7784,N_7571);
and U8324 (N_8324,N_7588,N_7576);
nor U8325 (N_8325,N_7972,N_7544);
nor U8326 (N_8326,N_7796,N_7696);
nor U8327 (N_8327,N_7849,N_7842);
or U8328 (N_8328,N_7965,N_7720);
or U8329 (N_8329,N_7962,N_7860);
or U8330 (N_8330,N_7650,N_7757);
or U8331 (N_8331,N_7716,N_7595);
nor U8332 (N_8332,N_7759,N_7881);
and U8333 (N_8333,N_7674,N_7798);
xnor U8334 (N_8334,N_7513,N_7626);
and U8335 (N_8335,N_7908,N_7851);
and U8336 (N_8336,N_7931,N_7787);
and U8337 (N_8337,N_7606,N_7679);
xor U8338 (N_8338,N_7610,N_7824);
or U8339 (N_8339,N_7622,N_7899);
nor U8340 (N_8340,N_7743,N_7761);
and U8341 (N_8341,N_7565,N_7857);
and U8342 (N_8342,N_7760,N_7578);
nor U8343 (N_8343,N_7957,N_7616);
xor U8344 (N_8344,N_7754,N_7763);
or U8345 (N_8345,N_7830,N_7989);
or U8346 (N_8346,N_7861,N_7764);
nand U8347 (N_8347,N_7660,N_7765);
or U8348 (N_8348,N_7537,N_7957);
nor U8349 (N_8349,N_7575,N_7991);
and U8350 (N_8350,N_7829,N_7853);
and U8351 (N_8351,N_7738,N_7896);
nand U8352 (N_8352,N_7711,N_7922);
and U8353 (N_8353,N_7947,N_7642);
nor U8354 (N_8354,N_7611,N_7798);
nor U8355 (N_8355,N_7887,N_7697);
nor U8356 (N_8356,N_7585,N_7997);
or U8357 (N_8357,N_7522,N_7574);
nand U8358 (N_8358,N_7938,N_7902);
nor U8359 (N_8359,N_7819,N_7841);
and U8360 (N_8360,N_7695,N_7830);
and U8361 (N_8361,N_7860,N_7784);
or U8362 (N_8362,N_7882,N_7843);
nand U8363 (N_8363,N_7792,N_7806);
nor U8364 (N_8364,N_7955,N_7676);
or U8365 (N_8365,N_7704,N_7690);
nand U8366 (N_8366,N_7860,N_7652);
nand U8367 (N_8367,N_7902,N_7701);
nor U8368 (N_8368,N_7912,N_7710);
nor U8369 (N_8369,N_7590,N_7664);
or U8370 (N_8370,N_7783,N_7860);
and U8371 (N_8371,N_7667,N_7826);
or U8372 (N_8372,N_7950,N_7635);
nand U8373 (N_8373,N_7694,N_7878);
nor U8374 (N_8374,N_7518,N_7799);
nor U8375 (N_8375,N_7640,N_7694);
nand U8376 (N_8376,N_7669,N_7973);
nand U8377 (N_8377,N_7859,N_7684);
xor U8378 (N_8378,N_7541,N_7693);
or U8379 (N_8379,N_7984,N_7939);
or U8380 (N_8380,N_7933,N_7826);
or U8381 (N_8381,N_7550,N_7987);
nand U8382 (N_8382,N_7753,N_7595);
nor U8383 (N_8383,N_7814,N_7784);
nor U8384 (N_8384,N_7563,N_7727);
and U8385 (N_8385,N_7971,N_7584);
or U8386 (N_8386,N_7923,N_7609);
and U8387 (N_8387,N_7681,N_7538);
and U8388 (N_8388,N_7735,N_7531);
nand U8389 (N_8389,N_7625,N_7763);
xor U8390 (N_8390,N_7554,N_7641);
and U8391 (N_8391,N_7723,N_7688);
and U8392 (N_8392,N_7731,N_7513);
and U8393 (N_8393,N_7577,N_7837);
nor U8394 (N_8394,N_7695,N_7588);
nor U8395 (N_8395,N_7745,N_7518);
and U8396 (N_8396,N_7551,N_7955);
or U8397 (N_8397,N_7940,N_7867);
nor U8398 (N_8398,N_7567,N_7612);
and U8399 (N_8399,N_7994,N_7876);
or U8400 (N_8400,N_7622,N_7681);
nor U8401 (N_8401,N_7831,N_7812);
nor U8402 (N_8402,N_7879,N_7696);
or U8403 (N_8403,N_7661,N_7778);
xor U8404 (N_8404,N_7958,N_7754);
or U8405 (N_8405,N_7597,N_7709);
xnor U8406 (N_8406,N_7758,N_7872);
nor U8407 (N_8407,N_7602,N_7860);
or U8408 (N_8408,N_7820,N_7883);
or U8409 (N_8409,N_7909,N_7858);
and U8410 (N_8410,N_7824,N_7599);
nor U8411 (N_8411,N_7706,N_7795);
and U8412 (N_8412,N_7700,N_7805);
and U8413 (N_8413,N_7808,N_7663);
xor U8414 (N_8414,N_7968,N_7705);
nand U8415 (N_8415,N_7668,N_7805);
or U8416 (N_8416,N_7983,N_7809);
and U8417 (N_8417,N_7872,N_7769);
and U8418 (N_8418,N_7870,N_7714);
nand U8419 (N_8419,N_7658,N_7506);
nand U8420 (N_8420,N_7798,N_7788);
and U8421 (N_8421,N_7625,N_7893);
xor U8422 (N_8422,N_7728,N_7743);
nand U8423 (N_8423,N_7695,N_7671);
nand U8424 (N_8424,N_7749,N_7555);
or U8425 (N_8425,N_7874,N_7660);
and U8426 (N_8426,N_7518,N_7713);
nand U8427 (N_8427,N_7607,N_7835);
nor U8428 (N_8428,N_7798,N_7992);
and U8429 (N_8429,N_7954,N_7836);
nor U8430 (N_8430,N_7965,N_7683);
nor U8431 (N_8431,N_7881,N_7858);
or U8432 (N_8432,N_7748,N_7820);
nor U8433 (N_8433,N_7738,N_7535);
nand U8434 (N_8434,N_7882,N_7938);
and U8435 (N_8435,N_7607,N_7558);
nor U8436 (N_8436,N_7762,N_7707);
xnor U8437 (N_8437,N_7500,N_7590);
nor U8438 (N_8438,N_7723,N_7912);
or U8439 (N_8439,N_7809,N_7938);
nand U8440 (N_8440,N_7672,N_7640);
and U8441 (N_8441,N_7800,N_7736);
or U8442 (N_8442,N_7567,N_7827);
and U8443 (N_8443,N_7820,N_7500);
nand U8444 (N_8444,N_7678,N_7952);
and U8445 (N_8445,N_7520,N_7878);
nor U8446 (N_8446,N_7839,N_7954);
or U8447 (N_8447,N_7921,N_7632);
nand U8448 (N_8448,N_7715,N_7925);
or U8449 (N_8449,N_7692,N_7518);
and U8450 (N_8450,N_7841,N_7901);
nand U8451 (N_8451,N_7722,N_7718);
and U8452 (N_8452,N_7706,N_7719);
nor U8453 (N_8453,N_7707,N_7872);
nor U8454 (N_8454,N_7670,N_7890);
nor U8455 (N_8455,N_7926,N_7551);
nand U8456 (N_8456,N_7912,N_7589);
nand U8457 (N_8457,N_7908,N_7682);
and U8458 (N_8458,N_7526,N_7557);
or U8459 (N_8459,N_7710,N_7605);
nor U8460 (N_8460,N_7807,N_7760);
nand U8461 (N_8461,N_7920,N_7619);
or U8462 (N_8462,N_7694,N_7760);
and U8463 (N_8463,N_7746,N_7778);
and U8464 (N_8464,N_7683,N_7622);
and U8465 (N_8465,N_7699,N_7513);
nor U8466 (N_8466,N_7894,N_7898);
or U8467 (N_8467,N_7868,N_7933);
and U8468 (N_8468,N_7976,N_7832);
and U8469 (N_8469,N_7865,N_7951);
or U8470 (N_8470,N_7946,N_7527);
and U8471 (N_8471,N_7764,N_7824);
and U8472 (N_8472,N_7882,N_7557);
nand U8473 (N_8473,N_7509,N_7626);
nand U8474 (N_8474,N_7500,N_7508);
xor U8475 (N_8475,N_7967,N_7531);
and U8476 (N_8476,N_7617,N_7750);
nand U8477 (N_8477,N_7596,N_7761);
or U8478 (N_8478,N_7613,N_7804);
nand U8479 (N_8479,N_7915,N_7896);
nand U8480 (N_8480,N_7952,N_7879);
or U8481 (N_8481,N_7875,N_7686);
or U8482 (N_8482,N_7661,N_7625);
and U8483 (N_8483,N_7743,N_7547);
xor U8484 (N_8484,N_7720,N_7964);
nor U8485 (N_8485,N_7621,N_7895);
nand U8486 (N_8486,N_7689,N_7592);
and U8487 (N_8487,N_7742,N_7646);
or U8488 (N_8488,N_7646,N_7840);
nor U8489 (N_8489,N_7565,N_7897);
nand U8490 (N_8490,N_7910,N_7814);
nor U8491 (N_8491,N_7921,N_7537);
and U8492 (N_8492,N_7803,N_7708);
or U8493 (N_8493,N_7670,N_7630);
nand U8494 (N_8494,N_7947,N_7538);
nand U8495 (N_8495,N_7859,N_7602);
or U8496 (N_8496,N_7891,N_7952);
and U8497 (N_8497,N_7780,N_7751);
and U8498 (N_8498,N_7948,N_7724);
nor U8499 (N_8499,N_7536,N_7631);
and U8500 (N_8500,N_8140,N_8168);
nand U8501 (N_8501,N_8110,N_8309);
nor U8502 (N_8502,N_8291,N_8256);
nand U8503 (N_8503,N_8451,N_8234);
or U8504 (N_8504,N_8406,N_8263);
or U8505 (N_8505,N_8359,N_8172);
nand U8506 (N_8506,N_8376,N_8498);
xnor U8507 (N_8507,N_8408,N_8214);
and U8508 (N_8508,N_8466,N_8308);
nand U8509 (N_8509,N_8370,N_8272);
nor U8510 (N_8510,N_8051,N_8289);
xor U8511 (N_8511,N_8392,N_8383);
and U8512 (N_8512,N_8008,N_8193);
nand U8513 (N_8513,N_8107,N_8056);
xnor U8514 (N_8514,N_8038,N_8298);
and U8515 (N_8515,N_8039,N_8029);
nor U8516 (N_8516,N_8266,N_8135);
xor U8517 (N_8517,N_8278,N_8178);
nor U8518 (N_8518,N_8350,N_8271);
and U8519 (N_8519,N_8077,N_8037);
xnor U8520 (N_8520,N_8373,N_8182);
or U8521 (N_8521,N_8415,N_8199);
or U8522 (N_8522,N_8353,N_8099);
xnor U8523 (N_8523,N_8185,N_8058);
nand U8524 (N_8524,N_8134,N_8343);
and U8525 (N_8525,N_8057,N_8103);
and U8526 (N_8526,N_8225,N_8102);
or U8527 (N_8527,N_8043,N_8418);
or U8528 (N_8528,N_8338,N_8106);
nand U8529 (N_8529,N_8410,N_8484);
nand U8530 (N_8530,N_8402,N_8421);
nand U8531 (N_8531,N_8048,N_8211);
nor U8532 (N_8532,N_8189,N_8206);
nand U8533 (N_8533,N_8380,N_8221);
or U8534 (N_8534,N_8310,N_8082);
nand U8535 (N_8535,N_8344,N_8327);
and U8536 (N_8536,N_8335,N_8479);
or U8537 (N_8537,N_8249,N_8478);
nand U8538 (N_8538,N_8012,N_8473);
and U8539 (N_8539,N_8024,N_8307);
nand U8540 (N_8540,N_8329,N_8313);
nand U8541 (N_8541,N_8210,N_8427);
and U8542 (N_8542,N_8398,N_8425);
and U8543 (N_8543,N_8433,N_8363);
nand U8544 (N_8544,N_8145,N_8397);
xor U8545 (N_8545,N_8286,N_8217);
and U8546 (N_8546,N_8460,N_8367);
nor U8547 (N_8547,N_8157,N_8318);
nor U8548 (N_8548,N_8416,N_8246);
nand U8549 (N_8549,N_8378,N_8042);
nor U8550 (N_8550,N_8238,N_8116);
nand U8551 (N_8551,N_8455,N_8068);
nor U8552 (N_8552,N_8482,N_8274);
nand U8553 (N_8553,N_8002,N_8026);
and U8554 (N_8554,N_8288,N_8203);
and U8555 (N_8555,N_8414,N_8073);
nand U8556 (N_8556,N_8314,N_8323);
nor U8557 (N_8557,N_8215,N_8171);
nor U8558 (N_8558,N_8142,N_8417);
and U8559 (N_8559,N_8248,N_8076);
nand U8560 (N_8560,N_8372,N_8340);
and U8561 (N_8561,N_8379,N_8305);
or U8562 (N_8562,N_8438,N_8216);
or U8563 (N_8563,N_8469,N_8449);
nand U8564 (N_8564,N_8162,N_8034);
or U8565 (N_8565,N_8296,N_8253);
xnor U8566 (N_8566,N_8081,N_8007);
or U8567 (N_8567,N_8066,N_8175);
or U8568 (N_8568,N_8493,N_8205);
xor U8569 (N_8569,N_8173,N_8192);
or U8570 (N_8570,N_8491,N_8282);
nor U8571 (N_8571,N_8164,N_8179);
xnor U8572 (N_8572,N_8407,N_8448);
and U8573 (N_8573,N_8485,N_8349);
nand U8574 (N_8574,N_8499,N_8022);
and U8575 (N_8575,N_8095,N_8317);
or U8576 (N_8576,N_8270,N_8019);
and U8577 (N_8577,N_8063,N_8129);
or U8578 (N_8578,N_8403,N_8496);
and U8579 (N_8579,N_8125,N_8244);
nand U8580 (N_8580,N_8444,N_8126);
nor U8581 (N_8581,N_8224,N_8094);
and U8582 (N_8582,N_8435,N_8459);
or U8583 (N_8583,N_8146,N_8463);
and U8584 (N_8584,N_8325,N_8446);
xor U8585 (N_8585,N_8465,N_8220);
or U8586 (N_8586,N_8388,N_8352);
and U8587 (N_8587,N_8117,N_8413);
and U8588 (N_8588,N_8277,N_8040);
or U8589 (N_8589,N_8165,N_8393);
xor U8590 (N_8590,N_8195,N_8003);
nor U8591 (N_8591,N_8454,N_8001);
and U8592 (N_8592,N_8052,N_8287);
and U8593 (N_8593,N_8059,N_8375);
or U8594 (N_8594,N_8232,N_8006);
nor U8595 (N_8595,N_8218,N_8490);
nand U8596 (N_8596,N_8275,N_8212);
and U8597 (N_8597,N_8100,N_8198);
or U8598 (N_8598,N_8194,N_8423);
nor U8599 (N_8599,N_8283,N_8025);
nor U8600 (N_8600,N_8497,N_8050);
or U8601 (N_8601,N_8437,N_8396);
or U8602 (N_8602,N_8268,N_8084);
nand U8603 (N_8603,N_8085,N_8108);
or U8604 (N_8604,N_8229,N_8404);
and U8605 (N_8605,N_8032,N_8295);
or U8606 (N_8606,N_8092,N_8269);
and U8607 (N_8607,N_8429,N_8045);
nor U8608 (N_8608,N_8345,N_8385);
nor U8609 (N_8609,N_8028,N_8492);
nor U8610 (N_8610,N_8202,N_8054);
xnor U8611 (N_8611,N_8080,N_8494);
nor U8612 (N_8612,N_8470,N_8382);
and U8613 (N_8613,N_8273,N_8401);
xnor U8614 (N_8614,N_8088,N_8369);
and U8615 (N_8615,N_8355,N_8487);
or U8616 (N_8616,N_8261,N_8097);
xor U8617 (N_8617,N_8264,N_8181);
and U8618 (N_8618,N_8412,N_8467);
xnor U8619 (N_8619,N_8009,N_8304);
nor U8620 (N_8620,N_8176,N_8368);
nor U8621 (N_8621,N_8347,N_8160);
or U8622 (N_8622,N_8285,N_8333);
nand U8623 (N_8623,N_8260,N_8062);
or U8624 (N_8624,N_8152,N_8148);
nor U8625 (N_8625,N_8137,N_8047);
or U8626 (N_8626,N_8128,N_8453);
xor U8627 (N_8627,N_8188,N_8120);
and U8628 (N_8628,N_8075,N_8381);
or U8629 (N_8629,N_8208,N_8141);
and U8630 (N_8630,N_8230,N_8197);
nor U8631 (N_8631,N_8311,N_8078);
xor U8632 (N_8632,N_8091,N_8070);
or U8633 (N_8633,N_8464,N_8055);
nor U8634 (N_8634,N_8332,N_8395);
nand U8635 (N_8635,N_8315,N_8130);
nand U8636 (N_8636,N_8133,N_8300);
nand U8637 (N_8637,N_8020,N_8098);
nand U8638 (N_8638,N_8462,N_8362);
and U8639 (N_8639,N_8239,N_8035);
nor U8640 (N_8640,N_8183,N_8326);
nor U8641 (N_8641,N_8104,N_8177);
nor U8642 (N_8642,N_8150,N_8456);
and U8643 (N_8643,N_8488,N_8155);
and U8644 (N_8644,N_8061,N_8219);
nor U8645 (N_8645,N_8374,N_8267);
or U8646 (N_8646,N_8013,N_8149);
nand U8647 (N_8647,N_8014,N_8036);
or U8648 (N_8648,N_8186,N_8017);
nand U8649 (N_8649,N_8357,N_8445);
xor U8650 (N_8650,N_8351,N_8004);
xnor U8651 (N_8651,N_8294,N_8292);
xor U8652 (N_8652,N_8144,N_8306);
nand U8653 (N_8653,N_8190,N_8167);
and U8654 (N_8654,N_8247,N_8365);
and U8655 (N_8655,N_8240,N_8236);
nor U8656 (N_8656,N_8143,N_8123);
or U8657 (N_8657,N_8342,N_8320);
nor U8658 (N_8658,N_8442,N_8472);
and U8659 (N_8659,N_8105,N_8439);
or U8660 (N_8660,N_8049,N_8330);
and U8661 (N_8661,N_8136,N_8187);
or U8662 (N_8662,N_8154,N_8151);
or U8663 (N_8663,N_8447,N_8113);
or U8664 (N_8664,N_8228,N_8293);
nor U8665 (N_8665,N_8428,N_8119);
or U8666 (N_8666,N_8301,N_8431);
nor U8667 (N_8667,N_8046,N_8452);
and U8668 (N_8668,N_8394,N_8476);
or U8669 (N_8669,N_8354,N_8419);
or U8670 (N_8670,N_8436,N_8245);
or U8671 (N_8671,N_8018,N_8204);
or U8672 (N_8672,N_8031,N_8321);
xor U8673 (N_8673,N_8259,N_8064);
or U8674 (N_8674,N_8132,N_8356);
nor U8675 (N_8675,N_8163,N_8441);
nor U8676 (N_8676,N_8458,N_8090);
nor U8677 (N_8677,N_8226,N_8312);
nor U8678 (N_8678,N_8252,N_8222);
nand U8679 (N_8679,N_8015,N_8118);
or U8680 (N_8680,N_8337,N_8339);
nor U8681 (N_8681,N_8213,N_8184);
and U8682 (N_8682,N_8169,N_8480);
nand U8683 (N_8683,N_8297,N_8079);
and U8684 (N_8684,N_8324,N_8074);
nand U8685 (N_8685,N_8434,N_8489);
and U8686 (N_8686,N_8432,N_8096);
and U8687 (N_8687,N_8389,N_8281);
nand U8688 (N_8688,N_8016,N_8166);
xnor U8689 (N_8689,N_8086,N_8109);
nor U8690 (N_8690,N_8360,N_8069);
nand U8691 (N_8691,N_8280,N_8147);
and U8692 (N_8692,N_8386,N_8377);
or U8693 (N_8693,N_8227,N_8364);
or U8694 (N_8694,N_8322,N_8457);
xnor U8695 (N_8695,N_8000,N_8200);
or U8696 (N_8696,N_8424,N_8241);
or U8697 (N_8697,N_8420,N_8279);
nand U8698 (N_8698,N_8284,N_8430);
or U8699 (N_8699,N_8384,N_8262);
nor U8700 (N_8700,N_8348,N_8089);
and U8701 (N_8701,N_8067,N_8461);
nor U8702 (N_8702,N_8409,N_8422);
nand U8703 (N_8703,N_8477,N_8153);
nand U8704 (N_8704,N_8302,N_8139);
and U8705 (N_8705,N_8112,N_8207);
nand U8706 (N_8706,N_8233,N_8156);
or U8707 (N_8707,N_8170,N_8471);
or U8708 (N_8708,N_8387,N_8101);
or U8709 (N_8709,N_8400,N_8065);
and U8710 (N_8710,N_8468,N_8411);
nand U8711 (N_8711,N_8242,N_8346);
nand U8712 (N_8712,N_8093,N_8191);
and U8713 (N_8713,N_8255,N_8196);
nor U8714 (N_8714,N_8334,N_8361);
nor U8715 (N_8715,N_8303,N_8011);
nand U8716 (N_8716,N_8180,N_8161);
and U8717 (N_8717,N_8174,N_8033);
xnor U8718 (N_8718,N_8083,N_8450);
and U8719 (N_8719,N_8486,N_8483);
nor U8720 (N_8720,N_8138,N_8481);
nor U8721 (N_8721,N_8426,N_8250);
and U8722 (N_8722,N_8114,N_8021);
and U8723 (N_8723,N_8044,N_8475);
nand U8724 (N_8724,N_8336,N_8257);
and U8725 (N_8725,N_8443,N_8071);
xor U8726 (N_8726,N_8474,N_8111);
and U8727 (N_8727,N_8235,N_8023);
nor U8728 (N_8728,N_8053,N_8087);
nor U8729 (N_8729,N_8258,N_8391);
and U8730 (N_8730,N_8331,N_8358);
nand U8731 (N_8731,N_8027,N_8201);
nand U8732 (N_8732,N_8159,N_8223);
nand U8733 (N_8733,N_8316,N_8371);
and U8734 (N_8734,N_8341,N_8237);
and U8735 (N_8735,N_8010,N_8005);
or U8736 (N_8736,N_8299,N_8122);
nor U8737 (N_8737,N_8328,N_8243);
and U8738 (N_8738,N_8209,N_8495);
and U8739 (N_8739,N_8276,N_8127);
nor U8740 (N_8740,N_8060,N_8041);
and U8741 (N_8741,N_8030,N_8405);
or U8742 (N_8742,N_8254,N_8366);
nand U8743 (N_8743,N_8121,N_8319);
nor U8744 (N_8744,N_8251,N_8290);
and U8745 (N_8745,N_8115,N_8158);
nand U8746 (N_8746,N_8440,N_8390);
xnor U8747 (N_8747,N_8131,N_8124);
nor U8748 (N_8748,N_8072,N_8231);
nor U8749 (N_8749,N_8265,N_8399);
xnor U8750 (N_8750,N_8350,N_8357);
and U8751 (N_8751,N_8144,N_8061);
or U8752 (N_8752,N_8434,N_8097);
nor U8753 (N_8753,N_8410,N_8458);
or U8754 (N_8754,N_8196,N_8090);
or U8755 (N_8755,N_8402,N_8198);
or U8756 (N_8756,N_8216,N_8469);
nor U8757 (N_8757,N_8208,N_8309);
nand U8758 (N_8758,N_8205,N_8303);
nand U8759 (N_8759,N_8222,N_8119);
nand U8760 (N_8760,N_8346,N_8323);
xnor U8761 (N_8761,N_8167,N_8238);
nor U8762 (N_8762,N_8326,N_8375);
and U8763 (N_8763,N_8405,N_8378);
and U8764 (N_8764,N_8271,N_8258);
nand U8765 (N_8765,N_8455,N_8301);
xnor U8766 (N_8766,N_8007,N_8207);
nand U8767 (N_8767,N_8324,N_8023);
nand U8768 (N_8768,N_8455,N_8093);
xor U8769 (N_8769,N_8365,N_8206);
xnor U8770 (N_8770,N_8225,N_8317);
nand U8771 (N_8771,N_8398,N_8140);
xor U8772 (N_8772,N_8328,N_8298);
and U8773 (N_8773,N_8285,N_8310);
and U8774 (N_8774,N_8085,N_8347);
nand U8775 (N_8775,N_8134,N_8467);
xor U8776 (N_8776,N_8340,N_8461);
nor U8777 (N_8777,N_8035,N_8204);
xnor U8778 (N_8778,N_8087,N_8011);
and U8779 (N_8779,N_8161,N_8013);
and U8780 (N_8780,N_8466,N_8396);
xnor U8781 (N_8781,N_8418,N_8286);
or U8782 (N_8782,N_8285,N_8453);
or U8783 (N_8783,N_8338,N_8416);
nand U8784 (N_8784,N_8221,N_8116);
xor U8785 (N_8785,N_8255,N_8284);
and U8786 (N_8786,N_8058,N_8483);
nor U8787 (N_8787,N_8042,N_8088);
nor U8788 (N_8788,N_8412,N_8367);
or U8789 (N_8789,N_8260,N_8193);
or U8790 (N_8790,N_8398,N_8405);
nor U8791 (N_8791,N_8491,N_8214);
nor U8792 (N_8792,N_8361,N_8032);
or U8793 (N_8793,N_8493,N_8333);
or U8794 (N_8794,N_8317,N_8413);
and U8795 (N_8795,N_8360,N_8473);
xnor U8796 (N_8796,N_8480,N_8378);
and U8797 (N_8797,N_8198,N_8266);
and U8798 (N_8798,N_8374,N_8275);
nor U8799 (N_8799,N_8489,N_8412);
or U8800 (N_8800,N_8001,N_8064);
nand U8801 (N_8801,N_8294,N_8487);
and U8802 (N_8802,N_8039,N_8425);
nor U8803 (N_8803,N_8208,N_8261);
and U8804 (N_8804,N_8007,N_8233);
and U8805 (N_8805,N_8057,N_8134);
nor U8806 (N_8806,N_8374,N_8148);
and U8807 (N_8807,N_8403,N_8140);
nor U8808 (N_8808,N_8233,N_8281);
and U8809 (N_8809,N_8353,N_8010);
xnor U8810 (N_8810,N_8325,N_8166);
nand U8811 (N_8811,N_8414,N_8205);
and U8812 (N_8812,N_8461,N_8366);
or U8813 (N_8813,N_8474,N_8462);
nand U8814 (N_8814,N_8118,N_8179);
or U8815 (N_8815,N_8239,N_8123);
xor U8816 (N_8816,N_8253,N_8455);
and U8817 (N_8817,N_8313,N_8254);
xor U8818 (N_8818,N_8116,N_8106);
nor U8819 (N_8819,N_8350,N_8010);
xor U8820 (N_8820,N_8126,N_8269);
nand U8821 (N_8821,N_8094,N_8483);
or U8822 (N_8822,N_8320,N_8317);
and U8823 (N_8823,N_8276,N_8176);
or U8824 (N_8824,N_8460,N_8142);
nand U8825 (N_8825,N_8459,N_8135);
nand U8826 (N_8826,N_8296,N_8266);
nor U8827 (N_8827,N_8049,N_8234);
and U8828 (N_8828,N_8020,N_8024);
or U8829 (N_8829,N_8135,N_8463);
or U8830 (N_8830,N_8380,N_8063);
xor U8831 (N_8831,N_8214,N_8109);
and U8832 (N_8832,N_8423,N_8400);
or U8833 (N_8833,N_8031,N_8290);
and U8834 (N_8834,N_8348,N_8168);
nor U8835 (N_8835,N_8342,N_8484);
nand U8836 (N_8836,N_8109,N_8020);
or U8837 (N_8837,N_8339,N_8426);
or U8838 (N_8838,N_8438,N_8098);
nor U8839 (N_8839,N_8094,N_8294);
nor U8840 (N_8840,N_8304,N_8171);
nor U8841 (N_8841,N_8313,N_8307);
and U8842 (N_8842,N_8222,N_8402);
and U8843 (N_8843,N_8325,N_8183);
or U8844 (N_8844,N_8205,N_8207);
nand U8845 (N_8845,N_8398,N_8143);
or U8846 (N_8846,N_8045,N_8113);
xnor U8847 (N_8847,N_8162,N_8388);
nand U8848 (N_8848,N_8060,N_8202);
nor U8849 (N_8849,N_8320,N_8452);
nor U8850 (N_8850,N_8150,N_8023);
xor U8851 (N_8851,N_8045,N_8196);
nand U8852 (N_8852,N_8459,N_8164);
nand U8853 (N_8853,N_8396,N_8009);
nor U8854 (N_8854,N_8078,N_8083);
nor U8855 (N_8855,N_8232,N_8019);
or U8856 (N_8856,N_8388,N_8463);
and U8857 (N_8857,N_8496,N_8283);
and U8858 (N_8858,N_8072,N_8419);
xor U8859 (N_8859,N_8305,N_8499);
and U8860 (N_8860,N_8204,N_8237);
nand U8861 (N_8861,N_8050,N_8137);
nor U8862 (N_8862,N_8013,N_8210);
and U8863 (N_8863,N_8428,N_8036);
nor U8864 (N_8864,N_8229,N_8490);
or U8865 (N_8865,N_8405,N_8044);
nor U8866 (N_8866,N_8183,N_8073);
nor U8867 (N_8867,N_8425,N_8098);
and U8868 (N_8868,N_8164,N_8188);
nand U8869 (N_8869,N_8494,N_8296);
or U8870 (N_8870,N_8476,N_8433);
or U8871 (N_8871,N_8250,N_8334);
nor U8872 (N_8872,N_8367,N_8009);
nor U8873 (N_8873,N_8286,N_8391);
nand U8874 (N_8874,N_8350,N_8051);
and U8875 (N_8875,N_8035,N_8482);
xor U8876 (N_8876,N_8432,N_8094);
nor U8877 (N_8877,N_8060,N_8313);
or U8878 (N_8878,N_8118,N_8488);
nor U8879 (N_8879,N_8420,N_8305);
xor U8880 (N_8880,N_8427,N_8454);
nand U8881 (N_8881,N_8036,N_8338);
nand U8882 (N_8882,N_8056,N_8050);
or U8883 (N_8883,N_8019,N_8224);
and U8884 (N_8884,N_8040,N_8448);
nand U8885 (N_8885,N_8476,N_8349);
nor U8886 (N_8886,N_8470,N_8223);
or U8887 (N_8887,N_8477,N_8467);
nand U8888 (N_8888,N_8149,N_8330);
or U8889 (N_8889,N_8349,N_8455);
nor U8890 (N_8890,N_8041,N_8486);
and U8891 (N_8891,N_8060,N_8151);
xnor U8892 (N_8892,N_8230,N_8199);
nor U8893 (N_8893,N_8104,N_8037);
and U8894 (N_8894,N_8455,N_8452);
nand U8895 (N_8895,N_8162,N_8220);
or U8896 (N_8896,N_8122,N_8475);
nor U8897 (N_8897,N_8312,N_8216);
or U8898 (N_8898,N_8430,N_8051);
or U8899 (N_8899,N_8459,N_8485);
nor U8900 (N_8900,N_8202,N_8015);
nand U8901 (N_8901,N_8035,N_8470);
nor U8902 (N_8902,N_8318,N_8444);
and U8903 (N_8903,N_8336,N_8488);
nor U8904 (N_8904,N_8298,N_8263);
nand U8905 (N_8905,N_8346,N_8104);
and U8906 (N_8906,N_8111,N_8317);
or U8907 (N_8907,N_8452,N_8469);
nor U8908 (N_8908,N_8245,N_8494);
and U8909 (N_8909,N_8136,N_8070);
or U8910 (N_8910,N_8383,N_8088);
and U8911 (N_8911,N_8048,N_8073);
nand U8912 (N_8912,N_8055,N_8297);
nand U8913 (N_8913,N_8001,N_8371);
or U8914 (N_8914,N_8402,N_8479);
xor U8915 (N_8915,N_8218,N_8141);
nand U8916 (N_8916,N_8302,N_8091);
nand U8917 (N_8917,N_8336,N_8367);
nor U8918 (N_8918,N_8362,N_8013);
and U8919 (N_8919,N_8165,N_8282);
and U8920 (N_8920,N_8143,N_8264);
and U8921 (N_8921,N_8260,N_8161);
and U8922 (N_8922,N_8322,N_8173);
nor U8923 (N_8923,N_8314,N_8489);
nor U8924 (N_8924,N_8303,N_8323);
and U8925 (N_8925,N_8059,N_8104);
nand U8926 (N_8926,N_8360,N_8064);
and U8927 (N_8927,N_8378,N_8023);
nand U8928 (N_8928,N_8084,N_8272);
nand U8929 (N_8929,N_8085,N_8372);
and U8930 (N_8930,N_8304,N_8114);
and U8931 (N_8931,N_8130,N_8416);
and U8932 (N_8932,N_8059,N_8312);
xor U8933 (N_8933,N_8035,N_8133);
or U8934 (N_8934,N_8266,N_8128);
and U8935 (N_8935,N_8055,N_8219);
or U8936 (N_8936,N_8482,N_8195);
and U8937 (N_8937,N_8087,N_8231);
and U8938 (N_8938,N_8143,N_8186);
nand U8939 (N_8939,N_8248,N_8152);
xnor U8940 (N_8940,N_8294,N_8373);
and U8941 (N_8941,N_8134,N_8403);
or U8942 (N_8942,N_8451,N_8492);
nand U8943 (N_8943,N_8131,N_8391);
xor U8944 (N_8944,N_8017,N_8285);
xnor U8945 (N_8945,N_8326,N_8241);
or U8946 (N_8946,N_8009,N_8038);
xnor U8947 (N_8947,N_8146,N_8202);
xor U8948 (N_8948,N_8345,N_8321);
nand U8949 (N_8949,N_8215,N_8032);
or U8950 (N_8950,N_8250,N_8287);
nand U8951 (N_8951,N_8366,N_8253);
nor U8952 (N_8952,N_8210,N_8272);
nor U8953 (N_8953,N_8320,N_8419);
and U8954 (N_8954,N_8497,N_8129);
nand U8955 (N_8955,N_8340,N_8243);
nor U8956 (N_8956,N_8123,N_8007);
nand U8957 (N_8957,N_8284,N_8055);
and U8958 (N_8958,N_8100,N_8193);
nand U8959 (N_8959,N_8109,N_8332);
and U8960 (N_8960,N_8465,N_8421);
and U8961 (N_8961,N_8120,N_8326);
and U8962 (N_8962,N_8323,N_8471);
or U8963 (N_8963,N_8254,N_8465);
nor U8964 (N_8964,N_8438,N_8260);
and U8965 (N_8965,N_8492,N_8388);
nand U8966 (N_8966,N_8096,N_8151);
nand U8967 (N_8967,N_8003,N_8088);
nor U8968 (N_8968,N_8062,N_8435);
nor U8969 (N_8969,N_8327,N_8481);
and U8970 (N_8970,N_8173,N_8318);
or U8971 (N_8971,N_8485,N_8256);
nand U8972 (N_8972,N_8362,N_8484);
or U8973 (N_8973,N_8241,N_8320);
xnor U8974 (N_8974,N_8385,N_8038);
nor U8975 (N_8975,N_8299,N_8400);
and U8976 (N_8976,N_8212,N_8083);
and U8977 (N_8977,N_8452,N_8082);
nor U8978 (N_8978,N_8005,N_8071);
nand U8979 (N_8979,N_8117,N_8417);
or U8980 (N_8980,N_8495,N_8474);
xor U8981 (N_8981,N_8072,N_8244);
nand U8982 (N_8982,N_8429,N_8042);
or U8983 (N_8983,N_8222,N_8155);
nor U8984 (N_8984,N_8011,N_8039);
nand U8985 (N_8985,N_8188,N_8233);
nand U8986 (N_8986,N_8407,N_8405);
nand U8987 (N_8987,N_8234,N_8027);
nor U8988 (N_8988,N_8388,N_8070);
nor U8989 (N_8989,N_8253,N_8089);
or U8990 (N_8990,N_8128,N_8006);
and U8991 (N_8991,N_8061,N_8201);
and U8992 (N_8992,N_8153,N_8369);
or U8993 (N_8993,N_8355,N_8212);
or U8994 (N_8994,N_8329,N_8410);
or U8995 (N_8995,N_8102,N_8432);
nor U8996 (N_8996,N_8484,N_8068);
or U8997 (N_8997,N_8157,N_8319);
nand U8998 (N_8998,N_8415,N_8166);
nor U8999 (N_8999,N_8199,N_8042);
or U9000 (N_9000,N_8690,N_8620);
nand U9001 (N_9001,N_8589,N_8987);
nor U9002 (N_9002,N_8972,N_8651);
and U9003 (N_9003,N_8902,N_8520);
and U9004 (N_9004,N_8527,N_8772);
or U9005 (N_9005,N_8901,N_8704);
nor U9006 (N_9006,N_8695,N_8908);
nand U9007 (N_9007,N_8819,N_8991);
nand U9008 (N_9008,N_8581,N_8788);
or U9009 (N_9009,N_8956,N_8674);
nand U9010 (N_9010,N_8750,N_8977);
nand U9011 (N_9011,N_8538,N_8687);
or U9012 (N_9012,N_8873,N_8967);
and U9013 (N_9013,N_8872,N_8613);
nor U9014 (N_9014,N_8910,N_8636);
or U9015 (N_9015,N_8714,N_8753);
xnor U9016 (N_9016,N_8610,N_8524);
nand U9017 (N_9017,N_8791,N_8707);
or U9018 (N_9018,N_8978,N_8778);
nor U9019 (N_9019,N_8507,N_8986);
and U9020 (N_9020,N_8775,N_8784);
and U9021 (N_9021,N_8523,N_8717);
nand U9022 (N_9022,N_8631,N_8734);
or U9023 (N_9023,N_8701,N_8746);
nor U9024 (N_9024,N_8948,N_8659);
nor U9025 (N_9025,N_8502,N_8737);
and U9026 (N_9026,N_8995,N_8592);
nor U9027 (N_9027,N_8799,N_8670);
or U9028 (N_9028,N_8839,N_8661);
and U9029 (N_9029,N_8993,N_8795);
nor U9030 (N_9030,N_8961,N_8685);
nand U9031 (N_9031,N_8899,N_8843);
and U9032 (N_9032,N_8833,N_8660);
nor U9033 (N_9033,N_8876,N_8877);
nor U9034 (N_9034,N_8745,N_8920);
nor U9035 (N_9035,N_8886,N_8878);
and U9036 (N_9036,N_8881,N_8890);
nor U9037 (N_9037,N_8529,N_8728);
xnor U9038 (N_9038,N_8990,N_8533);
and U9039 (N_9039,N_8758,N_8548);
nor U9040 (N_9040,N_8504,N_8710);
and U9041 (N_9041,N_8976,N_8582);
nand U9042 (N_9042,N_8935,N_8915);
and U9043 (N_9043,N_8852,N_8702);
and U9044 (N_9044,N_8535,N_8836);
nor U9045 (N_9045,N_8512,N_8882);
and U9046 (N_9046,N_8585,N_8733);
or U9047 (N_9047,N_8954,N_8681);
nor U9048 (N_9048,N_8834,N_8864);
and U9049 (N_9049,N_8642,N_8942);
nand U9050 (N_9050,N_8937,N_8835);
nor U9051 (N_9051,N_8676,N_8771);
nor U9052 (N_9052,N_8898,N_8511);
and U9053 (N_9053,N_8951,N_8632);
nand U9054 (N_9054,N_8801,N_8787);
and U9055 (N_9055,N_8906,N_8696);
nor U9056 (N_9056,N_8798,N_8828);
and U9057 (N_9057,N_8536,N_8938);
nand U9058 (N_9058,N_8974,N_8565);
or U9059 (N_9059,N_8561,N_8860);
or U9060 (N_9060,N_8541,N_8894);
or U9061 (N_9061,N_8970,N_8503);
or U9062 (N_9062,N_8577,N_8692);
nor U9063 (N_9063,N_8919,N_8576);
xor U9064 (N_9064,N_8516,N_8904);
and U9065 (N_9065,N_8999,N_8514);
nand U9066 (N_9066,N_8797,N_8715);
nand U9067 (N_9067,N_8664,N_8840);
and U9068 (N_9068,N_8587,N_8963);
nor U9069 (N_9069,N_8545,N_8558);
or U9070 (N_9070,N_8760,N_8542);
nor U9071 (N_9071,N_8985,N_8648);
nor U9072 (N_9072,N_8818,N_8764);
nor U9073 (N_9073,N_8614,N_8794);
and U9074 (N_9074,N_8907,N_8738);
or U9075 (N_9075,N_8781,N_8930);
nand U9076 (N_9076,N_8796,N_8622);
or U9077 (N_9077,N_8885,N_8824);
or U9078 (N_9078,N_8774,N_8591);
xor U9079 (N_9079,N_8950,N_8727);
and U9080 (N_9080,N_8996,N_8900);
nor U9081 (N_9081,N_8645,N_8735);
or U9082 (N_9082,N_8816,N_8669);
or U9083 (N_9083,N_8705,N_8983);
and U9084 (N_9084,N_8868,N_8509);
nand U9085 (N_9085,N_8875,N_8675);
or U9086 (N_9086,N_8556,N_8744);
and U9087 (N_9087,N_8962,N_8914);
nand U9088 (N_9088,N_8838,N_8643);
and U9089 (N_9089,N_8924,N_8629);
nand U9090 (N_9090,N_8953,N_8667);
and U9091 (N_9091,N_8747,N_8644);
or U9092 (N_9092,N_8709,N_8537);
or U9093 (N_9093,N_8992,N_8555);
nand U9094 (N_9094,N_8673,N_8525);
and U9095 (N_9095,N_8688,N_8552);
or U9096 (N_9096,N_8965,N_8566);
and U9097 (N_9097,N_8989,N_8815);
and U9098 (N_9098,N_8943,N_8739);
nand U9099 (N_9099,N_8652,N_8519);
or U9100 (N_9100,N_8742,N_8874);
nand U9101 (N_9101,N_8543,N_8599);
nor U9102 (N_9102,N_8813,N_8982);
xor U9103 (N_9103,N_8579,N_8934);
nor U9104 (N_9104,N_8889,N_8679);
nand U9105 (N_9105,N_8888,N_8949);
nand U9106 (N_9106,N_8699,N_8847);
or U9107 (N_9107,N_8724,N_8790);
and U9108 (N_9108,N_8909,N_8749);
or U9109 (N_9109,N_8647,N_8891);
nand U9110 (N_9110,N_8770,N_8553);
nor U9111 (N_9111,N_8827,N_8743);
or U9112 (N_9112,N_8947,N_8918);
xor U9113 (N_9113,N_8850,N_8812);
and U9114 (N_9114,N_8912,N_8626);
and U9115 (N_9115,N_8941,N_8522);
or U9116 (N_9116,N_8865,N_8789);
or U9117 (N_9117,N_8609,N_8571);
or U9118 (N_9118,N_8831,N_8929);
nand U9119 (N_9119,N_8557,N_8844);
and U9120 (N_9120,N_8546,N_8826);
or U9121 (N_9121,N_8741,N_8973);
nand U9122 (N_9122,N_8500,N_8646);
or U9123 (N_9123,N_8513,N_8731);
and U9124 (N_9124,N_8584,N_8586);
nor U9125 (N_9125,N_8800,N_8596);
or U9126 (N_9126,N_8637,N_8508);
nor U9127 (N_9127,N_8806,N_8672);
nand U9128 (N_9128,N_8867,N_8945);
and U9129 (N_9129,N_8928,N_8563);
or U9130 (N_9130,N_8720,N_8857);
xor U9131 (N_9131,N_8998,N_8805);
and U9132 (N_9132,N_8879,N_8666);
xor U9133 (N_9133,N_8602,N_8628);
and U9134 (N_9134,N_8649,N_8547);
or U9135 (N_9135,N_8922,N_8521);
or U9136 (N_9136,N_8600,N_8594);
or U9137 (N_9137,N_8767,N_8994);
and U9138 (N_9138,N_8944,N_8754);
xnor U9139 (N_9139,N_8638,N_8969);
nand U9140 (N_9140,N_8686,N_8780);
nand U9141 (N_9141,N_8939,N_8802);
and U9142 (N_9142,N_8958,N_8984);
xor U9143 (N_9143,N_8593,N_8940);
nand U9144 (N_9144,N_8856,N_8716);
nor U9145 (N_9145,N_8655,N_8708);
and U9146 (N_9146,N_8793,N_8682);
and U9147 (N_9147,N_8913,N_8751);
nand U9148 (N_9148,N_8884,N_8841);
nor U9149 (N_9149,N_8825,N_8678);
nor U9150 (N_9150,N_8763,N_8859);
or U9151 (N_9151,N_8641,N_8849);
nand U9152 (N_9152,N_8534,N_8830);
nor U9153 (N_9153,N_8663,N_8662);
or U9154 (N_9154,N_8677,N_8607);
nor U9155 (N_9155,N_8730,N_8615);
nor U9156 (N_9156,N_8765,N_8931);
and U9157 (N_9157,N_8554,N_8959);
xnor U9158 (N_9158,N_8808,N_8926);
nor U9159 (N_9159,N_8955,N_8532);
and U9160 (N_9160,N_8619,N_8777);
and U9161 (N_9161,N_8603,N_8568);
or U9162 (N_9162,N_8980,N_8927);
or U9163 (N_9163,N_8869,N_8779);
and U9164 (N_9164,N_8703,N_8654);
and U9165 (N_9165,N_8769,N_8700);
and U9166 (N_9166,N_8544,N_8570);
and U9167 (N_9167,N_8783,N_8505);
nand U9168 (N_9168,N_8979,N_8946);
or U9169 (N_9169,N_8729,N_8866);
and U9170 (N_9170,N_8625,N_8921);
nor U9171 (N_9171,N_8668,N_8761);
nor U9172 (N_9172,N_8905,N_8863);
or U9173 (N_9173,N_8851,N_8573);
nor U9174 (N_9174,N_8804,N_8639);
or U9175 (N_9175,N_8633,N_8706);
and U9176 (N_9176,N_8810,N_8698);
nand U9177 (N_9177,N_8575,N_8786);
nor U9178 (N_9178,N_8691,N_8526);
or U9179 (N_9179,N_8528,N_8694);
nand U9180 (N_9180,N_8846,N_8635);
nand U9181 (N_9181,N_8968,N_8721);
nor U9182 (N_9182,N_8932,N_8562);
and U9183 (N_9183,N_8680,N_8829);
or U9184 (N_9184,N_8768,N_8870);
xnor U9185 (N_9185,N_8848,N_8773);
nand U9186 (N_9186,N_8792,N_8854);
and U9187 (N_9187,N_8871,N_8740);
nor U9188 (N_9188,N_8853,N_8551);
nand U9189 (N_9189,N_8578,N_8975);
xnor U9190 (N_9190,N_8895,N_8506);
nand U9191 (N_9191,N_8736,N_8595);
nand U9192 (N_9192,N_8725,N_8823);
or U9193 (N_9193,N_8605,N_8640);
nor U9194 (N_9194,N_8693,N_8903);
nand U9195 (N_9195,N_8936,N_8539);
xnor U9196 (N_9196,N_8683,N_8712);
and U9197 (N_9197,N_8656,N_8684);
nand U9198 (N_9198,N_8757,N_8518);
and U9199 (N_9199,N_8583,N_8617);
nand U9200 (N_9200,N_8776,N_8722);
or U9201 (N_9201,N_8964,N_8892);
xor U9202 (N_9202,N_8897,N_8861);
nand U9203 (N_9203,N_8862,N_8650);
nor U9204 (N_9204,N_8837,N_8611);
or U9205 (N_9205,N_8665,N_8971);
or U9206 (N_9206,N_8569,N_8608);
nand U9207 (N_9207,N_8560,N_8820);
nand U9208 (N_9208,N_8814,N_8766);
nor U9209 (N_9209,N_8887,N_8621);
and U9210 (N_9210,N_8723,N_8726);
and U9211 (N_9211,N_8550,N_8574);
and U9212 (N_9212,N_8845,N_8785);
and U9213 (N_9213,N_8858,N_8671);
or U9214 (N_9214,N_8719,N_8917);
xnor U9215 (N_9215,N_8597,N_8606);
xnor U9216 (N_9216,N_8713,N_8822);
or U9217 (N_9217,N_8997,N_8634);
and U9218 (N_9218,N_8756,N_8653);
nand U9219 (N_9219,N_8925,N_8981);
nand U9220 (N_9220,N_8759,N_8697);
or U9221 (N_9221,N_8811,N_8817);
nor U9222 (N_9222,N_8515,N_8598);
nor U9223 (N_9223,N_8842,N_8896);
nand U9224 (N_9224,N_8782,N_8923);
nor U9225 (N_9225,N_8933,N_8624);
nor U9226 (N_9226,N_8517,N_8880);
and U9227 (N_9227,N_8689,N_8531);
nor U9228 (N_9228,N_8809,N_8572);
nor U9229 (N_9229,N_8893,N_8630);
and U9230 (N_9230,N_8952,N_8618);
nand U9231 (N_9231,N_8807,N_8752);
and U9232 (N_9232,N_8916,N_8530);
or U9233 (N_9233,N_8604,N_8658);
and U9234 (N_9234,N_8657,N_8748);
xnor U9235 (N_9235,N_8755,N_8616);
nor U9236 (N_9236,N_8623,N_8960);
or U9237 (N_9237,N_8559,N_8510);
or U9238 (N_9238,N_8612,N_8564);
and U9239 (N_9239,N_8732,N_8567);
or U9240 (N_9240,N_8988,N_8549);
nor U9241 (N_9241,N_8803,N_8627);
nor U9242 (N_9242,N_8601,N_8580);
nor U9243 (N_9243,N_8911,N_8501);
nand U9244 (N_9244,N_8821,N_8832);
or U9245 (N_9245,N_8588,N_8718);
nand U9246 (N_9246,N_8855,N_8590);
xnor U9247 (N_9247,N_8966,N_8540);
or U9248 (N_9248,N_8883,N_8957);
nand U9249 (N_9249,N_8762,N_8711);
nand U9250 (N_9250,N_8846,N_8802);
nand U9251 (N_9251,N_8940,N_8728);
and U9252 (N_9252,N_8993,N_8857);
or U9253 (N_9253,N_8610,N_8520);
and U9254 (N_9254,N_8963,N_8596);
xnor U9255 (N_9255,N_8511,N_8820);
or U9256 (N_9256,N_8845,N_8651);
and U9257 (N_9257,N_8576,N_8912);
xor U9258 (N_9258,N_8547,N_8647);
nor U9259 (N_9259,N_8928,N_8732);
nand U9260 (N_9260,N_8615,N_8670);
nor U9261 (N_9261,N_8976,N_8827);
and U9262 (N_9262,N_8532,N_8744);
nor U9263 (N_9263,N_8503,N_8641);
and U9264 (N_9264,N_8504,N_8756);
and U9265 (N_9265,N_8656,N_8540);
and U9266 (N_9266,N_8712,N_8804);
or U9267 (N_9267,N_8803,N_8625);
and U9268 (N_9268,N_8607,N_8857);
nor U9269 (N_9269,N_8990,N_8959);
nand U9270 (N_9270,N_8679,N_8528);
or U9271 (N_9271,N_8632,N_8762);
nor U9272 (N_9272,N_8768,N_8889);
nor U9273 (N_9273,N_8638,N_8822);
nor U9274 (N_9274,N_8942,N_8710);
and U9275 (N_9275,N_8500,N_8664);
and U9276 (N_9276,N_8966,N_8855);
nor U9277 (N_9277,N_8955,N_8920);
or U9278 (N_9278,N_8975,N_8967);
nand U9279 (N_9279,N_8991,N_8939);
xor U9280 (N_9280,N_8992,N_8859);
xnor U9281 (N_9281,N_8731,N_8659);
xor U9282 (N_9282,N_8623,N_8587);
nor U9283 (N_9283,N_8746,N_8846);
or U9284 (N_9284,N_8549,N_8759);
and U9285 (N_9285,N_8698,N_8523);
or U9286 (N_9286,N_8523,N_8623);
and U9287 (N_9287,N_8636,N_8672);
xor U9288 (N_9288,N_8899,N_8510);
nor U9289 (N_9289,N_8949,N_8722);
or U9290 (N_9290,N_8998,N_8806);
or U9291 (N_9291,N_8780,N_8642);
or U9292 (N_9292,N_8926,N_8979);
and U9293 (N_9293,N_8533,N_8965);
nand U9294 (N_9294,N_8893,N_8573);
or U9295 (N_9295,N_8848,N_8696);
or U9296 (N_9296,N_8943,N_8902);
and U9297 (N_9297,N_8885,N_8553);
xor U9298 (N_9298,N_8754,N_8727);
and U9299 (N_9299,N_8698,N_8671);
or U9300 (N_9300,N_8718,N_8965);
nand U9301 (N_9301,N_8865,N_8784);
nand U9302 (N_9302,N_8688,N_8648);
and U9303 (N_9303,N_8880,N_8727);
nor U9304 (N_9304,N_8968,N_8861);
xnor U9305 (N_9305,N_8517,N_8874);
or U9306 (N_9306,N_8995,N_8789);
and U9307 (N_9307,N_8627,N_8618);
and U9308 (N_9308,N_8799,N_8836);
or U9309 (N_9309,N_8693,N_8995);
or U9310 (N_9310,N_8967,N_8800);
nor U9311 (N_9311,N_8966,N_8981);
and U9312 (N_9312,N_8900,N_8699);
nand U9313 (N_9313,N_8906,N_8826);
nor U9314 (N_9314,N_8825,N_8587);
nor U9315 (N_9315,N_8982,N_8600);
nor U9316 (N_9316,N_8659,N_8907);
and U9317 (N_9317,N_8961,N_8641);
nand U9318 (N_9318,N_8530,N_8738);
and U9319 (N_9319,N_8567,N_8836);
xnor U9320 (N_9320,N_8563,N_8708);
and U9321 (N_9321,N_8935,N_8828);
nor U9322 (N_9322,N_8564,N_8680);
and U9323 (N_9323,N_8527,N_8875);
nand U9324 (N_9324,N_8786,N_8627);
or U9325 (N_9325,N_8708,N_8889);
and U9326 (N_9326,N_8829,N_8719);
nor U9327 (N_9327,N_8783,N_8905);
nand U9328 (N_9328,N_8771,N_8834);
xor U9329 (N_9329,N_8518,N_8921);
nor U9330 (N_9330,N_8998,N_8699);
or U9331 (N_9331,N_8631,N_8788);
and U9332 (N_9332,N_8552,N_8862);
xnor U9333 (N_9333,N_8861,N_8600);
nand U9334 (N_9334,N_8533,N_8524);
nand U9335 (N_9335,N_8913,N_8709);
and U9336 (N_9336,N_8543,N_8857);
nor U9337 (N_9337,N_8832,N_8815);
nand U9338 (N_9338,N_8694,N_8604);
or U9339 (N_9339,N_8503,N_8998);
nor U9340 (N_9340,N_8978,N_8594);
xnor U9341 (N_9341,N_8930,N_8915);
nor U9342 (N_9342,N_8691,N_8848);
nand U9343 (N_9343,N_8972,N_8514);
and U9344 (N_9344,N_8768,N_8848);
nand U9345 (N_9345,N_8682,N_8844);
nand U9346 (N_9346,N_8891,N_8677);
nand U9347 (N_9347,N_8906,N_8615);
nor U9348 (N_9348,N_8872,N_8585);
nor U9349 (N_9349,N_8632,N_8862);
or U9350 (N_9350,N_8942,N_8726);
nor U9351 (N_9351,N_8838,N_8819);
nand U9352 (N_9352,N_8795,N_8505);
nand U9353 (N_9353,N_8986,N_8855);
nand U9354 (N_9354,N_8559,N_8526);
and U9355 (N_9355,N_8583,N_8818);
or U9356 (N_9356,N_8991,N_8697);
or U9357 (N_9357,N_8574,N_8741);
nand U9358 (N_9358,N_8654,N_8628);
or U9359 (N_9359,N_8620,N_8635);
nand U9360 (N_9360,N_8567,N_8716);
and U9361 (N_9361,N_8527,N_8680);
and U9362 (N_9362,N_8755,N_8972);
or U9363 (N_9363,N_8746,N_8629);
or U9364 (N_9364,N_8738,N_8789);
or U9365 (N_9365,N_8842,N_8854);
and U9366 (N_9366,N_8708,N_8768);
or U9367 (N_9367,N_8840,N_8509);
xnor U9368 (N_9368,N_8735,N_8930);
nand U9369 (N_9369,N_8515,N_8881);
nor U9370 (N_9370,N_8525,N_8903);
and U9371 (N_9371,N_8730,N_8644);
nand U9372 (N_9372,N_8664,N_8763);
nor U9373 (N_9373,N_8700,N_8604);
and U9374 (N_9374,N_8821,N_8881);
and U9375 (N_9375,N_8705,N_8698);
nand U9376 (N_9376,N_8985,N_8723);
nand U9377 (N_9377,N_8648,N_8504);
nand U9378 (N_9378,N_8932,N_8757);
or U9379 (N_9379,N_8821,N_8955);
nand U9380 (N_9380,N_8600,N_8634);
nor U9381 (N_9381,N_8612,N_8885);
nor U9382 (N_9382,N_8796,N_8514);
nand U9383 (N_9383,N_8782,N_8973);
and U9384 (N_9384,N_8946,N_8955);
or U9385 (N_9385,N_8679,N_8589);
and U9386 (N_9386,N_8806,N_8994);
or U9387 (N_9387,N_8516,N_8937);
nor U9388 (N_9388,N_8813,N_8722);
or U9389 (N_9389,N_8596,N_8889);
xor U9390 (N_9390,N_8529,N_8982);
or U9391 (N_9391,N_8805,N_8578);
nor U9392 (N_9392,N_8833,N_8647);
or U9393 (N_9393,N_8864,N_8986);
nor U9394 (N_9394,N_8745,N_8532);
or U9395 (N_9395,N_8827,N_8529);
or U9396 (N_9396,N_8838,N_8534);
nor U9397 (N_9397,N_8500,N_8562);
nor U9398 (N_9398,N_8678,N_8649);
xnor U9399 (N_9399,N_8841,N_8856);
or U9400 (N_9400,N_8645,N_8666);
xnor U9401 (N_9401,N_8895,N_8936);
or U9402 (N_9402,N_8772,N_8656);
nor U9403 (N_9403,N_8851,N_8512);
nand U9404 (N_9404,N_8848,N_8981);
nor U9405 (N_9405,N_8989,N_8739);
xnor U9406 (N_9406,N_8574,N_8694);
nor U9407 (N_9407,N_8726,N_8806);
nor U9408 (N_9408,N_8522,N_8775);
nand U9409 (N_9409,N_8742,N_8837);
xnor U9410 (N_9410,N_8880,N_8977);
and U9411 (N_9411,N_8755,N_8768);
and U9412 (N_9412,N_8966,N_8953);
and U9413 (N_9413,N_8982,N_8876);
or U9414 (N_9414,N_8620,N_8876);
nand U9415 (N_9415,N_8641,N_8810);
nand U9416 (N_9416,N_8571,N_8870);
or U9417 (N_9417,N_8723,N_8627);
nand U9418 (N_9418,N_8889,N_8801);
and U9419 (N_9419,N_8666,N_8608);
nand U9420 (N_9420,N_8809,N_8915);
xnor U9421 (N_9421,N_8514,N_8636);
nor U9422 (N_9422,N_8754,N_8949);
nand U9423 (N_9423,N_8555,N_8673);
and U9424 (N_9424,N_8500,N_8560);
or U9425 (N_9425,N_8949,N_8730);
or U9426 (N_9426,N_8591,N_8655);
or U9427 (N_9427,N_8521,N_8773);
or U9428 (N_9428,N_8972,N_8976);
nand U9429 (N_9429,N_8868,N_8597);
nand U9430 (N_9430,N_8563,N_8631);
nor U9431 (N_9431,N_8848,N_8734);
nand U9432 (N_9432,N_8509,N_8577);
xnor U9433 (N_9433,N_8742,N_8938);
nand U9434 (N_9434,N_8671,N_8908);
or U9435 (N_9435,N_8939,N_8897);
nor U9436 (N_9436,N_8988,N_8697);
xor U9437 (N_9437,N_8800,N_8503);
nor U9438 (N_9438,N_8615,N_8599);
nor U9439 (N_9439,N_8863,N_8849);
or U9440 (N_9440,N_8667,N_8777);
xnor U9441 (N_9441,N_8965,N_8945);
and U9442 (N_9442,N_8988,N_8724);
and U9443 (N_9443,N_8739,N_8961);
nor U9444 (N_9444,N_8654,N_8633);
nor U9445 (N_9445,N_8756,N_8758);
nand U9446 (N_9446,N_8571,N_8851);
and U9447 (N_9447,N_8784,N_8820);
nand U9448 (N_9448,N_8878,N_8899);
and U9449 (N_9449,N_8515,N_8507);
and U9450 (N_9450,N_8971,N_8662);
or U9451 (N_9451,N_8671,N_8742);
nor U9452 (N_9452,N_8960,N_8966);
xnor U9453 (N_9453,N_8673,N_8957);
or U9454 (N_9454,N_8548,N_8527);
nand U9455 (N_9455,N_8554,N_8661);
or U9456 (N_9456,N_8665,N_8581);
nor U9457 (N_9457,N_8781,N_8987);
nor U9458 (N_9458,N_8795,N_8609);
nand U9459 (N_9459,N_8707,N_8743);
nor U9460 (N_9460,N_8871,N_8794);
nand U9461 (N_9461,N_8545,N_8888);
and U9462 (N_9462,N_8548,N_8811);
or U9463 (N_9463,N_8537,N_8846);
nor U9464 (N_9464,N_8990,N_8750);
nor U9465 (N_9465,N_8812,N_8694);
xnor U9466 (N_9466,N_8965,N_8724);
or U9467 (N_9467,N_8728,N_8566);
nand U9468 (N_9468,N_8566,N_8713);
nand U9469 (N_9469,N_8633,N_8506);
nor U9470 (N_9470,N_8512,N_8672);
and U9471 (N_9471,N_8919,N_8586);
and U9472 (N_9472,N_8923,N_8887);
nor U9473 (N_9473,N_8907,N_8793);
nor U9474 (N_9474,N_8930,N_8996);
nand U9475 (N_9475,N_8632,N_8883);
or U9476 (N_9476,N_8616,N_8853);
xor U9477 (N_9477,N_8869,N_8693);
xor U9478 (N_9478,N_8772,N_8840);
or U9479 (N_9479,N_8640,N_8639);
nor U9480 (N_9480,N_8835,N_8842);
nand U9481 (N_9481,N_8763,N_8657);
and U9482 (N_9482,N_8626,N_8523);
nor U9483 (N_9483,N_8526,N_8894);
nand U9484 (N_9484,N_8733,N_8763);
nand U9485 (N_9485,N_8770,N_8644);
nor U9486 (N_9486,N_8969,N_8636);
or U9487 (N_9487,N_8546,N_8547);
nor U9488 (N_9488,N_8515,N_8724);
nand U9489 (N_9489,N_8848,N_8727);
nor U9490 (N_9490,N_8981,N_8740);
and U9491 (N_9491,N_8516,N_8616);
nand U9492 (N_9492,N_8945,N_8596);
or U9493 (N_9493,N_8982,N_8720);
and U9494 (N_9494,N_8707,N_8888);
or U9495 (N_9495,N_8975,N_8503);
xnor U9496 (N_9496,N_8640,N_8586);
nand U9497 (N_9497,N_8919,N_8734);
or U9498 (N_9498,N_8922,N_8930);
and U9499 (N_9499,N_8511,N_8834);
and U9500 (N_9500,N_9068,N_9080);
or U9501 (N_9501,N_9369,N_9421);
and U9502 (N_9502,N_9201,N_9133);
or U9503 (N_9503,N_9339,N_9124);
or U9504 (N_9504,N_9443,N_9135);
and U9505 (N_9505,N_9405,N_9377);
or U9506 (N_9506,N_9086,N_9458);
and U9507 (N_9507,N_9448,N_9009);
and U9508 (N_9508,N_9276,N_9208);
nor U9509 (N_9509,N_9439,N_9084);
or U9510 (N_9510,N_9202,N_9365);
nand U9511 (N_9511,N_9088,N_9354);
xor U9512 (N_9512,N_9310,N_9416);
and U9513 (N_9513,N_9232,N_9452);
nor U9514 (N_9514,N_9332,N_9285);
nor U9515 (N_9515,N_9375,N_9497);
or U9516 (N_9516,N_9152,N_9122);
or U9517 (N_9517,N_9357,N_9238);
and U9518 (N_9518,N_9060,N_9438);
nand U9519 (N_9519,N_9412,N_9062);
xor U9520 (N_9520,N_9033,N_9266);
and U9521 (N_9521,N_9191,N_9142);
and U9522 (N_9522,N_9363,N_9250);
nor U9523 (N_9523,N_9102,N_9000);
or U9524 (N_9524,N_9333,N_9157);
nor U9525 (N_9525,N_9338,N_9057);
and U9526 (N_9526,N_9098,N_9308);
and U9527 (N_9527,N_9259,N_9200);
nand U9528 (N_9528,N_9241,N_9413);
or U9529 (N_9529,N_9240,N_9064);
and U9530 (N_9530,N_9367,N_9233);
nor U9531 (N_9531,N_9069,N_9175);
or U9532 (N_9532,N_9464,N_9454);
nand U9533 (N_9533,N_9059,N_9261);
and U9534 (N_9534,N_9426,N_9305);
or U9535 (N_9535,N_9028,N_9156);
or U9536 (N_9536,N_9113,N_9126);
or U9537 (N_9537,N_9170,N_9058);
nand U9538 (N_9538,N_9239,N_9029);
or U9539 (N_9539,N_9007,N_9445);
xnor U9540 (N_9540,N_9321,N_9316);
and U9541 (N_9541,N_9211,N_9195);
xor U9542 (N_9542,N_9118,N_9281);
nor U9543 (N_9543,N_9169,N_9273);
or U9544 (N_9544,N_9297,N_9143);
nor U9545 (N_9545,N_9341,N_9262);
or U9546 (N_9546,N_9117,N_9418);
nor U9547 (N_9547,N_9301,N_9465);
or U9548 (N_9548,N_9335,N_9155);
nor U9549 (N_9549,N_9425,N_9392);
nand U9550 (N_9550,N_9138,N_9132);
nand U9551 (N_9551,N_9032,N_9309);
and U9552 (N_9552,N_9486,N_9198);
nand U9553 (N_9553,N_9119,N_9437);
nand U9554 (N_9554,N_9427,N_9213);
and U9555 (N_9555,N_9353,N_9291);
or U9556 (N_9556,N_9167,N_9163);
and U9557 (N_9557,N_9356,N_9456);
or U9558 (N_9558,N_9026,N_9401);
nand U9559 (N_9559,N_9227,N_9078);
and U9560 (N_9560,N_9391,N_9130);
xnor U9561 (N_9561,N_9216,N_9121);
nor U9562 (N_9562,N_9073,N_9337);
nor U9563 (N_9563,N_9303,N_9011);
or U9564 (N_9564,N_9403,N_9090);
and U9565 (N_9565,N_9035,N_9151);
or U9566 (N_9566,N_9292,N_9436);
nand U9567 (N_9567,N_9450,N_9067);
nor U9568 (N_9568,N_9055,N_9433);
xor U9569 (N_9569,N_9346,N_9076);
and U9570 (N_9570,N_9269,N_9455);
and U9571 (N_9571,N_9477,N_9329);
xnor U9572 (N_9572,N_9253,N_9257);
nand U9573 (N_9573,N_9234,N_9236);
and U9574 (N_9574,N_9432,N_9225);
nand U9575 (N_9575,N_9300,N_9052);
and U9576 (N_9576,N_9063,N_9039);
or U9577 (N_9577,N_9129,N_9014);
nor U9578 (N_9578,N_9174,N_9484);
nor U9579 (N_9579,N_9447,N_9476);
and U9580 (N_9580,N_9277,N_9435);
and U9581 (N_9581,N_9214,N_9485);
and U9582 (N_9582,N_9429,N_9251);
nor U9583 (N_9583,N_9043,N_9324);
nand U9584 (N_9584,N_9255,N_9231);
nand U9585 (N_9585,N_9364,N_9323);
nor U9586 (N_9586,N_9244,N_9106);
and U9587 (N_9587,N_9220,N_9137);
and U9588 (N_9588,N_9087,N_9171);
or U9589 (N_9589,N_9289,N_9469);
nor U9590 (N_9590,N_9013,N_9495);
nand U9591 (N_9591,N_9298,N_9263);
and U9592 (N_9592,N_9109,N_9468);
and U9593 (N_9593,N_9472,N_9001);
xor U9594 (N_9594,N_9243,N_9114);
or U9595 (N_9595,N_9348,N_9389);
nand U9596 (N_9596,N_9399,N_9336);
and U9597 (N_9597,N_9409,N_9457);
or U9598 (N_9598,N_9038,N_9228);
and U9599 (N_9599,N_9187,N_9051);
or U9600 (N_9600,N_9177,N_9031);
xor U9601 (N_9601,N_9049,N_9320);
and U9602 (N_9602,N_9047,N_9085);
or U9603 (N_9603,N_9265,N_9154);
and U9604 (N_9604,N_9226,N_9473);
and U9605 (N_9605,N_9428,N_9207);
nand U9606 (N_9606,N_9217,N_9451);
or U9607 (N_9607,N_9070,N_9270);
and U9608 (N_9608,N_9296,N_9224);
and U9609 (N_9609,N_9145,N_9294);
and U9610 (N_9610,N_9105,N_9077);
nor U9611 (N_9611,N_9306,N_9467);
or U9612 (N_9612,N_9140,N_9150);
nand U9613 (N_9613,N_9284,N_9107);
nor U9614 (N_9614,N_9044,N_9302);
xnor U9615 (N_9615,N_9490,N_9350);
nand U9616 (N_9616,N_9164,N_9286);
or U9617 (N_9617,N_9111,N_9131);
and U9618 (N_9618,N_9494,N_9005);
and U9619 (N_9619,N_9134,N_9488);
or U9620 (N_9620,N_9349,N_9311);
nand U9621 (N_9621,N_9023,N_9071);
or U9622 (N_9622,N_9215,N_9492);
and U9623 (N_9623,N_9373,N_9441);
and U9624 (N_9624,N_9016,N_9319);
nand U9625 (N_9625,N_9293,N_9081);
and U9626 (N_9626,N_9393,N_9384);
or U9627 (N_9627,N_9158,N_9181);
and U9628 (N_9628,N_9082,N_9361);
nor U9629 (N_9629,N_9006,N_9021);
nor U9630 (N_9630,N_9371,N_9020);
nand U9631 (N_9631,N_9209,N_9193);
xnor U9632 (N_9632,N_9120,N_9288);
and U9633 (N_9633,N_9172,N_9342);
nand U9634 (N_9634,N_9101,N_9498);
or U9635 (N_9635,N_9414,N_9372);
nor U9636 (N_9636,N_9463,N_9094);
or U9637 (N_9637,N_9493,N_9304);
or U9638 (N_9638,N_9218,N_9491);
nor U9639 (N_9639,N_9274,N_9325);
or U9640 (N_9640,N_9173,N_9290);
nand U9641 (N_9641,N_9061,N_9344);
nand U9642 (N_9642,N_9318,N_9024);
nand U9643 (N_9643,N_9420,N_9358);
nand U9644 (N_9644,N_9017,N_9326);
xnor U9645 (N_9645,N_9222,N_9093);
nand U9646 (N_9646,N_9260,N_9431);
nand U9647 (N_9647,N_9278,N_9002);
nor U9648 (N_9648,N_9166,N_9127);
or U9649 (N_9649,N_9355,N_9136);
nand U9650 (N_9650,N_9203,N_9092);
and U9651 (N_9651,N_9280,N_9025);
or U9652 (N_9652,N_9386,N_9015);
or U9653 (N_9653,N_9307,N_9366);
nand U9654 (N_9654,N_9089,N_9475);
nor U9655 (N_9655,N_9499,N_9442);
xnor U9656 (N_9656,N_9190,N_9470);
nand U9657 (N_9657,N_9381,N_9205);
xor U9658 (N_9658,N_9390,N_9496);
nand U9659 (N_9659,N_9034,N_9100);
nand U9660 (N_9660,N_9045,N_9322);
and U9661 (N_9661,N_9219,N_9159);
nor U9662 (N_9662,N_9248,N_9148);
xor U9663 (N_9663,N_9430,N_9036);
nor U9664 (N_9664,N_9185,N_9128);
and U9665 (N_9665,N_9141,N_9419);
xor U9666 (N_9666,N_9400,N_9115);
and U9667 (N_9667,N_9197,N_9249);
nor U9668 (N_9668,N_9192,N_9388);
and U9669 (N_9669,N_9110,N_9327);
nor U9670 (N_9670,N_9398,N_9144);
and U9671 (N_9671,N_9378,N_9396);
nand U9672 (N_9672,N_9206,N_9165);
nor U9673 (N_9673,N_9066,N_9050);
xnor U9674 (N_9674,N_9314,N_9153);
or U9675 (N_9675,N_9010,N_9275);
or U9676 (N_9676,N_9008,N_9315);
and U9677 (N_9677,N_9230,N_9407);
and U9678 (N_9678,N_9099,N_9083);
nand U9679 (N_9679,N_9478,N_9379);
and U9680 (N_9680,N_9459,N_9108);
and U9681 (N_9681,N_9053,N_9188);
nand U9682 (N_9682,N_9168,N_9487);
nor U9683 (N_9683,N_9423,N_9097);
nand U9684 (N_9684,N_9112,N_9360);
and U9685 (N_9685,N_9056,N_9370);
or U9686 (N_9686,N_9210,N_9256);
or U9687 (N_9687,N_9264,N_9387);
xor U9688 (N_9688,N_9074,N_9212);
nand U9689 (N_9689,N_9096,N_9247);
nor U9690 (N_9690,N_9408,N_9162);
and U9691 (N_9691,N_9397,N_9415);
nand U9692 (N_9692,N_9054,N_9404);
and U9693 (N_9693,N_9482,N_9242);
nand U9694 (N_9694,N_9385,N_9125);
nand U9695 (N_9695,N_9196,N_9410);
nand U9696 (N_9696,N_9254,N_9139);
nor U9697 (N_9697,N_9347,N_9368);
or U9698 (N_9698,N_9022,N_9189);
nand U9699 (N_9699,N_9480,N_9453);
and U9700 (N_9700,N_9313,N_9194);
nand U9701 (N_9701,N_9411,N_9246);
or U9702 (N_9702,N_9283,N_9279);
or U9703 (N_9703,N_9434,N_9359);
or U9704 (N_9704,N_9103,N_9018);
and U9705 (N_9705,N_9382,N_9072);
nand U9706 (N_9706,N_9328,N_9079);
and U9707 (N_9707,N_9027,N_9221);
nand U9708 (N_9708,N_9252,N_9229);
or U9709 (N_9709,N_9440,N_9180);
nand U9710 (N_9710,N_9040,N_9489);
or U9711 (N_9711,N_9394,N_9042);
and U9712 (N_9712,N_9182,N_9104);
nand U9713 (N_9713,N_9204,N_9317);
nand U9714 (N_9714,N_9037,N_9267);
nor U9715 (N_9715,N_9012,N_9395);
and U9716 (N_9716,N_9186,N_9374);
nor U9717 (N_9717,N_9046,N_9483);
nor U9718 (N_9718,N_9479,N_9004);
or U9719 (N_9719,N_9380,N_9331);
and U9720 (N_9720,N_9449,N_9048);
xor U9721 (N_9721,N_9065,N_9424);
nor U9722 (N_9722,N_9149,N_9160);
or U9723 (N_9723,N_9030,N_9237);
nor U9724 (N_9724,N_9147,N_9406);
and U9725 (N_9725,N_9075,N_9268);
and U9726 (N_9726,N_9299,N_9176);
and U9727 (N_9727,N_9460,N_9199);
nor U9728 (N_9728,N_9041,N_9466);
and U9729 (N_9729,N_9287,N_9446);
and U9730 (N_9730,N_9183,N_9146);
or U9731 (N_9731,N_9462,N_9019);
xnor U9732 (N_9732,N_9295,N_9481);
and U9733 (N_9733,N_9417,N_9362);
or U9734 (N_9734,N_9312,N_9271);
or U9735 (N_9735,N_9471,N_9123);
nor U9736 (N_9736,N_9422,N_9178);
xor U9737 (N_9737,N_9091,N_9343);
nand U9738 (N_9738,N_9245,N_9258);
or U9739 (N_9739,N_9474,N_9272);
or U9740 (N_9740,N_9402,N_9351);
and U9741 (N_9741,N_9282,N_9116);
or U9742 (N_9742,N_9179,N_9376);
nor U9743 (N_9743,N_9223,N_9330);
nor U9744 (N_9744,N_9184,N_9340);
nor U9745 (N_9745,N_9461,N_9383);
nor U9746 (N_9746,N_9161,N_9095);
nand U9747 (N_9747,N_9003,N_9444);
xor U9748 (N_9748,N_9334,N_9345);
nand U9749 (N_9749,N_9235,N_9352);
xnor U9750 (N_9750,N_9391,N_9003);
xor U9751 (N_9751,N_9099,N_9440);
or U9752 (N_9752,N_9225,N_9401);
or U9753 (N_9753,N_9223,N_9030);
and U9754 (N_9754,N_9488,N_9171);
and U9755 (N_9755,N_9008,N_9088);
nand U9756 (N_9756,N_9120,N_9166);
nor U9757 (N_9757,N_9333,N_9080);
nor U9758 (N_9758,N_9212,N_9154);
or U9759 (N_9759,N_9098,N_9469);
nand U9760 (N_9760,N_9164,N_9180);
nor U9761 (N_9761,N_9115,N_9163);
nand U9762 (N_9762,N_9075,N_9388);
or U9763 (N_9763,N_9297,N_9411);
or U9764 (N_9764,N_9499,N_9133);
nor U9765 (N_9765,N_9390,N_9075);
nor U9766 (N_9766,N_9137,N_9131);
nand U9767 (N_9767,N_9317,N_9159);
or U9768 (N_9768,N_9229,N_9149);
and U9769 (N_9769,N_9439,N_9350);
nor U9770 (N_9770,N_9063,N_9379);
xnor U9771 (N_9771,N_9448,N_9270);
nand U9772 (N_9772,N_9466,N_9090);
nand U9773 (N_9773,N_9464,N_9144);
and U9774 (N_9774,N_9344,N_9430);
or U9775 (N_9775,N_9052,N_9368);
and U9776 (N_9776,N_9459,N_9498);
nor U9777 (N_9777,N_9227,N_9203);
nand U9778 (N_9778,N_9233,N_9234);
xor U9779 (N_9779,N_9439,N_9200);
or U9780 (N_9780,N_9486,N_9120);
xor U9781 (N_9781,N_9144,N_9037);
or U9782 (N_9782,N_9328,N_9065);
nor U9783 (N_9783,N_9314,N_9178);
nand U9784 (N_9784,N_9147,N_9489);
nand U9785 (N_9785,N_9472,N_9303);
and U9786 (N_9786,N_9410,N_9359);
nand U9787 (N_9787,N_9183,N_9127);
nor U9788 (N_9788,N_9056,N_9482);
and U9789 (N_9789,N_9070,N_9038);
nand U9790 (N_9790,N_9034,N_9047);
and U9791 (N_9791,N_9055,N_9326);
and U9792 (N_9792,N_9431,N_9127);
nor U9793 (N_9793,N_9356,N_9173);
nand U9794 (N_9794,N_9353,N_9203);
or U9795 (N_9795,N_9029,N_9155);
or U9796 (N_9796,N_9162,N_9131);
nand U9797 (N_9797,N_9336,N_9105);
nor U9798 (N_9798,N_9181,N_9062);
nand U9799 (N_9799,N_9271,N_9089);
nand U9800 (N_9800,N_9273,N_9393);
nand U9801 (N_9801,N_9184,N_9348);
xor U9802 (N_9802,N_9131,N_9119);
nand U9803 (N_9803,N_9052,N_9167);
nor U9804 (N_9804,N_9404,N_9439);
and U9805 (N_9805,N_9040,N_9246);
and U9806 (N_9806,N_9361,N_9310);
nor U9807 (N_9807,N_9204,N_9156);
or U9808 (N_9808,N_9227,N_9158);
and U9809 (N_9809,N_9267,N_9237);
and U9810 (N_9810,N_9097,N_9284);
and U9811 (N_9811,N_9289,N_9258);
nand U9812 (N_9812,N_9349,N_9327);
or U9813 (N_9813,N_9192,N_9392);
nor U9814 (N_9814,N_9373,N_9353);
nor U9815 (N_9815,N_9364,N_9053);
or U9816 (N_9816,N_9183,N_9035);
and U9817 (N_9817,N_9466,N_9447);
nor U9818 (N_9818,N_9034,N_9397);
nor U9819 (N_9819,N_9109,N_9228);
xor U9820 (N_9820,N_9191,N_9447);
nand U9821 (N_9821,N_9331,N_9354);
xnor U9822 (N_9822,N_9432,N_9205);
or U9823 (N_9823,N_9065,N_9186);
nand U9824 (N_9824,N_9383,N_9054);
or U9825 (N_9825,N_9360,N_9446);
and U9826 (N_9826,N_9057,N_9104);
nor U9827 (N_9827,N_9220,N_9287);
and U9828 (N_9828,N_9427,N_9058);
xnor U9829 (N_9829,N_9400,N_9182);
or U9830 (N_9830,N_9300,N_9361);
or U9831 (N_9831,N_9041,N_9396);
nor U9832 (N_9832,N_9043,N_9497);
nor U9833 (N_9833,N_9344,N_9305);
and U9834 (N_9834,N_9178,N_9432);
nand U9835 (N_9835,N_9204,N_9160);
xor U9836 (N_9836,N_9214,N_9029);
or U9837 (N_9837,N_9347,N_9082);
nor U9838 (N_9838,N_9044,N_9179);
nand U9839 (N_9839,N_9160,N_9255);
or U9840 (N_9840,N_9429,N_9417);
and U9841 (N_9841,N_9280,N_9358);
nand U9842 (N_9842,N_9344,N_9423);
nand U9843 (N_9843,N_9414,N_9355);
or U9844 (N_9844,N_9041,N_9245);
xnor U9845 (N_9845,N_9216,N_9395);
and U9846 (N_9846,N_9400,N_9343);
or U9847 (N_9847,N_9474,N_9112);
nand U9848 (N_9848,N_9361,N_9259);
nand U9849 (N_9849,N_9080,N_9447);
nor U9850 (N_9850,N_9153,N_9246);
or U9851 (N_9851,N_9493,N_9341);
nand U9852 (N_9852,N_9052,N_9341);
nor U9853 (N_9853,N_9092,N_9444);
nand U9854 (N_9854,N_9092,N_9452);
xor U9855 (N_9855,N_9082,N_9151);
nor U9856 (N_9856,N_9063,N_9265);
and U9857 (N_9857,N_9274,N_9267);
or U9858 (N_9858,N_9336,N_9473);
and U9859 (N_9859,N_9262,N_9426);
or U9860 (N_9860,N_9409,N_9317);
nor U9861 (N_9861,N_9274,N_9112);
nand U9862 (N_9862,N_9468,N_9316);
and U9863 (N_9863,N_9251,N_9471);
or U9864 (N_9864,N_9475,N_9034);
or U9865 (N_9865,N_9359,N_9383);
or U9866 (N_9866,N_9316,N_9152);
and U9867 (N_9867,N_9401,N_9446);
xnor U9868 (N_9868,N_9185,N_9254);
or U9869 (N_9869,N_9477,N_9230);
or U9870 (N_9870,N_9162,N_9100);
xnor U9871 (N_9871,N_9252,N_9065);
nand U9872 (N_9872,N_9475,N_9105);
or U9873 (N_9873,N_9167,N_9204);
nand U9874 (N_9874,N_9260,N_9479);
nand U9875 (N_9875,N_9304,N_9496);
nor U9876 (N_9876,N_9391,N_9366);
nand U9877 (N_9877,N_9476,N_9317);
nor U9878 (N_9878,N_9386,N_9372);
nor U9879 (N_9879,N_9031,N_9200);
nor U9880 (N_9880,N_9246,N_9293);
or U9881 (N_9881,N_9032,N_9124);
and U9882 (N_9882,N_9217,N_9166);
nand U9883 (N_9883,N_9037,N_9167);
and U9884 (N_9884,N_9135,N_9398);
nand U9885 (N_9885,N_9109,N_9415);
or U9886 (N_9886,N_9125,N_9182);
and U9887 (N_9887,N_9435,N_9250);
nand U9888 (N_9888,N_9151,N_9099);
nand U9889 (N_9889,N_9486,N_9091);
and U9890 (N_9890,N_9320,N_9074);
xor U9891 (N_9891,N_9237,N_9165);
and U9892 (N_9892,N_9325,N_9405);
or U9893 (N_9893,N_9480,N_9422);
nor U9894 (N_9894,N_9122,N_9427);
or U9895 (N_9895,N_9216,N_9495);
nor U9896 (N_9896,N_9201,N_9456);
and U9897 (N_9897,N_9435,N_9020);
or U9898 (N_9898,N_9150,N_9388);
and U9899 (N_9899,N_9001,N_9325);
nor U9900 (N_9900,N_9366,N_9394);
xnor U9901 (N_9901,N_9158,N_9230);
or U9902 (N_9902,N_9418,N_9381);
or U9903 (N_9903,N_9356,N_9405);
nand U9904 (N_9904,N_9201,N_9415);
nor U9905 (N_9905,N_9182,N_9229);
nand U9906 (N_9906,N_9191,N_9372);
nand U9907 (N_9907,N_9438,N_9074);
or U9908 (N_9908,N_9436,N_9414);
nand U9909 (N_9909,N_9451,N_9320);
or U9910 (N_9910,N_9325,N_9314);
xor U9911 (N_9911,N_9151,N_9031);
nand U9912 (N_9912,N_9009,N_9252);
nor U9913 (N_9913,N_9373,N_9150);
and U9914 (N_9914,N_9083,N_9076);
and U9915 (N_9915,N_9021,N_9387);
nand U9916 (N_9916,N_9136,N_9216);
nand U9917 (N_9917,N_9377,N_9242);
nand U9918 (N_9918,N_9099,N_9297);
nor U9919 (N_9919,N_9318,N_9157);
nand U9920 (N_9920,N_9322,N_9027);
and U9921 (N_9921,N_9179,N_9193);
xor U9922 (N_9922,N_9045,N_9003);
or U9923 (N_9923,N_9399,N_9237);
or U9924 (N_9924,N_9464,N_9078);
nor U9925 (N_9925,N_9187,N_9431);
nand U9926 (N_9926,N_9367,N_9281);
xor U9927 (N_9927,N_9304,N_9355);
xor U9928 (N_9928,N_9111,N_9312);
nor U9929 (N_9929,N_9026,N_9480);
nand U9930 (N_9930,N_9135,N_9234);
nor U9931 (N_9931,N_9106,N_9484);
nor U9932 (N_9932,N_9181,N_9239);
and U9933 (N_9933,N_9120,N_9454);
xor U9934 (N_9934,N_9195,N_9053);
nand U9935 (N_9935,N_9143,N_9127);
nor U9936 (N_9936,N_9138,N_9354);
nor U9937 (N_9937,N_9254,N_9289);
nor U9938 (N_9938,N_9402,N_9083);
xnor U9939 (N_9939,N_9014,N_9125);
or U9940 (N_9940,N_9358,N_9011);
xor U9941 (N_9941,N_9035,N_9228);
nand U9942 (N_9942,N_9007,N_9137);
nand U9943 (N_9943,N_9344,N_9002);
or U9944 (N_9944,N_9237,N_9210);
or U9945 (N_9945,N_9424,N_9092);
or U9946 (N_9946,N_9309,N_9391);
and U9947 (N_9947,N_9313,N_9007);
nand U9948 (N_9948,N_9053,N_9175);
or U9949 (N_9949,N_9057,N_9117);
xnor U9950 (N_9950,N_9313,N_9151);
nor U9951 (N_9951,N_9310,N_9422);
xnor U9952 (N_9952,N_9207,N_9028);
nand U9953 (N_9953,N_9002,N_9289);
xor U9954 (N_9954,N_9047,N_9334);
nor U9955 (N_9955,N_9336,N_9270);
nor U9956 (N_9956,N_9116,N_9349);
nor U9957 (N_9957,N_9045,N_9338);
xnor U9958 (N_9958,N_9053,N_9205);
or U9959 (N_9959,N_9404,N_9419);
nand U9960 (N_9960,N_9446,N_9349);
and U9961 (N_9961,N_9211,N_9385);
nand U9962 (N_9962,N_9112,N_9447);
nor U9963 (N_9963,N_9188,N_9349);
nor U9964 (N_9964,N_9393,N_9058);
and U9965 (N_9965,N_9293,N_9257);
nor U9966 (N_9966,N_9257,N_9381);
xor U9967 (N_9967,N_9252,N_9131);
nor U9968 (N_9968,N_9123,N_9336);
nor U9969 (N_9969,N_9373,N_9310);
nor U9970 (N_9970,N_9446,N_9475);
and U9971 (N_9971,N_9423,N_9365);
and U9972 (N_9972,N_9346,N_9211);
and U9973 (N_9973,N_9303,N_9323);
xnor U9974 (N_9974,N_9078,N_9158);
nand U9975 (N_9975,N_9411,N_9425);
and U9976 (N_9976,N_9325,N_9071);
nand U9977 (N_9977,N_9283,N_9374);
nand U9978 (N_9978,N_9172,N_9424);
nor U9979 (N_9979,N_9230,N_9269);
or U9980 (N_9980,N_9379,N_9216);
nand U9981 (N_9981,N_9373,N_9276);
nor U9982 (N_9982,N_9472,N_9479);
nor U9983 (N_9983,N_9256,N_9460);
or U9984 (N_9984,N_9043,N_9051);
or U9985 (N_9985,N_9344,N_9131);
or U9986 (N_9986,N_9223,N_9375);
or U9987 (N_9987,N_9188,N_9432);
and U9988 (N_9988,N_9404,N_9122);
and U9989 (N_9989,N_9179,N_9237);
nand U9990 (N_9990,N_9027,N_9014);
and U9991 (N_9991,N_9454,N_9099);
xor U9992 (N_9992,N_9474,N_9035);
and U9993 (N_9993,N_9005,N_9249);
nor U9994 (N_9994,N_9363,N_9496);
or U9995 (N_9995,N_9369,N_9198);
or U9996 (N_9996,N_9262,N_9176);
xnor U9997 (N_9997,N_9322,N_9413);
or U9998 (N_9998,N_9030,N_9089);
nor U9999 (N_9999,N_9222,N_9228);
or U10000 (N_10000,N_9690,N_9940);
nor U10001 (N_10001,N_9779,N_9966);
nand U10002 (N_10002,N_9506,N_9783);
nor U10003 (N_10003,N_9730,N_9986);
and U10004 (N_10004,N_9558,N_9835);
nor U10005 (N_10005,N_9815,N_9525);
nand U10006 (N_10006,N_9845,N_9792);
xor U10007 (N_10007,N_9703,N_9891);
nor U10008 (N_10008,N_9914,N_9911);
or U10009 (N_10009,N_9941,N_9546);
or U10010 (N_10010,N_9677,N_9538);
or U10011 (N_10011,N_9960,N_9515);
nor U10012 (N_10012,N_9858,N_9823);
xnor U10013 (N_10013,N_9624,N_9809);
or U10014 (N_10014,N_9755,N_9844);
nand U10015 (N_10015,N_9692,N_9832);
or U10016 (N_10016,N_9642,N_9671);
or U10017 (N_10017,N_9606,N_9925);
nor U10018 (N_10018,N_9859,N_9965);
nor U10019 (N_10019,N_9764,N_9843);
nand U10020 (N_10020,N_9898,N_9904);
nor U10021 (N_10021,N_9635,N_9666);
and U10022 (N_10022,N_9681,N_9957);
nand U10023 (N_10023,N_9753,N_9884);
and U10024 (N_10024,N_9534,N_9837);
and U10025 (N_10025,N_9789,N_9926);
nand U10026 (N_10026,N_9808,N_9722);
and U10027 (N_10027,N_9601,N_9948);
or U10028 (N_10028,N_9969,N_9587);
or U10029 (N_10029,N_9527,N_9613);
and U10030 (N_10030,N_9972,N_9933);
and U10031 (N_10031,N_9656,N_9597);
nor U10032 (N_10032,N_9710,N_9669);
nand U10033 (N_10033,N_9502,N_9906);
and U10034 (N_10034,N_9636,N_9605);
nand U10035 (N_10035,N_9556,N_9791);
nand U10036 (N_10036,N_9505,N_9923);
xor U10037 (N_10037,N_9640,N_9673);
nand U10038 (N_10038,N_9894,N_9707);
nor U10039 (N_10039,N_9616,N_9820);
nand U10040 (N_10040,N_9953,N_9594);
nor U10041 (N_10041,N_9934,N_9975);
nand U10042 (N_10042,N_9641,N_9874);
or U10043 (N_10043,N_9596,N_9973);
or U10044 (N_10044,N_9734,N_9617);
nand U10045 (N_10045,N_9687,N_9741);
nor U10046 (N_10046,N_9967,N_9510);
or U10047 (N_10047,N_9801,N_9622);
or U10048 (N_10048,N_9876,N_9739);
nand U10049 (N_10049,N_9705,N_9840);
nand U10050 (N_10050,N_9829,N_9757);
nand U10051 (N_10051,N_9699,N_9989);
nand U10052 (N_10052,N_9849,N_9970);
and U10053 (N_10053,N_9559,N_9821);
nand U10054 (N_10054,N_9649,N_9545);
nand U10055 (N_10055,N_9522,N_9626);
nor U10056 (N_10056,N_9991,N_9610);
xor U10057 (N_10057,N_9883,N_9943);
or U10058 (N_10058,N_9851,N_9961);
and U10059 (N_10059,N_9760,N_9544);
xor U10060 (N_10060,N_9786,N_9831);
or U10061 (N_10061,N_9763,N_9766);
nor U10062 (N_10062,N_9698,N_9803);
nor U10063 (N_10063,N_9680,N_9930);
or U10064 (N_10064,N_9650,N_9879);
or U10065 (N_10065,N_9566,N_9547);
nand U10066 (N_10066,N_9675,N_9910);
nor U10067 (N_10067,N_9903,N_9977);
nor U10068 (N_10068,N_9543,N_9530);
and U10069 (N_10069,N_9573,N_9578);
xnor U10070 (N_10070,N_9674,N_9773);
or U10071 (N_10071,N_9564,N_9682);
and U10072 (N_10072,N_9810,N_9598);
and U10073 (N_10073,N_9592,N_9694);
and U10074 (N_10074,N_9908,N_9655);
nand U10075 (N_10075,N_9591,N_9688);
xnor U10076 (N_10076,N_9775,N_9647);
or U10077 (N_10077,N_9890,N_9733);
and U10078 (N_10078,N_9738,N_9954);
nor U10079 (N_10079,N_9942,N_9672);
or U10080 (N_10080,N_9959,N_9863);
or U10081 (N_10081,N_9920,N_9634);
nor U10082 (N_10082,N_9718,N_9800);
nand U10083 (N_10083,N_9939,N_9731);
xor U10084 (N_10084,N_9643,N_9981);
nand U10085 (N_10085,N_9878,N_9870);
and U10086 (N_10086,N_9768,N_9631);
xor U10087 (N_10087,N_9569,N_9900);
and U10088 (N_10088,N_9551,N_9735);
nand U10089 (N_10089,N_9621,N_9772);
or U10090 (N_10090,N_9528,N_9976);
nor U10091 (N_10091,N_9913,N_9781);
and U10092 (N_10092,N_9728,N_9770);
nand U10093 (N_10093,N_9865,N_9664);
nor U10094 (N_10094,N_9974,N_9581);
nand U10095 (N_10095,N_9927,N_9813);
nor U10096 (N_10096,N_9955,N_9882);
and U10097 (N_10097,N_9589,N_9833);
or U10098 (N_10098,N_9552,N_9590);
and U10099 (N_10099,N_9549,N_9526);
or U10100 (N_10100,N_9509,N_9996);
xor U10101 (N_10101,N_9535,N_9542);
nor U10102 (N_10102,N_9866,N_9574);
xor U10103 (N_10103,N_9603,N_9872);
or U10104 (N_10104,N_9995,N_9839);
xnor U10105 (N_10105,N_9785,N_9554);
or U10106 (N_10106,N_9723,N_9877);
or U10107 (N_10107,N_9593,N_9614);
and U10108 (N_10108,N_9769,N_9689);
nor U10109 (N_10109,N_9612,N_9938);
nand U10110 (N_10110,N_9827,N_9576);
xor U10111 (N_10111,N_9714,N_9517);
nor U10112 (N_10112,N_9998,N_9716);
nor U10113 (N_10113,N_9787,N_9676);
and U10114 (N_10114,N_9794,N_9721);
or U10115 (N_10115,N_9881,N_9897);
or U10116 (N_10116,N_9529,N_9871);
nand U10117 (N_10117,N_9790,N_9956);
nor U10118 (N_10118,N_9946,N_9979);
nor U10119 (N_10119,N_9888,N_9711);
or U10120 (N_10120,N_9817,N_9696);
or U10121 (N_10121,N_9715,N_9873);
and U10122 (N_10122,N_9652,N_9765);
or U10123 (N_10123,N_9570,N_9788);
nand U10124 (N_10124,N_9701,N_9988);
nor U10125 (N_10125,N_9548,N_9653);
and U10126 (N_10126,N_9774,N_9567);
or U10127 (N_10127,N_9932,N_9987);
or U10128 (N_10128,N_9609,N_9747);
and U10129 (N_10129,N_9695,N_9795);
nor U10130 (N_10130,N_9654,N_9828);
nand U10131 (N_10131,N_9516,N_9958);
and U10132 (N_10132,N_9713,N_9825);
nand U10133 (N_10133,N_9629,N_9582);
xor U10134 (N_10134,N_9615,N_9984);
xnor U10135 (N_10135,N_9646,N_9912);
or U10136 (N_10136,N_9557,N_9706);
nand U10137 (N_10137,N_9964,N_9841);
or U10138 (N_10138,N_9563,N_9637);
nor U10139 (N_10139,N_9751,N_9907);
nor U10140 (N_10140,N_9868,N_9684);
or U10141 (N_10141,N_9892,N_9861);
or U10142 (N_10142,N_9504,N_9919);
or U10143 (N_10143,N_9793,N_9746);
nand U10144 (N_10144,N_9761,N_9905);
nand U10145 (N_10145,N_9999,N_9952);
nand U10146 (N_10146,N_9645,N_9944);
nor U10147 (N_10147,N_9816,N_9748);
xor U10148 (N_10148,N_9565,N_9830);
nand U10149 (N_10149,N_9658,N_9875);
nand U10150 (N_10150,N_9836,N_9571);
nand U10151 (N_10151,N_9651,N_9853);
or U10152 (N_10152,N_9889,N_9778);
and U10153 (N_10153,N_9814,N_9583);
nand U10154 (N_10154,N_9928,N_9886);
xnor U10155 (N_10155,N_9602,N_9804);
or U10156 (N_10156,N_9848,N_9595);
or U10157 (N_10157,N_9802,N_9740);
nand U10158 (N_10158,N_9806,N_9887);
and U10159 (N_10159,N_9686,N_9608);
and U10160 (N_10160,N_9811,N_9968);
and U10161 (N_10161,N_9648,N_9644);
or U10162 (N_10162,N_9500,N_9550);
nor U10163 (N_10163,N_9846,N_9850);
xor U10164 (N_10164,N_9501,N_9693);
nand U10165 (N_10165,N_9727,N_9963);
xor U10166 (N_10166,N_9798,N_9662);
nor U10167 (N_10167,N_9749,N_9860);
and U10168 (N_10168,N_9838,N_9679);
nand U10169 (N_10169,N_9562,N_9579);
xnor U10170 (N_10170,N_9560,N_9541);
and U10171 (N_10171,N_9936,N_9520);
nand U10172 (N_10172,N_9668,N_9799);
or U10173 (N_10173,N_9540,N_9555);
or U10174 (N_10174,N_9607,N_9660);
nand U10175 (N_10175,N_9902,N_9628);
and U10176 (N_10176,N_9797,N_9577);
nor U10177 (N_10177,N_9742,N_9536);
and U10178 (N_10178,N_9737,N_9762);
nor U10179 (N_10179,N_9869,N_9729);
nand U10180 (N_10180,N_9864,N_9750);
nor U10181 (N_10181,N_9657,N_9736);
nor U10182 (N_10182,N_9507,N_9901);
nand U10183 (N_10183,N_9584,N_9604);
or U10184 (N_10184,N_9611,N_9619);
and U10185 (N_10185,N_9661,N_9867);
nand U10186 (N_10186,N_9630,N_9588);
nor U10187 (N_10187,N_9922,N_9899);
and U10188 (N_10188,N_9708,N_9586);
nor U10189 (N_10189,N_9639,N_9776);
or U10190 (N_10190,N_9951,N_9725);
nor U10191 (N_10191,N_9531,N_9719);
nand U10192 (N_10192,N_9519,N_9880);
and U10193 (N_10193,N_9585,N_9937);
or U10194 (N_10194,N_9971,N_9709);
nand U10195 (N_10195,N_9712,N_9771);
nand U10196 (N_10196,N_9514,N_9513);
and U10197 (N_10197,N_9782,N_9777);
nor U10198 (N_10198,N_9659,N_9618);
nand U10199 (N_10199,N_9997,N_9896);
xor U10200 (N_10200,N_9992,N_9818);
nand U10201 (N_10201,N_9678,N_9994);
and U10202 (N_10202,N_9632,N_9599);
or U10203 (N_10203,N_9508,N_9667);
xor U10204 (N_10204,N_9980,N_9511);
or U10205 (N_10205,N_9796,N_9909);
nand U10206 (N_10206,N_9921,N_9726);
or U10207 (N_10207,N_9625,N_9935);
nor U10208 (N_10208,N_9697,N_9924);
and U10209 (N_10209,N_9580,N_9822);
nor U10210 (N_10210,N_9985,N_9756);
nor U10211 (N_10211,N_9600,N_9683);
or U10212 (N_10212,N_9518,N_9854);
nor U10213 (N_10213,N_9724,N_9537);
and U10214 (N_10214,N_9523,N_9950);
xor U10215 (N_10215,N_9539,N_9568);
and U10216 (N_10216,N_9620,N_9572);
and U10217 (N_10217,N_9812,N_9856);
nand U10218 (N_10218,N_9983,N_9752);
nand U10219 (N_10219,N_9524,N_9743);
nand U10220 (N_10220,N_9949,N_9978);
and U10221 (N_10221,N_9745,N_9857);
nor U10222 (N_10222,N_9633,N_9962);
or U10223 (N_10223,N_9754,N_9929);
xor U10224 (N_10224,N_9847,N_9834);
nor U10225 (N_10225,N_9826,N_9931);
nand U10226 (N_10226,N_9758,N_9700);
and U10227 (N_10227,N_9575,N_9532);
or U10228 (N_10228,N_9893,N_9717);
and U10229 (N_10229,N_9885,N_9627);
nand U10230 (N_10230,N_9561,N_9918);
nor U10231 (N_10231,N_9533,N_9807);
nand U10232 (N_10232,N_9691,N_9663);
and U10233 (N_10233,N_9862,N_9759);
and U10234 (N_10234,N_9805,N_9704);
nand U10235 (N_10235,N_9915,N_9993);
nor U10236 (N_10236,N_9685,N_9623);
or U10237 (N_10237,N_9732,N_9702);
nand U10238 (N_10238,N_9767,N_9982);
or U10239 (N_10239,N_9917,N_9842);
nand U10240 (N_10240,N_9945,N_9665);
and U10241 (N_10241,N_9780,N_9990);
or U10242 (N_10242,N_9895,N_9824);
xnor U10243 (N_10243,N_9744,N_9947);
and U10244 (N_10244,N_9855,N_9784);
or U10245 (N_10245,N_9819,N_9503);
xor U10246 (N_10246,N_9553,N_9720);
nor U10247 (N_10247,N_9916,N_9638);
xor U10248 (N_10248,N_9521,N_9852);
or U10249 (N_10249,N_9512,N_9670);
nand U10250 (N_10250,N_9963,N_9917);
and U10251 (N_10251,N_9617,N_9689);
xnor U10252 (N_10252,N_9733,N_9885);
or U10253 (N_10253,N_9861,N_9755);
xnor U10254 (N_10254,N_9761,N_9986);
nand U10255 (N_10255,N_9897,N_9837);
xor U10256 (N_10256,N_9791,N_9917);
and U10257 (N_10257,N_9907,N_9686);
nor U10258 (N_10258,N_9561,N_9807);
nand U10259 (N_10259,N_9800,N_9508);
nand U10260 (N_10260,N_9767,N_9650);
xnor U10261 (N_10261,N_9685,N_9962);
and U10262 (N_10262,N_9738,N_9772);
and U10263 (N_10263,N_9597,N_9548);
nand U10264 (N_10264,N_9910,N_9750);
nand U10265 (N_10265,N_9994,N_9569);
and U10266 (N_10266,N_9745,N_9697);
nand U10267 (N_10267,N_9950,N_9857);
xor U10268 (N_10268,N_9959,N_9711);
nor U10269 (N_10269,N_9804,N_9660);
nor U10270 (N_10270,N_9827,N_9701);
nor U10271 (N_10271,N_9597,N_9650);
xor U10272 (N_10272,N_9814,N_9578);
nand U10273 (N_10273,N_9501,N_9962);
nand U10274 (N_10274,N_9614,N_9717);
and U10275 (N_10275,N_9669,N_9960);
xor U10276 (N_10276,N_9595,N_9669);
or U10277 (N_10277,N_9655,N_9601);
or U10278 (N_10278,N_9885,N_9943);
nor U10279 (N_10279,N_9824,N_9843);
and U10280 (N_10280,N_9986,N_9616);
and U10281 (N_10281,N_9646,N_9851);
nand U10282 (N_10282,N_9573,N_9507);
and U10283 (N_10283,N_9565,N_9732);
or U10284 (N_10284,N_9656,N_9657);
or U10285 (N_10285,N_9723,N_9889);
or U10286 (N_10286,N_9691,N_9561);
xnor U10287 (N_10287,N_9719,N_9575);
and U10288 (N_10288,N_9506,N_9608);
or U10289 (N_10289,N_9645,N_9808);
nand U10290 (N_10290,N_9919,N_9737);
nand U10291 (N_10291,N_9863,N_9704);
and U10292 (N_10292,N_9510,N_9822);
and U10293 (N_10293,N_9897,N_9658);
and U10294 (N_10294,N_9536,N_9914);
or U10295 (N_10295,N_9923,N_9635);
nand U10296 (N_10296,N_9663,N_9563);
and U10297 (N_10297,N_9884,N_9947);
and U10298 (N_10298,N_9785,N_9887);
nand U10299 (N_10299,N_9654,N_9945);
nand U10300 (N_10300,N_9992,N_9641);
and U10301 (N_10301,N_9774,N_9656);
and U10302 (N_10302,N_9939,N_9699);
and U10303 (N_10303,N_9821,N_9599);
xnor U10304 (N_10304,N_9954,N_9911);
nand U10305 (N_10305,N_9762,N_9675);
nand U10306 (N_10306,N_9953,N_9758);
nand U10307 (N_10307,N_9724,N_9808);
and U10308 (N_10308,N_9891,N_9855);
and U10309 (N_10309,N_9857,N_9627);
or U10310 (N_10310,N_9762,N_9629);
and U10311 (N_10311,N_9693,N_9570);
and U10312 (N_10312,N_9510,N_9637);
nor U10313 (N_10313,N_9964,N_9511);
or U10314 (N_10314,N_9719,N_9580);
or U10315 (N_10315,N_9975,N_9712);
or U10316 (N_10316,N_9838,N_9836);
and U10317 (N_10317,N_9971,N_9596);
nand U10318 (N_10318,N_9952,N_9749);
nor U10319 (N_10319,N_9523,N_9734);
nand U10320 (N_10320,N_9626,N_9666);
nand U10321 (N_10321,N_9573,N_9876);
nand U10322 (N_10322,N_9572,N_9918);
nor U10323 (N_10323,N_9641,N_9760);
or U10324 (N_10324,N_9607,N_9640);
xor U10325 (N_10325,N_9911,N_9825);
or U10326 (N_10326,N_9560,N_9854);
and U10327 (N_10327,N_9597,N_9982);
nand U10328 (N_10328,N_9960,N_9546);
xnor U10329 (N_10329,N_9515,N_9902);
or U10330 (N_10330,N_9785,N_9929);
nand U10331 (N_10331,N_9596,N_9681);
nand U10332 (N_10332,N_9771,N_9553);
or U10333 (N_10333,N_9934,N_9558);
nand U10334 (N_10334,N_9953,N_9914);
and U10335 (N_10335,N_9769,N_9703);
xor U10336 (N_10336,N_9630,N_9582);
and U10337 (N_10337,N_9713,N_9519);
nor U10338 (N_10338,N_9560,N_9909);
nand U10339 (N_10339,N_9560,N_9978);
nor U10340 (N_10340,N_9715,N_9503);
nor U10341 (N_10341,N_9891,N_9894);
nand U10342 (N_10342,N_9776,N_9675);
nand U10343 (N_10343,N_9522,N_9974);
and U10344 (N_10344,N_9654,N_9955);
nand U10345 (N_10345,N_9580,N_9884);
and U10346 (N_10346,N_9919,N_9640);
xnor U10347 (N_10347,N_9672,N_9678);
and U10348 (N_10348,N_9564,N_9936);
nor U10349 (N_10349,N_9677,N_9660);
nand U10350 (N_10350,N_9889,N_9747);
nand U10351 (N_10351,N_9695,N_9776);
xor U10352 (N_10352,N_9817,N_9701);
or U10353 (N_10353,N_9917,N_9557);
and U10354 (N_10354,N_9949,N_9895);
and U10355 (N_10355,N_9557,N_9887);
xnor U10356 (N_10356,N_9654,N_9519);
or U10357 (N_10357,N_9676,N_9722);
nand U10358 (N_10358,N_9629,N_9700);
nor U10359 (N_10359,N_9660,N_9609);
or U10360 (N_10360,N_9651,N_9551);
or U10361 (N_10361,N_9725,N_9905);
nand U10362 (N_10362,N_9719,N_9896);
and U10363 (N_10363,N_9955,N_9881);
nor U10364 (N_10364,N_9764,N_9903);
nor U10365 (N_10365,N_9808,N_9531);
or U10366 (N_10366,N_9745,N_9579);
nor U10367 (N_10367,N_9739,N_9511);
nor U10368 (N_10368,N_9836,N_9650);
and U10369 (N_10369,N_9964,N_9692);
nand U10370 (N_10370,N_9872,N_9952);
and U10371 (N_10371,N_9550,N_9512);
or U10372 (N_10372,N_9877,N_9597);
nor U10373 (N_10373,N_9552,N_9583);
or U10374 (N_10374,N_9636,N_9603);
and U10375 (N_10375,N_9921,N_9611);
nor U10376 (N_10376,N_9911,N_9946);
and U10377 (N_10377,N_9719,N_9674);
or U10378 (N_10378,N_9983,N_9645);
and U10379 (N_10379,N_9564,N_9697);
nand U10380 (N_10380,N_9932,N_9548);
or U10381 (N_10381,N_9710,N_9702);
or U10382 (N_10382,N_9967,N_9937);
nand U10383 (N_10383,N_9588,N_9880);
nand U10384 (N_10384,N_9945,N_9756);
and U10385 (N_10385,N_9700,N_9540);
or U10386 (N_10386,N_9657,N_9876);
nor U10387 (N_10387,N_9659,N_9524);
nor U10388 (N_10388,N_9897,N_9933);
and U10389 (N_10389,N_9713,N_9939);
nor U10390 (N_10390,N_9526,N_9733);
nand U10391 (N_10391,N_9838,N_9637);
nor U10392 (N_10392,N_9664,N_9515);
nand U10393 (N_10393,N_9859,N_9639);
or U10394 (N_10394,N_9940,N_9892);
or U10395 (N_10395,N_9864,N_9754);
and U10396 (N_10396,N_9535,N_9794);
xnor U10397 (N_10397,N_9792,N_9576);
nor U10398 (N_10398,N_9659,N_9592);
nand U10399 (N_10399,N_9841,N_9729);
nor U10400 (N_10400,N_9724,N_9816);
nand U10401 (N_10401,N_9722,N_9564);
and U10402 (N_10402,N_9820,N_9592);
nor U10403 (N_10403,N_9996,N_9718);
and U10404 (N_10404,N_9911,N_9602);
or U10405 (N_10405,N_9657,N_9886);
and U10406 (N_10406,N_9557,N_9787);
nand U10407 (N_10407,N_9921,N_9793);
nor U10408 (N_10408,N_9802,N_9773);
nand U10409 (N_10409,N_9828,N_9549);
and U10410 (N_10410,N_9946,N_9891);
or U10411 (N_10411,N_9683,N_9510);
or U10412 (N_10412,N_9925,N_9617);
nor U10413 (N_10413,N_9721,N_9717);
nand U10414 (N_10414,N_9938,N_9757);
xnor U10415 (N_10415,N_9942,N_9510);
or U10416 (N_10416,N_9690,N_9771);
nor U10417 (N_10417,N_9795,N_9786);
nor U10418 (N_10418,N_9995,N_9758);
nand U10419 (N_10419,N_9657,N_9982);
nor U10420 (N_10420,N_9931,N_9730);
or U10421 (N_10421,N_9895,N_9879);
nor U10422 (N_10422,N_9715,N_9587);
nand U10423 (N_10423,N_9975,N_9816);
nand U10424 (N_10424,N_9594,N_9948);
nor U10425 (N_10425,N_9583,N_9926);
nor U10426 (N_10426,N_9878,N_9696);
nor U10427 (N_10427,N_9721,N_9723);
and U10428 (N_10428,N_9901,N_9561);
nand U10429 (N_10429,N_9782,N_9699);
nor U10430 (N_10430,N_9823,N_9582);
or U10431 (N_10431,N_9947,N_9824);
or U10432 (N_10432,N_9994,N_9625);
nand U10433 (N_10433,N_9886,N_9753);
and U10434 (N_10434,N_9591,N_9973);
or U10435 (N_10435,N_9710,N_9671);
xor U10436 (N_10436,N_9626,N_9594);
or U10437 (N_10437,N_9978,N_9534);
nand U10438 (N_10438,N_9807,N_9985);
or U10439 (N_10439,N_9509,N_9608);
nand U10440 (N_10440,N_9601,N_9911);
nor U10441 (N_10441,N_9866,N_9682);
nand U10442 (N_10442,N_9583,N_9842);
nor U10443 (N_10443,N_9572,N_9782);
and U10444 (N_10444,N_9603,N_9773);
xnor U10445 (N_10445,N_9847,N_9897);
or U10446 (N_10446,N_9953,N_9860);
nand U10447 (N_10447,N_9985,N_9519);
nand U10448 (N_10448,N_9893,N_9617);
nor U10449 (N_10449,N_9732,N_9919);
nand U10450 (N_10450,N_9590,N_9876);
nand U10451 (N_10451,N_9704,N_9955);
nor U10452 (N_10452,N_9706,N_9629);
xnor U10453 (N_10453,N_9691,N_9964);
nand U10454 (N_10454,N_9861,N_9542);
nand U10455 (N_10455,N_9714,N_9933);
nand U10456 (N_10456,N_9643,N_9581);
nand U10457 (N_10457,N_9894,N_9987);
or U10458 (N_10458,N_9553,N_9627);
xnor U10459 (N_10459,N_9691,N_9774);
and U10460 (N_10460,N_9548,N_9549);
nor U10461 (N_10461,N_9797,N_9678);
nor U10462 (N_10462,N_9975,N_9683);
or U10463 (N_10463,N_9701,N_9696);
nand U10464 (N_10464,N_9526,N_9981);
or U10465 (N_10465,N_9679,N_9938);
nor U10466 (N_10466,N_9726,N_9525);
xor U10467 (N_10467,N_9630,N_9930);
nor U10468 (N_10468,N_9549,N_9522);
nand U10469 (N_10469,N_9545,N_9834);
or U10470 (N_10470,N_9785,N_9625);
or U10471 (N_10471,N_9913,N_9979);
xnor U10472 (N_10472,N_9695,N_9612);
nand U10473 (N_10473,N_9759,N_9953);
nand U10474 (N_10474,N_9866,N_9856);
nor U10475 (N_10475,N_9654,N_9639);
and U10476 (N_10476,N_9662,N_9916);
xnor U10477 (N_10477,N_9995,N_9903);
nand U10478 (N_10478,N_9621,N_9655);
nand U10479 (N_10479,N_9654,N_9886);
xnor U10480 (N_10480,N_9713,N_9758);
and U10481 (N_10481,N_9980,N_9851);
and U10482 (N_10482,N_9952,N_9759);
nor U10483 (N_10483,N_9686,N_9876);
and U10484 (N_10484,N_9688,N_9820);
nand U10485 (N_10485,N_9677,N_9701);
and U10486 (N_10486,N_9842,N_9932);
nand U10487 (N_10487,N_9811,N_9662);
or U10488 (N_10488,N_9664,N_9692);
nor U10489 (N_10489,N_9813,N_9505);
nand U10490 (N_10490,N_9914,N_9626);
or U10491 (N_10491,N_9778,N_9794);
nand U10492 (N_10492,N_9898,N_9777);
nor U10493 (N_10493,N_9553,N_9915);
and U10494 (N_10494,N_9539,N_9858);
and U10495 (N_10495,N_9994,N_9689);
nor U10496 (N_10496,N_9806,N_9633);
xor U10497 (N_10497,N_9685,N_9856);
nand U10498 (N_10498,N_9723,N_9547);
or U10499 (N_10499,N_9668,N_9964);
nor U10500 (N_10500,N_10473,N_10207);
or U10501 (N_10501,N_10328,N_10379);
nand U10502 (N_10502,N_10415,N_10249);
and U10503 (N_10503,N_10324,N_10374);
and U10504 (N_10504,N_10134,N_10326);
nand U10505 (N_10505,N_10124,N_10406);
nor U10506 (N_10506,N_10270,N_10146);
xnor U10507 (N_10507,N_10192,N_10094);
or U10508 (N_10508,N_10010,N_10301);
xor U10509 (N_10509,N_10294,N_10407);
or U10510 (N_10510,N_10375,N_10442);
or U10511 (N_10511,N_10337,N_10269);
nand U10512 (N_10512,N_10239,N_10012);
nor U10513 (N_10513,N_10071,N_10232);
nand U10514 (N_10514,N_10230,N_10130);
and U10515 (N_10515,N_10104,N_10214);
and U10516 (N_10516,N_10266,N_10361);
and U10517 (N_10517,N_10248,N_10150);
or U10518 (N_10518,N_10236,N_10092);
or U10519 (N_10519,N_10009,N_10429);
and U10520 (N_10520,N_10359,N_10366);
nand U10521 (N_10521,N_10042,N_10342);
or U10522 (N_10522,N_10292,N_10199);
and U10523 (N_10523,N_10004,N_10434);
or U10524 (N_10524,N_10467,N_10055);
or U10525 (N_10525,N_10032,N_10077);
or U10526 (N_10526,N_10371,N_10451);
nand U10527 (N_10527,N_10123,N_10365);
or U10528 (N_10528,N_10325,N_10300);
or U10529 (N_10529,N_10212,N_10399);
nand U10530 (N_10530,N_10244,N_10441);
or U10531 (N_10531,N_10091,N_10408);
nand U10532 (N_10532,N_10430,N_10179);
nor U10533 (N_10533,N_10170,N_10193);
nor U10534 (N_10534,N_10386,N_10001);
nand U10535 (N_10535,N_10226,N_10242);
or U10536 (N_10536,N_10318,N_10385);
nor U10537 (N_10537,N_10404,N_10085);
nor U10538 (N_10538,N_10182,N_10126);
or U10539 (N_10539,N_10155,N_10414);
and U10540 (N_10540,N_10479,N_10353);
or U10541 (N_10541,N_10344,N_10175);
and U10542 (N_10542,N_10002,N_10422);
or U10543 (N_10543,N_10351,N_10078);
or U10544 (N_10544,N_10109,N_10265);
and U10545 (N_10545,N_10299,N_10162);
nand U10546 (N_10546,N_10168,N_10487);
or U10547 (N_10547,N_10247,N_10005);
or U10548 (N_10548,N_10343,N_10426);
or U10549 (N_10549,N_10086,N_10152);
nand U10550 (N_10550,N_10132,N_10115);
nor U10551 (N_10551,N_10202,N_10443);
or U10552 (N_10552,N_10433,N_10233);
nor U10553 (N_10553,N_10259,N_10453);
xor U10554 (N_10554,N_10056,N_10417);
nand U10555 (N_10555,N_10052,N_10348);
nor U10556 (N_10556,N_10469,N_10252);
or U10557 (N_10557,N_10000,N_10308);
nand U10558 (N_10558,N_10315,N_10218);
and U10559 (N_10559,N_10229,N_10332);
nor U10560 (N_10560,N_10100,N_10454);
or U10561 (N_10561,N_10046,N_10027);
or U10562 (N_10562,N_10234,N_10310);
or U10563 (N_10563,N_10050,N_10484);
or U10564 (N_10564,N_10497,N_10254);
nand U10565 (N_10565,N_10279,N_10006);
or U10566 (N_10566,N_10014,N_10195);
nor U10567 (N_10567,N_10224,N_10243);
nand U10568 (N_10568,N_10016,N_10447);
nand U10569 (N_10569,N_10278,N_10461);
and U10570 (N_10570,N_10147,N_10200);
xnor U10571 (N_10571,N_10311,N_10201);
and U10572 (N_10572,N_10380,N_10495);
nand U10573 (N_10573,N_10260,N_10312);
xnor U10574 (N_10574,N_10131,N_10045);
and U10575 (N_10575,N_10237,N_10142);
nor U10576 (N_10576,N_10107,N_10151);
nor U10577 (N_10577,N_10491,N_10476);
nor U10578 (N_10578,N_10297,N_10096);
nand U10579 (N_10579,N_10494,N_10076);
xnor U10580 (N_10580,N_10394,N_10320);
nor U10581 (N_10581,N_10456,N_10362);
xnor U10582 (N_10582,N_10220,N_10106);
or U10583 (N_10583,N_10390,N_10464);
or U10584 (N_10584,N_10177,N_10102);
nand U10585 (N_10585,N_10011,N_10127);
and U10586 (N_10586,N_10110,N_10022);
and U10587 (N_10587,N_10117,N_10145);
nand U10588 (N_10588,N_10373,N_10273);
and U10589 (N_10589,N_10338,N_10402);
and U10590 (N_10590,N_10079,N_10477);
or U10591 (N_10591,N_10120,N_10070);
nor U10592 (N_10592,N_10190,N_10166);
or U10593 (N_10593,N_10460,N_10144);
nor U10594 (N_10594,N_10309,N_10184);
or U10595 (N_10595,N_10432,N_10480);
nand U10596 (N_10596,N_10397,N_10267);
and U10597 (N_10597,N_10419,N_10423);
xor U10598 (N_10598,N_10061,N_10329);
nor U10599 (N_10599,N_10080,N_10008);
xor U10600 (N_10600,N_10222,N_10306);
or U10601 (N_10601,N_10053,N_10238);
nor U10602 (N_10602,N_10498,N_10274);
nand U10603 (N_10603,N_10468,N_10213);
and U10604 (N_10604,N_10221,N_10030);
and U10605 (N_10605,N_10240,N_10411);
nor U10606 (N_10606,N_10228,N_10277);
nor U10607 (N_10607,N_10262,N_10290);
nor U10608 (N_10608,N_10398,N_10119);
nor U10609 (N_10609,N_10223,N_10381);
and U10610 (N_10610,N_10227,N_10357);
or U10611 (N_10611,N_10246,N_10368);
xor U10612 (N_10612,N_10251,N_10478);
nor U10613 (N_10613,N_10256,N_10181);
and U10614 (N_10614,N_10438,N_10039);
nor U10615 (N_10615,N_10493,N_10158);
or U10616 (N_10616,N_10206,N_10302);
and U10617 (N_10617,N_10116,N_10336);
or U10618 (N_10618,N_10048,N_10041);
or U10619 (N_10619,N_10472,N_10172);
nand U10620 (N_10620,N_10098,N_10282);
or U10621 (N_10621,N_10471,N_10105);
nor U10622 (N_10622,N_10263,N_10153);
nor U10623 (N_10623,N_10340,N_10174);
nor U10624 (N_10624,N_10445,N_10331);
nor U10625 (N_10625,N_10463,N_10462);
nor U10626 (N_10626,N_10481,N_10210);
xnor U10627 (N_10627,N_10204,N_10341);
nand U10628 (N_10628,N_10424,N_10139);
and U10629 (N_10629,N_10316,N_10029);
xnor U10630 (N_10630,N_10436,N_10095);
and U10631 (N_10631,N_10093,N_10356);
and U10632 (N_10632,N_10349,N_10154);
nor U10633 (N_10633,N_10038,N_10412);
and U10634 (N_10634,N_10160,N_10088);
nand U10635 (N_10635,N_10176,N_10492);
nor U10636 (N_10636,N_10378,N_10285);
nand U10637 (N_10637,N_10196,N_10334);
nand U10638 (N_10638,N_10075,N_10031);
and U10639 (N_10639,N_10036,N_10215);
or U10640 (N_10640,N_10136,N_10090);
nand U10641 (N_10641,N_10217,N_10073);
nor U10642 (N_10642,N_10387,N_10287);
or U10643 (N_10643,N_10271,N_10125);
or U10644 (N_10644,N_10059,N_10191);
and U10645 (N_10645,N_10099,N_10013);
or U10646 (N_10646,N_10023,N_10446);
or U10647 (N_10647,N_10211,N_10347);
nor U10648 (N_10648,N_10482,N_10499);
or U10649 (N_10649,N_10490,N_10483);
and U10650 (N_10650,N_10017,N_10257);
nand U10651 (N_10651,N_10122,N_10288);
and U10652 (N_10652,N_10020,N_10466);
nor U10653 (N_10653,N_10143,N_10164);
nand U10654 (N_10654,N_10103,N_10035);
xnor U10655 (N_10655,N_10313,N_10037);
xnor U10656 (N_10656,N_10382,N_10448);
nand U10657 (N_10657,N_10431,N_10167);
nand U10658 (N_10658,N_10049,N_10437);
xor U10659 (N_10659,N_10264,N_10021);
nand U10660 (N_10660,N_10384,N_10465);
nand U10661 (N_10661,N_10084,N_10339);
xor U10662 (N_10662,N_10118,N_10040);
nor U10663 (N_10663,N_10025,N_10420);
and U10664 (N_10664,N_10372,N_10319);
nor U10665 (N_10665,N_10289,N_10401);
and U10666 (N_10666,N_10452,N_10409);
nor U10667 (N_10667,N_10486,N_10322);
or U10668 (N_10668,N_10111,N_10395);
or U10669 (N_10669,N_10389,N_10108);
or U10670 (N_10670,N_10369,N_10391);
nor U10671 (N_10671,N_10187,N_10064);
nor U10672 (N_10672,N_10296,N_10082);
and U10673 (N_10673,N_10138,N_10307);
or U10674 (N_10674,N_10364,N_10327);
xor U10675 (N_10675,N_10043,N_10425);
nand U10676 (N_10676,N_10067,N_10173);
and U10677 (N_10677,N_10161,N_10293);
xnor U10678 (N_10678,N_10485,N_10439);
or U10679 (N_10679,N_10097,N_10112);
xor U10680 (N_10680,N_10396,N_10074);
xnor U10681 (N_10681,N_10335,N_10028);
and U10682 (N_10682,N_10007,N_10241);
and U10683 (N_10683,N_10072,N_10253);
or U10684 (N_10684,N_10054,N_10458);
and U10685 (N_10685,N_10367,N_10148);
nand U10686 (N_10686,N_10457,N_10258);
nor U10687 (N_10687,N_10455,N_10189);
and U10688 (N_10688,N_10440,N_10169);
nor U10689 (N_10689,N_10129,N_10165);
nor U10690 (N_10690,N_10281,N_10488);
nand U10691 (N_10691,N_10280,N_10268);
nor U10692 (N_10692,N_10255,N_10083);
and U10693 (N_10693,N_10066,N_10283);
or U10694 (N_10694,N_10428,N_10163);
nand U10695 (N_10695,N_10418,N_10101);
or U10696 (N_10696,N_10459,N_10026);
nand U10697 (N_10697,N_10474,N_10358);
nor U10698 (N_10698,N_10034,N_10121);
nor U10699 (N_10699,N_10159,N_10323);
xor U10700 (N_10700,N_10276,N_10295);
and U10701 (N_10701,N_10197,N_10346);
nor U10702 (N_10702,N_10350,N_10033);
or U10703 (N_10703,N_10051,N_10156);
or U10704 (N_10704,N_10235,N_10449);
and U10705 (N_10705,N_10186,N_10180);
or U10706 (N_10706,N_10304,N_10370);
or U10707 (N_10707,N_10421,N_10089);
and U10708 (N_10708,N_10128,N_10377);
or U10709 (N_10709,N_10489,N_10149);
and U10710 (N_10710,N_10317,N_10225);
and U10711 (N_10711,N_10057,N_10393);
and U10712 (N_10712,N_10360,N_10137);
nor U10713 (N_10713,N_10496,N_10321);
xnor U10714 (N_10714,N_10470,N_10185);
nor U10715 (N_10715,N_10286,N_10140);
nor U10716 (N_10716,N_10298,N_10133);
or U10717 (N_10717,N_10403,N_10114);
nand U10718 (N_10718,N_10216,N_10245);
or U10719 (N_10719,N_10141,N_10392);
nor U10720 (N_10720,N_10305,N_10208);
and U10721 (N_10721,N_10015,N_10069);
and U10722 (N_10722,N_10400,N_10376);
nand U10723 (N_10723,N_10209,N_10354);
nor U10724 (N_10724,N_10178,N_10352);
or U10725 (N_10725,N_10219,N_10314);
nor U10726 (N_10726,N_10444,N_10171);
nor U10727 (N_10727,N_10194,N_10383);
and U10728 (N_10728,N_10413,N_10113);
nor U10729 (N_10729,N_10018,N_10231);
xnor U10730 (N_10730,N_10062,N_10410);
and U10731 (N_10731,N_10019,N_10333);
nand U10732 (N_10732,N_10044,N_10272);
or U10733 (N_10733,N_10205,N_10405);
xor U10734 (N_10734,N_10060,N_10081);
or U10735 (N_10735,N_10435,N_10135);
nand U10736 (N_10736,N_10416,N_10363);
and U10737 (N_10737,N_10330,N_10275);
nor U10738 (N_10738,N_10427,N_10203);
nand U10739 (N_10739,N_10157,N_10475);
or U10740 (N_10740,N_10087,N_10003);
nor U10741 (N_10741,N_10047,N_10183);
and U10742 (N_10742,N_10198,N_10068);
and U10743 (N_10743,N_10303,N_10261);
nor U10744 (N_10744,N_10355,N_10250);
nor U10745 (N_10745,N_10291,N_10065);
nor U10746 (N_10746,N_10450,N_10024);
nand U10747 (N_10747,N_10063,N_10284);
xnor U10748 (N_10748,N_10388,N_10058);
and U10749 (N_10749,N_10345,N_10188);
or U10750 (N_10750,N_10424,N_10463);
and U10751 (N_10751,N_10475,N_10423);
and U10752 (N_10752,N_10122,N_10416);
nor U10753 (N_10753,N_10046,N_10449);
nor U10754 (N_10754,N_10260,N_10064);
and U10755 (N_10755,N_10181,N_10146);
or U10756 (N_10756,N_10418,N_10037);
nor U10757 (N_10757,N_10009,N_10437);
nor U10758 (N_10758,N_10062,N_10058);
or U10759 (N_10759,N_10482,N_10139);
nor U10760 (N_10760,N_10250,N_10222);
xor U10761 (N_10761,N_10314,N_10404);
or U10762 (N_10762,N_10058,N_10164);
or U10763 (N_10763,N_10464,N_10300);
or U10764 (N_10764,N_10336,N_10207);
nand U10765 (N_10765,N_10413,N_10259);
nand U10766 (N_10766,N_10114,N_10318);
nor U10767 (N_10767,N_10031,N_10438);
and U10768 (N_10768,N_10438,N_10257);
xor U10769 (N_10769,N_10055,N_10263);
or U10770 (N_10770,N_10027,N_10374);
nand U10771 (N_10771,N_10147,N_10103);
nand U10772 (N_10772,N_10365,N_10274);
nand U10773 (N_10773,N_10225,N_10477);
nor U10774 (N_10774,N_10281,N_10366);
nor U10775 (N_10775,N_10042,N_10411);
nor U10776 (N_10776,N_10044,N_10228);
or U10777 (N_10777,N_10162,N_10126);
nand U10778 (N_10778,N_10141,N_10064);
nand U10779 (N_10779,N_10417,N_10067);
nand U10780 (N_10780,N_10294,N_10492);
nand U10781 (N_10781,N_10365,N_10369);
nor U10782 (N_10782,N_10215,N_10357);
nand U10783 (N_10783,N_10371,N_10165);
nor U10784 (N_10784,N_10089,N_10012);
xnor U10785 (N_10785,N_10363,N_10388);
or U10786 (N_10786,N_10039,N_10345);
xnor U10787 (N_10787,N_10149,N_10126);
nor U10788 (N_10788,N_10368,N_10033);
nand U10789 (N_10789,N_10158,N_10089);
and U10790 (N_10790,N_10397,N_10380);
xnor U10791 (N_10791,N_10096,N_10395);
nor U10792 (N_10792,N_10311,N_10296);
nor U10793 (N_10793,N_10059,N_10055);
and U10794 (N_10794,N_10473,N_10287);
nor U10795 (N_10795,N_10259,N_10048);
or U10796 (N_10796,N_10195,N_10317);
or U10797 (N_10797,N_10362,N_10349);
nor U10798 (N_10798,N_10083,N_10110);
nor U10799 (N_10799,N_10184,N_10418);
xnor U10800 (N_10800,N_10105,N_10438);
nor U10801 (N_10801,N_10177,N_10389);
and U10802 (N_10802,N_10062,N_10430);
nor U10803 (N_10803,N_10400,N_10240);
nor U10804 (N_10804,N_10380,N_10189);
nor U10805 (N_10805,N_10050,N_10409);
xor U10806 (N_10806,N_10063,N_10225);
or U10807 (N_10807,N_10340,N_10363);
or U10808 (N_10808,N_10397,N_10055);
nand U10809 (N_10809,N_10449,N_10154);
or U10810 (N_10810,N_10496,N_10373);
and U10811 (N_10811,N_10134,N_10243);
nor U10812 (N_10812,N_10044,N_10270);
or U10813 (N_10813,N_10254,N_10011);
xnor U10814 (N_10814,N_10187,N_10437);
nand U10815 (N_10815,N_10481,N_10016);
or U10816 (N_10816,N_10142,N_10380);
nor U10817 (N_10817,N_10464,N_10100);
xor U10818 (N_10818,N_10315,N_10043);
nor U10819 (N_10819,N_10063,N_10449);
nand U10820 (N_10820,N_10279,N_10165);
or U10821 (N_10821,N_10124,N_10049);
nor U10822 (N_10822,N_10391,N_10396);
nand U10823 (N_10823,N_10424,N_10338);
or U10824 (N_10824,N_10213,N_10322);
or U10825 (N_10825,N_10051,N_10050);
and U10826 (N_10826,N_10389,N_10360);
and U10827 (N_10827,N_10400,N_10222);
or U10828 (N_10828,N_10272,N_10351);
nor U10829 (N_10829,N_10346,N_10226);
or U10830 (N_10830,N_10007,N_10244);
xnor U10831 (N_10831,N_10084,N_10027);
nor U10832 (N_10832,N_10237,N_10233);
nor U10833 (N_10833,N_10360,N_10160);
nor U10834 (N_10834,N_10217,N_10385);
nand U10835 (N_10835,N_10288,N_10115);
nand U10836 (N_10836,N_10493,N_10315);
nand U10837 (N_10837,N_10285,N_10199);
or U10838 (N_10838,N_10139,N_10173);
nor U10839 (N_10839,N_10197,N_10371);
or U10840 (N_10840,N_10386,N_10013);
and U10841 (N_10841,N_10388,N_10107);
nor U10842 (N_10842,N_10421,N_10131);
or U10843 (N_10843,N_10193,N_10107);
or U10844 (N_10844,N_10236,N_10293);
or U10845 (N_10845,N_10074,N_10478);
and U10846 (N_10846,N_10212,N_10203);
nor U10847 (N_10847,N_10156,N_10305);
or U10848 (N_10848,N_10397,N_10175);
nand U10849 (N_10849,N_10390,N_10158);
or U10850 (N_10850,N_10193,N_10010);
and U10851 (N_10851,N_10358,N_10157);
and U10852 (N_10852,N_10177,N_10188);
or U10853 (N_10853,N_10266,N_10385);
nor U10854 (N_10854,N_10461,N_10155);
nor U10855 (N_10855,N_10443,N_10071);
nor U10856 (N_10856,N_10466,N_10272);
nand U10857 (N_10857,N_10041,N_10494);
nand U10858 (N_10858,N_10120,N_10413);
xor U10859 (N_10859,N_10287,N_10448);
xor U10860 (N_10860,N_10340,N_10457);
nand U10861 (N_10861,N_10269,N_10418);
xnor U10862 (N_10862,N_10462,N_10266);
xor U10863 (N_10863,N_10266,N_10289);
nor U10864 (N_10864,N_10497,N_10073);
and U10865 (N_10865,N_10407,N_10062);
or U10866 (N_10866,N_10010,N_10091);
or U10867 (N_10867,N_10470,N_10289);
nor U10868 (N_10868,N_10423,N_10325);
nor U10869 (N_10869,N_10287,N_10245);
and U10870 (N_10870,N_10458,N_10402);
nand U10871 (N_10871,N_10460,N_10098);
and U10872 (N_10872,N_10200,N_10337);
or U10873 (N_10873,N_10493,N_10323);
or U10874 (N_10874,N_10020,N_10169);
and U10875 (N_10875,N_10169,N_10038);
nor U10876 (N_10876,N_10090,N_10184);
or U10877 (N_10877,N_10439,N_10364);
or U10878 (N_10878,N_10273,N_10113);
and U10879 (N_10879,N_10040,N_10360);
xor U10880 (N_10880,N_10326,N_10449);
xnor U10881 (N_10881,N_10333,N_10080);
nor U10882 (N_10882,N_10453,N_10231);
nand U10883 (N_10883,N_10027,N_10162);
and U10884 (N_10884,N_10158,N_10482);
nor U10885 (N_10885,N_10207,N_10321);
nor U10886 (N_10886,N_10289,N_10021);
or U10887 (N_10887,N_10473,N_10162);
or U10888 (N_10888,N_10437,N_10301);
nor U10889 (N_10889,N_10243,N_10222);
nand U10890 (N_10890,N_10026,N_10217);
or U10891 (N_10891,N_10400,N_10381);
and U10892 (N_10892,N_10243,N_10039);
or U10893 (N_10893,N_10350,N_10013);
nor U10894 (N_10894,N_10312,N_10194);
or U10895 (N_10895,N_10057,N_10008);
and U10896 (N_10896,N_10078,N_10219);
xnor U10897 (N_10897,N_10351,N_10060);
nand U10898 (N_10898,N_10204,N_10157);
or U10899 (N_10899,N_10058,N_10242);
or U10900 (N_10900,N_10387,N_10317);
nor U10901 (N_10901,N_10353,N_10344);
and U10902 (N_10902,N_10494,N_10233);
and U10903 (N_10903,N_10397,N_10029);
or U10904 (N_10904,N_10493,N_10307);
nor U10905 (N_10905,N_10188,N_10242);
or U10906 (N_10906,N_10452,N_10495);
or U10907 (N_10907,N_10102,N_10041);
nand U10908 (N_10908,N_10485,N_10114);
nor U10909 (N_10909,N_10279,N_10244);
nand U10910 (N_10910,N_10125,N_10015);
nand U10911 (N_10911,N_10022,N_10196);
nor U10912 (N_10912,N_10063,N_10391);
and U10913 (N_10913,N_10445,N_10118);
nor U10914 (N_10914,N_10000,N_10222);
nor U10915 (N_10915,N_10264,N_10259);
nor U10916 (N_10916,N_10391,N_10124);
and U10917 (N_10917,N_10279,N_10203);
nand U10918 (N_10918,N_10067,N_10388);
and U10919 (N_10919,N_10408,N_10203);
xor U10920 (N_10920,N_10157,N_10299);
or U10921 (N_10921,N_10457,N_10292);
nand U10922 (N_10922,N_10067,N_10364);
nand U10923 (N_10923,N_10083,N_10456);
and U10924 (N_10924,N_10402,N_10470);
nand U10925 (N_10925,N_10421,N_10285);
nand U10926 (N_10926,N_10170,N_10034);
nand U10927 (N_10927,N_10382,N_10407);
nor U10928 (N_10928,N_10065,N_10262);
nor U10929 (N_10929,N_10245,N_10265);
or U10930 (N_10930,N_10399,N_10134);
nor U10931 (N_10931,N_10001,N_10024);
and U10932 (N_10932,N_10155,N_10382);
nand U10933 (N_10933,N_10218,N_10336);
nor U10934 (N_10934,N_10388,N_10454);
nor U10935 (N_10935,N_10026,N_10204);
nand U10936 (N_10936,N_10236,N_10475);
or U10937 (N_10937,N_10338,N_10107);
and U10938 (N_10938,N_10156,N_10091);
xnor U10939 (N_10939,N_10416,N_10358);
nand U10940 (N_10940,N_10475,N_10012);
xor U10941 (N_10941,N_10207,N_10267);
and U10942 (N_10942,N_10282,N_10326);
nand U10943 (N_10943,N_10249,N_10404);
and U10944 (N_10944,N_10092,N_10352);
xnor U10945 (N_10945,N_10429,N_10197);
nand U10946 (N_10946,N_10427,N_10279);
nand U10947 (N_10947,N_10199,N_10147);
nor U10948 (N_10948,N_10142,N_10074);
and U10949 (N_10949,N_10318,N_10232);
nor U10950 (N_10950,N_10179,N_10417);
or U10951 (N_10951,N_10114,N_10440);
xor U10952 (N_10952,N_10099,N_10499);
or U10953 (N_10953,N_10329,N_10416);
or U10954 (N_10954,N_10290,N_10415);
and U10955 (N_10955,N_10003,N_10496);
nand U10956 (N_10956,N_10336,N_10212);
nor U10957 (N_10957,N_10025,N_10071);
xnor U10958 (N_10958,N_10077,N_10022);
or U10959 (N_10959,N_10282,N_10394);
nor U10960 (N_10960,N_10427,N_10213);
nand U10961 (N_10961,N_10065,N_10071);
nor U10962 (N_10962,N_10131,N_10191);
nand U10963 (N_10963,N_10445,N_10438);
and U10964 (N_10964,N_10278,N_10313);
xnor U10965 (N_10965,N_10391,N_10208);
or U10966 (N_10966,N_10096,N_10416);
and U10967 (N_10967,N_10442,N_10283);
nand U10968 (N_10968,N_10029,N_10482);
or U10969 (N_10969,N_10270,N_10103);
nand U10970 (N_10970,N_10342,N_10231);
and U10971 (N_10971,N_10317,N_10365);
or U10972 (N_10972,N_10086,N_10130);
or U10973 (N_10973,N_10143,N_10088);
nor U10974 (N_10974,N_10078,N_10203);
or U10975 (N_10975,N_10403,N_10420);
xor U10976 (N_10976,N_10152,N_10407);
xnor U10977 (N_10977,N_10261,N_10005);
nor U10978 (N_10978,N_10185,N_10133);
xnor U10979 (N_10979,N_10222,N_10163);
or U10980 (N_10980,N_10181,N_10023);
nor U10981 (N_10981,N_10426,N_10492);
xor U10982 (N_10982,N_10154,N_10222);
or U10983 (N_10983,N_10149,N_10130);
or U10984 (N_10984,N_10118,N_10037);
or U10985 (N_10985,N_10369,N_10396);
nand U10986 (N_10986,N_10407,N_10155);
or U10987 (N_10987,N_10311,N_10254);
or U10988 (N_10988,N_10270,N_10357);
nor U10989 (N_10989,N_10239,N_10458);
nand U10990 (N_10990,N_10474,N_10493);
or U10991 (N_10991,N_10455,N_10228);
or U10992 (N_10992,N_10410,N_10430);
and U10993 (N_10993,N_10027,N_10358);
nor U10994 (N_10994,N_10337,N_10287);
or U10995 (N_10995,N_10033,N_10031);
and U10996 (N_10996,N_10018,N_10265);
nand U10997 (N_10997,N_10144,N_10209);
or U10998 (N_10998,N_10440,N_10092);
nand U10999 (N_10999,N_10253,N_10446);
nor U11000 (N_11000,N_10618,N_10528);
nand U11001 (N_11001,N_10999,N_10645);
nand U11002 (N_11002,N_10535,N_10769);
nor U11003 (N_11003,N_10792,N_10959);
nand U11004 (N_11004,N_10891,N_10894);
nor U11005 (N_11005,N_10990,N_10724);
and U11006 (N_11006,N_10865,N_10550);
xor U11007 (N_11007,N_10875,N_10907);
nand U11008 (N_11008,N_10937,N_10838);
xor U11009 (N_11009,N_10670,N_10938);
nand U11010 (N_11010,N_10939,N_10668);
xnor U11011 (N_11011,N_10658,N_10635);
nand U11012 (N_11012,N_10783,N_10915);
and U11013 (N_11013,N_10923,N_10630);
or U11014 (N_11014,N_10814,N_10788);
or U11015 (N_11015,N_10733,N_10772);
or U11016 (N_11016,N_10702,N_10958);
or U11017 (N_11017,N_10995,N_10538);
xnor U11018 (N_11018,N_10812,N_10912);
nand U11019 (N_11019,N_10977,N_10966);
nand U11020 (N_11020,N_10732,N_10597);
and U11021 (N_11021,N_10942,N_10968);
nor U11022 (N_11022,N_10614,N_10564);
nor U11023 (N_11023,N_10544,N_10862);
xnor U11024 (N_11024,N_10761,N_10619);
and U11025 (N_11025,N_10699,N_10613);
or U11026 (N_11026,N_10898,N_10830);
nand U11027 (N_11027,N_10636,N_10845);
or U11028 (N_11028,N_10980,N_10571);
nand U11029 (N_11029,N_10701,N_10957);
nor U11030 (N_11030,N_10657,N_10554);
nor U11031 (N_11031,N_10580,N_10688);
nor U11032 (N_11032,N_10622,N_10847);
and U11033 (N_11033,N_10671,N_10978);
nand U11034 (N_11034,N_10951,N_10866);
nor U11035 (N_11035,N_10893,N_10969);
xor U11036 (N_11036,N_10537,N_10527);
nor U11037 (N_11037,N_10900,N_10698);
nand U11038 (N_11038,N_10746,N_10950);
and U11039 (N_11039,N_10903,N_10648);
nand U11040 (N_11040,N_10642,N_10586);
and U11041 (N_11041,N_10581,N_10921);
nor U11042 (N_11042,N_10863,N_10762);
and U11043 (N_11043,N_10956,N_10821);
and U11044 (N_11044,N_10652,N_10567);
nand U11045 (N_11045,N_10722,N_10787);
nor U11046 (N_11046,N_10556,N_10555);
nor U11047 (N_11047,N_10974,N_10822);
or U11048 (N_11048,N_10515,N_10694);
nor U11049 (N_11049,N_10770,N_10578);
and U11050 (N_11050,N_10982,N_10911);
nand U11051 (N_11051,N_10935,N_10629);
and U11052 (N_11052,N_10771,N_10522);
nor U11053 (N_11053,N_10611,N_10596);
nand U11054 (N_11054,N_10773,N_10602);
or U11055 (N_11055,N_10692,N_10895);
nor U11056 (N_11056,N_10574,N_10712);
or U11057 (N_11057,N_10782,N_10885);
nand U11058 (N_11058,N_10612,N_10716);
nand U11059 (N_11059,N_10971,N_10810);
nor U11060 (N_11060,N_10967,N_10906);
nand U11061 (N_11061,N_10811,N_10638);
and U11062 (N_11062,N_10627,N_10615);
nor U11063 (N_11063,N_10815,N_10928);
nor U11064 (N_11064,N_10779,N_10690);
or U11065 (N_11065,N_10919,N_10726);
and U11066 (N_11066,N_10513,N_10637);
nand U11067 (N_11067,N_10632,N_10616);
nor U11068 (N_11068,N_10710,N_10641);
xnor U11069 (N_11069,N_10849,N_10674);
or U11070 (N_11070,N_10925,N_10667);
nor U11071 (N_11071,N_10867,N_10519);
nor U11072 (N_11072,N_10704,N_10888);
nand U11073 (N_11073,N_10665,N_10936);
nor U11074 (N_11074,N_10896,N_10708);
or U11075 (N_11075,N_10809,N_10512);
and U11076 (N_11076,N_10548,N_10856);
nand U11077 (N_11077,N_10709,N_10926);
or U11078 (N_11078,N_10504,N_10656);
nor U11079 (N_11079,N_10789,N_10514);
nor U11080 (N_11080,N_10557,N_10774);
nand U11081 (N_11081,N_10904,N_10598);
nand U11082 (N_11082,N_10947,N_10795);
and U11083 (N_11083,N_10836,N_10517);
and U11084 (N_11084,N_10687,N_10878);
nor U11085 (N_11085,N_10905,N_10521);
and U11086 (N_11086,N_10890,N_10643);
or U11087 (N_11087,N_10510,N_10520);
or U11088 (N_11088,N_10780,N_10981);
and U11089 (N_11089,N_10759,N_10591);
nor U11090 (N_11090,N_10543,N_10565);
and U11091 (N_11091,N_10914,N_10979);
and U11092 (N_11092,N_10502,N_10884);
nor U11093 (N_11093,N_10996,N_10531);
nand U11094 (N_11094,N_10559,N_10801);
and U11095 (N_11095,N_10837,N_10758);
and U11096 (N_11096,N_10786,N_10748);
xnor U11097 (N_11097,N_10998,N_10852);
and U11098 (N_11098,N_10620,N_10601);
or U11099 (N_11099,N_10902,N_10997);
nor U11100 (N_11100,N_10608,N_10575);
nor U11101 (N_11101,N_10857,N_10889);
nand U11102 (N_11102,N_10714,N_10719);
nor U11103 (N_11103,N_10546,N_10684);
or U11104 (N_11104,N_10853,N_10717);
or U11105 (N_11105,N_10595,N_10600);
nor U11106 (N_11106,N_10593,N_10713);
and U11107 (N_11107,N_10763,N_10539);
and U11108 (N_11108,N_10953,N_10844);
or U11109 (N_11109,N_10541,N_10963);
nor U11110 (N_11110,N_10775,N_10633);
nor U11111 (N_11111,N_10874,N_10932);
or U11112 (N_11112,N_10617,N_10877);
and U11113 (N_11113,N_10825,N_10561);
nor U11114 (N_11114,N_10587,N_10910);
nor U11115 (N_11115,N_10655,N_10695);
and U11116 (N_11116,N_10576,N_10827);
nor U11117 (N_11117,N_10609,N_10718);
and U11118 (N_11118,N_10745,N_10841);
nand U11119 (N_11119,N_10760,N_10946);
nor U11120 (N_11120,N_10983,N_10924);
nand U11121 (N_11121,N_10833,N_10854);
nor U11122 (N_11122,N_10834,N_10507);
or U11123 (N_11123,N_10785,N_10518);
and U11124 (N_11124,N_10679,N_10545);
nand U11125 (N_11125,N_10945,N_10736);
nand U11126 (N_11126,N_10964,N_10659);
or U11127 (N_11127,N_10603,N_10920);
or U11128 (N_11128,N_10835,N_10523);
nor U11129 (N_11129,N_10654,N_10840);
and U11130 (N_11130,N_10589,N_10858);
nand U11131 (N_11131,N_10917,N_10994);
nor U11132 (N_11132,N_10508,N_10828);
nor U11133 (N_11133,N_10563,N_10876);
and U11134 (N_11134,N_10634,N_10880);
nor U11135 (N_11135,N_10927,N_10560);
or U11136 (N_11136,N_10807,N_10682);
or U11137 (N_11137,N_10813,N_10738);
nand U11138 (N_11138,N_10913,N_10871);
nand U11139 (N_11139,N_10529,N_10664);
nand U11140 (N_11140,N_10992,N_10505);
or U11141 (N_11141,N_10816,N_10689);
xor U11142 (N_11142,N_10625,N_10826);
or U11143 (N_11143,N_10988,N_10952);
or U11144 (N_11144,N_10729,N_10700);
nor U11145 (N_11145,N_10703,N_10805);
nand U11146 (N_11146,N_10585,N_10842);
or U11147 (N_11147,N_10623,N_10931);
nand U11148 (N_11148,N_10594,N_10940);
and U11149 (N_11149,N_10540,N_10941);
xnor U11150 (N_11150,N_10954,N_10723);
or U11151 (N_11151,N_10933,N_10949);
and U11152 (N_11152,N_10678,N_10922);
xnor U11153 (N_11153,N_10588,N_10944);
or U11154 (N_11154,N_10778,N_10579);
nor U11155 (N_11155,N_10899,N_10943);
nand U11156 (N_11156,N_10647,N_10570);
and U11157 (N_11157,N_10989,N_10973);
or U11158 (N_11158,N_10735,N_10800);
and U11159 (N_11159,N_10551,N_10509);
or U11160 (N_11160,N_10864,N_10721);
and U11161 (N_11161,N_10605,N_10572);
or U11162 (N_11162,N_10511,N_10797);
nor U11163 (N_11163,N_10887,N_10839);
xnor U11164 (N_11164,N_10743,N_10848);
nor U11165 (N_11165,N_10651,N_10725);
and U11166 (N_11166,N_10534,N_10972);
and U11167 (N_11167,N_10882,N_10790);
and U11168 (N_11168,N_10530,N_10776);
and U11169 (N_11169,N_10532,N_10868);
or U11170 (N_11170,N_10742,N_10784);
nor U11171 (N_11171,N_10777,N_10639);
and U11172 (N_11172,N_10803,N_10820);
or U11173 (N_11173,N_10599,N_10650);
or U11174 (N_11174,N_10693,N_10558);
or U11175 (N_11175,N_10930,N_10987);
nor U11176 (N_11176,N_10646,N_10886);
or U11177 (N_11177,N_10621,N_10744);
and U11178 (N_11178,N_10960,N_10583);
nor U11179 (N_11179,N_10680,N_10881);
nand U11180 (N_11180,N_10962,N_10753);
nand U11181 (N_11181,N_10961,N_10796);
xnor U11182 (N_11182,N_10610,N_10749);
nor U11183 (N_11183,N_10955,N_10536);
and U11184 (N_11184,N_10542,N_10824);
and U11185 (N_11185,N_10756,N_10757);
nand U11186 (N_11186,N_10976,N_10644);
and U11187 (N_11187,N_10706,N_10901);
or U11188 (N_11188,N_10577,N_10985);
or U11189 (N_11189,N_10553,N_10851);
nand U11190 (N_11190,N_10663,N_10991);
nor U11191 (N_11191,N_10607,N_10737);
nand U11192 (N_11192,N_10666,N_10897);
nand U11193 (N_11193,N_10582,N_10802);
nor U11194 (N_11194,N_10547,N_10649);
or U11195 (N_11195,N_10503,N_10685);
xnor U11196 (N_11196,N_10506,N_10817);
nand U11197 (N_11197,N_10869,N_10566);
nand U11198 (N_11198,N_10873,N_10720);
or U11199 (N_11199,N_10752,N_10751);
nor U11200 (N_11200,N_10765,N_10677);
or U11201 (N_11201,N_10681,N_10855);
nor U11202 (N_11202,N_10740,N_10909);
xnor U11203 (N_11203,N_10916,N_10831);
or U11204 (N_11204,N_10755,N_10832);
nor U11205 (N_11205,N_10584,N_10918);
and U11206 (N_11206,N_10697,N_10970);
and U11207 (N_11207,N_10791,N_10569);
nand U11208 (N_11208,N_10766,N_10727);
nand U11209 (N_11209,N_10526,N_10846);
nor U11210 (N_11210,N_10662,N_10929);
and U11211 (N_11211,N_10683,N_10516);
nand U11212 (N_11212,N_10892,N_10843);
and U11213 (N_11213,N_10660,N_10606);
or U11214 (N_11214,N_10592,N_10715);
nand U11215 (N_11215,N_10500,N_10626);
nor U11216 (N_11216,N_10691,N_10879);
xor U11217 (N_11217,N_10806,N_10754);
nor U11218 (N_11218,N_10747,N_10804);
or U11219 (N_11219,N_10781,N_10908);
or U11220 (N_11220,N_10986,N_10562);
and U11221 (N_11221,N_10975,N_10823);
and U11222 (N_11222,N_10750,N_10861);
and U11223 (N_11223,N_10883,N_10794);
and U11224 (N_11224,N_10604,N_10533);
nand U11225 (N_11225,N_10669,N_10676);
nor U11226 (N_11226,N_10872,N_10984);
xor U11227 (N_11227,N_10696,N_10739);
nand U11228 (N_11228,N_10549,N_10799);
nand U11229 (N_11229,N_10730,N_10552);
xnor U11230 (N_11230,N_10628,N_10850);
nand U11231 (N_11231,N_10767,N_10573);
nand U11232 (N_11232,N_10798,N_10965);
nand U11233 (N_11233,N_10590,N_10675);
nor U11234 (N_11234,N_10859,N_10705);
and U11235 (N_11235,N_10818,N_10686);
xor U11236 (N_11236,N_10673,N_10764);
or U11237 (N_11237,N_10993,N_10734);
and U11238 (N_11238,N_10934,N_10731);
nor U11239 (N_11239,N_10829,N_10948);
and U11240 (N_11240,N_10860,N_10624);
nor U11241 (N_11241,N_10707,N_10640);
and U11242 (N_11242,N_10672,N_10501);
and U11243 (N_11243,N_10819,N_10568);
xor U11244 (N_11244,N_10525,N_10808);
or U11245 (N_11245,N_10768,N_10870);
or U11246 (N_11246,N_10793,N_10741);
nand U11247 (N_11247,N_10631,N_10711);
nor U11248 (N_11248,N_10728,N_10524);
or U11249 (N_11249,N_10661,N_10653);
nand U11250 (N_11250,N_10981,N_10684);
nand U11251 (N_11251,N_10990,N_10603);
nor U11252 (N_11252,N_10744,N_10807);
nand U11253 (N_11253,N_10892,N_10620);
or U11254 (N_11254,N_10766,N_10970);
or U11255 (N_11255,N_10505,N_10792);
nand U11256 (N_11256,N_10895,N_10951);
and U11257 (N_11257,N_10550,N_10683);
and U11258 (N_11258,N_10655,N_10631);
nor U11259 (N_11259,N_10726,N_10532);
or U11260 (N_11260,N_10896,N_10898);
nand U11261 (N_11261,N_10575,N_10639);
or U11262 (N_11262,N_10751,N_10730);
or U11263 (N_11263,N_10760,N_10986);
xnor U11264 (N_11264,N_10714,N_10794);
or U11265 (N_11265,N_10660,N_10735);
nand U11266 (N_11266,N_10608,N_10845);
nor U11267 (N_11267,N_10973,N_10942);
nor U11268 (N_11268,N_10516,N_10689);
nor U11269 (N_11269,N_10670,N_10502);
and U11270 (N_11270,N_10528,N_10873);
and U11271 (N_11271,N_10969,N_10902);
nand U11272 (N_11272,N_10868,N_10522);
xor U11273 (N_11273,N_10961,N_10797);
nor U11274 (N_11274,N_10934,N_10969);
or U11275 (N_11275,N_10926,N_10750);
nand U11276 (N_11276,N_10586,N_10887);
and U11277 (N_11277,N_10534,N_10882);
xor U11278 (N_11278,N_10946,N_10806);
and U11279 (N_11279,N_10652,N_10643);
or U11280 (N_11280,N_10841,N_10691);
nand U11281 (N_11281,N_10644,N_10576);
or U11282 (N_11282,N_10764,N_10913);
nand U11283 (N_11283,N_10952,N_10916);
or U11284 (N_11284,N_10594,N_10943);
nand U11285 (N_11285,N_10573,N_10774);
and U11286 (N_11286,N_10539,N_10737);
nor U11287 (N_11287,N_10511,N_10773);
and U11288 (N_11288,N_10528,N_10586);
and U11289 (N_11289,N_10962,N_10546);
nor U11290 (N_11290,N_10990,N_10829);
and U11291 (N_11291,N_10819,N_10692);
nor U11292 (N_11292,N_10733,N_10832);
and U11293 (N_11293,N_10644,N_10522);
nand U11294 (N_11294,N_10992,N_10643);
or U11295 (N_11295,N_10727,N_10969);
nor U11296 (N_11296,N_10654,N_10657);
nand U11297 (N_11297,N_10851,N_10948);
and U11298 (N_11298,N_10901,N_10507);
nor U11299 (N_11299,N_10947,N_10674);
nand U11300 (N_11300,N_10837,N_10874);
or U11301 (N_11301,N_10681,N_10973);
or U11302 (N_11302,N_10638,N_10850);
and U11303 (N_11303,N_10919,N_10678);
and U11304 (N_11304,N_10727,N_10504);
and U11305 (N_11305,N_10835,N_10647);
nand U11306 (N_11306,N_10584,N_10624);
and U11307 (N_11307,N_10693,N_10894);
xor U11308 (N_11308,N_10877,N_10999);
nor U11309 (N_11309,N_10893,N_10592);
and U11310 (N_11310,N_10812,N_10667);
nor U11311 (N_11311,N_10930,N_10831);
or U11312 (N_11312,N_10647,N_10848);
nor U11313 (N_11313,N_10791,N_10646);
or U11314 (N_11314,N_10916,N_10646);
nand U11315 (N_11315,N_10812,N_10838);
nand U11316 (N_11316,N_10697,N_10908);
or U11317 (N_11317,N_10672,N_10927);
or U11318 (N_11318,N_10697,N_10922);
nor U11319 (N_11319,N_10811,N_10835);
nor U11320 (N_11320,N_10633,N_10539);
or U11321 (N_11321,N_10731,N_10880);
xnor U11322 (N_11322,N_10772,N_10760);
or U11323 (N_11323,N_10883,N_10679);
and U11324 (N_11324,N_10515,N_10626);
and U11325 (N_11325,N_10645,N_10755);
and U11326 (N_11326,N_10726,N_10535);
nor U11327 (N_11327,N_10723,N_10629);
and U11328 (N_11328,N_10836,N_10599);
or U11329 (N_11329,N_10761,N_10743);
and U11330 (N_11330,N_10710,N_10996);
nand U11331 (N_11331,N_10854,N_10845);
nor U11332 (N_11332,N_10764,N_10759);
xor U11333 (N_11333,N_10826,N_10903);
or U11334 (N_11334,N_10760,N_10893);
or U11335 (N_11335,N_10643,N_10633);
xor U11336 (N_11336,N_10860,N_10602);
or U11337 (N_11337,N_10792,N_10860);
nand U11338 (N_11338,N_10735,N_10825);
nand U11339 (N_11339,N_10783,N_10949);
nor U11340 (N_11340,N_10853,N_10933);
nor U11341 (N_11341,N_10597,N_10898);
xnor U11342 (N_11342,N_10549,N_10539);
xnor U11343 (N_11343,N_10788,N_10736);
nor U11344 (N_11344,N_10962,N_10767);
nand U11345 (N_11345,N_10932,N_10852);
and U11346 (N_11346,N_10564,N_10632);
xor U11347 (N_11347,N_10616,N_10882);
nand U11348 (N_11348,N_10521,N_10800);
xor U11349 (N_11349,N_10713,N_10671);
nor U11350 (N_11350,N_10923,N_10985);
nor U11351 (N_11351,N_10804,N_10593);
xnor U11352 (N_11352,N_10546,N_10934);
nand U11353 (N_11353,N_10998,N_10753);
or U11354 (N_11354,N_10731,N_10695);
or U11355 (N_11355,N_10625,N_10987);
and U11356 (N_11356,N_10915,N_10650);
or U11357 (N_11357,N_10643,N_10742);
and U11358 (N_11358,N_10898,N_10953);
or U11359 (N_11359,N_10543,N_10556);
and U11360 (N_11360,N_10531,N_10649);
and U11361 (N_11361,N_10972,N_10641);
and U11362 (N_11362,N_10524,N_10809);
nand U11363 (N_11363,N_10929,N_10689);
nand U11364 (N_11364,N_10680,N_10797);
nor U11365 (N_11365,N_10618,N_10891);
and U11366 (N_11366,N_10631,N_10809);
xor U11367 (N_11367,N_10923,N_10824);
or U11368 (N_11368,N_10727,N_10633);
nand U11369 (N_11369,N_10675,N_10900);
and U11370 (N_11370,N_10819,N_10769);
nand U11371 (N_11371,N_10610,N_10670);
or U11372 (N_11372,N_10726,N_10906);
nor U11373 (N_11373,N_10575,N_10995);
and U11374 (N_11374,N_10781,N_10651);
xor U11375 (N_11375,N_10852,N_10918);
nand U11376 (N_11376,N_10822,N_10670);
nand U11377 (N_11377,N_10592,N_10857);
nor U11378 (N_11378,N_10767,N_10740);
xnor U11379 (N_11379,N_10621,N_10702);
or U11380 (N_11380,N_10752,N_10932);
and U11381 (N_11381,N_10944,N_10623);
and U11382 (N_11382,N_10615,N_10905);
nand U11383 (N_11383,N_10942,N_10791);
nor U11384 (N_11384,N_10619,N_10956);
or U11385 (N_11385,N_10699,N_10810);
and U11386 (N_11386,N_10977,N_10821);
and U11387 (N_11387,N_10896,N_10697);
or U11388 (N_11388,N_10932,N_10832);
or U11389 (N_11389,N_10629,N_10671);
nor U11390 (N_11390,N_10717,N_10809);
and U11391 (N_11391,N_10965,N_10739);
nand U11392 (N_11392,N_10615,N_10952);
nor U11393 (N_11393,N_10563,N_10998);
or U11394 (N_11394,N_10915,N_10592);
nor U11395 (N_11395,N_10547,N_10588);
or U11396 (N_11396,N_10825,N_10569);
and U11397 (N_11397,N_10822,N_10706);
and U11398 (N_11398,N_10520,N_10502);
and U11399 (N_11399,N_10517,N_10841);
or U11400 (N_11400,N_10654,N_10916);
nand U11401 (N_11401,N_10927,N_10627);
nor U11402 (N_11402,N_10646,N_10600);
or U11403 (N_11403,N_10998,N_10738);
or U11404 (N_11404,N_10846,N_10923);
nand U11405 (N_11405,N_10776,N_10578);
or U11406 (N_11406,N_10985,N_10668);
nor U11407 (N_11407,N_10883,N_10797);
or U11408 (N_11408,N_10984,N_10853);
nand U11409 (N_11409,N_10635,N_10750);
or U11410 (N_11410,N_10678,N_10905);
or U11411 (N_11411,N_10848,N_10892);
nor U11412 (N_11412,N_10716,N_10626);
xnor U11413 (N_11413,N_10818,N_10906);
or U11414 (N_11414,N_10797,N_10839);
nand U11415 (N_11415,N_10985,N_10616);
or U11416 (N_11416,N_10503,N_10837);
or U11417 (N_11417,N_10643,N_10989);
or U11418 (N_11418,N_10776,N_10664);
nand U11419 (N_11419,N_10893,N_10778);
and U11420 (N_11420,N_10819,N_10883);
nor U11421 (N_11421,N_10955,N_10869);
nand U11422 (N_11422,N_10576,N_10847);
nand U11423 (N_11423,N_10611,N_10653);
or U11424 (N_11424,N_10739,N_10794);
nand U11425 (N_11425,N_10548,N_10593);
or U11426 (N_11426,N_10816,N_10971);
nor U11427 (N_11427,N_10951,N_10724);
or U11428 (N_11428,N_10980,N_10638);
nor U11429 (N_11429,N_10708,N_10754);
nand U11430 (N_11430,N_10509,N_10822);
nor U11431 (N_11431,N_10742,N_10560);
and U11432 (N_11432,N_10630,N_10685);
nor U11433 (N_11433,N_10794,N_10930);
nor U11434 (N_11434,N_10749,N_10865);
and U11435 (N_11435,N_10877,N_10791);
and U11436 (N_11436,N_10734,N_10583);
nor U11437 (N_11437,N_10557,N_10865);
and U11438 (N_11438,N_10508,N_10558);
nor U11439 (N_11439,N_10975,N_10653);
or U11440 (N_11440,N_10558,N_10556);
or U11441 (N_11441,N_10625,N_10714);
or U11442 (N_11442,N_10941,N_10548);
nor U11443 (N_11443,N_10779,N_10659);
nor U11444 (N_11444,N_10861,N_10931);
nor U11445 (N_11445,N_10545,N_10876);
xor U11446 (N_11446,N_10703,N_10660);
nor U11447 (N_11447,N_10845,N_10605);
nand U11448 (N_11448,N_10630,N_10639);
nor U11449 (N_11449,N_10591,N_10930);
and U11450 (N_11450,N_10868,N_10937);
nor U11451 (N_11451,N_10773,N_10733);
and U11452 (N_11452,N_10973,N_10771);
nor U11453 (N_11453,N_10631,N_10714);
and U11454 (N_11454,N_10514,N_10991);
and U11455 (N_11455,N_10965,N_10549);
and U11456 (N_11456,N_10894,N_10853);
or U11457 (N_11457,N_10924,N_10968);
nand U11458 (N_11458,N_10683,N_10997);
or U11459 (N_11459,N_10552,N_10981);
and U11460 (N_11460,N_10955,N_10901);
and U11461 (N_11461,N_10550,N_10541);
or U11462 (N_11462,N_10870,N_10513);
nand U11463 (N_11463,N_10932,N_10563);
and U11464 (N_11464,N_10950,N_10849);
nor U11465 (N_11465,N_10987,N_10830);
and U11466 (N_11466,N_10875,N_10610);
or U11467 (N_11467,N_10938,N_10718);
nor U11468 (N_11468,N_10702,N_10668);
nor U11469 (N_11469,N_10765,N_10946);
xor U11470 (N_11470,N_10709,N_10625);
and U11471 (N_11471,N_10590,N_10657);
and U11472 (N_11472,N_10800,N_10986);
nand U11473 (N_11473,N_10506,N_10844);
or U11474 (N_11474,N_10795,N_10788);
nand U11475 (N_11475,N_10518,N_10650);
nor U11476 (N_11476,N_10828,N_10986);
or U11477 (N_11477,N_10962,N_10551);
and U11478 (N_11478,N_10834,N_10550);
nor U11479 (N_11479,N_10696,N_10672);
and U11480 (N_11480,N_10853,N_10595);
and U11481 (N_11481,N_10611,N_10671);
nand U11482 (N_11482,N_10984,N_10899);
and U11483 (N_11483,N_10508,N_10555);
and U11484 (N_11484,N_10997,N_10961);
nor U11485 (N_11485,N_10831,N_10758);
and U11486 (N_11486,N_10546,N_10837);
and U11487 (N_11487,N_10886,N_10772);
nor U11488 (N_11488,N_10537,N_10542);
xor U11489 (N_11489,N_10709,N_10509);
and U11490 (N_11490,N_10584,N_10606);
xor U11491 (N_11491,N_10572,N_10865);
nor U11492 (N_11492,N_10710,N_10776);
or U11493 (N_11493,N_10678,N_10516);
nand U11494 (N_11494,N_10953,N_10803);
or U11495 (N_11495,N_10867,N_10520);
or U11496 (N_11496,N_10682,N_10559);
nor U11497 (N_11497,N_10819,N_10724);
nand U11498 (N_11498,N_10520,N_10880);
nor U11499 (N_11499,N_10696,N_10716);
or U11500 (N_11500,N_11137,N_11256);
xnor U11501 (N_11501,N_11226,N_11412);
or U11502 (N_11502,N_11111,N_11090);
nor U11503 (N_11503,N_11307,N_11324);
and U11504 (N_11504,N_11127,N_11171);
or U11505 (N_11505,N_11318,N_11225);
or U11506 (N_11506,N_11378,N_11250);
nand U11507 (N_11507,N_11325,N_11148);
xnor U11508 (N_11508,N_11022,N_11163);
xnor U11509 (N_11509,N_11154,N_11195);
nor U11510 (N_11510,N_11006,N_11233);
nor U11511 (N_11511,N_11252,N_11169);
nor U11512 (N_11512,N_11160,N_11278);
or U11513 (N_11513,N_11141,N_11096);
nand U11514 (N_11514,N_11164,N_11286);
nor U11515 (N_11515,N_11176,N_11411);
nand U11516 (N_11516,N_11298,N_11395);
or U11517 (N_11517,N_11198,N_11317);
and U11518 (N_11518,N_11280,N_11194);
nand U11519 (N_11519,N_11049,N_11130);
or U11520 (N_11520,N_11266,N_11426);
nor U11521 (N_11521,N_11143,N_11467);
or U11522 (N_11522,N_11145,N_11190);
or U11523 (N_11523,N_11028,N_11429);
nand U11524 (N_11524,N_11000,N_11044);
nor U11525 (N_11525,N_11067,N_11264);
xnor U11526 (N_11526,N_11206,N_11421);
and U11527 (N_11527,N_11161,N_11249);
and U11528 (N_11528,N_11455,N_11401);
xnor U11529 (N_11529,N_11155,N_11251);
xnor U11530 (N_11530,N_11487,N_11201);
xor U11531 (N_11531,N_11413,N_11216);
nand U11532 (N_11532,N_11178,N_11191);
nand U11533 (N_11533,N_11323,N_11099);
or U11534 (N_11534,N_11053,N_11349);
nand U11535 (N_11535,N_11075,N_11045);
or U11536 (N_11536,N_11147,N_11149);
nor U11537 (N_11537,N_11026,N_11361);
nand U11538 (N_11538,N_11407,N_11446);
xnor U11539 (N_11539,N_11393,N_11156);
and U11540 (N_11540,N_11300,N_11210);
or U11541 (N_11541,N_11382,N_11268);
and U11542 (N_11542,N_11257,N_11105);
and U11543 (N_11543,N_11232,N_11065);
or U11544 (N_11544,N_11416,N_11061);
nand U11545 (N_11545,N_11261,N_11094);
and U11546 (N_11546,N_11348,N_11418);
and U11547 (N_11547,N_11379,N_11463);
nor U11548 (N_11548,N_11387,N_11299);
and U11549 (N_11549,N_11224,N_11010);
xor U11550 (N_11550,N_11084,N_11012);
nor U11551 (N_11551,N_11151,N_11255);
xor U11552 (N_11552,N_11482,N_11088);
nor U11553 (N_11553,N_11402,N_11024);
and U11554 (N_11554,N_11124,N_11309);
nand U11555 (N_11555,N_11409,N_11289);
nor U11556 (N_11556,N_11098,N_11396);
or U11557 (N_11557,N_11039,N_11265);
nand U11558 (N_11558,N_11474,N_11374);
and U11559 (N_11559,N_11048,N_11433);
and U11560 (N_11560,N_11177,N_11381);
and U11561 (N_11561,N_11112,N_11020);
nand U11562 (N_11562,N_11037,N_11306);
xor U11563 (N_11563,N_11436,N_11346);
nor U11564 (N_11564,N_11046,N_11362);
or U11565 (N_11565,N_11313,N_11495);
nor U11566 (N_11566,N_11092,N_11352);
nor U11567 (N_11567,N_11002,N_11437);
nor U11568 (N_11568,N_11340,N_11335);
or U11569 (N_11569,N_11471,N_11184);
nor U11570 (N_11570,N_11139,N_11050);
nand U11571 (N_11571,N_11218,N_11034);
and U11572 (N_11572,N_11469,N_11089);
and U11573 (N_11573,N_11312,N_11043);
or U11574 (N_11574,N_11366,N_11245);
nor U11575 (N_11575,N_11117,N_11449);
nor U11576 (N_11576,N_11447,N_11102);
or U11577 (N_11577,N_11167,N_11454);
or U11578 (N_11578,N_11125,N_11083);
and U11579 (N_11579,N_11027,N_11386);
nor U11580 (N_11580,N_11486,N_11247);
xnor U11581 (N_11581,N_11485,N_11244);
and U11582 (N_11582,N_11331,N_11473);
xor U11583 (N_11583,N_11142,N_11023);
nand U11584 (N_11584,N_11319,N_11439);
nand U11585 (N_11585,N_11337,N_11347);
nor U11586 (N_11586,N_11419,N_11234);
xor U11587 (N_11587,N_11015,N_11108);
nor U11588 (N_11588,N_11363,N_11458);
nor U11589 (N_11589,N_11276,N_11047);
nor U11590 (N_11590,N_11253,N_11456);
nand U11591 (N_11591,N_11399,N_11480);
or U11592 (N_11592,N_11284,N_11060);
and U11593 (N_11593,N_11059,N_11077);
xnor U11594 (N_11594,N_11263,N_11427);
and U11595 (N_11595,N_11484,N_11370);
and U11596 (N_11596,N_11078,N_11132);
or U11597 (N_11597,N_11259,N_11009);
or U11598 (N_11598,N_11172,N_11274);
nand U11599 (N_11599,N_11287,N_11041);
nor U11600 (N_11600,N_11272,N_11403);
and U11601 (N_11601,N_11466,N_11476);
xnor U11602 (N_11602,N_11380,N_11036);
nor U11603 (N_11603,N_11478,N_11062);
and U11604 (N_11604,N_11158,N_11301);
and U11605 (N_11605,N_11042,N_11377);
nor U11606 (N_11606,N_11129,N_11384);
and U11607 (N_11607,N_11071,N_11410);
nor U11608 (N_11608,N_11350,N_11074);
and U11609 (N_11609,N_11180,N_11038);
or U11610 (N_11610,N_11116,N_11351);
or U11611 (N_11611,N_11193,N_11293);
or U11612 (N_11612,N_11063,N_11070);
or U11613 (N_11613,N_11073,N_11223);
and U11614 (N_11614,N_11275,N_11087);
or U11615 (N_11615,N_11030,N_11248);
nor U11616 (N_11616,N_11270,N_11353);
or U11617 (N_11617,N_11296,N_11461);
and U11618 (N_11618,N_11457,N_11295);
nand U11619 (N_11619,N_11114,N_11425);
nor U11620 (N_11620,N_11031,N_11240);
or U11621 (N_11621,N_11336,N_11004);
nor U11622 (N_11622,N_11271,N_11103);
and U11623 (N_11623,N_11477,N_11435);
and U11624 (N_11624,N_11242,N_11133);
nor U11625 (N_11625,N_11122,N_11490);
and U11626 (N_11626,N_11290,N_11170);
or U11627 (N_11627,N_11267,N_11235);
or U11628 (N_11628,N_11007,N_11499);
or U11629 (N_11629,N_11135,N_11011);
nor U11630 (N_11630,N_11238,N_11262);
nand U11631 (N_11631,N_11442,N_11183);
nand U11632 (N_11632,N_11040,N_11021);
and U11633 (N_11633,N_11064,N_11231);
nor U11634 (N_11634,N_11364,N_11080);
nand U11635 (N_11635,N_11304,N_11450);
and U11636 (N_11636,N_11205,N_11221);
or U11637 (N_11637,N_11152,N_11339);
or U11638 (N_11638,N_11136,N_11097);
nor U11639 (N_11639,N_11391,N_11302);
and U11640 (N_11640,N_11315,N_11444);
nand U11641 (N_11641,N_11260,N_11372);
or U11642 (N_11642,N_11128,N_11294);
or U11643 (N_11643,N_11134,N_11157);
xnor U11644 (N_11644,N_11213,N_11175);
and U11645 (N_11645,N_11229,N_11441);
nor U11646 (N_11646,N_11375,N_11415);
or U11647 (N_11647,N_11373,N_11327);
or U11648 (N_11648,N_11222,N_11291);
nand U11649 (N_11649,N_11185,N_11292);
or U11650 (N_11650,N_11016,N_11123);
nand U11651 (N_11651,N_11118,N_11445);
or U11652 (N_11652,N_11470,N_11330);
nand U11653 (N_11653,N_11144,N_11192);
xor U11654 (N_11654,N_11334,N_11095);
and U11655 (N_11655,N_11008,N_11448);
nor U11656 (N_11656,N_11168,N_11239);
or U11657 (N_11657,N_11431,N_11109);
and U11658 (N_11658,N_11357,N_11138);
or U11659 (N_11659,N_11173,N_11342);
and U11660 (N_11660,N_11254,N_11199);
nand U11661 (N_11661,N_11121,N_11068);
xnor U11662 (N_11662,N_11269,N_11496);
nor U11663 (N_11663,N_11150,N_11406);
nor U11664 (N_11664,N_11033,N_11104);
and U11665 (N_11665,N_11032,N_11314);
nand U11666 (N_11666,N_11228,N_11475);
and U11667 (N_11667,N_11014,N_11243);
nand U11668 (N_11668,N_11390,N_11273);
nand U11669 (N_11669,N_11131,N_11430);
and U11670 (N_11670,N_11029,N_11054);
nor U11671 (N_11671,N_11333,N_11285);
and U11672 (N_11672,N_11303,N_11186);
nand U11673 (N_11673,N_11057,N_11432);
nand U11674 (N_11674,N_11187,N_11297);
or U11675 (N_11675,N_11283,N_11472);
and U11676 (N_11676,N_11069,N_11106);
or U11677 (N_11677,N_11417,N_11460);
nand U11678 (N_11678,N_11422,N_11019);
nor U11679 (N_11679,N_11072,N_11483);
nor U11680 (N_11680,N_11211,N_11440);
and U11681 (N_11681,N_11209,N_11326);
or U11682 (N_11682,N_11321,N_11491);
nor U11683 (N_11683,N_11498,N_11208);
nand U11684 (N_11684,N_11423,N_11214);
or U11685 (N_11685,N_11236,N_11207);
or U11686 (N_11686,N_11345,N_11196);
nor U11687 (N_11687,N_11497,N_11365);
nor U11688 (N_11688,N_11091,N_11146);
or U11689 (N_11689,N_11188,N_11489);
nor U11690 (N_11690,N_11126,N_11003);
nor U11691 (N_11691,N_11166,N_11197);
or U11692 (N_11692,N_11076,N_11343);
or U11693 (N_11693,N_11203,N_11189);
nor U11694 (N_11694,N_11093,N_11464);
nand U11695 (N_11695,N_11277,N_11025);
xor U11696 (N_11696,N_11165,N_11308);
nor U11697 (N_11697,N_11488,N_11389);
xor U11698 (N_11698,N_11465,N_11397);
nand U11699 (N_11699,N_11107,N_11359);
and U11700 (N_11700,N_11101,N_11215);
xor U11701 (N_11701,N_11282,N_11369);
nor U11702 (N_11702,N_11162,N_11428);
nor U11703 (N_11703,N_11241,N_11182);
nor U11704 (N_11704,N_11332,N_11305);
or U11705 (N_11705,N_11035,N_11005);
nand U11706 (N_11706,N_11311,N_11434);
or U11707 (N_11707,N_11204,N_11200);
nor U11708 (N_11708,N_11086,N_11338);
and U11709 (N_11709,N_11310,N_11328);
nand U11710 (N_11710,N_11341,N_11051);
and U11711 (N_11711,N_11358,N_11279);
and U11712 (N_11712,N_11494,N_11344);
xor U11713 (N_11713,N_11220,N_11159);
nor U11714 (N_11714,N_11082,N_11288);
nor U11715 (N_11715,N_11398,N_11281);
xor U11716 (N_11716,N_11081,N_11453);
nand U11717 (N_11717,N_11388,N_11120);
nand U11718 (N_11718,N_11451,N_11212);
nand U11719 (N_11719,N_11459,N_11376);
or U11720 (N_11720,N_11404,N_11153);
and U11721 (N_11721,N_11385,N_11230);
and U11722 (N_11722,N_11492,N_11079);
and U11723 (N_11723,N_11400,N_11320);
nand U11724 (N_11724,N_11356,N_11202);
nand U11725 (N_11725,N_11113,N_11452);
nand U11726 (N_11726,N_11219,N_11066);
xnor U11727 (N_11727,N_11258,N_11394);
nand U11728 (N_11728,N_11001,N_11414);
and U11729 (N_11729,N_11110,N_11462);
and U11730 (N_11730,N_11371,N_11179);
nand U11731 (N_11731,N_11443,N_11316);
nand U11732 (N_11732,N_11013,N_11392);
or U11733 (N_11733,N_11383,N_11174);
and U11734 (N_11734,N_11408,N_11237);
nor U11735 (N_11735,N_11115,N_11018);
or U11736 (N_11736,N_11368,N_11140);
and U11737 (N_11737,N_11056,N_11017);
and U11738 (N_11738,N_11355,N_11424);
nand U11739 (N_11739,N_11119,N_11085);
and U11740 (N_11740,N_11055,N_11181);
and U11741 (N_11741,N_11052,N_11227);
nand U11742 (N_11742,N_11405,N_11493);
nor U11743 (N_11743,N_11420,N_11322);
xnor U11744 (N_11744,N_11354,N_11479);
nor U11745 (N_11745,N_11438,N_11329);
or U11746 (N_11746,N_11468,N_11367);
or U11747 (N_11747,N_11058,N_11360);
or U11748 (N_11748,N_11481,N_11217);
or U11749 (N_11749,N_11100,N_11246);
and U11750 (N_11750,N_11265,N_11403);
nor U11751 (N_11751,N_11453,N_11063);
and U11752 (N_11752,N_11277,N_11497);
or U11753 (N_11753,N_11064,N_11426);
nor U11754 (N_11754,N_11102,N_11040);
or U11755 (N_11755,N_11351,N_11457);
or U11756 (N_11756,N_11247,N_11287);
xnor U11757 (N_11757,N_11386,N_11033);
and U11758 (N_11758,N_11451,N_11441);
and U11759 (N_11759,N_11290,N_11484);
xnor U11760 (N_11760,N_11219,N_11334);
nand U11761 (N_11761,N_11399,N_11195);
or U11762 (N_11762,N_11189,N_11367);
nand U11763 (N_11763,N_11306,N_11382);
and U11764 (N_11764,N_11442,N_11017);
nand U11765 (N_11765,N_11183,N_11329);
and U11766 (N_11766,N_11154,N_11021);
nand U11767 (N_11767,N_11357,N_11158);
nor U11768 (N_11768,N_11374,N_11057);
or U11769 (N_11769,N_11213,N_11454);
nor U11770 (N_11770,N_11131,N_11007);
nor U11771 (N_11771,N_11130,N_11090);
xor U11772 (N_11772,N_11355,N_11334);
and U11773 (N_11773,N_11025,N_11382);
and U11774 (N_11774,N_11013,N_11354);
nor U11775 (N_11775,N_11133,N_11083);
and U11776 (N_11776,N_11113,N_11083);
or U11777 (N_11777,N_11134,N_11094);
nand U11778 (N_11778,N_11129,N_11351);
nor U11779 (N_11779,N_11155,N_11137);
or U11780 (N_11780,N_11257,N_11090);
or U11781 (N_11781,N_11125,N_11208);
xor U11782 (N_11782,N_11379,N_11150);
nor U11783 (N_11783,N_11023,N_11117);
and U11784 (N_11784,N_11093,N_11105);
nand U11785 (N_11785,N_11470,N_11340);
and U11786 (N_11786,N_11024,N_11122);
nor U11787 (N_11787,N_11467,N_11119);
nor U11788 (N_11788,N_11329,N_11271);
nor U11789 (N_11789,N_11172,N_11486);
nand U11790 (N_11790,N_11039,N_11267);
or U11791 (N_11791,N_11394,N_11364);
nor U11792 (N_11792,N_11249,N_11091);
xor U11793 (N_11793,N_11439,N_11000);
or U11794 (N_11794,N_11116,N_11232);
and U11795 (N_11795,N_11209,N_11140);
nor U11796 (N_11796,N_11051,N_11001);
nand U11797 (N_11797,N_11171,N_11165);
nand U11798 (N_11798,N_11176,N_11236);
or U11799 (N_11799,N_11053,N_11481);
or U11800 (N_11800,N_11363,N_11022);
nand U11801 (N_11801,N_11026,N_11388);
and U11802 (N_11802,N_11324,N_11012);
nand U11803 (N_11803,N_11284,N_11275);
nand U11804 (N_11804,N_11145,N_11060);
and U11805 (N_11805,N_11410,N_11333);
nand U11806 (N_11806,N_11019,N_11014);
nand U11807 (N_11807,N_11057,N_11255);
xor U11808 (N_11808,N_11431,N_11274);
nor U11809 (N_11809,N_11114,N_11491);
xnor U11810 (N_11810,N_11390,N_11079);
nor U11811 (N_11811,N_11109,N_11025);
nor U11812 (N_11812,N_11429,N_11210);
or U11813 (N_11813,N_11201,N_11021);
or U11814 (N_11814,N_11010,N_11423);
nor U11815 (N_11815,N_11103,N_11386);
or U11816 (N_11816,N_11481,N_11391);
nor U11817 (N_11817,N_11375,N_11362);
nor U11818 (N_11818,N_11456,N_11189);
and U11819 (N_11819,N_11410,N_11055);
and U11820 (N_11820,N_11127,N_11378);
nor U11821 (N_11821,N_11466,N_11474);
nor U11822 (N_11822,N_11442,N_11206);
nor U11823 (N_11823,N_11291,N_11052);
nor U11824 (N_11824,N_11081,N_11454);
or U11825 (N_11825,N_11420,N_11252);
nand U11826 (N_11826,N_11267,N_11134);
nand U11827 (N_11827,N_11265,N_11004);
or U11828 (N_11828,N_11434,N_11099);
nor U11829 (N_11829,N_11225,N_11138);
and U11830 (N_11830,N_11284,N_11458);
or U11831 (N_11831,N_11134,N_11321);
or U11832 (N_11832,N_11436,N_11103);
and U11833 (N_11833,N_11490,N_11196);
nand U11834 (N_11834,N_11448,N_11316);
nand U11835 (N_11835,N_11383,N_11150);
nor U11836 (N_11836,N_11235,N_11360);
nor U11837 (N_11837,N_11168,N_11427);
nor U11838 (N_11838,N_11283,N_11081);
nand U11839 (N_11839,N_11361,N_11148);
and U11840 (N_11840,N_11206,N_11261);
and U11841 (N_11841,N_11322,N_11205);
nand U11842 (N_11842,N_11030,N_11134);
nand U11843 (N_11843,N_11238,N_11489);
and U11844 (N_11844,N_11311,N_11357);
nor U11845 (N_11845,N_11481,N_11469);
nor U11846 (N_11846,N_11436,N_11370);
or U11847 (N_11847,N_11105,N_11098);
nor U11848 (N_11848,N_11004,N_11426);
and U11849 (N_11849,N_11102,N_11199);
and U11850 (N_11850,N_11040,N_11011);
or U11851 (N_11851,N_11124,N_11126);
xnor U11852 (N_11852,N_11249,N_11228);
and U11853 (N_11853,N_11224,N_11024);
and U11854 (N_11854,N_11410,N_11036);
xnor U11855 (N_11855,N_11008,N_11096);
or U11856 (N_11856,N_11205,N_11389);
xnor U11857 (N_11857,N_11337,N_11039);
nor U11858 (N_11858,N_11477,N_11112);
xor U11859 (N_11859,N_11492,N_11069);
nor U11860 (N_11860,N_11189,N_11013);
nor U11861 (N_11861,N_11110,N_11263);
nand U11862 (N_11862,N_11036,N_11275);
and U11863 (N_11863,N_11114,N_11056);
nand U11864 (N_11864,N_11263,N_11103);
nand U11865 (N_11865,N_11190,N_11348);
xor U11866 (N_11866,N_11176,N_11189);
nor U11867 (N_11867,N_11254,N_11149);
nor U11868 (N_11868,N_11273,N_11411);
and U11869 (N_11869,N_11318,N_11115);
and U11870 (N_11870,N_11034,N_11190);
nand U11871 (N_11871,N_11448,N_11117);
nand U11872 (N_11872,N_11081,N_11366);
or U11873 (N_11873,N_11090,N_11148);
or U11874 (N_11874,N_11014,N_11480);
nand U11875 (N_11875,N_11394,N_11128);
or U11876 (N_11876,N_11281,N_11062);
nand U11877 (N_11877,N_11157,N_11167);
and U11878 (N_11878,N_11389,N_11431);
nor U11879 (N_11879,N_11163,N_11103);
nand U11880 (N_11880,N_11430,N_11085);
nand U11881 (N_11881,N_11083,N_11004);
and U11882 (N_11882,N_11209,N_11342);
or U11883 (N_11883,N_11416,N_11151);
and U11884 (N_11884,N_11215,N_11143);
nor U11885 (N_11885,N_11053,N_11176);
nor U11886 (N_11886,N_11058,N_11146);
or U11887 (N_11887,N_11470,N_11469);
nor U11888 (N_11888,N_11343,N_11015);
xor U11889 (N_11889,N_11393,N_11029);
nand U11890 (N_11890,N_11184,N_11172);
nand U11891 (N_11891,N_11239,N_11068);
nand U11892 (N_11892,N_11329,N_11156);
nor U11893 (N_11893,N_11224,N_11131);
nor U11894 (N_11894,N_11284,N_11449);
or U11895 (N_11895,N_11279,N_11005);
nand U11896 (N_11896,N_11066,N_11490);
and U11897 (N_11897,N_11222,N_11318);
nor U11898 (N_11898,N_11353,N_11059);
nand U11899 (N_11899,N_11255,N_11456);
nor U11900 (N_11900,N_11134,N_11004);
nand U11901 (N_11901,N_11083,N_11407);
or U11902 (N_11902,N_11109,N_11061);
nor U11903 (N_11903,N_11302,N_11063);
nor U11904 (N_11904,N_11389,N_11263);
and U11905 (N_11905,N_11462,N_11369);
nand U11906 (N_11906,N_11142,N_11208);
or U11907 (N_11907,N_11457,N_11028);
or U11908 (N_11908,N_11240,N_11382);
nand U11909 (N_11909,N_11259,N_11129);
nand U11910 (N_11910,N_11020,N_11032);
and U11911 (N_11911,N_11222,N_11422);
xor U11912 (N_11912,N_11290,N_11085);
and U11913 (N_11913,N_11360,N_11393);
or U11914 (N_11914,N_11018,N_11039);
nor U11915 (N_11915,N_11058,N_11045);
or U11916 (N_11916,N_11246,N_11260);
or U11917 (N_11917,N_11485,N_11258);
nand U11918 (N_11918,N_11286,N_11029);
or U11919 (N_11919,N_11396,N_11217);
nor U11920 (N_11920,N_11498,N_11377);
and U11921 (N_11921,N_11410,N_11198);
or U11922 (N_11922,N_11009,N_11121);
nand U11923 (N_11923,N_11344,N_11319);
nor U11924 (N_11924,N_11018,N_11110);
and U11925 (N_11925,N_11413,N_11272);
nor U11926 (N_11926,N_11367,N_11407);
and U11927 (N_11927,N_11368,N_11049);
nor U11928 (N_11928,N_11017,N_11321);
or U11929 (N_11929,N_11393,N_11152);
nor U11930 (N_11930,N_11259,N_11384);
or U11931 (N_11931,N_11312,N_11490);
xor U11932 (N_11932,N_11051,N_11211);
or U11933 (N_11933,N_11254,N_11074);
or U11934 (N_11934,N_11064,N_11016);
or U11935 (N_11935,N_11405,N_11351);
nor U11936 (N_11936,N_11097,N_11466);
nor U11937 (N_11937,N_11119,N_11134);
or U11938 (N_11938,N_11386,N_11298);
nand U11939 (N_11939,N_11451,N_11168);
nand U11940 (N_11940,N_11006,N_11052);
or U11941 (N_11941,N_11276,N_11477);
or U11942 (N_11942,N_11301,N_11397);
nand U11943 (N_11943,N_11310,N_11162);
and U11944 (N_11944,N_11431,N_11348);
nand U11945 (N_11945,N_11315,N_11155);
nand U11946 (N_11946,N_11198,N_11372);
or U11947 (N_11947,N_11143,N_11318);
and U11948 (N_11948,N_11025,N_11017);
nand U11949 (N_11949,N_11101,N_11018);
or U11950 (N_11950,N_11381,N_11076);
nand U11951 (N_11951,N_11321,N_11373);
nor U11952 (N_11952,N_11122,N_11282);
nand U11953 (N_11953,N_11204,N_11118);
nand U11954 (N_11954,N_11445,N_11191);
nand U11955 (N_11955,N_11236,N_11076);
or U11956 (N_11956,N_11233,N_11074);
or U11957 (N_11957,N_11048,N_11036);
or U11958 (N_11958,N_11332,N_11344);
nand U11959 (N_11959,N_11041,N_11198);
or U11960 (N_11960,N_11284,N_11327);
or U11961 (N_11961,N_11357,N_11026);
xor U11962 (N_11962,N_11160,N_11039);
nand U11963 (N_11963,N_11300,N_11092);
nor U11964 (N_11964,N_11204,N_11355);
nand U11965 (N_11965,N_11338,N_11260);
nor U11966 (N_11966,N_11256,N_11481);
and U11967 (N_11967,N_11291,N_11043);
and U11968 (N_11968,N_11430,N_11128);
and U11969 (N_11969,N_11482,N_11001);
nor U11970 (N_11970,N_11071,N_11067);
nor U11971 (N_11971,N_11046,N_11080);
or U11972 (N_11972,N_11443,N_11371);
or U11973 (N_11973,N_11488,N_11438);
nand U11974 (N_11974,N_11396,N_11257);
nand U11975 (N_11975,N_11008,N_11236);
nor U11976 (N_11976,N_11320,N_11194);
and U11977 (N_11977,N_11280,N_11210);
and U11978 (N_11978,N_11441,N_11194);
nor U11979 (N_11979,N_11343,N_11464);
or U11980 (N_11980,N_11146,N_11228);
nand U11981 (N_11981,N_11432,N_11331);
nand U11982 (N_11982,N_11129,N_11444);
or U11983 (N_11983,N_11011,N_11396);
and U11984 (N_11984,N_11042,N_11160);
or U11985 (N_11985,N_11231,N_11490);
nand U11986 (N_11986,N_11364,N_11194);
nand U11987 (N_11987,N_11383,N_11209);
nand U11988 (N_11988,N_11408,N_11458);
and U11989 (N_11989,N_11122,N_11001);
nand U11990 (N_11990,N_11240,N_11185);
nand U11991 (N_11991,N_11393,N_11355);
or U11992 (N_11992,N_11060,N_11287);
nor U11993 (N_11993,N_11414,N_11229);
or U11994 (N_11994,N_11328,N_11012);
nand U11995 (N_11995,N_11443,N_11463);
nor U11996 (N_11996,N_11134,N_11217);
nand U11997 (N_11997,N_11237,N_11456);
nor U11998 (N_11998,N_11167,N_11005);
nand U11999 (N_11999,N_11468,N_11454);
and U12000 (N_12000,N_11770,N_11606);
nor U12001 (N_12001,N_11631,N_11515);
or U12002 (N_12002,N_11500,N_11579);
nor U12003 (N_12003,N_11640,N_11540);
xnor U12004 (N_12004,N_11560,N_11543);
or U12005 (N_12005,N_11815,N_11521);
nand U12006 (N_12006,N_11690,N_11988);
nand U12007 (N_12007,N_11787,N_11747);
and U12008 (N_12008,N_11888,N_11875);
nand U12009 (N_12009,N_11971,N_11637);
xnor U12010 (N_12010,N_11677,N_11600);
nand U12011 (N_12011,N_11683,N_11975);
nand U12012 (N_12012,N_11907,N_11718);
nor U12013 (N_12013,N_11964,N_11555);
nor U12014 (N_12014,N_11726,N_11845);
and U12015 (N_12015,N_11750,N_11506);
or U12016 (N_12016,N_11922,N_11531);
or U12017 (N_12017,N_11928,N_11517);
or U12018 (N_12018,N_11742,N_11647);
nand U12019 (N_12019,N_11614,N_11778);
xnor U12020 (N_12020,N_11520,N_11666);
nand U12021 (N_12021,N_11705,N_11590);
and U12022 (N_12022,N_11923,N_11735);
nand U12023 (N_12023,N_11566,N_11648);
nand U12024 (N_12024,N_11977,N_11974);
or U12025 (N_12025,N_11986,N_11536);
and U12026 (N_12026,N_11908,N_11527);
and U12027 (N_12027,N_11684,N_11915);
nand U12028 (N_12028,N_11502,N_11550);
nand U12029 (N_12029,N_11645,N_11562);
nor U12030 (N_12030,N_11879,N_11938);
or U12031 (N_12031,N_11842,N_11693);
or U12032 (N_12032,N_11511,N_11834);
or U12033 (N_12033,N_11546,N_11811);
xor U12034 (N_12034,N_11903,N_11697);
nor U12035 (N_12035,N_11574,N_11594);
or U12036 (N_12036,N_11899,N_11840);
or U12037 (N_12037,N_11725,N_11777);
nand U12038 (N_12038,N_11706,N_11970);
nand U12039 (N_12039,N_11558,N_11931);
nand U12040 (N_12040,N_11769,N_11918);
and U12041 (N_12041,N_11618,N_11663);
or U12042 (N_12042,N_11681,N_11968);
xor U12043 (N_12043,N_11940,N_11837);
and U12044 (N_12044,N_11680,N_11696);
or U12045 (N_12045,N_11779,N_11675);
and U12046 (N_12046,N_11549,N_11982);
and U12047 (N_12047,N_11993,N_11623);
nand U12048 (N_12048,N_11987,N_11757);
nor U12049 (N_12049,N_11793,N_11951);
and U12050 (N_12050,N_11906,N_11597);
nor U12051 (N_12051,N_11700,N_11619);
and U12052 (N_12052,N_11821,N_11836);
and U12053 (N_12053,N_11796,N_11547);
nor U12054 (N_12054,N_11573,N_11810);
nor U12055 (N_12055,N_11716,N_11545);
nor U12056 (N_12056,N_11734,N_11900);
or U12057 (N_12057,N_11702,N_11665);
nand U12058 (N_12058,N_11801,N_11633);
xor U12059 (N_12059,N_11751,N_11676);
or U12060 (N_12060,N_11715,N_11865);
nor U12061 (N_12061,N_11638,N_11587);
nor U12062 (N_12062,N_11723,N_11823);
and U12063 (N_12063,N_11866,N_11630);
or U12064 (N_12064,N_11776,N_11501);
or U12065 (N_12065,N_11727,N_11695);
and U12066 (N_12066,N_11768,N_11744);
and U12067 (N_12067,N_11965,N_11952);
and U12068 (N_12068,N_11670,N_11992);
nand U12069 (N_12069,N_11892,N_11671);
nor U12070 (N_12070,N_11831,N_11529);
and U12071 (N_12071,N_11824,N_11598);
and U12072 (N_12072,N_11884,N_11516);
nand U12073 (N_12073,N_11858,N_11868);
or U12074 (N_12074,N_11891,N_11593);
nand U12075 (N_12075,N_11791,N_11848);
nor U12076 (N_12076,N_11651,N_11973);
nor U12077 (N_12077,N_11936,N_11841);
or U12078 (N_12078,N_11513,N_11958);
or U12079 (N_12079,N_11847,N_11689);
nor U12080 (N_12080,N_11911,N_11565);
nor U12081 (N_12081,N_11551,N_11771);
nor U12082 (N_12082,N_11781,N_11530);
and U12083 (N_12083,N_11518,N_11615);
and U12084 (N_12084,N_11621,N_11917);
xnor U12085 (N_12085,N_11902,N_11783);
nand U12086 (N_12086,N_11981,N_11962);
nor U12087 (N_12087,N_11584,N_11567);
nor U12088 (N_12088,N_11732,N_11758);
and U12089 (N_12089,N_11925,N_11800);
or U12090 (N_12090,N_11886,N_11883);
nor U12091 (N_12091,N_11978,N_11658);
nor U12092 (N_12092,N_11914,N_11814);
xnor U12093 (N_12093,N_11649,N_11904);
nand U12094 (N_12094,N_11660,N_11708);
xor U12095 (N_12095,N_11882,N_11743);
xnor U12096 (N_12096,N_11785,N_11577);
and U12097 (N_12097,N_11827,N_11818);
and U12098 (N_12098,N_11642,N_11997);
nor U12099 (N_12099,N_11844,N_11853);
nor U12100 (N_12100,N_11976,N_11504);
nor U12101 (N_12101,N_11678,N_11859);
nor U12102 (N_12102,N_11673,N_11712);
nand U12103 (N_12103,N_11953,N_11766);
xor U12104 (N_12104,N_11874,N_11804);
nor U12105 (N_12105,N_11701,N_11505);
nor U12106 (N_12106,N_11806,N_11763);
nand U12107 (N_12107,N_11581,N_11628);
or U12108 (N_12108,N_11654,N_11947);
xor U12109 (N_12109,N_11538,N_11912);
nand U12110 (N_12110,N_11755,N_11991);
or U12111 (N_12111,N_11659,N_11752);
or U12112 (N_12112,N_11887,N_11756);
or U12113 (N_12113,N_11950,N_11588);
and U12114 (N_12114,N_11578,N_11956);
and U12115 (N_12115,N_11881,N_11672);
nor U12116 (N_12116,N_11604,N_11568);
nand U12117 (N_12117,N_11780,N_11629);
nor U12118 (N_12118,N_11688,N_11998);
nor U12119 (N_12119,N_11507,N_11620);
nand U12120 (N_12120,N_11849,N_11905);
and U12121 (N_12121,N_11609,N_11720);
nand U12122 (N_12122,N_11709,N_11772);
and U12123 (N_12123,N_11786,N_11949);
or U12124 (N_12124,N_11765,N_11602);
nor U12125 (N_12125,N_11556,N_11897);
nor U12126 (N_12126,N_11599,N_11586);
or U12127 (N_12127,N_11959,N_11890);
nand U12128 (N_12128,N_11664,N_11661);
nand U12129 (N_12129,N_11924,N_11554);
and U12130 (N_12130,N_11961,N_11526);
nor U12131 (N_12131,N_11969,N_11534);
or U12132 (N_12132,N_11722,N_11807);
and U12133 (N_12133,N_11762,N_11559);
nand U12134 (N_12134,N_11731,N_11724);
or U12135 (N_12135,N_11963,N_11585);
nor U12136 (N_12136,N_11685,N_11605);
nor U12137 (N_12137,N_11601,N_11860);
and U12138 (N_12138,N_11730,N_11935);
nand U12139 (N_12139,N_11707,N_11512);
xnor U12140 (N_12140,N_11980,N_11764);
nand U12141 (N_12141,N_11533,N_11930);
nor U12142 (N_12142,N_11611,N_11850);
xor U12143 (N_12143,N_11896,N_11522);
and U12144 (N_12144,N_11563,N_11652);
xnor U12145 (N_12145,N_11608,N_11564);
nand U12146 (N_12146,N_11552,N_11535);
or U12147 (N_12147,N_11544,N_11561);
or U12148 (N_12148,N_11941,N_11851);
xnor U12149 (N_12149,N_11582,N_11916);
and U12150 (N_12150,N_11721,N_11622);
nand U12151 (N_12151,N_11873,N_11524);
nand U12152 (N_12152,N_11662,N_11537);
or U12153 (N_12153,N_11979,N_11740);
or U12154 (N_12154,N_11607,N_11862);
nor U12155 (N_12155,N_11939,N_11639);
and U12156 (N_12156,N_11603,N_11759);
nor U12157 (N_12157,N_11754,N_11713);
nor U12158 (N_12158,N_11798,N_11960);
nand U12159 (N_12159,N_11653,N_11532);
nand U12160 (N_12160,N_11643,N_11773);
nand U12161 (N_12161,N_11610,N_11632);
nand U12162 (N_12162,N_11767,N_11644);
and U12163 (N_12163,N_11945,N_11655);
xor U12164 (N_12164,N_11948,N_11878);
nor U12165 (N_12165,N_11870,N_11790);
nor U12166 (N_12166,N_11657,N_11839);
nor U12167 (N_12167,N_11760,N_11557);
nand U12168 (N_12168,N_11877,N_11825);
and U12169 (N_12169,N_11794,N_11797);
or U12170 (N_12170,N_11799,N_11710);
and U12171 (N_12171,N_11667,N_11596);
xnor U12172 (N_12172,N_11943,N_11782);
nor U12173 (N_12173,N_11817,N_11612);
nor U12174 (N_12174,N_11808,N_11719);
nand U12175 (N_12175,N_11833,N_11893);
and U12176 (N_12176,N_11944,N_11999);
nand U12177 (N_12177,N_11539,N_11548);
or U12178 (N_12178,N_11857,N_11894);
nand U12179 (N_12179,N_11933,N_11954);
nand U12180 (N_12180,N_11514,N_11937);
or U12181 (N_12181,N_11989,N_11576);
and U12182 (N_12182,N_11634,N_11803);
nand U12183 (N_12183,N_11957,N_11525);
nor U12184 (N_12184,N_11972,N_11703);
nand U12185 (N_12185,N_11869,N_11895);
and U12186 (N_12186,N_11946,N_11617);
nand U12187 (N_12187,N_11625,N_11854);
nand U12188 (N_12188,N_11699,N_11942);
or U12189 (N_12189,N_11816,N_11822);
or U12190 (N_12190,N_11985,N_11867);
and U12191 (N_12191,N_11813,N_11571);
nor U12192 (N_12192,N_11575,N_11909);
nor U12193 (N_12193,N_11635,N_11889);
and U12194 (N_12194,N_11692,N_11698);
and U12195 (N_12195,N_11627,N_11669);
xor U12196 (N_12196,N_11901,N_11880);
or U12197 (N_12197,N_11636,N_11927);
nor U12198 (N_12198,N_11809,N_11728);
or U12199 (N_12199,N_11528,N_11717);
and U12200 (N_12200,N_11592,N_11788);
nor U12201 (N_12201,N_11802,N_11852);
and U12202 (N_12202,N_11741,N_11861);
nand U12203 (N_12203,N_11774,N_11650);
and U12204 (N_12204,N_11921,N_11775);
and U12205 (N_12205,N_11838,N_11711);
xnor U12206 (N_12206,N_11668,N_11704);
and U12207 (N_12207,N_11828,N_11523);
and U12208 (N_12208,N_11674,N_11856);
xor U12209 (N_12209,N_11572,N_11714);
nand U12210 (N_12210,N_11553,N_11616);
nor U12211 (N_12211,N_11626,N_11580);
nand U12212 (N_12212,N_11736,N_11737);
or U12213 (N_12213,N_11843,N_11876);
or U12214 (N_12214,N_11846,N_11929);
and U12215 (N_12215,N_11795,N_11835);
or U12216 (N_12216,N_11913,N_11920);
nor U12217 (N_12217,N_11595,N_11784);
nor U12218 (N_12218,N_11910,N_11509);
xnor U12219 (N_12219,N_11994,N_11729);
nand U12220 (N_12220,N_11792,N_11682);
xnor U12221 (N_12221,N_11679,N_11805);
nor U12222 (N_12222,N_11733,N_11863);
nand U12223 (N_12223,N_11826,N_11955);
and U12224 (N_12224,N_11919,N_11934);
nor U12225 (N_12225,N_11541,N_11885);
nor U12226 (N_12226,N_11739,N_11966);
nor U12227 (N_12227,N_11832,N_11686);
and U12228 (N_12228,N_11589,N_11984);
nand U12229 (N_12229,N_11738,N_11761);
nand U12230 (N_12230,N_11898,N_11830);
xor U12231 (N_12231,N_11926,N_11591);
nor U12232 (N_12232,N_11872,N_11829);
nor U12233 (N_12233,N_11569,N_11691);
nand U12234 (N_12234,N_11990,N_11749);
or U12235 (N_12235,N_11746,N_11613);
and U12236 (N_12236,N_11995,N_11753);
and U12237 (N_12237,N_11871,N_11820);
nand U12238 (N_12238,N_11967,N_11687);
and U12239 (N_12239,N_11745,N_11641);
and U12240 (N_12240,N_11519,N_11789);
nor U12241 (N_12241,N_11570,N_11510);
or U12242 (N_12242,N_11624,N_11656);
nand U12243 (N_12243,N_11503,N_11855);
nor U12244 (N_12244,N_11932,N_11748);
nor U12245 (N_12245,N_11508,N_11694);
and U12246 (N_12246,N_11819,N_11542);
nand U12247 (N_12247,N_11864,N_11583);
nand U12248 (N_12248,N_11812,N_11996);
nand U12249 (N_12249,N_11646,N_11983);
nor U12250 (N_12250,N_11558,N_11871);
and U12251 (N_12251,N_11630,N_11700);
nand U12252 (N_12252,N_11618,N_11778);
and U12253 (N_12253,N_11736,N_11912);
and U12254 (N_12254,N_11900,N_11500);
nand U12255 (N_12255,N_11809,N_11913);
nor U12256 (N_12256,N_11701,N_11635);
xor U12257 (N_12257,N_11923,N_11716);
nor U12258 (N_12258,N_11770,N_11831);
or U12259 (N_12259,N_11674,N_11861);
or U12260 (N_12260,N_11806,N_11721);
xnor U12261 (N_12261,N_11748,N_11769);
and U12262 (N_12262,N_11542,N_11962);
xnor U12263 (N_12263,N_11975,N_11562);
nor U12264 (N_12264,N_11686,N_11662);
xnor U12265 (N_12265,N_11656,N_11579);
nand U12266 (N_12266,N_11977,N_11776);
and U12267 (N_12267,N_11645,N_11699);
nor U12268 (N_12268,N_11737,N_11742);
or U12269 (N_12269,N_11612,N_11706);
and U12270 (N_12270,N_11620,N_11875);
nor U12271 (N_12271,N_11796,N_11536);
nor U12272 (N_12272,N_11579,N_11631);
nand U12273 (N_12273,N_11987,N_11524);
xnor U12274 (N_12274,N_11564,N_11724);
or U12275 (N_12275,N_11861,N_11717);
or U12276 (N_12276,N_11773,N_11916);
and U12277 (N_12277,N_11512,N_11691);
and U12278 (N_12278,N_11512,N_11880);
nor U12279 (N_12279,N_11874,N_11678);
nand U12280 (N_12280,N_11745,N_11575);
nand U12281 (N_12281,N_11952,N_11586);
nor U12282 (N_12282,N_11631,N_11905);
or U12283 (N_12283,N_11894,N_11924);
xnor U12284 (N_12284,N_11950,N_11841);
and U12285 (N_12285,N_11804,N_11824);
nor U12286 (N_12286,N_11940,N_11738);
xnor U12287 (N_12287,N_11835,N_11712);
nand U12288 (N_12288,N_11961,N_11995);
and U12289 (N_12289,N_11553,N_11860);
or U12290 (N_12290,N_11993,N_11792);
and U12291 (N_12291,N_11971,N_11639);
and U12292 (N_12292,N_11833,N_11540);
nand U12293 (N_12293,N_11755,N_11580);
nor U12294 (N_12294,N_11775,N_11615);
and U12295 (N_12295,N_11698,N_11550);
or U12296 (N_12296,N_11563,N_11653);
or U12297 (N_12297,N_11981,N_11997);
nor U12298 (N_12298,N_11688,N_11557);
and U12299 (N_12299,N_11807,N_11780);
or U12300 (N_12300,N_11926,N_11955);
xor U12301 (N_12301,N_11643,N_11850);
and U12302 (N_12302,N_11681,N_11645);
xor U12303 (N_12303,N_11720,N_11780);
nand U12304 (N_12304,N_11885,N_11743);
and U12305 (N_12305,N_11622,N_11768);
or U12306 (N_12306,N_11875,N_11600);
nand U12307 (N_12307,N_11622,N_11683);
or U12308 (N_12308,N_11692,N_11836);
nor U12309 (N_12309,N_11885,N_11625);
nand U12310 (N_12310,N_11555,N_11838);
nand U12311 (N_12311,N_11877,N_11626);
and U12312 (N_12312,N_11859,N_11598);
or U12313 (N_12313,N_11952,N_11831);
or U12314 (N_12314,N_11814,N_11911);
or U12315 (N_12315,N_11987,N_11756);
nand U12316 (N_12316,N_11813,N_11977);
or U12317 (N_12317,N_11620,N_11721);
and U12318 (N_12318,N_11844,N_11998);
and U12319 (N_12319,N_11957,N_11630);
and U12320 (N_12320,N_11583,N_11522);
or U12321 (N_12321,N_11666,N_11698);
and U12322 (N_12322,N_11949,N_11900);
xnor U12323 (N_12323,N_11777,N_11861);
or U12324 (N_12324,N_11928,N_11865);
and U12325 (N_12325,N_11608,N_11542);
and U12326 (N_12326,N_11950,N_11877);
or U12327 (N_12327,N_11806,N_11893);
nor U12328 (N_12328,N_11788,N_11710);
nand U12329 (N_12329,N_11974,N_11758);
nand U12330 (N_12330,N_11856,N_11711);
xnor U12331 (N_12331,N_11525,N_11990);
nand U12332 (N_12332,N_11500,N_11533);
nand U12333 (N_12333,N_11540,N_11707);
and U12334 (N_12334,N_11818,N_11713);
nor U12335 (N_12335,N_11512,N_11958);
nor U12336 (N_12336,N_11512,N_11993);
or U12337 (N_12337,N_11958,N_11669);
nor U12338 (N_12338,N_11872,N_11667);
nor U12339 (N_12339,N_11953,N_11821);
and U12340 (N_12340,N_11684,N_11750);
and U12341 (N_12341,N_11985,N_11714);
or U12342 (N_12342,N_11874,N_11879);
nor U12343 (N_12343,N_11704,N_11666);
or U12344 (N_12344,N_11545,N_11791);
or U12345 (N_12345,N_11970,N_11840);
or U12346 (N_12346,N_11703,N_11647);
or U12347 (N_12347,N_11823,N_11511);
and U12348 (N_12348,N_11875,N_11659);
nand U12349 (N_12349,N_11774,N_11500);
and U12350 (N_12350,N_11548,N_11734);
and U12351 (N_12351,N_11815,N_11731);
nand U12352 (N_12352,N_11711,N_11914);
nand U12353 (N_12353,N_11749,N_11800);
and U12354 (N_12354,N_11713,N_11723);
nand U12355 (N_12355,N_11826,N_11881);
or U12356 (N_12356,N_11541,N_11802);
or U12357 (N_12357,N_11829,N_11562);
and U12358 (N_12358,N_11997,N_11770);
or U12359 (N_12359,N_11947,N_11573);
and U12360 (N_12360,N_11646,N_11514);
nor U12361 (N_12361,N_11750,N_11813);
or U12362 (N_12362,N_11763,N_11558);
nand U12363 (N_12363,N_11825,N_11991);
and U12364 (N_12364,N_11854,N_11609);
and U12365 (N_12365,N_11609,N_11624);
or U12366 (N_12366,N_11551,N_11866);
nor U12367 (N_12367,N_11756,N_11894);
and U12368 (N_12368,N_11525,N_11550);
nor U12369 (N_12369,N_11517,N_11700);
or U12370 (N_12370,N_11560,N_11792);
xnor U12371 (N_12371,N_11761,N_11874);
and U12372 (N_12372,N_11713,N_11533);
or U12373 (N_12373,N_11657,N_11607);
or U12374 (N_12374,N_11753,N_11947);
or U12375 (N_12375,N_11592,N_11528);
or U12376 (N_12376,N_11574,N_11625);
or U12377 (N_12377,N_11958,N_11746);
nor U12378 (N_12378,N_11987,N_11924);
or U12379 (N_12379,N_11646,N_11811);
nand U12380 (N_12380,N_11869,N_11965);
or U12381 (N_12381,N_11648,N_11782);
or U12382 (N_12382,N_11707,N_11931);
nor U12383 (N_12383,N_11547,N_11852);
or U12384 (N_12384,N_11657,N_11761);
nor U12385 (N_12385,N_11754,N_11938);
nand U12386 (N_12386,N_11941,N_11510);
or U12387 (N_12387,N_11813,N_11693);
or U12388 (N_12388,N_11646,N_11952);
xor U12389 (N_12389,N_11646,N_11889);
nand U12390 (N_12390,N_11874,N_11579);
nor U12391 (N_12391,N_11863,N_11987);
or U12392 (N_12392,N_11777,N_11907);
or U12393 (N_12393,N_11895,N_11718);
nand U12394 (N_12394,N_11759,N_11987);
xnor U12395 (N_12395,N_11704,N_11937);
nand U12396 (N_12396,N_11977,N_11985);
nand U12397 (N_12397,N_11532,N_11764);
and U12398 (N_12398,N_11938,N_11689);
or U12399 (N_12399,N_11918,N_11594);
nand U12400 (N_12400,N_11505,N_11977);
and U12401 (N_12401,N_11684,N_11930);
nor U12402 (N_12402,N_11644,N_11699);
and U12403 (N_12403,N_11909,N_11876);
and U12404 (N_12404,N_11688,N_11566);
xor U12405 (N_12405,N_11807,N_11854);
and U12406 (N_12406,N_11904,N_11823);
and U12407 (N_12407,N_11546,N_11986);
xnor U12408 (N_12408,N_11928,N_11842);
nand U12409 (N_12409,N_11854,N_11864);
nand U12410 (N_12410,N_11966,N_11845);
nor U12411 (N_12411,N_11994,N_11548);
nand U12412 (N_12412,N_11937,N_11763);
nand U12413 (N_12413,N_11609,N_11706);
or U12414 (N_12414,N_11948,N_11581);
or U12415 (N_12415,N_11917,N_11752);
and U12416 (N_12416,N_11542,N_11890);
nand U12417 (N_12417,N_11510,N_11560);
and U12418 (N_12418,N_11768,N_11934);
and U12419 (N_12419,N_11838,N_11953);
or U12420 (N_12420,N_11905,N_11972);
nor U12421 (N_12421,N_11700,N_11645);
or U12422 (N_12422,N_11941,N_11642);
nor U12423 (N_12423,N_11556,N_11661);
nand U12424 (N_12424,N_11806,N_11700);
and U12425 (N_12425,N_11779,N_11964);
or U12426 (N_12426,N_11536,N_11630);
nor U12427 (N_12427,N_11697,N_11905);
or U12428 (N_12428,N_11883,N_11703);
or U12429 (N_12429,N_11661,N_11574);
and U12430 (N_12430,N_11904,N_11789);
nor U12431 (N_12431,N_11783,N_11514);
xor U12432 (N_12432,N_11875,N_11907);
and U12433 (N_12433,N_11823,N_11745);
and U12434 (N_12434,N_11556,N_11500);
or U12435 (N_12435,N_11644,N_11806);
xnor U12436 (N_12436,N_11853,N_11509);
or U12437 (N_12437,N_11722,N_11867);
nand U12438 (N_12438,N_11786,N_11822);
nor U12439 (N_12439,N_11662,N_11606);
and U12440 (N_12440,N_11560,N_11953);
and U12441 (N_12441,N_11732,N_11931);
xnor U12442 (N_12442,N_11684,N_11759);
and U12443 (N_12443,N_11558,N_11844);
or U12444 (N_12444,N_11717,N_11702);
nor U12445 (N_12445,N_11945,N_11763);
nand U12446 (N_12446,N_11661,N_11929);
and U12447 (N_12447,N_11771,N_11529);
and U12448 (N_12448,N_11711,N_11720);
nor U12449 (N_12449,N_11998,N_11681);
nor U12450 (N_12450,N_11642,N_11644);
or U12451 (N_12451,N_11753,N_11615);
or U12452 (N_12452,N_11612,N_11988);
or U12453 (N_12453,N_11990,N_11790);
nor U12454 (N_12454,N_11889,N_11724);
xnor U12455 (N_12455,N_11668,N_11957);
nor U12456 (N_12456,N_11759,N_11931);
or U12457 (N_12457,N_11954,N_11916);
nand U12458 (N_12458,N_11676,N_11756);
xor U12459 (N_12459,N_11933,N_11791);
nand U12460 (N_12460,N_11855,N_11526);
xor U12461 (N_12461,N_11948,N_11819);
nor U12462 (N_12462,N_11708,N_11939);
nand U12463 (N_12463,N_11916,N_11619);
xnor U12464 (N_12464,N_11556,N_11939);
or U12465 (N_12465,N_11665,N_11626);
nor U12466 (N_12466,N_11874,N_11684);
nand U12467 (N_12467,N_11731,N_11561);
nor U12468 (N_12468,N_11938,N_11597);
and U12469 (N_12469,N_11570,N_11894);
nor U12470 (N_12470,N_11635,N_11755);
xor U12471 (N_12471,N_11793,N_11750);
and U12472 (N_12472,N_11621,N_11830);
or U12473 (N_12473,N_11691,N_11575);
nand U12474 (N_12474,N_11809,N_11617);
nand U12475 (N_12475,N_11881,N_11988);
nand U12476 (N_12476,N_11757,N_11519);
nor U12477 (N_12477,N_11868,N_11559);
nor U12478 (N_12478,N_11550,N_11569);
or U12479 (N_12479,N_11819,N_11962);
nor U12480 (N_12480,N_11866,N_11936);
nor U12481 (N_12481,N_11559,N_11618);
or U12482 (N_12482,N_11748,N_11922);
nand U12483 (N_12483,N_11655,N_11917);
nand U12484 (N_12484,N_11751,N_11868);
and U12485 (N_12485,N_11584,N_11751);
or U12486 (N_12486,N_11679,N_11519);
nor U12487 (N_12487,N_11849,N_11584);
and U12488 (N_12488,N_11727,N_11707);
nor U12489 (N_12489,N_11762,N_11955);
nor U12490 (N_12490,N_11587,N_11570);
and U12491 (N_12491,N_11869,N_11979);
xor U12492 (N_12492,N_11583,N_11671);
nor U12493 (N_12493,N_11626,N_11841);
or U12494 (N_12494,N_11770,N_11830);
or U12495 (N_12495,N_11718,N_11698);
and U12496 (N_12496,N_11582,N_11744);
and U12497 (N_12497,N_11798,N_11993);
nor U12498 (N_12498,N_11650,N_11875);
and U12499 (N_12499,N_11524,N_11559);
xnor U12500 (N_12500,N_12169,N_12197);
nor U12501 (N_12501,N_12287,N_12058);
nand U12502 (N_12502,N_12032,N_12281);
or U12503 (N_12503,N_12418,N_12141);
nand U12504 (N_12504,N_12127,N_12385);
and U12505 (N_12505,N_12095,N_12426);
or U12506 (N_12506,N_12099,N_12056);
nand U12507 (N_12507,N_12015,N_12443);
nand U12508 (N_12508,N_12463,N_12157);
nand U12509 (N_12509,N_12152,N_12117);
or U12510 (N_12510,N_12017,N_12452);
or U12511 (N_12511,N_12175,N_12033);
nand U12512 (N_12512,N_12469,N_12492);
and U12513 (N_12513,N_12499,N_12277);
or U12514 (N_12514,N_12477,N_12417);
or U12515 (N_12515,N_12147,N_12489);
and U12516 (N_12516,N_12104,N_12215);
and U12517 (N_12517,N_12007,N_12172);
or U12518 (N_12518,N_12202,N_12332);
nor U12519 (N_12519,N_12374,N_12247);
nor U12520 (N_12520,N_12055,N_12466);
or U12521 (N_12521,N_12128,N_12305);
and U12522 (N_12522,N_12438,N_12069);
nor U12523 (N_12523,N_12023,N_12354);
or U12524 (N_12524,N_12176,N_12498);
or U12525 (N_12525,N_12073,N_12491);
nand U12526 (N_12526,N_12327,N_12266);
and U12527 (N_12527,N_12401,N_12410);
nor U12528 (N_12528,N_12301,N_12420);
nand U12529 (N_12529,N_12046,N_12047);
or U12530 (N_12530,N_12029,N_12375);
nor U12531 (N_12531,N_12282,N_12143);
nor U12532 (N_12532,N_12276,N_12286);
and U12533 (N_12533,N_12495,N_12166);
and U12534 (N_12534,N_12138,N_12204);
or U12535 (N_12535,N_12363,N_12014);
nor U12536 (N_12536,N_12398,N_12206);
or U12537 (N_12537,N_12064,N_12432);
and U12538 (N_12538,N_12107,N_12246);
or U12539 (N_12539,N_12352,N_12037);
xnor U12540 (N_12540,N_12124,N_12254);
xnor U12541 (N_12541,N_12004,N_12194);
nor U12542 (N_12542,N_12497,N_12292);
xnor U12543 (N_12543,N_12271,N_12231);
nor U12544 (N_12544,N_12457,N_12181);
nor U12545 (N_12545,N_12249,N_12041);
nor U12546 (N_12546,N_12485,N_12284);
and U12547 (N_12547,N_12255,N_12446);
or U12548 (N_12548,N_12232,N_12154);
or U12549 (N_12549,N_12395,N_12196);
nor U12550 (N_12550,N_12326,N_12380);
nor U12551 (N_12551,N_12217,N_12031);
nand U12552 (N_12552,N_12061,N_12170);
or U12553 (N_12553,N_12010,N_12065);
and U12554 (N_12554,N_12213,N_12212);
nand U12555 (N_12555,N_12184,N_12221);
nand U12556 (N_12556,N_12296,N_12040);
xnor U12557 (N_12557,N_12075,N_12229);
xor U12558 (N_12558,N_12342,N_12150);
and U12559 (N_12559,N_12323,N_12289);
nor U12560 (N_12560,N_12487,N_12209);
nand U12561 (N_12561,N_12222,N_12114);
nor U12562 (N_12562,N_12449,N_12280);
xnor U12563 (N_12563,N_12011,N_12049);
nor U12564 (N_12564,N_12161,N_12230);
or U12565 (N_12565,N_12084,N_12493);
or U12566 (N_12566,N_12216,N_12074);
and U12567 (N_12567,N_12088,N_12465);
nand U12568 (N_12568,N_12076,N_12153);
xor U12569 (N_12569,N_12298,N_12470);
nor U12570 (N_12570,N_12399,N_12311);
xor U12571 (N_12571,N_12475,N_12260);
nor U12572 (N_12572,N_12455,N_12402);
and U12573 (N_12573,N_12494,N_12244);
or U12574 (N_12574,N_12453,N_12111);
xnor U12575 (N_12575,N_12490,N_12207);
nor U12576 (N_12576,N_12427,N_12362);
and U12577 (N_12577,N_12471,N_12331);
xor U12578 (N_12578,N_12191,N_12038);
nand U12579 (N_12579,N_12094,N_12087);
or U12580 (N_12580,N_12283,N_12123);
nor U12581 (N_12581,N_12434,N_12057);
nor U12582 (N_12582,N_12134,N_12310);
and U12583 (N_12583,N_12376,N_12160);
and U12584 (N_12584,N_12378,N_12383);
or U12585 (N_12585,N_12145,N_12067);
and U12586 (N_12586,N_12177,N_12256);
and U12587 (N_12587,N_12386,N_12109);
xor U12588 (N_12588,N_12297,N_12198);
nand U12589 (N_12589,N_12448,N_12328);
nand U12590 (N_12590,N_12472,N_12396);
nand U12591 (N_12591,N_12481,N_12042);
nor U12592 (N_12592,N_12101,N_12220);
nor U12593 (N_12593,N_12414,N_12190);
nand U12594 (N_12594,N_12113,N_12339);
or U12595 (N_12595,N_12462,N_12313);
nor U12596 (N_12596,N_12192,N_12008);
and U12597 (N_12597,N_12345,N_12158);
or U12598 (N_12598,N_12373,N_12259);
xnor U12599 (N_12599,N_12050,N_12388);
or U12600 (N_12600,N_12369,N_12164);
nand U12601 (N_12601,N_12187,N_12009);
nand U12602 (N_12602,N_12096,N_12408);
and U12603 (N_12603,N_12422,N_12146);
and U12604 (N_12604,N_12351,N_12306);
nand U12605 (N_12605,N_12319,N_12291);
nor U12606 (N_12606,N_12110,N_12350);
xor U12607 (N_12607,N_12450,N_12431);
nand U12608 (N_12608,N_12261,N_12242);
nand U12609 (N_12609,N_12288,N_12098);
xnor U12610 (N_12610,N_12295,N_12149);
and U12611 (N_12611,N_12265,N_12337);
xor U12612 (N_12612,N_12083,N_12182);
or U12613 (N_12613,N_12129,N_12173);
nor U12614 (N_12614,N_12444,N_12001);
nor U12615 (N_12615,N_12257,N_12341);
nand U12616 (N_12616,N_12137,N_12248);
nand U12617 (N_12617,N_12131,N_12382);
xor U12618 (N_12618,N_12142,N_12348);
and U12619 (N_12619,N_12413,N_12468);
nand U12620 (N_12620,N_12361,N_12241);
or U12621 (N_12621,N_12312,N_12294);
or U12622 (N_12622,N_12189,N_12002);
nor U12623 (N_12623,N_12325,N_12245);
or U12624 (N_12624,N_12316,N_12405);
nand U12625 (N_12625,N_12132,N_12372);
and U12626 (N_12626,N_12392,N_12022);
nand U12627 (N_12627,N_12018,N_12224);
and U12628 (N_12628,N_12479,N_12252);
and U12629 (N_12629,N_12262,N_12130);
nand U12630 (N_12630,N_12384,N_12437);
and U12631 (N_12631,N_12112,N_12293);
or U12632 (N_12632,N_12278,N_12336);
nand U12633 (N_12633,N_12307,N_12424);
nor U12634 (N_12634,N_12218,N_12086);
or U12635 (N_12635,N_12344,N_12126);
and U12636 (N_12636,N_12379,N_12148);
nand U12637 (N_12637,N_12121,N_12115);
nor U12638 (N_12638,N_12406,N_12179);
nand U12639 (N_12639,N_12108,N_12488);
nor U12640 (N_12640,N_12188,N_12024);
and U12641 (N_12641,N_12070,N_12279);
nand U12642 (N_12642,N_12394,N_12483);
nor U12643 (N_12643,N_12353,N_12036);
or U12644 (N_12644,N_12482,N_12054);
or U12645 (N_12645,N_12144,N_12000);
or U12646 (N_12646,N_12080,N_12407);
or U12647 (N_12647,N_12235,N_12303);
xor U12648 (N_12648,N_12030,N_12026);
and U12649 (N_12649,N_12411,N_12440);
and U12650 (N_12650,N_12005,N_12155);
and U12651 (N_12651,N_12251,N_12068);
nand U12652 (N_12652,N_12397,N_12151);
nor U12653 (N_12653,N_12458,N_12447);
and U12654 (N_12654,N_12039,N_12016);
xnor U12655 (N_12655,N_12171,N_12051);
nor U12656 (N_12656,N_12035,N_12300);
xnor U12657 (N_12657,N_12228,N_12178);
nor U12658 (N_12658,N_12356,N_12315);
and U12659 (N_12659,N_12347,N_12208);
nand U12660 (N_12660,N_12393,N_12106);
xor U12661 (N_12661,N_12210,N_12243);
or U12662 (N_12662,N_12340,N_12006);
or U12663 (N_12663,N_12233,N_12273);
and U12664 (N_12664,N_12140,N_12239);
or U12665 (N_12665,N_12486,N_12193);
nand U12666 (N_12666,N_12335,N_12387);
nor U12667 (N_12667,N_12441,N_12371);
or U12668 (N_12668,N_12250,N_12180);
nand U12669 (N_12669,N_12390,N_12118);
nand U12670 (N_12670,N_12072,N_12333);
nor U12671 (N_12671,N_12429,N_12122);
xnor U12672 (N_12672,N_12034,N_12476);
or U12673 (N_12673,N_12360,N_12451);
nand U12674 (N_12674,N_12219,N_12227);
or U12675 (N_12675,N_12366,N_12381);
nand U12676 (N_12676,N_12060,N_12105);
and U12677 (N_12677,N_12013,N_12019);
nand U12678 (N_12678,N_12093,N_12174);
nor U12679 (N_12679,N_12419,N_12162);
nand U12680 (N_12680,N_12433,N_12200);
and U12681 (N_12681,N_12133,N_12454);
and U12682 (N_12682,N_12400,N_12048);
xnor U12683 (N_12683,N_12436,N_12346);
and U12684 (N_12684,N_12139,N_12199);
or U12685 (N_12685,N_12357,N_12053);
nand U12686 (N_12686,N_12045,N_12082);
or U12687 (N_12687,N_12163,N_12059);
or U12688 (N_12688,N_12355,N_12090);
xnor U12689 (N_12689,N_12478,N_12321);
xor U12690 (N_12690,N_12268,N_12135);
or U12691 (N_12691,N_12195,N_12214);
or U12692 (N_12692,N_12116,N_12364);
nor U12693 (N_12693,N_12183,N_12238);
nand U12694 (N_12694,N_12125,N_12275);
and U12695 (N_12695,N_12304,N_12423);
xnor U12696 (N_12696,N_12085,N_12272);
and U12697 (N_12697,N_12021,N_12412);
or U12698 (N_12698,N_12338,N_12322);
xor U12699 (N_12699,N_12120,N_12027);
nor U12700 (N_12700,N_12003,N_12415);
nand U12701 (N_12701,N_12091,N_12156);
nor U12702 (N_12702,N_12302,N_12028);
or U12703 (N_12703,N_12225,N_12044);
nand U12704 (N_12704,N_12079,N_12285);
nor U12705 (N_12705,N_12185,N_12459);
and U12706 (N_12706,N_12203,N_12349);
or U12707 (N_12707,N_12223,N_12226);
nor U12708 (N_12708,N_12403,N_12205);
nor U12709 (N_12709,N_12370,N_12445);
nor U12710 (N_12710,N_12168,N_12416);
xor U12711 (N_12711,N_12330,N_12308);
nand U12712 (N_12712,N_12211,N_12329);
xor U12713 (N_12713,N_12167,N_12267);
and U12714 (N_12714,N_12234,N_12314);
nor U12715 (N_12715,N_12456,N_12464);
xor U12716 (N_12716,N_12263,N_12043);
or U12717 (N_12717,N_12428,N_12062);
or U12718 (N_12718,N_12081,N_12421);
nand U12719 (N_12719,N_12290,N_12439);
and U12720 (N_12720,N_12136,N_12186);
nor U12721 (N_12721,N_12430,N_12102);
nor U12722 (N_12722,N_12442,N_12474);
and U12723 (N_12723,N_12320,N_12324);
xnor U12724 (N_12724,N_12391,N_12343);
or U12725 (N_12725,N_12367,N_12359);
nor U12726 (N_12726,N_12063,N_12496);
xor U12727 (N_12727,N_12240,N_12460);
nand U12728 (N_12728,N_12020,N_12365);
xor U12729 (N_12729,N_12409,N_12269);
nand U12730 (N_12730,N_12461,N_12377);
and U12731 (N_12731,N_12025,N_12258);
xnor U12732 (N_12732,N_12066,N_12012);
nor U12733 (N_12733,N_12264,N_12368);
and U12734 (N_12734,N_12274,N_12480);
xnor U12735 (N_12735,N_12201,N_12425);
and U12736 (N_12736,N_12484,N_12165);
and U12737 (N_12737,N_12077,N_12334);
and U12738 (N_12738,N_12389,N_12159);
nor U12739 (N_12739,N_12071,N_12309);
nor U12740 (N_12740,N_12270,N_12435);
nor U12741 (N_12741,N_12404,N_12237);
nor U12742 (N_12742,N_12119,N_12467);
and U12743 (N_12743,N_12317,N_12100);
xnor U12744 (N_12744,N_12236,N_12318);
nand U12745 (N_12745,N_12103,N_12299);
nor U12746 (N_12746,N_12253,N_12097);
and U12747 (N_12747,N_12052,N_12358);
xor U12748 (N_12748,N_12078,N_12089);
xnor U12749 (N_12749,N_12092,N_12473);
nor U12750 (N_12750,N_12100,N_12174);
nand U12751 (N_12751,N_12053,N_12242);
or U12752 (N_12752,N_12105,N_12206);
nand U12753 (N_12753,N_12079,N_12016);
or U12754 (N_12754,N_12005,N_12069);
nor U12755 (N_12755,N_12362,N_12235);
or U12756 (N_12756,N_12463,N_12081);
nand U12757 (N_12757,N_12154,N_12053);
xnor U12758 (N_12758,N_12286,N_12064);
and U12759 (N_12759,N_12023,N_12416);
and U12760 (N_12760,N_12295,N_12409);
nand U12761 (N_12761,N_12129,N_12433);
nand U12762 (N_12762,N_12257,N_12499);
and U12763 (N_12763,N_12084,N_12051);
or U12764 (N_12764,N_12266,N_12320);
and U12765 (N_12765,N_12008,N_12332);
or U12766 (N_12766,N_12387,N_12188);
xor U12767 (N_12767,N_12150,N_12195);
xnor U12768 (N_12768,N_12185,N_12483);
and U12769 (N_12769,N_12351,N_12244);
nand U12770 (N_12770,N_12013,N_12364);
nor U12771 (N_12771,N_12349,N_12386);
or U12772 (N_12772,N_12048,N_12011);
nor U12773 (N_12773,N_12000,N_12481);
and U12774 (N_12774,N_12371,N_12167);
xor U12775 (N_12775,N_12147,N_12152);
nand U12776 (N_12776,N_12493,N_12134);
and U12777 (N_12777,N_12132,N_12111);
nand U12778 (N_12778,N_12064,N_12208);
or U12779 (N_12779,N_12406,N_12414);
or U12780 (N_12780,N_12071,N_12364);
nor U12781 (N_12781,N_12179,N_12245);
nand U12782 (N_12782,N_12156,N_12194);
and U12783 (N_12783,N_12478,N_12213);
xor U12784 (N_12784,N_12299,N_12224);
nand U12785 (N_12785,N_12404,N_12221);
nor U12786 (N_12786,N_12332,N_12281);
or U12787 (N_12787,N_12063,N_12221);
nor U12788 (N_12788,N_12182,N_12261);
nor U12789 (N_12789,N_12405,N_12469);
nor U12790 (N_12790,N_12079,N_12431);
nor U12791 (N_12791,N_12318,N_12329);
or U12792 (N_12792,N_12406,N_12028);
nand U12793 (N_12793,N_12340,N_12195);
or U12794 (N_12794,N_12317,N_12352);
nand U12795 (N_12795,N_12335,N_12481);
or U12796 (N_12796,N_12004,N_12329);
and U12797 (N_12797,N_12098,N_12265);
and U12798 (N_12798,N_12433,N_12046);
and U12799 (N_12799,N_12309,N_12297);
and U12800 (N_12800,N_12340,N_12178);
or U12801 (N_12801,N_12349,N_12048);
nand U12802 (N_12802,N_12007,N_12493);
nor U12803 (N_12803,N_12300,N_12468);
nor U12804 (N_12804,N_12066,N_12165);
xnor U12805 (N_12805,N_12021,N_12451);
or U12806 (N_12806,N_12373,N_12240);
nand U12807 (N_12807,N_12276,N_12339);
xnor U12808 (N_12808,N_12212,N_12123);
nor U12809 (N_12809,N_12041,N_12494);
nand U12810 (N_12810,N_12208,N_12074);
xor U12811 (N_12811,N_12197,N_12361);
nand U12812 (N_12812,N_12212,N_12446);
nand U12813 (N_12813,N_12189,N_12190);
nor U12814 (N_12814,N_12026,N_12219);
nand U12815 (N_12815,N_12454,N_12219);
or U12816 (N_12816,N_12322,N_12231);
nand U12817 (N_12817,N_12301,N_12144);
nor U12818 (N_12818,N_12107,N_12422);
or U12819 (N_12819,N_12144,N_12084);
or U12820 (N_12820,N_12330,N_12415);
nand U12821 (N_12821,N_12275,N_12176);
or U12822 (N_12822,N_12047,N_12358);
or U12823 (N_12823,N_12320,N_12433);
nand U12824 (N_12824,N_12438,N_12370);
nand U12825 (N_12825,N_12027,N_12336);
xnor U12826 (N_12826,N_12087,N_12211);
nand U12827 (N_12827,N_12125,N_12141);
nor U12828 (N_12828,N_12093,N_12300);
or U12829 (N_12829,N_12012,N_12176);
nor U12830 (N_12830,N_12174,N_12378);
nor U12831 (N_12831,N_12387,N_12223);
and U12832 (N_12832,N_12205,N_12429);
or U12833 (N_12833,N_12140,N_12355);
and U12834 (N_12834,N_12032,N_12310);
xor U12835 (N_12835,N_12194,N_12226);
nor U12836 (N_12836,N_12244,N_12282);
or U12837 (N_12837,N_12284,N_12460);
nor U12838 (N_12838,N_12245,N_12233);
nand U12839 (N_12839,N_12437,N_12203);
and U12840 (N_12840,N_12342,N_12086);
and U12841 (N_12841,N_12184,N_12002);
nor U12842 (N_12842,N_12419,N_12085);
xor U12843 (N_12843,N_12459,N_12449);
xor U12844 (N_12844,N_12092,N_12470);
nor U12845 (N_12845,N_12210,N_12327);
nand U12846 (N_12846,N_12027,N_12059);
or U12847 (N_12847,N_12278,N_12040);
or U12848 (N_12848,N_12421,N_12356);
nand U12849 (N_12849,N_12187,N_12339);
nand U12850 (N_12850,N_12143,N_12087);
or U12851 (N_12851,N_12219,N_12421);
or U12852 (N_12852,N_12493,N_12165);
xnor U12853 (N_12853,N_12145,N_12030);
or U12854 (N_12854,N_12029,N_12118);
or U12855 (N_12855,N_12128,N_12042);
nand U12856 (N_12856,N_12128,N_12279);
and U12857 (N_12857,N_12437,N_12147);
or U12858 (N_12858,N_12483,N_12322);
and U12859 (N_12859,N_12296,N_12021);
nand U12860 (N_12860,N_12472,N_12087);
nand U12861 (N_12861,N_12053,N_12360);
nor U12862 (N_12862,N_12087,N_12249);
xnor U12863 (N_12863,N_12269,N_12443);
nor U12864 (N_12864,N_12067,N_12438);
nand U12865 (N_12865,N_12150,N_12044);
xnor U12866 (N_12866,N_12458,N_12364);
and U12867 (N_12867,N_12116,N_12064);
and U12868 (N_12868,N_12308,N_12167);
xor U12869 (N_12869,N_12170,N_12480);
nand U12870 (N_12870,N_12024,N_12339);
and U12871 (N_12871,N_12321,N_12296);
nand U12872 (N_12872,N_12053,N_12008);
nand U12873 (N_12873,N_12123,N_12095);
and U12874 (N_12874,N_12199,N_12244);
or U12875 (N_12875,N_12295,N_12043);
and U12876 (N_12876,N_12163,N_12453);
or U12877 (N_12877,N_12092,N_12004);
nand U12878 (N_12878,N_12134,N_12127);
and U12879 (N_12879,N_12063,N_12045);
nand U12880 (N_12880,N_12229,N_12248);
nor U12881 (N_12881,N_12465,N_12314);
xnor U12882 (N_12882,N_12269,N_12414);
and U12883 (N_12883,N_12319,N_12463);
or U12884 (N_12884,N_12099,N_12185);
nor U12885 (N_12885,N_12045,N_12130);
nor U12886 (N_12886,N_12160,N_12471);
and U12887 (N_12887,N_12293,N_12075);
nand U12888 (N_12888,N_12130,N_12021);
xnor U12889 (N_12889,N_12104,N_12125);
and U12890 (N_12890,N_12157,N_12119);
or U12891 (N_12891,N_12395,N_12379);
xor U12892 (N_12892,N_12280,N_12300);
xor U12893 (N_12893,N_12227,N_12037);
and U12894 (N_12894,N_12104,N_12221);
nand U12895 (N_12895,N_12411,N_12259);
or U12896 (N_12896,N_12457,N_12012);
and U12897 (N_12897,N_12282,N_12121);
and U12898 (N_12898,N_12389,N_12037);
nand U12899 (N_12899,N_12210,N_12445);
nand U12900 (N_12900,N_12474,N_12493);
xor U12901 (N_12901,N_12283,N_12128);
xor U12902 (N_12902,N_12153,N_12315);
xor U12903 (N_12903,N_12083,N_12348);
nand U12904 (N_12904,N_12064,N_12086);
xor U12905 (N_12905,N_12126,N_12444);
or U12906 (N_12906,N_12087,N_12017);
or U12907 (N_12907,N_12463,N_12031);
nand U12908 (N_12908,N_12404,N_12045);
nor U12909 (N_12909,N_12463,N_12411);
and U12910 (N_12910,N_12453,N_12052);
nor U12911 (N_12911,N_12113,N_12420);
nand U12912 (N_12912,N_12443,N_12291);
nor U12913 (N_12913,N_12485,N_12033);
and U12914 (N_12914,N_12332,N_12183);
nor U12915 (N_12915,N_12341,N_12134);
or U12916 (N_12916,N_12362,N_12426);
and U12917 (N_12917,N_12208,N_12466);
nor U12918 (N_12918,N_12145,N_12453);
nor U12919 (N_12919,N_12047,N_12408);
or U12920 (N_12920,N_12134,N_12183);
xnor U12921 (N_12921,N_12125,N_12419);
xnor U12922 (N_12922,N_12007,N_12490);
or U12923 (N_12923,N_12170,N_12473);
or U12924 (N_12924,N_12199,N_12266);
and U12925 (N_12925,N_12371,N_12214);
nor U12926 (N_12926,N_12125,N_12011);
nand U12927 (N_12927,N_12223,N_12228);
and U12928 (N_12928,N_12136,N_12203);
nand U12929 (N_12929,N_12258,N_12196);
and U12930 (N_12930,N_12364,N_12267);
or U12931 (N_12931,N_12012,N_12438);
nand U12932 (N_12932,N_12452,N_12485);
xor U12933 (N_12933,N_12467,N_12470);
and U12934 (N_12934,N_12149,N_12202);
or U12935 (N_12935,N_12441,N_12151);
nor U12936 (N_12936,N_12175,N_12140);
or U12937 (N_12937,N_12494,N_12419);
nor U12938 (N_12938,N_12262,N_12307);
or U12939 (N_12939,N_12278,N_12356);
and U12940 (N_12940,N_12467,N_12013);
nor U12941 (N_12941,N_12069,N_12394);
xor U12942 (N_12942,N_12344,N_12230);
xnor U12943 (N_12943,N_12487,N_12218);
xnor U12944 (N_12944,N_12354,N_12252);
and U12945 (N_12945,N_12055,N_12468);
xnor U12946 (N_12946,N_12063,N_12182);
xor U12947 (N_12947,N_12014,N_12007);
or U12948 (N_12948,N_12078,N_12151);
nand U12949 (N_12949,N_12189,N_12066);
nor U12950 (N_12950,N_12066,N_12441);
nand U12951 (N_12951,N_12399,N_12305);
and U12952 (N_12952,N_12248,N_12425);
and U12953 (N_12953,N_12066,N_12427);
nor U12954 (N_12954,N_12260,N_12112);
or U12955 (N_12955,N_12128,N_12011);
nor U12956 (N_12956,N_12135,N_12465);
or U12957 (N_12957,N_12114,N_12412);
nand U12958 (N_12958,N_12209,N_12289);
nor U12959 (N_12959,N_12263,N_12030);
or U12960 (N_12960,N_12237,N_12346);
nor U12961 (N_12961,N_12117,N_12268);
or U12962 (N_12962,N_12377,N_12234);
nand U12963 (N_12963,N_12163,N_12049);
or U12964 (N_12964,N_12148,N_12146);
or U12965 (N_12965,N_12439,N_12209);
nor U12966 (N_12966,N_12304,N_12426);
or U12967 (N_12967,N_12222,N_12333);
or U12968 (N_12968,N_12336,N_12296);
or U12969 (N_12969,N_12457,N_12162);
nand U12970 (N_12970,N_12196,N_12282);
nand U12971 (N_12971,N_12461,N_12436);
nor U12972 (N_12972,N_12423,N_12229);
or U12973 (N_12973,N_12258,N_12233);
nor U12974 (N_12974,N_12413,N_12291);
xnor U12975 (N_12975,N_12391,N_12213);
or U12976 (N_12976,N_12498,N_12072);
or U12977 (N_12977,N_12370,N_12243);
and U12978 (N_12978,N_12455,N_12456);
and U12979 (N_12979,N_12318,N_12460);
and U12980 (N_12980,N_12323,N_12370);
nand U12981 (N_12981,N_12138,N_12222);
nand U12982 (N_12982,N_12274,N_12465);
and U12983 (N_12983,N_12369,N_12102);
or U12984 (N_12984,N_12012,N_12390);
or U12985 (N_12985,N_12251,N_12238);
nor U12986 (N_12986,N_12083,N_12086);
nor U12987 (N_12987,N_12471,N_12322);
and U12988 (N_12988,N_12297,N_12386);
or U12989 (N_12989,N_12380,N_12254);
or U12990 (N_12990,N_12113,N_12128);
and U12991 (N_12991,N_12139,N_12441);
or U12992 (N_12992,N_12098,N_12020);
nor U12993 (N_12993,N_12125,N_12071);
or U12994 (N_12994,N_12192,N_12480);
or U12995 (N_12995,N_12329,N_12226);
or U12996 (N_12996,N_12287,N_12486);
or U12997 (N_12997,N_12343,N_12120);
and U12998 (N_12998,N_12242,N_12097);
and U12999 (N_12999,N_12335,N_12415);
or U13000 (N_13000,N_12815,N_12632);
or U13001 (N_13001,N_12829,N_12714);
nand U13002 (N_13002,N_12669,N_12513);
or U13003 (N_13003,N_12610,N_12793);
xor U13004 (N_13004,N_12656,N_12700);
nand U13005 (N_13005,N_12986,N_12678);
and U13006 (N_13006,N_12847,N_12653);
or U13007 (N_13007,N_12781,N_12764);
or U13008 (N_13008,N_12587,N_12926);
and U13009 (N_13009,N_12701,N_12756);
nand U13010 (N_13010,N_12534,N_12602);
nor U13011 (N_13011,N_12642,N_12834);
or U13012 (N_13012,N_12574,N_12524);
and U13013 (N_13013,N_12579,N_12915);
or U13014 (N_13014,N_12633,N_12510);
xnor U13015 (N_13015,N_12641,N_12564);
or U13016 (N_13016,N_12997,N_12825);
or U13017 (N_13017,N_12888,N_12739);
or U13018 (N_13018,N_12902,N_12505);
nor U13019 (N_13019,N_12529,N_12725);
nand U13020 (N_13020,N_12999,N_12917);
or U13021 (N_13021,N_12639,N_12812);
nor U13022 (N_13022,N_12874,N_12811);
and U13023 (N_13023,N_12856,N_12891);
nand U13024 (N_13024,N_12671,N_12877);
or U13025 (N_13025,N_12692,N_12704);
and U13026 (N_13026,N_12777,N_12672);
or U13027 (N_13027,N_12562,N_12711);
or U13028 (N_13028,N_12814,N_12964);
nor U13029 (N_13029,N_12664,N_12567);
or U13030 (N_13030,N_12951,N_12962);
or U13031 (N_13031,N_12901,N_12861);
nor U13032 (N_13032,N_12988,N_12707);
and U13033 (N_13033,N_12979,N_12963);
and U13034 (N_13034,N_12871,N_12985);
and U13035 (N_13035,N_12643,N_12712);
and U13036 (N_13036,N_12740,N_12994);
nor U13037 (N_13037,N_12517,N_12876);
nand U13038 (N_13038,N_12600,N_12807);
nor U13039 (N_13039,N_12977,N_12978);
xor U13040 (N_13040,N_12818,N_12975);
and U13041 (N_13041,N_12854,N_12824);
nand U13042 (N_13042,N_12984,N_12762);
nor U13043 (N_13043,N_12931,N_12914);
and U13044 (N_13044,N_12850,N_12721);
and U13045 (N_13045,N_12973,N_12903);
nor U13046 (N_13046,N_12822,N_12682);
and U13047 (N_13047,N_12897,N_12735);
or U13048 (N_13048,N_12741,N_12925);
or U13049 (N_13049,N_12507,N_12661);
nor U13050 (N_13050,N_12890,N_12604);
xor U13051 (N_13051,N_12543,N_12606);
and U13052 (N_13052,N_12969,N_12621);
nor U13053 (N_13053,N_12865,N_12993);
nand U13054 (N_13054,N_12652,N_12511);
nor U13055 (N_13055,N_12583,N_12938);
or U13056 (N_13056,N_12677,N_12779);
or U13057 (N_13057,N_12763,N_12520);
or U13058 (N_13058,N_12631,N_12965);
nor U13059 (N_13059,N_12569,N_12803);
nand U13060 (N_13060,N_12957,N_12705);
and U13061 (N_13061,N_12713,N_12605);
and U13062 (N_13062,N_12668,N_12537);
or U13063 (N_13063,N_12676,N_12608);
nor U13064 (N_13064,N_12703,N_12559);
and U13065 (N_13065,N_12572,N_12727);
nand U13066 (N_13066,N_12571,N_12638);
nor U13067 (N_13067,N_12774,N_12835);
nand U13068 (N_13068,N_12519,N_12787);
xor U13069 (N_13069,N_12666,N_12637);
nor U13070 (N_13070,N_12589,N_12830);
and U13071 (N_13071,N_12684,N_12568);
and U13072 (N_13072,N_12949,N_12551);
nand U13073 (N_13073,N_12650,N_12670);
and U13074 (N_13074,N_12619,N_12972);
xnor U13075 (N_13075,N_12767,N_12745);
xnor U13076 (N_13076,N_12706,N_12930);
nor U13077 (N_13077,N_12581,N_12592);
and U13078 (N_13078,N_12504,N_12796);
nand U13079 (N_13079,N_12742,N_12748);
and U13080 (N_13080,N_12833,N_12772);
nor U13081 (N_13081,N_12565,N_12927);
or U13082 (N_13082,N_12823,N_12910);
and U13083 (N_13083,N_12771,N_12955);
or U13084 (N_13084,N_12776,N_12634);
nor U13085 (N_13085,N_12514,N_12734);
or U13086 (N_13086,N_12855,N_12853);
nor U13087 (N_13087,N_12699,N_12883);
and U13088 (N_13088,N_12523,N_12531);
nand U13089 (N_13089,N_12789,N_12868);
and U13090 (N_13090,N_12548,N_12674);
nor U13091 (N_13091,N_12819,N_12554);
or U13092 (N_13092,N_12765,N_12935);
and U13093 (N_13093,N_12909,N_12804);
nand U13094 (N_13094,N_12746,N_12760);
or U13095 (N_13095,N_12597,N_12550);
or U13096 (N_13096,N_12873,N_12696);
xor U13097 (N_13097,N_12743,N_12898);
nand U13098 (N_13098,N_12584,N_12797);
xor U13099 (N_13099,N_12724,N_12539);
or U13100 (N_13100,N_12546,N_12820);
or U13101 (N_13101,N_12882,N_12846);
and U13102 (N_13102,N_12593,N_12937);
nor U13103 (N_13103,N_12747,N_12545);
nand U13104 (N_13104,N_12726,N_12980);
and U13105 (N_13105,N_12996,N_12946);
nor U13106 (N_13106,N_12516,N_12595);
xor U13107 (N_13107,N_12733,N_12971);
nor U13108 (N_13108,N_12780,N_12576);
nor U13109 (N_13109,N_12751,N_12889);
nor U13110 (N_13110,N_12544,N_12547);
and U13111 (N_13111,N_12959,N_12785);
or U13112 (N_13112,N_12717,N_12950);
and U13113 (N_13113,N_12912,N_12867);
or U13114 (N_13114,N_12687,N_12794);
and U13115 (N_13115,N_12500,N_12922);
nor U13116 (N_13116,N_12613,N_12893);
xor U13117 (N_13117,N_12648,N_12626);
nand U13118 (N_13118,N_12885,N_12679);
nor U13119 (N_13119,N_12947,N_12782);
or U13120 (N_13120,N_12928,N_12612);
and U13121 (N_13121,N_12536,N_12693);
or U13122 (N_13122,N_12533,N_12786);
xnor U13123 (N_13123,N_12616,N_12770);
nor U13124 (N_13124,N_12738,N_12646);
xor U13125 (N_13125,N_12956,N_12702);
and U13126 (N_13126,N_12623,N_12525);
nand U13127 (N_13127,N_12960,N_12840);
nand U13128 (N_13128,N_12532,N_12872);
xnor U13129 (N_13129,N_12591,N_12647);
nand U13130 (N_13130,N_12755,N_12849);
xnor U13131 (N_13131,N_12821,N_12778);
or U13132 (N_13132,N_12508,N_12952);
xnor U13133 (N_13133,N_12802,N_12916);
nand U13134 (N_13134,N_12715,N_12618);
or U13135 (N_13135,N_12768,N_12769);
nand U13136 (N_13136,N_12654,N_12538);
nor U13137 (N_13137,N_12526,N_12869);
and U13138 (N_13138,N_12761,N_12683);
nor U13139 (N_13139,N_12837,N_12556);
nor U13140 (N_13140,N_12845,N_12673);
nand U13141 (N_13141,N_12660,N_12940);
nand U13142 (N_13142,N_12590,N_12982);
nand U13143 (N_13143,N_12575,N_12948);
or U13144 (N_13144,N_12753,N_12783);
xor U13145 (N_13145,N_12598,N_12578);
or U13146 (N_13146,N_12586,N_12798);
nand U13147 (N_13147,N_12918,N_12719);
nand U13148 (N_13148,N_12881,N_12603);
nand U13149 (N_13149,N_12838,N_12790);
or U13150 (N_13150,N_12983,N_12594);
nand U13151 (N_13151,N_12880,N_12685);
nor U13152 (N_13152,N_12981,N_12828);
nor U13153 (N_13153,N_12800,N_12506);
nand U13154 (N_13154,N_12601,N_12732);
nor U13155 (N_13155,N_12588,N_12878);
nand U13156 (N_13156,N_12939,N_12622);
and U13157 (N_13157,N_12635,N_12990);
or U13158 (N_13158,N_12624,N_12989);
and U13159 (N_13159,N_12919,N_12582);
nand U13160 (N_13160,N_12585,N_12691);
and U13161 (N_13161,N_12555,N_12809);
and U13162 (N_13162,N_12805,N_12766);
nor U13163 (N_13163,N_12908,N_12788);
and U13164 (N_13164,N_12627,N_12549);
or U13165 (N_13165,N_12784,N_12810);
nor U13166 (N_13166,N_12570,N_12967);
nand U13167 (N_13167,N_12958,N_12801);
nand U13168 (N_13168,N_12792,N_12904);
and U13169 (N_13169,N_12617,N_12954);
xor U13170 (N_13170,N_12929,N_12566);
xnor U13171 (N_13171,N_12528,N_12987);
nand U13172 (N_13172,N_12887,N_12832);
and U13173 (N_13173,N_12645,N_12710);
and U13174 (N_13174,N_12577,N_12563);
xnor U13175 (N_13175,N_12659,N_12558);
and U13176 (N_13176,N_12907,N_12799);
nor U13177 (N_13177,N_12737,N_12512);
and U13178 (N_13178,N_12813,N_12875);
nor U13179 (N_13179,N_12899,N_12857);
nand U13180 (N_13180,N_12863,N_12817);
or U13181 (N_13181,N_12895,N_12870);
nor U13182 (N_13182,N_12864,N_12709);
nor U13183 (N_13183,N_12791,N_12663);
nor U13184 (N_13184,N_12720,N_12503);
nand U13185 (N_13185,N_12806,N_12808);
nor U13186 (N_13186,N_12991,N_12961);
and U13187 (N_13187,N_12628,N_12518);
or U13188 (N_13188,N_12886,N_12974);
or U13189 (N_13189,N_12629,N_12723);
nand U13190 (N_13190,N_12858,N_12859);
or U13191 (N_13191,N_12686,N_12681);
xnor U13192 (N_13192,N_12970,N_12884);
nand U13193 (N_13193,N_12945,N_12611);
nand U13194 (N_13194,N_12560,N_12708);
or U13195 (N_13195,N_12649,N_12968);
or U13196 (N_13196,N_12879,N_12831);
and U13197 (N_13197,N_12573,N_12689);
nor U13198 (N_13198,N_12933,N_12557);
nor U13199 (N_13199,N_12680,N_12662);
nand U13200 (N_13200,N_12911,N_12501);
nand U13201 (N_13201,N_12657,N_12614);
nor U13202 (N_13202,N_12540,N_12942);
or U13203 (N_13203,N_12752,N_12754);
or U13204 (N_13204,N_12976,N_12827);
or U13205 (N_13205,N_12744,N_12561);
xor U13206 (N_13206,N_12736,N_12836);
or U13207 (N_13207,N_12943,N_12894);
nor U13208 (N_13208,N_12630,N_12992);
and U13209 (N_13209,N_12841,N_12905);
and U13210 (N_13210,N_12609,N_12521);
nand U13211 (N_13211,N_12900,N_12936);
xor U13212 (N_13212,N_12694,N_12750);
nand U13213 (N_13213,N_12795,N_12749);
nand U13214 (N_13214,N_12667,N_12932);
nor U13215 (N_13215,N_12923,N_12530);
or U13216 (N_13216,N_12842,N_12552);
and U13217 (N_13217,N_12941,N_12892);
nor U13218 (N_13218,N_12862,N_12698);
and U13219 (N_13219,N_12620,N_12651);
or U13220 (N_13220,N_12640,N_12759);
and U13221 (N_13221,N_12844,N_12851);
or U13222 (N_13222,N_12542,N_12625);
or U13223 (N_13223,N_12599,N_12728);
nor U13224 (N_13224,N_12775,N_12615);
nand U13225 (N_13225,N_12688,N_12722);
and U13226 (N_13226,N_12716,N_12515);
nand U13227 (N_13227,N_12944,N_12580);
nor U13228 (N_13228,N_12866,N_12527);
nand U13229 (N_13229,N_12860,N_12690);
nand U13230 (N_13230,N_12522,N_12773);
nor U13231 (N_13231,N_12636,N_12934);
nor U13232 (N_13232,N_12697,N_12509);
and U13233 (N_13233,N_12998,N_12655);
nand U13234 (N_13234,N_12695,N_12731);
nor U13235 (N_13235,N_12816,N_12644);
or U13236 (N_13236,N_12852,N_12924);
nor U13237 (N_13237,N_12596,N_12718);
and U13238 (N_13238,N_12541,N_12913);
and U13239 (N_13239,N_12729,N_12757);
or U13240 (N_13240,N_12921,N_12953);
nor U13241 (N_13241,N_12896,N_12675);
or U13242 (N_13242,N_12730,N_12906);
nor U13243 (N_13243,N_12502,N_12665);
nand U13244 (N_13244,N_12995,N_12553);
nand U13245 (N_13245,N_12920,N_12658);
or U13246 (N_13246,N_12607,N_12848);
xor U13247 (N_13247,N_12839,N_12826);
or U13248 (N_13248,N_12966,N_12535);
and U13249 (N_13249,N_12843,N_12758);
nand U13250 (N_13250,N_12955,N_12936);
nand U13251 (N_13251,N_12635,N_12610);
nor U13252 (N_13252,N_12922,N_12763);
nor U13253 (N_13253,N_12811,N_12833);
nand U13254 (N_13254,N_12976,N_12670);
or U13255 (N_13255,N_12703,N_12947);
xnor U13256 (N_13256,N_12768,N_12555);
xor U13257 (N_13257,N_12923,N_12675);
nor U13258 (N_13258,N_12962,N_12664);
nand U13259 (N_13259,N_12599,N_12534);
and U13260 (N_13260,N_12505,N_12703);
nand U13261 (N_13261,N_12700,N_12860);
xor U13262 (N_13262,N_12623,N_12808);
and U13263 (N_13263,N_12579,N_12827);
and U13264 (N_13264,N_12670,N_12566);
nor U13265 (N_13265,N_12507,N_12824);
or U13266 (N_13266,N_12934,N_12616);
xor U13267 (N_13267,N_12561,N_12873);
xor U13268 (N_13268,N_12848,N_12729);
and U13269 (N_13269,N_12809,N_12697);
and U13270 (N_13270,N_12927,N_12699);
or U13271 (N_13271,N_12668,N_12768);
nand U13272 (N_13272,N_12671,N_12990);
nand U13273 (N_13273,N_12685,N_12936);
nand U13274 (N_13274,N_12629,N_12526);
nor U13275 (N_13275,N_12766,N_12683);
nor U13276 (N_13276,N_12532,N_12546);
or U13277 (N_13277,N_12552,N_12874);
and U13278 (N_13278,N_12790,N_12900);
and U13279 (N_13279,N_12850,N_12650);
nor U13280 (N_13280,N_12929,N_12973);
and U13281 (N_13281,N_12919,N_12767);
or U13282 (N_13282,N_12878,N_12829);
nor U13283 (N_13283,N_12853,N_12819);
xor U13284 (N_13284,N_12624,N_12709);
nand U13285 (N_13285,N_12663,N_12826);
nor U13286 (N_13286,N_12944,N_12954);
nand U13287 (N_13287,N_12826,N_12977);
xor U13288 (N_13288,N_12988,N_12820);
or U13289 (N_13289,N_12985,N_12768);
and U13290 (N_13290,N_12845,N_12816);
nand U13291 (N_13291,N_12634,N_12862);
or U13292 (N_13292,N_12587,N_12717);
and U13293 (N_13293,N_12671,N_12779);
xnor U13294 (N_13294,N_12990,N_12743);
nor U13295 (N_13295,N_12783,N_12687);
nand U13296 (N_13296,N_12752,N_12653);
xor U13297 (N_13297,N_12710,N_12985);
nand U13298 (N_13298,N_12558,N_12832);
or U13299 (N_13299,N_12763,N_12811);
xor U13300 (N_13300,N_12891,N_12644);
or U13301 (N_13301,N_12672,N_12602);
xnor U13302 (N_13302,N_12782,N_12575);
and U13303 (N_13303,N_12723,N_12856);
or U13304 (N_13304,N_12705,N_12501);
and U13305 (N_13305,N_12646,N_12938);
xnor U13306 (N_13306,N_12902,N_12774);
and U13307 (N_13307,N_12860,N_12554);
xor U13308 (N_13308,N_12898,N_12607);
and U13309 (N_13309,N_12692,N_12606);
nor U13310 (N_13310,N_12889,N_12697);
nand U13311 (N_13311,N_12837,N_12503);
nand U13312 (N_13312,N_12529,N_12632);
or U13313 (N_13313,N_12908,N_12697);
or U13314 (N_13314,N_12684,N_12846);
nand U13315 (N_13315,N_12906,N_12568);
nand U13316 (N_13316,N_12922,N_12697);
and U13317 (N_13317,N_12920,N_12817);
or U13318 (N_13318,N_12507,N_12852);
nor U13319 (N_13319,N_12646,N_12873);
xnor U13320 (N_13320,N_12680,N_12763);
nor U13321 (N_13321,N_12631,N_12863);
and U13322 (N_13322,N_12590,N_12964);
nor U13323 (N_13323,N_12999,N_12636);
and U13324 (N_13324,N_12818,N_12592);
nor U13325 (N_13325,N_12682,N_12692);
and U13326 (N_13326,N_12564,N_12793);
and U13327 (N_13327,N_12655,N_12772);
nand U13328 (N_13328,N_12809,N_12892);
and U13329 (N_13329,N_12567,N_12766);
nand U13330 (N_13330,N_12861,N_12580);
nand U13331 (N_13331,N_12897,N_12957);
nand U13332 (N_13332,N_12746,N_12822);
or U13333 (N_13333,N_12991,N_12990);
nor U13334 (N_13334,N_12889,N_12789);
nand U13335 (N_13335,N_12782,N_12953);
nor U13336 (N_13336,N_12892,N_12672);
nor U13337 (N_13337,N_12956,N_12816);
nand U13338 (N_13338,N_12804,N_12674);
nand U13339 (N_13339,N_12911,N_12979);
and U13340 (N_13340,N_12605,N_12824);
and U13341 (N_13341,N_12844,N_12625);
or U13342 (N_13342,N_12893,N_12790);
nor U13343 (N_13343,N_12663,N_12944);
and U13344 (N_13344,N_12877,N_12581);
or U13345 (N_13345,N_12787,N_12719);
or U13346 (N_13346,N_12788,N_12533);
and U13347 (N_13347,N_12660,N_12918);
nand U13348 (N_13348,N_12510,N_12757);
nand U13349 (N_13349,N_12625,N_12919);
and U13350 (N_13350,N_12958,N_12749);
nor U13351 (N_13351,N_12696,N_12795);
or U13352 (N_13352,N_12678,N_12824);
xor U13353 (N_13353,N_12620,N_12554);
or U13354 (N_13354,N_12507,N_12767);
nor U13355 (N_13355,N_12878,N_12508);
nor U13356 (N_13356,N_12623,N_12731);
xnor U13357 (N_13357,N_12837,N_12976);
or U13358 (N_13358,N_12675,N_12701);
nor U13359 (N_13359,N_12562,N_12683);
nand U13360 (N_13360,N_12758,N_12809);
nand U13361 (N_13361,N_12798,N_12516);
nor U13362 (N_13362,N_12704,N_12808);
and U13363 (N_13363,N_12912,N_12646);
or U13364 (N_13364,N_12839,N_12838);
and U13365 (N_13365,N_12527,N_12707);
nand U13366 (N_13366,N_12643,N_12874);
and U13367 (N_13367,N_12779,N_12754);
nand U13368 (N_13368,N_12765,N_12620);
or U13369 (N_13369,N_12914,N_12532);
nand U13370 (N_13370,N_12570,N_12693);
and U13371 (N_13371,N_12685,N_12595);
nor U13372 (N_13372,N_12583,N_12785);
and U13373 (N_13373,N_12942,N_12734);
or U13374 (N_13374,N_12605,N_12998);
and U13375 (N_13375,N_12852,N_12931);
or U13376 (N_13376,N_12920,N_12644);
nor U13377 (N_13377,N_12975,N_12746);
and U13378 (N_13378,N_12756,N_12689);
nand U13379 (N_13379,N_12794,N_12796);
nand U13380 (N_13380,N_12613,N_12817);
and U13381 (N_13381,N_12786,N_12600);
or U13382 (N_13382,N_12992,N_12510);
nor U13383 (N_13383,N_12542,N_12768);
nand U13384 (N_13384,N_12604,N_12835);
nand U13385 (N_13385,N_12743,N_12728);
nand U13386 (N_13386,N_12969,N_12609);
nor U13387 (N_13387,N_12940,N_12765);
or U13388 (N_13388,N_12758,N_12750);
or U13389 (N_13389,N_12756,N_12781);
or U13390 (N_13390,N_12567,N_12939);
and U13391 (N_13391,N_12606,N_12999);
xnor U13392 (N_13392,N_12884,N_12920);
and U13393 (N_13393,N_12774,N_12900);
or U13394 (N_13394,N_12870,N_12936);
and U13395 (N_13395,N_12622,N_12722);
nand U13396 (N_13396,N_12682,N_12622);
and U13397 (N_13397,N_12876,N_12722);
or U13398 (N_13398,N_12721,N_12650);
nand U13399 (N_13399,N_12899,N_12695);
nor U13400 (N_13400,N_12504,N_12635);
and U13401 (N_13401,N_12532,N_12583);
nand U13402 (N_13402,N_12804,N_12660);
or U13403 (N_13403,N_12799,N_12716);
or U13404 (N_13404,N_12816,N_12597);
and U13405 (N_13405,N_12891,N_12518);
nand U13406 (N_13406,N_12704,N_12572);
or U13407 (N_13407,N_12684,N_12782);
or U13408 (N_13408,N_12886,N_12612);
or U13409 (N_13409,N_12694,N_12895);
or U13410 (N_13410,N_12718,N_12906);
xor U13411 (N_13411,N_12591,N_12951);
nor U13412 (N_13412,N_12697,N_12812);
nand U13413 (N_13413,N_12878,N_12912);
xor U13414 (N_13414,N_12954,N_12763);
or U13415 (N_13415,N_12881,N_12955);
nor U13416 (N_13416,N_12612,N_12644);
nor U13417 (N_13417,N_12704,N_12853);
or U13418 (N_13418,N_12973,N_12540);
and U13419 (N_13419,N_12505,N_12849);
or U13420 (N_13420,N_12513,N_12738);
nand U13421 (N_13421,N_12541,N_12955);
or U13422 (N_13422,N_12903,N_12582);
nor U13423 (N_13423,N_12865,N_12775);
xor U13424 (N_13424,N_12604,N_12599);
nor U13425 (N_13425,N_12776,N_12924);
nor U13426 (N_13426,N_12683,N_12519);
or U13427 (N_13427,N_12862,N_12607);
or U13428 (N_13428,N_12635,N_12621);
xor U13429 (N_13429,N_12926,N_12878);
xnor U13430 (N_13430,N_12924,N_12823);
nor U13431 (N_13431,N_12896,N_12748);
and U13432 (N_13432,N_12590,N_12825);
xnor U13433 (N_13433,N_12526,N_12964);
xnor U13434 (N_13434,N_12537,N_12638);
nand U13435 (N_13435,N_12791,N_12936);
or U13436 (N_13436,N_12631,N_12557);
nor U13437 (N_13437,N_12928,N_12513);
or U13438 (N_13438,N_12594,N_12949);
and U13439 (N_13439,N_12848,N_12684);
nor U13440 (N_13440,N_12884,N_12681);
nor U13441 (N_13441,N_12868,N_12921);
nor U13442 (N_13442,N_12613,N_12767);
nand U13443 (N_13443,N_12601,N_12964);
or U13444 (N_13444,N_12994,N_12884);
nor U13445 (N_13445,N_12694,N_12519);
xor U13446 (N_13446,N_12656,N_12574);
xnor U13447 (N_13447,N_12793,N_12812);
or U13448 (N_13448,N_12665,N_12896);
xor U13449 (N_13449,N_12654,N_12928);
or U13450 (N_13450,N_12695,N_12638);
nand U13451 (N_13451,N_12581,N_12513);
or U13452 (N_13452,N_12633,N_12883);
nand U13453 (N_13453,N_12994,N_12688);
nand U13454 (N_13454,N_12706,N_12657);
nor U13455 (N_13455,N_12883,N_12630);
nor U13456 (N_13456,N_12804,N_12646);
nand U13457 (N_13457,N_12872,N_12906);
nor U13458 (N_13458,N_12567,N_12604);
nor U13459 (N_13459,N_12871,N_12540);
or U13460 (N_13460,N_12816,N_12777);
nand U13461 (N_13461,N_12650,N_12814);
nor U13462 (N_13462,N_12503,N_12751);
and U13463 (N_13463,N_12866,N_12894);
xnor U13464 (N_13464,N_12747,N_12707);
and U13465 (N_13465,N_12699,N_12881);
nor U13466 (N_13466,N_12624,N_12610);
or U13467 (N_13467,N_12879,N_12603);
and U13468 (N_13468,N_12625,N_12680);
nand U13469 (N_13469,N_12587,N_12803);
or U13470 (N_13470,N_12591,N_12763);
and U13471 (N_13471,N_12838,N_12597);
nor U13472 (N_13472,N_12527,N_12812);
and U13473 (N_13473,N_12754,N_12682);
nand U13474 (N_13474,N_12962,N_12637);
xor U13475 (N_13475,N_12628,N_12830);
nand U13476 (N_13476,N_12902,N_12561);
or U13477 (N_13477,N_12626,N_12619);
or U13478 (N_13478,N_12678,N_12681);
and U13479 (N_13479,N_12616,N_12881);
or U13480 (N_13480,N_12762,N_12939);
nand U13481 (N_13481,N_12956,N_12540);
nand U13482 (N_13482,N_12507,N_12982);
xor U13483 (N_13483,N_12532,N_12707);
nand U13484 (N_13484,N_12768,N_12750);
or U13485 (N_13485,N_12674,N_12599);
and U13486 (N_13486,N_12989,N_12611);
or U13487 (N_13487,N_12892,N_12845);
nand U13488 (N_13488,N_12841,N_12891);
and U13489 (N_13489,N_12975,N_12847);
nand U13490 (N_13490,N_12927,N_12749);
xor U13491 (N_13491,N_12889,N_12900);
and U13492 (N_13492,N_12743,N_12708);
or U13493 (N_13493,N_12826,N_12925);
xnor U13494 (N_13494,N_12598,N_12775);
and U13495 (N_13495,N_12553,N_12915);
nor U13496 (N_13496,N_12626,N_12705);
nor U13497 (N_13497,N_12654,N_12708);
nand U13498 (N_13498,N_12750,N_12583);
nand U13499 (N_13499,N_12596,N_12661);
or U13500 (N_13500,N_13424,N_13419);
xor U13501 (N_13501,N_13026,N_13092);
nor U13502 (N_13502,N_13139,N_13364);
or U13503 (N_13503,N_13193,N_13072);
nor U13504 (N_13504,N_13440,N_13163);
nor U13505 (N_13505,N_13299,N_13421);
nor U13506 (N_13506,N_13089,N_13337);
nor U13507 (N_13507,N_13006,N_13395);
nor U13508 (N_13508,N_13159,N_13296);
nor U13509 (N_13509,N_13396,N_13399);
xor U13510 (N_13510,N_13214,N_13063);
and U13511 (N_13511,N_13207,N_13404);
or U13512 (N_13512,N_13410,N_13316);
nand U13513 (N_13513,N_13047,N_13438);
and U13514 (N_13514,N_13434,N_13075);
nor U13515 (N_13515,N_13258,N_13447);
nand U13516 (N_13516,N_13161,N_13441);
and U13517 (N_13517,N_13373,N_13336);
nand U13518 (N_13518,N_13050,N_13425);
or U13519 (N_13519,N_13433,N_13151);
nand U13520 (N_13520,N_13194,N_13169);
xnor U13521 (N_13521,N_13403,N_13414);
and U13522 (N_13522,N_13426,N_13381);
nor U13523 (N_13523,N_13230,N_13120);
or U13524 (N_13524,N_13067,N_13146);
xnor U13525 (N_13525,N_13321,N_13331);
or U13526 (N_13526,N_13107,N_13234);
nor U13527 (N_13527,N_13235,N_13097);
nand U13528 (N_13528,N_13477,N_13312);
xnor U13529 (N_13529,N_13480,N_13061);
nor U13530 (N_13530,N_13085,N_13117);
or U13531 (N_13531,N_13040,N_13225);
or U13532 (N_13532,N_13209,N_13211);
and U13533 (N_13533,N_13466,N_13429);
nand U13534 (N_13534,N_13221,N_13378);
or U13535 (N_13535,N_13273,N_13347);
or U13536 (N_13536,N_13228,N_13383);
or U13537 (N_13537,N_13152,N_13180);
and U13538 (N_13538,N_13079,N_13463);
nand U13539 (N_13539,N_13417,N_13288);
and U13540 (N_13540,N_13282,N_13494);
nand U13541 (N_13541,N_13239,N_13366);
or U13542 (N_13542,N_13392,N_13223);
and U13543 (N_13543,N_13432,N_13017);
nand U13544 (N_13544,N_13041,N_13135);
nand U13545 (N_13545,N_13363,N_13175);
nand U13546 (N_13546,N_13240,N_13226);
or U13547 (N_13547,N_13264,N_13053);
and U13548 (N_13548,N_13390,N_13314);
and U13549 (N_13549,N_13475,N_13087);
nor U13550 (N_13550,N_13397,N_13100);
xnor U13551 (N_13551,N_13317,N_13367);
and U13552 (N_13552,N_13188,N_13197);
nand U13553 (N_13553,N_13166,N_13110);
and U13554 (N_13554,N_13242,N_13405);
or U13555 (N_13555,N_13138,N_13099);
and U13556 (N_13556,N_13245,N_13150);
xor U13557 (N_13557,N_13157,N_13398);
xor U13558 (N_13558,N_13490,N_13122);
or U13559 (N_13559,N_13354,N_13095);
or U13560 (N_13560,N_13012,N_13307);
or U13561 (N_13561,N_13269,N_13034);
and U13562 (N_13562,N_13134,N_13431);
nand U13563 (N_13563,N_13492,N_13292);
or U13564 (N_13564,N_13465,N_13476);
nand U13565 (N_13565,N_13105,N_13220);
nor U13566 (N_13566,N_13196,N_13218);
or U13567 (N_13567,N_13439,N_13001);
nor U13568 (N_13568,N_13481,N_13145);
or U13569 (N_13569,N_13275,N_13411);
or U13570 (N_13570,N_13114,N_13037);
or U13571 (N_13571,N_13164,N_13078);
nor U13572 (N_13572,N_13015,N_13201);
xnor U13573 (N_13573,N_13177,N_13022);
or U13574 (N_13574,N_13020,N_13402);
and U13575 (N_13575,N_13204,N_13305);
or U13576 (N_13576,N_13147,N_13160);
and U13577 (N_13577,N_13136,N_13210);
and U13578 (N_13578,N_13200,N_13168);
or U13579 (N_13579,N_13348,N_13303);
nor U13580 (N_13580,N_13217,N_13249);
and U13581 (N_13581,N_13301,N_13064);
and U13582 (N_13582,N_13025,N_13371);
and U13583 (N_13583,N_13448,N_13167);
nor U13584 (N_13584,N_13370,N_13171);
and U13585 (N_13585,N_13250,N_13243);
nor U13586 (N_13586,N_13437,N_13073);
or U13587 (N_13587,N_13199,N_13495);
nand U13588 (N_13588,N_13387,N_13393);
or U13589 (N_13589,N_13076,N_13415);
nor U13590 (N_13590,N_13124,N_13340);
xnor U13591 (N_13591,N_13339,N_13335);
nor U13592 (N_13592,N_13016,N_13238);
and U13593 (N_13593,N_13290,N_13352);
nand U13594 (N_13594,N_13256,N_13057);
and U13595 (N_13595,N_13195,N_13450);
nor U13596 (N_13596,N_13007,N_13108);
and U13597 (N_13597,N_13345,N_13187);
or U13598 (N_13598,N_13189,N_13322);
nand U13599 (N_13599,N_13498,N_13010);
and U13600 (N_13600,N_13126,N_13133);
xnor U13601 (N_13601,N_13319,N_13236);
or U13602 (N_13602,N_13030,N_13130);
or U13603 (N_13603,N_13191,N_13036);
and U13604 (N_13604,N_13140,N_13461);
nand U13605 (N_13605,N_13077,N_13048);
nand U13606 (N_13606,N_13186,N_13311);
nor U13607 (N_13607,N_13384,N_13469);
or U13608 (N_13608,N_13179,N_13208);
nand U13609 (N_13609,N_13298,N_13070);
or U13610 (N_13610,N_13115,N_13054);
and U13611 (N_13611,N_13284,N_13062);
or U13612 (N_13612,N_13056,N_13278);
and U13613 (N_13613,N_13257,N_13005);
or U13614 (N_13614,N_13202,N_13153);
nand U13615 (N_13615,N_13148,N_13141);
and U13616 (N_13616,N_13129,N_13368);
xor U13617 (N_13617,N_13142,N_13013);
and U13618 (N_13618,N_13086,N_13111);
nand U13619 (N_13619,N_13467,N_13259);
nand U13620 (N_13620,N_13182,N_13262);
nand U13621 (N_13621,N_13444,N_13229);
or U13622 (N_13622,N_13241,N_13499);
nand U13623 (N_13623,N_13365,N_13325);
nand U13624 (N_13624,N_13281,N_13031);
nand U13625 (N_13625,N_13004,N_13183);
nand U13626 (N_13626,N_13318,N_13081);
or U13627 (N_13627,N_13266,N_13118);
or U13628 (N_13628,N_13400,N_13473);
and U13629 (N_13629,N_13423,N_13224);
and U13630 (N_13630,N_13216,N_13178);
and U13631 (N_13631,N_13009,N_13024);
nand U13632 (N_13632,N_13329,N_13125);
and U13633 (N_13633,N_13458,N_13029);
nand U13634 (N_13634,N_13049,N_13449);
xor U13635 (N_13635,N_13362,N_13309);
or U13636 (N_13636,N_13190,N_13462);
and U13637 (N_13637,N_13315,N_13091);
nand U13638 (N_13638,N_13289,N_13442);
nand U13639 (N_13639,N_13332,N_13185);
nor U13640 (N_13640,N_13341,N_13389);
nand U13641 (N_13641,N_13286,N_13069);
nand U13642 (N_13642,N_13413,N_13355);
and U13643 (N_13643,N_13394,N_13094);
or U13644 (N_13644,N_13386,N_13422);
or U13645 (N_13645,N_13102,N_13268);
nor U13646 (N_13646,N_13103,N_13478);
nor U13647 (N_13647,N_13101,N_13119);
and U13648 (N_13648,N_13082,N_13128);
or U13649 (N_13649,N_13039,N_13359);
nor U13650 (N_13650,N_13409,N_13008);
or U13651 (N_13651,N_13274,N_13104);
or U13652 (N_13652,N_13295,N_13059);
nor U13653 (N_13653,N_13088,N_13372);
xnor U13654 (N_13654,N_13412,N_13098);
nand U13655 (N_13655,N_13058,N_13472);
nor U13656 (N_13656,N_13260,N_13346);
or U13657 (N_13657,N_13497,N_13351);
and U13658 (N_13658,N_13283,N_13356);
nand U13659 (N_13659,N_13377,N_13358);
nor U13660 (N_13660,N_13028,N_13483);
nor U13661 (N_13661,N_13255,N_13454);
nor U13662 (N_13662,N_13109,N_13192);
and U13663 (N_13663,N_13326,N_13485);
nand U13664 (N_13664,N_13375,N_13173);
and U13665 (N_13665,N_13452,N_13215);
or U13666 (N_13666,N_13418,N_13172);
and U13667 (N_13667,N_13043,N_13493);
nand U13668 (N_13668,N_13174,N_13338);
or U13669 (N_13669,N_13093,N_13297);
or U13670 (N_13670,N_13032,N_13457);
or U13671 (N_13671,N_13276,N_13330);
nor U13672 (N_13672,N_13132,N_13045);
and U13673 (N_13673,N_13446,N_13113);
nor U13674 (N_13674,N_13486,N_13310);
or U13675 (N_13675,N_13206,N_13051);
nand U13676 (N_13676,N_13002,N_13158);
xnor U13677 (N_13677,N_13248,N_13237);
or U13678 (N_13678,N_13127,N_13451);
or U13679 (N_13679,N_13324,N_13406);
and U13680 (N_13680,N_13019,N_13123);
and U13681 (N_13681,N_13474,N_13154);
and U13682 (N_13682,N_13165,N_13033);
xnor U13683 (N_13683,N_13149,N_13388);
nor U13684 (N_13684,N_13408,N_13470);
or U13685 (N_13685,N_13181,N_13334);
xor U13686 (N_13686,N_13044,N_13277);
nand U13687 (N_13687,N_13323,N_13071);
and U13688 (N_13688,N_13251,N_13106);
nand U13689 (N_13689,N_13488,N_13000);
or U13690 (N_13690,N_13144,N_13263);
or U13691 (N_13691,N_13420,N_13084);
or U13692 (N_13692,N_13369,N_13407);
xnor U13693 (N_13693,N_13162,N_13270);
or U13694 (N_13694,N_13170,N_13300);
nor U13695 (N_13695,N_13304,N_13291);
and U13696 (N_13696,N_13279,N_13382);
or U13697 (N_13697,N_13333,N_13261);
nor U13698 (N_13698,N_13205,N_13460);
or U13699 (N_13699,N_13353,N_13385);
xnor U13700 (N_13700,N_13343,N_13083);
xor U13701 (N_13701,N_13023,N_13021);
or U13702 (N_13702,N_13436,N_13246);
or U13703 (N_13703,N_13137,N_13443);
nand U13704 (N_13704,N_13287,N_13052);
nor U13705 (N_13705,N_13468,N_13328);
nand U13706 (N_13706,N_13342,N_13184);
and U13707 (N_13707,N_13380,N_13046);
and U13708 (N_13708,N_13313,N_13066);
or U13709 (N_13709,N_13293,N_13265);
nor U13710 (N_13710,N_13121,N_13445);
nand U13711 (N_13711,N_13320,N_13038);
and U13712 (N_13712,N_13042,N_13489);
and U13713 (N_13713,N_13272,N_13011);
xnor U13714 (N_13714,N_13491,N_13456);
nor U13715 (N_13715,N_13280,N_13080);
nand U13716 (N_13716,N_13244,N_13227);
and U13717 (N_13717,N_13427,N_13294);
xor U13718 (N_13718,N_13203,N_13267);
or U13719 (N_13719,N_13096,N_13176);
or U13720 (N_13720,N_13360,N_13027);
or U13721 (N_13721,N_13379,N_13285);
nand U13722 (N_13722,N_13247,N_13401);
nor U13723 (N_13723,N_13484,N_13455);
or U13724 (N_13724,N_13232,N_13350);
or U13725 (N_13725,N_13035,N_13482);
and U13726 (N_13726,N_13302,N_13156);
and U13727 (N_13727,N_13376,N_13349);
nor U13728 (N_13728,N_13464,N_13306);
and U13729 (N_13729,N_13254,N_13252);
nor U13730 (N_13730,N_13131,N_13361);
nand U13731 (N_13731,N_13222,N_13219);
nor U13732 (N_13732,N_13213,N_13090);
and U13733 (N_13733,N_13430,N_13471);
or U13734 (N_13734,N_13487,N_13479);
or U13735 (N_13735,N_13391,N_13198);
or U13736 (N_13736,N_13074,N_13496);
nand U13737 (N_13737,N_13233,N_13416);
and U13738 (N_13738,N_13428,N_13374);
or U13739 (N_13739,N_13116,N_13143);
nand U13740 (N_13740,N_13231,N_13018);
and U13741 (N_13741,N_13344,N_13060);
and U13742 (N_13742,N_13357,N_13453);
nand U13743 (N_13743,N_13212,N_13327);
or U13744 (N_13744,N_13068,N_13065);
and U13745 (N_13745,N_13112,N_13308);
nand U13746 (N_13746,N_13459,N_13014);
or U13747 (N_13747,N_13055,N_13271);
nand U13748 (N_13748,N_13155,N_13253);
nor U13749 (N_13749,N_13435,N_13003);
nor U13750 (N_13750,N_13008,N_13436);
or U13751 (N_13751,N_13299,N_13221);
and U13752 (N_13752,N_13376,N_13039);
nor U13753 (N_13753,N_13334,N_13192);
or U13754 (N_13754,N_13262,N_13092);
nor U13755 (N_13755,N_13225,N_13471);
nand U13756 (N_13756,N_13189,N_13195);
nor U13757 (N_13757,N_13150,N_13047);
nor U13758 (N_13758,N_13238,N_13307);
or U13759 (N_13759,N_13328,N_13279);
nor U13760 (N_13760,N_13419,N_13008);
and U13761 (N_13761,N_13388,N_13014);
or U13762 (N_13762,N_13257,N_13343);
nor U13763 (N_13763,N_13445,N_13401);
nand U13764 (N_13764,N_13009,N_13040);
or U13765 (N_13765,N_13201,N_13412);
and U13766 (N_13766,N_13414,N_13265);
nor U13767 (N_13767,N_13212,N_13162);
nor U13768 (N_13768,N_13313,N_13483);
nand U13769 (N_13769,N_13186,N_13488);
xnor U13770 (N_13770,N_13032,N_13048);
nand U13771 (N_13771,N_13291,N_13341);
nor U13772 (N_13772,N_13346,N_13485);
nand U13773 (N_13773,N_13394,N_13363);
nor U13774 (N_13774,N_13436,N_13350);
nor U13775 (N_13775,N_13479,N_13064);
nand U13776 (N_13776,N_13225,N_13272);
and U13777 (N_13777,N_13139,N_13240);
nor U13778 (N_13778,N_13408,N_13458);
nand U13779 (N_13779,N_13473,N_13172);
xnor U13780 (N_13780,N_13132,N_13456);
and U13781 (N_13781,N_13196,N_13391);
and U13782 (N_13782,N_13429,N_13432);
or U13783 (N_13783,N_13408,N_13067);
nor U13784 (N_13784,N_13157,N_13041);
and U13785 (N_13785,N_13455,N_13237);
nor U13786 (N_13786,N_13248,N_13465);
nand U13787 (N_13787,N_13208,N_13438);
nor U13788 (N_13788,N_13339,N_13316);
nand U13789 (N_13789,N_13476,N_13399);
and U13790 (N_13790,N_13046,N_13487);
or U13791 (N_13791,N_13380,N_13170);
nand U13792 (N_13792,N_13222,N_13278);
nand U13793 (N_13793,N_13032,N_13361);
or U13794 (N_13794,N_13410,N_13472);
nand U13795 (N_13795,N_13487,N_13427);
and U13796 (N_13796,N_13145,N_13128);
or U13797 (N_13797,N_13276,N_13296);
nor U13798 (N_13798,N_13243,N_13180);
nand U13799 (N_13799,N_13315,N_13467);
nand U13800 (N_13800,N_13291,N_13479);
nand U13801 (N_13801,N_13449,N_13405);
nor U13802 (N_13802,N_13302,N_13418);
and U13803 (N_13803,N_13118,N_13202);
nand U13804 (N_13804,N_13438,N_13009);
or U13805 (N_13805,N_13123,N_13282);
nand U13806 (N_13806,N_13054,N_13283);
and U13807 (N_13807,N_13195,N_13073);
nor U13808 (N_13808,N_13334,N_13362);
and U13809 (N_13809,N_13261,N_13254);
nor U13810 (N_13810,N_13488,N_13440);
and U13811 (N_13811,N_13394,N_13199);
and U13812 (N_13812,N_13429,N_13032);
nor U13813 (N_13813,N_13435,N_13015);
nor U13814 (N_13814,N_13205,N_13428);
and U13815 (N_13815,N_13499,N_13322);
nor U13816 (N_13816,N_13142,N_13282);
nand U13817 (N_13817,N_13300,N_13064);
nand U13818 (N_13818,N_13409,N_13176);
nor U13819 (N_13819,N_13073,N_13484);
xor U13820 (N_13820,N_13067,N_13096);
and U13821 (N_13821,N_13477,N_13222);
nor U13822 (N_13822,N_13006,N_13075);
and U13823 (N_13823,N_13343,N_13452);
nand U13824 (N_13824,N_13310,N_13452);
nand U13825 (N_13825,N_13276,N_13143);
nor U13826 (N_13826,N_13048,N_13122);
or U13827 (N_13827,N_13098,N_13313);
nor U13828 (N_13828,N_13149,N_13407);
nand U13829 (N_13829,N_13339,N_13402);
and U13830 (N_13830,N_13191,N_13337);
nand U13831 (N_13831,N_13144,N_13009);
or U13832 (N_13832,N_13038,N_13247);
and U13833 (N_13833,N_13465,N_13490);
nand U13834 (N_13834,N_13457,N_13413);
nor U13835 (N_13835,N_13362,N_13163);
or U13836 (N_13836,N_13483,N_13367);
and U13837 (N_13837,N_13212,N_13474);
or U13838 (N_13838,N_13284,N_13430);
and U13839 (N_13839,N_13141,N_13409);
and U13840 (N_13840,N_13267,N_13245);
and U13841 (N_13841,N_13426,N_13275);
nand U13842 (N_13842,N_13492,N_13091);
xnor U13843 (N_13843,N_13247,N_13053);
or U13844 (N_13844,N_13329,N_13481);
or U13845 (N_13845,N_13236,N_13311);
nor U13846 (N_13846,N_13145,N_13491);
nor U13847 (N_13847,N_13369,N_13256);
nor U13848 (N_13848,N_13403,N_13001);
or U13849 (N_13849,N_13105,N_13050);
nand U13850 (N_13850,N_13154,N_13043);
and U13851 (N_13851,N_13474,N_13201);
xor U13852 (N_13852,N_13101,N_13473);
and U13853 (N_13853,N_13443,N_13083);
or U13854 (N_13854,N_13398,N_13322);
and U13855 (N_13855,N_13175,N_13093);
or U13856 (N_13856,N_13110,N_13041);
nor U13857 (N_13857,N_13366,N_13026);
and U13858 (N_13858,N_13421,N_13011);
or U13859 (N_13859,N_13478,N_13425);
nor U13860 (N_13860,N_13309,N_13037);
and U13861 (N_13861,N_13449,N_13493);
nand U13862 (N_13862,N_13409,N_13082);
nand U13863 (N_13863,N_13486,N_13408);
nand U13864 (N_13864,N_13249,N_13318);
nand U13865 (N_13865,N_13432,N_13453);
nand U13866 (N_13866,N_13190,N_13004);
xnor U13867 (N_13867,N_13472,N_13073);
or U13868 (N_13868,N_13476,N_13374);
and U13869 (N_13869,N_13104,N_13088);
nand U13870 (N_13870,N_13400,N_13102);
or U13871 (N_13871,N_13185,N_13087);
nand U13872 (N_13872,N_13447,N_13353);
nor U13873 (N_13873,N_13028,N_13098);
nor U13874 (N_13874,N_13048,N_13124);
or U13875 (N_13875,N_13164,N_13009);
and U13876 (N_13876,N_13266,N_13049);
nor U13877 (N_13877,N_13297,N_13164);
nor U13878 (N_13878,N_13087,N_13269);
and U13879 (N_13879,N_13163,N_13371);
and U13880 (N_13880,N_13188,N_13177);
nand U13881 (N_13881,N_13435,N_13403);
and U13882 (N_13882,N_13122,N_13100);
nor U13883 (N_13883,N_13031,N_13211);
and U13884 (N_13884,N_13076,N_13106);
xnor U13885 (N_13885,N_13359,N_13042);
and U13886 (N_13886,N_13454,N_13420);
xnor U13887 (N_13887,N_13474,N_13014);
nor U13888 (N_13888,N_13431,N_13243);
or U13889 (N_13889,N_13081,N_13246);
or U13890 (N_13890,N_13451,N_13073);
nand U13891 (N_13891,N_13121,N_13010);
or U13892 (N_13892,N_13383,N_13016);
and U13893 (N_13893,N_13182,N_13230);
nand U13894 (N_13894,N_13365,N_13371);
and U13895 (N_13895,N_13328,N_13079);
nand U13896 (N_13896,N_13401,N_13082);
nand U13897 (N_13897,N_13318,N_13403);
nand U13898 (N_13898,N_13404,N_13136);
nor U13899 (N_13899,N_13422,N_13244);
or U13900 (N_13900,N_13306,N_13355);
nor U13901 (N_13901,N_13086,N_13203);
and U13902 (N_13902,N_13135,N_13029);
nand U13903 (N_13903,N_13045,N_13237);
or U13904 (N_13904,N_13331,N_13305);
nand U13905 (N_13905,N_13197,N_13196);
or U13906 (N_13906,N_13207,N_13170);
xor U13907 (N_13907,N_13379,N_13220);
or U13908 (N_13908,N_13173,N_13320);
nor U13909 (N_13909,N_13133,N_13385);
or U13910 (N_13910,N_13199,N_13433);
and U13911 (N_13911,N_13024,N_13012);
nand U13912 (N_13912,N_13486,N_13249);
xor U13913 (N_13913,N_13185,N_13444);
nand U13914 (N_13914,N_13403,N_13205);
nand U13915 (N_13915,N_13420,N_13356);
nor U13916 (N_13916,N_13028,N_13153);
and U13917 (N_13917,N_13095,N_13496);
and U13918 (N_13918,N_13056,N_13285);
nand U13919 (N_13919,N_13065,N_13323);
xnor U13920 (N_13920,N_13485,N_13070);
nand U13921 (N_13921,N_13366,N_13331);
or U13922 (N_13922,N_13342,N_13252);
xor U13923 (N_13923,N_13266,N_13317);
nor U13924 (N_13924,N_13119,N_13472);
nor U13925 (N_13925,N_13027,N_13044);
and U13926 (N_13926,N_13231,N_13241);
and U13927 (N_13927,N_13375,N_13191);
or U13928 (N_13928,N_13406,N_13058);
nor U13929 (N_13929,N_13225,N_13159);
or U13930 (N_13930,N_13314,N_13182);
nor U13931 (N_13931,N_13381,N_13374);
or U13932 (N_13932,N_13163,N_13445);
xor U13933 (N_13933,N_13212,N_13381);
nand U13934 (N_13934,N_13158,N_13096);
nand U13935 (N_13935,N_13040,N_13073);
nand U13936 (N_13936,N_13084,N_13321);
nor U13937 (N_13937,N_13302,N_13056);
and U13938 (N_13938,N_13121,N_13036);
nor U13939 (N_13939,N_13228,N_13195);
or U13940 (N_13940,N_13338,N_13157);
nor U13941 (N_13941,N_13407,N_13123);
nand U13942 (N_13942,N_13109,N_13017);
xnor U13943 (N_13943,N_13175,N_13085);
xnor U13944 (N_13944,N_13258,N_13001);
and U13945 (N_13945,N_13129,N_13273);
and U13946 (N_13946,N_13057,N_13285);
and U13947 (N_13947,N_13239,N_13014);
or U13948 (N_13948,N_13175,N_13310);
nor U13949 (N_13949,N_13288,N_13249);
or U13950 (N_13950,N_13440,N_13127);
nor U13951 (N_13951,N_13463,N_13041);
or U13952 (N_13952,N_13057,N_13085);
or U13953 (N_13953,N_13059,N_13456);
nor U13954 (N_13954,N_13376,N_13233);
nand U13955 (N_13955,N_13183,N_13153);
and U13956 (N_13956,N_13297,N_13211);
nand U13957 (N_13957,N_13011,N_13414);
nand U13958 (N_13958,N_13150,N_13248);
nand U13959 (N_13959,N_13422,N_13060);
or U13960 (N_13960,N_13115,N_13155);
nor U13961 (N_13961,N_13474,N_13258);
nand U13962 (N_13962,N_13432,N_13444);
nand U13963 (N_13963,N_13198,N_13356);
nand U13964 (N_13964,N_13423,N_13398);
nor U13965 (N_13965,N_13112,N_13096);
and U13966 (N_13966,N_13109,N_13460);
or U13967 (N_13967,N_13355,N_13094);
and U13968 (N_13968,N_13297,N_13014);
nand U13969 (N_13969,N_13437,N_13153);
and U13970 (N_13970,N_13282,N_13154);
or U13971 (N_13971,N_13389,N_13375);
and U13972 (N_13972,N_13086,N_13282);
nor U13973 (N_13973,N_13433,N_13003);
and U13974 (N_13974,N_13467,N_13416);
xnor U13975 (N_13975,N_13047,N_13350);
or U13976 (N_13976,N_13007,N_13119);
nor U13977 (N_13977,N_13073,N_13248);
or U13978 (N_13978,N_13006,N_13127);
or U13979 (N_13979,N_13294,N_13279);
nand U13980 (N_13980,N_13068,N_13483);
nand U13981 (N_13981,N_13076,N_13097);
nand U13982 (N_13982,N_13333,N_13218);
nor U13983 (N_13983,N_13196,N_13247);
nor U13984 (N_13984,N_13158,N_13373);
and U13985 (N_13985,N_13078,N_13327);
or U13986 (N_13986,N_13026,N_13419);
and U13987 (N_13987,N_13264,N_13100);
nand U13988 (N_13988,N_13370,N_13367);
and U13989 (N_13989,N_13408,N_13054);
or U13990 (N_13990,N_13055,N_13151);
and U13991 (N_13991,N_13233,N_13333);
nand U13992 (N_13992,N_13055,N_13012);
nor U13993 (N_13993,N_13338,N_13042);
or U13994 (N_13994,N_13311,N_13105);
nor U13995 (N_13995,N_13005,N_13109);
nor U13996 (N_13996,N_13147,N_13417);
or U13997 (N_13997,N_13019,N_13112);
nand U13998 (N_13998,N_13003,N_13037);
and U13999 (N_13999,N_13200,N_13029);
and U14000 (N_14000,N_13569,N_13702);
nand U14001 (N_14001,N_13983,N_13874);
nor U14002 (N_14002,N_13704,N_13508);
and U14003 (N_14003,N_13553,N_13577);
and U14004 (N_14004,N_13899,N_13651);
nand U14005 (N_14005,N_13628,N_13610);
nand U14006 (N_14006,N_13908,N_13964);
or U14007 (N_14007,N_13841,N_13836);
xor U14008 (N_14008,N_13799,N_13753);
or U14009 (N_14009,N_13611,N_13898);
and U14010 (N_14010,N_13919,N_13878);
and U14011 (N_14011,N_13959,N_13670);
or U14012 (N_14012,N_13803,N_13656);
and U14013 (N_14013,N_13594,N_13905);
xnor U14014 (N_14014,N_13922,N_13510);
xnor U14015 (N_14015,N_13870,N_13539);
or U14016 (N_14016,N_13987,N_13957);
nand U14017 (N_14017,N_13906,N_13563);
nand U14018 (N_14018,N_13981,N_13666);
or U14019 (N_14019,N_13505,N_13746);
nand U14020 (N_14020,N_13572,N_13731);
or U14021 (N_14021,N_13686,N_13969);
nor U14022 (N_14022,N_13629,N_13661);
and U14023 (N_14023,N_13543,N_13848);
nand U14024 (N_14024,N_13769,N_13793);
xnor U14025 (N_14025,N_13607,N_13559);
nand U14026 (N_14026,N_13917,N_13837);
nor U14027 (N_14027,N_13744,N_13839);
and U14028 (N_14028,N_13672,N_13788);
nor U14029 (N_14029,N_13824,N_13787);
nand U14030 (N_14030,N_13972,N_13859);
nor U14031 (N_14031,N_13524,N_13897);
or U14032 (N_14032,N_13657,N_13915);
or U14033 (N_14033,N_13928,N_13778);
nand U14034 (N_14034,N_13631,N_13749);
and U14035 (N_14035,N_13502,N_13528);
and U14036 (N_14036,N_13944,N_13718);
nor U14037 (N_14037,N_13534,N_13893);
nand U14038 (N_14038,N_13679,N_13891);
or U14039 (N_14039,N_13568,N_13785);
xnor U14040 (N_14040,N_13624,N_13844);
xnor U14041 (N_14041,N_13766,N_13587);
nor U14042 (N_14042,N_13832,N_13912);
xor U14043 (N_14043,N_13556,N_13835);
nand U14044 (N_14044,N_13762,N_13834);
nor U14045 (N_14045,N_13984,N_13650);
nor U14046 (N_14046,N_13620,N_13740);
and U14047 (N_14047,N_13907,N_13940);
or U14048 (N_14048,N_13947,N_13723);
nor U14049 (N_14049,N_13576,N_13971);
nor U14050 (N_14050,N_13786,N_13732);
nand U14051 (N_14051,N_13939,N_13635);
nor U14052 (N_14052,N_13851,N_13843);
and U14053 (N_14053,N_13822,N_13700);
nand U14054 (N_14054,N_13688,N_13768);
nor U14055 (N_14055,N_13641,N_13767);
or U14056 (N_14056,N_13671,N_13750);
and U14057 (N_14057,N_13630,N_13782);
nor U14058 (N_14058,N_13717,N_13809);
or U14059 (N_14059,N_13578,N_13684);
and U14060 (N_14060,N_13888,N_13941);
nand U14061 (N_14061,N_13527,N_13862);
nand U14062 (N_14062,N_13789,N_13952);
nand U14063 (N_14063,N_13673,N_13660);
or U14064 (N_14064,N_13734,N_13930);
or U14065 (N_14065,N_13826,N_13975);
xnor U14066 (N_14066,N_13820,N_13810);
nand U14067 (N_14067,N_13927,N_13948);
nand U14068 (N_14068,N_13840,N_13754);
and U14069 (N_14069,N_13821,N_13573);
or U14070 (N_14070,N_13501,N_13982);
nand U14071 (N_14071,N_13701,N_13872);
or U14072 (N_14072,N_13612,N_13916);
xor U14073 (N_14073,N_13616,N_13604);
nor U14074 (N_14074,N_13733,N_13986);
xor U14075 (N_14075,N_13513,N_13558);
nand U14076 (N_14076,N_13581,N_13721);
xor U14077 (N_14077,N_13711,N_13649);
nor U14078 (N_14078,N_13950,N_13823);
nand U14079 (N_14079,N_13866,N_13997);
nor U14080 (N_14080,N_13910,N_13755);
nor U14081 (N_14081,N_13695,N_13980);
nand U14082 (N_14082,N_13989,N_13637);
and U14083 (N_14083,N_13640,N_13942);
and U14084 (N_14084,N_13595,N_13546);
xnor U14085 (N_14085,N_13998,N_13802);
and U14086 (N_14086,N_13691,N_13662);
xnor U14087 (N_14087,N_13901,N_13579);
nor U14088 (N_14088,N_13590,N_13690);
and U14089 (N_14089,N_13970,N_13920);
or U14090 (N_14090,N_13934,N_13596);
or U14091 (N_14091,N_13867,N_13693);
nand U14092 (N_14092,N_13668,N_13896);
xor U14093 (N_14093,N_13991,N_13511);
and U14094 (N_14094,N_13523,N_13623);
nand U14095 (N_14095,N_13938,N_13589);
and U14096 (N_14096,N_13993,N_13864);
nor U14097 (N_14097,N_13812,N_13949);
and U14098 (N_14098,N_13555,N_13730);
xnor U14099 (N_14099,N_13564,N_13936);
nor U14100 (N_14100,N_13902,N_13815);
nor U14101 (N_14101,N_13724,N_13760);
and U14102 (N_14102,N_13976,N_13707);
and U14103 (N_14103,N_13520,N_13894);
or U14104 (N_14104,N_13714,N_13542);
nor U14105 (N_14105,N_13638,N_13725);
nor U14106 (N_14106,N_13680,N_13654);
or U14107 (N_14107,N_13531,N_13847);
or U14108 (N_14108,N_13973,N_13665);
or U14109 (N_14109,N_13602,N_13667);
and U14110 (N_14110,N_13798,N_13842);
nand U14111 (N_14111,N_13593,N_13538);
and U14112 (N_14112,N_13882,N_13537);
nand U14113 (N_14113,N_13540,N_13655);
and U14114 (N_14114,N_13575,N_13692);
nand U14115 (N_14115,N_13549,N_13791);
and U14116 (N_14116,N_13833,N_13828);
nand U14117 (N_14117,N_13554,N_13876);
nand U14118 (N_14118,N_13658,N_13911);
or U14119 (N_14119,N_13644,N_13547);
nor U14120 (N_14120,N_13979,N_13988);
or U14121 (N_14121,N_13796,N_13779);
and U14122 (N_14122,N_13503,N_13951);
nand U14123 (N_14123,N_13921,N_13647);
nor U14124 (N_14124,N_13801,N_13817);
nand U14125 (N_14125,N_13929,N_13738);
nor U14126 (N_14126,N_13758,N_13884);
nand U14127 (N_14127,N_13999,N_13943);
nand U14128 (N_14128,N_13933,N_13525);
nor U14129 (N_14129,N_13591,N_13885);
or U14130 (N_14130,N_13518,N_13830);
nor U14131 (N_14131,N_13562,N_13974);
and U14132 (N_14132,N_13869,N_13530);
nand U14133 (N_14133,N_13825,N_13605);
xnor U14134 (N_14134,N_13565,N_13966);
and U14135 (N_14135,N_13727,N_13560);
nor U14136 (N_14136,N_13653,N_13715);
or U14137 (N_14137,N_13852,N_13804);
xor U14138 (N_14138,N_13506,N_13963);
nand U14139 (N_14139,N_13736,N_13516);
or U14140 (N_14140,N_13918,N_13705);
nand U14141 (N_14141,N_13773,N_13507);
nor U14142 (N_14142,N_13992,N_13892);
and U14143 (N_14143,N_13622,N_13625);
and U14144 (N_14144,N_13515,N_13926);
nand U14145 (N_14145,N_13858,N_13535);
or U14146 (N_14146,N_13584,N_13722);
or U14147 (N_14147,N_13741,N_13829);
and U14148 (N_14148,N_13855,N_13931);
or U14149 (N_14149,N_13532,N_13699);
and U14150 (N_14150,N_13886,N_13875);
or U14151 (N_14151,N_13677,N_13761);
nor U14152 (N_14152,N_13609,N_13621);
and U14153 (N_14153,N_13696,N_13648);
nand U14154 (N_14154,N_13945,N_13519);
and U14155 (N_14155,N_13923,N_13813);
and U14156 (N_14156,N_13978,N_13757);
nand U14157 (N_14157,N_13617,N_13889);
nand U14158 (N_14158,N_13639,N_13792);
and U14159 (N_14159,N_13827,N_13606);
nand U14160 (N_14160,N_13710,N_13694);
and U14161 (N_14161,N_13608,N_13808);
xnor U14162 (N_14162,N_13962,N_13509);
nor U14163 (N_14163,N_13853,N_13561);
nor U14164 (N_14164,N_13600,N_13689);
nor U14165 (N_14165,N_13687,N_13881);
and U14166 (N_14166,N_13582,N_13551);
or U14167 (N_14167,N_13883,N_13770);
nand U14168 (N_14168,N_13784,N_13681);
or U14169 (N_14169,N_13856,N_13706);
and U14170 (N_14170,N_13735,N_13720);
nand U14171 (N_14171,N_13529,N_13737);
and U14172 (N_14172,N_13583,N_13849);
nand U14173 (N_14173,N_13709,N_13863);
and U14174 (N_14174,N_13990,N_13965);
and U14175 (N_14175,N_13995,N_13548);
nand U14176 (N_14176,N_13713,N_13676);
nor U14177 (N_14177,N_13500,N_13586);
nand U14178 (N_14178,N_13504,N_13946);
and U14179 (N_14179,N_13937,N_13879);
or U14180 (N_14180,N_13729,N_13873);
nor U14181 (N_14181,N_13626,N_13985);
or U14182 (N_14182,N_13861,N_13967);
nand U14183 (N_14183,N_13712,N_13742);
nand U14184 (N_14184,N_13765,N_13790);
or U14185 (N_14185,N_13541,N_13663);
nor U14186 (N_14186,N_13592,N_13580);
xor U14187 (N_14187,N_13685,N_13968);
and U14188 (N_14188,N_13599,N_13845);
nand U14189 (N_14189,N_13683,N_13996);
or U14190 (N_14190,N_13536,N_13764);
or U14191 (N_14191,N_13924,N_13675);
or U14192 (N_14192,N_13961,N_13806);
and U14193 (N_14193,N_13614,N_13585);
or U14194 (N_14194,N_13756,N_13652);
and U14195 (N_14195,N_13954,N_13747);
nand U14196 (N_14196,N_13953,N_13634);
nor U14197 (N_14197,N_13752,N_13903);
nor U14198 (N_14198,N_13545,N_13636);
and U14199 (N_14199,N_13763,N_13805);
nand U14200 (N_14200,N_13566,N_13567);
and U14201 (N_14201,N_13783,N_13748);
nand U14202 (N_14202,N_13645,N_13800);
or U14203 (N_14203,N_13719,N_13743);
and U14204 (N_14204,N_13517,N_13552);
or U14205 (N_14205,N_13574,N_13774);
or U14206 (N_14206,N_13659,N_13708);
and U14207 (N_14207,N_13698,N_13643);
and U14208 (N_14208,N_13550,N_13913);
or U14209 (N_14209,N_13814,N_13646);
or U14210 (N_14210,N_13588,N_13781);
and U14211 (N_14211,N_13914,N_13925);
nand U14212 (N_14212,N_13818,N_13977);
nor U14213 (N_14213,N_13775,N_13571);
and U14214 (N_14214,N_13890,N_13514);
or U14215 (N_14215,N_13598,N_13745);
or U14216 (N_14216,N_13871,N_13838);
or U14217 (N_14217,N_13726,N_13728);
or U14218 (N_14218,N_13960,N_13797);
and U14219 (N_14219,N_13904,N_13759);
nor U14220 (N_14220,N_13627,N_13682);
and U14221 (N_14221,N_13850,N_13860);
and U14222 (N_14222,N_13831,N_13512);
or U14223 (N_14223,N_13865,N_13909);
nor U14224 (N_14224,N_13615,N_13674);
or U14225 (N_14225,N_13618,N_13526);
or U14226 (N_14226,N_13664,N_13772);
or U14227 (N_14227,N_13544,N_13854);
nor U14228 (N_14228,N_13868,N_13807);
or U14229 (N_14229,N_13522,N_13771);
or U14230 (N_14230,N_13994,N_13603);
xnor U14231 (N_14231,N_13958,N_13857);
or U14232 (N_14232,N_13900,N_13816);
nand U14233 (N_14233,N_13819,N_13570);
and U14234 (N_14234,N_13703,N_13895);
nor U14235 (N_14235,N_13751,N_13956);
or U14236 (N_14236,N_13697,N_13880);
nor U14237 (N_14237,N_13533,N_13669);
and U14238 (N_14238,N_13619,N_13776);
nor U14239 (N_14239,N_13613,N_13633);
or U14240 (N_14240,N_13795,N_13739);
nand U14241 (N_14241,N_13777,N_13521);
nor U14242 (N_14242,N_13642,N_13601);
xor U14243 (N_14243,N_13811,N_13632);
and U14244 (N_14244,N_13877,N_13932);
and U14245 (N_14245,N_13887,N_13935);
or U14246 (N_14246,N_13794,N_13557);
nand U14247 (N_14247,N_13716,N_13780);
nor U14248 (N_14248,N_13597,N_13955);
nor U14249 (N_14249,N_13678,N_13846);
or U14250 (N_14250,N_13696,N_13710);
and U14251 (N_14251,N_13844,N_13548);
or U14252 (N_14252,N_13525,N_13716);
or U14253 (N_14253,N_13902,N_13586);
xnor U14254 (N_14254,N_13767,N_13728);
and U14255 (N_14255,N_13736,N_13535);
and U14256 (N_14256,N_13943,N_13503);
nand U14257 (N_14257,N_13910,N_13741);
or U14258 (N_14258,N_13630,N_13763);
nand U14259 (N_14259,N_13869,N_13579);
nor U14260 (N_14260,N_13844,N_13874);
or U14261 (N_14261,N_13512,N_13698);
nand U14262 (N_14262,N_13870,N_13622);
or U14263 (N_14263,N_13851,N_13759);
and U14264 (N_14264,N_13995,N_13814);
nor U14265 (N_14265,N_13833,N_13903);
and U14266 (N_14266,N_13837,N_13625);
nand U14267 (N_14267,N_13855,N_13563);
nand U14268 (N_14268,N_13842,N_13847);
or U14269 (N_14269,N_13535,N_13546);
nand U14270 (N_14270,N_13802,N_13514);
or U14271 (N_14271,N_13514,N_13836);
and U14272 (N_14272,N_13973,N_13917);
xnor U14273 (N_14273,N_13668,N_13899);
or U14274 (N_14274,N_13553,N_13995);
and U14275 (N_14275,N_13619,N_13872);
and U14276 (N_14276,N_13981,N_13964);
and U14277 (N_14277,N_13521,N_13755);
xnor U14278 (N_14278,N_13960,N_13627);
and U14279 (N_14279,N_13640,N_13661);
nor U14280 (N_14280,N_13580,N_13746);
or U14281 (N_14281,N_13732,N_13607);
or U14282 (N_14282,N_13894,N_13586);
or U14283 (N_14283,N_13515,N_13848);
xnor U14284 (N_14284,N_13890,N_13723);
xor U14285 (N_14285,N_13530,N_13913);
and U14286 (N_14286,N_13883,N_13673);
and U14287 (N_14287,N_13696,N_13677);
and U14288 (N_14288,N_13717,N_13860);
nand U14289 (N_14289,N_13507,N_13525);
xnor U14290 (N_14290,N_13559,N_13556);
nand U14291 (N_14291,N_13808,N_13525);
xor U14292 (N_14292,N_13816,N_13684);
xnor U14293 (N_14293,N_13586,N_13899);
nor U14294 (N_14294,N_13727,N_13849);
nor U14295 (N_14295,N_13549,N_13588);
nand U14296 (N_14296,N_13743,N_13519);
and U14297 (N_14297,N_13976,N_13690);
xor U14298 (N_14298,N_13840,N_13796);
or U14299 (N_14299,N_13706,N_13757);
nand U14300 (N_14300,N_13998,N_13529);
nand U14301 (N_14301,N_13689,N_13519);
or U14302 (N_14302,N_13772,N_13807);
and U14303 (N_14303,N_13535,N_13873);
and U14304 (N_14304,N_13993,N_13843);
and U14305 (N_14305,N_13794,N_13533);
nor U14306 (N_14306,N_13721,N_13906);
or U14307 (N_14307,N_13525,N_13880);
or U14308 (N_14308,N_13611,N_13708);
nor U14309 (N_14309,N_13617,N_13534);
nor U14310 (N_14310,N_13645,N_13935);
and U14311 (N_14311,N_13608,N_13918);
nor U14312 (N_14312,N_13759,N_13573);
nor U14313 (N_14313,N_13608,N_13749);
nor U14314 (N_14314,N_13718,N_13997);
nand U14315 (N_14315,N_13987,N_13572);
or U14316 (N_14316,N_13661,N_13556);
nand U14317 (N_14317,N_13534,N_13737);
and U14318 (N_14318,N_13938,N_13896);
nor U14319 (N_14319,N_13506,N_13646);
xor U14320 (N_14320,N_13654,N_13932);
nor U14321 (N_14321,N_13673,N_13965);
and U14322 (N_14322,N_13964,N_13930);
nand U14323 (N_14323,N_13536,N_13767);
nor U14324 (N_14324,N_13510,N_13687);
xor U14325 (N_14325,N_13708,N_13903);
and U14326 (N_14326,N_13868,N_13671);
nand U14327 (N_14327,N_13592,N_13958);
or U14328 (N_14328,N_13661,N_13718);
or U14329 (N_14329,N_13523,N_13755);
nand U14330 (N_14330,N_13663,N_13896);
xnor U14331 (N_14331,N_13592,N_13719);
nand U14332 (N_14332,N_13554,N_13985);
and U14333 (N_14333,N_13532,N_13569);
nor U14334 (N_14334,N_13790,N_13778);
nor U14335 (N_14335,N_13929,N_13613);
xnor U14336 (N_14336,N_13657,N_13621);
or U14337 (N_14337,N_13592,N_13775);
and U14338 (N_14338,N_13523,N_13541);
nand U14339 (N_14339,N_13920,N_13950);
nand U14340 (N_14340,N_13842,N_13737);
xor U14341 (N_14341,N_13738,N_13703);
nand U14342 (N_14342,N_13697,N_13598);
and U14343 (N_14343,N_13986,N_13947);
and U14344 (N_14344,N_13701,N_13759);
or U14345 (N_14345,N_13727,N_13974);
and U14346 (N_14346,N_13526,N_13646);
nand U14347 (N_14347,N_13695,N_13710);
nor U14348 (N_14348,N_13976,N_13845);
nor U14349 (N_14349,N_13539,N_13930);
nor U14350 (N_14350,N_13994,N_13722);
xnor U14351 (N_14351,N_13637,N_13826);
and U14352 (N_14352,N_13894,N_13661);
or U14353 (N_14353,N_13753,N_13617);
and U14354 (N_14354,N_13804,N_13621);
or U14355 (N_14355,N_13855,N_13847);
nor U14356 (N_14356,N_13956,N_13623);
nand U14357 (N_14357,N_13929,N_13563);
nand U14358 (N_14358,N_13845,N_13996);
or U14359 (N_14359,N_13681,N_13835);
and U14360 (N_14360,N_13750,N_13797);
xor U14361 (N_14361,N_13826,N_13688);
nand U14362 (N_14362,N_13776,N_13555);
nand U14363 (N_14363,N_13968,N_13993);
xnor U14364 (N_14364,N_13657,N_13820);
nor U14365 (N_14365,N_13618,N_13807);
nand U14366 (N_14366,N_13716,N_13619);
xnor U14367 (N_14367,N_13987,N_13595);
nand U14368 (N_14368,N_13589,N_13804);
and U14369 (N_14369,N_13957,N_13882);
nor U14370 (N_14370,N_13580,N_13801);
xnor U14371 (N_14371,N_13566,N_13695);
nor U14372 (N_14372,N_13892,N_13774);
nor U14373 (N_14373,N_13821,N_13764);
and U14374 (N_14374,N_13917,N_13931);
nor U14375 (N_14375,N_13601,N_13986);
nand U14376 (N_14376,N_13908,N_13600);
and U14377 (N_14377,N_13663,N_13632);
or U14378 (N_14378,N_13978,N_13949);
or U14379 (N_14379,N_13892,N_13825);
xor U14380 (N_14380,N_13683,N_13648);
nor U14381 (N_14381,N_13860,N_13809);
nand U14382 (N_14382,N_13884,N_13625);
and U14383 (N_14383,N_13837,N_13881);
nor U14384 (N_14384,N_13540,N_13939);
or U14385 (N_14385,N_13764,N_13592);
and U14386 (N_14386,N_13957,N_13748);
or U14387 (N_14387,N_13897,N_13849);
nand U14388 (N_14388,N_13817,N_13914);
or U14389 (N_14389,N_13895,N_13783);
or U14390 (N_14390,N_13943,N_13686);
nand U14391 (N_14391,N_13706,N_13839);
or U14392 (N_14392,N_13980,N_13908);
or U14393 (N_14393,N_13661,N_13665);
and U14394 (N_14394,N_13869,N_13503);
and U14395 (N_14395,N_13929,N_13916);
and U14396 (N_14396,N_13933,N_13592);
nor U14397 (N_14397,N_13542,N_13732);
and U14398 (N_14398,N_13587,N_13673);
or U14399 (N_14399,N_13649,N_13769);
xor U14400 (N_14400,N_13675,N_13522);
and U14401 (N_14401,N_13609,N_13982);
or U14402 (N_14402,N_13597,N_13573);
and U14403 (N_14403,N_13897,N_13925);
nand U14404 (N_14404,N_13572,N_13574);
nand U14405 (N_14405,N_13873,N_13719);
or U14406 (N_14406,N_13694,N_13548);
or U14407 (N_14407,N_13670,N_13895);
or U14408 (N_14408,N_13584,N_13817);
xnor U14409 (N_14409,N_13611,N_13533);
or U14410 (N_14410,N_13739,N_13755);
nand U14411 (N_14411,N_13795,N_13991);
and U14412 (N_14412,N_13900,N_13796);
or U14413 (N_14413,N_13834,N_13941);
or U14414 (N_14414,N_13707,N_13724);
nor U14415 (N_14415,N_13830,N_13800);
and U14416 (N_14416,N_13778,N_13508);
xnor U14417 (N_14417,N_13561,N_13696);
or U14418 (N_14418,N_13869,N_13696);
nand U14419 (N_14419,N_13664,N_13724);
nand U14420 (N_14420,N_13674,N_13909);
or U14421 (N_14421,N_13695,N_13574);
nor U14422 (N_14422,N_13911,N_13840);
nor U14423 (N_14423,N_13834,N_13686);
or U14424 (N_14424,N_13965,N_13715);
xor U14425 (N_14425,N_13893,N_13786);
or U14426 (N_14426,N_13690,N_13609);
nand U14427 (N_14427,N_13722,N_13801);
or U14428 (N_14428,N_13991,N_13860);
nor U14429 (N_14429,N_13778,N_13564);
and U14430 (N_14430,N_13721,N_13780);
or U14431 (N_14431,N_13832,N_13824);
or U14432 (N_14432,N_13998,N_13975);
nand U14433 (N_14433,N_13943,N_13743);
nor U14434 (N_14434,N_13702,N_13996);
or U14435 (N_14435,N_13958,N_13794);
nor U14436 (N_14436,N_13643,N_13854);
nand U14437 (N_14437,N_13646,N_13963);
xnor U14438 (N_14438,N_13681,N_13992);
nor U14439 (N_14439,N_13777,N_13800);
or U14440 (N_14440,N_13990,N_13815);
and U14441 (N_14441,N_13605,N_13814);
and U14442 (N_14442,N_13787,N_13747);
or U14443 (N_14443,N_13888,N_13959);
xor U14444 (N_14444,N_13731,N_13632);
or U14445 (N_14445,N_13552,N_13627);
nand U14446 (N_14446,N_13919,N_13786);
xnor U14447 (N_14447,N_13927,N_13844);
and U14448 (N_14448,N_13769,N_13694);
nand U14449 (N_14449,N_13888,N_13737);
or U14450 (N_14450,N_13988,N_13621);
and U14451 (N_14451,N_13977,N_13605);
or U14452 (N_14452,N_13857,N_13647);
nor U14453 (N_14453,N_13752,N_13753);
or U14454 (N_14454,N_13608,N_13525);
nor U14455 (N_14455,N_13602,N_13944);
nor U14456 (N_14456,N_13530,N_13722);
nor U14457 (N_14457,N_13617,N_13891);
nand U14458 (N_14458,N_13969,N_13649);
nand U14459 (N_14459,N_13646,N_13945);
nor U14460 (N_14460,N_13727,N_13862);
or U14461 (N_14461,N_13511,N_13690);
nor U14462 (N_14462,N_13627,N_13952);
and U14463 (N_14463,N_13573,N_13630);
nand U14464 (N_14464,N_13924,N_13587);
or U14465 (N_14465,N_13545,N_13549);
nand U14466 (N_14466,N_13709,N_13956);
and U14467 (N_14467,N_13676,N_13624);
nor U14468 (N_14468,N_13904,N_13963);
or U14469 (N_14469,N_13913,N_13681);
and U14470 (N_14470,N_13919,N_13805);
nand U14471 (N_14471,N_13843,N_13972);
nand U14472 (N_14472,N_13773,N_13577);
nand U14473 (N_14473,N_13565,N_13951);
or U14474 (N_14474,N_13939,N_13593);
and U14475 (N_14475,N_13826,N_13985);
nor U14476 (N_14476,N_13623,N_13684);
nor U14477 (N_14477,N_13546,N_13553);
and U14478 (N_14478,N_13541,N_13964);
or U14479 (N_14479,N_13842,N_13917);
or U14480 (N_14480,N_13887,N_13872);
or U14481 (N_14481,N_13674,N_13616);
nor U14482 (N_14482,N_13641,N_13721);
nor U14483 (N_14483,N_13688,N_13865);
nor U14484 (N_14484,N_13503,N_13532);
xor U14485 (N_14485,N_13904,N_13654);
xnor U14486 (N_14486,N_13940,N_13725);
nor U14487 (N_14487,N_13803,N_13855);
nor U14488 (N_14488,N_13856,N_13506);
or U14489 (N_14489,N_13583,N_13641);
and U14490 (N_14490,N_13513,N_13856);
nand U14491 (N_14491,N_13544,N_13508);
or U14492 (N_14492,N_13787,N_13989);
nand U14493 (N_14493,N_13948,N_13776);
and U14494 (N_14494,N_13662,N_13922);
nand U14495 (N_14495,N_13541,N_13669);
and U14496 (N_14496,N_13916,N_13634);
or U14497 (N_14497,N_13854,N_13949);
nor U14498 (N_14498,N_13999,N_13554);
nand U14499 (N_14499,N_13766,N_13568);
nand U14500 (N_14500,N_14248,N_14376);
xor U14501 (N_14501,N_14106,N_14401);
nand U14502 (N_14502,N_14490,N_14460);
xor U14503 (N_14503,N_14304,N_14125);
and U14504 (N_14504,N_14273,N_14305);
nand U14505 (N_14505,N_14452,N_14255);
nor U14506 (N_14506,N_14236,N_14225);
nand U14507 (N_14507,N_14339,N_14166);
nand U14508 (N_14508,N_14213,N_14066);
or U14509 (N_14509,N_14353,N_14456);
or U14510 (N_14510,N_14115,N_14061);
or U14511 (N_14511,N_14408,N_14204);
or U14512 (N_14512,N_14285,N_14244);
and U14513 (N_14513,N_14214,N_14040);
or U14514 (N_14514,N_14479,N_14447);
xnor U14515 (N_14515,N_14381,N_14357);
xor U14516 (N_14516,N_14471,N_14494);
and U14517 (N_14517,N_14393,N_14011);
nand U14518 (N_14518,N_14349,N_14152);
or U14519 (N_14519,N_14052,N_14022);
or U14520 (N_14520,N_14287,N_14361);
xnor U14521 (N_14521,N_14030,N_14084);
nand U14522 (N_14522,N_14492,N_14375);
xor U14523 (N_14523,N_14462,N_14228);
nor U14524 (N_14524,N_14094,N_14390);
nand U14525 (N_14525,N_14174,N_14006);
or U14526 (N_14526,N_14135,N_14158);
xor U14527 (N_14527,N_14189,N_14445);
and U14528 (N_14528,N_14055,N_14378);
or U14529 (N_14529,N_14137,N_14283);
or U14530 (N_14530,N_14433,N_14301);
or U14531 (N_14531,N_14466,N_14407);
xnor U14532 (N_14532,N_14120,N_14076);
or U14533 (N_14533,N_14418,N_14139);
and U14534 (N_14534,N_14156,N_14141);
and U14535 (N_14535,N_14288,N_14050);
nand U14536 (N_14536,N_14253,N_14063);
xor U14537 (N_14537,N_14464,N_14208);
nand U14538 (N_14538,N_14387,N_14033);
or U14539 (N_14539,N_14315,N_14146);
nand U14540 (N_14540,N_14048,N_14319);
nor U14541 (N_14541,N_14184,N_14270);
nor U14542 (N_14542,N_14252,N_14355);
or U14543 (N_14543,N_14123,N_14332);
nor U14544 (N_14544,N_14016,N_14099);
xnor U14545 (N_14545,N_14254,N_14493);
nand U14546 (N_14546,N_14019,N_14463);
or U14547 (N_14547,N_14303,N_14427);
xnor U14548 (N_14548,N_14042,N_14176);
or U14549 (N_14549,N_14110,N_14070);
nand U14550 (N_14550,N_14364,N_14198);
or U14551 (N_14551,N_14185,N_14018);
nor U14552 (N_14552,N_14369,N_14109);
nand U14553 (N_14553,N_14343,N_14468);
or U14554 (N_14554,N_14440,N_14275);
and U14555 (N_14555,N_14346,N_14154);
nor U14556 (N_14556,N_14437,N_14274);
or U14557 (N_14557,N_14177,N_14132);
and U14558 (N_14558,N_14151,N_14413);
or U14559 (N_14559,N_14075,N_14484);
nand U14560 (N_14560,N_14320,N_14021);
or U14561 (N_14561,N_14167,N_14017);
and U14562 (N_14562,N_14374,N_14327);
nand U14563 (N_14563,N_14264,N_14370);
xor U14564 (N_14564,N_14020,N_14444);
nand U14565 (N_14565,N_14197,N_14299);
or U14566 (N_14566,N_14009,N_14281);
and U14567 (N_14567,N_14068,N_14302);
nor U14568 (N_14568,N_14103,N_14180);
nor U14569 (N_14569,N_14086,N_14196);
or U14570 (N_14570,N_14163,N_14005);
and U14571 (N_14571,N_14219,N_14087);
and U14572 (N_14572,N_14350,N_14144);
nand U14573 (N_14573,N_14495,N_14414);
nor U14574 (N_14574,N_14307,N_14477);
xor U14575 (N_14575,N_14010,N_14382);
nand U14576 (N_14576,N_14227,N_14316);
and U14577 (N_14577,N_14206,N_14426);
and U14578 (N_14578,N_14238,N_14291);
nand U14579 (N_14579,N_14266,N_14015);
nand U14580 (N_14580,N_14483,N_14341);
nor U14581 (N_14581,N_14379,N_14239);
and U14582 (N_14582,N_14229,N_14113);
and U14583 (N_14583,N_14127,N_14140);
nor U14584 (N_14584,N_14187,N_14124);
nand U14585 (N_14585,N_14432,N_14191);
nand U14586 (N_14586,N_14164,N_14162);
nor U14587 (N_14587,N_14080,N_14342);
xnor U14588 (N_14588,N_14251,N_14182);
nand U14589 (N_14589,N_14212,N_14322);
nor U14590 (N_14590,N_14259,N_14446);
and U14591 (N_14591,N_14458,N_14027);
nand U14592 (N_14592,N_14358,N_14380);
nand U14593 (N_14593,N_14435,N_14143);
and U14594 (N_14594,N_14023,N_14114);
nand U14595 (N_14595,N_14280,N_14313);
nor U14596 (N_14596,N_14035,N_14395);
and U14597 (N_14597,N_14450,N_14488);
xor U14598 (N_14598,N_14107,N_14069);
nand U14599 (N_14599,N_14297,N_14039);
nor U14600 (N_14600,N_14203,N_14134);
or U14601 (N_14601,N_14088,N_14480);
or U14602 (N_14602,N_14294,N_14478);
nor U14603 (N_14603,N_14454,N_14383);
or U14604 (N_14604,N_14059,N_14279);
nor U14605 (N_14605,N_14205,N_14360);
xor U14606 (N_14606,N_14058,N_14108);
or U14607 (N_14607,N_14241,N_14249);
or U14608 (N_14608,N_14008,N_14377);
or U14609 (N_14609,N_14218,N_14474);
or U14610 (N_14610,N_14155,N_14062);
nand U14611 (N_14611,N_14153,N_14100);
nor U14612 (N_14612,N_14041,N_14138);
nor U14613 (N_14613,N_14260,N_14003);
nor U14614 (N_14614,N_14095,N_14311);
nor U14615 (N_14615,N_14425,N_14193);
or U14616 (N_14616,N_14060,N_14220);
or U14617 (N_14617,N_14194,N_14046);
or U14618 (N_14618,N_14476,N_14324);
nand U14619 (N_14619,N_14424,N_14118);
xor U14620 (N_14620,N_14000,N_14415);
nor U14621 (N_14621,N_14243,N_14293);
nor U14622 (N_14622,N_14234,N_14047);
and U14623 (N_14623,N_14178,N_14130);
xnor U14624 (N_14624,N_14429,N_14145);
or U14625 (N_14625,N_14306,N_14286);
nor U14626 (N_14626,N_14133,N_14049);
and U14627 (N_14627,N_14232,N_14221);
nand U14628 (N_14628,N_14072,N_14200);
and U14629 (N_14629,N_14053,N_14417);
nor U14630 (N_14630,N_14290,N_14356);
or U14631 (N_14631,N_14338,N_14334);
or U14632 (N_14632,N_14400,N_14029);
xnor U14633 (N_14633,N_14131,N_14065);
nor U14634 (N_14634,N_14263,N_14430);
nor U14635 (N_14635,N_14171,N_14037);
nor U14636 (N_14636,N_14237,N_14481);
nand U14637 (N_14637,N_14173,N_14186);
or U14638 (N_14638,N_14412,N_14295);
nand U14639 (N_14639,N_14201,N_14034);
or U14640 (N_14640,N_14001,N_14215);
nor U14641 (N_14641,N_14265,N_14347);
nor U14642 (N_14642,N_14129,N_14128);
nor U14643 (N_14643,N_14292,N_14312);
or U14644 (N_14644,N_14475,N_14309);
and U14645 (N_14645,N_14328,N_14121);
nor U14646 (N_14646,N_14199,N_14465);
and U14647 (N_14647,N_14392,N_14271);
or U14648 (N_14648,N_14261,N_14181);
nand U14649 (N_14649,N_14386,N_14160);
and U14650 (N_14650,N_14246,N_14406);
nor U14651 (N_14651,N_14366,N_14165);
nor U14652 (N_14652,N_14074,N_14496);
nand U14653 (N_14653,N_14233,N_14067);
nand U14654 (N_14654,N_14004,N_14344);
nor U14655 (N_14655,N_14242,N_14489);
and U14656 (N_14656,N_14148,N_14276);
nor U14657 (N_14657,N_14073,N_14278);
nor U14658 (N_14658,N_14256,N_14397);
or U14659 (N_14659,N_14404,N_14335);
and U14660 (N_14660,N_14116,N_14472);
nand U14661 (N_14661,N_14470,N_14428);
or U14662 (N_14662,N_14368,N_14031);
nor U14663 (N_14663,N_14365,N_14399);
nor U14664 (N_14664,N_14025,N_14410);
or U14665 (N_14665,N_14222,N_14269);
nor U14666 (N_14666,N_14459,N_14223);
and U14667 (N_14667,N_14321,N_14240);
nand U14668 (N_14668,N_14211,N_14331);
nand U14669 (N_14669,N_14102,N_14455);
and U14670 (N_14670,N_14056,N_14032);
nor U14671 (N_14671,N_14284,N_14230);
and U14672 (N_14672,N_14434,N_14351);
nor U14673 (N_14673,N_14363,N_14117);
nand U14674 (N_14674,N_14389,N_14258);
and U14675 (N_14675,N_14391,N_14416);
nand U14676 (N_14676,N_14439,N_14420);
nor U14677 (N_14677,N_14217,N_14482);
nor U14678 (N_14678,N_14498,N_14409);
nor U14679 (N_14679,N_14354,N_14448);
nand U14680 (N_14680,N_14345,N_14012);
nor U14681 (N_14681,N_14192,N_14089);
nor U14682 (N_14682,N_14314,N_14308);
nor U14683 (N_14683,N_14325,N_14441);
nor U14684 (N_14684,N_14300,N_14169);
and U14685 (N_14685,N_14403,N_14150);
nor U14686 (N_14686,N_14096,N_14026);
and U14687 (N_14687,N_14337,N_14333);
or U14688 (N_14688,N_14396,N_14497);
nor U14689 (N_14689,N_14385,N_14226);
and U14690 (N_14690,N_14310,N_14298);
nand U14691 (N_14691,N_14443,N_14336);
and U14692 (N_14692,N_14002,N_14262);
and U14693 (N_14693,N_14216,N_14436);
or U14694 (N_14694,N_14467,N_14045);
or U14695 (N_14695,N_14159,N_14207);
nor U14696 (N_14696,N_14451,N_14161);
and U14697 (N_14697,N_14028,N_14272);
or U14698 (N_14698,N_14421,N_14296);
or U14699 (N_14699,N_14112,N_14122);
and U14700 (N_14700,N_14091,N_14422);
nand U14701 (N_14701,N_14352,N_14277);
and U14702 (N_14702,N_14317,N_14398);
or U14703 (N_14703,N_14326,N_14082);
and U14704 (N_14704,N_14209,N_14486);
nor U14705 (N_14705,N_14323,N_14188);
and U14706 (N_14706,N_14231,N_14372);
nor U14707 (N_14707,N_14104,N_14268);
nand U14708 (N_14708,N_14013,N_14172);
xor U14709 (N_14709,N_14057,N_14289);
and U14710 (N_14710,N_14195,N_14064);
or U14711 (N_14711,N_14473,N_14394);
nor U14712 (N_14712,N_14168,N_14051);
or U14713 (N_14713,N_14157,N_14078);
or U14714 (N_14714,N_14149,N_14442);
nand U14715 (N_14715,N_14147,N_14202);
or U14716 (N_14716,N_14092,N_14348);
xnor U14717 (N_14717,N_14438,N_14257);
or U14718 (N_14718,N_14098,N_14101);
or U14719 (N_14719,N_14081,N_14077);
nand U14720 (N_14720,N_14014,N_14499);
nor U14721 (N_14721,N_14043,N_14318);
or U14722 (N_14722,N_14097,N_14190);
or U14723 (N_14723,N_14419,N_14175);
nor U14724 (N_14724,N_14105,N_14136);
or U14725 (N_14725,N_14402,N_14457);
and U14726 (N_14726,N_14085,N_14487);
nor U14727 (N_14727,N_14038,N_14126);
xnor U14728 (N_14728,N_14423,N_14384);
or U14729 (N_14729,N_14071,N_14371);
or U14730 (N_14730,N_14179,N_14411);
nand U14731 (N_14731,N_14405,N_14329);
nand U14732 (N_14732,N_14373,N_14469);
or U14733 (N_14733,N_14340,N_14079);
nand U14734 (N_14734,N_14431,N_14485);
or U14735 (N_14735,N_14330,N_14367);
or U14736 (N_14736,N_14235,N_14036);
and U14737 (N_14737,N_14044,N_14111);
nand U14738 (N_14738,N_14362,N_14224);
nor U14739 (N_14739,N_14090,N_14170);
nor U14740 (N_14740,N_14183,N_14491);
or U14741 (N_14741,N_14453,N_14250);
nor U14742 (N_14742,N_14007,N_14247);
and U14743 (N_14743,N_14083,N_14388);
xor U14744 (N_14744,N_14054,N_14245);
or U14745 (N_14745,N_14142,N_14282);
xor U14746 (N_14746,N_14267,N_14024);
nand U14747 (N_14747,N_14093,N_14210);
xor U14748 (N_14748,N_14119,N_14449);
and U14749 (N_14749,N_14359,N_14461);
and U14750 (N_14750,N_14424,N_14397);
nor U14751 (N_14751,N_14494,N_14057);
nor U14752 (N_14752,N_14336,N_14020);
nand U14753 (N_14753,N_14220,N_14379);
xnor U14754 (N_14754,N_14141,N_14345);
and U14755 (N_14755,N_14164,N_14405);
or U14756 (N_14756,N_14270,N_14428);
nand U14757 (N_14757,N_14353,N_14282);
nand U14758 (N_14758,N_14171,N_14142);
nor U14759 (N_14759,N_14377,N_14467);
nor U14760 (N_14760,N_14188,N_14135);
xor U14761 (N_14761,N_14391,N_14076);
nand U14762 (N_14762,N_14214,N_14267);
nor U14763 (N_14763,N_14302,N_14143);
nor U14764 (N_14764,N_14050,N_14015);
and U14765 (N_14765,N_14100,N_14210);
or U14766 (N_14766,N_14485,N_14466);
and U14767 (N_14767,N_14397,N_14057);
nand U14768 (N_14768,N_14355,N_14130);
or U14769 (N_14769,N_14172,N_14304);
nand U14770 (N_14770,N_14062,N_14068);
or U14771 (N_14771,N_14050,N_14496);
nor U14772 (N_14772,N_14468,N_14361);
or U14773 (N_14773,N_14184,N_14354);
and U14774 (N_14774,N_14408,N_14475);
xor U14775 (N_14775,N_14329,N_14241);
xor U14776 (N_14776,N_14447,N_14461);
or U14777 (N_14777,N_14265,N_14190);
nor U14778 (N_14778,N_14347,N_14118);
and U14779 (N_14779,N_14126,N_14307);
or U14780 (N_14780,N_14349,N_14459);
and U14781 (N_14781,N_14229,N_14163);
nor U14782 (N_14782,N_14266,N_14295);
xor U14783 (N_14783,N_14088,N_14233);
xnor U14784 (N_14784,N_14400,N_14090);
nand U14785 (N_14785,N_14168,N_14425);
or U14786 (N_14786,N_14207,N_14137);
or U14787 (N_14787,N_14476,N_14465);
nand U14788 (N_14788,N_14386,N_14325);
and U14789 (N_14789,N_14482,N_14145);
nor U14790 (N_14790,N_14077,N_14212);
xor U14791 (N_14791,N_14172,N_14492);
or U14792 (N_14792,N_14129,N_14110);
and U14793 (N_14793,N_14181,N_14490);
nand U14794 (N_14794,N_14281,N_14176);
xnor U14795 (N_14795,N_14420,N_14479);
and U14796 (N_14796,N_14342,N_14042);
and U14797 (N_14797,N_14400,N_14356);
or U14798 (N_14798,N_14341,N_14373);
nand U14799 (N_14799,N_14124,N_14019);
nor U14800 (N_14800,N_14109,N_14455);
nand U14801 (N_14801,N_14286,N_14168);
nor U14802 (N_14802,N_14133,N_14211);
or U14803 (N_14803,N_14317,N_14341);
nor U14804 (N_14804,N_14370,N_14142);
nand U14805 (N_14805,N_14468,N_14375);
nor U14806 (N_14806,N_14349,N_14287);
xnor U14807 (N_14807,N_14273,N_14339);
and U14808 (N_14808,N_14471,N_14156);
nand U14809 (N_14809,N_14476,N_14005);
or U14810 (N_14810,N_14176,N_14283);
or U14811 (N_14811,N_14293,N_14098);
nor U14812 (N_14812,N_14384,N_14035);
nand U14813 (N_14813,N_14062,N_14358);
and U14814 (N_14814,N_14385,N_14189);
and U14815 (N_14815,N_14446,N_14191);
and U14816 (N_14816,N_14257,N_14332);
nor U14817 (N_14817,N_14038,N_14452);
and U14818 (N_14818,N_14113,N_14070);
xnor U14819 (N_14819,N_14252,N_14275);
nor U14820 (N_14820,N_14396,N_14464);
nor U14821 (N_14821,N_14482,N_14491);
nand U14822 (N_14822,N_14325,N_14104);
nand U14823 (N_14823,N_14296,N_14103);
or U14824 (N_14824,N_14306,N_14052);
or U14825 (N_14825,N_14105,N_14143);
nand U14826 (N_14826,N_14144,N_14254);
xnor U14827 (N_14827,N_14173,N_14145);
xnor U14828 (N_14828,N_14483,N_14452);
nand U14829 (N_14829,N_14389,N_14257);
or U14830 (N_14830,N_14052,N_14271);
nand U14831 (N_14831,N_14383,N_14145);
and U14832 (N_14832,N_14142,N_14241);
and U14833 (N_14833,N_14468,N_14117);
nor U14834 (N_14834,N_14416,N_14077);
or U14835 (N_14835,N_14483,N_14386);
nor U14836 (N_14836,N_14218,N_14204);
xor U14837 (N_14837,N_14055,N_14108);
nor U14838 (N_14838,N_14402,N_14266);
or U14839 (N_14839,N_14357,N_14176);
nor U14840 (N_14840,N_14042,N_14317);
nor U14841 (N_14841,N_14090,N_14469);
nor U14842 (N_14842,N_14372,N_14415);
nand U14843 (N_14843,N_14396,N_14483);
and U14844 (N_14844,N_14128,N_14024);
and U14845 (N_14845,N_14305,N_14123);
or U14846 (N_14846,N_14121,N_14076);
nor U14847 (N_14847,N_14357,N_14207);
nor U14848 (N_14848,N_14360,N_14213);
and U14849 (N_14849,N_14056,N_14287);
or U14850 (N_14850,N_14379,N_14365);
nand U14851 (N_14851,N_14059,N_14114);
nand U14852 (N_14852,N_14169,N_14143);
nand U14853 (N_14853,N_14423,N_14382);
and U14854 (N_14854,N_14347,N_14426);
and U14855 (N_14855,N_14015,N_14383);
xor U14856 (N_14856,N_14246,N_14327);
or U14857 (N_14857,N_14119,N_14029);
or U14858 (N_14858,N_14173,N_14076);
nor U14859 (N_14859,N_14090,N_14475);
and U14860 (N_14860,N_14069,N_14430);
nand U14861 (N_14861,N_14401,N_14055);
or U14862 (N_14862,N_14133,N_14170);
nor U14863 (N_14863,N_14491,N_14363);
nor U14864 (N_14864,N_14029,N_14244);
nand U14865 (N_14865,N_14475,N_14448);
and U14866 (N_14866,N_14300,N_14402);
nand U14867 (N_14867,N_14049,N_14299);
nand U14868 (N_14868,N_14440,N_14130);
and U14869 (N_14869,N_14395,N_14231);
and U14870 (N_14870,N_14316,N_14014);
or U14871 (N_14871,N_14075,N_14000);
nand U14872 (N_14872,N_14128,N_14349);
and U14873 (N_14873,N_14338,N_14456);
and U14874 (N_14874,N_14323,N_14088);
or U14875 (N_14875,N_14298,N_14363);
nand U14876 (N_14876,N_14305,N_14130);
nor U14877 (N_14877,N_14138,N_14159);
or U14878 (N_14878,N_14196,N_14260);
or U14879 (N_14879,N_14123,N_14310);
nor U14880 (N_14880,N_14400,N_14115);
and U14881 (N_14881,N_14278,N_14251);
nand U14882 (N_14882,N_14391,N_14195);
nor U14883 (N_14883,N_14138,N_14198);
xnor U14884 (N_14884,N_14139,N_14279);
and U14885 (N_14885,N_14320,N_14130);
nor U14886 (N_14886,N_14149,N_14045);
and U14887 (N_14887,N_14241,N_14038);
nand U14888 (N_14888,N_14237,N_14437);
or U14889 (N_14889,N_14455,N_14333);
and U14890 (N_14890,N_14260,N_14164);
or U14891 (N_14891,N_14109,N_14346);
or U14892 (N_14892,N_14059,N_14062);
or U14893 (N_14893,N_14164,N_14025);
or U14894 (N_14894,N_14175,N_14203);
nand U14895 (N_14895,N_14312,N_14351);
nor U14896 (N_14896,N_14096,N_14070);
and U14897 (N_14897,N_14147,N_14096);
nand U14898 (N_14898,N_14429,N_14017);
nor U14899 (N_14899,N_14309,N_14224);
xor U14900 (N_14900,N_14444,N_14210);
nor U14901 (N_14901,N_14443,N_14360);
nor U14902 (N_14902,N_14089,N_14439);
or U14903 (N_14903,N_14448,N_14405);
xnor U14904 (N_14904,N_14158,N_14369);
nand U14905 (N_14905,N_14345,N_14414);
xnor U14906 (N_14906,N_14142,N_14207);
nand U14907 (N_14907,N_14065,N_14032);
nand U14908 (N_14908,N_14485,N_14432);
xnor U14909 (N_14909,N_14028,N_14296);
or U14910 (N_14910,N_14418,N_14320);
nand U14911 (N_14911,N_14102,N_14046);
or U14912 (N_14912,N_14085,N_14050);
or U14913 (N_14913,N_14361,N_14339);
and U14914 (N_14914,N_14195,N_14366);
xor U14915 (N_14915,N_14108,N_14459);
and U14916 (N_14916,N_14272,N_14288);
and U14917 (N_14917,N_14018,N_14260);
nor U14918 (N_14918,N_14017,N_14307);
and U14919 (N_14919,N_14117,N_14206);
or U14920 (N_14920,N_14234,N_14006);
nand U14921 (N_14921,N_14285,N_14413);
xnor U14922 (N_14922,N_14474,N_14472);
nor U14923 (N_14923,N_14338,N_14430);
and U14924 (N_14924,N_14409,N_14336);
and U14925 (N_14925,N_14327,N_14063);
or U14926 (N_14926,N_14151,N_14157);
or U14927 (N_14927,N_14470,N_14133);
and U14928 (N_14928,N_14212,N_14179);
and U14929 (N_14929,N_14101,N_14484);
or U14930 (N_14930,N_14398,N_14006);
nand U14931 (N_14931,N_14157,N_14267);
and U14932 (N_14932,N_14238,N_14115);
nor U14933 (N_14933,N_14332,N_14027);
or U14934 (N_14934,N_14069,N_14030);
or U14935 (N_14935,N_14382,N_14371);
nand U14936 (N_14936,N_14008,N_14292);
nor U14937 (N_14937,N_14045,N_14321);
or U14938 (N_14938,N_14098,N_14413);
and U14939 (N_14939,N_14475,N_14323);
xor U14940 (N_14940,N_14266,N_14099);
nand U14941 (N_14941,N_14131,N_14365);
nor U14942 (N_14942,N_14489,N_14248);
and U14943 (N_14943,N_14274,N_14388);
nand U14944 (N_14944,N_14018,N_14329);
or U14945 (N_14945,N_14073,N_14116);
xor U14946 (N_14946,N_14331,N_14219);
nor U14947 (N_14947,N_14209,N_14087);
or U14948 (N_14948,N_14404,N_14135);
or U14949 (N_14949,N_14103,N_14312);
nand U14950 (N_14950,N_14238,N_14443);
nand U14951 (N_14951,N_14165,N_14245);
xor U14952 (N_14952,N_14440,N_14344);
and U14953 (N_14953,N_14199,N_14076);
nor U14954 (N_14954,N_14395,N_14096);
nor U14955 (N_14955,N_14173,N_14243);
and U14956 (N_14956,N_14424,N_14028);
nand U14957 (N_14957,N_14129,N_14381);
nor U14958 (N_14958,N_14317,N_14220);
xnor U14959 (N_14959,N_14400,N_14443);
nand U14960 (N_14960,N_14196,N_14362);
or U14961 (N_14961,N_14435,N_14482);
nand U14962 (N_14962,N_14499,N_14124);
and U14963 (N_14963,N_14404,N_14125);
nand U14964 (N_14964,N_14487,N_14228);
or U14965 (N_14965,N_14194,N_14030);
or U14966 (N_14966,N_14190,N_14020);
or U14967 (N_14967,N_14200,N_14160);
and U14968 (N_14968,N_14347,N_14144);
xnor U14969 (N_14969,N_14172,N_14008);
xnor U14970 (N_14970,N_14430,N_14409);
and U14971 (N_14971,N_14317,N_14202);
or U14972 (N_14972,N_14383,N_14167);
nor U14973 (N_14973,N_14333,N_14078);
and U14974 (N_14974,N_14084,N_14001);
nand U14975 (N_14975,N_14244,N_14037);
nor U14976 (N_14976,N_14165,N_14369);
nand U14977 (N_14977,N_14484,N_14088);
and U14978 (N_14978,N_14108,N_14126);
or U14979 (N_14979,N_14033,N_14401);
or U14980 (N_14980,N_14302,N_14252);
or U14981 (N_14981,N_14308,N_14180);
xnor U14982 (N_14982,N_14433,N_14313);
nand U14983 (N_14983,N_14196,N_14018);
nor U14984 (N_14984,N_14144,N_14353);
nor U14985 (N_14985,N_14186,N_14232);
nand U14986 (N_14986,N_14422,N_14041);
or U14987 (N_14987,N_14442,N_14153);
nor U14988 (N_14988,N_14081,N_14291);
nand U14989 (N_14989,N_14346,N_14330);
and U14990 (N_14990,N_14485,N_14230);
or U14991 (N_14991,N_14300,N_14420);
and U14992 (N_14992,N_14442,N_14013);
and U14993 (N_14993,N_14377,N_14281);
nor U14994 (N_14994,N_14092,N_14239);
and U14995 (N_14995,N_14186,N_14378);
or U14996 (N_14996,N_14239,N_14166);
nor U14997 (N_14997,N_14394,N_14039);
nor U14998 (N_14998,N_14495,N_14074);
and U14999 (N_14999,N_14251,N_14317);
or UO_0 (O_0,N_14611,N_14687);
or UO_1 (O_1,N_14582,N_14524);
or UO_2 (O_2,N_14844,N_14558);
nor UO_3 (O_3,N_14994,N_14652);
or UO_4 (O_4,N_14911,N_14672);
or UO_5 (O_5,N_14602,N_14834);
nand UO_6 (O_6,N_14995,N_14860);
xor UO_7 (O_7,N_14557,N_14545);
nand UO_8 (O_8,N_14610,N_14749);
and UO_9 (O_9,N_14768,N_14746);
nand UO_10 (O_10,N_14991,N_14638);
and UO_11 (O_11,N_14907,N_14806);
or UO_12 (O_12,N_14777,N_14579);
nand UO_13 (O_13,N_14724,N_14893);
and UO_14 (O_14,N_14862,N_14967);
or UO_15 (O_15,N_14658,N_14581);
nand UO_16 (O_16,N_14644,N_14521);
nor UO_17 (O_17,N_14881,N_14641);
and UO_18 (O_18,N_14504,N_14739);
nor UO_19 (O_19,N_14536,N_14629);
nor UO_20 (O_20,N_14964,N_14717);
and UO_21 (O_21,N_14515,N_14925);
nor UO_22 (O_22,N_14503,N_14999);
or UO_23 (O_23,N_14510,N_14904);
xor UO_24 (O_24,N_14623,N_14661);
nor UO_25 (O_25,N_14670,N_14526);
nor UO_26 (O_26,N_14896,N_14952);
nand UO_27 (O_27,N_14955,N_14659);
and UO_28 (O_28,N_14795,N_14802);
and UO_29 (O_29,N_14772,N_14851);
and UO_30 (O_30,N_14981,N_14666);
nor UO_31 (O_31,N_14554,N_14722);
nor UO_32 (O_32,N_14946,N_14702);
nand UO_33 (O_33,N_14756,N_14514);
or UO_34 (O_34,N_14870,N_14742);
and UO_35 (O_35,N_14609,N_14842);
nor UO_36 (O_36,N_14520,N_14616);
and UO_37 (O_37,N_14958,N_14596);
nor UO_38 (O_38,N_14797,N_14636);
nand UO_39 (O_39,N_14729,N_14978);
nand UO_40 (O_40,N_14854,N_14956);
or UO_41 (O_41,N_14940,N_14643);
or UO_42 (O_42,N_14732,N_14827);
xnor UO_43 (O_43,N_14556,N_14892);
xor UO_44 (O_44,N_14605,N_14875);
xor UO_45 (O_45,N_14776,N_14818);
or UO_46 (O_46,N_14678,N_14538);
and UO_47 (O_47,N_14712,N_14752);
or UO_48 (O_48,N_14968,N_14608);
nand UO_49 (O_49,N_14976,N_14511);
nand UO_50 (O_50,N_14668,N_14762);
nor UO_51 (O_51,N_14576,N_14792);
nand UO_52 (O_52,N_14790,N_14694);
and UO_53 (O_53,N_14548,N_14998);
nand UO_54 (O_54,N_14954,N_14509);
nand UO_55 (O_55,N_14778,N_14810);
nand UO_56 (O_56,N_14690,N_14734);
or UO_57 (O_57,N_14552,N_14866);
and UO_58 (O_58,N_14537,N_14513);
nor UO_59 (O_59,N_14615,N_14915);
nor UO_60 (O_60,N_14848,N_14764);
or UO_61 (O_61,N_14714,N_14603);
or UO_62 (O_62,N_14905,N_14938);
or UO_63 (O_63,N_14728,N_14950);
nor UO_64 (O_64,N_14760,N_14523);
nand UO_65 (O_65,N_14721,N_14698);
nor UO_66 (O_66,N_14829,N_14787);
or UO_67 (O_67,N_14727,N_14701);
or UO_68 (O_68,N_14689,N_14990);
and UO_69 (O_69,N_14750,N_14540);
and UO_70 (O_70,N_14805,N_14933);
xnor UO_71 (O_71,N_14757,N_14819);
nor UO_72 (O_72,N_14686,N_14913);
nand UO_73 (O_73,N_14944,N_14949);
nand UO_74 (O_74,N_14912,N_14997);
or UO_75 (O_75,N_14826,N_14630);
nand UO_76 (O_76,N_14989,N_14931);
xnor UO_77 (O_77,N_14561,N_14679);
xor UO_78 (O_78,N_14709,N_14879);
or UO_79 (O_79,N_14830,N_14909);
or UO_80 (O_80,N_14871,N_14535);
or UO_81 (O_81,N_14857,N_14974);
nand UO_82 (O_82,N_14707,N_14917);
xnor UO_83 (O_83,N_14626,N_14841);
and UO_84 (O_84,N_14799,N_14584);
xor UO_85 (O_85,N_14745,N_14662);
or UO_86 (O_86,N_14985,N_14527);
and UO_87 (O_87,N_14575,N_14634);
nand UO_88 (O_88,N_14858,N_14577);
and UO_89 (O_89,N_14885,N_14651);
and UO_90 (O_90,N_14755,N_14657);
and UO_91 (O_91,N_14977,N_14720);
nand UO_92 (O_92,N_14785,N_14606);
or UO_93 (O_93,N_14780,N_14895);
nand UO_94 (O_94,N_14519,N_14861);
nand UO_95 (O_95,N_14637,N_14649);
xnor UO_96 (O_96,N_14867,N_14684);
and UO_97 (O_97,N_14525,N_14864);
nor UO_98 (O_98,N_14716,N_14766);
or UO_99 (O_99,N_14595,N_14664);
and UO_100 (O_100,N_14803,N_14617);
and UO_101 (O_101,N_14840,N_14839);
and UO_102 (O_102,N_14823,N_14965);
and UO_103 (O_103,N_14683,N_14816);
or UO_104 (O_104,N_14673,N_14979);
or UO_105 (O_105,N_14969,N_14522);
nor UO_106 (O_106,N_14599,N_14927);
or UO_107 (O_107,N_14531,N_14770);
nand UO_108 (O_108,N_14922,N_14835);
and UO_109 (O_109,N_14568,N_14972);
xor UO_110 (O_110,N_14975,N_14753);
nand UO_111 (O_111,N_14593,N_14831);
or UO_112 (O_112,N_14551,N_14783);
and UO_113 (O_113,N_14718,N_14902);
or UO_114 (O_114,N_14982,N_14853);
nand UO_115 (O_115,N_14529,N_14500);
nand UO_116 (O_116,N_14663,N_14627);
nor UO_117 (O_117,N_14656,N_14872);
or UO_118 (O_118,N_14733,N_14624);
or UO_119 (O_119,N_14594,N_14894);
nor UO_120 (O_120,N_14947,N_14685);
nand UO_121 (O_121,N_14639,N_14948);
nor UO_122 (O_122,N_14889,N_14920);
nor UO_123 (O_123,N_14587,N_14801);
xor UO_124 (O_124,N_14983,N_14674);
or UO_125 (O_125,N_14758,N_14695);
or UO_126 (O_126,N_14773,N_14546);
nand UO_127 (O_127,N_14725,N_14574);
nor UO_128 (O_128,N_14993,N_14859);
nor UO_129 (O_129,N_14719,N_14597);
and UO_130 (O_130,N_14846,N_14754);
nor UO_131 (O_131,N_14507,N_14887);
nand UO_132 (O_132,N_14929,N_14980);
and UO_133 (O_133,N_14761,N_14696);
and UO_134 (O_134,N_14843,N_14618);
or UO_135 (O_135,N_14547,N_14622);
nor UO_136 (O_136,N_14585,N_14880);
or UO_137 (O_137,N_14660,N_14533);
nor UO_138 (O_138,N_14992,N_14647);
xnor UO_139 (O_139,N_14650,N_14808);
nor UO_140 (O_140,N_14788,N_14731);
nor UO_141 (O_141,N_14555,N_14934);
nor UO_142 (O_142,N_14607,N_14769);
nand UO_143 (O_143,N_14781,N_14693);
and UO_144 (O_144,N_14804,N_14868);
nor UO_145 (O_145,N_14563,N_14936);
or UO_146 (O_146,N_14910,N_14899);
nor UO_147 (O_147,N_14916,N_14648);
nor UO_148 (O_148,N_14655,N_14665);
or UO_149 (O_149,N_14821,N_14502);
or UO_150 (O_150,N_14580,N_14653);
or UO_151 (O_151,N_14759,N_14633);
nor UO_152 (O_152,N_14744,N_14971);
and UO_153 (O_153,N_14682,N_14571);
nand UO_154 (O_154,N_14970,N_14619);
and UO_155 (O_155,N_14713,N_14614);
nor UO_156 (O_156,N_14937,N_14628);
and UO_157 (O_157,N_14621,N_14751);
or UO_158 (O_158,N_14506,N_14923);
and UO_159 (O_159,N_14960,N_14932);
nand UO_160 (O_160,N_14850,N_14836);
or UO_161 (O_161,N_14539,N_14681);
nor UO_162 (O_162,N_14996,N_14908);
and UO_163 (O_163,N_14570,N_14530);
nand UO_164 (O_164,N_14706,N_14919);
nand UO_165 (O_165,N_14784,N_14847);
xnor UO_166 (O_166,N_14833,N_14849);
or UO_167 (O_167,N_14928,N_14914);
and UO_168 (O_168,N_14508,N_14926);
and UO_169 (O_169,N_14988,N_14640);
or UO_170 (O_170,N_14863,N_14562);
xor UO_171 (O_171,N_14737,N_14874);
xnor UO_172 (O_172,N_14765,N_14962);
nor UO_173 (O_173,N_14884,N_14959);
and UO_174 (O_174,N_14957,N_14815);
xnor UO_175 (O_175,N_14898,N_14945);
and UO_176 (O_176,N_14730,N_14569);
nand UO_177 (O_177,N_14921,N_14900);
and UO_178 (O_178,N_14961,N_14505);
and UO_179 (O_179,N_14812,N_14883);
and UO_180 (O_180,N_14817,N_14735);
and UO_181 (O_181,N_14501,N_14855);
and UO_182 (O_182,N_14986,N_14963);
and UO_183 (O_183,N_14924,N_14930);
nor UO_184 (O_184,N_14943,N_14631);
or UO_185 (O_185,N_14973,N_14567);
nor UO_186 (O_186,N_14612,N_14676);
nand UO_187 (O_187,N_14942,N_14680);
nor UO_188 (O_188,N_14691,N_14748);
nor UO_189 (O_189,N_14856,N_14573);
nand UO_190 (O_190,N_14620,N_14953);
and UO_191 (O_191,N_14796,N_14590);
nor UO_192 (O_192,N_14700,N_14632);
or UO_193 (O_193,N_14869,N_14743);
nand UO_194 (O_194,N_14786,N_14542);
xor UO_195 (O_195,N_14708,N_14791);
nand UO_196 (O_196,N_14876,N_14534);
and UO_197 (O_197,N_14688,N_14935);
or UO_198 (O_198,N_14873,N_14891);
nand UO_199 (O_199,N_14793,N_14877);
nor UO_200 (O_200,N_14984,N_14888);
nand UO_201 (O_201,N_14583,N_14820);
nor UO_202 (O_202,N_14794,N_14882);
or UO_203 (O_203,N_14771,N_14966);
nand UO_204 (O_204,N_14782,N_14565);
nor UO_205 (O_205,N_14604,N_14951);
or UO_206 (O_206,N_14941,N_14711);
or UO_207 (O_207,N_14901,N_14591);
nor UO_208 (O_208,N_14897,N_14903);
or UO_209 (O_209,N_14738,N_14890);
xnor UO_210 (O_210,N_14852,N_14559);
nand UO_211 (O_211,N_14800,N_14763);
and UO_212 (O_212,N_14811,N_14517);
nand UO_213 (O_213,N_14838,N_14550);
and UO_214 (O_214,N_14532,N_14704);
xor UO_215 (O_215,N_14518,N_14886);
nor UO_216 (O_216,N_14807,N_14588);
nand UO_217 (O_217,N_14809,N_14592);
nor UO_218 (O_218,N_14814,N_14825);
or UO_219 (O_219,N_14705,N_14699);
nand UO_220 (O_220,N_14822,N_14645);
xnor UO_221 (O_221,N_14779,N_14544);
nand UO_222 (O_222,N_14723,N_14703);
xnor UO_223 (O_223,N_14560,N_14528);
and UO_224 (O_224,N_14667,N_14516);
nor UO_225 (O_225,N_14669,N_14837);
or UO_226 (O_226,N_14878,N_14543);
and UO_227 (O_227,N_14767,N_14813);
and UO_228 (O_228,N_14613,N_14541);
or UO_229 (O_229,N_14601,N_14635);
nand UO_230 (O_230,N_14600,N_14747);
nand UO_231 (O_231,N_14987,N_14589);
nor UO_232 (O_232,N_14646,N_14906);
and UO_233 (O_233,N_14715,N_14671);
nand UO_234 (O_234,N_14845,N_14586);
xnor UO_235 (O_235,N_14572,N_14774);
and UO_236 (O_236,N_14512,N_14710);
and UO_237 (O_237,N_14775,N_14654);
and UO_238 (O_238,N_14789,N_14798);
and UO_239 (O_239,N_14832,N_14824);
nand UO_240 (O_240,N_14578,N_14564);
and UO_241 (O_241,N_14939,N_14549);
nor UO_242 (O_242,N_14553,N_14697);
and UO_243 (O_243,N_14625,N_14740);
or UO_244 (O_244,N_14677,N_14736);
nand UO_245 (O_245,N_14741,N_14566);
or UO_246 (O_246,N_14675,N_14726);
nor UO_247 (O_247,N_14828,N_14865);
or UO_248 (O_248,N_14642,N_14692);
and UO_249 (O_249,N_14598,N_14918);
or UO_250 (O_250,N_14851,N_14771);
or UO_251 (O_251,N_14829,N_14904);
nand UO_252 (O_252,N_14829,N_14600);
or UO_253 (O_253,N_14975,N_14676);
and UO_254 (O_254,N_14893,N_14604);
nand UO_255 (O_255,N_14726,N_14759);
xor UO_256 (O_256,N_14731,N_14724);
xor UO_257 (O_257,N_14632,N_14959);
nand UO_258 (O_258,N_14547,N_14781);
nor UO_259 (O_259,N_14605,N_14937);
or UO_260 (O_260,N_14983,N_14570);
and UO_261 (O_261,N_14744,N_14812);
or UO_262 (O_262,N_14789,N_14554);
nand UO_263 (O_263,N_14523,N_14679);
nand UO_264 (O_264,N_14558,N_14565);
and UO_265 (O_265,N_14787,N_14519);
or UO_266 (O_266,N_14719,N_14634);
nand UO_267 (O_267,N_14709,N_14764);
or UO_268 (O_268,N_14929,N_14711);
xor UO_269 (O_269,N_14982,N_14785);
and UO_270 (O_270,N_14664,N_14931);
nand UO_271 (O_271,N_14880,N_14752);
and UO_272 (O_272,N_14796,N_14953);
nor UO_273 (O_273,N_14936,N_14692);
nand UO_274 (O_274,N_14879,N_14972);
nand UO_275 (O_275,N_14622,N_14958);
nor UO_276 (O_276,N_14837,N_14676);
nor UO_277 (O_277,N_14918,N_14731);
or UO_278 (O_278,N_14571,N_14725);
and UO_279 (O_279,N_14553,N_14668);
nand UO_280 (O_280,N_14676,N_14719);
nand UO_281 (O_281,N_14677,N_14955);
and UO_282 (O_282,N_14873,N_14961);
or UO_283 (O_283,N_14601,N_14667);
or UO_284 (O_284,N_14995,N_14800);
nor UO_285 (O_285,N_14657,N_14674);
nor UO_286 (O_286,N_14964,N_14734);
or UO_287 (O_287,N_14631,N_14893);
or UO_288 (O_288,N_14639,N_14675);
nand UO_289 (O_289,N_14741,N_14534);
and UO_290 (O_290,N_14636,N_14685);
nand UO_291 (O_291,N_14981,N_14610);
nand UO_292 (O_292,N_14973,N_14680);
or UO_293 (O_293,N_14592,N_14693);
nand UO_294 (O_294,N_14851,N_14995);
nor UO_295 (O_295,N_14862,N_14692);
and UO_296 (O_296,N_14533,N_14560);
nand UO_297 (O_297,N_14550,N_14708);
or UO_298 (O_298,N_14619,N_14921);
xor UO_299 (O_299,N_14574,N_14654);
and UO_300 (O_300,N_14794,N_14644);
or UO_301 (O_301,N_14787,N_14690);
nor UO_302 (O_302,N_14745,N_14645);
or UO_303 (O_303,N_14586,N_14782);
or UO_304 (O_304,N_14518,N_14907);
and UO_305 (O_305,N_14510,N_14823);
xnor UO_306 (O_306,N_14962,N_14699);
and UO_307 (O_307,N_14940,N_14911);
xor UO_308 (O_308,N_14766,N_14810);
nor UO_309 (O_309,N_14764,N_14628);
or UO_310 (O_310,N_14816,N_14896);
xor UO_311 (O_311,N_14583,N_14877);
or UO_312 (O_312,N_14785,N_14592);
and UO_313 (O_313,N_14915,N_14538);
or UO_314 (O_314,N_14956,N_14539);
and UO_315 (O_315,N_14938,N_14876);
nor UO_316 (O_316,N_14756,N_14853);
nand UO_317 (O_317,N_14634,N_14715);
nor UO_318 (O_318,N_14988,N_14762);
nand UO_319 (O_319,N_14538,N_14509);
nand UO_320 (O_320,N_14685,N_14961);
nor UO_321 (O_321,N_14701,N_14625);
nor UO_322 (O_322,N_14959,N_14523);
xor UO_323 (O_323,N_14868,N_14867);
nand UO_324 (O_324,N_14882,N_14890);
or UO_325 (O_325,N_14969,N_14795);
nand UO_326 (O_326,N_14906,N_14984);
and UO_327 (O_327,N_14615,N_14916);
nand UO_328 (O_328,N_14812,N_14941);
nor UO_329 (O_329,N_14928,N_14649);
and UO_330 (O_330,N_14821,N_14762);
nor UO_331 (O_331,N_14895,N_14659);
or UO_332 (O_332,N_14913,N_14788);
nand UO_333 (O_333,N_14805,N_14903);
and UO_334 (O_334,N_14875,N_14704);
and UO_335 (O_335,N_14784,N_14740);
nor UO_336 (O_336,N_14710,N_14596);
nand UO_337 (O_337,N_14991,N_14518);
xnor UO_338 (O_338,N_14549,N_14763);
nand UO_339 (O_339,N_14988,N_14930);
xnor UO_340 (O_340,N_14640,N_14925);
and UO_341 (O_341,N_14813,N_14838);
nand UO_342 (O_342,N_14921,N_14920);
nand UO_343 (O_343,N_14569,N_14508);
or UO_344 (O_344,N_14743,N_14977);
nand UO_345 (O_345,N_14682,N_14615);
or UO_346 (O_346,N_14742,N_14762);
nand UO_347 (O_347,N_14681,N_14652);
nand UO_348 (O_348,N_14787,N_14761);
nor UO_349 (O_349,N_14805,N_14544);
or UO_350 (O_350,N_14781,N_14590);
nor UO_351 (O_351,N_14657,N_14843);
and UO_352 (O_352,N_14517,N_14787);
nand UO_353 (O_353,N_14526,N_14517);
and UO_354 (O_354,N_14680,N_14593);
or UO_355 (O_355,N_14681,N_14830);
or UO_356 (O_356,N_14509,N_14686);
nor UO_357 (O_357,N_14958,N_14985);
nor UO_358 (O_358,N_14851,N_14528);
and UO_359 (O_359,N_14620,N_14667);
nor UO_360 (O_360,N_14890,N_14930);
xnor UO_361 (O_361,N_14641,N_14774);
and UO_362 (O_362,N_14507,N_14716);
or UO_363 (O_363,N_14862,N_14508);
xor UO_364 (O_364,N_14737,N_14970);
or UO_365 (O_365,N_14987,N_14583);
or UO_366 (O_366,N_14776,N_14555);
and UO_367 (O_367,N_14705,N_14698);
or UO_368 (O_368,N_14629,N_14906);
xnor UO_369 (O_369,N_14529,N_14783);
xnor UO_370 (O_370,N_14819,N_14577);
and UO_371 (O_371,N_14641,N_14555);
nand UO_372 (O_372,N_14649,N_14690);
or UO_373 (O_373,N_14690,N_14955);
nor UO_374 (O_374,N_14605,N_14518);
nor UO_375 (O_375,N_14931,N_14638);
nor UO_376 (O_376,N_14761,N_14862);
nor UO_377 (O_377,N_14859,N_14525);
nor UO_378 (O_378,N_14564,N_14764);
and UO_379 (O_379,N_14888,N_14852);
nand UO_380 (O_380,N_14629,N_14524);
or UO_381 (O_381,N_14885,N_14807);
nor UO_382 (O_382,N_14970,N_14667);
xor UO_383 (O_383,N_14699,N_14716);
xor UO_384 (O_384,N_14742,N_14930);
xnor UO_385 (O_385,N_14716,N_14926);
nand UO_386 (O_386,N_14888,N_14948);
nand UO_387 (O_387,N_14870,N_14734);
nand UO_388 (O_388,N_14684,N_14784);
xor UO_389 (O_389,N_14717,N_14639);
nand UO_390 (O_390,N_14774,N_14734);
and UO_391 (O_391,N_14928,N_14623);
and UO_392 (O_392,N_14515,N_14501);
or UO_393 (O_393,N_14569,N_14928);
nor UO_394 (O_394,N_14534,N_14644);
and UO_395 (O_395,N_14619,N_14768);
and UO_396 (O_396,N_14664,N_14841);
nand UO_397 (O_397,N_14945,N_14869);
nor UO_398 (O_398,N_14961,N_14569);
nor UO_399 (O_399,N_14986,N_14720);
nand UO_400 (O_400,N_14761,N_14519);
nand UO_401 (O_401,N_14763,N_14911);
or UO_402 (O_402,N_14832,N_14701);
and UO_403 (O_403,N_14690,N_14856);
nand UO_404 (O_404,N_14785,N_14543);
and UO_405 (O_405,N_14534,N_14613);
nand UO_406 (O_406,N_14537,N_14927);
nand UO_407 (O_407,N_14788,N_14510);
nor UO_408 (O_408,N_14703,N_14789);
and UO_409 (O_409,N_14590,N_14777);
nand UO_410 (O_410,N_14807,N_14672);
nor UO_411 (O_411,N_14767,N_14569);
xor UO_412 (O_412,N_14547,N_14964);
and UO_413 (O_413,N_14509,N_14849);
or UO_414 (O_414,N_14997,N_14601);
nor UO_415 (O_415,N_14835,N_14526);
nand UO_416 (O_416,N_14623,N_14756);
nand UO_417 (O_417,N_14609,N_14714);
nor UO_418 (O_418,N_14809,N_14509);
or UO_419 (O_419,N_14712,N_14806);
and UO_420 (O_420,N_14962,N_14719);
nand UO_421 (O_421,N_14909,N_14770);
nand UO_422 (O_422,N_14680,N_14641);
nand UO_423 (O_423,N_14678,N_14671);
nor UO_424 (O_424,N_14892,N_14715);
nor UO_425 (O_425,N_14658,N_14710);
nand UO_426 (O_426,N_14759,N_14594);
or UO_427 (O_427,N_14660,N_14767);
xnor UO_428 (O_428,N_14715,N_14569);
or UO_429 (O_429,N_14826,N_14774);
nor UO_430 (O_430,N_14646,N_14853);
and UO_431 (O_431,N_14691,N_14811);
nor UO_432 (O_432,N_14775,N_14810);
nor UO_433 (O_433,N_14706,N_14691);
and UO_434 (O_434,N_14673,N_14899);
nand UO_435 (O_435,N_14695,N_14770);
or UO_436 (O_436,N_14980,N_14635);
or UO_437 (O_437,N_14920,N_14806);
xor UO_438 (O_438,N_14893,N_14925);
and UO_439 (O_439,N_14816,N_14941);
nand UO_440 (O_440,N_14544,N_14711);
nand UO_441 (O_441,N_14628,N_14558);
and UO_442 (O_442,N_14500,N_14919);
nand UO_443 (O_443,N_14552,N_14830);
nand UO_444 (O_444,N_14677,N_14860);
nand UO_445 (O_445,N_14600,N_14882);
or UO_446 (O_446,N_14814,N_14813);
nand UO_447 (O_447,N_14591,N_14877);
and UO_448 (O_448,N_14758,N_14869);
nand UO_449 (O_449,N_14855,N_14657);
nor UO_450 (O_450,N_14732,N_14863);
or UO_451 (O_451,N_14794,N_14838);
or UO_452 (O_452,N_14655,N_14656);
xnor UO_453 (O_453,N_14525,N_14722);
and UO_454 (O_454,N_14800,N_14930);
or UO_455 (O_455,N_14853,N_14882);
or UO_456 (O_456,N_14694,N_14677);
and UO_457 (O_457,N_14530,N_14575);
nor UO_458 (O_458,N_14879,N_14922);
nand UO_459 (O_459,N_14962,N_14984);
and UO_460 (O_460,N_14749,N_14501);
and UO_461 (O_461,N_14558,N_14692);
nor UO_462 (O_462,N_14963,N_14953);
nand UO_463 (O_463,N_14681,N_14819);
or UO_464 (O_464,N_14616,N_14702);
nand UO_465 (O_465,N_14936,N_14965);
and UO_466 (O_466,N_14881,N_14546);
nand UO_467 (O_467,N_14803,N_14519);
nor UO_468 (O_468,N_14625,N_14561);
nor UO_469 (O_469,N_14702,N_14818);
and UO_470 (O_470,N_14790,N_14863);
and UO_471 (O_471,N_14555,N_14862);
and UO_472 (O_472,N_14820,N_14722);
xnor UO_473 (O_473,N_14757,N_14810);
nor UO_474 (O_474,N_14743,N_14598);
nand UO_475 (O_475,N_14591,N_14857);
and UO_476 (O_476,N_14774,N_14807);
or UO_477 (O_477,N_14891,N_14505);
nand UO_478 (O_478,N_14950,N_14511);
and UO_479 (O_479,N_14631,N_14829);
xor UO_480 (O_480,N_14715,N_14511);
or UO_481 (O_481,N_14755,N_14830);
and UO_482 (O_482,N_14953,N_14830);
nand UO_483 (O_483,N_14516,N_14868);
nand UO_484 (O_484,N_14513,N_14968);
and UO_485 (O_485,N_14974,N_14955);
nor UO_486 (O_486,N_14588,N_14962);
nor UO_487 (O_487,N_14956,N_14585);
or UO_488 (O_488,N_14717,N_14676);
or UO_489 (O_489,N_14745,N_14516);
nand UO_490 (O_490,N_14641,N_14893);
and UO_491 (O_491,N_14501,N_14733);
or UO_492 (O_492,N_14617,N_14795);
and UO_493 (O_493,N_14795,N_14997);
nand UO_494 (O_494,N_14744,N_14730);
and UO_495 (O_495,N_14562,N_14855);
xnor UO_496 (O_496,N_14697,N_14765);
xnor UO_497 (O_497,N_14817,N_14613);
or UO_498 (O_498,N_14639,N_14602);
or UO_499 (O_499,N_14529,N_14597);
or UO_500 (O_500,N_14595,N_14785);
and UO_501 (O_501,N_14678,N_14654);
nand UO_502 (O_502,N_14942,N_14752);
xor UO_503 (O_503,N_14756,N_14604);
nor UO_504 (O_504,N_14987,N_14962);
xnor UO_505 (O_505,N_14538,N_14650);
or UO_506 (O_506,N_14730,N_14941);
or UO_507 (O_507,N_14949,N_14579);
and UO_508 (O_508,N_14918,N_14742);
or UO_509 (O_509,N_14932,N_14828);
or UO_510 (O_510,N_14855,N_14616);
nand UO_511 (O_511,N_14723,N_14781);
or UO_512 (O_512,N_14716,N_14735);
nor UO_513 (O_513,N_14969,N_14851);
nand UO_514 (O_514,N_14924,N_14800);
xor UO_515 (O_515,N_14858,N_14882);
nor UO_516 (O_516,N_14509,N_14725);
and UO_517 (O_517,N_14636,N_14887);
nand UO_518 (O_518,N_14804,N_14803);
or UO_519 (O_519,N_14603,N_14720);
or UO_520 (O_520,N_14772,N_14545);
or UO_521 (O_521,N_14911,N_14552);
nor UO_522 (O_522,N_14838,N_14859);
and UO_523 (O_523,N_14633,N_14891);
nand UO_524 (O_524,N_14801,N_14781);
nand UO_525 (O_525,N_14731,N_14945);
and UO_526 (O_526,N_14769,N_14834);
xor UO_527 (O_527,N_14732,N_14635);
or UO_528 (O_528,N_14574,N_14886);
nand UO_529 (O_529,N_14837,N_14532);
or UO_530 (O_530,N_14746,N_14958);
nand UO_531 (O_531,N_14781,N_14606);
or UO_532 (O_532,N_14626,N_14714);
nor UO_533 (O_533,N_14744,N_14993);
or UO_534 (O_534,N_14587,N_14629);
nor UO_535 (O_535,N_14859,N_14545);
or UO_536 (O_536,N_14787,N_14974);
nor UO_537 (O_537,N_14592,N_14751);
or UO_538 (O_538,N_14831,N_14788);
nor UO_539 (O_539,N_14805,N_14681);
nand UO_540 (O_540,N_14533,N_14905);
nand UO_541 (O_541,N_14960,N_14966);
and UO_542 (O_542,N_14556,N_14842);
or UO_543 (O_543,N_14839,N_14896);
xnor UO_544 (O_544,N_14715,N_14888);
nand UO_545 (O_545,N_14512,N_14560);
xnor UO_546 (O_546,N_14943,N_14720);
nand UO_547 (O_547,N_14631,N_14572);
or UO_548 (O_548,N_14846,N_14944);
nor UO_549 (O_549,N_14805,N_14524);
or UO_550 (O_550,N_14707,N_14797);
nor UO_551 (O_551,N_14617,N_14573);
nor UO_552 (O_552,N_14844,N_14858);
nor UO_553 (O_553,N_14505,N_14810);
xor UO_554 (O_554,N_14574,N_14778);
nor UO_555 (O_555,N_14554,N_14693);
or UO_556 (O_556,N_14838,N_14809);
nand UO_557 (O_557,N_14792,N_14687);
or UO_558 (O_558,N_14738,N_14730);
and UO_559 (O_559,N_14569,N_14971);
and UO_560 (O_560,N_14617,N_14970);
or UO_561 (O_561,N_14583,N_14631);
nand UO_562 (O_562,N_14996,N_14729);
or UO_563 (O_563,N_14554,N_14670);
and UO_564 (O_564,N_14728,N_14769);
nor UO_565 (O_565,N_14585,N_14523);
xnor UO_566 (O_566,N_14643,N_14914);
nor UO_567 (O_567,N_14808,N_14680);
nand UO_568 (O_568,N_14744,N_14619);
nor UO_569 (O_569,N_14776,N_14728);
and UO_570 (O_570,N_14654,N_14622);
nand UO_571 (O_571,N_14777,N_14780);
or UO_572 (O_572,N_14553,N_14736);
and UO_573 (O_573,N_14583,N_14659);
or UO_574 (O_574,N_14688,N_14660);
or UO_575 (O_575,N_14523,N_14526);
or UO_576 (O_576,N_14694,N_14946);
or UO_577 (O_577,N_14880,N_14847);
nand UO_578 (O_578,N_14716,N_14800);
nor UO_579 (O_579,N_14879,N_14647);
and UO_580 (O_580,N_14799,N_14581);
or UO_581 (O_581,N_14542,N_14884);
or UO_582 (O_582,N_14643,N_14636);
nand UO_583 (O_583,N_14867,N_14658);
nand UO_584 (O_584,N_14802,N_14755);
xor UO_585 (O_585,N_14533,N_14880);
nand UO_586 (O_586,N_14936,N_14699);
and UO_587 (O_587,N_14542,N_14847);
nand UO_588 (O_588,N_14645,N_14810);
nor UO_589 (O_589,N_14658,N_14531);
nand UO_590 (O_590,N_14524,N_14541);
nor UO_591 (O_591,N_14864,N_14579);
and UO_592 (O_592,N_14995,N_14964);
and UO_593 (O_593,N_14793,N_14767);
and UO_594 (O_594,N_14925,N_14514);
or UO_595 (O_595,N_14913,N_14968);
and UO_596 (O_596,N_14585,N_14602);
and UO_597 (O_597,N_14702,N_14717);
or UO_598 (O_598,N_14827,N_14690);
or UO_599 (O_599,N_14952,N_14982);
and UO_600 (O_600,N_14956,N_14819);
and UO_601 (O_601,N_14580,N_14804);
xor UO_602 (O_602,N_14833,N_14513);
nor UO_603 (O_603,N_14995,N_14763);
and UO_604 (O_604,N_14868,N_14687);
nand UO_605 (O_605,N_14594,N_14643);
nand UO_606 (O_606,N_14588,N_14566);
and UO_607 (O_607,N_14826,N_14996);
nor UO_608 (O_608,N_14778,N_14840);
or UO_609 (O_609,N_14934,N_14624);
and UO_610 (O_610,N_14577,N_14980);
nor UO_611 (O_611,N_14908,N_14912);
or UO_612 (O_612,N_14956,N_14820);
xnor UO_613 (O_613,N_14819,N_14794);
nand UO_614 (O_614,N_14758,N_14741);
or UO_615 (O_615,N_14915,N_14995);
nor UO_616 (O_616,N_14739,N_14585);
and UO_617 (O_617,N_14760,N_14951);
nor UO_618 (O_618,N_14935,N_14940);
and UO_619 (O_619,N_14504,N_14822);
or UO_620 (O_620,N_14955,N_14895);
or UO_621 (O_621,N_14605,N_14748);
nand UO_622 (O_622,N_14746,N_14788);
nor UO_623 (O_623,N_14946,N_14722);
or UO_624 (O_624,N_14516,N_14883);
and UO_625 (O_625,N_14788,N_14708);
nand UO_626 (O_626,N_14887,N_14968);
nand UO_627 (O_627,N_14526,N_14764);
and UO_628 (O_628,N_14663,N_14563);
nor UO_629 (O_629,N_14673,N_14749);
nor UO_630 (O_630,N_14592,N_14739);
xnor UO_631 (O_631,N_14619,N_14845);
xnor UO_632 (O_632,N_14562,N_14748);
nand UO_633 (O_633,N_14696,N_14908);
and UO_634 (O_634,N_14727,N_14630);
or UO_635 (O_635,N_14939,N_14920);
or UO_636 (O_636,N_14975,N_14669);
and UO_637 (O_637,N_14770,N_14796);
nand UO_638 (O_638,N_14958,N_14773);
nand UO_639 (O_639,N_14749,N_14641);
xnor UO_640 (O_640,N_14500,N_14545);
nor UO_641 (O_641,N_14594,N_14538);
nor UO_642 (O_642,N_14974,N_14845);
nand UO_643 (O_643,N_14699,N_14737);
nor UO_644 (O_644,N_14887,N_14896);
and UO_645 (O_645,N_14736,N_14729);
or UO_646 (O_646,N_14760,N_14649);
and UO_647 (O_647,N_14937,N_14983);
and UO_648 (O_648,N_14791,N_14503);
nand UO_649 (O_649,N_14637,N_14720);
nor UO_650 (O_650,N_14688,N_14924);
or UO_651 (O_651,N_14633,N_14796);
xnor UO_652 (O_652,N_14605,N_14637);
nor UO_653 (O_653,N_14895,N_14879);
and UO_654 (O_654,N_14816,N_14715);
nor UO_655 (O_655,N_14746,N_14569);
nand UO_656 (O_656,N_14888,N_14592);
xor UO_657 (O_657,N_14604,N_14593);
or UO_658 (O_658,N_14896,N_14578);
nor UO_659 (O_659,N_14856,N_14807);
or UO_660 (O_660,N_14512,N_14635);
and UO_661 (O_661,N_14661,N_14563);
nor UO_662 (O_662,N_14692,N_14532);
and UO_663 (O_663,N_14831,N_14763);
and UO_664 (O_664,N_14948,N_14637);
and UO_665 (O_665,N_14786,N_14721);
xor UO_666 (O_666,N_14768,N_14901);
nand UO_667 (O_667,N_14883,N_14767);
nor UO_668 (O_668,N_14767,N_14694);
or UO_669 (O_669,N_14925,N_14902);
and UO_670 (O_670,N_14765,N_14776);
and UO_671 (O_671,N_14833,N_14662);
and UO_672 (O_672,N_14655,N_14525);
nor UO_673 (O_673,N_14606,N_14748);
and UO_674 (O_674,N_14589,N_14870);
xnor UO_675 (O_675,N_14927,N_14614);
nor UO_676 (O_676,N_14605,N_14811);
nand UO_677 (O_677,N_14549,N_14925);
nor UO_678 (O_678,N_14906,N_14869);
nor UO_679 (O_679,N_14750,N_14547);
and UO_680 (O_680,N_14868,N_14743);
xor UO_681 (O_681,N_14677,N_14931);
nand UO_682 (O_682,N_14982,N_14731);
or UO_683 (O_683,N_14583,N_14822);
nand UO_684 (O_684,N_14916,N_14834);
and UO_685 (O_685,N_14662,N_14932);
nand UO_686 (O_686,N_14917,N_14533);
and UO_687 (O_687,N_14854,N_14516);
and UO_688 (O_688,N_14762,N_14604);
nor UO_689 (O_689,N_14517,N_14846);
and UO_690 (O_690,N_14618,N_14559);
or UO_691 (O_691,N_14536,N_14979);
nor UO_692 (O_692,N_14929,N_14960);
and UO_693 (O_693,N_14698,N_14552);
or UO_694 (O_694,N_14761,N_14599);
nor UO_695 (O_695,N_14916,N_14792);
and UO_696 (O_696,N_14542,N_14632);
nor UO_697 (O_697,N_14551,N_14534);
nor UO_698 (O_698,N_14907,N_14627);
or UO_699 (O_699,N_14728,N_14913);
nand UO_700 (O_700,N_14791,N_14942);
nand UO_701 (O_701,N_14977,N_14910);
nand UO_702 (O_702,N_14648,N_14920);
or UO_703 (O_703,N_14752,N_14776);
and UO_704 (O_704,N_14821,N_14630);
or UO_705 (O_705,N_14675,N_14501);
and UO_706 (O_706,N_14759,N_14853);
and UO_707 (O_707,N_14617,N_14717);
nor UO_708 (O_708,N_14702,N_14730);
nor UO_709 (O_709,N_14636,N_14628);
and UO_710 (O_710,N_14856,N_14667);
xor UO_711 (O_711,N_14757,N_14591);
or UO_712 (O_712,N_14859,N_14596);
and UO_713 (O_713,N_14515,N_14687);
nor UO_714 (O_714,N_14553,N_14986);
nor UO_715 (O_715,N_14707,N_14548);
or UO_716 (O_716,N_14541,N_14849);
nand UO_717 (O_717,N_14961,N_14776);
and UO_718 (O_718,N_14716,N_14583);
or UO_719 (O_719,N_14906,N_14831);
nor UO_720 (O_720,N_14860,N_14974);
and UO_721 (O_721,N_14904,N_14697);
nand UO_722 (O_722,N_14772,N_14697);
or UO_723 (O_723,N_14638,N_14983);
nand UO_724 (O_724,N_14833,N_14726);
nor UO_725 (O_725,N_14968,N_14849);
and UO_726 (O_726,N_14666,N_14528);
and UO_727 (O_727,N_14582,N_14790);
nor UO_728 (O_728,N_14993,N_14756);
nor UO_729 (O_729,N_14523,N_14716);
nor UO_730 (O_730,N_14969,N_14950);
and UO_731 (O_731,N_14570,N_14505);
nor UO_732 (O_732,N_14803,N_14907);
nand UO_733 (O_733,N_14678,N_14598);
or UO_734 (O_734,N_14726,N_14766);
or UO_735 (O_735,N_14750,N_14622);
and UO_736 (O_736,N_14819,N_14864);
nand UO_737 (O_737,N_14911,N_14698);
and UO_738 (O_738,N_14944,N_14972);
or UO_739 (O_739,N_14927,N_14831);
nand UO_740 (O_740,N_14924,N_14806);
or UO_741 (O_741,N_14716,N_14864);
nor UO_742 (O_742,N_14848,N_14797);
nand UO_743 (O_743,N_14857,N_14882);
or UO_744 (O_744,N_14563,N_14735);
or UO_745 (O_745,N_14546,N_14905);
nor UO_746 (O_746,N_14930,N_14665);
or UO_747 (O_747,N_14689,N_14837);
or UO_748 (O_748,N_14634,N_14755);
or UO_749 (O_749,N_14583,N_14710);
and UO_750 (O_750,N_14954,N_14898);
or UO_751 (O_751,N_14764,N_14909);
xor UO_752 (O_752,N_14547,N_14502);
xnor UO_753 (O_753,N_14948,N_14814);
and UO_754 (O_754,N_14740,N_14599);
or UO_755 (O_755,N_14892,N_14666);
and UO_756 (O_756,N_14835,N_14758);
or UO_757 (O_757,N_14734,N_14652);
or UO_758 (O_758,N_14888,N_14928);
xor UO_759 (O_759,N_14902,N_14699);
nand UO_760 (O_760,N_14620,N_14660);
nor UO_761 (O_761,N_14943,N_14635);
nor UO_762 (O_762,N_14614,N_14982);
or UO_763 (O_763,N_14911,N_14808);
xnor UO_764 (O_764,N_14943,N_14707);
and UO_765 (O_765,N_14575,N_14929);
nor UO_766 (O_766,N_14987,N_14543);
xor UO_767 (O_767,N_14583,N_14789);
or UO_768 (O_768,N_14598,N_14751);
nand UO_769 (O_769,N_14737,N_14845);
nand UO_770 (O_770,N_14542,N_14902);
nor UO_771 (O_771,N_14933,N_14551);
nor UO_772 (O_772,N_14827,N_14956);
nor UO_773 (O_773,N_14516,N_14774);
and UO_774 (O_774,N_14972,N_14755);
nand UO_775 (O_775,N_14657,N_14574);
and UO_776 (O_776,N_14759,N_14933);
nor UO_777 (O_777,N_14766,N_14679);
nor UO_778 (O_778,N_14821,N_14961);
nand UO_779 (O_779,N_14918,N_14944);
and UO_780 (O_780,N_14832,N_14514);
xnor UO_781 (O_781,N_14606,N_14647);
nand UO_782 (O_782,N_14864,N_14943);
and UO_783 (O_783,N_14563,N_14612);
or UO_784 (O_784,N_14726,N_14801);
nand UO_785 (O_785,N_14509,N_14855);
nand UO_786 (O_786,N_14820,N_14775);
or UO_787 (O_787,N_14830,N_14780);
nand UO_788 (O_788,N_14946,N_14785);
and UO_789 (O_789,N_14772,N_14947);
nand UO_790 (O_790,N_14996,N_14868);
and UO_791 (O_791,N_14767,N_14789);
and UO_792 (O_792,N_14664,N_14818);
nor UO_793 (O_793,N_14822,N_14687);
or UO_794 (O_794,N_14545,N_14566);
or UO_795 (O_795,N_14840,N_14510);
nor UO_796 (O_796,N_14815,N_14709);
nor UO_797 (O_797,N_14680,N_14793);
nand UO_798 (O_798,N_14936,N_14755);
and UO_799 (O_799,N_14879,N_14852);
nor UO_800 (O_800,N_14980,N_14851);
and UO_801 (O_801,N_14537,N_14610);
or UO_802 (O_802,N_14907,N_14517);
and UO_803 (O_803,N_14704,N_14812);
and UO_804 (O_804,N_14885,N_14762);
xnor UO_805 (O_805,N_14631,N_14721);
xor UO_806 (O_806,N_14810,N_14628);
nand UO_807 (O_807,N_14631,N_14816);
or UO_808 (O_808,N_14879,N_14560);
or UO_809 (O_809,N_14925,N_14999);
and UO_810 (O_810,N_14845,N_14663);
nand UO_811 (O_811,N_14862,N_14573);
xnor UO_812 (O_812,N_14828,N_14592);
nor UO_813 (O_813,N_14708,N_14581);
nor UO_814 (O_814,N_14999,N_14892);
and UO_815 (O_815,N_14509,N_14864);
and UO_816 (O_816,N_14878,N_14846);
xor UO_817 (O_817,N_14771,N_14548);
xnor UO_818 (O_818,N_14780,N_14676);
xnor UO_819 (O_819,N_14759,N_14897);
and UO_820 (O_820,N_14992,N_14646);
or UO_821 (O_821,N_14516,N_14703);
nand UO_822 (O_822,N_14525,N_14868);
nand UO_823 (O_823,N_14967,N_14943);
or UO_824 (O_824,N_14757,N_14785);
and UO_825 (O_825,N_14905,N_14902);
nand UO_826 (O_826,N_14543,N_14909);
xor UO_827 (O_827,N_14800,N_14746);
and UO_828 (O_828,N_14899,N_14594);
nand UO_829 (O_829,N_14679,N_14964);
nor UO_830 (O_830,N_14872,N_14578);
nand UO_831 (O_831,N_14578,N_14899);
nand UO_832 (O_832,N_14706,N_14934);
xor UO_833 (O_833,N_14719,N_14991);
nor UO_834 (O_834,N_14718,N_14743);
nor UO_835 (O_835,N_14500,N_14841);
and UO_836 (O_836,N_14976,N_14657);
and UO_837 (O_837,N_14669,N_14981);
and UO_838 (O_838,N_14909,N_14659);
or UO_839 (O_839,N_14956,N_14949);
nor UO_840 (O_840,N_14721,N_14821);
or UO_841 (O_841,N_14938,N_14891);
or UO_842 (O_842,N_14707,N_14695);
or UO_843 (O_843,N_14649,N_14728);
nand UO_844 (O_844,N_14795,N_14816);
xnor UO_845 (O_845,N_14827,N_14719);
nand UO_846 (O_846,N_14688,N_14501);
and UO_847 (O_847,N_14720,N_14804);
nor UO_848 (O_848,N_14547,N_14976);
xor UO_849 (O_849,N_14639,N_14692);
and UO_850 (O_850,N_14876,N_14745);
or UO_851 (O_851,N_14999,N_14794);
nand UO_852 (O_852,N_14575,N_14940);
or UO_853 (O_853,N_14524,N_14512);
or UO_854 (O_854,N_14818,N_14687);
and UO_855 (O_855,N_14955,N_14920);
or UO_856 (O_856,N_14776,N_14579);
nand UO_857 (O_857,N_14786,N_14579);
nand UO_858 (O_858,N_14760,N_14934);
or UO_859 (O_859,N_14710,N_14875);
nand UO_860 (O_860,N_14780,N_14693);
or UO_861 (O_861,N_14730,N_14910);
xnor UO_862 (O_862,N_14784,N_14663);
and UO_863 (O_863,N_14523,N_14855);
nand UO_864 (O_864,N_14810,N_14610);
nand UO_865 (O_865,N_14894,N_14854);
or UO_866 (O_866,N_14627,N_14577);
and UO_867 (O_867,N_14903,N_14576);
nand UO_868 (O_868,N_14724,N_14854);
nor UO_869 (O_869,N_14556,N_14855);
and UO_870 (O_870,N_14780,N_14840);
xor UO_871 (O_871,N_14925,N_14870);
or UO_872 (O_872,N_14847,N_14884);
and UO_873 (O_873,N_14760,N_14805);
nand UO_874 (O_874,N_14797,N_14640);
xor UO_875 (O_875,N_14624,N_14997);
or UO_876 (O_876,N_14718,N_14641);
or UO_877 (O_877,N_14644,N_14650);
or UO_878 (O_878,N_14741,N_14865);
or UO_879 (O_879,N_14578,N_14813);
or UO_880 (O_880,N_14693,N_14593);
or UO_881 (O_881,N_14999,N_14653);
nor UO_882 (O_882,N_14722,N_14851);
or UO_883 (O_883,N_14977,N_14563);
nor UO_884 (O_884,N_14899,N_14620);
nand UO_885 (O_885,N_14784,N_14862);
or UO_886 (O_886,N_14900,N_14629);
nor UO_887 (O_887,N_14530,N_14930);
and UO_888 (O_888,N_14974,N_14633);
and UO_889 (O_889,N_14812,N_14808);
nor UO_890 (O_890,N_14688,N_14511);
or UO_891 (O_891,N_14700,N_14856);
nand UO_892 (O_892,N_14514,N_14682);
nor UO_893 (O_893,N_14990,N_14852);
or UO_894 (O_894,N_14930,N_14982);
nand UO_895 (O_895,N_14555,N_14846);
nor UO_896 (O_896,N_14969,N_14563);
xnor UO_897 (O_897,N_14989,N_14913);
or UO_898 (O_898,N_14501,N_14803);
xor UO_899 (O_899,N_14598,N_14895);
xnor UO_900 (O_900,N_14758,N_14907);
or UO_901 (O_901,N_14757,N_14822);
nor UO_902 (O_902,N_14681,N_14513);
nor UO_903 (O_903,N_14990,N_14765);
and UO_904 (O_904,N_14536,N_14839);
and UO_905 (O_905,N_14583,N_14623);
nor UO_906 (O_906,N_14966,N_14516);
and UO_907 (O_907,N_14781,N_14507);
nand UO_908 (O_908,N_14954,N_14741);
and UO_909 (O_909,N_14635,N_14781);
nor UO_910 (O_910,N_14587,N_14742);
nand UO_911 (O_911,N_14797,N_14773);
and UO_912 (O_912,N_14578,N_14537);
or UO_913 (O_913,N_14746,N_14859);
and UO_914 (O_914,N_14976,N_14679);
nand UO_915 (O_915,N_14633,N_14940);
xor UO_916 (O_916,N_14798,N_14944);
nand UO_917 (O_917,N_14693,N_14907);
nor UO_918 (O_918,N_14687,N_14971);
or UO_919 (O_919,N_14782,N_14554);
and UO_920 (O_920,N_14662,N_14563);
and UO_921 (O_921,N_14781,N_14628);
and UO_922 (O_922,N_14703,N_14624);
or UO_923 (O_923,N_14670,N_14830);
nor UO_924 (O_924,N_14835,N_14653);
nand UO_925 (O_925,N_14505,N_14925);
nand UO_926 (O_926,N_14567,N_14759);
and UO_927 (O_927,N_14990,N_14653);
or UO_928 (O_928,N_14907,N_14697);
or UO_929 (O_929,N_14698,N_14667);
xor UO_930 (O_930,N_14792,N_14940);
nand UO_931 (O_931,N_14662,N_14877);
or UO_932 (O_932,N_14718,N_14958);
or UO_933 (O_933,N_14628,N_14683);
xor UO_934 (O_934,N_14801,N_14695);
nor UO_935 (O_935,N_14862,N_14680);
nor UO_936 (O_936,N_14799,N_14718);
nand UO_937 (O_937,N_14563,N_14931);
and UO_938 (O_938,N_14931,N_14707);
nor UO_939 (O_939,N_14913,N_14666);
or UO_940 (O_940,N_14596,N_14674);
xor UO_941 (O_941,N_14835,N_14810);
nand UO_942 (O_942,N_14902,N_14733);
nor UO_943 (O_943,N_14680,N_14626);
and UO_944 (O_944,N_14716,N_14843);
and UO_945 (O_945,N_14558,N_14589);
nand UO_946 (O_946,N_14704,N_14862);
nor UO_947 (O_947,N_14514,N_14960);
or UO_948 (O_948,N_14943,N_14548);
xnor UO_949 (O_949,N_14585,N_14923);
xnor UO_950 (O_950,N_14766,N_14671);
nand UO_951 (O_951,N_14564,N_14503);
or UO_952 (O_952,N_14597,N_14999);
xnor UO_953 (O_953,N_14776,N_14755);
or UO_954 (O_954,N_14756,N_14860);
or UO_955 (O_955,N_14785,N_14555);
or UO_956 (O_956,N_14617,N_14975);
nor UO_957 (O_957,N_14588,N_14855);
or UO_958 (O_958,N_14760,N_14691);
nor UO_959 (O_959,N_14846,N_14766);
and UO_960 (O_960,N_14540,N_14795);
nor UO_961 (O_961,N_14717,N_14638);
and UO_962 (O_962,N_14618,N_14866);
nor UO_963 (O_963,N_14808,N_14523);
and UO_964 (O_964,N_14631,N_14995);
and UO_965 (O_965,N_14582,N_14719);
and UO_966 (O_966,N_14599,N_14826);
nand UO_967 (O_967,N_14555,N_14913);
nand UO_968 (O_968,N_14929,N_14534);
or UO_969 (O_969,N_14941,N_14671);
and UO_970 (O_970,N_14785,N_14899);
or UO_971 (O_971,N_14745,N_14512);
or UO_972 (O_972,N_14693,N_14856);
nand UO_973 (O_973,N_14711,N_14718);
or UO_974 (O_974,N_14640,N_14792);
and UO_975 (O_975,N_14759,N_14596);
xnor UO_976 (O_976,N_14836,N_14566);
or UO_977 (O_977,N_14654,N_14949);
nor UO_978 (O_978,N_14814,N_14922);
and UO_979 (O_979,N_14693,N_14832);
nand UO_980 (O_980,N_14970,N_14785);
nor UO_981 (O_981,N_14520,N_14931);
or UO_982 (O_982,N_14710,N_14989);
or UO_983 (O_983,N_14874,N_14605);
nor UO_984 (O_984,N_14783,N_14552);
and UO_985 (O_985,N_14570,N_14643);
and UO_986 (O_986,N_14660,N_14915);
nand UO_987 (O_987,N_14932,N_14881);
or UO_988 (O_988,N_14689,N_14789);
or UO_989 (O_989,N_14713,N_14678);
and UO_990 (O_990,N_14792,N_14649);
nor UO_991 (O_991,N_14922,N_14988);
xor UO_992 (O_992,N_14751,N_14865);
and UO_993 (O_993,N_14588,N_14732);
nand UO_994 (O_994,N_14629,N_14553);
nor UO_995 (O_995,N_14814,N_14549);
nand UO_996 (O_996,N_14556,N_14610);
nand UO_997 (O_997,N_14882,N_14939);
and UO_998 (O_998,N_14567,N_14704);
nand UO_999 (O_999,N_14764,N_14916);
or UO_1000 (O_1000,N_14727,N_14517);
nor UO_1001 (O_1001,N_14530,N_14600);
nor UO_1002 (O_1002,N_14835,N_14692);
or UO_1003 (O_1003,N_14551,N_14927);
or UO_1004 (O_1004,N_14851,N_14895);
or UO_1005 (O_1005,N_14811,N_14869);
nor UO_1006 (O_1006,N_14766,N_14899);
nand UO_1007 (O_1007,N_14733,N_14748);
and UO_1008 (O_1008,N_14581,N_14722);
and UO_1009 (O_1009,N_14781,N_14658);
nor UO_1010 (O_1010,N_14812,N_14724);
and UO_1011 (O_1011,N_14589,N_14819);
and UO_1012 (O_1012,N_14865,N_14851);
nor UO_1013 (O_1013,N_14565,N_14627);
or UO_1014 (O_1014,N_14754,N_14568);
nor UO_1015 (O_1015,N_14637,N_14711);
nand UO_1016 (O_1016,N_14731,N_14583);
nand UO_1017 (O_1017,N_14878,N_14790);
or UO_1018 (O_1018,N_14940,N_14985);
xnor UO_1019 (O_1019,N_14854,N_14519);
nor UO_1020 (O_1020,N_14754,N_14619);
xor UO_1021 (O_1021,N_14848,N_14867);
xnor UO_1022 (O_1022,N_14760,N_14747);
and UO_1023 (O_1023,N_14774,N_14757);
and UO_1024 (O_1024,N_14504,N_14962);
nor UO_1025 (O_1025,N_14795,N_14681);
nand UO_1026 (O_1026,N_14886,N_14548);
nor UO_1027 (O_1027,N_14838,N_14692);
nand UO_1028 (O_1028,N_14946,N_14953);
nand UO_1029 (O_1029,N_14595,N_14931);
or UO_1030 (O_1030,N_14617,N_14875);
xor UO_1031 (O_1031,N_14892,N_14639);
nor UO_1032 (O_1032,N_14639,N_14759);
or UO_1033 (O_1033,N_14849,N_14621);
nor UO_1034 (O_1034,N_14655,N_14710);
or UO_1035 (O_1035,N_14629,N_14961);
nor UO_1036 (O_1036,N_14853,N_14637);
nor UO_1037 (O_1037,N_14603,N_14821);
or UO_1038 (O_1038,N_14542,N_14524);
xor UO_1039 (O_1039,N_14769,N_14920);
or UO_1040 (O_1040,N_14721,N_14805);
and UO_1041 (O_1041,N_14952,N_14885);
nand UO_1042 (O_1042,N_14504,N_14634);
or UO_1043 (O_1043,N_14578,N_14737);
xnor UO_1044 (O_1044,N_14672,N_14681);
nand UO_1045 (O_1045,N_14642,N_14887);
nand UO_1046 (O_1046,N_14570,N_14865);
nand UO_1047 (O_1047,N_14922,N_14625);
or UO_1048 (O_1048,N_14727,N_14515);
nor UO_1049 (O_1049,N_14938,N_14840);
nand UO_1050 (O_1050,N_14935,N_14938);
nor UO_1051 (O_1051,N_14508,N_14693);
and UO_1052 (O_1052,N_14650,N_14988);
or UO_1053 (O_1053,N_14515,N_14679);
or UO_1054 (O_1054,N_14663,N_14634);
and UO_1055 (O_1055,N_14879,N_14671);
or UO_1056 (O_1056,N_14797,N_14676);
nor UO_1057 (O_1057,N_14647,N_14620);
nor UO_1058 (O_1058,N_14635,N_14875);
and UO_1059 (O_1059,N_14750,N_14726);
xnor UO_1060 (O_1060,N_14865,N_14630);
or UO_1061 (O_1061,N_14591,N_14561);
nand UO_1062 (O_1062,N_14976,N_14500);
nand UO_1063 (O_1063,N_14686,N_14874);
xor UO_1064 (O_1064,N_14687,N_14536);
or UO_1065 (O_1065,N_14758,N_14639);
and UO_1066 (O_1066,N_14680,N_14519);
nand UO_1067 (O_1067,N_14690,N_14587);
nand UO_1068 (O_1068,N_14957,N_14743);
nand UO_1069 (O_1069,N_14526,N_14591);
xnor UO_1070 (O_1070,N_14565,N_14724);
and UO_1071 (O_1071,N_14535,N_14859);
nand UO_1072 (O_1072,N_14613,N_14740);
and UO_1073 (O_1073,N_14834,N_14812);
xor UO_1074 (O_1074,N_14695,N_14511);
nor UO_1075 (O_1075,N_14909,N_14915);
nand UO_1076 (O_1076,N_14777,N_14723);
nand UO_1077 (O_1077,N_14954,N_14653);
and UO_1078 (O_1078,N_14953,N_14662);
or UO_1079 (O_1079,N_14573,N_14655);
nor UO_1080 (O_1080,N_14966,N_14809);
or UO_1081 (O_1081,N_14731,N_14944);
and UO_1082 (O_1082,N_14698,N_14749);
or UO_1083 (O_1083,N_14741,N_14689);
nor UO_1084 (O_1084,N_14979,N_14801);
nor UO_1085 (O_1085,N_14995,N_14730);
or UO_1086 (O_1086,N_14965,N_14845);
nor UO_1087 (O_1087,N_14639,N_14912);
xor UO_1088 (O_1088,N_14866,N_14737);
nor UO_1089 (O_1089,N_14762,N_14869);
nand UO_1090 (O_1090,N_14913,N_14824);
or UO_1091 (O_1091,N_14883,N_14722);
or UO_1092 (O_1092,N_14887,N_14706);
nand UO_1093 (O_1093,N_14750,N_14863);
nor UO_1094 (O_1094,N_14568,N_14978);
nor UO_1095 (O_1095,N_14632,N_14930);
nand UO_1096 (O_1096,N_14963,N_14985);
xor UO_1097 (O_1097,N_14785,N_14858);
nand UO_1098 (O_1098,N_14561,N_14687);
nand UO_1099 (O_1099,N_14966,N_14609);
and UO_1100 (O_1100,N_14542,N_14782);
or UO_1101 (O_1101,N_14999,N_14507);
or UO_1102 (O_1102,N_14884,N_14938);
nor UO_1103 (O_1103,N_14962,N_14538);
and UO_1104 (O_1104,N_14588,N_14528);
nand UO_1105 (O_1105,N_14675,N_14722);
or UO_1106 (O_1106,N_14808,N_14655);
nand UO_1107 (O_1107,N_14647,N_14605);
or UO_1108 (O_1108,N_14546,N_14589);
and UO_1109 (O_1109,N_14752,N_14833);
nor UO_1110 (O_1110,N_14969,N_14976);
nor UO_1111 (O_1111,N_14530,N_14963);
and UO_1112 (O_1112,N_14643,N_14926);
or UO_1113 (O_1113,N_14913,N_14724);
or UO_1114 (O_1114,N_14846,N_14508);
and UO_1115 (O_1115,N_14973,N_14806);
or UO_1116 (O_1116,N_14695,N_14976);
nand UO_1117 (O_1117,N_14536,N_14632);
nor UO_1118 (O_1118,N_14678,N_14860);
and UO_1119 (O_1119,N_14725,N_14699);
nand UO_1120 (O_1120,N_14890,N_14921);
or UO_1121 (O_1121,N_14514,N_14623);
and UO_1122 (O_1122,N_14738,N_14536);
xnor UO_1123 (O_1123,N_14749,N_14782);
and UO_1124 (O_1124,N_14966,N_14756);
nor UO_1125 (O_1125,N_14857,N_14993);
or UO_1126 (O_1126,N_14501,N_14807);
and UO_1127 (O_1127,N_14973,N_14629);
xor UO_1128 (O_1128,N_14569,N_14720);
or UO_1129 (O_1129,N_14629,N_14948);
nand UO_1130 (O_1130,N_14972,N_14750);
nand UO_1131 (O_1131,N_14910,N_14584);
or UO_1132 (O_1132,N_14903,N_14861);
xnor UO_1133 (O_1133,N_14702,N_14923);
and UO_1134 (O_1134,N_14649,N_14564);
nor UO_1135 (O_1135,N_14561,N_14670);
nor UO_1136 (O_1136,N_14951,N_14810);
or UO_1137 (O_1137,N_14832,N_14697);
nor UO_1138 (O_1138,N_14732,N_14525);
or UO_1139 (O_1139,N_14792,N_14897);
or UO_1140 (O_1140,N_14621,N_14691);
nor UO_1141 (O_1141,N_14787,N_14625);
nor UO_1142 (O_1142,N_14708,N_14677);
and UO_1143 (O_1143,N_14697,N_14548);
nor UO_1144 (O_1144,N_14803,N_14933);
nor UO_1145 (O_1145,N_14681,N_14917);
and UO_1146 (O_1146,N_14605,N_14643);
or UO_1147 (O_1147,N_14931,N_14995);
nor UO_1148 (O_1148,N_14909,N_14743);
nor UO_1149 (O_1149,N_14866,N_14612);
and UO_1150 (O_1150,N_14668,N_14745);
xor UO_1151 (O_1151,N_14564,N_14604);
nor UO_1152 (O_1152,N_14592,N_14624);
nor UO_1153 (O_1153,N_14758,N_14746);
and UO_1154 (O_1154,N_14778,N_14766);
and UO_1155 (O_1155,N_14502,N_14993);
or UO_1156 (O_1156,N_14997,N_14659);
and UO_1157 (O_1157,N_14632,N_14985);
nor UO_1158 (O_1158,N_14630,N_14664);
or UO_1159 (O_1159,N_14702,N_14888);
xnor UO_1160 (O_1160,N_14895,N_14700);
or UO_1161 (O_1161,N_14821,N_14507);
nand UO_1162 (O_1162,N_14729,N_14527);
nand UO_1163 (O_1163,N_14930,N_14701);
nand UO_1164 (O_1164,N_14733,N_14895);
nor UO_1165 (O_1165,N_14552,N_14702);
or UO_1166 (O_1166,N_14557,N_14561);
nand UO_1167 (O_1167,N_14579,N_14521);
nor UO_1168 (O_1168,N_14507,N_14977);
nand UO_1169 (O_1169,N_14609,N_14515);
nand UO_1170 (O_1170,N_14771,N_14857);
nor UO_1171 (O_1171,N_14793,N_14715);
and UO_1172 (O_1172,N_14953,N_14600);
and UO_1173 (O_1173,N_14951,N_14948);
and UO_1174 (O_1174,N_14769,N_14818);
nand UO_1175 (O_1175,N_14942,N_14890);
or UO_1176 (O_1176,N_14500,N_14640);
nand UO_1177 (O_1177,N_14852,N_14928);
and UO_1178 (O_1178,N_14579,N_14565);
nor UO_1179 (O_1179,N_14648,N_14969);
nor UO_1180 (O_1180,N_14745,N_14529);
nor UO_1181 (O_1181,N_14912,N_14837);
nand UO_1182 (O_1182,N_14897,N_14545);
or UO_1183 (O_1183,N_14784,N_14506);
nor UO_1184 (O_1184,N_14896,N_14958);
or UO_1185 (O_1185,N_14825,N_14668);
nor UO_1186 (O_1186,N_14854,N_14627);
and UO_1187 (O_1187,N_14897,N_14901);
nor UO_1188 (O_1188,N_14721,N_14987);
or UO_1189 (O_1189,N_14504,N_14523);
and UO_1190 (O_1190,N_14929,N_14582);
or UO_1191 (O_1191,N_14805,N_14915);
or UO_1192 (O_1192,N_14642,N_14639);
nor UO_1193 (O_1193,N_14547,N_14862);
nor UO_1194 (O_1194,N_14831,N_14861);
nand UO_1195 (O_1195,N_14781,N_14669);
or UO_1196 (O_1196,N_14602,N_14522);
nand UO_1197 (O_1197,N_14917,N_14595);
or UO_1198 (O_1198,N_14898,N_14863);
nand UO_1199 (O_1199,N_14788,N_14949);
or UO_1200 (O_1200,N_14826,N_14676);
and UO_1201 (O_1201,N_14930,N_14710);
and UO_1202 (O_1202,N_14919,N_14908);
nor UO_1203 (O_1203,N_14839,N_14738);
or UO_1204 (O_1204,N_14665,N_14709);
and UO_1205 (O_1205,N_14715,N_14604);
and UO_1206 (O_1206,N_14920,N_14935);
nor UO_1207 (O_1207,N_14987,N_14599);
nor UO_1208 (O_1208,N_14978,N_14610);
xnor UO_1209 (O_1209,N_14790,N_14557);
nand UO_1210 (O_1210,N_14841,N_14569);
or UO_1211 (O_1211,N_14507,N_14568);
nor UO_1212 (O_1212,N_14571,N_14938);
or UO_1213 (O_1213,N_14998,N_14889);
or UO_1214 (O_1214,N_14549,N_14684);
and UO_1215 (O_1215,N_14942,N_14608);
nand UO_1216 (O_1216,N_14765,N_14913);
or UO_1217 (O_1217,N_14647,N_14974);
or UO_1218 (O_1218,N_14653,N_14650);
nor UO_1219 (O_1219,N_14784,N_14949);
and UO_1220 (O_1220,N_14575,N_14758);
nand UO_1221 (O_1221,N_14529,N_14941);
nand UO_1222 (O_1222,N_14747,N_14581);
and UO_1223 (O_1223,N_14957,N_14569);
and UO_1224 (O_1224,N_14761,N_14726);
or UO_1225 (O_1225,N_14871,N_14530);
or UO_1226 (O_1226,N_14996,N_14734);
nor UO_1227 (O_1227,N_14895,N_14981);
and UO_1228 (O_1228,N_14822,N_14740);
nand UO_1229 (O_1229,N_14501,N_14929);
nor UO_1230 (O_1230,N_14698,N_14633);
nand UO_1231 (O_1231,N_14808,N_14698);
or UO_1232 (O_1232,N_14958,N_14780);
and UO_1233 (O_1233,N_14960,N_14699);
nor UO_1234 (O_1234,N_14765,N_14815);
or UO_1235 (O_1235,N_14869,N_14910);
nand UO_1236 (O_1236,N_14732,N_14654);
xnor UO_1237 (O_1237,N_14955,N_14705);
or UO_1238 (O_1238,N_14756,N_14954);
nand UO_1239 (O_1239,N_14812,N_14516);
xor UO_1240 (O_1240,N_14709,N_14985);
and UO_1241 (O_1241,N_14819,N_14787);
nor UO_1242 (O_1242,N_14580,N_14799);
or UO_1243 (O_1243,N_14799,N_14986);
or UO_1244 (O_1244,N_14971,N_14937);
or UO_1245 (O_1245,N_14943,N_14969);
or UO_1246 (O_1246,N_14611,N_14715);
and UO_1247 (O_1247,N_14653,N_14839);
or UO_1248 (O_1248,N_14706,N_14777);
xor UO_1249 (O_1249,N_14844,N_14645);
nor UO_1250 (O_1250,N_14932,N_14842);
xor UO_1251 (O_1251,N_14964,N_14557);
nand UO_1252 (O_1252,N_14614,N_14676);
nand UO_1253 (O_1253,N_14707,N_14582);
nor UO_1254 (O_1254,N_14984,N_14961);
nor UO_1255 (O_1255,N_14883,N_14622);
nand UO_1256 (O_1256,N_14560,N_14946);
and UO_1257 (O_1257,N_14522,N_14841);
nor UO_1258 (O_1258,N_14619,N_14882);
nand UO_1259 (O_1259,N_14669,N_14794);
nand UO_1260 (O_1260,N_14851,N_14967);
nand UO_1261 (O_1261,N_14503,N_14627);
nand UO_1262 (O_1262,N_14915,N_14793);
xnor UO_1263 (O_1263,N_14951,N_14507);
nor UO_1264 (O_1264,N_14882,N_14973);
or UO_1265 (O_1265,N_14925,N_14617);
nor UO_1266 (O_1266,N_14579,N_14811);
and UO_1267 (O_1267,N_14968,N_14762);
nand UO_1268 (O_1268,N_14769,N_14500);
and UO_1269 (O_1269,N_14538,N_14701);
and UO_1270 (O_1270,N_14671,N_14912);
nor UO_1271 (O_1271,N_14684,N_14898);
nand UO_1272 (O_1272,N_14565,N_14962);
nand UO_1273 (O_1273,N_14836,N_14995);
or UO_1274 (O_1274,N_14696,N_14953);
nor UO_1275 (O_1275,N_14840,N_14757);
or UO_1276 (O_1276,N_14859,N_14732);
or UO_1277 (O_1277,N_14924,N_14512);
and UO_1278 (O_1278,N_14518,N_14818);
nand UO_1279 (O_1279,N_14786,N_14964);
nand UO_1280 (O_1280,N_14627,N_14530);
or UO_1281 (O_1281,N_14943,N_14523);
and UO_1282 (O_1282,N_14890,N_14926);
or UO_1283 (O_1283,N_14746,N_14879);
or UO_1284 (O_1284,N_14795,N_14731);
and UO_1285 (O_1285,N_14948,N_14706);
nand UO_1286 (O_1286,N_14963,N_14882);
and UO_1287 (O_1287,N_14604,N_14768);
nand UO_1288 (O_1288,N_14965,N_14804);
and UO_1289 (O_1289,N_14762,N_14682);
nor UO_1290 (O_1290,N_14640,N_14882);
and UO_1291 (O_1291,N_14698,N_14619);
and UO_1292 (O_1292,N_14606,N_14763);
nor UO_1293 (O_1293,N_14691,N_14698);
nand UO_1294 (O_1294,N_14982,N_14645);
nor UO_1295 (O_1295,N_14522,N_14843);
nand UO_1296 (O_1296,N_14801,N_14898);
nand UO_1297 (O_1297,N_14557,N_14862);
nor UO_1298 (O_1298,N_14846,N_14785);
or UO_1299 (O_1299,N_14982,N_14672);
or UO_1300 (O_1300,N_14567,N_14927);
nor UO_1301 (O_1301,N_14685,N_14800);
nand UO_1302 (O_1302,N_14903,N_14620);
xor UO_1303 (O_1303,N_14613,N_14955);
nand UO_1304 (O_1304,N_14509,N_14592);
xor UO_1305 (O_1305,N_14718,N_14746);
nor UO_1306 (O_1306,N_14867,N_14712);
nand UO_1307 (O_1307,N_14731,N_14542);
xnor UO_1308 (O_1308,N_14880,N_14928);
or UO_1309 (O_1309,N_14905,N_14811);
nor UO_1310 (O_1310,N_14941,N_14909);
nor UO_1311 (O_1311,N_14912,N_14508);
nor UO_1312 (O_1312,N_14786,N_14627);
nand UO_1313 (O_1313,N_14823,N_14995);
xnor UO_1314 (O_1314,N_14542,N_14895);
nand UO_1315 (O_1315,N_14992,N_14764);
nand UO_1316 (O_1316,N_14611,N_14921);
xor UO_1317 (O_1317,N_14638,N_14813);
nand UO_1318 (O_1318,N_14791,N_14991);
and UO_1319 (O_1319,N_14884,N_14914);
and UO_1320 (O_1320,N_14694,N_14914);
nand UO_1321 (O_1321,N_14722,N_14842);
or UO_1322 (O_1322,N_14754,N_14766);
and UO_1323 (O_1323,N_14808,N_14888);
and UO_1324 (O_1324,N_14843,N_14760);
nor UO_1325 (O_1325,N_14783,N_14602);
nor UO_1326 (O_1326,N_14688,N_14763);
nor UO_1327 (O_1327,N_14702,N_14654);
and UO_1328 (O_1328,N_14626,N_14856);
or UO_1329 (O_1329,N_14678,N_14882);
and UO_1330 (O_1330,N_14705,N_14811);
and UO_1331 (O_1331,N_14919,N_14730);
nor UO_1332 (O_1332,N_14728,N_14742);
nor UO_1333 (O_1333,N_14882,N_14673);
nand UO_1334 (O_1334,N_14656,N_14770);
nand UO_1335 (O_1335,N_14987,N_14806);
nand UO_1336 (O_1336,N_14503,N_14710);
or UO_1337 (O_1337,N_14886,N_14809);
nand UO_1338 (O_1338,N_14720,N_14793);
nand UO_1339 (O_1339,N_14506,N_14665);
nand UO_1340 (O_1340,N_14501,N_14747);
or UO_1341 (O_1341,N_14521,N_14509);
nor UO_1342 (O_1342,N_14844,N_14840);
nand UO_1343 (O_1343,N_14865,N_14984);
nor UO_1344 (O_1344,N_14980,N_14691);
and UO_1345 (O_1345,N_14693,N_14798);
nand UO_1346 (O_1346,N_14962,N_14532);
and UO_1347 (O_1347,N_14575,N_14982);
nor UO_1348 (O_1348,N_14640,N_14903);
xor UO_1349 (O_1349,N_14642,N_14732);
nor UO_1350 (O_1350,N_14603,N_14544);
or UO_1351 (O_1351,N_14971,N_14761);
nand UO_1352 (O_1352,N_14770,N_14502);
xor UO_1353 (O_1353,N_14998,N_14739);
or UO_1354 (O_1354,N_14714,N_14993);
or UO_1355 (O_1355,N_14659,N_14546);
and UO_1356 (O_1356,N_14990,N_14866);
nand UO_1357 (O_1357,N_14962,N_14632);
nand UO_1358 (O_1358,N_14622,N_14509);
xnor UO_1359 (O_1359,N_14829,N_14518);
or UO_1360 (O_1360,N_14699,N_14516);
nor UO_1361 (O_1361,N_14973,N_14641);
nor UO_1362 (O_1362,N_14733,N_14874);
nor UO_1363 (O_1363,N_14778,N_14568);
nor UO_1364 (O_1364,N_14705,N_14831);
and UO_1365 (O_1365,N_14743,N_14926);
nor UO_1366 (O_1366,N_14552,N_14944);
nor UO_1367 (O_1367,N_14669,N_14510);
nor UO_1368 (O_1368,N_14907,N_14715);
nand UO_1369 (O_1369,N_14870,N_14640);
nor UO_1370 (O_1370,N_14782,N_14887);
and UO_1371 (O_1371,N_14603,N_14956);
nand UO_1372 (O_1372,N_14940,N_14624);
and UO_1373 (O_1373,N_14815,N_14955);
nand UO_1374 (O_1374,N_14860,N_14608);
and UO_1375 (O_1375,N_14972,N_14725);
nand UO_1376 (O_1376,N_14645,N_14552);
nor UO_1377 (O_1377,N_14629,N_14872);
nor UO_1378 (O_1378,N_14723,N_14561);
and UO_1379 (O_1379,N_14642,N_14934);
and UO_1380 (O_1380,N_14651,N_14692);
nor UO_1381 (O_1381,N_14807,N_14664);
nand UO_1382 (O_1382,N_14557,N_14703);
nor UO_1383 (O_1383,N_14619,N_14824);
nand UO_1384 (O_1384,N_14989,N_14702);
xor UO_1385 (O_1385,N_14565,N_14945);
nand UO_1386 (O_1386,N_14909,N_14577);
nand UO_1387 (O_1387,N_14879,N_14820);
or UO_1388 (O_1388,N_14502,N_14787);
nand UO_1389 (O_1389,N_14857,N_14536);
or UO_1390 (O_1390,N_14936,N_14786);
and UO_1391 (O_1391,N_14882,N_14848);
nand UO_1392 (O_1392,N_14507,N_14557);
nand UO_1393 (O_1393,N_14505,N_14803);
nand UO_1394 (O_1394,N_14778,N_14755);
nand UO_1395 (O_1395,N_14859,N_14688);
and UO_1396 (O_1396,N_14709,N_14962);
or UO_1397 (O_1397,N_14716,N_14598);
xnor UO_1398 (O_1398,N_14803,N_14796);
nor UO_1399 (O_1399,N_14689,N_14769);
nand UO_1400 (O_1400,N_14892,N_14928);
nor UO_1401 (O_1401,N_14952,N_14699);
or UO_1402 (O_1402,N_14536,N_14811);
or UO_1403 (O_1403,N_14926,N_14784);
nor UO_1404 (O_1404,N_14897,N_14976);
nor UO_1405 (O_1405,N_14503,N_14855);
and UO_1406 (O_1406,N_14957,N_14962);
or UO_1407 (O_1407,N_14752,N_14569);
and UO_1408 (O_1408,N_14775,N_14964);
or UO_1409 (O_1409,N_14610,N_14689);
nand UO_1410 (O_1410,N_14592,N_14951);
or UO_1411 (O_1411,N_14667,N_14934);
or UO_1412 (O_1412,N_14572,N_14610);
xor UO_1413 (O_1413,N_14746,N_14728);
nor UO_1414 (O_1414,N_14903,N_14799);
nand UO_1415 (O_1415,N_14849,N_14612);
and UO_1416 (O_1416,N_14762,N_14708);
xor UO_1417 (O_1417,N_14742,N_14835);
and UO_1418 (O_1418,N_14928,N_14514);
and UO_1419 (O_1419,N_14704,N_14896);
nor UO_1420 (O_1420,N_14819,N_14911);
and UO_1421 (O_1421,N_14992,N_14511);
nand UO_1422 (O_1422,N_14699,N_14851);
and UO_1423 (O_1423,N_14712,N_14723);
nor UO_1424 (O_1424,N_14923,N_14980);
and UO_1425 (O_1425,N_14520,N_14993);
nor UO_1426 (O_1426,N_14771,N_14883);
or UO_1427 (O_1427,N_14830,N_14520);
nand UO_1428 (O_1428,N_14970,N_14795);
nor UO_1429 (O_1429,N_14961,N_14922);
or UO_1430 (O_1430,N_14575,N_14896);
nor UO_1431 (O_1431,N_14554,N_14589);
and UO_1432 (O_1432,N_14588,N_14819);
or UO_1433 (O_1433,N_14976,N_14520);
and UO_1434 (O_1434,N_14619,N_14684);
and UO_1435 (O_1435,N_14823,N_14668);
nand UO_1436 (O_1436,N_14635,N_14627);
nor UO_1437 (O_1437,N_14576,N_14710);
nand UO_1438 (O_1438,N_14760,N_14821);
nor UO_1439 (O_1439,N_14508,N_14756);
nand UO_1440 (O_1440,N_14556,N_14700);
and UO_1441 (O_1441,N_14725,N_14802);
xnor UO_1442 (O_1442,N_14827,N_14553);
or UO_1443 (O_1443,N_14758,N_14875);
or UO_1444 (O_1444,N_14745,N_14697);
nand UO_1445 (O_1445,N_14815,N_14810);
nand UO_1446 (O_1446,N_14532,N_14871);
nand UO_1447 (O_1447,N_14992,N_14996);
and UO_1448 (O_1448,N_14912,N_14727);
and UO_1449 (O_1449,N_14513,N_14530);
and UO_1450 (O_1450,N_14680,N_14792);
and UO_1451 (O_1451,N_14901,N_14823);
nand UO_1452 (O_1452,N_14978,N_14776);
nand UO_1453 (O_1453,N_14881,N_14656);
nand UO_1454 (O_1454,N_14877,N_14981);
nor UO_1455 (O_1455,N_14933,N_14672);
nor UO_1456 (O_1456,N_14841,N_14556);
xor UO_1457 (O_1457,N_14721,N_14664);
nor UO_1458 (O_1458,N_14716,N_14954);
nand UO_1459 (O_1459,N_14963,N_14923);
nor UO_1460 (O_1460,N_14842,N_14817);
or UO_1461 (O_1461,N_14794,N_14977);
or UO_1462 (O_1462,N_14602,N_14687);
and UO_1463 (O_1463,N_14809,N_14955);
or UO_1464 (O_1464,N_14860,N_14932);
nor UO_1465 (O_1465,N_14615,N_14868);
or UO_1466 (O_1466,N_14752,N_14773);
nand UO_1467 (O_1467,N_14974,N_14545);
nor UO_1468 (O_1468,N_14584,N_14571);
nor UO_1469 (O_1469,N_14818,N_14633);
nand UO_1470 (O_1470,N_14642,N_14967);
nand UO_1471 (O_1471,N_14907,N_14799);
xor UO_1472 (O_1472,N_14611,N_14925);
nor UO_1473 (O_1473,N_14729,N_14642);
or UO_1474 (O_1474,N_14884,N_14784);
nand UO_1475 (O_1475,N_14607,N_14698);
or UO_1476 (O_1476,N_14790,N_14543);
or UO_1477 (O_1477,N_14680,N_14617);
xnor UO_1478 (O_1478,N_14933,N_14609);
xor UO_1479 (O_1479,N_14607,N_14672);
or UO_1480 (O_1480,N_14787,N_14721);
nor UO_1481 (O_1481,N_14658,N_14588);
xnor UO_1482 (O_1482,N_14697,N_14669);
nor UO_1483 (O_1483,N_14617,N_14850);
nor UO_1484 (O_1484,N_14868,N_14852);
and UO_1485 (O_1485,N_14772,N_14521);
and UO_1486 (O_1486,N_14630,N_14540);
nand UO_1487 (O_1487,N_14829,N_14842);
and UO_1488 (O_1488,N_14750,N_14925);
or UO_1489 (O_1489,N_14656,N_14810);
xnor UO_1490 (O_1490,N_14918,N_14599);
or UO_1491 (O_1491,N_14612,N_14906);
nand UO_1492 (O_1492,N_14501,N_14601);
and UO_1493 (O_1493,N_14742,N_14722);
or UO_1494 (O_1494,N_14561,N_14790);
xor UO_1495 (O_1495,N_14985,N_14682);
and UO_1496 (O_1496,N_14834,N_14748);
and UO_1497 (O_1497,N_14930,N_14671);
or UO_1498 (O_1498,N_14768,N_14652);
and UO_1499 (O_1499,N_14887,N_14839);
or UO_1500 (O_1500,N_14583,N_14597);
or UO_1501 (O_1501,N_14582,N_14523);
nor UO_1502 (O_1502,N_14867,N_14956);
nor UO_1503 (O_1503,N_14919,N_14528);
or UO_1504 (O_1504,N_14963,N_14504);
and UO_1505 (O_1505,N_14762,N_14871);
xnor UO_1506 (O_1506,N_14648,N_14874);
or UO_1507 (O_1507,N_14687,N_14856);
and UO_1508 (O_1508,N_14616,N_14559);
nor UO_1509 (O_1509,N_14627,N_14975);
and UO_1510 (O_1510,N_14668,N_14888);
and UO_1511 (O_1511,N_14977,N_14540);
nor UO_1512 (O_1512,N_14890,N_14512);
nor UO_1513 (O_1513,N_14996,N_14520);
nor UO_1514 (O_1514,N_14994,N_14548);
nand UO_1515 (O_1515,N_14987,N_14896);
xor UO_1516 (O_1516,N_14607,N_14688);
or UO_1517 (O_1517,N_14836,N_14867);
nand UO_1518 (O_1518,N_14966,N_14543);
and UO_1519 (O_1519,N_14992,N_14853);
nor UO_1520 (O_1520,N_14619,N_14785);
or UO_1521 (O_1521,N_14968,N_14590);
nand UO_1522 (O_1522,N_14573,N_14672);
nor UO_1523 (O_1523,N_14661,N_14729);
or UO_1524 (O_1524,N_14792,N_14779);
or UO_1525 (O_1525,N_14704,N_14860);
nor UO_1526 (O_1526,N_14696,N_14512);
nor UO_1527 (O_1527,N_14535,N_14734);
and UO_1528 (O_1528,N_14978,N_14987);
or UO_1529 (O_1529,N_14791,N_14643);
nor UO_1530 (O_1530,N_14881,N_14675);
nand UO_1531 (O_1531,N_14888,N_14935);
and UO_1532 (O_1532,N_14579,N_14984);
or UO_1533 (O_1533,N_14660,N_14686);
nor UO_1534 (O_1534,N_14915,N_14634);
nand UO_1535 (O_1535,N_14742,N_14767);
nand UO_1536 (O_1536,N_14811,N_14593);
nand UO_1537 (O_1537,N_14826,N_14750);
xnor UO_1538 (O_1538,N_14504,N_14847);
nand UO_1539 (O_1539,N_14820,N_14510);
and UO_1540 (O_1540,N_14590,N_14771);
or UO_1541 (O_1541,N_14592,N_14563);
nand UO_1542 (O_1542,N_14953,N_14781);
nand UO_1543 (O_1543,N_14699,N_14951);
nand UO_1544 (O_1544,N_14655,N_14700);
nand UO_1545 (O_1545,N_14515,N_14857);
nand UO_1546 (O_1546,N_14624,N_14974);
or UO_1547 (O_1547,N_14691,N_14823);
and UO_1548 (O_1548,N_14964,N_14898);
nor UO_1549 (O_1549,N_14869,N_14943);
nand UO_1550 (O_1550,N_14670,N_14671);
nand UO_1551 (O_1551,N_14508,N_14958);
nor UO_1552 (O_1552,N_14942,N_14881);
and UO_1553 (O_1553,N_14933,N_14522);
and UO_1554 (O_1554,N_14860,N_14854);
xor UO_1555 (O_1555,N_14901,N_14892);
nor UO_1556 (O_1556,N_14604,N_14618);
and UO_1557 (O_1557,N_14512,N_14766);
and UO_1558 (O_1558,N_14567,N_14583);
nor UO_1559 (O_1559,N_14778,N_14583);
or UO_1560 (O_1560,N_14791,N_14770);
nor UO_1561 (O_1561,N_14998,N_14787);
nand UO_1562 (O_1562,N_14551,N_14567);
or UO_1563 (O_1563,N_14894,N_14619);
nand UO_1564 (O_1564,N_14826,N_14594);
and UO_1565 (O_1565,N_14548,N_14564);
or UO_1566 (O_1566,N_14852,N_14823);
or UO_1567 (O_1567,N_14771,N_14703);
and UO_1568 (O_1568,N_14575,N_14803);
and UO_1569 (O_1569,N_14642,N_14726);
nor UO_1570 (O_1570,N_14933,N_14569);
nor UO_1571 (O_1571,N_14650,N_14589);
nor UO_1572 (O_1572,N_14538,N_14838);
nor UO_1573 (O_1573,N_14541,N_14940);
and UO_1574 (O_1574,N_14644,N_14720);
or UO_1575 (O_1575,N_14655,N_14760);
and UO_1576 (O_1576,N_14972,N_14674);
or UO_1577 (O_1577,N_14931,N_14600);
nor UO_1578 (O_1578,N_14568,N_14516);
or UO_1579 (O_1579,N_14700,N_14710);
and UO_1580 (O_1580,N_14567,N_14975);
nor UO_1581 (O_1581,N_14854,N_14746);
xor UO_1582 (O_1582,N_14623,N_14730);
nand UO_1583 (O_1583,N_14947,N_14889);
and UO_1584 (O_1584,N_14934,N_14767);
and UO_1585 (O_1585,N_14748,N_14663);
and UO_1586 (O_1586,N_14835,N_14878);
nor UO_1587 (O_1587,N_14853,N_14520);
xor UO_1588 (O_1588,N_14977,N_14824);
or UO_1589 (O_1589,N_14886,N_14989);
nor UO_1590 (O_1590,N_14859,N_14925);
or UO_1591 (O_1591,N_14946,N_14797);
or UO_1592 (O_1592,N_14633,N_14989);
or UO_1593 (O_1593,N_14752,N_14620);
and UO_1594 (O_1594,N_14643,N_14769);
or UO_1595 (O_1595,N_14628,N_14700);
and UO_1596 (O_1596,N_14510,N_14796);
or UO_1597 (O_1597,N_14852,N_14791);
or UO_1598 (O_1598,N_14623,N_14770);
nand UO_1599 (O_1599,N_14684,N_14666);
or UO_1600 (O_1600,N_14944,N_14750);
or UO_1601 (O_1601,N_14889,N_14609);
nor UO_1602 (O_1602,N_14812,N_14531);
or UO_1603 (O_1603,N_14742,N_14674);
or UO_1604 (O_1604,N_14592,N_14789);
nand UO_1605 (O_1605,N_14622,N_14672);
and UO_1606 (O_1606,N_14841,N_14876);
xnor UO_1607 (O_1607,N_14773,N_14894);
nor UO_1608 (O_1608,N_14865,N_14660);
nand UO_1609 (O_1609,N_14758,N_14888);
nand UO_1610 (O_1610,N_14814,N_14808);
nand UO_1611 (O_1611,N_14676,N_14791);
nand UO_1612 (O_1612,N_14949,N_14538);
nand UO_1613 (O_1613,N_14812,N_14535);
xnor UO_1614 (O_1614,N_14711,N_14884);
nand UO_1615 (O_1615,N_14704,N_14717);
nand UO_1616 (O_1616,N_14855,N_14552);
and UO_1617 (O_1617,N_14883,N_14577);
nor UO_1618 (O_1618,N_14840,N_14560);
nor UO_1619 (O_1619,N_14594,N_14637);
nor UO_1620 (O_1620,N_14945,N_14649);
and UO_1621 (O_1621,N_14858,N_14544);
and UO_1622 (O_1622,N_14817,N_14510);
nand UO_1623 (O_1623,N_14930,N_14778);
and UO_1624 (O_1624,N_14563,N_14710);
nor UO_1625 (O_1625,N_14819,N_14823);
xnor UO_1626 (O_1626,N_14875,N_14978);
and UO_1627 (O_1627,N_14914,N_14761);
and UO_1628 (O_1628,N_14578,N_14536);
and UO_1629 (O_1629,N_14743,N_14644);
xnor UO_1630 (O_1630,N_14940,N_14659);
nor UO_1631 (O_1631,N_14849,N_14892);
nand UO_1632 (O_1632,N_14619,N_14944);
or UO_1633 (O_1633,N_14525,N_14563);
nor UO_1634 (O_1634,N_14540,N_14980);
and UO_1635 (O_1635,N_14961,N_14531);
or UO_1636 (O_1636,N_14605,N_14556);
or UO_1637 (O_1637,N_14911,N_14682);
xor UO_1638 (O_1638,N_14879,N_14639);
nand UO_1639 (O_1639,N_14977,N_14922);
nor UO_1640 (O_1640,N_14955,N_14594);
and UO_1641 (O_1641,N_14851,N_14592);
and UO_1642 (O_1642,N_14995,N_14527);
or UO_1643 (O_1643,N_14878,N_14734);
or UO_1644 (O_1644,N_14710,N_14572);
and UO_1645 (O_1645,N_14548,N_14950);
and UO_1646 (O_1646,N_14540,N_14534);
nand UO_1647 (O_1647,N_14811,N_14847);
xor UO_1648 (O_1648,N_14996,N_14569);
nand UO_1649 (O_1649,N_14709,N_14537);
nand UO_1650 (O_1650,N_14786,N_14794);
nand UO_1651 (O_1651,N_14816,N_14901);
nor UO_1652 (O_1652,N_14603,N_14672);
nor UO_1653 (O_1653,N_14570,N_14817);
nor UO_1654 (O_1654,N_14907,N_14573);
nand UO_1655 (O_1655,N_14811,N_14650);
or UO_1656 (O_1656,N_14770,N_14515);
nand UO_1657 (O_1657,N_14906,N_14666);
or UO_1658 (O_1658,N_14606,N_14522);
nor UO_1659 (O_1659,N_14965,N_14504);
nor UO_1660 (O_1660,N_14512,N_14793);
nand UO_1661 (O_1661,N_14764,N_14979);
xnor UO_1662 (O_1662,N_14943,N_14530);
or UO_1663 (O_1663,N_14653,N_14643);
and UO_1664 (O_1664,N_14622,N_14642);
and UO_1665 (O_1665,N_14587,N_14939);
nand UO_1666 (O_1666,N_14875,N_14829);
and UO_1667 (O_1667,N_14858,N_14974);
nand UO_1668 (O_1668,N_14943,N_14747);
nor UO_1669 (O_1669,N_14510,N_14864);
xnor UO_1670 (O_1670,N_14790,N_14728);
nand UO_1671 (O_1671,N_14834,N_14928);
xnor UO_1672 (O_1672,N_14615,N_14715);
or UO_1673 (O_1673,N_14879,N_14550);
nand UO_1674 (O_1674,N_14515,N_14745);
nand UO_1675 (O_1675,N_14833,N_14864);
nand UO_1676 (O_1676,N_14512,N_14780);
nor UO_1677 (O_1677,N_14775,N_14534);
and UO_1678 (O_1678,N_14852,N_14779);
nand UO_1679 (O_1679,N_14759,N_14504);
nand UO_1680 (O_1680,N_14719,N_14611);
nor UO_1681 (O_1681,N_14533,N_14695);
nand UO_1682 (O_1682,N_14723,N_14975);
or UO_1683 (O_1683,N_14712,N_14745);
or UO_1684 (O_1684,N_14966,N_14813);
nand UO_1685 (O_1685,N_14824,N_14793);
nand UO_1686 (O_1686,N_14705,N_14867);
xnor UO_1687 (O_1687,N_14862,N_14632);
nor UO_1688 (O_1688,N_14535,N_14710);
nor UO_1689 (O_1689,N_14642,N_14844);
and UO_1690 (O_1690,N_14974,N_14646);
nand UO_1691 (O_1691,N_14909,N_14565);
nand UO_1692 (O_1692,N_14891,N_14732);
nor UO_1693 (O_1693,N_14687,N_14824);
or UO_1694 (O_1694,N_14579,N_14528);
nor UO_1695 (O_1695,N_14799,N_14611);
nand UO_1696 (O_1696,N_14582,N_14630);
xnor UO_1697 (O_1697,N_14586,N_14983);
and UO_1698 (O_1698,N_14557,N_14933);
xnor UO_1699 (O_1699,N_14650,N_14985);
and UO_1700 (O_1700,N_14567,N_14688);
or UO_1701 (O_1701,N_14968,N_14827);
or UO_1702 (O_1702,N_14755,N_14964);
or UO_1703 (O_1703,N_14721,N_14674);
and UO_1704 (O_1704,N_14894,N_14989);
and UO_1705 (O_1705,N_14990,N_14722);
and UO_1706 (O_1706,N_14976,N_14578);
nand UO_1707 (O_1707,N_14954,N_14683);
and UO_1708 (O_1708,N_14600,N_14533);
or UO_1709 (O_1709,N_14743,N_14875);
and UO_1710 (O_1710,N_14563,N_14981);
and UO_1711 (O_1711,N_14897,N_14628);
or UO_1712 (O_1712,N_14644,N_14792);
nand UO_1713 (O_1713,N_14958,N_14748);
nand UO_1714 (O_1714,N_14821,N_14755);
or UO_1715 (O_1715,N_14526,N_14631);
nor UO_1716 (O_1716,N_14546,N_14701);
and UO_1717 (O_1717,N_14682,N_14802);
nand UO_1718 (O_1718,N_14758,N_14751);
nor UO_1719 (O_1719,N_14612,N_14626);
or UO_1720 (O_1720,N_14931,N_14817);
nand UO_1721 (O_1721,N_14873,N_14505);
and UO_1722 (O_1722,N_14605,N_14844);
nor UO_1723 (O_1723,N_14622,N_14588);
nor UO_1724 (O_1724,N_14791,N_14838);
or UO_1725 (O_1725,N_14620,N_14637);
and UO_1726 (O_1726,N_14690,N_14746);
and UO_1727 (O_1727,N_14916,N_14760);
nand UO_1728 (O_1728,N_14822,N_14519);
and UO_1729 (O_1729,N_14615,N_14832);
nor UO_1730 (O_1730,N_14974,N_14654);
nor UO_1731 (O_1731,N_14741,N_14691);
nor UO_1732 (O_1732,N_14832,N_14720);
or UO_1733 (O_1733,N_14751,N_14723);
nand UO_1734 (O_1734,N_14830,N_14750);
xor UO_1735 (O_1735,N_14718,N_14808);
nand UO_1736 (O_1736,N_14976,N_14987);
and UO_1737 (O_1737,N_14798,N_14838);
or UO_1738 (O_1738,N_14662,N_14534);
nand UO_1739 (O_1739,N_14889,N_14994);
or UO_1740 (O_1740,N_14728,N_14604);
nor UO_1741 (O_1741,N_14743,N_14887);
and UO_1742 (O_1742,N_14779,N_14722);
xnor UO_1743 (O_1743,N_14525,N_14890);
and UO_1744 (O_1744,N_14773,N_14796);
nand UO_1745 (O_1745,N_14832,N_14913);
and UO_1746 (O_1746,N_14977,N_14636);
nor UO_1747 (O_1747,N_14521,N_14916);
nand UO_1748 (O_1748,N_14687,N_14973);
and UO_1749 (O_1749,N_14858,N_14881);
or UO_1750 (O_1750,N_14822,N_14659);
or UO_1751 (O_1751,N_14500,N_14606);
and UO_1752 (O_1752,N_14946,N_14561);
nand UO_1753 (O_1753,N_14740,N_14847);
nor UO_1754 (O_1754,N_14811,N_14750);
or UO_1755 (O_1755,N_14911,N_14741);
xnor UO_1756 (O_1756,N_14685,N_14749);
nand UO_1757 (O_1757,N_14669,N_14867);
or UO_1758 (O_1758,N_14719,N_14755);
and UO_1759 (O_1759,N_14725,N_14988);
xor UO_1760 (O_1760,N_14933,N_14649);
or UO_1761 (O_1761,N_14828,N_14656);
nor UO_1762 (O_1762,N_14920,N_14621);
nand UO_1763 (O_1763,N_14710,N_14849);
nor UO_1764 (O_1764,N_14537,N_14780);
nand UO_1765 (O_1765,N_14582,N_14567);
and UO_1766 (O_1766,N_14901,N_14618);
and UO_1767 (O_1767,N_14977,N_14664);
and UO_1768 (O_1768,N_14600,N_14913);
or UO_1769 (O_1769,N_14744,N_14536);
xnor UO_1770 (O_1770,N_14733,N_14824);
nor UO_1771 (O_1771,N_14821,N_14609);
xnor UO_1772 (O_1772,N_14584,N_14970);
nand UO_1773 (O_1773,N_14962,N_14998);
nor UO_1774 (O_1774,N_14604,N_14707);
nor UO_1775 (O_1775,N_14797,N_14595);
and UO_1776 (O_1776,N_14515,N_14514);
or UO_1777 (O_1777,N_14859,N_14597);
and UO_1778 (O_1778,N_14779,N_14738);
and UO_1779 (O_1779,N_14566,N_14578);
nand UO_1780 (O_1780,N_14864,N_14939);
nor UO_1781 (O_1781,N_14785,N_14783);
or UO_1782 (O_1782,N_14547,N_14777);
and UO_1783 (O_1783,N_14819,N_14877);
and UO_1784 (O_1784,N_14583,N_14895);
nand UO_1785 (O_1785,N_14720,N_14638);
nor UO_1786 (O_1786,N_14926,N_14898);
nand UO_1787 (O_1787,N_14902,N_14598);
and UO_1788 (O_1788,N_14829,N_14603);
nand UO_1789 (O_1789,N_14705,N_14584);
and UO_1790 (O_1790,N_14598,N_14828);
nand UO_1791 (O_1791,N_14592,N_14835);
xor UO_1792 (O_1792,N_14691,N_14502);
nand UO_1793 (O_1793,N_14957,N_14788);
or UO_1794 (O_1794,N_14950,N_14636);
nand UO_1795 (O_1795,N_14762,N_14532);
or UO_1796 (O_1796,N_14713,N_14787);
nor UO_1797 (O_1797,N_14948,N_14856);
or UO_1798 (O_1798,N_14874,N_14635);
xor UO_1799 (O_1799,N_14636,N_14578);
or UO_1800 (O_1800,N_14691,N_14749);
or UO_1801 (O_1801,N_14700,N_14964);
nor UO_1802 (O_1802,N_14848,N_14827);
nor UO_1803 (O_1803,N_14783,N_14808);
and UO_1804 (O_1804,N_14780,N_14839);
or UO_1805 (O_1805,N_14612,N_14871);
nand UO_1806 (O_1806,N_14986,N_14500);
nor UO_1807 (O_1807,N_14708,N_14783);
nor UO_1808 (O_1808,N_14619,N_14746);
nor UO_1809 (O_1809,N_14598,N_14520);
nor UO_1810 (O_1810,N_14540,N_14662);
nand UO_1811 (O_1811,N_14883,N_14845);
nand UO_1812 (O_1812,N_14672,N_14764);
or UO_1813 (O_1813,N_14589,N_14949);
or UO_1814 (O_1814,N_14577,N_14800);
or UO_1815 (O_1815,N_14681,N_14650);
xnor UO_1816 (O_1816,N_14562,N_14654);
or UO_1817 (O_1817,N_14929,N_14967);
and UO_1818 (O_1818,N_14699,N_14927);
xnor UO_1819 (O_1819,N_14907,N_14903);
and UO_1820 (O_1820,N_14927,N_14616);
xnor UO_1821 (O_1821,N_14723,N_14748);
and UO_1822 (O_1822,N_14857,N_14532);
nor UO_1823 (O_1823,N_14509,N_14985);
and UO_1824 (O_1824,N_14874,N_14610);
nor UO_1825 (O_1825,N_14961,N_14912);
or UO_1826 (O_1826,N_14836,N_14842);
and UO_1827 (O_1827,N_14783,N_14565);
nor UO_1828 (O_1828,N_14859,N_14899);
nand UO_1829 (O_1829,N_14642,N_14564);
nor UO_1830 (O_1830,N_14689,N_14586);
nand UO_1831 (O_1831,N_14519,N_14557);
and UO_1832 (O_1832,N_14865,N_14532);
nand UO_1833 (O_1833,N_14995,N_14787);
or UO_1834 (O_1834,N_14851,N_14524);
and UO_1835 (O_1835,N_14517,N_14759);
and UO_1836 (O_1836,N_14952,N_14872);
nand UO_1837 (O_1837,N_14757,N_14743);
nand UO_1838 (O_1838,N_14855,N_14511);
nor UO_1839 (O_1839,N_14557,N_14886);
nor UO_1840 (O_1840,N_14946,N_14730);
or UO_1841 (O_1841,N_14969,N_14562);
nor UO_1842 (O_1842,N_14998,N_14519);
xor UO_1843 (O_1843,N_14813,N_14869);
nor UO_1844 (O_1844,N_14880,N_14711);
nand UO_1845 (O_1845,N_14862,N_14965);
xnor UO_1846 (O_1846,N_14965,N_14531);
and UO_1847 (O_1847,N_14794,N_14875);
nor UO_1848 (O_1848,N_14742,N_14562);
nand UO_1849 (O_1849,N_14788,N_14611);
nand UO_1850 (O_1850,N_14970,N_14653);
nor UO_1851 (O_1851,N_14534,N_14984);
or UO_1852 (O_1852,N_14869,N_14876);
xor UO_1853 (O_1853,N_14960,N_14956);
and UO_1854 (O_1854,N_14758,N_14861);
nand UO_1855 (O_1855,N_14937,N_14885);
and UO_1856 (O_1856,N_14642,N_14545);
and UO_1857 (O_1857,N_14816,N_14522);
nand UO_1858 (O_1858,N_14528,N_14529);
or UO_1859 (O_1859,N_14786,N_14533);
nor UO_1860 (O_1860,N_14926,N_14618);
nor UO_1861 (O_1861,N_14884,N_14709);
nor UO_1862 (O_1862,N_14854,N_14880);
nand UO_1863 (O_1863,N_14886,N_14713);
nor UO_1864 (O_1864,N_14523,N_14511);
nand UO_1865 (O_1865,N_14937,N_14729);
nor UO_1866 (O_1866,N_14749,N_14518);
nand UO_1867 (O_1867,N_14682,N_14935);
nand UO_1868 (O_1868,N_14877,N_14684);
and UO_1869 (O_1869,N_14555,N_14992);
xnor UO_1870 (O_1870,N_14767,N_14548);
nand UO_1871 (O_1871,N_14787,N_14654);
nand UO_1872 (O_1872,N_14632,N_14532);
and UO_1873 (O_1873,N_14604,N_14519);
nand UO_1874 (O_1874,N_14906,N_14966);
or UO_1875 (O_1875,N_14919,N_14634);
and UO_1876 (O_1876,N_14947,N_14871);
and UO_1877 (O_1877,N_14798,N_14814);
and UO_1878 (O_1878,N_14981,N_14965);
or UO_1879 (O_1879,N_14796,N_14984);
or UO_1880 (O_1880,N_14591,N_14550);
or UO_1881 (O_1881,N_14711,N_14545);
nand UO_1882 (O_1882,N_14556,N_14648);
nand UO_1883 (O_1883,N_14575,N_14887);
or UO_1884 (O_1884,N_14813,N_14505);
xnor UO_1885 (O_1885,N_14757,N_14999);
or UO_1886 (O_1886,N_14641,N_14748);
or UO_1887 (O_1887,N_14568,N_14648);
and UO_1888 (O_1888,N_14897,N_14526);
or UO_1889 (O_1889,N_14820,N_14832);
nor UO_1890 (O_1890,N_14719,N_14592);
nand UO_1891 (O_1891,N_14524,N_14740);
or UO_1892 (O_1892,N_14732,N_14976);
nand UO_1893 (O_1893,N_14684,N_14502);
nand UO_1894 (O_1894,N_14512,N_14830);
xnor UO_1895 (O_1895,N_14882,N_14852);
and UO_1896 (O_1896,N_14612,N_14585);
and UO_1897 (O_1897,N_14613,N_14830);
or UO_1898 (O_1898,N_14530,N_14535);
nand UO_1899 (O_1899,N_14969,N_14703);
and UO_1900 (O_1900,N_14582,N_14955);
xnor UO_1901 (O_1901,N_14741,N_14900);
and UO_1902 (O_1902,N_14905,N_14893);
or UO_1903 (O_1903,N_14946,N_14630);
nand UO_1904 (O_1904,N_14648,N_14675);
and UO_1905 (O_1905,N_14772,N_14784);
and UO_1906 (O_1906,N_14800,N_14512);
nand UO_1907 (O_1907,N_14610,N_14690);
or UO_1908 (O_1908,N_14597,N_14814);
nand UO_1909 (O_1909,N_14984,N_14716);
or UO_1910 (O_1910,N_14577,N_14792);
and UO_1911 (O_1911,N_14943,N_14760);
nor UO_1912 (O_1912,N_14899,N_14636);
or UO_1913 (O_1913,N_14742,N_14596);
nor UO_1914 (O_1914,N_14995,N_14828);
nand UO_1915 (O_1915,N_14942,N_14790);
nor UO_1916 (O_1916,N_14863,N_14988);
or UO_1917 (O_1917,N_14797,N_14855);
nor UO_1918 (O_1918,N_14585,N_14952);
nor UO_1919 (O_1919,N_14752,N_14764);
and UO_1920 (O_1920,N_14698,N_14709);
xnor UO_1921 (O_1921,N_14980,N_14911);
xnor UO_1922 (O_1922,N_14910,N_14974);
nand UO_1923 (O_1923,N_14895,N_14926);
nand UO_1924 (O_1924,N_14899,N_14985);
or UO_1925 (O_1925,N_14593,N_14998);
and UO_1926 (O_1926,N_14785,N_14904);
nor UO_1927 (O_1927,N_14603,N_14670);
and UO_1928 (O_1928,N_14525,N_14520);
nand UO_1929 (O_1929,N_14567,N_14873);
or UO_1930 (O_1930,N_14559,N_14725);
and UO_1931 (O_1931,N_14754,N_14805);
nor UO_1932 (O_1932,N_14795,N_14783);
nor UO_1933 (O_1933,N_14906,N_14668);
xor UO_1934 (O_1934,N_14735,N_14575);
nor UO_1935 (O_1935,N_14903,N_14807);
nand UO_1936 (O_1936,N_14779,N_14778);
and UO_1937 (O_1937,N_14776,N_14851);
nor UO_1938 (O_1938,N_14518,N_14684);
and UO_1939 (O_1939,N_14535,N_14942);
or UO_1940 (O_1940,N_14747,N_14643);
and UO_1941 (O_1941,N_14880,N_14521);
and UO_1942 (O_1942,N_14826,N_14684);
nand UO_1943 (O_1943,N_14830,N_14805);
nand UO_1944 (O_1944,N_14800,N_14628);
xor UO_1945 (O_1945,N_14711,N_14517);
nand UO_1946 (O_1946,N_14985,N_14778);
xnor UO_1947 (O_1947,N_14689,N_14911);
and UO_1948 (O_1948,N_14957,N_14505);
and UO_1949 (O_1949,N_14622,N_14876);
and UO_1950 (O_1950,N_14637,N_14945);
nand UO_1951 (O_1951,N_14637,N_14561);
xor UO_1952 (O_1952,N_14792,N_14877);
xor UO_1953 (O_1953,N_14826,N_14563);
xor UO_1954 (O_1954,N_14547,N_14647);
nand UO_1955 (O_1955,N_14579,N_14539);
and UO_1956 (O_1956,N_14597,N_14587);
nor UO_1957 (O_1957,N_14830,N_14539);
nor UO_1958 (O_1958,N_14651,N_14809);
nand UO_1959 (O_1959,N_14513,N_14840);
or UO_1960 (O_1960,N_14763,N_14958);
nor UO_1961 (O_1961,N_14777,N_14862);
nor UO_1962 (O_1962,N_14748,N_14822);
or UO_1963 (O_1963,N_14759,N_14912);
nand UO_1964 (O_1964,N_14778,N_14740);
nor UO_1965 (O_1965,N_14996,N_14672);
or UO_1966 (O_1966,N_14555,N_14800);
nor UO_1967 (O_1967,N_14833,N_14772);
or UO_1968 (O_1968,N_14899,N_14994);
nor UO_1969 (O_1969,N_14884,N_14714);
and UO_1970 (O_1970,N_14995,N_14540);
nor UO_1971 (O_1971,N_14593,N_14586);
nand UO_1972 (O_1972,N_14595,N_14674);
or UO_1973 (O_1973,N_14613,N_14940);
nor UO_1974 (O_1974,N_14908,N_14737);
nand UO_1975 (O_1975,N_14723,N_14698);
and UO_1976 (O_1976,N_14962,N_14754);
nand UO_1977 (O_1977,N_14734,N_14601);
nor UO_1978 (O_1978,N_14564,N_14983);
or UO_1979 (O_1979,N_14869,N_14589);
or UO_1980 (O_1980,N_14927,N_14877);
and UO_1981 (O_1981,N_14563,N_14906);
nand UO_1982 (O_1982,N_14804,N_14715);
nand UO_1983 (O_1983,N_14512,N_14708);
nor UO_1984 (O_1984,N_14726,N_14720);
xor UO_1985 (O_1985,N_14820,N_14536);
nand UO_1986 (O_1986,N_14765,N_14907);
xnor UO_1987 (O_1987,N_14882,N_14932);
and UO_1988 (O_1988,N_14723,N_14876);
or UO_1989 (O_1989,N_14835,N_14552);
and UO_1990 (O_1990,N_14607,N_14832);
nor UO_1991 (O_1991,N_14778,N_14671);
xor UO_1992 (O_1992,N_14872,N_14665);
nand UO_1993 (O_1993,N_14856,N_14704);
and UO_1994 (O_1994,N_14940,N_14571);
nor UO_1995 (O_1995,N_14685,N_14940);
xnor UO_1996 (O_1996,N_14851,N_14811);
or UO_1997 (O_1997,N_14970,N_14638);
and UO_1998 (O_1998,N_14871,N_14948);
and UO_1999 (O_1999,N_14791,N_14994);
endmodule