module basic_1500_15000_2000_30_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_146,In_30);
nor U1 (N_1,In_62,In_1007);
and U2 (N_2,In_348,In_547);
or U3 (N_3,In_463,In_950);
nor U4 (N_4,In_1236,In_944);
and U5 (N_5,In_585,In_1112);
and U6 (N_6,In_374,In_921);
nand U7 (N_7,In_508,In_1443);
xnor U8 (N_8,In_1111,In_1263);
nand U9 (N_9,In_1071,In_928);
nand U10 (N_10,In_1070,In_229);
or U11 (N_11,In_534,In_1259);
or U12 (N_12,In_973,In_175);
or U13 (N_13,In_1093,In_1412);
nor U14 (N_14,In_1434,In_1358);
nor U15 (N_15,In_65,In_37);
nand U16 (N_16,In_717,In_92);
nand U17 (N_17,In_600,In_1401);
or U18 (N_18,In_1425,In_616);
nor U19 (N_19,In_510,In_842);
and U20 (N_20,In_595,In_98);
xnor U21 (N_21,In_50,In_527);
or U22 (N_22,In_380,In_1229);
and U23 (N_23,In_1058,In_957);
nor U24 (N_24,In_16,In_1035);
or U25 (N_25,In_912,In_704);
and U26 (N_26,In_59,In_919);
xor U27 (N_27,In_1329,In_556);
nand U28 (N_28,In_1497,In_896);
xnor U29 (N_29,In_856,In_138);
or U30 (N_30,In_1364,In_284);
xor U31 (N_31,In_642,In_975);
and U32 (N_32,In_464,In_851);
and U33 (N_33,In_837,In_605);
nand U34 (N_34,In_750,In_1140);
xor U35 (N_35,In_95,In_1281);
and U36 (N_36,In_1465,In_264);
nor U37 (N_37,In_208,In_805);
nand U38 (N_38,In_291,In_143);
and U39 (N_39,In_447,In_583);
and U40 (N_40,In_772,In_309);
nand U41 (N_41,In_783,In_343);
xnor U42 (N_42,In_860,In_763);
and U43 (N_43,In_1261,In_158);
xnor U44 (N_44,In_659,In_573);
and U45 (N_45,In_360,In_259);
xor U46 (N_46,In_757,In_133);
or U47 (N_47,In_849,In_293);
xnor U48 (N_48,In_1242,In_410);
and U49 (N_49,In_1078,In_361);
or U50 (N_50,In_1493,In_793);
nand U51 (N_51,In_394,In_1410);
nand U52 (N_52,In_1210,In_330);
xnor U53 (N_53,In_1139,In_1415);
or U54 (N_54,In_370,In_1197);
or U55 (N_55,In_993,In_1137);
or U56 (N_56,In_1393,In_313);
nand U57 (N_57,In_375,In_416);
xnor U58 (N_58,In_674,In_771);
and U59 (N_59,In_115,In_672);
xnor U60 (N_60,In_1119,In_586);
nand U61 (N_61,In_415,In_577);
nor U62 (N_62,In_978,In_884);
or U63 (N_63,In_156,In_1349);
nand U64 (N_64,In_946,In_454);
and U65 (N_65,In_724,In_1160);
nand U66 (N_66,In_1278,In_269);
nor U67 (N_67,In_201,In_18);
and U68 (N_68,In_328,In_1190);
nor U69 (N_69,In_1082,In_575);
and U70 (N_70,In_1048,In_329);
nand U71 (N_71,In_1244,In_377);
nor U72 (N_72,In_1251,In_766);
and U73 (N_73,In_1227,In_1192);
xor U74 (N_74,In_632,In_404);
nand U75 (N_75,In_1057,In_446);
and U76 (N_76,In_1471,In_500);
and U77 (N_77,In_923,In_45);
nand U78 (N_78,In_644,In_352);
and U79 (N_79,In_714,In_916);
xor U80 (N_80,In_443,In_272);
nor U81 (N_81,In_637,In_738);
and U82 (N_82,In_211,In_1086);
xor U83 (N_83,In_1123,In_760);
nor U84 (N_84,In_384,In_1422);
or U85 (N_85,In_824,In_137);
and U86 (N_86,In_8,In_1310);
nand U87 (N_87,In_1447,In_1306);
xnor U88 (N_88,In_572,In_1234);
xnor U89 (N_89,In_273,In_1464);
nand U90 (N_90,In_1323,In_762);
and U91 (N_91,In_1146,In_816);
and U92 (N_92,In_233,In_578);
and U93 (N_93,In_807,In_867);
xnor U94 (N_94,In_283,In_13);
and U95 (N_95,In_1260,In_287);
and U96 (N_96,In_650,In_698);
nand U97 (N_97,In_207,In_1159);
or U98 (N_98,In_319,In_61);
and U99 (N_99,In_821,In_275);
and U100 (N_100,In_202,In_1025);
nor U101 (N_101,In_551,In_589);
nor U102 (N_102,In_46,In_1388);
nand U103 (N_103,In_883,In_186);
xnor U104 (N_104,In_524,In_1428);
and U105 (N_105,In_1418,In_1353);
nand U106 (N_106,In_231,In_88);
nor U107 (N_107,In_1013,In_480);
or U108 (N_108,In_1094,In_459);
nand U109 (N_109,In_693,In_1461);
and U110 (N_110,In_587,In_295);
nor U111 (N_111,In_70,In_1390);
and U112 (N_112,In_989,In_1382);
and U113 (N_113,In_132,In_1377);
nand U114 (N_114,In_362,In_200);
and U115 (N_115,In_943,In_1356);
or U116 (N_116,In_35,In_400);
nor U117 (N_117,In_890,In_1079);
nor U118 (N_118,In_103,In_1193);
xor U119 (N_119,In_533,In_1084);
xnor U120 (N_120,In_286,In_1352);
nand U121 (N_121,In_1335,In_20);
xnor U122 (N_122,In_703,In_1436);
nand U123 (N_123,In_1301,In_758);
and U124 (N_124,In_382,In_94);
or U125 (N_125,In_1168,In_838);
xor U126 (N_126,In_1188,In_880);
xor U127 (N_127,In_185,In_535);
nand U128 (N_128,In_241,In_876);
or U129 (N_129,In_184,In_696);
and U130 (N_130,In_429,In_811);
nor U131 (N_131,In_1402,In_326);
or U132 (N_132,In_280,In_746);
and U133 (N_133,In_1098,In_1017);
or U134 (N_134,In_615,In_685);
and U135 (N_135,In_297,In_176);
xnor U136 (N_136,In_1001,In_669);
and U137 (N_137,In_1470,In_761);
and U138 (N_138,In_188,In_791);
nor U139 (N_139,In_312,In_1172);
xor U140 (N_140,In_1099,In_633);
xor U141 (N_141,In_42,In_651);
nor U142 (N_142,In_647,In_1065);
nand U143 (N_143,In_658,In_1457);
and U144 (N_144,In_1296,In_920);
or U145 (N_145,In_89,In_435);
xor U146 (N_146,In_1423,In_260);
or U147 (N_147,In_308,In_141);
nor U148 (N_148,In_321,In_496);
or U149 (N_149,In_1325,In_356);
xor U150 (N_150,In_1435,In_1265);
nor U151 (N_151,In_423,In_1297);
or U152 (N_152,In_933,In_1004);
and U153 (N_153,In_1472,In_5);
nor U154 (N_154,In_433,In_1042);
nor U155 (N_155,In_827,In_870);
xor U156 (N_156,In_378,In_774);
nand U157 (N_157,In_419,In_1161);
and U158 (N_158,In_549,In_203);
or U159 (N_159,In_1187,In_187);
xnor U160 (N_160,In_351,In_740);
xor U161 (N_161,In_1459,In_1037);
or U162 (N_162,In_335,In_492);
and U163 (N_163,In_1338,In_1432);
nand U164 (N_164,In_952,In_1373);
xnor U165 (N_165,In_1487,In_931);
xor U166 (N_166,In_1419,In_1149);
xor U167 (N_167,In_1092,In_624);
nand U168 (N_168,In_1274,In_1273);
nand U169 (N_169,In_1134,In_408);
and U170 (N_170,In_1406,In_1468);
nor U171 (N_171,In_246,In_521);
nor U172 (N_172,In_1305,In_1153);
nor U173 (N_173,In_1262,In_1087);
xor U174 (N_174,In_691,In_179);
nand U175 (N_175,In_1315,In_582);
xnor U176 (N_176,In_1345,In_1346);
xor U177 (N_177,In_1043,In_1431);
and U178 (N_178,In_1330,In_213);
or U179 (N_179,In_1199,In_662);
xnor U180 (N_180,In_266,In_1289);
xnor U181 (N_181,In_610,In_28);
nand U182 (N_182,In_546,In_990);
or U183 (N_183,In_1176,In_1253);
or U184 (N_184,In_236,In_889);
and U185 (N_185,In_972,In_550);
or U186 (N_186,In_317,In_116);
xor U187 (N_187,In_739,In_1113);
or U188 (N_188,In_265,In_281);
nor U189 (N_189,In_1005,In_1298);
nand U190 (N_190,In_1152,In_1022);
and U191 (N_191,In_53,In_707);
xnor U192 (N_192,In_609,In_1238);
and U193 (N_193,In_1361,In_1075);
and U194 (N_194,In_1342,In_153);
nor U195 (N_195,In_965,In_336);
and U196 (N_196,In_548,In_1339);
xor U197 (N_197,In_695,In_1209);
nor U198 (N_198,In_392,In_801);
xor U199 (N_199,In_819,In_561);
and U200 (N_200,In_56,In_4);
xnor U201 (N_201,In_372,In_413);
or U202 (N_202,In_1453,In_1105);
and U203 (N_203,In_748,In_1135);
nor U204 (N_204,In_1375,In_1291);
nor U205 (N_205,In_31,In_1129);
nand U206 (N_206,In_1174,In_1029);
nor U207 (N_207,In_537,In_412);
nand U208 (N_208,In_205,In_77);
or U209 (N_209,In_1055,In_14);
and U210 (N_210,In_618,In_671);
nor U211 (N_211,In_1317,In_1398);
and U212 (N_212,In_249,In_1286);
and U213 (N_213,In_430,In_1151);
nor U214 (N_214,In_307,In_1107);
and U215 (N_215,In_723,In_894);
or U216 (N_216,In_1433,In_421);
and U217 (N_217,In_7,In_1072);
nand U218 (N_218,In_652,In_709);
nor U219 (N_219,In_1038,In_15);
nor U220 (N_220,In_1252,In_539);
or U221 (N_221,In_1407,In_1458);
xnor U222 (N_222,In_344,In_778);
and U223 (N_223,In_1002,In_230);
or U224 (N_224,In_84,In_134);
xor U225 (N_225,In_1378,In_514);
nand U226 (N_226,In_457,In_574);
nor U227 (N_227,In_892,In_840);
nor U228 (N_228,In_1277,In_171);
or U229 (N_229,In_694,In_545);
xor U230 (N_230,In_75,In_123);
nor U231 (N_231,In_914,In_555);
and U232 (N_232,In_1125,In_515);
or U233 (N_233,In_562,In_1491);
and U234 (N_234,In_441,In_903);
or U235 (N_235,In_663,In_1343);
nand U236 (N_236,In_1056,In_478);
or U237 (N_237,In_1040,In_263);
or U238 (N_238,In_1416,In_497);
nand U239 (N_239,In_544,In_794);
or U240 (N_240,In_718,In_768);
and U241 (N_241,In_985,In_994);
or U242 (N_242,In_861,In_87);
and U243 (N_243,In_974,In_1223);
and U244 (N_244,In_1327,In_1429);
nor U245 (N_245,In_962,In_1308);
nor U246 (N_246,In_210,In_1336);
nand U247 (N_247,In_887,In_10);
and U248 (N_248,In_522,In_225);
or U249 (N_249,In_1316,In_1130);
nand U250 (N_250,In_1050,In_9);
or U251 (N_251,In_212,In_949);
nand U252 (N_252,In_64,In_1387);
nand U253 (N_253,In_398,In_1167);
or U254 (N_254,In_221,In_216);
xnor U255 (N_255,In_571,In_345);
or U256 (N_256,In_773,In_1163);
xnor U257 (N_257,In_301,In_1103);
nand U258 (N_258,In_409,In_1304);
nor U259 (N_259,In_1359,In_756);
and U260 (N_260,In_40,In_466);
and U261 (N_261,In_1276,In_741);
xnor U262 (N_262,In_1053,In_1489);
and U263 (N_263,In_63,In_1031);
and U264 (N_264,In_67,In_11);
xor U265 (N_265,In_683,In_487);
nor U266 (N_266,In_190,In_596);
and U267 (N_267,In_44,In_970);
nand U268 (N_268,In_1269,In_822);
and U269 (N_269,In_787,In_646);
nand U270 (N_270,In_523,In_73);
nor U271 (N_271,In_125,In_204);
and U272 (N_272,In_1404,In_479);
or U273 (N_273,In_969,In_1488);
or U274 (N_274,In_238,In_1138);
or U275 (N_275,In_366,In_243);
and U276 (N_276,In_611,In_1030);
or U277 (N_277,In_135,In_486);
or U278 (N_278,In_701,In_834);
nand U279 (N_279,In_802,In_1181);
xor U280 (N_280,In_667,In_1397);
xor U281 (N_281,In_1104,In_954);
or U282 (N_282,In_491,In_854);
or U283 (N_283,In_414,In_630);
and U284 (N_284,In_1391,In_1196);
nand U285 (N_285,In_1219,In_648);
nand U286 (N_286,In_1462,In_355);
or U287 (N_287,In_924,In_909);
xnor U288 (N_288,In_159,In_654);
or U289 (N_289,In_407,In_489);
xor U290 (N_290,In_1108,In_399);
nand U291 (N_291,In_1365,In_961);
or U292 (N_292,In_237,In_1367);
and U293 (N_293,In_1283,In_966);
and U294 (N_294,In_729,In_730);
nand U295 (N_295,In_784,In_782);
and U296 (N_296,In_1486,In_1456);
or U297 (N_297,In_641,In_96);
or U298 (N_298,In_1216,In_1062);
or U299 (N_299,In_1073,In_769);
and U300 (N_300,In_476,In_918);
or U301 (N_301,In_1085,In_1191);
or U302 (N_302,In_980,In_113);
nor U303 (N_303,In_905,In_1148);
nor U304 (N_304,In_1214,In_482);
or U305 (N_305,In_1426,In_277);
or U306 (N_306,In_679,In_566);
xnor U307 (N_307,In_367,In_258);
and U308 (N_308,In_104,In_626);
xor U309 (N_309,In_1424,In_311);
and U310 (N_310,In_450,In_222);
nor U311 (N_311,In_604,In_684);
nor U312 (N_312,In_458,In_1246);
xor U313 (N_313,In_350,In_196);
nor U314 (N_314,In_1376,In_41);
and U315 (N_315,In_1088,In_1201);
or U316 (N_316,In_737,In_431);
xor U317 (N_317,In_1386,In_1309);
or U318 (N_318,In_1240,In_559);
or U319 (N_319,In_720,In_417);
nor U320 (N_320,In_149,In_371);
or U321 (N_321,In_1155,In_1385);
nand U322 (N_322,In_178,In_625);
nand U323 (N_323,In_795,In_1446);
nand U324 (N_324,In_942,In_1028);
and U325 (N_325,In_560,In_1363);
nor U326 (N_326,In_1403,In_682);
xnor U327 (N_327,In_937,In_434);
nand U328 (N_328,In_47,In_438);
and U329 (N_329,In_51,In_1469);
xnor U330 (N_330,In_468,In_661);
nor U331 (N_331,In_437,In_987);
and U332 (N_332,In_710,In_1200);
nand U333 (N_333,In_726,In_1354);
xor U334 (N_334,In_456,In_1019);
or U335 (N_335,In_1067,In_1369);
nand U336 (N_336,In_316,In_192);
nor U337 (N_337,In_906,In_529);
and U338 (N_338,In_655,In_1206);
nor U339 (N_339,In_1097,In_908);
and U340 (N_340,In_217,In_553);
or U341 (N_341,In_797,In_557);
xnor U342 (N_342,In_1280,In_494);
nand U343 (N_343,In_499,In_744);
xor U344 (N_344,In_991,In_1101);
and U345 (N_345,In_488,In_1466);
nor U346 (N_346,In_91,In_675);
nand U347 (N_347,In_292,In_697);
xor U348 (N_348,In_1384,In_907);
nor U349 (N_349,In_227,In_1215);
xor U350 (N_350,In_588,In_99);
nor U351 (N_351,In_379,In_1454);
xnor U352 (N_352,In_1408,In_580);
nand U353 (N_353,In_1449,In_107);
nor U354 (N_354,In_1485,In_779);
xnor U355 (N_355,In_988,In_953);
and U356 (N_356,In_365,In_393);
or U357 (N_357,In_39,In_1165);
nor U358 (N_358,In_182,In_34);
and U359 (N_359,In_1221,In_747);
nor U360 (N_360,In_341,In_1066);
or U361 (N_361,In_608,In_1313);
and U362 (N_362,In_242,In_340);
and U363 (N_363,In_245,In_1496);
nor U364 (N_364,In_1026,In_80);
nand U365 (N_365,In_1083,In_114);
nor U366 (N_366,In_855,In_79);
nand U367 (N_367,In_564,In_52);
nor U368 (N_368,In_1347,In_623);
and U369 (N_369,In_823,In_1194);
or U370 (N_370,In_670,In_1145);
xor U371 (N_371,In_964,In_531);
xnor U372 (N_372,In_590,In_131);
or U373 (N_373,In_228,In_955);
nand U374 (N_374,In_1178,In_247);
nor U375 (N_375,In_60,In_676);
or U376 (N_376,In_579,In_613);
nor U377 (N_377,In_1195,In_959);
nor U378 (N_378,In_1318,In_1324);
and U379 (N_379,In_152,In_38);
xnor U380 (N_380,In_29,In_893);
xnor U381 (N_381,In_1383,In_2);
or U382 (N_382,In_622,In_305);
nand U383 (N_383,In_460,In_294);
or U384 (N_384,In_353,In_1293);
nor U385 (N_385,In_917,In_299);
or U386 (N_386,In_424,In_567);
and U387 (N_387,In_518,In_879);
nand U388 (N_388,In_841,In_25);
or U389 (N_389,In_925,In_1302);
and U390 (N_390,In_358,In_1250);
or U391 (N_391,In_935,In_1015);
nand U392 (N_392,In_945,In_1414);
or U393 (N_393,In_1355,In_1245);
xnor U394 (N_394,In_664,In_1256);
nor U395 (N_395,In_81,In_1226);
nor U396 (N_396,In_1344,In_93);
nand U397 (N_397,In_922,In_183);
nor U398 (N_398,In_904,In_490);
nand U399 (N_399,In_144,In_1012);
xnor U400 (N_400,In_167,In_252);
nand U401 (N_401,In_677,In_1467);
xnor U402 (N_402,In_1440,In_1096);
nor U403 (N_403,In_984,In_495);
and U404 (N_404,In_689,In_285);
nand U405 (N_405,In_215,In_570);
nand U406 (N_406,In_1060,In_1483);
nor U407 (N_407,In_369,In_342);
xor U408 (N_408,In_23,In_325);
xnor U409 (N_409,In_498,In_1437);
nor U410 (N_410,In_767,In_310);
xnor U411 (N_411,In_1039,In_711);
nand U412 (N_412,In_898,In_770);
and U413 (N_413,In_1258,In_678);
and U414 (N_414,In_17,In_406);
xnor U415 (N_415,In_1303,In_139);
and U416 (N_416,In_727,In_591);
or U417 (N_417,In_552,In_1184);
or U418 (N_418,In_0,In_1064);
nand U419 (N_419,In_798,In_1292);
xnor U420 (N_420,In_349,In_1164);
nor U421 (N_421,In_160,In_72);
and U422 (N_422,In_452,In_828);
xor U423 (N_423,In_858,In_157);
or U424 (N_424,In_1224,In_716);
and U425 (N_425,In_124,In_532);
nor U426 (N_426,In_173,In_1285);
nor U427 (N_427,In_1047,In_1158);
nand U428 (N_428,In_373,In_318);
or U429 (N_429,In_174,In_1090);
nor U430 (N_430,In_765,In_472);
nand U431 (N_431,In_1332,In_1290);
xor U432 (N_432,In_220,In_83);
nand U433 (N_433,In_1212,In_992);
nand U434 (N_434,In_886,In_752);
and U435 (N_435,In_810,In_1198);
nand U436 (N_436,In_331,In_298);
nor U437 (N_437,In_1186,In_69);
nand U438 (N_438,In_1257,In_692);
xor U439 (N_439,In_815,In_1473);
or U440 (N_440,In_712,In_536);
or U441 (N_441,In_736,In_958);
nor U442 (N_442,In_1270,In_719);
nor U443 (N_443,In_599,In_279);
and U444 (N_444,In_812,In_1089);
nand U445 (N_445,In_323,In_733);
xor U446 (N_446,In_1170,In_785);
nor U447 (N_447,In_1314,In_592);
and U448 (N_448,In_1395,In_930);
nor U449 (N_449,In_1220,In_97);
nand U450 (N_450,In_68,In_1116);
and U451 (N_451,In_934,In_1463);
nor U452 (N_452,In_857,In_1307);
nor U453 (N_453,In_657,In_118);
xnor U454 (N_454,In_402,In_383);
nand U455 (N_455,In_565,In_1452);
nor U456 (N_456,In_108,In_1020);
nand U457 (N_457,In_289,In_859);
and U458 (N_458,In_198,In_830);
or U459 (N_459,In_983,In_197);
and U460 (N_460,In_645,In_1156);
nor U461 (N_461,In_90,In_1076);
nor U462 (N_462,In_558,In_977);
or U463 (N_463,In_1441,In_150);
and U464 (N_464,In_526,In_1173);
or U465 (N_465,In_274,In_913);
and U466 (N_466,In_168,In_866);
or U467 (N_467,In_130,In_1118);
nand U468 (N_468,In_1249,In_926);
or U469 (N_469,In_71,In_120);
nor U470 (N_470,In_449,In_806);
and U471 (N_471,In_799,In_1451);
or U472 (N_472,In_839,In_376);
or U473 (N_473,In_1427,In_620);
xnor U474 (N_474,In_1430,In_43);
nor U475 (N_475,In_1455,In_927);
or U476 (N_476,In_956,In_1366);
nor U477 (N_477,In_1008,In_538);
and U478 (N_478,In_528,In_1069);
and U479 (N_479,In_638,In_327);
xnor U480 (N_480,In_688,In_734);
nand U481 (N_481,In_3,In_1166);
nor U482 (N_482,In_475,In_938);
xor U483 (N_483,In_1208,In_951);
nor U484 (N_484,In_440,In_1032);
and U485 (N_485,In_877,In_1420);
and U486 (N_486,In_520,In_1009);
xnor U487 (N_487,In_147,In_296);
nand U488 (N_488,In_936,In_792);
nor U489 (N_489,In_1018,In_1484);
or U490 (N_490,In_1222,In_1237);
xnor U491 (N_491,In_1312,In_971);
or U492 (N_492,In_483,In_1045);
or U493 (N_493,In_554,In_902);
and U494 (N_494,In_254,In_395);
nor U495 (N_495,In_1442,In_1326);
nor U496 (N_496,In_1157,In_1490);
nor U497 (N_497,In_1109,In_1063);
nand U498 (N_498,In_915,In_1122);
and U499 (N_499,In_363,In_85);
xnor U500 (N_500,N_55,In_833);
nor U501 (N_501,In_232,N_325);
xor U502 (N_502,N_397,N_123);
nor U503 (N_503,N_89,N_31);
and U504 (N_504,In_875,N_283);
or U505 (N_505,N_68,N_497);
nor U506 (N_506,In_728,In_825);
nand U507 (N_507,N_227,In_453);
and U508 (N_508,N_212,In_255);
or U509 (N_509,N_475,N_157);
nand U510 (N_510,N_461,In_603);
and U511 (N_511,In_27,In_507);
and U512 (N_512,In_432,N_271);
or U513 (N_513,N_464,N_298);
xor U514 (N_514,N_113,N_71);
nand U515 (N_515,N_446,In_122);
nor U516 (N_516,N_57,In_708);
nand U517 (N_517,In_66,N_63);
and U518 (N_518,In_74,In_381);
and U519 (N_519,N_85,N_306);
nand U520 (N_520,N_178,In_881);
or U521 (N_521,In_885,N_20);
xor U522 (N_522,In_477,In_1254);
nand U523 (N_523,In_850,N_378);
xor U524 (N_524,In_1203,In_700);
and U525 (N_525,In_1478,In_1218);
or U526 (N_526,In_1255,In_177);
or U527 (N_527,In_397,In_161);
and U528 (N_528,In_148,In_389);
nor U529 (N_529,In_1341,N_204);
xnor U530 (N_530,N_303,N_53);
or U531 (N_531,In_1439,N_405);
or U532 (N_532,N_307,N_483);
nand U533 (N_533,N_67,In_1110);
nand U534 (N_534,N_291,In_1143);
or U535 (N_535,In_1479,In_627);
xnor U536 (N_536,In_1328,N_239);
nand U537 (N_537,N_290,N_442);
nand U538 (N_538,In_420,In_1077);
or U539 (N_539,In_1333,In_1337);
xor U540 (N_540,N_209,In_1474);
xor U541 (N_541,N_468,N_379);
or U542 (N_542,N_169,In_929);
xnor U543 (N_543,N_328,In_21);
and U544 (N_544,In_117,N_219);
nand U545 (N_545,In_223,N_134);
or U546 (N_546,In_872,In_78);
xor U547 (N_547,In_346,In_33);
xnor U548 (N_548,In_948,N_177);
xnor U549 (N_549,N_376,N_100);
nor U550 (N_550,N_214,N_234);
xnor U551 (N_551,In_428,N_5);
nor U552 (N_552,In_368,N_380);
or U553 (N_553,N_498,In_1154);
or U554 (N_554,N_355,N_324);
nand U555 (N_555,N_494,In_1272);
nand U556 (N_556,In_509,In_1127);
and U557 (N_557,N_79,N_462);
xor U558 (N_558,N_454,In_776);
nor U559 (N_559,In_1348,N_259);
and U560 (N_560,In_1340,N_285);
and U561 (N_561,In_112,N_488);
and U562 (N_562,N_215,In_1438);
nand U563 (N_563,N_81,N_149);
or U564 (N_564,In_1179,N_297);
and U565 (N_565,In_614,In_493);
xnor U566 (N_566,N_481,N_162);
xor U567 (N_567,In_194,In_54);
nor U568 (N_568,N_315,N_312);
nand U569 (N_569,N_491,In_322);
nor U570 (N_570,N_457,In_530);
or U571 (N_571,In_1000,In_219);
nor U572 (N_572,N_345,In_628);
nor U573 (N_573,N_484,N_64);
nor U574 (N_574,N_459,In_199);
and U575 (N_575,N_411,N_171);
nor U576 (N_576,N_479,In_270);
nand U577 (N_577,In_1231,In_502);
nor U578 (N_578,In_848,In_1106);
nand U579 (N_579,N_410,In_947);
nand U580 (N_580,N_409,N_24);
and U581 (N_581,In_789,N_407);
or U582 (N_582,N_168,In_649);
xnor U583 (N_583,N_106,N_116);
and U584 (N_584,In_110,In_1080);
or U585 (N_585,In_268,In_1027);
or U586 (N_586,In_722,In_941);
and U587 (N_587,In_1074,N_294);
nand U588 (N_588,In_781,N_29);
xor U589 (N_589,In_214,In_1011);
or U590 (N_590,N_66,In_332);
nor U591 (N_591,In_444,In_1264);
and U592 (N_592,In_940,N_301);
and U593 (N_593,N_318,In_339);
and U594 (N_594,In_981,N_34);
nand U595 (N_595,N_220,N_309);
xor U596 (N_596,N_16,N_363);
and U597 (N_597,In_660,In_12);
and U598 (N_598,N_404,N_438);
nor U599 (N_599,N_377,N_490);
nor U600 (N_600,N_286,In_470);
xor U601 (N_601,N_231,In_304);
nor U602 (N_602,In_218,In_818);
or U603 (N_603,N_384,In_844);
or U604 (N_604,N_279,In_804);
nand U605 (N_605,N_211,In_636);
and U606 (N_606,In_775,N_319);
nand U607 (N_607,N_458,In_1482);
nor U608 (N_608,In_576,N_323);
nand U609 (N_609,N_158,In_846);
nor U610 (N_610,In_1117,N_197);
xnor U611 (N_611,In_1126,N_87);
or U612 (N_612,In_999,In_864);
nor U613 (N_613,N_159,N_224);
and U614 (N_614,In_1182,In_1068);
or U615 (N_615,In_759,N_201);
or U616 (N_616,N_101,In_364);
xnor U617 (N_617,N_27,N_439);
or U618 (N_618,In_1175,N_469);
and U619 (N_619,In_1034,In_1334);
and U620 (N_620,In_982,In_895);
nand U621 (N_621,In_829,In_1169);
and U622 (N_622,N_449,N_332);
and U623 (N_623,N_73,N_186);
nand U624 (N_624,N_248,N_416);
nand U625 (N_625,N_75,In_1360);
xnor U626 (N_626,In_1010,In_735);
nor U627 (N_627,N_173,In_1217);
nor U628 (N_628,N_256,In_891);
or U629 (N_629,N_13,N_51);
or U630 (N_630,In_869,N_32);
and U631 (N_631,N_111,In_796);
xnor U632 (N_632,In_901,N_445);
nor U633 (N_633,N_15,In_786);
xor U634 (N_634,In_411,N_128);
xor U635 (N_635,In_455,N_262);
nor U636 (N_636,In_731,N_167);
nand U637 (N_637,In_597,In_584);
nand U638 (N_638,N_487,In_1295);
nand U639 (N_639,N_76,In_334);
nand U640 (N_640,N_225,In_1185);
xor U641 (N_641,In_163,N_130);
or U642 (N_642,N_499,N_147);
and U643 (N_643,N_473,In_826);
nand U644 (N_644,N_249,In_354);
xor U645 (N_645,N_496,N_391);
or U646 (N_646,N_402,In_832);
xor U647 (N_647,N_78,In_788);
nand U648 (N_648,N_143,N_389);
xor U649 (N_649,In_1396,N_174);
or U650 (N_650,In_1205,N_188);
and U651 (N_651,N_273,In_910);
or U652 (N_652,N_276,In_900);
or U653 (N_653,N_194,In_1033);
nor U654 (N_654,In_1021,In_1);
nor U655 (N_655,In_845,N_141);
nand U656 (N_656,N_436,N_199);
and U657 (N_657,N_47,N_403);
or U658 (N_658,N_435,N_69);
and U659 (N_659,N_299,N_295);
nor U660 (N_660,In_1409,N_396);
or U661 (N_661,In_1202,In_22);
xnor U662 (N_662,In_1311,In_1294);
or U663 (N_663,In_997,In_82);
xnor U664 (N_664,In_673,In_388);
nand U665 (N_665,In_813,In_1228);
nand U666 (N_666,In_963,N_181);
xor U667 (N_667,N_46,In_1357);
or U668 (N_668,N_62,N_243);
nor U669 (N_669,N_288,In_387);
xor U670 (N_670,In_142,In_1279);
xor U671 (N_671,N_421,In_180);
xor U672 (N_672,N_482,N_125);
or U673 (N_673,N_260,In_1495);
xor U674 (N_674,In_1460,N_360);
nand U675 (N_675,In_101,N_180);
and U676 (N_676,In_1372,In_1036);
and U677 (N_677,N_202,N_10);
nor U678 (N_678,In_1207,In_1091);
nand U679 (N_679,N_493,In_504);
xor U680 (N_680,N_210,N_118);
nand U681 (N_681,N_191,In_1183);
and U682 (N_682,N_444,In_814);
or U683 (N_683,In_598,N_151);
nand U684 (N_684,In_26,In_1180);
nand U685 (N_685,In_111,N_321);
xor U686 (N_686,In_852,In_1477);
nor U687 (N_687,In_154,N_49);
or U688 (N_688,In_612,In_911);
and U689 (N_689,In_235,In_418);
nand U690 (N_690,In_541,In_619);
nand U691 (N_691,N_59,N_369);
or U692 (N_692,N_337,In_448);
xor U693 (N_693,N_93,N_467);
xor U694 (N_694,In_878,N_278);
nor U695 (N_695,In_288,N_292);
xnor U696 (N_696,N_333,N_472);
nand U697 (N_697,N_423,N_373);
nand U698 (N_698,N_105,N_452);
xnor U699 (N_699,N_184,In_278);
or U700 (N_700,In_1476,N_0);
and U701 (N_701,N_140,In_1379);
or U702 (N_702,In_1371,In_639);
xor U703 (N_703,N_305,N_155);
nor U704 (N_704,In_1114,N_165);
nor U705 (N_705,N_183,N_386);
xnor U706 (N_706,N_182,In_871);
nand U707 (N_707,N_284,N_395);
nand U708 (N_708,N_103,In_1141);
and U709 (N_709,In_248,In_1150);
nor U710 (N_710,N_261,In_749);
nand U711 (N_711,In_445,N_175);
nor U712 (N_712,In_862,In_1322);
xor U713 (N_713,N_48,In_189);
or U714 (N_714,N_372,N_1);
and U715 (N_715,In_581,N_86);
nand U716 (N_716,In_1006,In_803);
nor U717 (N_717,In_338,N_23);
nand U718 (N_718,In_653,In_240);
nand U719 (N_719,N_451,N_80);
or U720 (N_720,In_385,In_1494);
or U721 (N_721,N_196,In_1132);
xor U722 (N_722,N_14,In_1044);
nor U723 (N_723,N_401,In_1400);
or U724 (N_724,N_145,In_1023);
and U725 (N_725,In_76,In_686);
xor U726 (N_726,In_193,In_725);
nand U727 (N_727,In_1267,In_306);
nand U728 (N_728,N_144,N_107);
xor U729 (N_729,N_353,In_1380);
xnor U730 (N_730,In_140,N_41);
xor U731 (N_731,In_1230,In_665);
nor U732 (N_732,N_195,N_172);
nor U733 (N_733,In_820,N_198);
xnor U734 (N_734,N_466,N_342);
xor U735 (N_735,In_271,In_865);
and U736 (N_736,N_440,In_1204);
nand U737 (N_737,In_155,N_223);
nor U738 (N_738,In_1239,N_361);
and U739 (N_739,In_635,In_742);
nor U740 (N_740,N_218,In_568);
nor U741 (N_741,In_126,N_136);
and U742 (N_742,In_897,In_1131);
or U743 (N_743,In_629,N_420);
and U744 (N_744,In_808,N_8);
nand U745 (N_745,N_357,In_606);
nand U746 (N_746,In_873,In_543);
nor U747 (N_747,In_119,N_17);
nor U748 (N_748,N_139,In_391);
xnor U749 (N_749,In_939,In_1481);
or U750 (N_750,N_344,In_503);
nand U751 (N_751,N_275,In_668);
nor U752 (N_752,N_33,N_121);
nand U753 (N_753,N_40,In_601);
or U754 (N_754,N_161,In_451);
nor U755 (N_755,In_602,N_25);
nand U756 (N_756,In_181,In_853);
and U757 (N_757,N_280,N_266);
nand U758 (N_758,N_368,In_1284);
and U759 (N_759,N_351,In_1405);
xor U760 (N_760,In_347,N_94);
nor U761 (N_761,N_138,N_250);
nor U762 (N_762,In_426,N_170);
xnor U763 (N_763,In_105,N_406);
nand U764 (N_764,In_690,N_229);
xor U765 (N_765,N_44,In_234);
or U766 (N_766,In_49,N_336);
nand U767 (N_767,N_109,In_569);
and U768 (N_768,N_207,N_392);
and U769 (N_769,In_513,N_365);
nand U770 (N_770,N_370,In_425);
xor U771 (N_771,N_264,N_115);
or U772 (N_772,In_1445,N_399);
nor U773 (N_773,In_1016,In_1241);
or U774 (N_774,N_2,N_470);
nand U775 (N_775,In_465,In_1171);
nor U776 (N_776,In_250,N_456);
xor U777 (N_777,In_6,N_253);
nand U778 (N_778,In_1046,N_329);
nor U779 (N_779,N_350,N_477);
nand U780 (N_780,N_364,N_426);
nor U781 (N_781,In_1232,N_70);
or U782 (N_782,In_436,In_471);
nand U783 (N_783,In_1243,N_430);
nor U784 (N_784,In_226,N_320);
and U785 (N_785,N_117,N_460);
nand U786 (N_786,N_54,In_162);
or U787 (N_787,In_764,In_55);
and U788 (N_788,N_308,In_109);
nand U789 (N_789,N_120,N_382);
nor U790 (N_790,N_492,N_232);
and U791 (N_791,N_471,N_91);
nand U792 (N_792,N_408,N_455);
xnor U793 (N_793,N_428,N_119);
nand U794 (N_794,N_108,In_1248);
nand U795 (N_795,N_18,N_255);
nor U796 (N_796,N_434,In_1421);
xnor U797 (N_797,N_281,N_114);
xnor U798 (N_798,N_65,In_1133);
xnor U799 (N_799,N_163,N_50);
xnor U800 (N_800,In_128,In_1499);
nor U801 (N_801,N_390,N_152);
or U802 (N_802,In_396,In_1235);
nor U803 (N_803,In_1331,In_1350);
nand U804 (N_804,In_467,N_43);
nand U805 (N_805,N_433,N_431);
and U806 (N_806,N_289,In_1275);
xor U807 (N_807,N_437,In_607);
xnor U808 (N_808,In_976,In_800);
or U809 (N_809,In_1128,In_1370);
and U810 (N_810,In_315,In_1321);
and U811 (N_811,N_257,N_427);
or U812 (N_812,N_374,In_745);
nor U813 (N_813,In_687,In_1448);
or U814 (N_814,In_1392,N_61);
or U815 (N_815,N_270,In_1052);
and U816 (N_816,In_1320,In_1374);
nor U817 (N_817,N_221,N_131);
xor U818 (N_818,N_189,N_441);
xnor U819 (N_819,N_447,N_6);
xnor U820 (N_820,In_979,In_681);
nor U821 (N_821,In_58,N_269);
xnor U822 (N_822,In_357,In_151);
nor U823 (N_823,In_48,N_343);
xnor U824 (N_824,N_205,In_239);
nor U825 (N_825,N_154,N_35);
xor U826 (N_826,N_331,N_465);
nor U827 (N_827,In_505,In_1381);
and U828 (N_828,N_104,N_450);
and U829 (N_829,N_153,N_132);
nand U830 (N_830,In_1233,N_110);
nor U831 (N_831,N_274,In_932);
nor U832 (N_832,N_267,In_743);
and U833 (N_833,N_254,In_1142);
nand U834 (N_834,In_631,N_453);
nand U835 (N_835,In_1282,N_238);
nor U836 (N_836,In_1049,N_340);
nor U837 (N_837,N_45,In_1136);
nand U838 (N_838,In_1120,In_713);
xor U839 (N_839,N_99,N_160);
xnor U840 (N_840,In_835,N_417);
nor U841 (N_841,N_230,N_359);
nor U842 (N_842,N_11,In_484);
or U843 (N_843,N_90,N_300);
nor U844 (N_844,In_359,In_512);
nand U845 (N_845,In_1300,In_501);
or U846 (N_846,In_754,N_226);
nand U847 (N_847,In_1299,N_425);
nor U848 (N_848,In_314,In_439);
nor U849 (N_849,In_1211,N_52);
or U850 (N_850,In_1095,In_401);
and U851 (N_851,N_98,In_511);
nor U852 (N_852,N_166,N_322);
and U853 (N_853,N_12,N_246);
nand U854 (N_854,N_244,In_656);
nor U855 (N_855,N_247,N_293);
nand U856 (N_856,In_594,N_313);
or U857 (N_857,N_56,N_348);
and U858 (N_858,N_489,N_432);
and U859 (N_859,N_77,In_1444);
and U860 (N_860,In_617,N_265);
and U861 (N_861,In_715,In_1124);
nor U862 (N_862,N_422,N_150);
or U863 (N_863,N_9,In_481);
xor U864 (N_864,N_7,In_100);
nor U865 (N_865,N_277,N_448);
xnor U866 (N_866,In_1051,N_38);
nand U867 (N_867,In_256,N_240);
nor U868 (N_868,In_831,N_95);
xor U869 (N_869,N_415,In_121);
and U870 (N_870,In_1287,In_986);
or U871 (N_871,N_413,In_680);
and U872 (N_872,In_261,In_166);
xor U873 (N_873,In_1411,In_145);
and U874 (N_874,N_381,In_257);
and U875 (N_875,N_179,In_422);
nand U876 (N_876,N_317,N_200);
nor U877 (N_877,N_366,In_1177);
nand U878 (N_878,N_463,In_427);
xor U879 (N_879,In_102,N_478);
or U880 (N_880,N_272,N_375);
nor U881 (N_881,In_753,N_235);
nor U882 (N_882,N_133,In_324);
and U883 (N_883,In_1480,In_282);
or U884 (N_884,In_1061,In_755);
nand U885 (N_885,In_863,N_127);
xnor U886 (N_886,In_998,N_122);
nor U887 (N_887,In_888,In_209);
or U888 (N_888,N_358,In_1121);
nor U889 (N_889,N_241,In_517);
or U890 (N_890,In_1394,In_643);
or U891 (N_891,In_169,In_790);
nand U892 (N_892,In_1399,N_335);
nor U893 (N_893,In_206,In_1268);
or U894 (N_894,In_1413,N_208);
nand U895 (N_895,N_30,In_843);
nand U896 (N_896,N_330,In_1144);
nand U897 (N_897,N_341,N_102);
nand U898 (N_898,N_217,N_346);
and U899 (N_899,In_1059,N_314);
xnor U900 (N_900,N_414,In_699);
nand U901 (N_901,In_563,N_36);
nor U902 (N_902,In_525,N_310);
nand U903 (N_903,In_461,N_316);
nor U904 (N_904,N_185,In_251);
nor U905 (N_905,N_21,In_836);
and U906 (N_906,In_666,In_1041);
or U907 (N_907,In_303,In_253);
nor U908 (N_908,N_258,In_1288);
and U909 (N_909,N_338,N_187);
nor U910 (N_910,N_58,In_1362);
and U911 (N_911,In_519,N_385);
and U912 (N_912,N_124,In_874);
nor U913 (N_913,In_1102,N_268);
or U914 (N_914,N_362,In_1492);
nor U915 (N_915,In_968,In_469);
and U916 (N_916,N_356,In_540);
and U917 (N_917,In_1014,In_1162);
nor U918 (N_918,N_28,N_296);
nor U919 (N_919,N_112,N_88);
nand U920 (N_920,In_403,In_129);
and U921 (N_921,In_267,In_136);
nand U922 (N_922,In_995,N_42);
xor U923 (N_923,N_302,N_164);
or U924 (N_924,In_868,N_213);
nor U925 (N_925,N_398,N_387);
or U926 (N_926,In_485,N_135);
and U927 (N_927,N_203,In_473);
or U928 (N_928,In_86,In_462);
nor U929 (N_929,N_394,N_26);
and U930 (N_930,N_3,N_216);
nor U931 (N_931,N_237,In_1247);
or U932 (N_932,N_476,N_352);
nand U933 (N_933,In_705,In_300);
or U934 (N_934,N_418,N_222);
xor U935 (N_935,In_1266,N_339);
and U936 (N_936,In_32,N_412);
xnor U937 (N_937,In_19,In_262);
nand U938 (N_938,In_996,In_1498);
xor U939 (N_939,In_847,N_486);
or U940 (N_940,In_1054,In_224);
or U941 (N_941,In_276,N_311);
nand U942 (N_942,In_640,N_22);
nor U943 (N_943,N_474,In_1115);
nand U944 (N_944,N_424,In_593);
nand U945 (N_945,In_320,N_242);
and U946 (N_946,N_37,N_383);
xor U947 (N_947,In_244,N_176);
nor U948 (N_948,N_19,In_1368);
or U949 (N_949,In_1417,N_349);
and U950 (N_950,N_192,In_634);
nor U951 (N_951,N_252,N_233);
xor U952 (N_952,In_899,In_127);
and U953 (N_953,In_386,N_72);
nand U954 (N_954,In_1351,N_347);
nand U955 (N_955,In_442,In_777);
or U956 (N_956,In_751,In_967);
nand U957 (N_957,In_780,In_506);
and U958 (N_958,In_1100,N_251);
nor U959 (N_959,In_1225,In_516);
nor U960 (N_960,In_809,N_193);
or U961 (N_961,In_1475,N_263);
nor U962 (N_962,N_39,N_156);
or U963 (N_963,In_191,In_1271);
nand U964 (N_964,In_1389,N_327);
nor U965 (N_965,N_74,N_137);
xor U966 (N_966,In_290,N_129);
or U967 (N_967,N_126,N_388);
xnor U968 (N_968,N_367,N_60);
nor U969 (N_969,N_400,In_1024);
nand U970 (N_970,In_1213,N_142);
or U971 (N_971,N_148,In_333);
xnor U972 (N_972,In_390,In_542);
and U973 (N_973,N_146,In_24);
and U974 (N_974,In_474,In_732);
or U975 (N_975,In_36,In_721);
xor U976 (N_976,In_337,N_97);
or U977 (N_977,N_495,In_106);
nand U978 (N_978,N_282,In_1450);
nor U979 (N_979,In_882,N_429);
nor U980 (N_980,In_1081,In_172);
nand U981 (N_981,N_354,N_443);
xnor U982 (N_982,N_92,In_57);
nand U983 (N_983,N_84,In_706);
xor U984 (N_984,In_1189,N_480);
nor U985 (N_985,In_164,N_326);
nand U986 (N_986,In_170,In_302);
nand U987 (N_987,N_287,In_702);
nand U988 (N_988,N_228,In_960);
and U989 (N_989,N_419,N_4);
xor U990 (N_990,In_817,N_190);
nand U991 (N_991,N_83,In_405);
xor U992 (N_992,N_96,N_485);
and U993 (N_993,N_371,N_334);
nor U994 (N_994,In_1003,In_195);
nor U995 (N_995,In_621,N_245);
nor U996 (N_996,In_1147,N_393);
or U997 (N_997,N_304,In_165);
and U998 (N_998,In_1319,N_206);
nor U999 (N_999,N_236,N_82);
xnor U1000 (N_1000,N_963,N_841);
or U1001 (N_1001,N_915,N_891);
nor U1002 (N_1002,N_560,N_702);
xnor U1003 (N_1003,N_661,N_708);
or U1004 (N_1004,N_548,N_959);
xnor U1005 (N_1005,N_730,N_558);
xnor U1006 (N_1006,N_551,N_636);
nor U1007 (N_1007,N_545,N_852);
nand U1008 (N_1008,N_534,N_678);
nand U1009 (N_1009,N_821,N_918);
or U1010 (N_1010,N_921,N_693);
xnor U1011 (N_1011,N_904,N_872);
and U1012 (N_1012,N_553,N_762);
nand U1013 (N_1013,N_979,N_931);
or U1014 (N_1014,N_945,N_562);
nand U1015 (N_1015,N_621,N_700);
and U1016 (N_1016,N_801,N_861);
and U1017 (N_1017,N_863,N_719);
and U1018 (N_1018,N_751,N_660);
xor U1019 (N_1019,N_817,N_576);
nor U1020 (N_1020,N_758,N_722);
nand U1021 (N_1021,N_855,N_783);
or U1022 (N_1022,N_639,N_640);
xor U1023 (N_1023,N_528,N_793);
nor U1024 (N_1024,N_772,N_582);
nor U1025 (N_1025,N_713,N_820);
nor U1026 (N_1026,N_780,N_992);
and U1027 (N_1027,N_644,N_657);
nor U1028 (N_1028,N_724,N_687);
or U1029 (N_1029,N_973,N_796);
nor U1030 (N_1030,N_508,N_927);
and U1031 (N_1031,N_543,N_969);
nor U1032 (N_1032,N_716,N_692);
or U1033 (N_1033,N_857,N_658);
or U1034 (N_1034,N_734,N_706);
nand U1035 (N_1035,N_526,N_961);
xnor U1036 (N_1036,N_810,N_981);
and U1037 (N_1037,N_802,N_809);
and U1038 (N_1038,N_889,N_769);
nand U1039 (N_1039,N_797,N_847);
and U1040 (N_1040,N_749,N_711);
and U1041 (N_1041,N_954,N_837);
xor U1042 (N_1042,N_926,N_928);
xnor U1043 (N_1043,N_903,N_570);
nor U1044 (N_1044,N_788,N_890);
or U1045 (N_1045,N_691,N_873);
nand U1046 (N_1046,N_947,N_836);
or U1047 (N_1047,N_964,N_659);
nor U1048 (N_1048,N_573,N_698);
nand U1049 (N_1049,N_624,N_625);
nand U1050 (N_1050,N_830,N_760);
or U1051 (N_1051,N_675,N_842);
nand U1052 (N_1052,N_977,N_906);
and U1053 (N_1053,N_853,N_643);
and U1054 (N_1054,N_787,N_631);
xor U1055 (N_1055,N_613,N_627);
nand U1056 (N_1056,N_934,N_984);
or U1057 (N_1057,N_633,N_816);
or U1058 (N_1058,N_666,N_667);
or U1059 (N_1059,N_759,N_888);
xnor U1060 (N_1060,N_727,N_533);
and U1061 (N_1061,N_912,N_745);
nor U1062 (N_1062,N_506,N_884);
or U1063 (N_1063,N_744,N_850);
nand U1064 (N_1064,N_507,N_768);
xor U1065 (N_1065,N_606,N_647);
or U1066 (N_1066,N_930,N_846);
or U1067 (N_1067,N_944,N_999);
nand U1068 (N_1068,N_909,N_567);
xnor U1069 (N_1069,N_808,N_572);
and U1070 (N_1070,N_653,N_747);
nand U1071 (N_1071,N_529,N_843);
nand U1072 (N_1072,N_579,N_822);
or U1073 (N_1073,N_940,N_826);
and U1074 (N_1074,N_645,N_869);
nand U1075 (N_1075,N_900,N_654);
nor U1076 (N_1076,N_806,N_602);
xor U1077 (N_1077,N_733,N_557);
xor U1078 (N_1078,N_723,N_831);
and U1079 (N_1079,N_587,N_868);
nand U1080 (N_1080,N_514,N_752);
nand U1081 (N_1081,N_967,N_677);
nand U1082 (N_1082,N_513,N_886);
and U1083 (N_1083,N_575,N_592);
and U1084 (N_1084,N_966,N_717);
and U1085 (N_1085,N_544,N_935);
and U1086 (N_1086,N_845,N_766);
xnor U1087 (N_1087,N_581,N_585);
nand U1088 (N_1088,N_971,N_827);
nor U1089 (N_1089,N_811,N_595);
or U1090 (N_1090,N_807,N_916);
xnor U1091 (N_1091,N_630,N_518);
and U1092 (N_1092,N_804,N_763);
xor U1093 (N_1093,N_538,N_832);
xor U1094 (N_1094,N_781,N_799);
or U1095 (N_1095,N_858,N_829);
and U1096 (N_1096,N_883,N_565);
or U1097 (N_1097,N_583,N_569);
xnor U1098 (N_1098,N_870,N_597);
nand U1099 (N_1099,N_591,N_761);
xor U1100 (N_1100,N_665,N_834);
nand U1101 (N_1101,N_958,N_955);
nor U1102 (N_1102,N_839,N_782);
or U1103 (N_1103,N_814,N_878);
or U1104 (N_1104,N_974,N_705);
nand U1105 (N_1105,N_532,N_683);
xnor U1106 (N_1106,N_509,N_785);
and U1107 (N_1107,N_892,N_527);
and U1108 (N_1108,N_756,N_738);
and U1109 (N_1109,N_957,N_860);
nand U1110 (N_1110,N_925,N_689);
xor U1111 (N_1111,N_978,N_995);
nor U1112 (N_1112,N_688,N_972);
xnor U1113 (N_1113,N_965,N_594);
nor U1114 (N_1114,N_503,N_901);
and U1115 (N_1115,N_662,N_523);
and U1116 (N_1116,N_776,N_684);
or U1117 (N_1117,N_517,N_616);
nor U1118 (N_1118,N_881,N_764);
xnor U1119 (N_1119,N_571,N_701);
and U1120 (N_1120,N_755,N_652);
nor U1121 (N_1121,N_664,N_704);
nand U1122 (N_1122,N_976,N_985);
nor U1123 (N_1123,N_501,N_771);
xor U1124 (N_1124,N_608,N_859);
nand U1125 (N_1125,N_651,N_598);
xor U1126 (N_1126,N_586,N_628);
and U1127 (N_1127,N_865,N_670);
or U1128 (N_1128,N_867,N_686);
and U1129 (N_1129,N_894,N_770);
nand U1130 (N_1130,N_696,N_531);
xor U1131 (N_1131,N_779,N_993);
and U1132 (N_1132,N_611,N_709);
xor U1133 (N_1133,N_521,N_962);
xor U1134 (N_1134,N_599,N_986);
nor U1135 (N_1135,N_735,N_540);
xor U1136 (N_1136,N_753,N_897);
or U1137 (N_1137,N_646,N_946);
nand U1138 (N_1138,N_968,N_876);
xor U1139 (N_1139,N_874,N_911);
nor U1140 (N_1140,N_823,N_511);
or U1141 (N_1141,N_980,N_987);
xnor U1142 (N_1142,N_714,N_712);
nor U1143 (N_1143,N_694,N_690);
and U1144 (N_1144,N_546,N_838);
nor U1145 (N_1145,N_556,N_710);
nor U1146 (N_1146,N_564,N_748);
or U1147 (N_1147,N_536,N_637);
nand U1148 (N_1148,N_933,N_794);
and U1149 (N_1149,N_924,N_610);
and U1150 (N_1150,N_887,N_603);
nor U1151 (N_1151,N_798,N_680);
or U1152 (N_1152,N_619,N_877);
and U1153 (N_1153,N_996,N_988);
xor U1154 (N_1154,N_939,N_648);
or U1155 (N_1155,N_784,N_975);
nand U1156 (N_1156,N_584,N_673);
and U1157 (N_1157,N_994,N_685);
and U1158 (N_1158,N_908,N_697);
nand U1159 (N_1159,N_537,N_866);
nor U1160 (N_1160,N_917,N_668);
and U1161 (N_1161,N_590,N_559);
and U1162 (N_1162,N_525,N_656);
nor U1163 (N_1163,N_905,N_910);
and U1164 (N_1164,N_505,N_504);
xor U1165 (N_1165,N_681,N_754);
nand U1166 (N_1166,N_825,N_638);
nor U1167 (N_1167,N_746,N_805);
and U1168 (N_1168,N_948,N_737);
nor U1169 (N_1169,N_923,N_998);
and U1170 (N_1170,N_672,N_561);
nor U1171 (N_1171,N_813,N_600);
and U1172 (N_1172,N_615,N_726);
or U1173 (N_1173,N_899,N_535);
nor U1174 (N_1174,N_942,N_932);
nand U1175 (N_1175,N_844,N_898);
xor U1176 (N_1176,N_835,N_626);
nor U1177 (N_1177,N_541,N_703);
and U1178 (N_1178,N_902,N_642);
nor U1179 (N_1179,N_552,N_907);
nand U1180 (N_1180,N_729,N_914);
nand U1181 (N_1181,N_563,N_520);
or U1182 (N_1182,N_718,N_663);
or U1183 (N_1183,N_767,N_919);
or U1184 (N_1184,N_893,N_943);
or U1185 (N_1185,N_812,N_549);
or U1186 (N_1186,N_851,N_913);
nand U1187 (N_1187,N_676,N_707);
or U1188 (N_1188,N_815,N_765);
and U1189 (N_1189,N_609,N_941);
or U1190 (N_1190,N_792,N_715);
or U1191 (N_1191,N_922,N_588);
xor U1192 (N_1192,N_953,N_635);
nand U1193 (N_1193,N_936,N_773);
nand U1194 (N_1194,N_989,N_790);
xnor U1195 (N_1195,N_596,N_632);
nor U1196 (N_1196,N_856,N_728);
nand U1197 (N_1197,N_824,N_896);
nor U1198 (N_1198,N_818,N_990);
or U1199 (N_1199,N_510,N_671);
nand U1200 (N_1200,N_566,N_828);
nand U1201 (N_1201,N_614,N_929);
xor U1202 (N_1202,N_519,N_871);
xor U1203 (N_1203,N_864,N_885);
or U1204 (N_1204,N_550,N_956);
xnor U1205 (N_1205,N_840,N_634);
or U1206 (N_1206,N_970,N_778);
nand U1207 (N_1207,N_516,N_741);
and U1208 (N_1208,N_951,N_952);
xnor U1209 (N_1209,N_791,N_695);
nand U1210 (N_1210,N_522,N_895);
or U1211 (N_1211,N_542,N_669);
and U1212 (N_1212,N_512,N_607);
or U1213 (N_1213,N_622,N_750);
or U1214 (N_1214,N_879,N_736);
and U1215 (N_1215,N_547,N_612);
xnor U1216 (N_1216,N_795,N_502);
or U1217 (N_1217,N_555,N_880);
or U1218 (N_1218,N_739,N_740);
xnor U1219 (N_1219,N_997,N_774);
or U1220 (N_1220,N_530,N_983);
and U1221 (N_1221,N_649,N_568);
nor U1222 (N_1222,N_777,N_775);
nor U1223 (N_1223,N_500,N_854);
and U1224 (N_1224,N_757,N_589);
xnor U1225 (N_1225,N_991,N_515);
and U1226 (N_1226,N_650,N_604);
nand U1227 (N_1227,N_731,N_849);
or U1228 (N_1228,N_641,N_819);
and U1229 (N_1229,N_524,N_960);
nor U1230 (N_1230,N_580,N_800);
nand U1231 (N_1231,N_833,N_786);
or U1232 (N_1232,N_682,N_950);
xnor U1233 (N_1233,N_938,N_655);
or U1234 (N_1234,N_617,N_574);
xor U1235 (N_1235,N_618,N_620);
nand U1236 (N_1236,N_721,N_743);
or U1237 (N_1237,N_742,N_593);
nand U1238 (N_1238,N_982,N_920);
or U1239 (N_1239,N_937,N_949);
nand U1240 (N_1240,N_789,N_679);
and U1241 (N_1241,N_554,N_629);
nor U1242 (N_1242,N_848,N_699);
nand U1243 (N_1243,N_803,N_882);
nor U1244 (N_1244,N_674,N_875);
nand U1245 (N_1245,N_725,N_605);
nor U1246 (N_1246,N_720,N_577);
and U1247 (N_1247,N_539,N_623);
or U1248 (N_1248,N_862,N_732);
xor U1249 (N_1249,N_578,N_601);
or U1250 (N_1250,N_532,N_600);
nor U1251 (N_1251,N_885,N_670);
or U1252 (N_1252,N_610,N_775);
or U1253 (N_1253,N_814,N_887);
or U1254 (N_1254,N_676,N_784);
or U1255 (N_1255,N_760,N_821);
nand U1256 (N_1256,N_992,N_546);
nor U1257 (N_1257,N_864,N_866);
and U1258 (N_1258,N_596,N_940);
nor U1259 (N_1259,N_944,N_597);
nor U1260 (N_1260,N_503,N_668);
and U1261 (N_1261,N_834,N_632);
xor U1262 (N_1262,N_901,N_944);
xnor U1263 (N_1263,N_652,N_575);
or U1264 (N_1264,N_725,N_864);
nor U1265 (N_1265,N_622,N_623);
xor U1266 (N_1266,N_824,N_702);
nor U1267 (N_1267,N_867,N_818);
or U1268 (N_1268,N_545,N_794);
and U1269 (N_1269,N_601,N_723);
xnor U1270 (N_1270,N_908,N_536);
xnor U1271 (N_1271,N_842,N_507);
or U1272 (N_1272,N_693,N_939);
or U1273 (N_1273,N_937,N_943);
nor U1274 (N_1274,N_799,N_555);
nand U1275 (N_1275,N_914,N_778);
nor U1276 (N_1276,N_802,N_856);
nor U1277 (N_1277,N_950,N_931);
nor U1278 (N_1278,N_671,N_765);
nor U1279 (N_1279,N_911,N_902);
nor U1280 (N_1280,N_597,N_568);
and U1281 (N_1281,N_504,N_617);
nand U1282 (N_1282,N_796,N_752);
or U1283 (N_1283,N_632,N_715);
and U1284 (N_1284,N_867,N_906);
nor U1285 (N_1285,N_934,N_918);
nor U1286 (N_1286,N_944,N_502);
and U1287 (N_1287,N_686,N_912);
xor U1288 (N_1288,N_605,N_878);
xnor U1289 (N_1289,N_555,N_921);
nand U1290 (N_1290,N_571,N_607);
nand U1291 (N_1291,N_927,N_614);
nor U1292 (N_1292,N_693,N_915);
or U1293 (N_1293,N_786,N_855);
and U1294 (N_1294,N_837,N_535);
nor U1295 (N_1295,N_520,N_598);
xor U1296 (N_1296,N_887,N_669);
nand U1297 (N_1297,N_943,N_618);
xor U1298 (N_1298,N_854,N_800);
or U1299 (N_1299,N_921,N_955);
xnor U1300 (N_1300,N_661,N_700);
nor U1301 (N_1301,N_997,N_582);
xnor U1302 (N_1302,N_791,N_804);
xor U1303 (N_1303,N_793,N_805);
nor U1304 (N_1304,N_992,N_756);
or U1305 (N_1305,N_703,N_770);
and U1306 (N_1306,N_856,N_557);
and U1307 (N_1307,N_746,N_955);
nand U1308 (N_1308,N_907,N_674);
and U1309 (N_1309,N_839,N_675);
or U1310 (N_1310,N_648,N_823);
nand U1311 (N_1311,N_625,N_998);
and U1312 (N_1312,N_873,N_666);
or U1313 (N_1313,N_630,N_728);
and U1314 (N_1314,N_565,N_542);
nor U1315 (N_1315,N_848,N_548);
nor U1316 (N_1316,N_830,N_698);
and U1317 (N_1317,N_637,N_938);
or U1318 (N_1318,N_824,N_628);
and U1319 (N_1319,N_597,N_918);
xor U1320 (N_1320,N_880,N_619);
nand U1321 (N_1321,N_641,N_960);
nor U1322 (N_1322,N_876,N_931);
nor U1323 (N_1323,N_835,N_719);
and U1324 (N_1324,N_852,N_814);
and U1325 (N_1325,N_575,N_508);
xor U1326 (N_1326,N_529,N_722);
nand U1327 (N_1327,N_507,N_717);
nand U1328 (N_1328,N_714,N_601);
and U1329 (N_1329,N_803,N_924);
xor U1330 (N_1330,N_556,N_582);
or U1331 (N_1331,N_627,N_823);
nand U1332 (N_1332,N_553,N_747);
nand U1333 (N_1333,N_737,N_856);
or U1334 (N_1334,N_834,N_694);
nor U1335 (N_1335,N_552,N_909);
nand U1336 (N_1336,N_730,N_743);
xor U1337 (N_1337,N_976,N_851);
nor U1338 (N_1338,N_829,N_677);
nor U1339 (N_1339,N_903,N_901);
xnor U1340 (N_1340,N_706,N_989);
xor U1341 (N_1341,N_999,N_755);
or U1342 (N_1342,N_575,N_907);
xor U1343 (N_1343,N_554,N_885);
nor U1344 (N_1344,N_548,N_505);
xnor U1345 (N_1345,N_721,N_659);
xor U1346 (N_1346,N_814,N_796);
xor U1347 (N_1347,N_913,N_582);
nor U1348 (N_1348,N_837,N_963);
and U1349 (N_1349,N_963,N_746);
or U1350 (N_1350,N_742,N_928);
and U1351 (N_1351,N_847,N_913);
or U1352 (N_1352,N_768,N_504);
and U1353 (N_1353,N_533,N_934);
or U1354 (N_1354,N_713,N_903);
nor U1355 (N_1355,N_700,N_674);
nor U1356 (N_1356,N_613,N_897);
xnor U1357 (N_1357,N_707,N_866);
and U1358 (N_1358,N_749,N_775);
or U1359 (N_1359,N_889,N_551);
xor U1360 (N_1360,N_819,N_812);
or U1361 (N_1361,N_571,N_992);
nand U1362 (N_1362,N_688,N_915);
xor U1363 (N_1363,N_803,N_752);
or U1364 (N_1364,N_568,N_636);
nor U1365 (N_1365,N_540,N_697);
xor U1366 (N_1366,N_523,N_729);
nor U1367 (N_1367,N_514,N_627);
nor U1368 (N_1368,N_815,N_802);
nor U1369 (N_1369,N_554,N_827);
and U1370 (N_1370,N_594,N_976);
nor U1371 (N_1371,N_546,N_870);
nor U1372 (N_1372,N_797,N_521);
xnor U1373 (N_1373,N_743,N_578);
or U1374 (N_1374,N_928,N_850);
and U1375 (N_1375,N_871,N_862);
and U1376 (N_1376,N_594,N_572);
nand U1377 (N_1377,N_617,N_762);
and U1378 (N_1378,N_746,N_572);
nand U1379 (N_1379,N_956,N_650);
or U1380 (N_1380,N_909,N_751);
nand U1381 (N_1381,N_607,N_773);
or U1382 (N_1382,N_904,N_697);
or U1383 (N_1383,N_730,N_899);
and U1384 (N_1384,N_532,N_755);
and U1385 (N_1385,N_652,N_903);
or U1386 (N_1386,N_803,N_616);
nand U1387 (N_1387,N_610,N_664);
nor U1388 (N_1388,N_950,N_872);
nand U1389 (N_1389,N_827,N_869);
nor U1390 (N_1390,N_953,N_750);
or U1391 (N_1391,N_725,N_718);
and U1392 (N_1392,N_569,N_840);
xor U1393 (N_1393,N_863,N_595);
and U1394 (N_1394,N_753,N_761);
xor U1395 (N_1395,N_655,N_826);
nor U1396 (N_1396,N_513,N_651);
nand U1397 (N_1397,N_697,N_634);
nand U1398 (N_1398,N_667,N_509);
nor U1399 (N_1399,N_681,N_833);
xnor U1400 (N_1400,N_529,N_814);
xnor U1401 (N_1401,N_682,N_742);
nand U1402 (N_1402,N_693,N_948);
and U1403 (N_1403,N_779,N_799);
nor U1404 (N_1404,N_586,N_803);
nand U1405 (N_1405,N_997,N_789);
nor U1406 (N_1406,N_983,N_936);
or U1407 (N_1407,N_561,N_941);
nand U1408 (N_1408,N_666,N_779);
nor U1409 (N_1409,N_588,N_635);
or U1410 (N_1410,N_857,N_817);
nand U1411 (N_1411,N_827,N_908);
nand U1412 (N_1412,N_987,N_817);
nor U1413 (N_1413,N_829,N_847);
nor U1414 (N_1414,N_952,N_515);
and U1415 (N_1415,N_965,N_604);
xnor U1416 (N_1416,N_746,N_574);
or U1417 (N_1417,N_836,N_800);
xor U1418 (N_1418,N_506,N_504);
nand U1419 (N_1419,N_791,N_923);
or U1420 (N_1420,N_524,N_836);
nand U1421 (N_1421,N_832,N_978);
xnor U1422 (N_1422,N_538,N_889);
and U1423 (N_1423,N_779,N_883);
or U1424 (N_1424,N_928,N_919);
nor U1425 (N_1425,N_886,N_665);
nand U1426 (N_1426,N_866,N_995);
xnor U1427 (N_1427,N_798,N_871);
nor U1428 (N_1428,N_511,N_555);
xnor U1429 (N_1429,N_521,N_968);
and U1430 (N_1430,N_773,N_669);
nand U1431 (N_1431,N_799,N_994);
nor U1432 (N_1432,N_910,N_929);
nand U1433 (N_1433,N_735,N_698);
or U1434 (N_1434,N_762,N_515);
nor U1435 (N_1435,N_622,N_503);
nand U1436 (N_1436,N_895,N_583);
and U1437 (N_1437,N_937,N_676);
and U1438 (N_1438,N_992,N_634);
or U1439 (N_1439,N_769,N_672);
or U1440 (N_1440,N_621,N_869);
xnor U1441 (N_1441,N_666,N_526);
xnor U1442 (N_1442,N_941,N_890);
xnor U1443 (N_1443,N_777,N_684);
nand U1444 (N_1444,N_776,N_575);
and U1445 (N_1445,N_683,N_655);
or U1446 (N_1446,N_916,N_668);
nor U1447 (N_1447,N_977,N_926);
or U1448 (N_1448,N_827,N_754);
and U1449 (N_1449,N_909,N_743);
xor U1450 (N_1450,N_928,N_715);
and U1451 (N_1451,N_991,N_628);
xnor U1452 (N_1452,N_968,N_552);
nand U1453 (N_1453,N_780,N_760);
or U1454 (N_1454,N_970,N_904);
xnor U1455 (N_1455,N_818,N_748);
and U1456 (N_1456,N_584,N_603);
and U1457 (N_1457,N_795,N_517);
xor U1458 (N_1458,N_894,N_692);
nand U1459 (N_1459,N_892,N_899);
or U1460 (N_1460,N_557,N_891);
xnor U1461 (N_1461,N_500,N_900);
or U1462 (N_1462,N_692,N_978);
or U1463 (N_1463,N_627,N_822);
nand U1464 (N_1464,N_560,N_596);
nor U1465 (N_1465,N_683,N_701);
xnor U1466 (N_1466,N_552,N_640);
and U1467 (N_1467,N_931,N_655);
nor U1468 (N_1468,N_520,N_731);
nor U1469 (N_1469,N_875,N_879);
nor U1470 (N_1470,N_676,N_539);
nand U1471 (N_1471,N_707,N_938);
nor U1472 (N_1472,N_687,N_999);
nand U1473 (N_1473,N_932,N_983);
xor U1474 (N_1474,N_666,N_596);
nand U1475 (N_1475,N_612,N_762);
nor U1476 (N_1476,N_674,N_981);
nor U1477 (N_1477,N_836,N_562);
and U1478 (N_1478,N_931,N_692);
nor U1479 (N_1479,N_639,N_915);
or U1480 (N_1480,N_857,N_599);
nand U1481 (N_1481,N_967,N_602);
nand U1482 (N_1482,N_895,N_652);
xor U1483 (N_1483,N_524,N_730);
nand U1484 (N_1484,N_606,N_517);
and U1485 (N_1485,N_754,N_699);
xor U1486 (N_1486,N_509,N_535);
nand U1487 (N_1487,N_632,N_521);
nand U1488 (N_1488,N_608,N_526);
nor U1489 (N_1489,N_666,N_855);
nand U1490 (N_1490,N_568,N_527);
nor U1491 (N_1491,N_778,N_709);
xor U1492 (N_1492,N_692,N_829);
nor U1493 (N_1493,N_737,N_845);
nor U1494 (N_1494,N_512,N_832);
xor U1495 (N_1495,N_552,N_769);
nor U1496 (N_1496,N_748,N_528);
xor U1497 (N_1497,N_792,N_688);
xor U1498 (N_1498,N_619,N_623);
and U1499 (N_1499,N_523,N_710);
nor U1500 (N_1500,N_1048,N_1174);
nor U1501 (N_1501,N_1030,N_1348);
xnor U1502 (N_1502,N_1419,N_1051);
nand U1503 (N_1503,N_1110,N_1192);
or U1504 (N_1504,N_1295,N_1431);
or U1505 (N_1505,N_1134,N_1376);
xnor U1506 (N_1506,N_1396,N_1077);
or U1507 (N_1507,N_1093,N_1023);
xor U1508 (N_1508,N_1132,N_1316);
and U1509 (N_1509,N_1344,N_1096);
xnor U1510 (N_1510,N_1177,N_1219);
nor U1511 (N_1511,N_1176,N_1355);
and U1512 (N_1512,N_1401,N_1322);
or U1513 (N_1513,N_1411,N_1223);
nor U1514 (N_1514,N_1474,N_1349);
and U1515 (N_1515,N_1080,N_1095);
or U1516 (N_1516,N_1391,N_1189);
nand U1517 (N_1517,N_1392,N_1178);
nor U1518 (N_1518,N_1480,N_1155);
or U1519 (N_1519,N_1338,N_1086);
and U1520 (N_1520,N_1307,N_1124);
or U1521 (N_1521,N_1196,N_1242);
and U1522 (N_1522,N_1033,N_1424);
or U1523 (N_1523,N_1193,N_1246);
or U1524 (N_1524,N_1404,N_1267);
nor U1525 (N_1525,N_1187,N_1430);
or U1526 (N_1526,N_1206,N_1118);
nand U1527 (N_1527,N_1125,N_1087);
xnor U1528 (N_1528,N_1180,N_1388);
or U1529 (N_1529,N_1153,N_1004);
and U1530 (N_1530,N_1014,N_1248);
or U1531 (N_1531,N_1444,N_1166);
or U1532 (N_1532,N_1353,N_1022);
and U1533 (N_1533,N_1390,N_1420);
nor U1534 (N_1534,N_1179,N_1498);
nor U1535 (N_1535,N_1276,N_1243);
xnor U1536 (N_1536,N_1122,N_1136);
and U1537 (N_1537,N_1143,N_1367);
or U1538 (N_1538,N_1101,N_1190);
and U1539 (N_1539,N_1137,N_1212);
or U1540 (N_1540,N_1321,N_1144);
nand U1541 (N_1541,N_1319,N_1207);
nand U1542 (N_1542,N_1294,N_1363);
and U1543 (N_1543,N_1078,N_1071);
nand U1544 (N_1544,N_1462,N_1194);
or U1545 (N_1545,N_1074,N_1170);
or U1546 (N_1546,N_1290,N_1374);
xnor U1547 (N_1547,N_1465,N_1441);
and U1548 (N_1548,N_1335,N_1476);
or U1549 (N_1549,N_1495,N_1262);
or U1550 (N_1550,N_1156,N_1375);
or U1551 (N_1551,N_1050,N_1112);
and U1552 (N_1552,N_1039,N_1247);
and U1553 (N_1553,N_1326,N_1133);
nand U1554 (N_1554,N_1450,N_1043);
nand U1555 (N_1555,N_1020,N_1075);
or U1556 (N_1556,N_1362,N_1198);
xnor U1557 (N_1557,N_1008,N_1052);
nor U1558 (N_1558,N_1415,N_1029);
nor U1559 (N_1559,N_1293,N_1397);
and U1560 (N_1560,N_1257,N_1456);
and U1561 (N_1561,N_1324,N_1005);
nand U1562 (N_1562,N_1461,N_1369);
nor U1563 (N_1563,N_1479,N_1205);
or U1564 (N_1564,N_1309,N_1183);
nor U1565 (N_1565,N_1076,N_1395);
nor U1566 (N_1566,N_1208,N_1073);
or U1567 (N_1567,N_1302,N_1266);
and U1568 (N_1568,N_1100,N_1184);
nand U1569 (N_1569,N_1440,N_1346);
and U1570 (N_1570,N_1454,N_1060);
and U1571 (N_1571,N_1313,N_1280);
nor U1572 (N_1572,N_1241,N_1382);
nor U1573 (N_1573,N_1164,N_1237);
nand U1574 (N_1574,N_1062,N_1064);
xor U1575 (N_1575,N_1378,N_1249);
xor U1576 (N_1576,N_1364,N_1090);
nor U1577 (N_1577,N_1002,N_1473);
and U1578 (N_1578,N_1470,N_1059);
or U1579 (N_1579,N_1109,N_1482);
nor U1580 (N_1580,N_1305,N_1417);
nand U1581 (N_1581,N_1497,N_1046);
xor U1582 (N_1582,N_1055,N_1467);
nor U1583 (N_1583,N_1057,N_1458);
xor U1584 (N_1584,N_1270,N_1412);
or U1585 (N_1585,N_1334,N_1149);
nor U1586 (N_1586,N_1127,N_1306);
nor U1587 (N_1587,N_1494,N_1220);
and U1588 (N_1588,N_1094,N_1373);
xnor U1589 (N_1589,N_1282,N_1105);
or U1590 (N_1590,N_1496,N_1379);
nand U1591 (N_1591,N_1263,N_1332);
and U1592 (N_1592,N_1146,N_1056);
nor U1593 (N_1593,N_1469,N_1017);
or U1594 (N_1594,N_1161,N_1032);
nor U1595 (N_1595,N_1471,N_1477);
xnor U1596 (N_1596,N_1021,N_1227);
nor U1597 (N_1597,N_1359,N_1235);
or U1598 (N_1598,N_1026,N_1010);
or U1599 (N_1599,N_1387,N_1377);
or U1600 (N_1600,N_1492,N_1157);
and U1601 (N_1601,N_1296,N_1162);
nand U1602 (N_1602,N_1366,N_1258);
and U1603 (N_1603,N_1016,N_1277);
nor U1604 (N_1604,N_1013,N_1451);
xor U1605 (N_1605,N_1084,N_1489);
nand U1606 (N_1606,N_1422,N_1082);
or U1607 (N_1607,N_1384,N_1402);
and U1608 (N_1608,N_1434,N_1197);
xnor U1609 (N_1609,N_1141,N_1210);
nand U1610 (N_1610,N_1435,N_1288);
nand U1611 (N_1611,N_1217,N_1209);
xor U1612 (N_1612,N_1152,N_1231);
or U1613 (N_1613,N_1036,N_1218);
nor U1614 (N_1614,N_1314,N_1350);
nand U1615 (N_1615,N_1466,N_1114);
nor U1616 (N_1616,N_1347,N_1195);
and U1617 (N_1617,N_1038,N_1403);
xor U1618 (N_1618,N_1394,N_1345);
nor U1619 (N_1619,N_1460,N_1234);
and U1620 (N_1620,N_1148,N_1203);
or U1621 (N_1621,N_1091,N_1286);
or U1622 (N_1622,N_1233,N_1236);
nand U1623 (N_1623,N_1172,N_1279);
xor U1624 (N_1624,N_1006,N_1045);
xnor U1625 (N_1625,N_1027,N_1040);
xor U1626 (N_1626,N_1323,N_1167);
or U1627 (N_1627,N_1478,N_1447);
or U1628 (N_1628,N_1072,N_1493);
and U1629 (N_1629,N_1371,N_1264);
nand U1630 (N_1630,N_1421,N_1151);
or U1631 (N_1631,N_1214,N_1425);
or U1632 (N_1632,N_1251,N_1418);
and U1633 (N_1633,N_1455,N_1273);
and U1634 (N_1634,N_1000,N_1131);
xor U1635 (N_1635,N_1423,N_1410);
nand U1636 (N_1636,N_1271,N_1191);
nor U1637 (N_1637,N_1464,N_1287);
or U1638 (N_1638,N_1140,N_1486);
nand U1639 (N_1639,N_1330,N_1047);
and U1640 (N_1640,N_1115,N_1119);
nand U1641 (N_1641,N_1452,N_1436);
xnor U1642 (N_1642,N_1188,N_1063);
and U1643 (N_1643,N_1001,N_1199);
nor U1644 (N_1644,N_1413,N_1135);
nand U1645 (N_1645,N_1092,N_1108);
nand U1646 (N_1646,N_1201,N_1230);
nor U1647 (N_1647,N_1386,N_1175);
or U1648 (N_1648,N_1037,N_1240);
nor U1649 (N_1649,N_1031,N_1416);
nor U1650 (N_1650,N_1088,N_1147);
or U1651 (N_1651,N_1304,N_1414);
nand U1652 (N_1652,N_1459,N_1099);
xnor U1653 (N_1653,N_1491,N_1275);
nor U1654 (N_1654,N_1487,N_1303);
nand U1655 (N_1655,N_1224,N_1300);
xor U1656 (N_1656,N_1438,N_1102);
and U1657 (N_1657,N_1216,N_1272);
nand U1658 (N_1658,N_1400,N_1485);
and U1659 (N_1659,N_1238,N_1007);
xnor U1660 (N_1660,N_1009,N_1383);
xnor U1661 (N_1661,N_1292,N_1204);
xor U1662 (N_1662,N_1154,N_1121);
or U1663 (N_1663,N_1284,N_1012);
or U1664 (N_1664,N_1499,N_1185);
or U1665 (N_1665,N_1126,N_1336);
or U1666 (N_1666,N_1483,N_1278);
nor U1667 (N_1667,N_1085,N_1142);
and U1668 (N_1668,N_1299,N_1318);
or U1669 (N_1669,N_1213,N_1281);
nor U1670 (N_1670,N_1357,N_1439);
nor U1671 (N_1671,N_1221,N_1361);
and U1672 (N_1672,N_1065,N_1405);
nand U1673 (N_1673,N_1200,N_1352);
nand U1674 (N_1674,N_1106,N_1381);
xor U1675 (N_1675,N_1182,N_1232);
nand U1676 (N_1676,N_1310,N_1222);
nor U1677 (N_1677,N_1261,N_1067);
and U1678 (N_1678,N_1173,N_1340);
or U1679 (N_1679,N_1442,N_1331);
nor U1680 (N_1680,N_1445,N_1358);
nor U1681 (N_1681,N_1116,N_1446);
or U1682 (N_1682,N_1488,N_1228);
and U1683 (N_1683,N_1372,N_1035);
nand U1684 (N_1684,N_1297,N_1186);
nand U1685 (N_1685,N_1432,N_1245);
xnor U1686 (N_1686,N_1490,N_1239);
and U1687 (N_1687,N_1069,N_1229);
nor U1688 (N_1688,N_1111,N_1448);
nor U1689 (N_1689,N_1370,N_1327);
nor U1690 (N_1690,N_1393,N_1259);
nor U1691 (N_1691,N_1068,N_1408);
xnor U1692 (N_1692,N_1308,N_1165);
nand U1693 (N_1693,N_1160,N_1107);
nor U1694 (N_1694,N_1312,N_1070);
nand U1695 (N_1695,N_1254,N_1181);
nand U1696 (N_1696,N_1311,N_1024);
xnor U1697 (N_1697,N_1163,N_1315);
or U1698 (N_1698,N_1484,N_1342);
nor U1699 (N_1699,N_1274,N_1368);
and U1700 (N_1700,N_1406,N_1252);
xnor U1701 (N_1701,N_1468,N_1003);
or U1702 (N_1702,N_1356,N_1171);
and U1703 (N_1703,N_1089,N_1320);
nand U1704 (N_1704,N_1301,N_1283);
nand U1705 (N_1705,N_1018,N_1129);
nand U1706 (N_1706,N_1042,N_1011);
or U1707 (N_1707,N_1225,N_1341);
nor U1708 (N_1708,N_1285,N_1079);
and U1709 (N_1709,N_1269,N_1054);
or U1710 (N_1710,N_1265,N_1475);
nor U1711 (N_1711,N_1211,N_1202);
nand U1712 (N_1712,N_1015,N_1098);
and U1713 (N_1713,N_1255,N_1428);
nor U1714 (N_1714,N_1463,N_1103);
nor U1715 (N_1715,N_1168,N_1291);
nand U1716 (N_1716,N_1337,N_1268);
xor U1717 (N_1717,N_1385,N_1130);
and U1718 (N_1718,N_1138,N_1481);
xor U1719 (N_1719,N_1289,N_1158);
xnor U1720 (N_1720,N_1081,N_1427);
xnor U1721 (N_1721,N_1260,N_1351);
or U1722 (N_1722,N_1380,N_1328);
and U1723 (N_1723,N_1250,N_1034);
nand U1724 (N_1724,N_1053,N_1253);
xnor U1725 (N_1725,N_1041,N_1083);
or U1726 (N_1726,N_1433,N_1120);
and U1727 (N_1727,N_1457,N_1117);
and U1728 (N_1728,N_1028,N_1343);
nor U1729 (N_1729,N_1407,N_1058);
and U1730 (N_1730,N_1472,N_1398);
nor U1731 (N_1731,N_1139,N_1329);
nor U1732 (N_1732,N_1409,N_1066);
nand U1733 (N_1733,N_1226,N_1443);
or U1734 (N_1734,N_1333,N_1044);
nor U1735 (N_1735,N_1123,N_1429);
nor U1736 (N_1736,N_1025,N_1256);
or U1737 (N_1737,N_1453,N_1215);
and U1738 (N_1738,N_1325,N_1019);
and U1739 (N_1739,N_1049,N_1317);
nand U1740 (N_1740,N_1360,N_1097);
nor U1741 (N_1741,N_1449,N_1113);
nor U1742 (N_1742,N_1426,N_1104);
nand U1743 (N_1743,N_1061,N_1437);
or U1744 (N_1744,N_1145,N_1298);
nand U1745 (N_1745,N_1244,N_1150);
xnor U1746 (N_1746,N_1169,N_1365);
nor U1747 (N_1747,N_1354,N_1389);
and U1748 (N_1748,N_1399,N_1159);
and U1749 (N_1749,N_1128,N_1339);
or U1750 (N_1750,N_1382,N_1363);
nor U1751 (N_1751,N_1370,N_1495);
xnor U1752 (N_1752,N_1159,N_1206);
and U1753 (N_1753,N_1194,N_1357);
nor U1754 (N_1754,N_1058,N_1113);
nand U1755 (N_1755,N_1196,N_1389);
and U1756 (N_1756,N_1327,N_1372);
xnor U1757 (N_1757,N_1465,N_1383);
nand U1758 (N_1758,N_1466,N_1191);
or U1759 (N_1759,N_1049,N_1345);
nand U1760 (N_1760,N_1198,N_1038);
or U1761 (N_1761,N_1319,N_1426);
nor U1762 (N_1762,N_1038,N_1200);
and U1763 (N_1763,N_1234,N_1338);
nand U1764 (N_1764,N_1291,N_1207);
nor U1765 (N_1765,N_1228,N_1246);
or U1766 (N_1766,N_1298,N_1328);
or U1767 (N_1767,N_1252,N_1210);
nor U1768 (N_1768,N_1294,N_1164);
or U1769 (N_1769,N_1177,N_1139);
and U1770 (N_1770,N_1050,N_1367);
or U1771 (N_1771,N_1045,N_1019);
xor U1772 (N_1772,N_1199,N_1042);
nor U1773 (N_1773,N_1372,N_1382);
xor U1774 (N_1774,N_1469,N_1055);
and U1775 (N_1775,N_1336,N_1384);
or U1776 (N_1776,N_1147,N_1461);
or U1777 (N_1777,N_1239,N_1155);
nor U1778 (N_1778,N_1299,N_1121);
nand U1779 (N_1779,N_1202,N_1371);
xor U1780 (N_1780,N_1128,N_1055);
and U1781 (N_1781,N_1095,N_1262);
and U1782 (N_1782,N_1171,N_1227);
nand U1783 (N_1783,N_1347,N_1206);
nand U1784 (N_1784,N_1416,N_1058);
nor U1785 (N_1785,N_1240,N_1258);
and U1786 (N_1786,N_1144,N_1074);
or U1787 (N_1787,N_1068,N_1386);
nand U1788 (N_1788,N_1043,N_1230);
nand U1789 (N_1789,N_1256,N_1279);
xor U1790 (N_1790,N_1176,N_1140);
nor U1791 (N_1791,N_1447,N_1452);
xnor U1792 (N_1792,N_1069,N_1231);
nand U1793 (N_1793,N_1182,N_1129);
and U1794 (N_1794,N_1271,N_1327);
xnor U1795 (N_1795,N_1487,N_1128);
nor U1796 (N_1796,N_1044,N_1434);
and U1797 (N_1797,N_1192,N_1484);
nor U1798 (N_1798,N_1100,N_1049);
xnor U1799 (N_1799,N_1498,N_1307);
nor U1800 (N_1800,N_1287,N_1434);
nand U1801 (N_1801,N_1383,N_1434);
and U1802 (N_1802,N_1018,N_1386);
xnor U1803 (N_1803,N_1176,N_1041);
xnor U1804 (N_1804,N_1057,N_1183);
nor U1805 (N_1805,N_1444,N_1437);
nand U1806 (N_1806,N_1321,N_1291);
xnor U1807 (N_1807,N_1428,N_1416);
xnor U1808 (N_1808,N_1010,N_1182);
nand U1809 (N_1809,N_1262,N_1211);
nor U1810 (N_1810,N_1337,N_1144);
nor U1811 (N_1811,N_1020,N_1485);
xnor U1812 (N_1812,N_1083,N_1475);
and U1813 (N_1813,N_1338,N_1035);
xor U1814 (N_1814,N_1407,N_1246);
nand U1815 (N_1815,N_1121,N_1451);
nand U1816 (N_1816,N_1296,N_1266);
xor U1817 (N_1817,N_1070,N_1232);
and U1818 (N_1818,N_1241,N_1189);
nor U1819 (N_1819,N_1205,N_1071);
nand U1820 (N_1820,N_1055,N_1333);
xor U1821 (N_1821,N_1464,N_1217);
and U1822 (N_1822,N_1468,N_1153);
nor U1823 (N_1823,N_1180,N_1143);
nor U1824 (N_1824,N_1435,N_1218);
and U1825 (N_1825,N_1015,N_1272);
nor U1826 (N_1826,N_1279,N_1287);
and U1827 (N_1827,N_1399,N_1289);
xnor U1828 (N_1828,N_1054,N_1248);
or U1829 (N_1829,N_1075,N_1065);
xor U1830 (N_1830,N_1012,N_1064);
nand U1831 (N_1831,N_1150,N_1492);
xor U1832 (N_1832,N_1194,N_1228);
nor U1833 (N_1833,N_1363,N_1277);
nor U1834 (N_1834,N_1061,N_1029);
or U1835 (N_1835,N_1065,N_1121);
or U1836 (N_1836,N_1186,N_1029);
nand U1837 (N_1837,N_1349,N_1273);
nand U1838 (N_1838,N_1142,N_1231);
nand U1839 (N_1839,N_1206,N_1290);
and U1840 (N_1840,N_1288,N_1105);
nor U1841 (N_1841,N_1155,N_1186);
xnor U1842 (N_1842,N_1244,N_1421);
nor U1843 (N_1843,N_1173,N_1353);
and U1844 (N_1844,N_1204,N_1211);
nand U1845 (N_1845,N_1240,N_1178);
nand U1846 (N_1846,N_1362,N_1471);
nor U1847 (N_1847,N_1039,N_1487);
xnor U1848 (N_1848,N_1435,N_1051);
or U1849 (N_1849,N_1134,N_1314);
nand U1850 (N_1850,N_1185,N_1112);
xor U1851 (N_1851,N_1285,N_1386);
and U1852 (N_1852,N_1272,N_1164);
or U1853 (N_1853,N_1216,N_1205);
xnor U1854 (N_1854,N_1045,N_1208);
or U1855 (N_1855,N_1096,N_1343);
or U1856 (N_1856,N_1379,N_1114);
nor U1857 (N_1857,N_1472,N_1118);
nand U1858 (N_1858,N_1180,N_1161);
xnor U1859 (N_1859,N_1335,N_1178);
or U1860 (N_1860,N_1262,N_1440);
nor U1861 (N_1861,N_1122,N_1059);
nor U1862 (N_1862,N_1450,N_1432);
nor U1863 (N_1863,N_1177,N_1215);
nand U1864 (N_1864,N_1480,N_1058);
and U1865 (N_1865,N_1300,N_1118);
xor U1866 (N_1866,N_1137,N_1117);
nor U1867 (N_1867,N_1068,N_1038);
nor U1868 (N_1868,N_1216,N_1264);
xnor U1869 (N_1869,N_1182,N_1421);
xnor U1870 (N_1870,N_1174,N_1434);
nor U1871 (N_1871,N_1210,N_1043);
nand U1872 (N_1872,N_1100,N_1224);
or U1873 (N_1873,N_1053,N_1396);
nand U1874 (N_1874,N_1025,N_1143);
and U1875 (N_1875,N_1108,N_1452);
or U1876 (N_1876,N_1002,N_1036);
nor U1877 (N_1877,N_1146,N_1455);
nor U1878 (N_1878,N_1397,N_1150);
xnor U1879 (N_1879,N_1287,N_1186);
nor U1880 (N_1880,N_1085,N_1329);
nand U1881 (N_1881,N_1257,N_1067);
and U1882 (N_1882,N_1225,N_1188);
and U1883 (N_1883,N_1224,N_1452);
nor U1884 (N_1884,N_1262,N_1373);
nor U1885 (N_1885,N_1174,N_1030);
and U1886 (N_1886,N_1432,N_1087);
and U1887 (N_1887,N_1327,N_1262);
nor U1888 (N_1888,N_1014,N_1379);
or U1889 (N_1889,N_1345,N_1195);
and U1890 (N_1890,N_1104,N_1275);
xor U1891 (N_1891,N_1479,N_1443);
and U1892 (N_1892,N_1201,N_1339);
nand U1893 (N_1893,N_1274,N_1498);
and U1894 (N_1894,N_1171,N_1102);
or U1895 (N_1895,N_1163,N_1131);
or U1896 (N_1896,N_1149,N_1039);
nor U1897 (N_1897,N_1351,N_1342);
nor U1898 (N_1898,N_1296,N_1412);
nand U1899 (N_1899,N_1335,N_1143);
and U1900 (N_1900,N_1421,N_1339);
nand U1901 (N_1901,N_1422,N_1102);
nand U1902 (N_1902,N_1410,N_1468);
and U1903 (N_1903,N_1119,N_1020);
or U1904 (N_1904,N_1341,N_1265);
nand U1905 (N_1905,N_1499,N_1341);
nand U1906 (N_1906,N_1006,N_1405);
or U1907 (N_1907,N_1006,N_1071);
nand U1908 (N_1908,N_1145,N_1305);
and U1909 (N_1909,N_1445,N_1071);
and U1910 (N_1910,N_1051,N_1033);
or U1911 (N_1911,N_1345,N_1496);
nand U1912 (N_1912,N_1396,N_1169);
nor U1913 (N_1913,N_1309,N_1366);
or U1914 (N_1914,N_1423,N_1087);
and U1915 (N_1915,N_1073,N_1163);
or U1916 (N_1916,N_1280,N_1297);
nor U1917 (N_1917,N_1434,N_1278);
and U1918 (N_1918,N_1091,N_1073);
nor U1919 (N_1919,N_1170,N_1441);
or U1920 (N_1920,N_1279,N_1273);
nand U1921 (N_1921,N_1094,N_1398);
and U1922 (N_1922,N_1278,N_1062);
nor U1923 (N_1923,N_1002,N_1412);
or U1924 (N_1924,N_1117,N_1034);
and U1925 (N_1925,N_1203,N_1447);
xnor U1926 (N_1926,N_1202,N_1353);
nand U1927 (N_1927,N_1212,N_1308);
nand U1928 (N_1928,N_1378,N_1391);
nand U1929 (N_1929,N_1124,N_1182);
and U1930 (N_1930,N_1087,N_1328);
nor U1931 (N_1931,N_1238,N_1211);
nand U1932 (N_1932,N_1243,N_1311);
xnor U1933 (N_1933,N_1387,N_1487);
or U1934 (N_1934,N_1458,N_1255);
or U1935 (N_1935,N_1277,N_1188);
nand U1936 (N_1936,N_1325,N_1278);
and U1937 (N_1937,N_1397,N_1152);
or U1938 (N_1938,N_1280,N_1041);
nor U1939 (N_1939,N_1255,N_1378);
xnor U1940 (N_1940,N_1185,N_1474);
xnor U1941 (N_1941,N_1031,N_1427);
and U1942 (N_1942,N_1098,N_1459);
nand U1943 (N_1943,N_1106,N_1479);
nand U1944 (N_1944,N_1422,N_1441);
nor U1945 (N_1945,N_1072,N_1475);
nand U1946 (N_1946,N_1398,N_1124);
or U1947 (N_1947,N_1468,N_1114);
nand U1948 (N_1948,N_1254,N_1399);
or U1949 (N_1949,N_1014,N_1013);
xnor U1950 (N_1950,N_1215,N_1068);
or U1951 (N_1951,N_1322,N_1389);
nand U1952 (N_1952,N_1231,N_1431);
or U1953 (N_1953,N_1262,N_1115);
or U1954 (N_1954,N_1148,N_1007);
nand U1955 (N_1955,N_1308,N_1409);
xor U1956 (N_1956,N_1182,N_1077);
nor U1957 (N_1957,N_1441,N_1153);
or U1958 (N_1958,N_1309,N_1383);
nor U1959 (N_1959,N_1143,N_1035);
nand U1960 (N_1960,N_1055,N_1269);
nor U1961 (N_1961,N_1000,N_1296);
or U1962 (N_1962,N_1172,N_1257);
and U1963 (N_1963,N_1237,N_1441);
and U1964 (N_1964,N_1378,N_1165);
and U1965 (N_1965,N_1455,N_1119);
xnor U1966 (N_1966,N_1409,N_1234);
nand U1967 (N_1967,N_1106,N_1057);
nor U1968 (N_1968,N_1028,N_1015);
nor U1969 (N_1969,N_1411,N_1023);
xor U1970 (N_1970,N_1395,N_1450);
or U1971 (N_1971,N_1124,N_1376);
and U1972 (N_1972,N_1151,N_1242);
or U1973 (N_1973,N_1234,N_1079);
nor U1974 (N_1974,N_1129,N_1349);
nand U1975 (N_1975,N_1480,N_1405);
and U1976 (N_1976,N_1081,N_1073);
xor U1977 (N_1977,N_1291,N_1360);
nor U1978 (N_1978,N_1389,N_1092);
xor U1979 (N_1979,N_1392,N_1186);
nor U1980 (N_1980,N_1479,N_1013);
and U1981 (N_1981,N_1333,N_1345);
or U1982 (N_1982,N_1220,N_1394);
xor U1983 (N_1983,N_1118,N_1137);
and U1984 (N_1984,N_1185,N_1062);
xor U1985 (N_1985,N_1417,N_1366);
nor U1986 (N_1986,N_1047,N_1337);
or U1987 (N_1987,N_1494,N_1077);
and U1988 (N_1988,N_1372,N_1482);
xnor U1989 (N_1989,N_1184,N_1131);
and U1990 (N_1990,N_1241,N_1045);
nand U1991 (N_1991,N_1428,N_1002);
nor U1992 (N_1992,N_1401,N_1009);
nand U1993 (N_1993,N_1118,N_1024);
nand U1994 (N_1994,N_1289,N_1483);
and U1995 (N_1995,N_1255,N_1442);
and U1996 (N_1996,N_1183,N_1149);
nand U1997 (N_1997,N_1013,N_1097);
or U1998 (N_1998,N_1372,N_1155);
nand U1999 (N_1999,N_1258,N_1191);
nand U2000 (N_2000,N_1608,N_1650);
and U2001 (N_2001,N_1508,N_1934);
xnor U2002 (N_2002,N_1577,N_1639);
xnor U2003 (N_2003,N_1759,N_1788);
and U2004 (N_2004,N_1837,N_1509);
xor U2005 (N_2005,N_1894,N_1814);
nand U2006 (N_2006,N_1998,N_1529);
or U2007 (N_2007,N_1825,N_1584);
or U2008 (N_2008,N_1751,N_1607);
and U2009 (N_2009,N_1510,N_1642);
nand U2010 (N_2010,N_1747,N_1551);
nand U2011 (N_2011,N_1739,N_1878);
and U2012 (N_2012,N_1968,N_1810);
or U2013 (N_2013,N_1775,N_1920);
and U2014 (N_2014,N_1909,N_1807);
and U2015 (N_2015,N_1595,N_1827);
nand U2016 (N_2016,N_1734,N_1724);
and U2017 (N_2017,N_1627,N_1873);
nor U2018 (N_2018,N_1527,N_1903);
or U2019 (N_2019,N_1728,N_1717);
and U2020 (N_2020,N_1944,N_1780);
and U2021 (N_2021,N_1783,N_1645);
nand U2022 (N_2022,N_1541,N_1581);
xor U2023 (N_2023,N_1742,N_1950);
or U2024 (N_2024,N_1953,N_1905);
nor U2025 (N_2025,N_1557,N_1779);
xor U2026 (N_2026,N_1749,N_1987);
and U2027 (N_2027,N_1578,N_1802);
nand U2028 (N_2028,N_1815,N_1988);
xor U2029 (N_2029,N_1892,N_1659);
nand U2030 (N_2030,N_1971,N_1567);
nor U2031 (N_2031,N_1633,N_1689);
and U2032 (N_2032,N_1958,N_1915);
or U2033 (N_2033,N_1593,N_1952);
and U2034 (N_2034,N_1670,N_1580);
and U2035 (N_2035,N_1757,N_1564);
nor U2036 (N_2036,N_1525,N_1682);
or U2037 (N_2037,N_1907,N_1705);
nand U2038 (N_2038,N_1972,N_1696);
nor U2039 (N_2039,N_1517,N_1543);
and U2040 (N_2040,N_1756,N_1974);
nor U2041 (N_2041,N_1748,N_1550);
nor U2042 (N_2042,N_1686,N_1745);
and U2043 (N_2043,N_1694,N_1701);
and U2044 (N_2044,N_1594,N_1874);
nand U2045 (N_2045,N_1755,N_1722);
and U2046 (N_2046,N_1604,N_1771);
xnor U2047 (N_2047,N_1855,N_1600);
nand U2048 (N_2048,N_1621,N_1610);
nor U2049 (N_2049,N_1927,N_1678);
and U2050 (N_2050,N_1785,N_1723);
xor U2051 (N_2051,N_1556,N_1570);
and U2052 (N_2052,N_1673,N_1546);
or U2053 (N_2053,N_1991,N_1753);
or U2054 (N_2054,N_1959,N_1769);
xor U2055 (N_2055,N_1778,N_1799);
and U2056 (N_2056,N_1711,N_1962);
nand U2057 (N_2057,N_1663,N_1926);
xnor U2058 (N_2058,N_1754,N_1982);
or U2059 (N_2059,N_1812,N_1572);
nand U2060 (N_2060,N_1822,N_1583);
or U2061 (N_2061,N_1830,N_1811);
and U2062 (N_2062,N_1922,N_1851);
xor U2063 (N_2063,N_1538,N_1699);
xnor U2064 (N_2064,N_1895,N_1654);
nand U2065 (N_2065,N_1619,N_1626);
xnor U2066 (N_2066,N_1732,N_1881);
and U2067 (N_2067,N_1667,N_1537);
and U2068 (N_2068,N_1648,N_1863);
nor U2069 (N_2069,N_1816,N_1957);
nor U2070 (N_2070,N_1932,N_1976);
nand U2071 (N_2071,N_1929,N_1609);
xor U2072 (N_2072,N_1871,N_1866);
or U2073 (N_2073,N_1782,N_1946);
and U2074 (N_2074,N_1676,N_1504);
nor U2075 (N_2075,N_1582,N_1542);
nand U2076 (N_2076,N_1938,N_1908);
xnor U2077 (N_2077,N_1949,N_1970);
nor U2078 (N_2078,N_1733,N_1801);
nand U2079 (N_2079,N_1930,N_1875);
nor U2080 (N_2080,N_1836,N_1777);
nand U2081 (N_2081,N_1740,N_1679);
nor U2082 (N_2082,N_1960,N_1591);
nor U2083 (N_2083,N_1692,N_1576);
xnor U2084 (N_2084,N_1973,N_1620);
nor U2085 (N_2085,N_1804,N_1977);
nand U2086 (N_2086,N_1884,N_1640);
nor U2087 (N_2087,N_1945,N_1710);
nor U2088 (N_2088,N_1687,N_1603);
xnor U2089 (N_2089,N_1616,N_1993);
nor U2090 (N_2090,N_1649,N_1554);
or U2091 (N_2091,N_1513,N_1916);
nand U2092 (N_2092,N_1688,N_1684);
nand U2093 (N_2093,N_1773,N_1843);
and U2094 (N_2094,N_1937,N_1795);
or U2095 (N_2095,N_1713,N_1984);
nand U2096 (N_2096,N_1760,N_1540);
xor U2097 (N_2097,N_1997,N_1752);
xor U2098 (N_2098,N_1897,N_1887);
or U2099 (N_2099,N_1790,N_1715);
nand U2100 (N_2100,N_1768,N_1992);
or U2101 (N_2101,N_1501,N_1899);
nand U2102 (N_2102,N_1622,N_1856);
nor U2103 (N_2103,N_1911,N_1906);
xor U2104 (N_2104,N_1615,N_1956);
xnor U2105 (N_2105,N_1560,N_1561);
or U2106 (N_2106,N_1628,N_1794);
nand U2107 (N_2107,N_1872,N_1625);
xnor U2108 (N_2108,N_1720,N_1512);
and U2109 (N_2109,N_1826,N_1562);
and U2110 (N_2110,N_1921,N_1936);
nor U2111 (N_2111,N_1672,N_1526);
nor U2112 (N_2112,N_1571,N_1889);
and U2113 (N_2113,N_1664,N_1941);
or U2114 (N_2114,N_1716,N_1511);
and U2115 (N_2115,N_1796,N_1879);
xor U2116 (N_2116,N_1803,N_1961);
nor U2117 (N_2117,N_1985,N_1566);
xor U2118 (N_2118,N_1900,N_1712);
or U2119 (N_2119,N_1709,N_1690);
nor U2120 (N_2120,N_1635,N_1661);
or U2121 (N_2121,N_1767,N_1821);
nand U2122 (N_2122,N_1763,N_1736);
nand U2123 (N_2123,N_1939,N_1677);
nand U2124 (N_2124,N_1784,N_1641);
nor U2125 (N_2125,N_1555,N_1935);
or U2126 (N_2126,N_1611,N_1902);
and U2127 (N_2127,N_1854,N_1986);
nor U2128 (N_2128,N_1657,N_1806);
nor U2129 (N_2129,N_1592,N_1698);
and U2130 (N_2130,N_1703,N_1589);
nand U2131 (N_2131,N_1617,N_1853);
nor U2132 (N_2132,N_1634,N_1738);
and U2133 (N_2133,N_1762,N_1590);
nand U2134 (N_2134,N_1612,N_1776);
or U2135 (N_2135,N_1868,N_1652);
nand U2136 (N_2136,N_1817,N_1597);
and U2137 (N_2137,N_1864,N_1893);
or U2138 (N_2138,N_1861,N_1516);
nand U2139 (N_2139,N_1500,N_1823);
and U2140 (N_2140,N_1841,N_1613);
nor U2141 (N_2141,N_1539,N_1840);
or U2142 (N_2142,N_1766,N_1727);
nand U2143 (N_2143,N_1587,N_1898);
nor U2144 (N_2144,N_1585,N_1791);
and U2145 (N_2145,N_1913,N_1521);
xor U2146 (N_2146,N_1813,N_1553);
and U2147 (N_2147,N_1990,N_1618);
nor U2148 (N_2148,N_1919,N_1725);
or U2149 (N_2149,N_1805,N_1636);
or U2150 (N_2150,N_1744,N_1505);
xnor U2151 (N_2151,N_1629,N_1928);
or U2152 (N_2152,N_1731,N_1808);
nand U2153 (N_2153,N_1647,N_1523);
and U2154 (N_2154,N_1832,N_1844);
nor U2155 (N_2155,N_1979,N_1774);
and U2156 (N_2156,N_1859,N_1552);
and U2157 (N_2157,N_1666,N_1644);
nand U2158 (N_2158,N_1786,N_1781);
nor U2159 (N_2159,N_1519,N_1573);
nor U2160 (N_2160,N_1846,N_1707);
nand U2161 (N_2161,N_1995,N_1917);
nand U2162 (N_2162,N_1602,N_1730);
nand U2163 (N_2163,N_1865,N_1877);
or U2164 (N_2164,N_1924,N_1758);
xor U2165 (N_2165,N_1849,N_1764);
xnor U2166 (N_2166,N_1518,N_1850);
nor U2167 (N_2167,N_1965,N_1520);
xnor U2168 (N_2168,N_1901,N_1630);
nor U2169 (N_2169,N_1914,N_1721);
xor U2170 (N_2170,N_1536,N_1503);
and U2171 (N_2171,N_1656,N_1923);
xnor U2172 (N_2172,N_1870,N_1624);
xor U2173 (N_2173,N_1506,N_1704);
nand U2174 (N_2174,N_1691,N_1708);
or U2175 (N_2175,N_1706,N_1588);
and U2176 (N_2176,N_1798,N_1789);
nor U2177 (N_2177,N_1535,N_1896);
nor U2178 (N_2178,N_1770,N_1833);
xor U2179 (N_2179,N_1829,N_1955);
nor U2180 (N_2180,N_1606,N_1533);
nor U2181 (N_2181,N_1680,N_1981);
nor U2182 (N_2182,N_1765,N_1876);
or U2183 (N_2183,N_1668,N_1651);
and U2184 (N_2184,N_1869,N_1662);
xnor U2185 (N_2185,N_1653,N_1835);
or U2186 (N_2186,N_1983,N_1940);
nand U2187 (N_2187,N_1596,N_1507);
nor U2188 (N_2188,N_1999,N_1514);
xor U2189 (N_2189,N_1632,N_1559);
or U2190 (N_2190,N_1532,N_1834);
and U2191 (N_2191,N_1809,N_1681);
and U2192 (N_2192,N_1643,N_1947);
and U2193 (N_2193,N_1729,N_1714);
nor U2194 (N_2194,N_1671,N_1693);
and U2195 (N_2195,N_1631,N_1820);
nor U2196 (N_2196,N_1646,N_1669);
or U2197 (N_2197,N_1867,N_1746);
nor U2198 (N_2198,N_1792,N_1989);
nand U2199 (N_2199,N_1658,N_1954);
nor U2200 (N_2200,N_1951,N_1980);
or U2201 (N_2201,N_1967,N_1996);
nor U2202 (N_2202,N_1918,N_1761);
and U2203 (N_2203,N_1697,N_1601);
nor U2204 (N_2204,N_1530,N_1549);
xor U2205 (N_2205,N_1568,N_1569);
nor U2206 (N_2206,N_1531,N_1660);
and U2207 (N_2207,N_1515,N_1637);
nor U2208 (N_2208,N_1528,N_1824);
or U2209 (N_2209,N_1638,N_1737);
and U2210 (N_2210,N_1857,N_1838);
and U2211 (N_2211,N_1623,N_1675);
and U2212 (N_2212,N_1547,N_1735);
or U2213 (N_2213,N_1793,N_1545);
and U2214 (N_2214,N_1858,N_1502);
xor U2215 (N_2215,N_1524,N_1978);
or U2216 (N_2216,N_1655,N_1800);
xnor U2217 (N_2217,N_1888,N_1586);
xnor U2218 (N_2218,N_1994,N_1674);
xor U2219 (N_2219,N_1522,N_1614);
and U2220 (N_2220,N_1852,N_1548);
nor U2221 (N_2221,N_1750,N_1904);
nand U2222 (N_2222,N_1719,N_1565);
or U2223 (N_2223,N_1885,N_1579);
nor U2224 (N_2224,N_1563,N_1700);
nor U2225 (N_2225,N_1695,N_1683);
and U2226 (N_2226,N_1845,N_1743);
and U2227 (N_2227,N_1842,N_1599);
nand U2228 (N_2228,N_1741,N_1910);
and U2229 (N_2229,N_1797,N_1558);
and U2230 (N_2230,N_1702,N_1891);
and U2231 (N_2231,N_1819,N_1726);
and U2232 (N_2232,N_1943,N_1818);
or U2233 (N_2233,N_1605,N_1948);
xnor U2234 (N_2234,N_1860,N_1847);
and U2235 (N_2235,N_1925,N_1882);
nor U2236 (N_2236,N_1574,N_1975);
or U2237 (N_2237,N_1969,N_1862);
nand U2238 (N_2238,N_1963,N_1831);
and U2239 (N_2239,N_1665,N_1883);
or U2240 (N_2240,N_1828,N_1718);
nor U2241 (N_2241,N_1544,N_1964);
and U2242 (N_2242,N_1685,N_1966);
nand U2243 (N_2243,N_1942,N_1839);
or U2244 (N_2244,N_1912,N_1787);
xnor U2245 (N_2245,N_1931,N_1886);
xor U2246 (N_2246,N_1890,N_1575);
nand U2247 (N_2247,N_1848,N_1534);
xor U2248 (N_2248,N_1933,N_1772);
nand U2249 (N_2249,N_1598,N_1880);
xor U2250 (N_2250,N_1823,N_1899);
xor U2251 (N_2251,N_1714,N_1906);
xor U2252 (N_2252,N_1528,N_1825);
xor U2253 (N_2253,N_1543,N_1963);
xor U2254 (N_2254,N_1731,N_1655);
nor U2255 (N_2255,N_1602,N_1864);
xor U2256 (N_2256,N_1579,N_1561);
nor U2257 (N_2257,N_1748,N_1938);
xor U2258 (N_2258,N_1527,N_1955);
and U2259 (N_2259,N_1570,N_1863);
and U2260 (N_2260,N_1648,N_1722);
xor U2261 (N_2261,N_1959,N_1509);
or U2262 (N_2262,N_1841,N_1521);
xor U2263 (N_2263,N_1609,N_1786);
or U2264 (N_2264,N_1547,N_1759);
or U2265 (N_2265,N_1810,N_1958);
xor U2266 (N_2266,N_1901,N_1912);
nor U2267 (N_2267,N_1576,N_1547);
nor U2268 (N_2268,N_1578,N_1503);
and U2269 (N_2269,N_1761,N_1534);
or U2270 (N_2270,N_1727,N_1769);
or U2271 (N_2271,N_1690,N_1997);
or U2272 (N_2272,N_1683,N_1648);
xnor U2273 (N_2273,N_1717,N_1610);
or U2274 (N_2274,N_1540,N_1987);
nand U2275 (N_2275,N_1603,N_1975);
and U2276 (N_2276,N_1642,N_1543);
or U2277 (N_2277,N_1812,N_1948);
and U2278 (N_2278,N_1692,N_1687);
and U2279 (N_2279,N_1712,N_1635);
or U2280 (N_2280,N_1522,N_1709);
or U2281 (N_2281,N_1939,N_1585);
or U2282 (N_2282,N_1547,N_1737);
nand U2283 (N_2283,N_1656,N_1932);
nor U2284 (N_2284,N_1703,N_1916);
nor U2285 (N_2285,N_1730,N_1982);
or U2286 (N_2286,N_1916,N_1641);
and U2287 (N_2287,N_1979,N_1933);
nand U2288 (N_2288,N_1664,N_1644);
xor U2289 (N_2289,N_1908,N_1813);
xor U2290 (N_2290,N_1887,N_1751);
or U2291 (N_2291,N_1524,N_1780);
xor U2292 (N_2292,N_1907,N_1667);
nor U2293 (N_2293,N_1510,N_1507);
nor U2294 (N_2294,N_1691,N_1625);
or U2295 (N_2295,N_1543,N_1554);
or U2296 (N_2296,N_1803,N_1926);
nor U2297 (N_2297,N_1613,N_1896);
xnor U2298 (N_2298,N_1503,N_1667);
xnor U2299 (N_2299,N_1769,N_1534);
nor U2300 (N_2300,N_1953,N_1883);
or U2301 (N_2301,N_1831,N_1823);
or U2302 (N_2302,N_1653,N_1920);
and U2303 (N_2303,N_1970,N_1987);
xnor U2304 (N_2304,N_1545,N_1962);
nand U2305 (N_2305,N_1664,N_1812);
and U2306 (N_2306,N_1904,N_1579);
or U2307 (N_2307,N_1653,N_1720);
or U2308 (N_2308,N_1811,N_1502);
and U2309 (N_2309,N_1607,N_1932);
nor U2310 (N_2310,N_1973,N_1931);
nor U2311 (N_2311,N_1716,N_1976);
nand U2312 (N_2312,N_1778,N_1942);
xor U2313 (N_2313,N_1855,N_1999);
and U2314 (N_2314,N_1519,N_1541);
and U2315 (N_2315,N_1704,N_1745);
nor U2316 (N_2316,N_1685,N_1680);
and U2317 (N_2317,N_1525,N_1553);
nor U2318 (N_2318,N_1655,N_1600);
xnor U2319 (N_2319,N_1751,N_1508);
or U2320 (N_2320,N_1580,N_1726);
nor U2321 (N_2321,N_1996,N_1577);
or U2322 (N_2322,N_1743,N_1728);
and U2323 (N_2323,N_1574,N_1892);
nand U2324 (N_2324,N_1750,N_1888);
or U2325 (N_2325,N_1867,N_1580);
or U2326 (N_2326,N_1633,N_1825);
nor U2327 (N_2327,N_1970,N_1581);
and U2328 (N_2328,N_1528,N_1862);
xor U2329 (N_2329,N_1633,N_1987);
nand U2330 (N_2330,N_1935,N_1964);
nand U2331 (N_2331,N_1944,N_1770);
and U2332 (N_2332,N_1653,N_1826);
nor U2333 (N_2333,N_1557,N_1693);
nand U2334 (N_2334,N_1617,N_1644);
nand U2335 (N_2335,N_1896,N_1655);
or U2336 (N_2336,N_1636,N_1683);
xnor U2337 (N_2337,N_1746,N_1982);
or U2338 (N_2338,N_1505,N_1845);
and U2339 (N_2339,N_1527,N_1636);
and U2340 (N_2340,N_1769,N_1983);
nor U2341 (N_2341,N_1521,N_1685);
nand U2342 (N_2342,N_1587,N_1677);
nor U2343 (N_2343,N_1543,N_1831);
nor U2344 (N_2344,N_1929,N_1664);
and U2345 (N_2345,N_1662,N_1644);
nor U2346 (N_2346,N_1849,N_1629);
and U2347 (N_2347,N_1595,N_1737);
and U2348 (N_2348,N_1981,N_1922);
and U2349 (N_2349,N_1705,N_1692);
and U2350 (N_2350,N_1660,N_1838);
or U2351 (N_2351,N_1511,N_1831);
and U2352 (N_2352,N_1507,N_1629);
and U2353 (N_2353,N_1555,N_1981);
nor U2354 (N_2354,N_1909,N_1845);
nand U2355 (N_2355,N_1835,N_1896);
nand U2356 (N_2356,N_1603,N_1613);
xor U2357 (N_2357,N_1714,N_1856);
nor U2358 (N_2358,N_1783,N_1810);
xor U2359 (N_2359,N_1815,N_1885);
or U2360 (N_2360,N_1703,N_1812);
or U2361 (N_2361,N_1503,N_1898);
or U2362 (N_2362,N_1929,N_1700);
xnor U2363 (N_2363,N_1687,N_1675);
and U2364 (N_2364,N_1554,N_1560);
or U2365 (N_2365,N_1902,N_1595);
nor U2366 (N_2366,N_1969,N_1630);
nand U2367 (N_2367,N_1966,N_1642);
and U2368 (N_2368,N_1840,N_1760);
nand U2369 (N_2369,N_1901,N_1780);
or U2370 (N_2370,N_1652,N_1644);
and U2371 (N_2371,N_1665,N_1714);
nor U2372 (N_2372,N_1779,N_1981);
nor U2373 (N_2373,N_1902,N_1935);
or U2374 (N_2374,N_1654,N_1752);
and U2375 (N_2375,N_1592,N_1566);
and U2376 (N_2376,N_1971,N_1915);
or U2377 (N_2377,N_1550,N_1733);
and U2378 (N_2378,N_1930,N_1518);
nor U2379 (N_2379,N_1757,N_1840);
xor U2380 (N_2380,N_1759,N_1959);
xnor U2381 (N_2381,N_1931,N_1725);
and U2382 (N_2382,N_1683,N_1947);
xnor U2383 (N_2383,N_1574,N_1772);
and U2384 (N_2384,N_1902,N_1523);
and U2385 (N_2385,N_1785,N_1636);
nor U2386 (N_2386,N_1959,N_1594);
xnor U2387 (N_2387,N_1801,N_1687);
or U2388 (N_2388,N_1558,N_1512);
nor U2389 (N_2389,N_1636,N_1778);
xor U2390 (N_2390,N_1653,N_1567);
and U2391 (N_2391,N_1926,N_1826);
or U2392 (N_2392,N_1609,N_1921);
xor U2393 (N_2393,N_1542,N_1833);
nor U2394 (N_2394,N_1520,N_1726);
nand U2395 (N_2395,N_1561,N_1617);
nor U2396 (N_2396,N_1743,N_1805);
nor U2397 (N_2397,N_1825,N_1886);
xnor U2398 (N_2398,N_1684,N_1708);
and U2399 (N_2399,N_1899,N_1588);
and U2400 (N_2400,N_1767,N_1592);
nand U2401 (N_2401,N_1618,N_1753);
or U2402 (N_2402,N_1744,N_1595);
nor U2403 (N_2403,N_1684,N_1545);
nand U2404 (N_2404,N_1529,N_1980);
nor U2405 (N_2405,N_1561,N_1778);
nand U2406 (N_2406,N_1806,N_1961);
or U2407 (N_2407,N_1641,N_1613);
or U2408 (N_2408,N_1816,N_1893);
or U2409 (N_2409,N_1660,N_1690);
or U2410 (N_2410,N_1787,N_1967);
and U2411 (N_2411,N_1925,N_1704);
nor U2412 (N_2412,N_1933,N_1969);
and U2413 (N_2413,N_1829,N_1631);
xor U2414 (N_2414,N_1966,N_1854);
or U2415 (N_2415,N_1744,N_1596);
or U2416 (N_2416,N_1539,N_1664);
nand U2417 (N_2417,N_1620,N_1707);
or U2418 (N_2418,N_1692,N_1570);
and U2419 (N_2419,N_1700,N_1503);
or U2420 (N_2420,N_1635,N_1607);
and U2421 (N_2421,N_1677,N_1632);
xnor U2422 (N_2422,N_1866,N_1927);
or U2423 (N_2423,N_1701,N_1612);
nor U2424 (N_2424,N_1979,N_1519);
xnor U2425 (N_2425,N_1603,N_1825);
nor U2426 (N_2426,N_1726,N_1845);
nor U2427 (N_2427,N_1851,N_1623);
or U2428 (N_2428,N_1872,N_1888);
or U2429 (N_2429,N_1543,N_1600);
nand U2430 (N_2430,N_1984,N_1658);
or U2431 (N_2431,N_1705,N_1727);
xor U2432 (N_2432,N_1651,N_1663);
xor U2433 (N_2433,N_1569,N_1761);
nor U2434 (N_2434,N_1893,N_1831);
xor U2435 (N_2435,N_1861,N_1913);
nor U2436 (N_2436,N_1710,N_1910);
and U2437 (N_2437,N_1693,N_1998);
nand U2438 (N_2438,N_1762,N_1588);
nor U2439 (N_2439,N_1957,N_1992);
nor U2440 (N_2440,N_1610,N_1830);
and U2441 (N_2441,N_1500,N_1868);
nor U2442 (N_2442,N_1722,N_1638);
or U2443 (N_2443,N_1660,N_1632);
or U2444 (N_2444,N_1521,N_1931);
nand U2445 (N_2445,N_1607,N_1544);
nor U2446 (N_2446,N_1987,N_1864);
or U2447 (N_2447,N_1939,N_1757);
or U2448 (N_2448,N_1778,N_1758);
nor U2449 (N_2449,N_1800,N_1907);
nand U2450 (N_2450,N_1841,N_1652);
nand U2451 (N_2451,N_1770,N_1909);
and U2452 (N_2452,N_1987,N_1998);
or U2453 (N_2453,N_1826,N_1640);
nand U2454 (N_2454,N_1741,N_1795);
or U2455 (N_2455,N_1912,N_1702);
and U2456 (N_2456,N_1710,N_1967);
and U2457 (N_2457,N_1544,N_1711);
or U2458 (N_2458,N_1839,N_1703);
nor U2459 (N_2459,N_1907,N_1966);
nand U2460 (N_2460,N_1873,N_1506);
nand U2461 (N_2461,N_1678,N_1687);
nor U2462 (N_2462,N_1946,N_1544);
and U2463 (N_2463,N_1781,N_1506);
and U2464 (N_2464,N_1624,N_1600);
xor U2465 (N_2465,N_1514,N_1905);
xnor U2466 (N_2466,N_1776,N_1815);
nor U2467 (N_2467,N_1834,N_1779);
xor U2468 (N_2468,N_1885,N_1660);
and U2469 (N_2469,N_1770,N_1695);
nand U2470 (N_2470,N_1879,N_1858);
or U2471 (N_2471,N_1664,N_1681);
nand U2472 (N_2472,N_1732,N_1791);
xnor U2473 (N_2473,N_1726,N_1899);
nor U2474 (N_2474,N_1661,N_1848);
and U2475 (N_2475,N_1537,N_1656);
nand U2476 (N_2476,N_1743,N_1868);
or U2477 (N_2477,N_1612,N_1743);
or U2478 (N_2478,N_1797,N_1521);
nand U2479 (N_2479,N_1764,N_1854);
and U2480 (N_2480,N_1658,N_1807);
nor U2481 (N_2481,N_1915,N_1738);
or U2482 (N_2482,N_1894,N_1594);
or U2483 (N_2483,N_1948,N_1749);
nor U2484 (N_2484,N_1922,N_1756);
or U2485 (N_2485,N_1687,N_1833);
nor U2486 (N_2486,N_1867,N_1912);
nor U2487 (N_2487,N_1881,N_1728);
or U2488 (N_2488,N_1584,N_1812);
nor U2489 (N_2489,N_1690,N_1821);
nor U2490 (N_2490,N_1761,N_1919);
xnor U2491 (N_2491,N_1770,N_1605);
and U2492 (N_2492,N_1955,N_1935);
nand U2493 (N_2493,N_1590,N_1741);
xor U2494 (N_2494,N_1780,N_1605);
or U2495 (N_2495,N_1679,N_1850);
xnor U2496 (N_2496,N_1823,N_1632);
nor U2497 (N_2497,N_1754,N_1933);
nand U2498 (N_2498,N_1840,N_1548);
xnor U2499 (N_2499,N_1632,N_1884);
or U2500 (N_2500,N_2051,N_2095);
xor U2501 (N_2501,N_2307,N_2458);
or U2502 (N_2502,N_2204,N_2322);
and U2503 (N_2503,N_2323,N_2304);
nand U2504 (N_2504,N_2468,N_2412);
nand U2505 (N_2505,N_2014,N_2108);
nor U2506 (N_2506,N_2290,N_2033);
nand U2507 (N_2507,N_2371,N_2081);
and U2508 (N_2508,N_2293,N_2182);
nand U2509 (N_2509,N_2274,N_2329);
and U2510 (N_2510,N_2202,N_2038);
nand U2511 (N_2511,N_2024,N_2223);
or U2512 (N_2512,N_2076,N_2395);
nor U2513 (N_2513,N_2111,N_2421);
xor U2514 (N_2514,N_2214,N_2338);
nor U2515 (N_2515,N_2445,N_2093);
nand U2516 (N_2516,N_2449,N_2391);
and U2517 (N_2517,N_2281,N_2004);
nand U2518 (N_2518,N_2492,N_2339);
nor U2519 (N_2519,N_2297,N_2150);
or U2520 (N_2520,N_2061,N_2369);
nor U2521 (N_2521,N_2074,N_2244);
and U2522 (N_2522,N_2013,N_2264);
or U2523 (N_2523,N_2349,N_2473);
xor U2524 (N_2524,N_2393,N_2071);
nand U2525 (N_2525,N_2318,N_2390);
nor U2526 (N_2526,N_2341,N_2016);
or U2527 (N_2527,N_2464,N_2092);
nand U2528 (N_2528,N_2163,N_2463);
or U2529 (N_2529,N_2428,N_2087);
or U2530 (N_2530,N_2450,N_2257);
and U2531 (N_2531,N_2226,N_2357);
nor U2532 (N_2532,N_2165,N_2188);
xor U2533 (N_2533,N_2285,N_2288);
nand U2534 (N_2534,N_2020,N_2403);
and U2535 (N_2535,N_2132,N_2229);
xnor U2536 (N_2536,N_2175,N_2139);
xnor U2537 (N_2537,N_2496,N_2106);
and U2538 (N_2538,N_2153,N_2373);
and U2539 (N_2539,N_2306,N_2439);
nor U2540 (N_2540,N_2177,N_2392);
nand U2541 (N_2541,N_2089,N_2030);
xor U2542 (N_2542,N_2054,N_2027);
xnor U2543 (N_2543,N_2101,N_2317);
or U2544 (N_2544,N_2408,N_2258);
or U2545 (N_2545,N_2047,N_2032);
nand U2546 (N_2546,N_2401,N_2495);
nor U2547 (N_2547,N_2066,N_2220);
and U2548 (N_2548,N_2482,N_2007);
and U2549 (N_2549,N_2319,N_2480);
or U2550 (N_2550,N_2140,N_2266);
nand U2551 (N_2551,N_2242,N_2079);
nand U2552 (N_2552,N_2372,N_2042);
and U2553 (N_2553,N_2159,N_2134);
nor U2554 (N_2554,N_2174,N_2298);
xnor U2555 (N_2555,N_2368,N_2173);
xnor U2556 (N_2556,N_2295,N_2299);
nand U2557 (N_2557,N_2073,N_2096);
and U2558 (N_2558,N_2351,N_2481);
nand U2559 (N_2559,N_2107,N_2334);
xnor U2560 (N_2560,N_2055,N_2219);
nor U2561 (N_2561,N_2147,N_2465);
nor U2562 (N_2562,N_2197,N_2354);
nor U2563 (N_2563,N_2353,N_2275);
xor U2564 (N_2564,N_2327,N_2417);
or U2565 (N_2565,N_2470,N_2386);
nand U2566 (N_2566,N_2179,N_2387);
or U2567 (N_2567,N_2355,N_2454);
or U2568 (N_2568,N_2120,N_2234);
or U2569 (N_2569,N_2041,N_2447);
xor U2570 (N_2570,N_2186,N_2017);
nor U2571 (N_2571,N_2483,N_2021);
nor U2572 (N_2572,N_2494,N_2067);
and U2573 (N_2573,N_2337,N_2268);
xor U2574 (N_2574,N_2194,N_2365);
xnor U2575 (N_2575,N_2034,N_2015);
nor U2576 (N_2576,N_2171,N_2037);
xnor U2577 (N_2577,N_2131,N_2077);
or U2578 (N_2578,N_2453,N_2011);
xor U2579 (N_2579,N_2286,N_2397);
and U2580 (N_2580,N_2452,N_2446);
nor U2581 (N_2581,N_2098,N_2080);
nand U2582 (N_2582,N_2321,N_2313);
or U2583 (N_2583,N_2099,N_2343);
and U2584 (N_2584,N_2315,N_2415);
and U2585 (N_2585,N_2200,N_2406);
nor U2586 (N_2586,N_2206,N_2151);
xor U2587 (N_2587,N_2455,N_2090);
nand U2588 (N_2588,N_2126,N_2023);
nor U2589 (N_2589,N_2130,N_2053);
and U2590 (N_2590,N_2058,N_2169);
xor U2591 (N_2591,N_2438,N_2196);
or U2592 (N_2592,N_2324,N_2102);
and U2593 (N_2593,N_2426,N_2172);
and U2594 (N_2594,N_2233,N_2057);
and U2595 (N_2595,N_2314,N_2457);
xnor U2596 (N_2596,N_2199,N_2409);
nand U2597 (N_2597,N_2072,N_2156);
and U2598 (N_2598,N_2484,N_2479);
and U2599 (N_2599,N_2003,N_2084);
and U2600 (N_2600,N_2394,N_2208);
nor U2601 (N_2601,N_2344,N_2049);
nor U2602 (N_2602,N_2279,N_2209);
nor U2603 (N_2603,N_2191,N_2442);
xor U2604 (N_2604,N_2471,N_2261);
nand U2605 (N_2605,N_2375,N_2245);
and U2606 (N_2606,N_2180,N_2222);
nor U2607 (N_2607,N_2142,N_2121);
nand U2608 (N_2608,N_2012,N_2148);
nand U2609 (N_2609,N_2019,N_2377);
nand U2610 (N_2610,N_2282,N_2138);
nand U2611 (N_2611,N_2486,N_2149);
or U2612 (N_2612,N_2062,N_2292);
xor U2613 (N_2613,N_2462,N_2348);
nand U2614 (N_2614,N_2434,N_2133);
or U2615 (N_2615,N_2340,N_2193);
and U2616 (N_2616,N_2152,N_2316);
nand U2617 (N_2617,N_2161,N_2000);
and U2618 (N_2618,N_2311,N_2384);
nor U2619 (N_2619,N_2215,N_2410);
xnor U2620 (N_2620,N_2256,N_2398);
nor U2621 (N_2621,N_2122,N_2082);
xnor U2622 (N_2622,N_2239,N_2145);
and U2623 (N_2623,N_2361,N_2001);
xnor U2624 (N_2624,N_2094,N_2181);
nor U2625 (N_2625,N_2070,N_2396);
or U2626 (N_2626,N_2028,N_2228);
and U2627 (N_2627,N_2056,N_2364);
nor U2628 (N_2628,N_2356,N_2225);
nor U2629 (N_2629,N_2157,N_2262);
and U2630 (N_2630,N_2002,N_2416);
or U2631 (N_2631,N_2010,N_2413);
xor U2632 (N_2632,N_2088,N_2493);
nor U2633 (N_2633,N_2259,N_2437);
nand U2634 (N_2634,N_2078,N_2432);
nor U2635 (N_2635,N_2238,N_2043);
or U2636 (N_2636,N_2291,N_2289);
and U2637 (N_2637,N_2388,N_2221);
xor U2638 (N_2638,N_2411,N_2497);
or U2639 (N_2639,N_2063,N_2272);
or U2640 (N_2640,N_2459,N_2269);
nor U2641 (N_2641,N_2376,N_2499);
and U2642 (N_2642,N_2490,N_2280);
nand U2643 (N_2643,N_2472,N_2052);
xor U2644 (N_2644,N_2296,N_2247);
xnor U2645 (N_2645,N_2212,N_2183);
nor U2646 (N_2646,N_2127,N_2105);
xnor U2647 (N_2647,N_2489,N_2125);
xor U2648 (N_2648,N_2124,N_2065);
or U2649 (N_2649,N_2230,N_2205);
nand U2650 (N_2650,N_2083,N_2213);
nand U2651 (N_2651,N_2302,N_2383);
nand U2652 (N_2652,N_2162,N_2270);
and U2653 (N_2653,N_2326,N_2170);
and U2654 (N_2654,N_2301,N_2422);
nor U2655 (N_2655,N_2389,N_2460);
or U2656 (N_2656,N_2109,N_2320);
and U2657 (N_2657,N_2190,N_2069);
nand U2658 (N_2658,N_2345,N_2166);
and U2659 (N_2659,N_2425,N_2436);
xor U2660 (N_2660,N_2342,N_2064);
or U2661 (N_2661,N_2407,N_2155);
xor U2662 (N_2662,N_2435,N_2026);
or U2663 (N_2663,N_2006,N_2277);
nand U2664 (N_2664,N_2379,N_2018);
or U2665 (N_2665,N_2231,N_2227);
or U2666 (N_2666,N_2431,N_2267);
and U2667 (N_2667,N_2086,N_2456);
nand U2668 (N_2668,N_2333,N_2469);
nor U2669 (N_2669,N_2117,N_2240);
or U2670 (N_2670,N_2059,N_2176);
nor U2671 (N_2671,N_2232,N_2119);
nand U2672 (N_2672,N_2305,N_2048);
nand U2673 (N_2673,N_2441,N_2309);
and U2674 (N_2674,N_2260,N_2444);
or U2675 (N_2675,N_2184,N_2068);
nor U2676 (N_2676,N_2129,N_2367);
xnor U2677 (N_2677,N_2252,N_2236);
nand U2678 (N_2678,N_2115,N_2287);
and U2679 (N_2679,N_2418,N_2381);
and U2680 (N_2680,N_2331,N_2187);
nand U2681 (N_2681,N_2207,N_2347);
and U2682 (N_2682,N_2031,N_2241);
xnor U2683 (N_2683,N_2100,N_2029);
nor U2684 (N_2684,N_2350,N_2402);
xor U2685 (N_2685,N_2185,N_2104);
or U2686 (N_2686,N_2036,N_2136);
and U2687 (N_2687,N_2308,N_2224);
and U2688 (N_2688,N_2467,N_2022);
nand U2689 (N_2689,N_2294,N_2237);
nand U2690 (N_2690,N_2443,N_2146);
nor U2691 (N_2691,N_2251,N_2328);
nor U2692 (N_2692,N_2370,N_2135);
and U2693 (N_2693,N_2203,N_2414);
nand U2694 (N_2694,N_2440,N_2276);
and U2695 (N_2695,N_2346,N_2123);
nor U2696 (N_2696,N_2352,N_2374);
and U2697 (N_2697,N_2097,N_2243);
or U2698 (N_2698,N_2263,N_2363);
nand U2699 (N_2699,N_2330,N_2366);
and U2700 (N_2700,N_2312,N_2336);
nor U2701 (N_2701,N_2118,N_2378);
or U2702 (N_2702,N_2448,N_2110);
nor U2703 (N_2703,N_2466,N_2380);
xnor U2704 (N_2704,N_2362,N_2424);
or U2705 (N_2705,N_2216,N_2235);
nor U2706 (N_2706,N_2246,N_2385);
and U2707 (N_2707,N_2075,N_2451);
xor U2708 (N_2708,N_2218,N_2103);
or U2709 (N_2709,N_2478,N_2154);
or U2710 (N_2710,N_2060,N_2278);
nor U2711 (N_2711,N_2160,N_2168);
nor U2712 (N_2712,N_2271,N_2400);
nand U2713 (N_2713,N_2035,N_2141);
or U2714 (N_2714,N_2427,N_2210);
nor U2715 (N_2715,N_2491,N_2114);
nand U2716 (N_2716,N_2477,N_2419);
and U2717 (N_2717,N_2498,N_2045);
and U2718 (N_2718,N_2195,N_2433);
and U2719 (N_2719,N_2250,N_2474);
or U2720 (N_2720,N_2143,N_2005);
and U2721 (N_2721,N_2358,N_2335);
and U2722 (N_2722,N_2085,N_2488);
xor U2723 (N_2723,N_2461,N_2420);
nor U2724 (N_2724,N_2044,N_2189);
and U2725 (N_2725,N_2404,N_2128);
nor U2726 (N_2726,N_2112,N_2178);
nor U2727 (N_2727,N_2039,N_2249);
and U2728 (N_2728,N_2025,N_2144);
xnor U2729 (N_2729,N_2423,N_2040);
nor U2730 (N_2730,N_2429,N_2325);
nor U2731 (N_2731,N_2008,N_2303);
xnor U2732 (N_2732,N_2046,N_2050);
and U2733 (N_2733,N_2091,N_2158);
nor U2734 (N_2734,N_2167,N_2487);
and U2735 (N_2735,N_2475,N_2265);
and U2736 (N_2736,N_2360,N_2254);
xor U2737 (N_2737,N_2399,N_2359);
nand U2738 (N_2738,N_2217,N_2332);
xor U2739 (N_2739,N_2405,N_2284);
and U2740 (N_2740,N_2253,N_2283);
xnor U2741 (N_2741,N_2382,N_2116);
or U2742 (N_2742,N_2476,N_2164);
nand U2743 (N_2743,N_2192,N_2009);
xor U2744 (N_2744,N_2485,N_2137);
nand U2745 (N_2745,N_2113,N_2198);
or U2746 (N_2746,N_2248,N_2300);
nand U2747 (N_2747,N_2273,N_2430);
nand U2748 (N_2748,N_2310,N_2211);
or U2749 (N_2749,N_2201,N_2255);
and U2750 (N_2750,N_2376,N_2207);
nor U2751 (N_2751,N_2364,N_2445);
xnor U2752 (N_2752,N_2207,N_2081);
xnor U2753 (N_2753,N_2357,N_2345);
or U2754 (N_2754,N_2196,N_2298);
nand U2755 (N_2755,N_2049,N_2333);
or U2756 (N_2756,N_2156,N_2063);
nand U2757 (N_2757,N_2151,N_2049);
or U2758 (N_2758,N_2493,N_2295);
or U2759 (N_2759,N_2078,N_2255);
and U2760 (N_2760,N_2068,N_2153);
nand U2761 (N_2761,N_2332,N_2166);
xor U2762 (N_2762,N_2132,N_2313);
and U2763 (N_2763,N_2421,N_2151);
nand U2764 (N_2764,N_2046,N_2386);
and U2765 (N_2765,N_2007,N_2182);
nand U2766 (N_2766,N_2328,N_2420);
nand U2767 (N_2767,N_2474,N_2221);
xor U2768 (N_2768,N_2172,N_2143);
and U2769 (N_2769,N_2153,N_2044);
xnor U2770 (N_2770,N_2144,N_2032);
nor U2771 (N_2771,N_2016,N_2057);
or U2772 (N_2772,N_2066,N_2137);
xor U2773 (N_2773,N_2140,N_2302);
nand U2774 (N_2774,N_2473,N_2314);
or U2775 (N_2775,N_2325,N_2029);
or U2776 (N_2776,N_2304,N_2460);
nand U2777 (N_2777,N_2433,N_2007);
xor U2778 (N_2778,N_2175,N_2022);
or U2779 (N_2779,N_2491,N_2460);
xnor U2780 (N_2780,N_2036,N_2022);
and U2781 (N_2781,N_2174,N_2372);
or U2782 (N_2782,N_2482,N_2251);
nor U2783 (N_2783,N_2173,N_2058);
and U2784 (N_2784,N_2466,N_2209);
and U2785 (N_2785,N_2423,N_2333);
and U2786 (N_2786,N_2233,N_2400);
nand U2787 (N_2787,N_2039,N_2230);
or U2788 (N_2788,N_2436,N_2495);
or U2789 (N_2789,N_2235,N_2375);
xnor U2790 (N_2790,N_2423,N_2009);
xnor U2791 (N_2791,N_2167,N_2032);
or U2792 (N_2792,N_2333,N_2370);
or U2793 (N_2793,N_2182,N_2062);
or U2794 (N_2794,N_2343,N_2489);
or U2795 (N_2795,N_2173,N_2240);
or U2796 (N_2796,N_2196,N_2481);
xnor U2797 (N_2797,N_2186,N_2293);
nand U2798 (N_2798,N_2445,N_2349);
xnor U2799 (N_2799,N_2069,N_2106);
and U2800 (N_2800,N_2125,N_2083);
nand U2801 (N_2801,N_2093,N_2382);
xnor U2802 (N_2802,N_2058,N_2458);
xor U2803 (N_2803,N_2169,N_2176);
or U2804 (N_2804,N_2257,N_2433);
or U2805 (N_2805,N_2014,N_2433);
nor U2806 (N_2806,N_2303,N_2451);
nor U2807 (N_2807,N_2067,N_2386);
nand U2808 (N_2808,N_2204,N_2089);
or U2809 (N_2809,N_2365,N_2034);
and U2810 (N_2810,N_2244,N_2007);
nor U2811 (N_2811,N_2182,N_2231);
nand U2812 (N_2812,N_2338,N_2057);
and U2813 (N_2813,N_2134,N_2265);
nand U2814 (N_2814,N_2460,N_2285);
nor U2815 (N_2815,N_2337,N_2157);
and U2816 (N_2816,N_2312,N_2196);
or U2817 (N_2817,N_2360,N_2150);
and U2818 (N_2818,N_2321,N_2402);
xor U2819 (N_2819,N_2356,N_2354);
xor U2820 (N_2820,N_2360,N_2395);
or U2821 (N_2821,N_2226,N_2067);
xnor U2822 (N_2822,N_2472,N_2360);
and U2823 (N_2823,N_2290,N_2285);
xor U2824 (N_2824,N_2037,N_2352);
nor U2825 (N_2825,N_2301,N_2195);
xnor U2826 (N_2826,N_2443,N_2400);
and U2827 (N_2827,N_2354,N_2222);
nand U2828 (N_2828,N_2042,N_2380);
nand U2829 (N_2829,N_2388,N_2277);
and U2830 (N_2830,N_2036,N_2041);
and U2831 (N_2831,N_2245,N_2113);
or U2832 (N_2832,N_2098,N_2263);
nand U2833 (N_2833,N_2382,N_2027);
nand U2834 (N_2834,N_2241,N_2237);
xor U2835 (N_2835,N_2153,N_2122);
nor U2836 (N_2836,N_2457,N_2330);
or U2837 (N_2837,N_2402,N_2482);
and U2838 (N_2838,N_2127,N_2317);
nand U2839 (N_2839,N_2344,N_2032);
xor U2840 (N_2840,N_2324,N_2489);
or U2841 (N_2841,N_2299,N_2057);
and U2842 (N_2842,N_2103,N_2256);
nor U2843 (N_2843,N_2200,N_2441);
or U2844 (N_2844,N_2497,N_2368);
xor U2845 (N_2845,N_2414,N_2280);
or U2846 (N_2846,N_2471,N_2370);
and U2847 (N_2847,N_2478,N_2094);
and U2848 (N_2848,N_2290,N_2414);
or U2849 (N_2849,N_2103,N_2127);
or U2850 (N_2850,N_2066,N_2007);
or U2851 (N_2851,N_2180,N_2273);
nor U2852 (N_2852,N_2181,N_2160);
or U2853 (N_2853,N_2192,N_2185);
nor U2854 (N_2854,N_2482,N_2255);
or U2855 (N_2855,N_2140,N_2024);
xor U2856 (N_2856,N_2201,N_2039);
nand U2857 (N_2857,N_2440,N_2485);
and U2858 (N_2858,N_2129,N_2441);
nor U2859 (N_2859,N_2476,N_2253);
and U2860 (N_2860,N_2448,N_2099);
nand U2861 (N_2861,N_2052,N_2268);
nand U2862 (N_2862,N_2444,N_2096);
nand U2863 (N_2863,N_2373,N_2047);
xor U2864 (N_2864,N_2164,N_2203);
xor U2865 (N_2865,N_2076,N_2016);
or U2866 (N_2866,N_2215,N_2243);
nor U2867 (N_2867,N_2219,N_2019);
nand U2868 (N_2868,N_2329,N_2129);
nor U2869 (N_2869,N_2470,N_2083);
nand U2870 (N_2870,N_2455,N_2204);
nand U2871 (N_2871,N_2202,N_2057);
xor U2872 (N_2872,N_2434,N_2018);
or U2873 (N_2873,N_2479,N_2011);
nand U2874 (N_2874,N_2464,N_2051);
nand U2875 (N_2875,N_2119,N_2021);
nand U2876 (N_2876,N_2246,N_2264);
nand U2877 (N_2877,N_2181,N_2226);
or U2878 (N_2878,N_2103,N_2101);
and U2879 (N_2879,N_2366,N_2253);
or U2880 (N_2880,N_2246,N_2392);
nor U2881 (N_2881,N_2283,N_2421);
and U2882 (N_2882,N_2477,N_2467);
nor U2883 (N_2883,N_2245,N_2496);
nor U2884 (N_2884,N_2029,N_2383);
nand U2885 (N_2885,N_2132,N_2077);
and U2886 (N_2886,N_2194,N_2142);
xnor U2887 (N_2887,N_2114,N_2444);
nor U2888 (N_2888,N_2175,N_2094);
nand U2889 (N_2889,N_2295,N_2021);
xor U2890 (N_2890,N_2205,N_2454);
nand U2891 (N_2891,N_2073,N_2334);
nor U2892 (N_2892,N_2413,N_2361);
nand U2893 (N_2893,N_2137,N_2075);
nor U2894 (N_2894,N_2018,N_2004);
nor U2895 (N_2895,N_2305,N_2112);
or U2896 (N_2896,N_2425,N_2491);
and U2897 (N_2897,N_2237,N_2105);
or U2898 (N_2898,N_2483,N_2036);
nor U2899 (N_2899,N_2032,N_2355);
and U2900 (N_2900,N_2476,N_2029);
and U2901 (N_2901,N_2229,N_2071);
or U2902 (N_2902,N_2253,N_2351);
or U2903 (N_2903,N_2134,N_2443);
and U2904 (N_2904,N_2169,N_2117);
xor U2905 (N_2905,N_2154,N_2406);
xor U2906 (N_2906,N_2469,N_2183);
nand U2907 (N_2907,N_2000,N_2038);
xor U2908 (N_2908,N_2369,N_2072);
and U2909 (N_2909,N_2366,N_2020);
xor U2910 (N_2910,N_2302,N_2272);
or U2911 (N_2911,N_2238,N_2414);
nand U2912 (N_2912,N_2307,N_2058);
nand U2913 (N_2913,N_2048,N_2121);
nand U2914 (N_2914,N_2492,N_2371);
nand U2915 (N_2915,N_2365,N_2139);
nor U2916 (N_2916,N_2282,N_2035);
and U2917 (N_2917,N_2416,N_2485);
xnor U2918 (N_2918,N_2117,N_2064);
and U2919 (N_2919,N_2433,N_2125);
nor U2920 (N_2920,N_2155,N_2153);
nor U2921 (N_2921,N_2386,N_2251);
or U2922 (N_2922,N_2120,N_2309);
xor U2923 (N_2923,N_2477,N_2246);
nor U2924 (N_2924,N_2494,N_2024);
or U2925 (N_2925,N_2447,N_2327);
xor U2926 (N_2926,N_2394,N_2081);
nor U2927 (N_2927,N_2413,N_2461);
xnor U2928 (N_2928,N_2247,N_2435);
xor U2929 (N_2929,N_2273,N_2256);
xor U2930 (N_2930,N_2468,N_2300);
or U2931 (N_2931,N_2186,N_2363);
or U2932 (N_2932,N_2113,N_2038);
nor U2933 (N_2933,N_2018,N_2390);
nor U2934 (N_2934,N_2056,N_2492);
nor U2935 (N_2935,N_2210,N_2384);
and U2936 (N_2936,N_2181,N_2496);
nand U2937 (N_2937,N_2154,N_2178);
nand U2938 (N_2938,N_2008,N_2442);
and U2939 (N_2939,N_2071,N_2273);
and U2940 (N_2940,N_2291,N_2491);
nor U2941 (N_2941,N_2049,N_2108);
and U2942 (N_2942,N_2424,N_2046);
nor U2943 (N_2943,N_2380,N_2481);
xnor U2944 (N_2944,N_2050,N_2249);
or U2945 (N_2945,N_2494,N_2204);
or U2946 (N_2946,N_2488,N_2382);
and U2947 (N_2947,N_2416,N_2139);
or U2948 (N_2948,N_2095,N_2428);
or U2949 (N_2949,N_2371,N_2381);
and U2950 (N_2950,N_2364,N_2044);
nand U2951 (N_2951,N_2308,N_2032);
nand U2952 (N_2952,N_2311,N_2048);
nand U2953 (N_2953,N_2446,N_2289);
nor U2954 (N_2954,N_2259,N_2153);
xor U2955 (N_2955,N_2174,N_2064);
nor U2956 (N_2956,N_2382,N_2067);
nand U2957 (N_2957,N_2382,N_2392);
nand U2958 (N_2958,N_2147,N_2474);
nand U2959 (N_2959,N_2387,N_2196);
nor U2960 (N_2960,N_2096,N_2192);
xor U2961 (N_2961,N_2040,N_2226);
nor U2962 (N_2962,N_2430,N_2058);
and U2963 (N_2963,N_2177,N_2010);
xor U2964 (N_2964,N_2069,N_2141);
nor U2965 (N_2965,N_2081,N_2003);
and U2966 (N_2966,N_2075,N_2454);
xnor U2967 (N_2967,N_2146,N_2181);
xnor U2968 (N_2968,N_2231,N_2194);
xnor U2969 (N_2969,N_2099,N_2490);
and U2970 (N_2970,N_2240,N_2370);
xor U2971 (N_2971,N_2097,N_2452);
xor U2972 (N_2972,N_2181,N_2084);
nor U2973 (N_2973,N_2434,N_2181);
or U2974 (N_2974,N_2495,N_2015);
xor U2975 (N_2975,N_2485,N_2262);
xnor U2976 (N_2976,N_2485,N_2267);
nand U2977 (N_2977,N_2318,N_2195);
nand U2978 (N_2978,N_2055,N_2283);
xnor U2979 (N_2979,N_2192,N_2099);
and U2980 (N_2980,N_2436,N_2230);
nand U2981 (N_2981,N_2172,N_2445);
and U2982 (N_2982,N_2427,N_2063);
xor U2983 (N_2983,N_2441,N_2319);
and U2984 (N_2984,N_2490,N_2159);
nand U2985 (N_2985,N_2049,N_2309);
nor U2986 (N_2986,N_2428,N_2442);
xnor U2987 (N_2987,N_2264,N_2356);
or U2988 (N_2988,N_2430,N_2380);
xor U2989 (N_2989,N_2055,N_2312);
and U2990 (N_2990,N_2259,N_2326);
and U2991 (N_2991,N_2126,N_2365);
xnor U2992 (N_2992,N_2400,N_2379);
or U2993 (N_2993,N_2206,N_2480);
xor U2994 (N_2994,N_2485,N_2322);
and U2995 (N_2995,N_2221,N_2214);
nor U2996 (N_2996,N_2323,N_2069);
and U2997 (N_2997,N_2277,N_2230);
xnor U2998 (N_2998,N_2494,N_2207);
nand U2999 (N_2999,N_2187,N_2086);
and U3000 (N_3000,N_2549,N_2853);
or U3001 (N_3001,N_2662,N_2629);
nor U3002 (N_3002,N_2664,N_2537);
and U3003 (N_3003,N_2739,N_2598);
xnor U3004 (N_3004,N_2890,N_2733);
or U3005 (N_3005,N_2951,N_2746);
nor U3006 (N_3006,N_2904,N_2894);
nand U3007 (N_3007,N_2703,N_2886);
and U3008 (N_3008,N_2609,N_2881);
nand U3009 (N_3009,N_2658,N_2837);
nor U3010 (N_3010,N_2657,N_2965);
or U3011 (N_3011,N_2915,N_2942);
and U3012 (N_3012,N_2758,N_2948);
nand U3013 (N_3013,N_2668,N_2999);
nor U3014 (N_3014,N_2763,N_2792);
xor U3015 (N_3015,N_2954,N_2719);
nor U3016 (N_3016,N_2632,N_2995);
or U3017 (N_3017,N_2591,N_2568);
nand U3018 (N_3018,N_2585,N_2626);
nand U3019 (N_3019,N_2876,N_2829);
or U3020 (N_3020,N_2927,N_2660);
and U3021 (N_3021,N_2516,N_2822);
nor U3022 (N_3022,N_2742,N_2912);
and U3023 (N_3023,N_2646,N_2956);
nor U3024 (N_3024,N_2860,N_2540);
or U3025 (N_3025,N_2985,N_2637);
and U3026 (N_3026,N_2774,N_2892);
nor U3027 (N_3027,N_2762,N_2922);
and U3028 (N_3028,N_2541,N_2771);
or U3029 (N_3029,N_2652,N_2882);
nor U3030 (N_3030,N_2845,N_2712);
xor U3031 (N_3031,N_2640,N_2786);
nor U3032 (N_3032,N_2799,N_2911);
nand U3033 (N_3033,N_2982,N_2789);
xor U3034 (N_3034,N_2548,N_2615);
or U3035 (N_3035,N_2717,N_2914);
xor U3036 (N_3036,N_2984,N_2744);
nand U3037 (N_3037,N_2694,N_2800);
xnor U3038 (N_3038,N_2749,N_2899);
nor U3039 (N_3039,N_2950,N_2913);
and U3040 (N_3040,N_2817,N_2634);
xnor U3041 (N_3041,N_2543,N_2674);
and U3042 (N_3042,N_2700,N_2811);
nand U3043 (N_3043,N_2635,N_2716);
nor U3044 (N_3044,N_2610,N_2940);
or U3045 (N_3045,N_2967,N_2961);
and U3046 (N_3046,N_2679,N_2697);
nor U3047 (N_3047,N_2692,N_2907);
nor U3048 (N_3048,N_2530,N_2727);
nor U3049 (N_3049,N_2592,N_2975);
nor U3050 (N_3050,N_2848,N_2636);
nand U3051 (N_3051,N_2520,N_2849);
and U3052 (N_3052,N_2676,N_2900);
xnor U3053 (N_3053,N_2823,N_2870);
nor U3054 (N_3054,N_2843,N_2600);
and U3055 (N_3055,N_2624,N_2879);
or U3056 (N_3056,N_2695,N_2671);
nand U3057 (N_3057,N_2866,N_2651);
xor U3058 (N_3058,N_2526,N_2846);
xnor U3059 (N_3059,N_2693,N_2937);
nor U3060 (N_3060,N_2794,N_2593);
nor U3061 (N_3061,N_2734,N_2648);
xor U3062 (N_3062,N_2989,N_2687);
nor U3063 (N_3063,N_2723,N_2562);
and U3064 (N_3064,N_2683,N_2514);
and U3065 (N_3065,N_2711,N_2839);
nand U3066 (N_3066,N_2567,N_2542);
nand U3067 (N_3067,N_2770,N_2945);
xor U3068 (N_3068,N_2825,N_2536);
and U3069 (N_3069,N_2602,N_2828);
nor U3070 (N_3070,N_2990,N_2737);
xor U3071 (N_3071,N_2873,N_2962);
nand U3072 (N_3072,N_2670,N_2788);
xnor U3073 (N_3073,N_2643,N_2960);
or U3074 (N_3074,N_2747,N_2628);
xor U3075 (N_3075,N_2709,N_2986);
nand U3076 (N_3076,N_2906,N_2896);
nor U3077 (N_3077,N_2686,N_2688);
or U3078 (N_3078,N_2889,N_2519);
or U3079 (N_3079,N_2966,N_2745);
or U3080 (N_3080,N_2813,N_2597);
and U3081 (N_3081,N_2752,N_2809);
nand U3082 (N_3082,N_2714,N_2805);
nand U3083 (N_3083,N_2659,N_2777);
nand U3084 (N_3084,N_2521,N_2645);
and U3085 (N_3085,N_2833,N_2509);
and U3086 (N_3086,N_2768,N_2702);
xor U3087 (N_3087,N_2618,N_2773);
nand U3088 (N_3088,N_2623,N_2827);
nor U3089 (N_3089,N_2832,N_2769);
nand U3090 (N_3090,N_2826,N_2836);
or U3091 (N_3091,N_2563,N_2844);
or U3092 (N_3092,N_2528,N_2955);
and U3093 (N_3093,N_2917,N_2798);
xnor U3094 (N_3094,N_2724,N_2754);
nor U3095 (N_3095,N_2755,N_2925);
and U3096 (N_3096,N_2790,N_2880);
and U3097 (N_3097,N_2994,N_2554);
or U3098 (N_3098,N_2958,N_2920);
xor U3099 (N_3099,N_2731,N_2617);
xnor U3100 (N_3100,N_2564,N_2667);
and U3101 (N_3101,N_2572,N_2550);
nor U3102 (N_3102,N_2863,N_2620);
or U3103 (N_3103,N_2625,N_2932);
and U3104 (N_3104,N_2685,N_2582);
and U3105 (N_3105,N_2533,N_2614);
or U3106 (N_3106,N_2689,N_2748);
or U3107 (N_3107,N_2997,N_2782);
nor U3108 (N_3108,N_2513,N_2574);
nor U3109 (N_3109,N_2797,N_2921);
xnor U3110 (N_3110,N_2661,N_2976);
xor U3111 (N_3111,N_2633,N_2583);
nor U3112 (N_3112,N_2715,N_2783);
xor U3113 (N_3113,N_2547,N_2840);
nor U3114 (N_3114,N_2611,N_2818);
or U3115 (N_3115,N_2808,N_2918);
and U3116 (N_3116,N_2729,N_2964);
nor U3117 (N_3117,N_2761,N_2518);
and U3118 (N_3118,N_2577,N_2713);
and U3119 (N_3119,N_2728,N_2772);
nor U3120 (N_3120,N_2857,N_2622);
nor U3121 (N_3121,N_2814,N_2968);
and U3122 (N_3122,N_2802,N_2821);
nand U3123 (N_3123,N_2963,N_2517);
xor U3124 (N_3124,N_2561,N_2505);
nor U3125 (N_3125,N_2696,N_2718);
and U3126 (N_3126,N_2998,N_2656);
and U3127 (N_3127,N_2551,N_2952);
or U3128 (N_3128,N_2861,N_2938);
nor U3129 (N_3129,N_2501,N_2949);
xnor U3130 (N_3130,N_2902,N_2793);
and U3131 (N_3131,N_2581,N_2690);
or U3132 (N_3132,N_2515,N_2673);
nor U3133 (N_3133,N_2936,N_2887);
nor U3134 (N_3134,N_2874,N_2767);
xnor U3135 (N_3135,N_2803,N_2511);
xor U3136 (N_3136,N_2534,N_2820);
or U3137 (N_3137,N_2557,N_2862);
nor U3138 (N_3138,N_2981,N_2590);
nor U3139 (N_3139,N_2531,N_2571);
xor U3140 (N_3140,N_2750,N_2864);
nand U3141 (N_3141,N_2850,N_2831);
xor U3142 (N_3142,N_2791,N_2573);
nor U3143 (N_3143,N_2738,N_2684);
nor U3144 (N_3144,N_2710,N_2926);
or U3145 (N_3145,N_2875,N_2638);
or U3146 (N_3146,N_2779,N_2720);
nor U3147 (N_3147,N_2556,N_2631);
and U3148 (N_3148,N_2895,N_2512);
or U3149 (N_3149,N_2835,N_2604);
xnor U3150 (N_3150,N_2705,N_2878);
nand U3151 (N_3151,N_2957,N_2898);
nor U3152 (N_3152,N_2947,N_2816);
or U3153 (N_3153,N_2586,N_2877);
xor U3154 (N_3154,N_2871,N_2740);
or U3155 (N_3155,N_2678,N_2991);
xor U3156 (N_3156,N_2854,N_2672);
or U3157 (N_3157,N_2570,N_2939);
nand U3158 (N_3158,N_2812,N_2544);
nand U3159 (N_3159,N_2579,N_2741);
or U3160 (N_3160,N_2508,N_2775);
nand U3161 (N_3161,N_2653,N_2819);
or U3162 (N_3162,N_2919,N_2677);
or U3163 (N_3163,N_2580,N_2841);
xnor U3164 (N_3164,N_2980,N_2959);
nor U3165 (N_3165,N_2650,N_2996);
or U3166 (N_3166,N_2905,N_2972);
nand U3167 (N_3167,N_2759,N_2566);
nand U3168 (N_3168,N_2977,N_2893);
nand U3169 (N_3169,N_2736,N_2644);
and U3170 (N_3170,N_2507,N_2974);
nor U3171 (N_3171,N_2613,N_2934);
and U3172 (N_3172,N_2522,N_2612);
nand U3173 (N_3173,N_2647,N_2756);
nor U3174 (N_3174,N_2884,N_2908);
nand U3175 (N_3175,N_2654,N_2560);
or U3176 (N_3176,N_2606,N_2524);
or U3177 (N_3177,N_2847,N_2834);
and U3178 (N_3178,N_2682,N_2663);
nand U3179 (N_3179,N_2764,N_2859);
and U3180 (N_3180,N_2732,N_2642);
and U3181 (N_3181,N_2675,N_2933);
nor U3182 (N_3182,N_2796,N_2973);
nand U3183 (N_3183,N_2891,N_2584);
nor U3184 (N_3184,N_2680,N_2924);
nor U3185 (N_3185,N_2681,N_2901);
and U3186 (N_3186,N_2721,N_2838);
and U3187 (N_3187,N_2869,N_2807);
nor U3188 (N_3188,N_2706,N_2776);
nor U3189 (N_3189,N_2970,N_2855);
and U3190 (N_3190,N_2503,N_2559);
xor U3191 (N_3191,N_2795,N_2743);
nor U3192 (N_3192,N_2824,N_2804);
and U3193 (N_3193,N_2785,N_2842);
and U3194 (N_3194,N_2669,N_2558);
nor U3195 (N_3195,N_2931,N_2510);
nor U3196 (N_3196,N_2865,N_2532);
and U3197 (N_3197,N_2897,N_2529);
or U3198 (N_3198,N_2766,N_2704);
nor U3199 (N_3199,N_2701,N_2500);
xor U3200 (N_3200,N_2988,N_2993);
nor U3201 (N_3201,N_2888,N_2971);
or U3202 (N_3202,N_2607,N_2923);
or U3203 (N_3203,N_2753,N_2929);
nor U3204 (N_3204,N_2730,N_2699);
nor U3205 (N_3205,N_2655,N_2851);
nand U3206 (N_3206,N_2608,N_2596);
nand U3207 (N_3207,N_2760,N_2555);
or U3208 (N_3208,N_2916,N_2603);
nand U3209 (N_3209,N_2801,N_2641);
and U3210 (N_3210,N_2539,N_2757);
and U3211 (N_3211,N_2969,N_2616);
nand U3212 (N_3212,N_2502,N_2525);
xor U3213 (N_3213,N_2725,N_2504);
xor U3214 (N_3214,N_2806,N_2930);
and U3215 (N_3215,N_2953,N_2944);
or U3216 (N_3216,N_2992,N_2872);
nor U3217 (N_3217,N_2605,N_2665);
xnor U3218 (N_3218,N_2858,N_2639);
or U3219 (N_3219,N_2576,N_2552);
nor U3220 (N_3220,N_2781,N_2852);
nor U3221 (N_3221,N_2538,N_2707);
and U3222 (N_3222,N_2726,N_2868);
nor U3223 (N_3223,N_2778,N_2780);
xnor U3224 (N_3224,N_2885,N_2627);
or U3225 (N_3225,N_2594,N_2708);
xor U3226 (N_3226,N_2527,N_2978);
nor U3227 (N_3227,N_2979,N_2935);
xor U3228 (N_3228,N_2546,N_2523);
nor U3229 (N_3229,N_2928,N_2784);
or U3230 (N_3230,N_2751,N_2565);
and U3231 (N_3231,N_2588,N_2630);
nor U3232 (N_3232,N_2946,N_2649);
nand U3233 (N_3233,N_2589,N_2578);
nor U3234 (N_3234,N_2910,N_2810);
or U3235 (N_3235,N_2903,N_2815);
and U3236 (N_3236,N_2666,N_2575);
nor U3237 (N_3237,N_2621,N_2735);
nand U3238 (N_3238,N_2983,N_2553);
and U3239 (N_3239,N_2595,N_2722);
nor U3240 (N_3240,N_2601,N_2535);
xnor U3241 (N_3241,N_2943,N_2941);
nor U3242 (N_3242,N_2787,N_2883);
and U3243 (N_3243,N_2691,N_2909);
or U3244 (N_3244,N_2830,N_2856);
nor U3245 (N_3245,N_2987,N_2569);
or U3246 (N_3246,N_2506,N_2765);
or U3247 (N_3247,N_2867,N_2619);
or U3248 (N_3248,N_2587,N_2545);
nand U3249 (N_3249,N_2698,N_2599);
and U3250 (N_3250,N_2578,N_2918);
nand U3251 (N_3251,N_2939,N_2739);
and U3252 (N_3252,N_2501,N_2670);
xor U3253 (N_3253,N_2943,N_2881);
xnor U3254 (N_3254,N_2855,N_2814);
or U3255 (N_3255,N_2899,N_2577);
nand U3256 (N_3256,N_2675,N_2527);
nand U3257 (N_3257,N_2893,N_2537);
nor U3258 (N_3258,N_2896,N_2501);
nand U3259 (N_3259,N_2888,N_2840);
and U3260 (N_3260,N_2959,N_2892);
or U3261 (N_3261,N_2829,N_2711);
and U3262 (N_3262,N_2622,N_2882);
nand U3263 (N_3263,N_2557,N_2732);
xnor U3264 (N_3264,N_2860,N_2563);
and U3265 (N_3265,N_2990,N_2834);
nor U3266 (N_3266,N_2630,N_2946);
or U3267 (N_3267,N_2746,N_2847);
and U3268 (N_3268,N_2654,N_2917);
and U3269 (N_3269,N_2658,N_2554);
or U3270 (N_3270,N_2924,N_2602);
xor U3271 (N_3271,N_2503,N_2980);
nor U3272 (N_3272,N_2520,N_2569);
nor U3273 (N_3273,N_2708,N_2605);
or U3274 (N_3274,N_2660,N_2683);
or U3275 (N_3275,N_2670,N_2746);
nand U3276 (N_3276,N_2877,N_2851);
nor U3277 (N_3277,N_2740,N_2617);
or U3278 (N_3278,N_2594,N_2573);
xor U3279 (N_3279,N_2512,N_2988);
nand U3280 (N_3280,N_2622,N_2787);
xor U3281 (N_3281,N_2562,N_2912);
or U3282 (N_3282,N_2982,N_2816);
and U3283 (N_3283,N_2852,N_2522);
xor U3284 (N_3284,N_2897,N_2969);
nand U3285 (N_3285,N_2999,N_2944);
nor U3286 (N_3286,N_2978,N_2779);
nor U3287 (N_3287,N_2695,N_2637);
xnor U3288 (N_3288,N_2633,N_2933);
or U3289 (N_3289,N_2522,N_2876);
nor U3290 (N_3290,N_2585,N_2509);
or U3291 (N_3291,N_2831,N_2653);
or U3292 (N_3292,N_2940,N_2623);
and U3293 (N_3293,N_2598,N_2829);
nand U3294 (N_3294,N_2757,N_2651);
nor U3295 (N_3295,N_2868,N_2527);
nand U3296 (N_3296,N_2695,N_2912);
and U3297 (N_3297,N_2577,N_2833);
nand U3298 (N_3298,N_2523,N_2601);
and U3299 (N_3299,N_2683,N_2958);
xnor U3300 (N_3300,N_2808,N_2624);
nor U3301 (N_3301,N_2987,N_2676);
xor U3302 (N_3302,N_2800,N_2739);
nor U3303 (N_3303,N_2817,N_2749);
nor U3304 (N_3304,N_2919,N_2539);
or U3305 (N_3305,N_2920,N_2695);
or U3306 (N_3306,N_2745,N_2550);
nor U3307 (N_3307,N_2660,N_2928);
or U3308 (N_3308,N_2513,N_2962);
nor U3309 (N_3309,N_2830,N_2813);
nor U3310 (N_3310,N_2612,N_2671);
and U3311 (N_3311,N_2655,N_2742);
and U3312 (N_3312,N_2752,N_2626);
nor U3313 (N_3313,N_2829,N_2752);
nand U3314 (N_3314,N_2550,N_2721);
xor U3315 (N_3315,N_2553,N_2982);
xnor U3316 (N_3316,N_2837,N_2958);
and U3317 (N_3317,N_2954,N_2640);
nor U3318 (N_3318,N_2845,N_2620);
nand U3319 (N_3319,N_2739,N_2837);
or U3320 (N_3320,N_2502,N_2966);
nand U3321 (N_3321,N_2638,N_2680);
nand U3322 (N_3322,N_2524,N_2571);
or U3323 (N_3323,N_2692,N_2506);
nand U3324 (N_3324,N_2855,N_2845);
nand U3325 (N_3325,N_2501,N_2532);
nand U3326 (N_3326,N_2853,N_2771);
nor U3327 (N_3327,N_2899,N_2886);
xnor U3328 (N_3328,N_2755,N_2918);
or U3329 (N_3329,N_2517,N_2531);
nand U3330 (N_3330,N_2826,N_2889);
nand U3331 (N_3331,N_2720,N_2753);
nand U3332 (N_3332,N_2886,N_2545);
or U3333 (N_3333,N_2740,N_2795);
and U3334 (N_3334,N_2658,N_2678);
nand U3335 (N_3335,N_2629,N_2899);
nor U3336 (N_3336,N_2717,N_2934);
or U3337 (N_3337,N_2507,N_2523);
nor U3338 (N_3338,N_2662,N_2708);
xor U3339 (N_3339,N_2518,N_2940);
or U3340 (N_3340,N_2855,N_2748);
xnor U3341 (N_3341,N_2862,N_2988);
and U3342 (N_3342,N_2570,N_2998);
or U3343 (N_3343,N_2801,N_2661);
nand U3344 (N_3344,N_2804,N_2875);
nor U3345 (N_3345,N_2676,N_2988);
nand U3346 (N_3346,N_2503,N_2775);
and U3347 (N_3347,N_2754,N_2681);
nor U3348 (N_3348,N_2567,N_2701);
nand U3349 (N_3349,N_2509,N_2992);
or U3350 (N_3350,N_2557,N_2692);
nor U3351 (N_3351,N_2712,N_2627);
nor U3352 (N_3352,N_2940,N_2502);
or U3353 (N_3353,N_2896,N_2793);
xnor U3354 (N_3354,N_2856,N_2533);
or U3355 (N_3355,N_2920,N_2562);
or U3356 (N_3356,N_2786,N_2636);
and U3357 (N_3357,N_2730,N_2935);
or U3358 (N_3358,N_2755,N_2965);
and U3359 (N_3359,N_2525,N_2583);
or U3360 (N_3360,N_2972,N_2967);
or U3361 (N_3361,N_2553,N_2987);
xor U3362 (N_3362,N_2643,N_2991);
xnor U3363 (N_3363,N_2977,N_2998);
and U3364 (N_3364,N_2781,N_2788);
xnor U3365 (N_3365,N_2982,N_2786);
and U3366 (N_3366,N_2938,N_2847);
and U3367 (N_3367,N_2915,N_2861);
nor U3368 (N_3368,N_2537,N_2672);
nand U3369 (N_3369,N_2993,N_2822);
nand U3370 (N_3370,N_2507,N_2538);
and U3371 (N_3371,N_2540,N_2786);
nor U3372 (N_3372,N_2750,N_2755);
nand U3373 (N_3373,N_2779,N_2793);
nand U3374 (N_3374,N_2817,N_2810);
xor U3375 (N_3375,N_2830,N_2938);
nor U3376 (N_3376,N_2545,N_2510);
nor U3377 (N_3377,N_2764,N_2653);
or U3378 (N_3378,N_2672,N_2649);
nand U3379 (N_3379,N_2964,N_2947);
and U3380 (N_3380,N_2546,N_2871);
nand U3381 (N_3381,N_2602,N_2616);
or U3382 (N_3382,N_2823,N_2743);
nand U3383 (N_3383,N_2832,N_2830);
or U3384 (N_3384,N_2636,N_2745);
xor U3385 (N_3385,N_2786,N_2677);
nand U3386 (N_3386,N_2581,N_2755);
nor U3387 (N_3387,N_2955,N_2936);
nand U3388 (N_3388,N_2670,N_2838);
and U3389 (N_3389,N_2762,N_2857);
and U3390 (N_3390,N_2913,N_2916);
and U3391 (N_3391,N_2673,N_2684);
nor U3392 (N_3392,N_2658,N_2922);
or U3393 (N_3393,N_2609,N_2559);
xor U3394 (N_3394,N_2886,N_2817);
nand U3395 (N_3395,N_2674,N_2668);
or U3396 (N_3396,N_2601,N_2512);
and U3397 (N_3397,N_2518,N_2632);
nand U3398 (N_3398,N_2916,N_2921);
and U3399 (N_3399,N_2744,N_2597);
xor U3400 (N_3400,N_2914,N_2655);
or U3401 (N_3401,N_2617,N_2631);
nor U3402 (N_3402,N_2773,N_2753);
nor U3403 (N_3403,N_2826,N_2854);
xor U3404 (N_3404,N_2717,N_2978);
xnor U3405 (N_3405,N_2693,N_2879);
xor U3406 (N_3406,N_2775,N_2557);
and U3407 (N_3407,N_2856,N_2773);
nor U3408 (N_3408,N_2577,N_2749);
nor U3409 (N_3409,N_2522,N_2875);
nand U3410 (N_3410,N_2886,N_2544);
and U3411 (N_3411,N_2897,N_2516);
nor U3412 (N_3412,N_2548,N_2920);
and U3413 (N_3413,N_2640,N_2791);
nor U3414 (N_3414,N_2945,N_2737);
and U3415 (N_3415,N_2904,N_2932);
nand U3416 (N_3416,N_2942,N_2595);
xor U3417 (N_3417,N_2533,N_2715);
and U3418 (N_3418,N_2604,N_2745);
nand U3419 (N_3419,N_2703,N_2656);
or U3420 (N_3420,N_2677,N_2885);
nor U3421 (N_3421,N_2517,N_2514);
xnor U3422 (N_3422,N_2722,N_2615);
or U3423 (N_3423,N_2867,N_2520);
nand U3424 (N_3424,N_2980,N_2559);
or U3425 (N_3425,N_2589,N_2981);
or U3426 (N_3426,N_2555,N_2653);
nand U3427 (N_3427,N_2504,N_2613);
or U3428 (N_3428,N_2854,N_2665);
xnor U3429 (N_3429,N_2589,N_2982);
xor U3430 (N_3430,N_2756,N_2708);
nor U3431 (N_3431,N_2693,N_2753);
nor U3432 (N_3432,N_2809,N_2857);
or U3433 (N_3433,N_2918,N_2967);
and U3434 (N_3434,N_2987,N_2812);
and U3435 (N_3435,N_2704,N_2668);
nand U3436 (N_3436,N_2669,N_2519);
and U3437 (N_3437,N_2690,N_2984);
or U3438 (N_3438,N_2589,N_2639);
nor U3439 (N_3439,N_2807,N_2558);
and U3440 (N_3440,N_2804,N_2898);
nor U3441 (N_3441,N_2662,N_2719);
or U3442 (N_3442,N_2979,N_2640);
or U3443 (N_3443,N_2971,N_2566);
xnor U3444 (N_3444,N_2873,N_2887);
nand U3445 (N_3445,N_2721,N_2708);
nor U3446 (N_3446,N_2787,N_2634);
or U3447 (N_3447,N_2513,N_2538);
nor U3448 (N_3448,N_2775,N_2553);
nor U3449 (N_3449,N_2667,N_2595);
nand U3450 (N_3450,N_2805,N_2822);
xnor U3451 (N_3451,N_2596,N_2909);
nand U3452 (N_3452,N_2905,N_2565);
or U3453 (N_3453,N_2746,N_2637);
xnor U3454 (N_3454,N_2850,N_2628);
and U3455 (N_3455,N_2635,N_2922);
xor U3456 (N_3456,N_2969,N_2985);
or U3457 (N_3457,N_2995,N_2918);
nand U3458 (N_3458,N_2688,N_2872);
and U3459 (N_3459,N_2504,N_2998);
and U3460 (N_3460,N_2586,N_2874);
and U3461 (N_3461,N_2511,N_2941);
nor U3462 (N_3462,N_2953,N_2587);
nand U3463 (N_3463,N_2812,N_2888);
nor U3464 (N_3464,N_2864,N_2710);
and U3465 (N_3465,N_2965,N_2945);
or U3466 (N_3466,N_2642,N_2550);
and U3467 (N_3467,N_2877,N_2982);
xor U3468 (N_3468,N_2530,N_2505);
or U3469 (N_3469,N_2906,N_2562);
or U3470 (N_3470,N_2987,N_2932);
or U3471 (N_3471,N_2938,N_2700);
or U3472 (N_3472,N_2727,N_2519);
nand U3473 (N_3473,N_2616,N_2701);
nor U3474 (N_3474,N_2523,N_2879);
nor U3475 (N_3475,N_2984,N_2736);
and U3476 (N_3476,N_2717,N_2621);
and U3477 (N_3477,N_2768,N_2676);
and U3478 (N_3478,N_2632,N_2849);
nand U3479 (N_3479,N_2985,N_2921);
nor U3480 (N_3480,N_2807,N_2863);
and U3481 (N_3481,N_2596,N_2668);
nor U3482 (N_3482,N_2893,N_2632);
and U3483 (N_3483,N_2803,N_2697);
nand U3484 (N_3484,N_2595,N_2614);
nor U3485 (N_3485,N_2893,N_2531);
nand U3486 (N_3486,N_2831,N_2560);
and U3487 (N_3487,N_2575,N_2746);
xnor U3488 (N_3488,N_2716,N_2662);
xor U3489 (N_3489,N_2625,N_2629);
nor U3490 (N_3490,N_2959,N_2835);
nor U3491 (N_3491,N_2838,N_2648);
nor U3492 (N_3492,N_2516,N_2774);
or U3493 (N_3493,N_2682,N_2614);
nand U3494 (N_3494,N_2843,N_2626);
nor U3495 (N_3495,N_2996,N_2613);
xnor U3496 (N_3496,N_2938,N_2655);
xor U3497 (N_3497,N_2768,N_2854);
xnor U3498 (N_3498,N_2976,N_2603);
nor U3499 (N_3499,N_2904,N_2967);
and U3500 (N_3500,N_3434,N_3250);
and U3501 (N_3501,N_3172,N_3084);
nor U3502 (N_3502,N_3159,N_3060);
xnor U3503 (N_3503,N_3321,N_3268);
or U3504 (N_3504,N_3439,N_3028);
and U3505 (N_3505,N_3129,N_3251);
nand U3506 (N_3506,N_3153,N_3341);
nor U3507 (N_3507,N_3393,N_3026);
nor U3508 (N_3508,N_3347,N_3135);
nand U3509 (N_3509,N_3040,N_3451);
xnor U3510 (N_3510,N_3269,N_3215);
nor U3511 (N_3511,N_3199,N_3273);
nand U3512 (N_3512,N_3192,N_3460);
nand U3513 (N_3513,N_3041,N_3021);
nand U3514 (N_3514,N_3487,N_3063);
nand U3515 (N_3515,N_3307,N_3286);
nor U3516 (N_3516,N_3177,N_3406);
nor U3517 (N_3517,N_3488,N_3107);
nand U3518 (N_3518,N_3476,N_3225);
and U3519 (N_3519,N_3113,N_3367);
nand U3520 (N_3520,N_3164,N_3398);
nor U3521 (N_3521,N_3018,N_3285);
xnor U3522 (N_3522,N_3138,N_3163);
nor U3523 (N_3523,N_3370,N_3205);
xnor U3524 (N_3524,N_3196,N_3110);
nand U3525 (N_3525,N_3124,N_3381);
nand U3526 (N_3526,N_3049,N_3275);
or U3527 (N_3527,N_3012,N_3183);
xor U3528 (N_3528,N_3234,N_3233);
xor U3529 (N_3529,N_3038,N_3042);
nor U3530 (N_3530,N_3281,N_3384);
nor U3531 (N_3531,N_3086,N_3459);
nand U3532 (N_3532,N_3206,N_3477);
xor U3533 (N_3533,N_3161,N_3009);
or U3534 (N_3534,N_3463,N_3166);
xnor U3535 (N_3535,N_3264,N_3475);
or U3536 (N_3536,N_3472,N_3249);
nand U3537 (N_3537,N_3061,N_3377);
or U3538 (N_3538,N_3180,N_3080);
or U3539 (N_3539,N_3213,N_3355);
xor U3540 (N_3540,N_3221,N_3154);
nor U3541 (N_3541,N_3141,N_3426);
xnor U3542 (N_3542,N_3142,N_3240);
or U3543 (N_3543,N_3365,N_3146);
xor U3544 (N_3544,N_3470,N_3311);
nand U3545 (N_3545,N_3150,N_3246);
nor U3546 (N_3546,N_3415,N_3447);
xnor U3547 (N_3547,N_3057,N_3013);
and U3548 (N_3548,N_3364,N_3072);
nand U3549 (N_3549,N_3003,N_3202);
xor U3550 (N_3550,N_3125,N_3191);
nor U3551 (N_3551,N_3007,N_3320);
and U3552 (N_3552,N_3111,N_3430);
nand U3553 (N_3553,N_3333,N_3046);
and U3554 (N_3554,N_3066,N_3462);
or U3555 (N_3555,N_3395,N_3235);
nand U3556 (N_3556,N_3027,N_3294);
and U3557 (N_3557,N_3308,N_3145);
xor U3558 (N_3558,N_3485,N_3337);
xor U3559 (N_3559,N_3397,N_3278);
and U3560 (N_3560,N_3318,N_3017);
or U3561 (N_3561,N_3376,N_3179);
nand U3562 (N_3562,N_3372,N_3212);
nor U3563 (N_3563,N_3020,N_3282);
nand U3564 (N_3564,N_3022,N_3468);
and U3565 (N_3565,N_3039,N_3494);
and U3566 (N_3566,N_3139,N_3496);
or U3567 (N_3567,N_3015,N_3416);
and U3568 (N_3568,N_3214,N_3170);
nor U3569 (N_3569,N_3217,N_3375);
nor U3570 (N_3570,N_3326,N_3252);
xnor U3571 (N_3571,N_3152,N_3241);
nand U3572 (N_3572,N_3002,N_3185);
or U3573 (N_3573,N_3108,N_3062);
nor U3574 (N_3574,N_3243,N_3357);
and U3575 (N_3575,N_3469,N_3391);
and U3576 (N_3576,N_3036,N_3174);
and U3577 (N_3577,N_3343,N_3137);
nand U3578 (N_3578,N_3033,N_3228);
xor U3579 (N_3579,N_3330,N_3300);
and U3580 (N_3580,N_3483,N_3369);
xnor U3581 (N_3581,N_3272,N_3328);
nor U3582 (N_3582,N_3335,N_3405);
or U3583 (N_3583,N_3077,N_3000);
xor U3584 (N_3584,N_3133,N_3350);
xnor U3585 (N_3585,N_3474,N_3032);
and U3586 (N_3586,N_3407,N_3043);
nor U3587 (N_3587,N_3271,N_3186);
or U3588 (N_3588,N_3093,N_3418);
xor U3589 (N_3589,N_3280,N_3493);
nor U3590 (N_3590,N_3053,N_3495);
nand U3591 (N_3591,N_3076,N_3218);
or U3592 (N_3592,N_3413,N_3356);
xor U3593 (N_3593,N_3336,N_3081);
nor U3594 (N_3594,N_3155,N_3290);
nand U3595 (N_3595,N_3410,N_3193);
nand U3596 (N_3596,N_3237,N_3298);
nand U3597 (N_3597,N_3445,N_3200);
nor U3598 (N_3598,N_3008,N_3097);
and U3599 (N_3599,N_3480,N_3429);
and U3600 (N_3600,N_3121,N_3226);
nand U3601 (N_3601,N_3473,N_3329);
or U3602 (N_3602,N_3396,N_3197);
or U3603 (N_3603,N_3498,N_3014);
or U3604 (N_3604,N_3359,N_3448);
nor U3605 (N_3605,N_3323,N_3070);
xnor U3606 (N_3606,N_3244,N_3056);
nand U3607 (N_3607,N_3385,N_3047);
xor U3608 (N_3608,N_3283,N_3140);
or U3609 (N_3609,N_3310,N_3064);
or U3610 (N_3610,N_3059,N_3402);
nor U3611 (N_3611,N_3147,N_3342);
nor U3612 (N_3612,N_3016,N_3334);
nor U3613 (N_3613,N_3052,N_3001);
xor U3614 (N_3614,N_3253,N_3119);
xor U3615 (N_3615,N_3490,N_3340);
and U3616 (N_3616,N_3446,N_3112);
or U3617 (N_3617,N_3387,N_3464);
xor U3618 (N_3618,N_3207,N_3096);
and U3619 (N_3619,N_3037,N_3313);
nand U3620 (N_3620,N_3383,N_3123);
xnor U3621 (N_3621,N_3087,N_3044);
nor U3622 (N_3622,N_3288,N_3149);
xnor U3623 (N_3623,N_3079,N_3148);
or U3624 (N_3624,N_3453,N_3344);
nor U3625 (N_3625,N_3263,N_3019);
and U3626 (N_3626,N_3386,N_3169);
and U3627 (N_3627,N_3189,N_3303);
nor U3628 (N_3628,N_3380,N_3222);
xnor U3629 (N_3629,N_3167,N_3031);
or U3630 (N_3630,N_3262,N_3465);
xnor U3631 (N_3631,N_3363,N_3419);
xnor U3632 (N_3632,N_3412,N_3223);
and U3633 (N_3633,N_3486,N_3088);
nor U3634 (N_3634,N_3131,N_3181);
or U3635 (N_3635,N_3443,N_3437);
xnor U3636 (N_3636,N_3100,N_3083);
nor U3637 (N_3637,N_3069,N_3302);
and U3638 (N_3638,N_3030,N_3399);
nand U3639 (N_3639,N_3208,N_3274);
and U3640 (N_3640,N_3297,N_3284);
xor U3641 (N_3641,N_3195,N_3312);
and U3642 (N_3642,N_3051,N_3127);
nor U3643 (N_3643,N_3231,N_3075);
or U3644 (N_3644,N_3368,N_3292);
and U3645 (N_3645,N_3435,N_3394);
or U3646 (N_3646,N_3258,N_3482);
nand U3647 (N_3647,N_3184,N_3442);
xor U3648 (N_3648,N_3073,N_3085);
xnor U3649 (N_3649,N_3165,N_3414);
xnor U3650 (N_3650,N_3242,N_3401);
xnor U3651 (N_3651,N_3287,N_3024);
or U3652 (N_3652,N_3455,N_3102);
and U3653 (N_3653,N_3409,N_3309);
and U3654 (N_3654,N_3373,N_3256);
nand U3655 (N_3655,N_3230,N_3417);
xor U3656 (N_3656,N_3204,N_3104);
and U3657 (N_3657,N_3101,N_3325);
nor U3658 (N_3658,N_3160,N_3245);
nand U3659 (N_3659,N_3029,N_3499);
or U3660 (N_3660,N_3348,N_3130);
and U3661 (N_3661,N_3098,N_3236);
nand U3662 (N_3662,N_3117,N_3366);
and U3663 (N_3663,N_3099,N_3045);
nor U3664 (N_3664,N_3058,N_3425);
xor U3665 (N_3665,N_3456,N_3050);
nand U3666 (N_3666,N_3450,N_3420);
or U3667 (N_3667,N_3411,N_3317);
and U3668 (N_3668,N_3427,N_3362);
or U3669 (N_3669,N_3338,N_3339);
nor U3670 (N_3670,N_3305,N_3182);
xor U3671 (N_3671,N_3109,N_3345);
nor U3672 (N_3672,N_3289,N_3227);
nand U3673 (N_3673,N_3248,N_3265);
nand U3674 (N_3674,N_3006,N_3216);
or U3675 (N_3675,N_3188,N_3010);
nor U3676 (N_3676,N_3094,N_3034);
nor U3677 (N_3677,N_3301,N_3144);
and U3678 (N_3678,N_3322,N_3378);
nand U3679 (N_3679,N_3071,N_3162);
or U3680 (N_3680,N_3404,N_3408);
nand U3681 (N_3681,N_3209,N_3260);
and U3682 (N_3682,N_3319,N_3438);
nand U3683 (N_3683,N_3054,N_3315);
xor U3684 (N_3684,N_3238,N_3481);
nand U3685 (N_3685,N_3440,N_3126);
or U3686 (N_3686,N_3224,N_3279);
xor U3687 (N_3687,N_3324,N_3316);
and U3688 (N_3688,N_3095,N_3115);
or U3689 (N_3689,N_3444,N_3171);
xnor U3690 (N_3690,N_3428,N_3074);
or U3691 (N_3691,N_3390,N_3089);
xnor U3692 (N_3692,N_3361,N_3025);
and U3693 (N_3693,N_3198,N_3210);
nor U3694 (N_3694,N_3422,N_3122);
or U3695 (N_3695,N_3304,N_3277);
or U3696 (N_3696,N_3471,N_3232);
nor U3697 (N_3697,N_3346,N_3035);
and U3698 (N_3698,N_3255,N_3379);
or U3699 (N_3699,N_3492,N_3266);
nand U3700 (N_3700,N_3023,N_3479);
nor U3701 (N_3701,N_3327,N_3299);
nand U3702 (N_3702,N_3353,N_3132);
or U3703 (N_3703,N_3187,N_3331);
nor U3704 (N_3704,N_3067,N_3423);
nor U3705 (N_3705,N_3467,N_3424);
or U3706 (N_3706,N_3203,N_3421);
and U3707 (N_3707,N_3004,N_3461);
nor U3708 (N_3708,N_3114,N_3374);
and U3709 (N_3709,N_3332,N_3005);
nand U3710 (N_3710,N_3201,N_3190);
xnor U3711 (N_3711,N_3259,N_3349);
xor U3712 (N_3712,N_3151,N_3220);
or U3713 (N_3713,N_3143,N_3293);
nor U3714 (N_3714,N_3403,N_3314);
or U3715 (N_3715,N_3178,N_3351);
nor U3716 (N_3716,N_3382,N_3267);
or U3717 (N_3717,N_3484,N_3400);
or U3718 (N_3718,N_3106,N_3432);
xnor U3719 (N_3719,N_3431,N_3173);
xor U3720 (N_3720,N_3276,N_3388);
nand U3721 (N_3721,N_3257,N_3103);
or U3722 (N_3722,N_3295,N_3219);
nor U3723 (N_3723,N_3136,N_3082);
nand U3724 (N_3724,N_3068,N_3352);
nor U3725 (N_3725,N_3158,N_3116);
nor U3726 (N_3726,N_3449,N_3118);
nor U3727 (N_3727,N_3128,N_3229);
and U3728 (N_3728,N_3254,N_3048);
xnor U3729 (N_3729,N_3247,N_3090);
or U3730 (N_3730,N_3296,N_3011);
nand U3731 (N_3731,N_3354,N_3091);
and U3732 (N_3732,N_3458,N_3436);
xnor U3733 (N_3733,N_3454,N_3157);
xor U3734 (N_3734,N_3358,N_3389);
and U3735 (N_3735,N_3457,N_3360);
nand U3736 (N_3736,N_3156,N_3092);
nand U3737 (N_3737,N_3176,N_3433);
and U3738 (N_3738,N_3371,N_3134);
and U3739 (N_3739,N_3194,N_3120);
xor U3740 (N_3740,N_3175,N_3392);
or U3741 (N_3741,N_3055,N_3441);
nand U3742 (N_3742,N_3489,N_3239);
nand U3743 (N_3743,N_3211,N_3291);
and U3744 (N_3744,N_3466,N_3452);
and U3745 (N_3745,N_3168,N_3306);
or U3746 (N_3746,N_3261,N_3105);
or U3747 (N_3747,N_3078,N_3491);
xor U3748 (N_3748,N_3478,N_3065);
nand U3749 (N_3749,N_3270,N_3497);
xnor U3750 (N_3750,N_3424,N_3384);
and U3751 (N_3751,N_3275,N_3349);
and U3752 (N_3752,N_3184,N_3169);
nand U3753 (N_3753,N_3048,N_3044);
xor U3754 (N_3754,N_3110,N_3031);
and U3755 (N_3755,N_3017,N_3397);
and U3756 (N_3756,N_3344,N_3368);
nor U3757 (N_3757,N_3248,N_3383);
xnor U3758 (N_3758,N_3287,N_3104);
nand U3759 (N_3759,N_3104,N_3193);
and U3760 (N_3760,N_3178,N_3068);
nor U3761 (N_3761,N_3082,N_3200);
or U3762 (N_3762,N_3015,N_3214);
nand U3763 (N_3763,N_3049,N_3126);
and U3764 (N_3764,N_3298,N_3277);
nor U3765 (N_3765,N_3068,N_3313);
nand U3766 (N_3766,N_3192,N_3247);
nand U3767 (N_3767,N_3000,N_3317);
and U3768 (N_3768,N_3474,N_3361);
nor U3769 (N_3769,N_3329,N_3257);
nor U3770 (N_3770,N_3329,N_3350);
xnor U3771 (N_3771,N_3128,N_3119);
nor U3772 (N_3772,N_3423,N_3418);
or U3773 (N_3773,N_3260,N_3173);
nand U3774 (N_3774,N_3251,N_3465);
and U3775 (N_3775,N_3195,N_3277);
and U3776 (N_3776,N_3398,N_3262);
and U3777 (N_3777,N_3495,N_3047);
and U3778 (N_3778,N_3083,N_3438);
nand U3779 (N_3779,N_3124,N_3183);
xor U3780 (N_3780,N_3131,N_3411);
nand U3781 (N_3781,N_3414,N_3297);
nor U3782 (N_3782,N_3102,N_3096);
and U3783 (N_3783,N_3471,N_3264);
or U3784 (N_3784,N_3374,N_3461);
nand U3785 (N_3785,N_3339,N_3191);
nand U3786 (N_3786,N_3057,N_3144);
nor U3787 (N_3787,N_3302,N_3257);
or U3788 (N_3788,N_3142,N_3104);
nand U3789 (N_3789,N_3227,N_3492);
and U3790 (N_3790,N_3021,N_3219);
nand U3791 (N_3791,N_3245,N_3101);
nor U3792 (N_3792,N_3376,N_3242);
xor U3793 (N_3793,N_3344,N_3172);
nor U3794 (N_3794,N_3316,N_3377);
xor U3795 (N_3795,N_3069,N_3375);
nor U3796 (N_3796,N_3279,N_3252);
or U3797 (N_3797,N_3301,N_3323);
xnor U3798 (N_3798,N_3203,N_3036);
nand U3799 (N_3799,N_3262,N_3194);
and U3800 (N_3800,N_3478,N_3111);
nand U3801 (N_3801,N_3327,N_3489);
nor U3802 (N_3802,N_3203,N_3224);
xnor U3803 (N_3803,N_3276,N_3199);
and U3804 (N_3804,N_3006,N_3058);
or U3805 (N_3805,N_3122,N_3097);
and U3806 (N_3806,N_3071,N_3130);
or U3807 (N_3807,N_3046,N_3177);
nand U3808 (N_3808,N_3428,N_3070);
and U3809 (N_3809,N_3332,N_3358);
nor U3810 (N_3810,N_3352,N_3045);
or U3811 (N_3811,N_3275,N_3168);
nor U3812 (N_3812,N_3133,N_3171);
nor U3813 (N_3813,N_3104,N_3497);
xor U3814 (N_3814,N_3413,N_3138);
and U3815 (N_3815,N_3353,N_3296);
or U3816 (N_3816,N_3279,N_3093);
xor U3817 (N_3817,N_3455,N_3365);
nor U3818 (N_3818,N_3011,N_3472);
nor U3819 (N_3819,N_3132,N_3346);
nand U3820 (N_3820,N_3102,N_3048);
or U3821 (N_3821,N_3331,N_3385);
xor U3822 (N_3822,N_3376,N_3319);
or U3823 (N_3823,N_3470,N_3394);
and U3824 (N_3824,N_3259,N_3330);
or U3825 (N_3825,N_3152,N_3064);
nand U3826 (N_3826,N_3299,N_3247);
or U3827 (N_3827,N_3477,N_3414);
and U3828 (N_3828,N_3365,N_3159);
and U3829 (N_3829,N_3071,N_3096);
nor U3830 (N_3830,N_3089,N_3261);
or U3831 (N_3831,N_3080,N_3078);
or U3832 (N_3832,N_3307,N_3489);
or U3833 (N_3833,N_3372,N_3044);
xnor U3834 (N_3834,N_3482,N_3239);
or U3835 (N_3835,N_3344,N_3373);
or U3836 (N_3836,N_3163,N_3370);
nor U3837 (N_3837,N_3055,N_3179);
or U3838 (N_3838,N_3400,N_3211);
xnor U3839 (N_3839,N_3261,N_3281);
xnor U3840 (N_3840,N_3199,N_3390);
and U3841 (N_3841,N_3395,N_3348);
xor U3842 (N_3842,N_3213,N_3278);
xor U3843 (N_3843,N_3461,N_3188);
or U3844 (N_3844,N_3420,N_3242);
nor U3845 (N_3845,N_3277,N_3463);
nor U3846 (N_3846,N_3156,N_3400);
and U3847 (N_3847,N_3189,N_3270);
nor U3848 (N_3848,N_3114,N_3255);
xnor U3849 (N_3849,N_3314,N_3145);
and U3850 (N_3850,N_3388,N_3499);
xnor U3851 (N_3851,N_3338,N_3022);
nand U3852 (N_3852,N_3488,N_3008);
and U3853 (N_3853,N_3386,N_3396);
xor U3854 (N_3854,N_3018,N_3310);
and U3855 (N_3855,N_3415,N_3020);
or U3856 (N_3856,N_3041,N_3166);
nor U3857 (N_3857,N_3001,N_3470);
and U3858 (N_3858,N_3236,N_3312);
nor U3859 (N_3859,N_3386,N_3175);
or U3860 (N_3860,N_3389,N_3119);
nor U3861 (N_3861,N_3396,N_3211);
or U3862 (N_3862,N_3220,N_3066);
nor U3863 (N_3863,N_3278,N_3027);
or U3864 (N_3864,N_3026,N_3236);
xnor U3865 (N_3865,N_3066,N_3309);
and U3866 (N_3866,N_3206,N_3324);
nand U3867 (N_3867,N_3478,N_3492);
or U3868 (N_3868,N_3076,N_3469);
nand U3869 (N_3869,N_3487,N_3169);
nor U3870 (N_3870,N_3201,N_3141);
or U3871 (N_3871,N_3085,N_3335);
or U3872 (N_3872,N_3021,N_3080);
and U3873 (N_3873,N_3168,N_3043);
and U3874 (N_3874,N_3471,N_3065);
xnor U3875 (N_3875,N_3306,N_3461);
nor U3876 (N_3876,N_3031,N_3392);
nand U3877 (N_3877,N_3258,N_3397);
or U3878 (N_3878,N_3106,N_3151);
or U3879 (N_3879,N_3103,N_3453);
or U3880 (N_3880,N_3486,N_3352);
and U3881 (N_3881,N_3166,N_3141);
or U3882 (N_3882,N_3060,N_3220);
xor U3883 (N_3883,N_3336,N_3361);
nor U3884 (N_3884,N_3073,N_3063);
nand U3885 (N_3885,N_3427,N_3469);
nor U3886 (N_3886,N_3104,N_3448);
xnor U3887 (N_3887,N_3245,N_3038);
nor U3888 (N_3888,N_3307,N_3014);
and U3889 (N_3889,N_3390,N_3421);
or U3890 (N_3890,N_3100,N_3184);
nand U3891 (N_3891,N_3194,N_3431);
and U3892 (N_3892,N_3455,N_3016);
xnor U3893 (N_3893,N_3264,N_3397);
xor U3894 (N_3894,N_3242,N_3065);
and U3895 (N_3895,N_3496,N_3259);
nor U3896 (N_3896,N_3444,N_3273);
and U3897 (N_3897,N_3111,N_3141);
nor U3898 (N_3898,N_3255,N_3374);
xor U3899 (N_3899,N_3422,N_3264);
or U3900 (N_3900,N_3312,N_3059);
nor U3901 (N_3901,N_3001,N_3035);
xor U3902 (N_3902,N_3224,N_3317);
and U3903 (N_3903,N_3210,N_3168);
or U3904 (N_3904,N_3349,N_3428);
and U3905 (N_3905,N_3350,N_3164);
or U3906 (N_3906,N_3265,N_3066);
or U3907 (N_3907,N_3414,N_3401);
and U3908 (N_3908,N_3367,N_3028);
nand U3909 (N_3909,N_3025,N_3098);
or U3910 (N_3910,N_3080,N_3084);
nor U3911 (N_3911,N_3060,N_3032);
nor U3912 (N_3912,N_3193,N_3497);
and U3913 (N_3913,N_3369,N_3253);
nand U3914 (N_3914,N_3179,N_3142);
and U3915 (N_3915,N_3103,N_3237);
or U3916 (N_3916,N_3299,N_3295);
and U3917 (N_3917,N_3312,N_3353);
and U3918 (N_3918,N_3025,N_3075);
and U3919 (N_3919,N_3025,N_3170);
nand U3920 (N_3920,N_3254,N_3266);
xnor U3921 (N_3921,N_3098,N_3053);
or U3922 (N_3922,N_3403,N_3193);
nor U3923 (N_3923,N_3408,N_3245);
nor U3924 (N_3924,N_3055,N_3336);
nor U3925 (N_3925,N_3299,N_3171);
and U3926 (N_3926,N_3239,N_3301);
nor U3927 (N_3927,N_3428,N_3136);
nor U3928 (N_3928,N_3328,N_3240);
xnor U3929 (N_3929,N_3100,N_3186);
xor U3930 (N_3930,N_3328,N_3046);
and U3931 (N_3931,N_3341,N_3239);
nor U3932 (N_3932,N_3333,N_3077);
xor U3933 (N_3933,N_3299,N_3309);
xnor U3934 (N_3934,N_3330,N_3382);
or U3935 (N_3935,N_3055,N_3414);
or U3936 (N_3936,N_3481,N_3085);
or U3937 (N_3937,N_3356,N_3468);
nand U3938 (N_3938,N_3318,N_3038);
and U3939 (N_3939,N_3403,N_3166);
xnor U3940 (N_3940,N_3035,N_3369);
or U3941 (N_3941,N_3340,N_3177);
xnor U3942 (N_3942,N_3431,N_3000);
nor U3943 (N_3943,N_3427,N_3088);
and U3944 (N_3944,N_3424,N_3062);
and U3945 (N_3945,N_3335,N_3071);
nor U3946 (N_3946,N_3414,N_3240);
and U3947 (N_3947,N_3460,N_3223);
or U3948 (N_3948,N_3095,N_3449);
and U3949 (N_3949,N_3470,N_3207);
nand U3950 (N_3950,N_3205,N_3418);
or U3951 (N_3951,N_3004,N_3281);
or U3952 (N_3952,N_3323,N_3124);
and U3953 (N_3953,N_3420,N_3434);
and U3954 (N_3954,N_3499,N_3116);
xnor U3955 (N_3955,N_3170,N_3222);
nor U3956 (N_3956,N_3097,N_3296);
and U3957 (N_3957,N_3420,N_3326);
and U3958 (N_3958,N_3236,N_3126);
nand U3959 (N_3959,N_3161,N_3287);
and U3960 (N_3960,N_3206,N_3093);
nor U3961 (N_3961,N_3342,N_3052);
or U3962 (N_3962,N_3116,N_3459);
and U3963 (N_3963,N_3022,N_3137);
and U3964 (N_3964,N_3107,N_3054);
nand U3965 (N_3965,N_3451,N_3499);
nor U3966 (N_3966,N_3301,N_3210);
and U3967 (N_3967,N_3323,N_3108);
nand U3968 (N_3968,N_3062,N_3475);
nand U3969 (N_3969,N_3438,N_3311);
xnor U3970 (N_3970,N_3493,N_3149);
nor U3971 (N_3971,N_3231,N_3207);
and U3972 (N_3972,N_3125,N_3130);
nand U3973 (N_3973,N_3327,N_3125);
or U3974 (N_3974,N_3034,N_3475);
or U3975 (N_3975,N_3447,N_3328);
xor U3976 (N_3976,N_3360,N_3016);
and U3977 (N_3977,N_3491,N_3318);
and U3978 (N_3978,N_3184,N_3123);
and U3979 (N_3979,N_3100,N_3394);
xor U3980 (N_3980,N_3133,N_3064);
and U3981 (N_3981,N_3418,N_3334);
nand U3982 (N_3982,N_3158,N_3167);
and U3983 (N_3983,N_3015,N_3000);
and U3984 (N_3984,N_3436,N_3092);
or U3985 (N_3985,N_3040,N_3104);
nand U3986 (N_3986,N_3200,N_3310);
xor U3987 (N_3987,N_3214,N_3353);
nand U3988 (N_3988,N_3390,N_3118);
xor U3989 (N_3989,N_3410,N_3286);
or U3990 (N_3990,N_3054,N_3142);
or U3991 (N_3991,N_3367,N_3075);
nand U3992 (N_3992,N_3031,N_3083);
xor U3993 (N_3993,N_3105,N_3054);
or U3994 (N_3994,N_3299,N_3217);
and U3995 (N_3995,N_3003,N_3021);
nand U3996 (N_3996,N_3247,N_3040);
or U3997 (N_3997,N_3347,N_3066);
nand U3998 (N_3998,N_3026,N_3363);
or U3999 (N_3999,N_3109,N_3103);
or U4000 (N_4000,N_3660,N_3991);
xnor U4001 (N_4001,N_3894,N_3607);
xnor U4002 (N_4002,N_3711,N_3682);
or U4003 (N_4003,N_3520,N_3988);
xor U4004 (N_4004,N_3788,N_3935);
and U4005 (N_4005,N_3547,N_3752);
nand U4006 (N_4006,N_3539,N_3951);
nand U4007 (N_4007,N_3865,N_3965);
nand U4008 (N_4008,N_3784,N_3576);
nand U4009 (N_4009,N_3958,N_3675);
nor U4010 (N_4010,N_3756,N_3623);
xor U4011 (N_4011,N_3727,N_3587);
or U4012 (N_4012,N_3797,N_3507);
xnor U4013 (N_4013,N_3963,N_3923);
and U4014 (N_4014,N_3810,N_3613);
nand U4015 (N_4015,N_3673,N_3892);
and U4016 (N_4016,N_3853,N_3553);
and U4017 (N_4017,N_3896,N_3580);
xor U4018 (N_4018,N_3969,N_3645);
or U4019 (N_4019,N_3719,N_3976);
or U4020 (N_4020,N_3781,N_3642);
or U4021 (N_4021,N_3689,N_3891);
nand U4022 (N_4022,N_3629,N_3852);
nor U4023 (N_4023,N_3888,N_3605);
or U4024 (N_4024,N_3811,N_3981);
xor U4025 (N_4025,N_3943,N_3582);
xor U4026 (N_4026,N_3674,N_3595);
or U4027 (N_4027,N_3728,N_3750);
and U4028 (N_4028,N_3989,N_3790);
nor U4029 (N_4029,N_3535,N_3816);
nand U4030 (N_4030,N_3872,N_3566);
or U4031 (N_4031,N_3834,N_3759);
xnor U4032 (N_4032,N_3622,N_3786);
or U4033 (N_4033,N_3597,N_3821);
xnor U4034 (N_4034,N_3505,N_3835);
nand U4035 (N_4035,N_3650,N_3792);
and U4036 (N_4036,N_3628,N_3959);
xor U4037 (N_4037,N_3747,N_3990);
nor U4038 (N_4038,N_3742,N_3905);
and U4039 (N_4039,N_3569,N_3700);
nor U4040 (N_4040,N_3545,N_3731);
nand U4041 (N_4041,N_3726,N_3699);
nor U4042 (N_4042,N_3718,N_3616);
xnor U4043 (N_4043,N_3909,N_3528);
xnor U4044 (N_4044,N_3533,N_3670);
or U4045 (N_4045,N_3679,N_3836);
and U4046 (N_4046,N_3926,N_3575);
and U4047 (N_4047,N_3739,N_3802);
nand U4048 (N_4048,N_3634,N_3820);
xor U4049 (N_4049,N_3666,N_3911);
nor U4050 (N_4050,N_3920,N_3663);
nand U4051 (N_4051,N_3655,N_3626);
and U4052 (N_4052,N_3778,N_3721);
or U4053 (N_4053,N_3832,N_3997);
nor U4054 (N_4054,N_3515,N_3644);
and U4055 (N_4055,N_3695,N_3823);
xnor U4056 (N_4056,N_3783,N_3680);
nor U4057 (N_4057,N_3858,N_3662);
nand U4058 (N_4058,N_3782,N_3600);
nand U4059 (N_4059,N_3702,N_3937);
nand U4060 (N_4060,N_3803,N_3620);
nor U4061 (N_4061,N_3516,N_3860);
or U4062 (N_4062,N_3966,N_3972);
nor U4063 (N_4063,N_3636,N_3824);
nor U4064 (N_4064,N_3771,N_3912);
or U4065 (N_4065,N_3665,N_3766);
nand U4066 (N_4066,N_3598,N_3574);
and U4067 (N_4067,N_3948,N_3931);
nor U4068 (N_4068,N_3971,N_3900);
or U4069 (N_4069,N_3698,N_3866);
and U4070 (N_4070,N_3714,N_3720);
nand U4071 (N_4071,N_3585,N_3627);
or U4072 (N_4072,N_3930,N_3913);
or U4073 (N_4073,N_3640,N_3678);
xor U4074 (N_4074,N_3631,N_3667);
nor U4075 (N_4075,N_3939,N_3744);
and U4076 (N_4076,N_3651,N_3929);
and U4077 (N_4077,N_3557,N_3643);
xor U4078 (N_4078,N_3796,N_3915);
nand U4079 (N_4079,N_3985,N_3813);
xnor U4080 (N_4080,N_3579,N_3761);
nor U4081 (N_4081,N_3710,N_3549);
and U4082 (N_4082,N_3639,N_3565);
nor U4083 (N_4083,N_3854,N_3876);
and U4084 (N_4084,N_3996,N_3558);
xor U4085 (N_4085,N_3837,N_3632);
nor U4086 (N_4086,N_3513,N_3998);
or U4087 (N_4087,N_3849,N_3691);
and U4088 (N_4088,N_3671,N_3737);
nor U4089 (N_4089,N_3509,N_3583);
nand U4090 (N_4090,N_3812,N_3502);
and U4091 (N_4091,N_3897,N_3561);
xor U4092 (N_4092,N_3530,N_3946);
nand U4093 (N_4093,N_3864,N_3952);
or U4094 (N_4094,N_3540,N_3577);
and U4095 (N_4095,N_3992,N_3503);
or U4096 (N_4096,N_3850,N_3704);
and U4097 (N_4097,N_3567,N_3536);
nor U4098 (N_4098,N_3975,N_3770);
xor U4099 (N_4099,N_3571,N_3922);
nand U4100 (N_4100,N_3725,N_3610);
xnor U4101 (N_4101,N_3621,N_3588);
nor U4102 (N_4102,N_3983,N_3517);
and U4103 (N_4103,N_3659,N_3995);
xnor U4104 (N_4104,N_3551,N_3870);
and U4105 (N_4105,N_3510,N_3572);
or U4106 (N_4106,N_3791,N_3984);
xor U4107 (N_4107,N_3809,N_3732);
nand U4108 (N_4108,N_3570,N_3871);
nor U4109 (N_4109,N_3706,N_3690);
nand U4110 (N_4110,N_3833,N_3962);
nand U4111 (N_4111,N_3844,N_3521);
or U4112 (N_4112,N_3548,N_3822);
xor U4113 (N_4113,N_3648,N_3859);
xor U4114 (N_4114,N_3688,N_3668);
nand U4115 (N_4115,N_3800,N_3608);
or U4116 (N_4116,N_3942,N_3534);
and U4117 (N_4117,N_3907,N_3889);
xor U4118 (N_4118,N_3735,N_3947);
nor U4119 (N_4119,N_3960,N_3685);
or U4120 (N_4120,N_3635,N_3977);
nor U4121 (N_4121,N_3776,N_3514);
nor U4122 (N_4122,N_3869,N_3618);
xor U4123 (N_4123,N_3581,N_3980);
xor U4124 (N_4124,N_3885,N_3707);
nand U4125 (N_4125,N_3795,N_3921);
or U4126 (N_4126,N_3729,N_3881);
xor U4127 (N_4127,N_3902,N_3649);
nand U4128 (N_4128,N_3532,N_3949);
nand U4129 (N_4129,N_3838,N_3654);
nand U4130 (N_4130,N_3760,N_3694);
nand U4131 (N_4131,N_3775,N_3772);
and U4132 (N_4132,N_3954,N_3664);
xnor U4133 (N_4133,N_3882,N_3681);
xnor U4134 (N_4134,N_3774,N_3831);
or U4135 (N_4135,N_3573,N_3855);
and U4136 (N_4136,N_3601,N_3712);
and U4137 (N_4137,N_3841,N_3780);
and U4138 (N_4138,N_3856,N_3550);
nor U4139 (N_4139,N_3504,N_3918);
nor U4140 (N_4140,N_3611,N_3697);
xor U4141 (N_4141,N_3693,N_3619);
xnor U4142 (N_4142,N_3722,N_3878);
nor U4143 (N_4143,N_3819,N_3519);
nor U4144 (N_4144,N_3687,N_3677);
xnor U4145 (N_4145,N_3908,N_3542);
or U4146 (N_4146,N_3589,N_3877);
or U4147 (N_4147,N_3967,N_3827);
or U4148 (N_4148,N_3749,N_3842);
and U4149 (N_4149,N_3511,N_3746);
xor U4150 (N_4150,N_3932,N_3646);
or U4151 (N_4151,N_3925,N_3979);
and U4152 (N_4152,N_3506,N_3596);
xor U4153 (N_4153,N_3846,N_3686);
nand U4154 (N_4154,N_3578,N_3763);
xor U4155 (N_4155,N_3652,N_3789);
xor U4156 (N_4156,N_3705,N_3713);
nand U4157 (N_4157,N_3936,N_3653);
and U4158 (N_4158,N_3993,N_3906);
nand U4159 (N_4159,N_3564,N_3556);
nand U4160 (N_4160,N_3968,N_3753);
and U4161 (N_4161,N_3825,N_3875);
xor U4162 (N_4162,N_3748,N_3741);
and U4163 (N_4163,N_3716,N_3754);
and U4164 (N_4164,N_3609,N_3893);
xnor U4165 (N_4165,N_3987,N_3798);
or U4166 (N_4166,N_3543,N_3683);
xnor U4167 (N_4167,N_3630,N_3839);
nand U4168 (N_4168,N_3916,N_3730);
nand U4169 (N_4169,N_3669,N_3898);
or U4170 (N_4170,N_3944,N_3563);
xnor U4171 (N_4171,N_3594,N_3590);
or U4172 (N_4172,N_3895,N_3938);
or U4173 (N_4173,N_3562,N_3523);
xor U4174 (N_4174,N_3779,N_3879);
or U4175 (N_4175,N_3733,N_3787);
or U4176 (N_4176,N_3901,N_3501);
or U4177 (N_4177,N_3522,N_3956);
and U4178 (N_4178,N_3941,N_3890);
nor U4179 (N_4179,N_3538,N_3606);
nor U4180 (N_4180,N_3518,N_3999);
nor U4181 (N_4181,N_3874,N_3961);
or U4182 (N_4182,N_3757,N_3830);
nand U4183 (N_4183,N_3927,N_3934);
or U4184 (N_4184,N_3970,N_3637);
xnor U4185 (N_4185,N_3676,N_3724);
and U4186 (N_4186,N_3641,N_3814);
and U4187 (N_4187,N_3696,N_3828);
xor U4188 (N_4188,N_3692,N_3751);
and U4189 (N_4189,N_3806,N_3848);
and U4190 (N_4190,N_3883,N_3886);
xor U4191 (N_4191,N_3843,N_3857);
nor U4192 (N_4192,N_3829,N_3978);
xor U4193 (N_4193,N_3529,N_3591);
xnor U4194 (N_4194,N_3773,N_3762);
or U4195 (N_4195,N_3512,N_3526);
and U4196 (N_4196,N_3604,N_3982);
and U4197 (N_4197,N_3955,N_3862);
or U4198 (N_4198,N_3840,N_3986);
nand U4199 (N_4199,N_3868,N_3793);
nor U4200 (N_4200,N_3861,N_3624);
nor U4201 (N_4201,N_3745,N_3658);
and U4202 (N_4202,N_3568,N_3544);
xor U4203 (N_4203,N_3817,N_3586);
and U4204 (N_4204,N_3701,N_3863);
nor U4205 (N_4205,N_3994,N_3801);
nor U4206 (N_4206,N_3917,N_3950);
xor U4207 (N_4207,N_3924,N_3612);
xor U4208 (N_4208,N_3656,N_3884);
and U4209 (N_4209,N_3738,N_3537);
nor U4210 (N_4210,N_3717,N_3851);
xor U4211 (N_4211,N_3880,N_3715);
or U4212 (N_4212,N_3555,N_3815);
nand U4213 (N_4213,N_3867,N_3887);
nor U4214 (N_4214,N_3541,N_3899);
nand U4215 (N_4215,N_3767,N_3661);
or U4216 (N_4216,N_3953,N_3599);
nand U4217 (N_4217,N_3531,N_3777);
or U4218 (N_4218,N_3684,N_3914);
and U4219 (N_4219,N_3617,N_3638);
xnor U4220 (N_4220,N_3808,N_3740);
xor U4221 (N_4221,N_3603,N_3964);
or U4222 (N_4222,N_3552,N_3945);
xor U4223 (N_4223,N_3957,N_3758);
nand U4224 (N_4224,N_3615,N_3799);
xnor U4225 (N_4225,N_3709,N_3764);
or U4226 (N_4226,N_3818,N_3768);
and U4227 (N_4227,N_3584,N_3633);
and U4228 (N_4228,N_3602,N_3973);
nand U4229 (N_4229,N_3559,N_3625);
nor U4230 (N_4230,N_3593,N_3904);
xor U4231 (N_4231,N_3765,N_3500);
or U4232 (N_4232,N_3847,N_3873);
nor U4233 (N_4233,N_3614,N_3919);
nor U4234 (N_4234,N_3524,N_3647);
and U4235 (N_4235,N_3527,N_3794);
and U4236 (N_4236,N_3769,N_3974);
nor U4237 (N_4237,N_3554,N_3736);
nor U4238 (N_4238,N_3933,N_3940);
and U4239 (N_4239,N_3560,N_3785);
xnor U4240 (N_4240,N_3734,N_3508);
nor U4241 (N_4241,N_3928,N_3546);
xor U4242 (N_4242,N_3845,N_3657);
nor U4243 (N_4243,N_3525,N_3723);
or U4244 (N_4244,N_3592,N_3708);
xnor U4245 (N_4245,N_3672,N_3910);
xor U4246 (N_4246,N_3755,N_3805);
xor U4247 (N_4247,N_3743,N_3826);
and U4248 (N_4248,N_3804,N_3703);
and U4249 (N_4249,N_3903,N_3807);
and U4250 (N_4250,N_3899,N_3925);
or U4251 (N_4251,N_3923,N_3677);
xor U4252 (N_4252,N_3755,N_3659);
nand U4253 (N_4253,N_3613,N_3790);
xor U4254 (N_4254,N_3872,N_3924);
xor U4255 (N_4255,N_3704,N_3899);
nor U4256 (N_4256,N_3709,N_3651);
and U4257 (N_4257,N_3800,N_3665);
or U4258 (N_4258,N_3887,N_3621);
xor U4259 (N_4259,N_3913,N_3854);
and U4260 (N_4260,N_3848,N_3605);
or U4261 (N_4261,N_3870,N_3843);
nor U4262 (N_4262,N_3539,N_3538);
xnor U4263 (N_4263,N_3868,N_3620);
xnor U4264 (N_4264,N_3957,N_3608);
xnor U4265 (N_4265,N_3735,N_3556);
xor U4266 (N_4266,N_3929,N_3903);
or U4267 (N_4267,N_3784,N_3564);
nor U4268 (N_4268,N_3577,N_3942);
nand U4269 (N_4269,N_3580,N_3638);
or U4270 (N_4270,N_3628,N_3540);
xor U4271 (N_4271,N_3726,N_3600);
nor U4272 (N_4272,N_3998,N_3842);
and U4273 (N_4273,N_3578,N_3633);
or U4274 (N_4274,N_3791,N_3880);
nand U4275 (N_4275,N_3856,N_3905);
nor U4276 (N_4276,N_3677,N_3544);
or U4277 (N_4277,N_3575,N_3510);
or U4278 (N_4278,N_3751,N_3910);
xor U4279 (N_4279,N_3759,N_3678);
xor U4280 (N_4280,N_3809,N_3701);
and U4281 (N_4281,N_3860,N_3638);
or U4282 (N_4282,N_3517,N_3749);
and U4283 (N_4283,N_3633,N_3690);
nand U4284 (N_4284,N_3939,N_3891);
and U4285 (N_4285,N_3868,N_3654);
or U4286 (N_4286,N_3690,N_3694);
and U4287 (N_4287,N_3571,N_3856);
xnor U4288 (N_4288,N_3949,N_3845);
or U4289 (N_4289,N_3692,N_3918);
or U4290 (N_4290,N_3960,N_3539);
nor U4291 (N_4291,N_3533,N_3904);
nand U4292 (N_4292,N_3649,N_3799);
nor U4293 (N_4293,N_3957,N_3659);
and U4294 (N_4294,N_3542,N_3663);
nor U4295 (N_4295,N_3902,N_3653);
and U4296 (N_4296,N_3566,N_3989);
xnor U4297 (N_4297,N_3589,N_3587);
xor U4298 (N_4298,N_3687,N_3507);
or U4299 (N_4299,N_3914,N_3973);
and U4300 (N_4300,N_3585,N_3511);
and U4301 (N_4301,N_3600,N_3516);
xnor U4302 (N_4302,N_3985,N_3983);
or U4303 (N_4303,N_3796,N_3638);
or U4304 (N_4304,N_3914,N_3890);
and U4305 (N_4305,N_3773,N_3620);
nand U4306 (N_4306,N_3634,N_3816);
nand U4307 (N_4307,N_3770,N_3740);
xnor U4308 (N_4308,N_3879,N_3513);
nor U4309 (N_4309,N_3669,N_3810);
nand U4310 (N_4310,N_3960,N_3605);
nand U4311 (N_4311,N_3788,N_3623);
xnor U4312 (N_4312,N_3996,N_3549);
and U4313 (N_4313,N_3565,N_3540);
xnor U4314 (N_4314,N_3973,N_3967);
nand U4315 (N_4315,N_3787,N_3528);
and U4316 (N_4316,N_3551,N_3806);
nand U4317 (N_4317,N_3910,N_3969);
nand U4318 (N_4318,N_3606,N_3515);
and U4319 (N_4319,N_3739,N_3648);
nor U4320 (N_4320,N_3619,N_3743);
nand U4321 (N_4321,N_3560,N_3783);
and U4322 (N_4322,N_3743,N_3591);
nand U4323 (N_4323,N_3878,N_3731);
and U4324 (N_4324,N_3951,N_3866);
and U4325 (N_4325,N_3582,N_3847);
nand U4326 (N_4326,N_3890,N_3788);
and U4327 (N_4327,N_3756,N_3629);
nor U4328 (N_4328,N_3923,N_3723);
and U4329 (N_4329,N_3953,N_3635);
nor U4330 (N_4330,N_3678,N_3942);
nor U4331 (N_4331,N_3656,N_3890);
nor U4332 (N_4332,N_3771,N_3789);
xnor U4333 (N_4333,N_3806,N_3849);
and U4334 (N_4334,N_3564,N_3618);
nor U4335 (N_4335,N_3698,N_3730);
nor U4336 (N_4336,N_3964,N_3884);
nand U4337 (N_4337,N_3551,N_3922);
xor U4338 (N_4338,N_3950,N_3518);
nand U4339 (N_4339,N_3651,N_3941);
xnor U4340 (N_4340,N_3896,N_3547);
xnor U4341 (N_4341,N_3991,N_3958);
or U4342 (N_4342,N_3932,N_3555);
nor U4343 (N_4343,N_3628,N_3726);
nand U4344 (N_4344,N_3869,N_3851);
nor U4345 (N_4345,N_3517,N_3979);
or U4346 (N_4346,N_3833,N_3890);
and U4347 (N_4347,N_3570,N_3656);
nor U4348 (N_4348,N_3625,N_3875);
nor U4349 (N_4349,N_3758,N_3910);
nor U4350 (N_4350,N_3905,N_3584);
nand U4351 (N_4351,N_3693,N_3523);
xnor U4352 (N_4352,N_3836,N_3896);
and U4353 (N_4353,N_3569,N_3548);
or U4354 (N_4354,N_3818,N_3869);
and U4355 (N_4355,N_3525,N_3731);
xnor U4356 (N_4356,N_3714,N_3756);
xor U4357 (N_4357,N_3807,N_3668);
and U4358 (N_4358,N_3800,N_3715);
nand U4359 (N_4359,N_3969,N_3728);
nand U4360 (N_4360,N_3888,N_3953);
nand U4361 (N_4361,N_3785,N_3577);
nor U4362 (N_4362,N_3948,N_3899);
and U4363 (N_4363,N_3851,N_3544);
xnor U4364 (N_4364,N_3975,N_3919);
nand U4365 (N_4365,N_3946,N_3511);
and U4366 (N_4366,N_3617,N_3656);
xnor U4367 (N_4367,N_3768,N_3723);
or U4368 (N_4368,N_3667,N_3791);
and U4369 (N_4369,N_3648,N_3557);
nand U4370 (N_4370,N_3629,N_3624);
or U4371 (N_4371,N_3510,N_3869);
xnor U4372 (N_4372,N_3905,N_3665);
nand U4373 (N_4373,N_3951,N_3774);
xnor U4374 (N_4374,N_3587,N_3707);
xnor U4375 (N_4375,N_3664,N_3617);
nand U4376 (N_4376,N_3688,N_3719);
xnor U4377 (N_4377,N_3788,N_3664);
or U4378 (N_4378,N_3635,N_3514);
nor U4379 (N_4379,N_3962,N_3507);
and U4380 (N_4380,N_3552,N_3596);
or U4381 (N_4381,N_3630,N_3840);
nand U4382 (N_4382,N_3671,N_3616);
nand U4383 (N_4383,N_3706,N_3589);
or U4384 (N_4384,N_3535,N_3957);
nand U4385 (N_4385,N_3983,N_3818);
nand U4386 (N_4386,N_3801,N_3763);
and U4387 (N_4387,N_3724,N_3971);
or U4388 (N_4388,N_3879,N_3516);
nand U4389 (N_4389,N_3592,N_3759);
nor U4390 (N_4390,N_3770,N_3982);
or U4391 (N_4391,N_3972,N_3529);
or U4392 (N_4392,N_3807,N_3535);
nor U4393 (N_4393,N_3731,N_3934);
and U4394 (N_4394,N_3581,N_3560);
nor U4395 (N_4395,N_3651,N_3913);
and U4396 (N_4396,N_3518,N_3709);
nor U4397 (N_4397,N_3511,N_3718);
nor U4398 (N_4398,N_3970,N_3993);
nand U4399 (N_4399,N_3564,N_3630);
nand U4400 (N_4400,N_3559,N_3848);
nand U4401 (N_4401,N_3535,N_3908);
and U4402 (N_4402,N_3729,N_3774);
or U4403 (N_4403,N_3731,N_3724);
or U4404 (N_4404,N_3590,N_3683);
nand U4405 (N_4405,N_3995,N_3955);
or U4406 (N_4406,N_3886,N_3900);
nor U4407 (N_4407,N_3939,N_3906);
nand U4408 (N_4408,N_3626,N_3674);
and U4409 (N_4409,N_3718,N_3777);
nor U4410 (N_4410,N_3565,N_3762);
or U4411 (N_4411,N_3599,N_3703);
nand U4412 (N_4412,N_3963,N_3737);
nor U4413 (N_4413,N_3708,N_3516);
and U4414 (N_4414,N_3577,N_3853);
or U4415 (N_4415,N_3823,N_3824);
nor U4416 (N_4416,N_3907,N_3617);
and U4417 (N_4417,N_3639,N_3728);
and U4418 (N_4418,N_3709,N_3800);
and U4419 (N_4419,N_3930,N_3744);
and U4420 (N_4420,N_3511,N_3611);
nand U4421 (N_4421,N_3663,N_3981);
nand U4422 (N_4422,N_3812,N_3967);
or U4423 (N_4423,N_3606,N_3712);
xor U4424 (N_4424,N_3588,N_3954);
xor U4425 (N_4425,N_3510,N_3636);
nor U4426 (N_4426,N_3539,N_3572);
nand U4427 (N_4427,N_3581,N_3516);
nor U4428 (N_4428,N_3510,N_3882);
and U4429 (N_4429,N_3972,N_3607);
and U4430 (N_4430,N_3965,N_3885);
or U4431 (N_4431,N_3795,N_3920);
nand U4432 (N_4432,N_3959,N_3626);
and U4433 (N_4433,N_3851,N_3826);
xor U4434 (N_4434,N_3856,N_3815);
xnor U4435 (N_4435,N_3515,N_3829);
and U4436 (N_4436,N_3847,N_3905);
and U4437 (N_4437,N_3871,N_3839);
or U4438 (N_4438,N_3953,N_3656);
nor U4439 (N_4439,N_3908,N_3750);
nor U4440 (N_4440,N_3535,N_3720);
and U4441 (N_4441,N_3612,N_3876);
nand U4442 (N_4442,N_3634,N_3948);
and U4443 (N_4443,N_3585,N_3581);
nand U4444 (N_4444,N_3820,N_3538);
xnor U4445 (N_4445,N_3535,N_3796);
nand U4446 (N_4446,N_3802,N_3513);
and U4447 (N_4447,N_3569,N_3535);
xnor U4448 (N_4448,N_3675,N_3574);
or U4449 (N_4449,N_3612,N_3735);
or U4450 (N_4450,N_3503,N_3945);
and U4451 (N_4451,N_3913,N_3786);
or U4452 (N_4452,N_3534,N_3535);
xor U4453 (N_4453,N_3928,N_3939);
and U4454 (N_4454,N_3957,N_3850);
nor U4455 (N_4455,N_3667,N_3542);
and U4456 (N_4456,N_3731,N_3983);
xnor U4457 (N_4457,N_3754,N_3572);
nor U4458 (N_4458,N_3624,N_3523);
xnor U4459 (N_4459,N_3596,N_3682);
nand U4460 (N_4460,N_3747,N_3624);
nand U4461 (N_4461,N_3730,N_3594);
nor U4462 (N_4462,N_3527,N_3804);
xnor U4463 (N_4463,N_3529,N_3726);
or U4464 (N_4464,N_3583,N_3652);
or U4465 (N_4465,N_3551,N_3938);
xnor U4466 (N_4466,N_3926,N_3548);
and U4467 (N_4467,N_3840,N_3734);
xor U4468 (N_4468,N_3832,N_3601);
nor U4469 (N_4469,N_3979,N_3532);
xnor U4470 (N_4470,N_3686,N_3609);
xnor U4471 (N_4471,N_3711,N_3969);
nand U4472 (N_4472,N_3714,N_3612);
xnor U4473 (N_4473,N_3524,N_3899);
xor U4474 (N_4474,N_3785,N_3861);
nor U4475 (N_4475,N_3636,N_3895);
and U4476 (N_4476,N_3944,N_3569);
and U4477 (N_4477,N_3602,N_3537);
or U4478 (N_4478,N_3631,N_3956);
nand U4479 (N_4479,N_3515,N_3879);
nor U4480 (N_4480,N_3693,N_3584);
nor U4481 (N_4481,N_3608,N_3558);
nand U4482 (N_4482,N_3853,N_3889);
xor U4483 (N_4483,N_3778,N_3685);
nor U4484 (N_4484,N_3708,N_3627);
and U4485 (N_4485,N_3539,N_3778);
nand U4486 (N_4486,N_3666,N_3734);
or U4487 (N_4487,N_3884,N_3571);
xor U4488 (N_4488,N_3958,N_3757);
xor U4489 (N_4489,N_3843,N_3933);
xor U4490 (N_4490,N_3548,N_3607);
xnor U4491 (N_4491,N_3857,N_3806);
nor U4492 (N_4492,N_3637,N_3869);
nor U4493 (N_4493,N_3816,N_3604);
nor U4494 (N_4494,N_3927,N_3729);
and U4495 (N_4495,N_3598,N_3500);
and U4496 (N_4496,N_3869,N_3904);
and U4497 (N_4497,N_3857,N_3723);
nor U4498 (N_4498,N_3714,N_3530);
or U4499 (N_4499,N_3863,N_3615);
or U4500 (N_4500,N_4280,N_4062);
nand U4501 (N_4501,N_4286,N_4096);
and U4502 (N_4502,N_4180,N_4246);
xnor U4503 (N_4503,N_4453,N_4176);
or U4504 (N_4504,N_4348,N_4224);
and U4505 (N_4505,N_4311,N_4105);
nand U4506 (N_4506,N_4217,N_4335);
or U4507 (N_4507,N_4011,N_4173);
xnor U4508 (N_4508,N_4029,N_4076);
nand U4509 (N_4509,N_4387,N_4287);
nand U4510 (N_4510,N_4263,N_4002);
and U4511 (N_4511,N_4279,N_4141);
nor U4512 (N_4512,N_4075,N_4313);
or U4513 (N_4513,N_4033,N_4168);
nand U4514 (N_4514,N_4393,N_4219);
and U4515 (N_4515,N_4451,N_4183);
xnor U4516 (N_4516,N_4111,N_4237);
or U4517 (N_4517,N_4007,N_4023);
nor U4518 (N_4518,N_4154,N_4157);
and U4519 (N_4519,N_4388,N_4301);
nor U4520 (N_4520,N_4175,N_4347);
and U4521 (N_4521,N_4384,N_4123);
xor U4522 (N_4522,N_4249,N_4350);
or U4523 (N_4523,N_4427,N_4116);
or U4524 (N_4524,N_4412,N_4413);
xor U4525 (N_4525,N_4159,N_4385);
or U4526 (N_4526,N_4245,N_4359);
nand U4527 (N_4527,N_4061,N_4372);
xnor U4528 (N_4528,N_4035,N_4403);
nor U4529 (N_4529,N_4129,N_4333);
nor U4530 (N_4530,N_4461,N_4285);
or U4531 (N_4531,N_4155,N_4079);
xnor U4532 (N_4532,N_4126,N_4468);
xor U4533 (N_4533,N_4356,N_4473);
nor U4534 (N_4534,N_4460,N_4408);
xnor U4535 (N_4535,N_4475,N_4499);
or U4536 (N_4536,N_4143,N_4315);
or U4537 (N_4537,N_4381,N_4124);
nor U4538 (N_4538,N_4277,N_4289);
and U4539 (N_4539,N_4378,N_4088);
xor U4540 (N_4540,N_4373,N_4380);
xnor U4541 (N_4541,N_4272,N_4262);
xor U4542 (N_4542,N_4179,N_4320);
and U4543 (N_4543,N_4095,N_4044);
nor U4544 (N_4544,N_4360,N_4274);
nor U4545 (N_4545,N_4382,N_4165);
and U4546 (N_4546,N_4300,N_4196);
nand U4547 (N_4547,N_4107,N_4034);
and U4548 (N_4548,N_4200,N_4312);
nor U4549 (N_4549,N_4325,N_4156);
xor U4550 (N_4550,N_4045,N_4128);
xnor U4551 (N_4551,N_4308,N_4296);
nor U4552 (N_4552,N_4250,N_4069);
and U4553 (N_4553,N_4243,N_4239);
or U4554 (N_4554,N_4205,N_4085);
xnor U4555 (N_4555,N_4367,N_4115);
and U4556 (N_4556,N_4423,N_4189);
nor U4557 (N_4557,N_4073,N_4486);
or U4558 (N_4558,N_4211,N_4299);
nand U4559 (N_4559,N_4476,N_4055);
nand U4560 (N_4560,N_4112,N_4424);
and U4561 (N_4561,N_4419,N_4125);
or U4562 (N_4562,N_4178,N_4005);
nor U4563 (N_4563,N_4247,N_4471);
or U4564 (N_4564,N_4009,N_4227);
nand U4565 (N_4565,N_4118,N_4036);
xor U4566 (N_4566,N_4188,N_4150);
xor U4567 (N_4567,N_4240,N_4093);
and U4568 (N_4568,N_4317,N_4014);
nand U4569 (N_4569,N_4142,N_4006);
and U4570 (N_4570,N_4420,N_4267);
or U4571 (N_4571,N_4358,N_4341);
and U4572 (N_4572,N_4332,N_4158);
and U4573 (N_4573,N_4092,N_4363);
nand U4574 (N_4574,N_4236,N_4462);
xor U4575 (N_4575,N_4059,N_4162);
and U4576 (N_4576,N_4153,N_4037);
nor U4577 (N_4577,N_4282,N_4307);
xor U4578 (N_4578,N_4192,N_4319);
nand U4579 (N_4579,N_4309,N_4172);
nand U4580 (N_4580,N_4411,N_4106);
nor U4581 (N_4581,N_4397,N_4102);
xor U4582 (N_4582,N_4003,N_4213);
xor U4583 (N_4583,N_4255,N_4013);
nand U4584 (N_4584,N_4422,N_4480);
nor U4585 (N_4585,N_4060,N_4435);
nand U4586 (N_4586,N_4113,N_4264);
nor U4587 (N_4587,N_4483,N_4470);
nand U4588 (N_4588,N_4004,N_4232);
or U4589 (N_4589,N_4104,N_4316);
nor U4590 (N_4590,N_4398,N_4321);
or U4591 (N_4591,N_4138,N_4428);
xor U4592 (N_4592,N_4407,N_4493);
xor U4593 (N_4593,N_4432,N_4099);
xor U4594 (N_4594,N_4357,N_4027);
xnor U4595 (N_4595,N_4310,N_4436);
or U4596 (N_4596,N_4024,N_4489);
or U4597 (N_4597,N_4261,N_4297);
or U4598 (N_4598,N_4064,N_4041);
nand U4599 (N_4599,N_4409,N_4108);
nand U4600 (N_4600,N_4242,N_4230);
nand U4601 (N_4601,N_4117,N_4353);
nor U4602 (N_4602,N_4314,N_4330);
and U4603 (N_4603,N_4140,N_4253);
nand U4604 (N_4604,N_4052,N_4194);
nor U4605 (N_4605,N_4087,N_4038);
nor U4606 (N_4606,N_4049,N_4446);
nand U4607 (N_4607,N_4414,N_4371);
and U4608 (N_4608,N_4342,N_4001);
xnor U4609 (N_4609,N_4438,N_4094);
xor U4610 (N_4610,N_4334,N_4000);
nor U4611 (N_4611,N_4395,N_4229);
nor U4612 (N_4612,N_4210,N_4071);
nand U4613 (N_4613,N_4439,N_4429);
nand U4614 (N_4614,N_4191,N_4131);
nor U4615 (N_4615,N_4120,N_4058);
and U4616 (N_4616,N_4269,N_4295);
nor U4617 (N_4617,N_4271,N_4352);
and U4618 (N_4618,N_4465,N_4083);
xor U4619 (N_4619,N_4195,N_4410);
or U4620 (N_4620,N_4366,N_4455);
nor U4621 (N_4621,N_4235,N_4345);
or U4622 (N_4622,N_4233,N_4127);
nor U4623 (N_4623,N_4097,N_4303);
xor U4624 (N_4624,N_4067,N_4008);
or U4625 (N_4625,N_4268,N_4103);
and U4626 (N_4626,N_4101,N_4441);
nand U4627 (N_4627,N_4349,N_4291);
nor U4628 (N_4628,N_4132,N_4326);
and U4629 (N_4629,N_4053,N_4212);
nor U4630 (N_4630,N_4447,N_4032);
and U4631 (N_4631,N_4169,N_4021);
or U4632 (N_4632,N_4066,N_4238);
and U4633 (N_4633,N_4374,N_4405);
and U4634 (N_4634,N_4077,N_4391);
nor U4635 (N_4635,N_4376,N_4479);
nor U4636 (N_4636,N_4344,N_4415);
nor U4637 (N_4637,N_4361,N_4355);
xor U4638 (N_4638,N_4278,N_4051);
or U4639 (N_4639,N_4478,N_4431);
and U4640 (N_4640,N_4351,N_4221);
nor U4641 (N_4641,N_4495,N_4228);
and U4642 (N_4642,N_4340,N_4260);
nor U4643 (N_4643,N_4456,N_4498);
or U4644 (N_4644,N_4281,N_4474);
xor U4645 (N_4645,N_4134,N_4450);
nand U4646 (N_4646,N_4394,N_4098);
and U4647 (N_4647,N_4327,N_4234);
or U4648 (N_4648,N_4110,N_4458);
xnor U4649 (N_4649,N_4050,N_4084);
nor U4650 (N_4650,N_4399,N_4145);
nand U4651 (N_4651,N_4404,N_4137);
nor U4652 (N_4652,N_4331,N_4026);
nand U4653 (N_4653,N_4294,N_4418);
or U4654 (N_4654,N_4390,N_4089);
and U4655 (N_4655,N_4100,N_4290);
and U4656 (N_4656,N_4302,N_4223);
nand U4657 (N_4657,N_4226,N_4248);
and U4658 (N_4658,N_4186,N_4146);
or U4659 (N_4659,N_4338,N_4421);
or U4660 (N_4660,N_4170,N_4485);
nor U4661 (N_4661,N_4222,N_4204);
nor U4662 (N_4662,N_4121,N_4199);
or U4663 (N_4663,N_4437,N_4063);
and U4664 (N_4664,N_4136,N_4177);
and U4665 (N_4665,N_4028,N_4020);
nand U4666 (N_4666,N_4482,N_4171);
nand U4667 (N_4667,N_4434,N_4257);
nor U4668 (N_4668,N_4392,N_4151);
nand U4669 (N_4669,N_4090,N_4464);
and U4670 (N_4670,N_4417,N_4467);
and U4671 (N_4671,N_4426,N_4369);
xnor U4672 (N_4672,N_4220,N_4364);
and U4673 (N_4673,N_4048,N_4365);
xor U4674 (N_4674,N_4216,N_4074);
nand U4675 (N_4675,N_4270,N_4119);
xor U4676 (N_4676,N_4047,N_4016);
and U4677 (N_4677,N_4133,N_4425);
and U4678 (N_4678,N_4284,N_4368);
nor U4679 (N_4679,N_4144,N_4068);
nor U4680 (N_4680,N_4042,N_4266);
nor U4681 (N_4681,N_4305,N_4244);
xor U4682 (N_4682,N_4491,N_4457);
and U4683 (N_4683,N_4396,N_4275);
and U4684 (N_4684,N_4201,N_4197);
or U4685 (N_4685,N_4207,N_4362);
nor U4686 (N_4686,N_4401,N_4256);
or U4687 (N_4687,N_4402,N_4190);
or U4688 (N_4688,N_4040,N_4182);
nor U4689 (N_4689,N_4383,N_4057);
nor U4690 (N_4690,N_4147,N_4298);
xor U4691 (N_4691,N_4109,N_4185);
or U4692 (N_4692,N_4161,N_4181);
nor U4693 (N_4693,N_4288,N_4046);
or U4694 (N_4694,N_4463,N_4322);
nand U4695 (N_4695,N_4139,N_4377);
or U4696 (N_4696,N_4160,N_4167);
nor U4697 (N_4697,N_4225,N_4148);
and U4698 (N_4698,N_4086,N_4241);
xnor U4699 (N_4699,N_4252,N_4215);
nor U4700 (N_4700,N_4043,N_4163);
xnor U4701 (N_4701,N_4442,N_4487);
nor U4702 (N_4702,N_4494,N_4054);
xor U4703 (N_4703,N_4306,N_4354);
nand U4704 (N_4704,N_4135,N_4452);
and U4705 (N_4705,N_4445,N_4070);
nor U4706 (N_4706,N_4193,N_4273);
or U4707 (N_4707,N_4430,N_4443);
xnor U4708 (N_4708,N_4206,N_4080);
or U4709 (N_4709,N_4448,N_4400);
and U4710 (N_4710,N_4015,N_4440);
or U4711 (N_4711,N_4336,N_4496);
nor U4712 (N_4712,N_4472,N_4454);
xor U4713 (N_4713,N_4488,N_4433);
nor U4714 (N_4714,N_4208,N_4386);
xor U4715 (N_4715,N_4019,N_4081);
nand U4716 (N_4716,N_4346,N_4328);
nor U4717 (N_4717,N_4010,N_4078);
or U4718 (N_4718,N_4304,N_4283);
nor U4719 (N_4719,N_4406,N_4254);
or U4720 (N_4720,N_4072,N_4492);
nand U4721 (N_4721,N_4214,N_4039);
nand U4722 (N_4722,N_4293,N_4469);
or U4723 (N_4723,N_4375,N_4218);
nor U4724 (N_4724,N_4324,N_4318);
and U4725 (N_4725,N_4082,N_4329);
nor U4726 (N_4726,N_4370,N_4018);
nand U4727 (N_4727,N_4209,N_4292);
or U4728 (N_4728,N_4477,N_4481);
xnor U4729 (N_4729,N_4323,N_4203);
nand U4730 (N_4730,N_4466,N_4130);
nand U4731 (N_4731,N_4065,N_4164);
nand U4732 (N_4732,N_4459,N_4231);
nand U4733 (N_4733,N_4258,N_4444);
xnor U4734 (N_4734,N_4114,N_4166);
xor U4735 (N_4735,N_4276,N_4259);
xnor U4736 (N_4736,N_4022,N_4251);
or U4737 (N_4737,N_4122,N_4416);
xnor U4738 (N_4738,N_4265,N_4184);
or U4739 (N_4739,N_4031,N_4030);
xnor U4740 (N_4740,N_4202,N_4343);
xor U4741 (N_4741,N_4149,N_4337);
nand U4742 (N_4742,N_4339,N_4091);
and U4743 (N_4743,N_4152,N_4389);
and U4744 (N_4744,N_4497,N_4490);
xnor U4745 (N_4745,N_4017,N_4025);
nand U4746 (N_4746,N_4187,N_4012);
nand U4747 (N_4747,N_4174,N_4379);
xor U4748 (N_4748,N_4484,N_4056);
nor U4749 (N_4749,N_4198,N_4449);
and U4750 (N_4750,N_4209,N_4377);
xnor U4751 (N_4751,N_4165,N_4186);
and U4752 (N_4752,N_4264,N_4182);
xor U4753 (N_4753,N_4199,N_4404);
and U4754 (N_4754,N_4475,N_4085);
nand U4755 (N_4755,N_4083,N_4430);
nor U4756 (N_4756,N_4036,N_4323);
nand U4757 (N_4757,N_4242,N_4007);
nor U4758 (N_4758,N_4027,N_4288);
xnor U4759 (N_4759,N_4201,N_4499);
and U4760 (N_4760,N_4179,N_4475);
xnor U4761 (N_4761,N_4062,N_4480);
and U4762 (N_4762,N_4088,N_4455);
or U4763 (N_4763,N_4444,N_4282);
nand U4764 (N_4764,N_4049,N_4430);
nor U4765 (N_4765,N_4123,N_4086);
nor U4766 (N_4766,N_4043,N_4419);
or U4767 (N_4767,N_4329,N_4242);
nor U4768 (N_4768,N_4423,N_4490);
xnor U4769 (N_4769,N_4469,N_4487);
and U4770 (N_4770,N_4078,N_4499);
or U4771 (N_4771,N_4258,N_4171);
xor U4772 (N_4772,N_4266,N_4401);
xor U4773 (N_4773,N_4141,N_4077);
and U4774 (N_4774,N_4180,N_4326);
nand U4775 (N_4775,N_4192,N_4228);
xor U4776 (N_4776,N_4119,N_4109);
and U4777 (N_4777,N_4397,N_4310);
xor U4778 (N_4778,N_4010,N_4138);
xor U4779 (N_4779,N_4192,N_4146);
nand U4780 (N_4780,N_4194,N_4004);
and U4781 (N_4781,N_4213,N_4234);
and U4782 (N_4782,N_4271,N_4342);
nor U4783 (N_4783,N_4399,N_4296);
or U4784 (N_4784,N_4442,N_4374);
and U4785 (N_4785,N_4131,N_4354);
or U4786 (N_4786,N_4227,N_4193);
nand U4787 (N_4787,N_4332,N_4134);
or U4788 (N_4788,N_4497,N_4462);
xor U4789 (N_4789,N_4494,N_4126);
nor U4790 (N_4790,N_4021,N_4138);
nor U4791 (N_4791,N_4121,N_4420);
nor U4792 (N_4792,N_4393,N_4045);
and U4793 (N_4793,N_4298,N_4070);
nor U4794 (N_4794,N_4263,N_4133);
nand U4795 (N_4795,N_4033,N_4221);
or U4796 (N_4796,N_4140,N_4044);
nor U4797 (N_4797,N_4340,N_4481);
nor U4798 (N_4798,N_4389,N_4453);
nand U4799 (N_4799,N_4168,N_4297);
nor U4800 (N_4800,N_4174,N_4112);
and U4801 (N_4801,N_4378,N_4472);
or U4802 (N_4802,N_4213,N_4129);
or U4803 (N_4803,N_4109,N_4082);
nand U4804 (N_4804,N_4103,N_4070);
nand U4805 (N_4805,N_4311,N_4301);
nor U4806 (N_4806,N_4056,N_4313);
nand U4807 (N_4807,N_4272,N_4439);
and U4808 (N_4808,N_4058,N_4049);
xor U4809 (N_4809,N_4179,N_4346);
or U4810 (N_4810,N_4237,N_4316);
and U4811 (N_4811,N_4037,N_4363);
and U4812 (N_4812,N_4012,N_4467);
nand U4813 (N_4813,N_4463,N_4058);
and U4814 (N_4814,N_4358,N_4181);
or U4815 (N_4815,N_4152,N_4100);
and U4816 (N_4816,N_4017,N_4262);
nor U4817 (N_4817,N_4081,N_4485);
nor U4818 (N_4818,N_4374,N_4208);
or U4819 (N_4819,N_4268,N_4164);
nand U4820 (N_4820,N_4071,N_4131);
or U4821 (N_4821,N_4315,N_4490);
and U4822 (N_4822,N_4162,N_4038);
and U4823 (N_4823,N_4259,N_4103);
nand U4824 (N_4824,N_4298,N_4491);
xor U4825 (N_4825,N_4284,N_4449);
xnor U4826 (N_4826,N_4134,N_4421);
xnor U4827 (N_4827,N_4065,N_4368);
or U4828 (N_4828,N_4051,N_4090);
and U4829 (N_4829,N_4086,N_4238);
xor U4830 (N_4830,N_4069,N_4461);
nor U4831 (N_4831,N_4082,N_4300);
xor U4832 (N_4832,N_4462,N_4004);
nand U4833 (N_4833,N_4019,N_4004);
nand U4834 (N_4834,N_4203,N_4189);
and U4835 (N_4835,N_4494,N_4065);
nor U4836 (N_4836,N_4221,N_4117);
nand U4837 (N_4837,N_4369,N_4432);
nor U4838 (N_4838,N_4101,N_4418);
or U4839 (N_4839,N_4223,N_4305);
xnor U4840 (N_4840,N_4382,N_4374);
and U4841 (N_4841,N_4406,N_4067);
nor U4842 (N_4842,N_4244,N_4287);
nand U4843 (N_4843,N_4304,N_4141);
nand U4844 (N_4844,N_4028,N_4413);
nor U4845 (N_4845,N_4388,N_4468);
or U4846 (N_4846,N_4336,N_4106);
and U4847 (N_4847,N_4017,N_4400);
or U4848 (N_4848,N_4034,N_4329);
nand U4849 (N_4849,N_4058,N_4056);
nand U4850 (N_4850,N_4099,N_4387);
or U4851 (N_4851,N_4150,N_4045);
nand U4852 (N_4852,N_4343,N_4065);
and U4853 (N_4853,N_4243,N_4064);
and U4854 (N_4854,N_4067,N_4416);
or U4855 (N_4855,N_4488,N_4088);
and U4856 (N_4856,N_4289,N_4307);
nor U4857 (N_4857,N_4211,N_4127);
nand U4858 (N_4858,N_4216,N_4012);
nand U4859 (N_4859,N_4269,N_4079);
or U4860 (N_4860,N_4489,N_4266);
xor U4861 (N_4861,N_4008,N_4127);
or U4862 (N_4862,N_4473,N_4407);
nor U4863 (N_4863,N_4161,N_4490);
nand U4864 (N_4864,N_4417,N_4089);
nand U4865 (N_4865,N_4446,N_4276);
nor U4866 (N_4866,N_4409,N_4073);
or U4867 (N_4867,N_4021,N_4072);
xor U4868 (N_4868,N_4073,N_4414);
and U4869 (N_4869,N_4440,N_4144);
xnor U4870 (N_4870,N_4336,N_4064);
nand U4871 (N_4871,N_4191,N_4422);
xor U4872 (N_4872,N_4034,N_4497);
and U4873 (N_4873,N_4125,N_4472);
nand U4874 (N_4874,N_4053,N_4031);
nor U4875 (N_4875,N_4337,N_4468);
and U4876 (N_4876,N_4377,N_4031);
xnor U4877 (N_4877,N_4295,N_4371);
and U4878 (N_4878,N_4001,N_4458);
or U4879 (N_4879,N_4381,N_4077);
nor U4880 (N_4880,N_4085,N_4310);
nand U4881 (N_4881,N_4022,N_4427);
and U4882 (N_4882,N_4161,N_4397);
nor U4883 (N_4883,N_4140,N_4074);
nand U4884 (N_4884,N_4175,N_4065);
nor U4885 (N_4885,N_4089,N_4275);
and U4886 (N_4886,N_4409,N_4168);
or U4887 (N_4887,N_4233,N_4348);
nor U4888 (N_4888,N_4399,N_4294);
nor U4889 (N_4889,N_4180,N_4026);
nand U4890 (N_4890,N_4343,N_4022);
xor U4891 (N_4891,N_4234,N_4270);
or U4892 (N_4892,N_4484,N_4053);
nand U4893 (N_4893,N_4313,N_4157);
nor U4894 (N_4894,N_4037,N_4358);
nand U4895 (N_4895,N_4453,N_4260);
and U4896 (N_4896,N_4049,N_4157);
xnor U4897 (N_4897,N_4147,N_4352);
nand U4898 (N_4898,N_4349,N_4026);
xor U4899 (N_4899,N_4168,N_4369);
and U4900 (N_4900,N_4012,N_4379);
nand U4901 (N_4901,N_4216,N_4336);
or U4902 (N_4902,N_4016,N_4041);
xnor U4903 (N_4903,N_4279,N_4241);
nor U4904 (N_4904,N_4089,N_4132);
or U4905 (N_4905,N_4071,N_4003);
or U4906 (N_4906,N_4380,N_4103);
xnor U4907 (N_4907,N_4096,N_4244);
and U4908 (N_4908,N_4299,N_4027);
or U4909 (N_4909,N_4325,N_4241);
nor U4910 (N_4910,N_4156,N_4427);
xor U4911 (N_4911,N_4370,N_4440);
nor U4912 (N_4912,N_4114,N_4414);
nand U4913 (N_4913,N_4374,N_4300);
or U4914 (N_4914,N_4499,N_4243);
and U4915 (N_4915,N_4314,N_4475);
xor U4916 (N_4916,N_4070,N_4019);
and U4917 (N_4917,N_4499,N_4238);
xor U4918 (N_4918,N_4409,N_4197);
and U4919 (N_4919,N_4385,N_4215);
and U4920 (N_4920,N_4302,N_4317);
nand U4921 (N_4921,N_4114,N_4120);
nand U4922 (N_4922,N_4036,N_4369);
nand U4923 (N_4923,N_4343,N_4332);
and U4924 (N_4924,N_4074,N_4445);
nor U4925 (N_4925,N_4356,N_4168);
xor U4926 (N_4926,N_4217,N_4496);
xor U4927 (N_4927,N_4417,N_4256);
and U4928 (N_4928,N_4157,N_4031);
nand U4929 (N_4929,N_4052,N_4266);
or U4930 (N_4930,N_4102,N_4211);
or U4931 (N_4931,N_4311,N_4294);
nor U4932 (N_4932,N_4029,N_4077);
nand U4933 (N_4933,N_4063,N_4026);
nor U4934 (N_4934,N_4224,N_4203);
or U4935 (N_4935,N_4483,N_4161);
xor U4936 (N_4936,N_4217,N_4199);
or U4937 (N_4937,N_4358,N_4376);
and U4938 (N_4938,N_4438,N_4080);
and U4939 (N_4939,N_4301,N_4379);
nand U4940 (N_4940,N_4151,N_4159);
or U4941 (N_4941,N_4366,N_4022);
or U4942 (N_4942,N_4323,N_4028);
nand U4943 (N_4943,N_4160,N_4472);
nand U4944 (N_4944,N_4041,N_4435);
or U4945 (N_4945,N_4088,N_4349);
or U4946 (N_4946,N_4182,N_4416);
nor U4947 (N_4947,N_4478,N_4128);
xor U4948 (N_4948,N_4156,N_4134);
xnor U4949 (N_4949,N_4218,N_4062);
nor U4950 (N_4950,N_4246,N_4418);
or U4951 (N_4951,N_4204,N_4124);
nand U4952 (N_4952,N_4185,N_4222);
and U4953 (N_4953,N_4178,N_4333);
nor U4954 (N_4954,N_4152,N_4179);
xor U4955 (N_4955,N_4249,N_4389);
nor U4956 (N_4956,N_4338,N_4369);
xnor U4957 (N_4957,N_4107,N_4310);
or U4958 (N_4958,N_4072,N_4215);
nor U4959 (N_4959,N_4182,N_4171);
or U4960 (N_4960,N_4219,N_4100);
or U4961 (N_4961,N_4196,N_4467);
nand U4962 (N_4962,N_4473,N_4104);
or U4963 (N_4963,N_4216,N_4289);
and U4964 (N_4964,N_4135,N_4033);
nor U4965 (N_4965,N_4406,N_4342);
nand U4966 (N_4966,N_4433,N_4469);
or U4967 (N_4967,N_4439,N_4009);
and U4968 (N_4968,N_4255,N_4227);
nand U4969 (N_4969,N_4051,N_4281);
xor U4970 (N_4970,N_4239,N_4223);
and U4971 (N_4971,N_4274,N_4021);
and U4972 (N_4972,N_4445,N_4250);
nor U4973 (N_4973,N_4173,N_4136);
and U4974 (N_4974,N_4269,N_4420);
and U4975 (N_4975,N_4006,N_4169);
nand U4976 (N_4976,N_4442,N_4326);
xnor U4977 (N_4977,N_4356,N_4222);
and U4978 (N_4978,N_4033,N_4152);
xor U4979 (N_4979,N_4110,N_4372);
and U4980 (N_4980,N_4448,N_4382);
nor U4981 (N_4981,N_4364,N_4323);
nand U4982 (N_4982,N_4392,N_4443);
nand U4983 (N_4983,N_4323,N_4152);
nand U4984 (N_4984,N_4070,N_4336);
xnor U4985 (N_4985,N_4410,N_4032);
nor U4986 (N_4986,N_4215,N_4074);
or U4987 (N_4987,N_4435,N_4280);
nor U4988 (N_4988,N_4291,N_4404);
nor U4989 (N_4989,N_4301,N_4213);
xor U4990 (N_4990,N_4184,N_4250);
nor U4991 (N_4991,N_4383,N_4266);
nor U4992 (N_4992,N_4271,N_4404);
nand U4993 (N_4993,N_4233,N_4241);
nor U4994 (N_4994,N_4277,N_4295);
xor U4995 (N_4995,N_4062,N_4077);
or U4996 (N_4996,N_4039,N_4447);
nor U4997 (N_4997,N_4162,N_4236);
nor U4998 (N_4998,N_4096,N_4168);
xor U4999 (N_4999,N_4386,N_4094);
nor U5000 (N_5000,N_4628,N_4903);
nor U5001 (N_5001,N_4834,N_4641);
or U5002 (N_5002,N_4572,N_4924);
nor U5003 (N_5003,N_4993,N_4828);
and U5004 (N_5004,N_4700,N_4586);
xor U5005 (N_5005,N_4733,N_4520);
or U5006 (N_5006,N_4537,N_4593);
and U5007 (N_5007,N_4670,N_4772);
nor U5008 (N_5008,N_4998,N_4757);
xnor U5009 (N_5009,N_4879,N_4944);
or U5010 (N_5010,N_4697,N_4888);
or U5011 (N_5011,N_4929,N_4869);
or U5012 (N_5012,N_4878,N_4827);
nand U5013 (N_5013,N_4769,N_4590);
or U5014 (N_5014,N_4504,N_4802);
nand U5015 (N_5015,N_4809,N_4594);
xor U5016 (N_5016,N_4626,N_4996);
nor U5017 (N_5017,N_4574,N_4543);
and U5018 (N_5018,N_4611,N_4730);
or U5019 (N_5019,N_4844,N_4583);
and U5020 (N_5020,N_4814,N_4560);
xnor U5021 (N_5021,N_4555,N_4618);
xor U5022 (N_5022,N_4876,N_4692);
and U5023 (N_5023,N_4835,N_4523);
and U5024 (N_5024,N_4542,N_4801);
and U5025 (N_5025,N_4660,N_4630);
nor U5026 (N_5026,N_4875,N_4767);
xnor U5027 (N_5027,N_4860,N_4525);
and U5028 (N_5028,N_4535,N_4912);
xor U5029 (N_5029,N_4620,N_4527);
nor U5030 (N_5030,N_4779,N_4857);
xnor U5031 (N_5031,N_4717,N_4647);
or U5032 (N_5032,N_4976,N_4732);
or U5033 (N_5033,N_4648,N_4868);
xnor U5034 (N_5034,N_4665,N_4913);
xnor U5035 (N_5035,N_4679,N_4725);
xor U5036 (N_5036,N_4710,N_4643);
and U5037 (N_5037,N_4726,N_4663);
xor U5038 (N_5038,N_4877,N_4753);
or U5039 (N_5039,N_4724,N_4926);
nor U5040 (N_5040,N_4609,N_4515);
xnor U5041 (N_5041,N_4962,N_4920);
or U5042 (N_5042,N_4748,N_4536);
nor U5043 (N_5043,N_4681,N_4501);
nor U5044 (N_5044,N_4738,N_4969);
or U5045 (N_5045,N_4608,N_4659);
nand U5046 (N_5046,N_4902,N_4634);
xnor U5047 (N_5047,N_4636,N_4615);
and U5048 (N_5048,N_4874,N_4723);
or U5049 (N_5049,N_4596,N_4921);
nand U5050 (N_5050,N_4999,N_4745);
or U5051 (N_5051,N_4683,N_4990);
nand U5052 (N_5052,N_4581,N_4949);
nor U5053 (N_5053,N_4882,N_4736);
or U5054 (N_5054,N_4642,N_4919);
xor U5055 (N_5055,N_4832,N_4859);
or U5056 (N_5056,N_4526,N_4896);
xnor U5057 (N_5057,N_4598,N_4904);
xnor U5058 (N_5058,N_4770,N_4908);
and U5059 (N_5059,N_4979,N_4631);
and U5060 (N_5060,N_4833,N_4782);
or U5061 (N_5061,N_4972,N_4507);
xnor U5062 (N_5062,N_4780,N_4985);
or U5063 (N_5063,N_4553,N_4592);
nor U5064 (N_5064,N_4629,N_4939);
and U5065 (N_5065,N_4941,N_4807);
nand U5066 (N_5066,N_4855,N_4865);
and U5067 (N_5067,N_4668,N_4777);
nor U5068 (N_5068,N_4749,N_4937);
xnor U5069 (N_5069,N_4691,N_4811);
nor U5070 (N_5070,N_4587,N_4701);
xor U5071 (N_5071,N_4530,N_4933);
xnor U5072 (N_5072,N_4940,N_4714);
and U5073 (N_5073,N_4931,N_4722);
nand U5074 (N_5074,N_4682,N_4644);
or U5075 (N_5075,N_4699,N_4974);
or U5076 (N_5076,N_4971,N_4565);
nor U5077 (N_5077,N_4640,N_4787);
or U5078 (N_5078,N_4823,N_4545);
xnor U5079 (N_5079,N_4562,N_4977);
nor U5080 (N_5080,N_4754,N_4584);
xnor U5081 (N_5081,N_4915,N_4622);
xnor U5082 (N_5082,N_4747,N_4961);
and U5083 (N_5083,N_4975,N_4863);
or U5084 (N_5084,N_4597,N_4804);
or U5085 (N_5085,N_4705,N_4702);
and U5086 (N_5086,N_4667,N_4610);
or U5087 (N_5087,N_4824,N_4656);
nand U5088 (N_5088,N_4651,N_4694);
nor U5089 (N_5089,N_4517,N_4817);
nand U5090 (N_5090,N_4711,N_4946);
or U5091 (N_5091,N_4649,N_4718);
nor U5092 (N_5092,N_4664,N_4843);
nand U5093 (N_5093,N_4938,N_4698);
xor U5094 (N_5094,N_4576,N_4816);
or U5095 (N_5095,N_4554,N_4819);
nor U5096 (N_5096,N_4883,N_4935);
and U5097 (N_5097,N_4911,N_4778);
nor U5098 (N_5098,N_4546,N_4632);
nor U5099 (N_5099,N_4830,N_4708);
and U5100 (N_5100,N_4842,N_4513);
and U5101 (N_5101,N_4502,N_4715);
and U5102 (N_5102,N_4740,N_4564);
and U5103 (N_5103,N_4758,N_4529);
or U5104 (N_5104,N_4541,N_4764);
nor U5105 (N_5105,N_4791,N_4989);
xor U5106 (N_5106,N_4760,N_4957);
nand U5107 (N_5107,N_4947,N_4930);
nand U5108 (N_5108,N_4783,N_4897);
or U5109 (N_5109,N_4788,N_4739);
nand U5110 (N_5110,N_4964,N_4800);
and U5111 (N_5111,N_4968,N_4601);
and U5112 (N_5112,N_4959,N_4812);
nand U5113 (N_5113,N_4614,N_4786);
nor U5114 (N_5114,N_4591,N_4559);
xnor U5115 (N_5115,N_4885,N_4567);
nor U5116 (N_5116,N_4566,N_4988);
nand U5117 (N_5117,N_4943,N_4666);
and U5118 (N_5118,N_4849,N_4704);
xor U5119 (N_5119,N_4687,N_4728);
xnor U5120 (N_5120,N_4625,N_4552);
and U5121 (N_5121,N_4646,N_4785);
nand U5122 (N_5122,N_4673,N_4890);
nor U5123 (N_5123,N_4942,N_4602);
and U5124 (N_5124,N_4661,N_4690);
nor U5125 (N_5125,N_4936,N_4895);
nand U5126 (N_5126,N_4674,N_4680);
and U5127 (N_5127,N_4508,N_4509);
nand U5128 (N_5128,N_4900,N_4752);
and U5129 (N_5129,N_4803,N_4645);
xor U5130 (N_5130,N_4635,N_4505);
nand U5131 (N_5131,N_4899,N_4599);
and U5132 (N_5132,N_4578,N_4612);
xnor U5133 (N_5133,N_4893,N_4870);
nor U5134 (N_5134,N_4506,N_4986);
and U5135 (N_5135,N_4677,N_4831);
and U5136 (N_5136,N_4538,N_4652);
and U5137 (N_5137,N_4846,N_4925);
nand U5138 (N_5138,N_4881,N_4952);
and U5139 (N_5139,N_4540,N_4751);
or U5140 (N_5140,N_4798,N_4633);
nor U5141 (N_5141,N_4512,N_4503);
nor U5142 (N_5142,N_4675,N_4838);
and U5143 (N_5143,N_4954,N_4991);
or U5144 (N_5144,N_4514,N_4982);
nor U5145 (N_5145,N_4826,N_4686);
xnor U5146 (N_5146,N_4852,N_4637);
nand U5147 (N_5147,N_4746,N_4638);
nand U5148 (N_5148,N_4500,N_4556);
xor U5149 (N_5149,N_4889,N_4918);
or U5150 (N_5150,N_4923,N_4573);
or U5151 (N_5151,N_4729,N_4678);
nand U5152 (N_5152,N_4789,N_4624);
nor U5153 (N_5153,N_4695,N_4953);
nand U5154 (N_5154,N_4582,N_4856);
nor U5155 (N_5155,N_4676,N_4966);
nor U5156 (N_5156,N_4534,N_4524);
or U5157 (N_5157,N_4914,N_4539);
and U5158 (N_5158,N_4588,N_4922);
or U5159 (N_5159,N_4887,N_4706);
nor U5160 (N_5160,N_4518,N_4808);
or U5161 (N_5161,N_4848,N_4685);
xor U5162 (N_5162,N_4841,N_4821);
xor U5163 (N_5163,N_4776,N_4984);
and U5164 (N_5164,N_4796,N_4873);
nand U5165 (N_5165,N_4616,N_4750);
xor U5166 (N_5166,N_4766,N_4847);
nand U5167 (N_5167,N_4763,N_4579);
or U5168 (N_5168,N_4575,N_4654);
xor U5169 (N_5169,N_4532,N_4557);
and U5170 (N_5170,N_4519,N_4916);
xor U5171 (N_5171,N_4605,N_4910);
xor U5172 (N_5172,N_4773,N_4765);
or U5173 (N_5173,N_4741,N_4669);
nor U5174 (N_5174,N_4528,N_4511);
nor U5175 (N_5175,N_4837,N_4853);
nor U5176 (N_5176,N_4805,N_4716);
nor U5177 (N_5177,N_4547,N_4619);
nor U5178 (N_5178,N_4713,N_4688);
nand U5179 (N_5179,N_4737,N_4898);
nor U5180 (N_5180,N_4613,N_4712);
or U5181 (N_5181,N_4549,N_4603);
and U5182 (N_5182,N_4840,N_4983);
and U5183 (N_5183,N_4662,N_4797);
nor U5184 (N_5184,N_4759,N_4871);
or U5185 (N_5185,N_4994,N_4799);
or U5186 (N_5186,N_4522,N_4658);
nor U5187 (N_5187,N_4995,N_4815);
xor U5188 (N_5188,N_4951,N_4720);
and U5189 (N_5189,N_4550,N_4719);
nor U5190 (N_5190,N_4606,N_4531);
nand U5191 (N_5191,N_4570,N_4784);
or U5192 (N_5192,N_4639,N_4987);
or U5193 (N_5193,N_4934,N_4568);
and U5194 (N_5194,N_4703,N_4945);
and U5195 (N_5195,N_4905,N_4696);
and U5196 (N_5196,N_4854,N_4978);
xnor U5197 (N_5197,N_4861,N_4607);
and U5198 (N_5198,N_4761,N_4617);
nand U5199 (N_5199,N_4810,N_4650);
nor U5200 (N_5200,N_4781,N_4981);
and U5201 (N_5201,N_4901,N_4735);
or U5202 (N_5202,N_4839,N_4992);
and U5203 (N_5203,N_4762,N_4533);
and U5204 (N_5204,N_4820,N_4891);
xor U5205 (N_5205,N_4756,N_4774);
or U5206 (N_5206,N_4672,N_4742);
nand U5207 (N_5207,N_4707,N_4963);
nor U5208 (N_5208,N_4689,N_4755);
and U5209 (N_5209,N_4721,N_4653);
nor U5210 (N_5210,N_4768,N_4866);
and U5211 (N_5211,N_4806,N_4825);
xor U5212 (N_5212,N_4544,N_4822);
xnor U5213 (N_5213,N_4932,N_4892);
xnor U5214 (N_5214,N_4948,N_4850);
nand U5215 (N_5215,N_4967,N_4950);
or U5216 (N_5216,N_4958,N_4864);
nor U5217 (N_5217,N_4793,N_4973);
and U5218 (N_5218,N_4862,N_4600);
and U5219 (N_5219,N_4884,N_4775);
or U5220 (N_5220,N_4551,N_4548);
nor U5221 (N_5221,N_4693,N_4595);
xor U5222 (N_5222,N_4970,N_4709);
nand U5223 (N_5223,N_4627,N_4684);
or U5224 (N_5224,N_4561,N_4795);
nand U5225 (N_5225,N_4909,N_4955);
or U5226 (N_5226,N_4563,N_4965);
or U5227 (N_5227,N_4997,N_4960);
nand U5228 (N_5228,N_4858,N_4577);
nor U5229 (N_5229,N_4851,N_4907);
xnor U5230 (N_5230,N_4794,N_4818);
and U5231 (N_5231,N_4872,N_4790);
and U5232 (N_5232,N_4569,N_4906);
and U5233 (N_5233,N_4867,N_4928);
xor U5234 (N_5234,N_4623,N_4894);
nor U5235 (N_5235,N_4731,N_4657);
and U5236 (N_5236,N_4845,N_4829);
xnor U5237 (N_5237,N_4743,N_4880);
nor U5238 (N_5238,N_4516,N_4836);
nor U5239 (N_5239,N_4744,N_4727);
or U5240 (N_5240,N_4886,N_4585);
nor U5241 (N_5241,N_4604,N_4771);
nand U5242 (N_5242,N_4734,N_4621);
and U5243 (N_5243,N_4521,N_4980);
or U5244 (N_5244,N_4510,N_4792);
nand U5245 (N_5245,N_4927,N_4571);
nand U5246 (N_5246,N_4558,N_4917);
and U5247 (N_5247,N_4956,N_4655);
xor U5248 (N_5248,N_4580,N_4813);
xor U5249 (N_5249,N_4671,N_4589);
and U5250 (N_5250,N_4961,N_4581);
nor U5251 (N_5251,N_4957,N_4713);
or U5252 (N_5252,N_4936,N_4618);
nor U5253 (N_5253,N_4811,N_4640);
xnor U5254 (N_5254,N_4583,N_4719);
and U5255 (N_5255,N_4519,N_4546);
nor U5256 (N_5256,N_4828,N_4947);
nand U5257 (N_5257,N_4521,N_4643);
xor U5258 (N_5258,N_4757,N_4892);
xor U5259 (N_5259,N_4756,N_4683);
xor U5260 (N_5260,N_4672,N_4949);
xor U5261 (N_5261,N_4752,N_4615);
xnor U5262 (N_5262,N_4629,N_4635);
nor U5263 (N_5263,N_4959,N_4916);
and U5264 (N_5264,N_4911,N_4792);
nand U5265 (N_5265,N_4715,N_4817);
or U5266 (N_5266,N_4982,N_4930);
nand U5267 (N_5267,N_4765,N_4606);
nand U5268 (N_5268,N_4847,N_4719);
nor U5269 (N_5269,N_4715,N_4643);
or U5270 (N_5270,N_4563,N_4693);
and U5271 (N_5271,N_4838,N_4948);
nand U5272 (N_5272,N_4537,N_4877);
and U5273 (N_5273,N_4747,N_4533);
and U5274 (N_5274,N_4689,N_4715);
nand U5275 (N_5275,N_4779,N_4540);
nor U5276 (N_5276,N_4771,N_4791);
or U5277 (N_5277,N_4988,N_4509);
xnor U5278 (N_5278,N_4542,N_4848);
xnor U5279 (N_5279,N_4611,N_4913);
or U5280 (N_5280,N_4522,N_4896);
and U5281 (N_5281,N_4759,N_4951);
nor U5282 (N_5282,N_4882,N_4713);
nand U5283 (N_5283,N_4808,N_4605);
or U5284 (N_5284,N_4806,N_4993);
xnor U5285 (N_5285,N_4510,N_4951);
nand U5286 (N_5286,N_4921,N_4710);
or U5287 (N_5287,N_4607,N_4986);
xnor U5288 (N_5288,N_4676,N_4968);
xor U5289 (N_5289,N_4998,N_4921);
and U5290 (N_5290,N_4616,N_4780);
nand U5291 (N_5291,N_4565,N_4873);
or U5292 (N_5292,N_4737,N_4920);
and U5293 (N_5293,N_4734,N_4745);
nor U5294 (N_5294,N_4809,N_4833);
nand U5295 (N_5295,N_4951,N_4523);
or U5296 (N_5296,N_4733,N_4903);
and U5297 (N_5297,N_4766,N_4773);
nor U5298 (N_5298,N_4759,N_4548);
or U5299 (N_5299,N_4835,N_4988);
xnor U5300 (N_5300,N_4900,N_4883);
and U5301 (N_5301,N_4816,N_4691);
nor U5302 (N_5302,N_4707,N_4552);
nand U5303 (N_5303,N_4947,N_4580);
and U5304 (N_5304,N_4637,N_4920);
xor U5305 (N_5305,N_4548,N_4876);
nand U5306 (N_5306,N_4957,N_4949);
nand U5307 (N_5307,N_4866,N_4762);
or U5308 (N_5308,N_4855,N_4561);
nor U5309 (N_5309,N_4841,N_4663);
xor U5310 (N_5310,N_4979,N_4985);
xor U5311 (N_5311,N_4836,N_4556);
nor U5312 (N_5312,N_4770,N_4709);
xnor U5313 (N_5313,N_4568,N_4584);
nor U5314 (N_5314,N_4578,N_4763);
or U5315 (N_5315,N_4906,N_4605);
nand U5316 (N_5316,N_4652,N_4531);
or U5317 (N_5317,N_4703,N_4847);
xnor U5318 (N_5318,N_4852,N_4533);
xor U5319 (N_5319,N_4626,N_4533);
xor U5320 (N_5320,N_4986,N_4543);
or U5321 (N_5321,N_4953,N_4996);
xor U5322 (N_5322,N_4974,N_4933);
xor U5323 (N_5323,N_4964,N_4644);
nor U5324 (N_5324,N_4547,N_4715);
nor U5325 (N_5325,N_4896,N_4917);
or U5326 (N_5326,N_4714,N_4554);
nor U5327 (N_5327,N_4576,N_4660);
or U5328 (N_5328,N_4994,N_4554);
and U5329 (N_5329,N_4944,N_4928);
or U5330 (N_5330,N_4921,N_4976);
nor U5331 (N_5331,N_4643,N_4862);
xor U5332 (N_5332,N_4853,N_4999);
and U5333 (N_5333,N_4504,N_4521);
nand U5334 (N_5334,N_4709,N_4740);
and U5335 (N_5335,N_4905,N_4890);
xnor U5336 (N_5336,N_4622,N_4994);
and U5337 (N_5337,N_4576,N_4541);
nor U5338 (N_5338,N_4828,N_4959);
nor U5339 (N_5339,N_4851,N_4772);
or U5340 (N_5340,N_4926,N_4832);
and U5341 (N_5341,N_4914,N_4560);
and U5342 (N_5342,N_4783,N_4823);
nand U5343 (N_5343,N_4691,N_4797);
and U5344 (N_5344,N_4619,N_4707);
nand U5345 (N_5345,N_4722,N_4598);
and U5346 (N_5346,N_4708,N_4883);
and U5347 (N_5347,N_4977,N_4618);
xor U5348 (N_5348,N_4927,N_4742);
and U5349 (N_5349,N_4733,N_4864);
or U5350 (N_5350,N_4682,N_4622);
or U5351 (N_5351,N_4736,N_4827);
or U5352 (N_5352,N_4538,N_4707);
nand U5353 (N_5353,N_4599,N_4640);
and U5354 (N_5354,N_4950,N_4956);
nand U5355 (N_5355,N_4824,N_4751);
xor U5356 (N_5356,N_4861,N_4670);
xor U5357 (N_5357,N_4629,N_4884);
and U5358 (N_5358,N_4627,N_4613);
xor U5359 (N_5359,N_4650,N_4823);
nand U5360 (N_5360,N_4981,N_4638);
nor U5361 (N_5361,N_4805,N_4845);
or U5362 (N_5362,N_4665,N_4732);
or U5363 (N_5363,N_4528,N_4846);
and U5364 (N_5364,N_4997,N_4595);
nand U5365 (N_5365,N_4637,N_4651);
nor U5366 (N_5366,N_4918,N_4551);
nor U5367 (N_5367,N_4867,N_4974);
or U5368 (N_5368,N_4691,N_4900);
and U5369 (N_5369,N_4978,N_4986);
nor U5370 (N_5370,N_4837,N_4729);
nor U5371 (N_5371,N_4674,N_4924);
nor U5372 (N_5372,N_4686,N_4589);
nand U5373 (N_5373,N_4892,N_4827);
nand U5374 (N_5374,N_4679,N_4877);
and U5375 (N_5375,N_4528,N_4597);
nand U5376 (N_5376,N_4655,N_4921);
and U5377 (N_5377,N_4980,N_4593);
xor U5378 (N_5378,N_4795,N_4737);
xnor U5379 (N_5379,N_4704,N_4785);
and U5380 (N_5380,N_4720,N_4638);
or U5381 (N_5381,N_4944,N_4903);
and U5382 (N_5382,N_4760,N_4799);
xnor U5383 (N_5383,N_4757,N_4932);
xor U5384 (N_5384,N_4922,N_4535);
xnor U5385 (N_5385,N_4614,N_4930);
or U5386 (N_5386,N_4983,N_4852);
nor U5387 (N_5387,N_4935,N_4950);
nor U5388 (N_5388,N_4936,N_4953);
or U5389 (N_5389,N_4544,N_4848);
or U5390 (N_5390,N_4843,N_4950);
or U5391 (N_5391,N_4940,N_4750);
or U5392 (N_5392,N_4683,N_4696);
nand U5393 (N_5393,N_4811,N_4837);
xor U5394 (N_5394,N_4878,N_4893);
nand U5395 (N_5395,N_4626,N_4565);
or U5396 (N_5396,N_4959,N_4598);
nand U5397 (N_5397,N_4528,N_4951);
and U5398 (N_5398,N_4867,N_4805);
and U5399 (N_5399,N_4675,N_4713);
and U5400 (N_5400,N_4708,N_4625);
or U5401 (N_5401,N_4884,N_4859);
or U5402 (N_5402,N_4887,N_4741);
nand U5403 (N_5403,N_4928,N_4646);
xnor U5404 (N_5404,N_4936,N_4796);
and U5405 (N_5405,N_4824,N_4834);
nor U5406 (N_5406,N_4659,N_4898);
or U5407 (N_5407,N_4787,N_4840);
or U5408 (N_5408,N_4831,N_4628);
xnor U5409 (N_5409,N_4887,N_4960);
and U5410 (N_5410,N_4733,N_4538);
xor U5411 (N_5411,N_4655,N_4710);
nand U5412 (N_5412,N_4809,N_4634);
or U5413 (N_5413,N_4856,N_4765);
or U5414 (N_5414,N_4634,N_4886);
or U5415 (N_5415,N_4660,N_4927);
nand U5416 (N_5416,N_4650,N_4791);
nor U5417 (N_5417,N_4808,N_4782);
xnor U5418 (N_5418,N_4666,N_4859);
nor U5419 (N_5419,N_4760,N_4763);
xnor U5420 (N_5420,N_4586,N_4719);
and U5421 (N_5421,N_4653,N_4937);
or U5422 (N_5422,N_4566,N_4852);
nand U5423 (N_5423,N_4587,N_4794);
nand U5424 (N_5424,N_4793,N_4685);
xor U5425 (N_5425,N_4703,N_4849);
nand U5426 (N_5426,N_4563,N_4900);
nor U5427 (N_5427,N_4960,N_4942);
or U5428 (N_5428,N_4541,N_4530);
nand U5429 (N_5429,N_4743,N_4905);
xnor U5430 (N_5430,N_4623,N_4656);
nand U5431 (N_5431,N_4618,N_4512);
nor U5432 (N_5432,N_4543,N_4729);
nand U5433 (N_5433,N_4853,N_4974);
nor U5434 (N_5434,N_4844,N_4723);
nor U5435 (N_5435,N_4877,N_4924);
nor U5436 (N_5436,N_4840,N_4767);
nand U5437 (N_5437,N_4942,N_4500);
or U5438 (N_5438,N_4608,N_4648);
nand U5439 (N_5439,N_4746,N_4800);
nor U5440 (N_5440,N_4616,N_4690);
or U5441 (N_5441,N_4776,N_4652);
nor U5442 (N_5442,N_4601,N_4729);
or U5443 (N_5443,N_4712,N_4617);
nand U5444 (N_5444,N_4887,N_4983);
xor U5445 (N_5445,N_4997,N_4998);
and U5446 (N_5446,N_4693,N_4724);
or U5447 (N_5447,N_4650,N_4722);
xor U5448 (N_5448,N_4509,N_4684);
and U5449 (N_5449,N_4745,N_4981);
nand U5450 (N_5450,N_4769,N_4525);
xor U5451 (N_5451,N_4605,N_4834);
and U5452 (N_5452,N_4820,N_4501);
nor U5453 (N_5453,N_4879,N_4702);
and U5454 (N_5454,N_4616,N_4781);
and U5455 (N_5455,N_4893,N_4767);
and U5456 (N_5456,N_4960,N_4949);
nor U5457 (N_5457,N_4803,N_4581);
nand U5458 (N_5458,N_4784,N_4650);
or U5459 (N_5459,N_4795,N_4855);
nor U5460 (N_5460,N_4578,N_4757);
and U5461 (N_5461,N_4560,N_4686);
or U5462 (N_5462,N_4527,N_4804);
nor U5463 (N_5463,N_4562,N_4990);
xor U5464 (N_5464,N_4775,N_4727);
nor U5465 (N_5465,N_4535,N_4910);
or U5466 (N_5466,N_4895,N_4982);
nor U5467 (N_5467,N_4618,N_4607);
or U5468 (N_5468,N_4656,N_4709);
nand U5469 (N_5469,N_4586,N_4500);
nand U5470 (N_5470,N_4584,N_4625);
xor U5471 (N_5471,N_4851,N_4969);
nand U5472 (N_5472,N_4544,N_4524);
or U5473 (N_5473,N_4557,N_4594);
or U5474 (N_5474,N_4664,N_4728);
and U5475 (N_5475,N_4877,N_4614);
nor U5476 (N_5476,N_4885,N_4880);
xor U5477 (N_5477,N_4613,N_4990);
nand U5478 (N_5478,N_4946,N_4618);
and U5479 (N_5479,N_4876,N_4913);
nand U5480 (N_5480,N_4785,N_4544);
nor U5481 (N_5481,N_4647,N_4943);
or U5482 (N_5482,N_4518,N_4576);
or U5483 (N_5483,N_4506,N_4569);
nand U5484 (N_5484,N_4955,N_4941);
or U5485 (N_5485,N_4676,N_4599);
or U5486 (N_5486,N_4880,N_4676);
nand U5487 (N_5487,N_4921,N_4553);
nor U5488 (N_5488,N_4757,N_4563);
and U5489 (N_5489,N_4971,N_4517);
nor U5490 (N_5490,N_4588,N_4698);
and U5491 (N_5491,N_4795,N_4809);
and U5492 (N_5492,N_4782,N_4797);
or U5493 (N_5493,N_4595,N_4631);
nand U5494 (N_5494,N_4807,N_4551);
and U5495 (N_5495,N_4714,N_4612);
xor U5496 (N_5496,N_4722,N_4961);
xnor U5497 (N_5497,N_4600,N_4895);
nand U5498 (N_5498,N_4677,N_4689);
nand U5499 (N_5499,N_4808,N_4841);
or U5500 (N_5500,N_5256,N_5166);
xor U5501 (N_5501,N_5091,N_5325);
xor U5502 (N_5502,N_5261,N_5454);
or U5503 (N_5503,N_5418,N_5046);
or U5504 (N_5504,N_5191,N_5410);
nand U5505 (N_5505,N_5376,N_5407);
nor U5506 (N_5506,N_5182,N_5270);
nand U5507 (N_5507,N_5035,N_5496);
or U5508 (N_5508,N_5115,N_5415);
nor U5509 (N_5509,N_5289,N_5312);
nand U5510 (N_5510,N_5277,N_5023);
nor U5511 (N_5511,N_5252,N_5194);
and U5512 (N_5512,N_5498,N_5017);
or U5513 (N_5513,N_5335,N_5127);
nand U5514 (N_5514,N_5011,N_5111);
and U5515 (N_5515,N_5220,N_5374);
nor U5516 (N_5516,N_5026,N_5358);
and U5517 (N_5517,N_5329,N_5367);
nand U5518 (N_5518,N_5061,N_5467);
and U5519 (N_5519,N_5390,N_5002);
and U5520 (N_5520,N_5004,N_5196);
nand U5521 (N_5521,N_5079,N_5269);
nand U5522 (N_5522,N_5326,N_5014);
xor U5523 (N_5523,N_5413,N_5143);
nor U5524 (N_5524,N_5207,N_5200);
and U5525 (N_5525,N_5491,N_5223);
or U5526 (N_5526,N_5279,N_5040);
or U5527 (N_5527,N_5384,N_5487);
or U5528 (N_5528,N_5016,N_5007);
xnor U5529 (N_5529,N_5424,N_5118);
or U5530 (N_5530,N_5383,N_5055);
or U5531 (N_5531,N_5113,N_5402);
xnor U5532 (N_5532,N_5062,N_5226);
and U5533 (N_5533,N_5097,N_5259);
and U5534 (N_5534,N_5396,N_5343);
or U5535 (N_5535,N_5032,N_5419);
nand U5536 (N_5536,N_5034,N_5095);
nand U5537 (N_5537,N_5075,N_5398);
nor U5538 (N_5538,N_5400,N_5368);
and U5539 (N_5539,N_5492,N_5020);
and U5540 (N_5540,N_5485,N_5058);
nor U5541 (N_5541,N_5322,N_5109);
xor U5542 (N_5542,N_5070,N_5336);
or U5543 (N_5543,N_5015,N_5059);
and U5544 (N_5544,N_5077,N_5481);
nor U5545 (N_5545,N_5366,N_5029);
and U5546 (N_5546,N_5484,N_5489);
xor U5547 (N_5547,N_5137,N_5170);
nor U5548 (N_5548,N_5293,N_5294);
nor U5549 (N_5549,N_5445,N_5010);
or U5550 (N_5550,N_5250,N_5416);
xnor U5551 (N_5551,N_5102,N_5056);
and U5552 (N_5552,N_5320,N_5169);
nand U5553 (N_5553,N_5447,N_5262);
nand U5554 (N_5554,N_5060,N_5180);
nor U5555 (N_5555,N_5126,N_5443);
nor U5556 (N_5556,N_5100,N_5471);
nor U5557 (N_5557,N_5494,N_5309);
xor U5558 (N_5558,N_5231,N_5209);
and U5559 (N_5559,N_5080,N_5283);
nand U5560 (N_5560,N_5131,N_5296);
xor U5561 (N_5561,N_5244,N_5064);
or U5562 (N_5562,N_5006,N_5151);
xor U5563 (N_5563,N_5328,N_5455);
and U5564 (N_5564,N_5292,N_5462);
nor U5565 (N_5565,N_5409,N_5371);
xnor U5566 (N_5566,N_5202,N_5365);
and U5567 (N_5567,N_5159,N_5218);
and U5568 (N_5568,N_5355,N_5225);
and U5569 (N_5569,N_5266,N_5043);
or U5570 (N_5570,N_5315,N_5473);
nand U5571 (N_5571,N_5307,N_5162);
or U5572 (N_5572,N_5107,N_5360);
and U5573 (N_5573,N_5123,N_5213);
nor U5574 (N_5574,N_5027,N_5012);
nor U5575 (N_5575,N_5228,N_5397);
nor U5576 (N_5576,N_5067,N_5372);
xnor U5577 (N_5577,N_5392,N_5304);
or U5578 (N_5578,N_5235,N_5068);
nand U5579 (N_5579,N_5050,N_5163);
xnor U5580 (N_5580,N_5156,N_5076);
xnor U5581 (N_5581,N_5242,N_5057);
nand U5582 (N_5582,N_5105,N_5089);
nand U5583 (N_5583,N_5421,N_5476);
xnor U5584 (N_5584,N_5391,N_5299);
nand U5585 (N_5585,N_5395,N_5480);
nand U5586 (N_5586,N_5423,N_5041);
and U5587 (N_5587,N_5426,N_5042);
and U5588 (N_5588,N_5098,N_5394);
or U5589 (N_5589,N_5275,N_5205);
and U5590 (N_5590,N_5351,N_5090);
xor U5591 (N_5591,N_5263,N_5211);
nand U5592 (N_5592,N_5092,N_5073);
xor U5593 (N_5593,N_5297,N_5441);
xnor U5594 (N_5594,N_5387,N_5350);
nand U5595 (N_5595,N_5033,N_5472);
xor U5596 (N_5596,N_5286,N_5239);
xnor U5597 (N_5597,N_5378,N_5183);
nand U5598 (N_5598,N_5248,N_5380);
nand U5599 (N_5599,N_5364,N_5175);
xor U5600 (N_5600,N_5065,N_5347);
and U5601 (N_5601,N_5303,N_5341);
nor U5602 (N_5602,N_5417,N_5458);
or U5603 (N_5603,N_5340,N_5393);
xnor U5604 (N_5604,N_5128,N_5074);
nor U5605 (N_5605,N_5408,N_5434);
nor U5606 (N_5606,N_5373,N_5094);
and U5607 (N_5607,N_5139,N_5449);
xnor U5608 (N_5608,N_5184,N_5363);
and U5609 (N_5609,N_5466,N_5192);
or U5610 (N_5610,N_5142,N_5499);
xnor U5611 (N_5611,N_5199,N_5339);
nand U5612 (N_5612,N_5179,N_5291);
and U5613 (N_5613,N_5132,N_5287);
or U5614 (N_5614,N_5167,N_5136);
or U5615 (N_5615,N_5108,N_5138);
or U5616 (N_5616,N_5323,N_5087);
nor U5617 (N_5617,N_5356,N_5246);
nor U5618 (N_5618,N_5044,N_5104);
nand U5619 (N_5619,N_5324,N_5052);
nor U5620 (N_5620,N_5161,N_5405);
and U5621 (N_5621,N_5099,N_5025);
xnor U5622 (N_5622,N_5227,N_5134);
xor U5623 (N_5623,N_5464,N_5451);
xnor U5624 (N_5624,N_5298,N_5063);
nand U5625 (N_5625,N_5411,N_5450);
nor U5626 (N_5626,N_5215,N_5190);
and U5627 (N_5627,N_5439,N_5222);
and U5628 (N_5628,N_5117,N_5038);
or U5629 (N_5629,N_5308,N_5216);
and U5630 (N_5630,N_5479,N_5129);
xnor U5631 (N_5631,N_5030,N_5463);
nor U5632 (N_5632,N_5490,N_5440);
nand U5633 (N_5633,N_5317,N_5406);
and U5634 (N_5634,N_5316,N_5278);
xnor U5635 (N_5635,N_5428,N_5497);
nand U5636 (N_5636,N_5332,N_5185);
or U5637 (N_5637,N_5310,N_5150);
nand U5638 (N_5638,N_5255,N_5446);
nand U5639 (N_5639,N_5154,N_5168);
and U5640 (N_5640,N_5236,N_5045);
and U5641 (N_5641,N_5477,N_5195);
xnor U5642 (N_5642,N_5149,N_5334);
and U5643 (N_5643,N_5253,N_5212);
nand U5644 (N_5644,N_5327,N_5053);
and U5645 (N_5645,N_5164,N_5217);
nand U5646 (N_5646,N_5110,N_5171);
nand U5647 (N_5647,N_5039,N_5272);
or U5648 (N_5648,N_5188,N_5385);
or U5649 (N_5649,N_5344,N_5054);
nor U5650 (N_5650,N_5247,N_5486);
nand U5651 (N_5651,N_5133,N_5456);
or U5652 (N_5652,N_5243,N_5436);
nor U5653 (N_5653,N_5233,N_5198);
or U5654 (N_5654,N_5282,N_5468);
nand U5655 (N_5655,N_5230,N_5422);
nand U5656 (N_5656,N_5386,N_5093);
or U5657 (N_5657,N_5280,N_5488);
nor U5658 (N_5658,N_5146,N_5357);
and U5659 (N_5659,N_5444,N_5201);
nand U5660 (N_5660,N_5290,N_5346);
nand U5661 (N_5661,N_5021,N_5271);
nand U5662 (N_5662,N_5082,N_5013);
xor U5663 (N_5663,N_5288,N_5001);
xor U5664 (N_5664,N_5249,N_5333);
nand U5665 (N_5665,N_5197,N_5321);
xor U5666 (N_5666,N_5148,N_5210);
nor U5667 (N_5667,N_5338,N_5369);
xor U5668 (N_5668,N_5022,N_5106);
nor U5669 (N_5669,N_5379,N_5483);
xor U5670 (N_5670,N_5155,N_5051);
nand U5671 (N_5671,N_5008,N_5177);
nand U5672 (N_5672,N_5474,N_5281);
or U5673 (N_5673,N_5047,N_5302);
nor U5674 (N_5674,N_5234,N_5314);
or U5675 (N_5675,N_5187,N_5066);
or U5676 (N_5676,N_5125,N_5457);
nand U5677 (N_5677,N_5219,N_5024);
or U5678 (N_5678,N_5224,N_5452);
and U5679 (N_5679,N_5482,N_5313);
nand U5680 (N_5680,N_5354,N_5193);
nor U5681 (N_5681,N_5425,N_5186);
xnor U5682 (N_5682,N_5005,N_5412);
nand U5683 (N_5683,N_5305,N_5414);
xor U5684 (N_5684,N_5221,N_5088);
and U5685 (N_5685,N_5254,N_5361);
nand U5686 (N_5686,N_5433,N_5267);
nand U5687 (N_5687,N_5083,N_5475);
and U5688 (N_5688,N_5157,N_5189);
nor U5689 (N_5689,N_5174,N_5069);
and U5690 (N_5690,N_5009,N_5112);
or U5691 (N_5691,N_5116,N_5158);
and U5692 (N_5692,N_5260,N_5399);
and U5693 (N_5693,N_5176,N_5318);
nor U5694 (N_5694,N_5019,N_5382);
or U5695 (N_5695,N_5460,N_5495);
nor U5696 (N_5696,N_5229,N_5438);
nor U5697 (N_5697,N_5078,N_5359);
or U5698 (N_5698,N_5096,N_5265);
and U5699 (N_5699,N_5214,N_5086);
and U5700 (N_5700,N_5469,N_5437);
or U5701 (N_5701,N_5206,N_5160);
or U5702 (N_5702,N_5493,N_5470);
nand U5703 (N_5703,N_5204,N_5145);
nor U5704 (N_5704,N_5306,N_5141);
or U5705 (N_5705,N_5144,N_5353);
and U5706 (N_5706,N_5028,N_5345);
nor U5707 (N_5707,N_5420,N_5071);
nor U5708 (N_5708,N_5048,N_5130);
nand U5709 (N_5709,N_5319,N_5153);
and U5710 (N_5710,N_5258,N_5430);
or U5711 (N_5711,N_5352,N_5003);
xor U5712 (N_5712,N_5203,N_5276);
and U5713 (N_5713,N_5461,N_5342);
nand U5714 (N_5714,N_5401,N_5284);
or U5715 (N_5715,N_5181,N_5165);
xnor U5716 (N_5716,N_5331,N_5337);
xor U5717 (N_5717,N_5330,N_5348);
and U5718 (N_5718,N_5377,N_5018);
nor U5719 (N_5719,N_5349,N_5232);
and U5720 (N_5720,N_5238,N_5124);
or U5721 (N_5721,N_5427,N_5000);
nor U5722 (N_5722,N_5121,N_5257);
nand U5723 (N_5723,N_5459,N_5140);
nor U5724 (N_5724,N_5101,N_5072);
xor U5725 (N_5725,N_5173,N_5432);
xnor U5726 (N_5726,N_5295,N_5152);
or U5727 (N_5727,N_5429,N_5037);
and U5728 (N_5728,N_5085,N_5135);
and U5729 (N_5729,N_5300,N_5245);
and U5730 (N_5730,N_5122,N_5172);
nand U5731 (N_5731,N_5388,N_5240);
xor U5732 (N_5732,N_5031,N_5268);
or U5733 (N_5733,N_5285,N_5453);
or U5734 (N_5734,N_5431,N_5036);
xor U5735 (N_5735,N_5465,N_5103);
nand U5736 (N_5736,N_5237,N_5049);
or U5737 (N_5737,N_5084,N_5311);
or U5738 (N_5738,N_5208,N_5081);
or U5739 (N_5739,N_5435,N_5448);
nand U5740 (N_5740,N_5362,N_5404);
nand U5741 (N_5741,N_5301,N_5274);
and U5742 (N_5742,N_5114,N_5389);
nor U5743 (N_5743,N_5273,N_5381);
and U5744 (N_5744,N_5241,N_5478);
xnor U5745 (N_5745,N_5251,N_5119);
nor U5746 (N_5746,N_5370,N_5375);
nand U5747 (N_5747,N_5178,N_5120);
nor U5748 (N_5748,N_5403,N_5264);
and U5749 (N_5749,N_5147,N_5442);
or U5750 (N_5750,N_5076,N_5005);
nor U5751 (N_5751,N_5138,N_5404);
and U5752 (N_5752,N_5231,N_5208);
xnor U5753 (N_5753,N_5137,N_5136);
or U5754 (N_5754,N_5115,N_5327);
nand U5755 (N_5755,N_5443,N_5398);
or U5756 (N_5756,N_5238,N_5393);
or U5757 (N_5757,N_5160,N_5030);
and U5758 (N_5758,N_5198,N_5118);
and U5759 (N_5759,N_5322,N_5438);
and U5760 (N_5760,N_5075,N_5382);
xor U5761 (N_5761,N_5148,N_5281);
nand U5762 (N_5762,N_5075,N_5304);
or U5763 (N_5763,N_5475,N_5288);
nor U5764 (N_5764,N_5466,N_5226);
or U5765 (N_5765,N_5214,N_5113);
xor U5766 (N_5766,N_5187,N_5486);
nand U5767 (N_5767,N_5254,N_5283);
or U5768 (N_5768,N_5264,N_5119);
xor U5769 (N_5769,N_5100,N_5097);
nand U5770 (N_5770,N_5256,N_5229);
nor U5771 (N_5771,N_5168,N_5022);
xor U5772 (N_5772,N_5237,N_5166);
xnor U5773 (N_5773,N_5132,N_5196);
or U5774 (N_5774,N_5259,N_5180);
nor U5775 (N_5775,N_5142,N_5306);
nand U5776 (N_5776,N_5464,N_5366);
or U5777 (N_5777,N_5357,N_5168);
nor U5778 (N_5778,N_5033,N_5309);
or U5779 (N_5779,N_5477,N_5161);
nor U5780 (N_5780,N_5359,N_5353);
and U5781 (N_5781,N_5129,N_5203);
and U5782 (N_5782,N_5243,N_5160);
xnor U5783 (N_5783,N_5395,N_5063);
or U5784 (N_5784,N_5101,N_5416);
xor U5785 (N_5785,N_5186,N_5083);
xor U5786 (N_5786,N_5220,N_5399);
nand U5787 (N_5787,N_5196,N_5077);
and U5788 (N_5788,N_5157,N_5170);
and U5789 (N_5789,N_5350,N_5276);
xnor U5790 (N_5790,N_5471,N_5272);
xor U5791 (N_5791,N_5248,N_5041);
xnor U5792 (N_5792,N_5090,N_5254);
nand U5793 (N_5793,N_5200,N_5345);
xor U5794 (N_5794,N_5108,N_5152);
xnor U5795 (N_5795,N_5029,N_5169);
nand U5796 (N_5796,N_5326,N_5266);
nor U5797 (N_5797,N_5272,N_5187);
or U5798 (N_5798,N_5315,N_5092);
nor U5799 (N_5799,N_5009,N_5174);
nand U5800 (N_5800,N_5330,N_5409);
nor U5801 (N_5801,N_5230,N_5245);
or U5802 (N_5802,N_5445,N_5075);
or U5803 (N_5803,N_5177,N_5220);
nor U5804 (N_5804,N_5469,N_5179);
nand U5805 (N_5805,N_5023,N_5191);
nand U5806 (N_5806,N_5218,N_5046);
nor U5807 (N_5807,N_5151,N_5260);
nor U5808 (N_5808,N_5327,N_5021);
nor U5809 (N_5809,N_5456,N_5075);
or U5810 (N_5810,N_5238,N_5310);
and U5811 (N_5811,N_5167,N_5395);
nor U5812 (N_5812,N_5253,N_5122);
xnor U5813 (N_5813,N_5293,N_5353);
xnor U5814 (N_5814,N_5477,N_5319);
nand U5815 (N_5815,N_5164,N_5393);
xnor U5816 (N_5816,N_5453,N_5421);
xnor U5817 (N_5817,N_5214,N_5276);
xor U5818 (N_5818,N_5266,N_5468);
nor U5819 (N_5819,N_5068,N_5455);
nand U5820 (N_5820,N_5287,N_5463);
or U5821 (N_5821,N_5094,N_5236);
xnor U5822 (N_5822,N_5468,N_5013);
and U5823 (N_5823,N_5178,N_5252);
nand U5824 (N_5824,N_5169,N_5427);
and U5825 (N_5825,N_5376,N_5359);
or U5826 (N_5826,N_5343,N_5361);
xor U5827 (N_5827,N_5393,N_5008);
or U5828 (N_5828,N_5267,N_5125);
nand U5829 (N_5829,N_5311,N_5270);
and U5830 (N_5830,N_5386,N_5227);
nor U5831 (N_5831,N_5420,N_5132);
and U5832 (N_5832,N_5100,N_5340);
and U5833 (N_5833,N_5354,N_5148);
and U5834 (N_5834,N_5269,N_5337);
nand U5835 (N_5835,N_5323,N_5190);
xor U5836 (N_5836,N_5068,N_5093);
nand U5837 (N_5837,N_5029,N_5086);
nor U5838 (N_5838,N_5064,N_5361);
nor U5839 (N_5839,N_5490,N_5002);
xor U5840 (N_5840,N_5001,N_5396);
nor U5841 (N_5841,N_5455,N_5329);
or U5842 (N_5842,N_5023,N_5322);
xor U5843 (N_5843,N_5323,N_5271);
and U5844 (N_5844,N_5117,N_5317);
xor U5845 (N_5845,N_5180,N_5401);
nor U5846 (N_5846,N_5331,N_5399);
nor U5847 (N_5847,N_5253,N_5174);
nand U5848 (N_5848,N_5193,N_5078);
xnor U5849 (N_5849,N_5489,N_5210);
xnor U5850 (N_5850,N_5073,N_5046);
nor U5851 (N_5851,N_5255,N_5113);
xnor U5852 (N_5852,N_5278,N_5012);
nand U5853 (N_5853,N_5439,N_5308);
xor U5854 (N_5854,N_5102,N_5058);
nor U5855 (N_5855,N_5323,N_5380);
nor U5856 (N_5856,N_5212,N_5389);
or U5857 (N_5857,N_5485,N_5022);
xor U5858 (N_5858,N_5342,N_5031);
nor U5859 (N_5859,N_5049,N_5231);
nor U5860 (N_5860,N_5329,N_5109);
nor U5861 (N_5861,N_5356,N_5429);
and U5862 (N_5862,N_5192,N_5124);
or U5863 (N_5863,N_5155,N_5393);
xor U5864 (N_5864,N_5014,N_5039);
xor U5865 (N_5865,N_5373,N_5315);
nand U5866 (N_5866,N_5153,N_5364);
or U5867 (N_5867,N_5339,N_5203);
or U5868 (N_5868,N_5137,N_5243);
nor U5869 (N_5869,N_5458,N_5189);
nor U5870 (N_5870,N_5468,N_5070);
nor U5871 (N_5871,N_5114,N_5444);
xor U5872 (N_5872,N_5090,N_5330);
and U5873 (N_5873,N_5418,N_5156);
or U5874 (N_5874,N_5273,N_5290);
xor U5875 (N_5875,N_5067,N_5470);
nand U5876 (N_5876,N_5133,N_5174);
and U5877 (N_5877,N_5447,N_5337);
or U5878 (N_5878,N_5095,N_5411);
or U5879 (N_5879,N_5213,N_5063);
and U5880 (N_5880,N_5210,N_5453);
nor U5881 (N_5881,N_5214,N_5463);
nor U5882 (N_5882,N_5273,N_5392);
and U5883 (N_5883,N_5150,N_5477);
nor U5884 (N_5884,N_5122,N_5137);
and U5885 (N_5885,N_5258,N_5376);
xor U5886 (N_5886,N_5303,N_5238);
xor U5887 (N_5887,N_5317,N_5404);
or U5888 (N_5888,N_5308,N_5394);
or U5889 (N_5889,N_5325,N_5194);
xor U5890 (N_5890,N_5431,N_5240);
nor U5891 (N_5891,N_5039,N_5204);
xor U5892 (N_5892,N_5300,N_5054);
xor U5893 (N_5893,N_5037,N_5419);
nor U5894 (N_5894,N_5358,N_5469);
nand U5895 (N_5895,N_5483,N_5494);
nand U5896 (N_5896,N_5374,N_5170);
or U5897 (N_5897,N_5040,N_5495);
and U5898 (N_5898,N_5070,N_5240);
nand U5899 (N_5899,N_5094,N_5204);
or U5900 (N_5900,N_5299,N_5353);
nor U5901 (N_5901,N_5203,N_5385);
or U5902 (N_5902,N_5413,N_5458);
and U5903 (N_5903,N_5360,N_5475);
nand U5904 (N_5904,N_5234,N_5312);
nand U5905 (N_5905,N_5266,N_5144);
nor U5906 (N_5906,N_5197,N_5471);
and U5907 (N_5907,N_5457,N_5354);
or U5908 (N_5908,N_5325,N_5030);
and U5909 (N_5909,N_5216,N_5353);
xor U5910 (N_5910,N_5151,N_5345);
or U5911 (N_5911,N_5436,N_5226);
nor U5912 (N_5912,N_5174,N_5427);
nand U5913 (N_5913,N_5129,N_5277);
xnor U5914 (N_5914,N_5313,N_5377);
and U5915 (N_5915,N_5275,N_5078);
nor U5916 (N_5916,N_5463,N_5419);
nand U5917 (N_5917,N_5499,N_5144);
or U5918 (N_5918,N_5097,N_5099);
nor U5919 (N_5919,N_5014,N_5457);
nand U5920 (N_5920,N_5150,N_5300);
or U5921 (N_5921,N_5392,N_5197);
xor U5922 (N_5922,N_5078,N_5376);
or U5923 (N_5923,N_5320,N_5457);
and U5924 (N_5924,N_5391,N_5338);
xnor U5925 (N_5925,N_5458,N_5441);
nand U5926 (N_5926,N_5244,N_5190);
nor U5927 (N_5927,N_5481,N_5468);
nor U5928 (N_5928,N_5448,N_5412);
nor U5929 (N_5929,N_5352,N_5455);
or U5930 (N_5930,N_5053,N_5394);
nor U5931 (N_5931,N_5068,N_5053);
xnor U5932 (N_5932,N_5360,N_5427);
and U5933 (N_5933,N_5392,N_5443);
xor U5934 (N_5934,N_5323,N_5333);
nor U5935 (N_5935,N_5409,N_5212);
nand U5936 (N_5936,N_5360,N_5006);
and U5937 (N_5937,N_5407,N_5106);
xor U5938 (N_5938,N_5028,N_5440);
and U5939 (N_5939,N_5370,N_5140);
nor U5940 (N_5940,N_5441,N_5300);
and U5941 (N_5941,N_5127,N_5019);
or U5942 (N_5942,N_5295,N_5067);
or U5943 (N_5943,N_5190,N_5178);
nand U5944 (N_5944,N_5108,N_5250);
xor U5945 (N_5945,N_5362,N_5052);
nand U5946 (N_5946,N_5163,N_5305);
nor U5947 (N_5947,N_5161,N_5071);
or U5948 (N_5948,N_5101,N_5105);
nor U5949 (N_5949,N_5397,N_5412);
xnor U5950 (N_5950,N_5389,N_5323);
xnor U5951 (N_5951,N_5492,N_5132);
or U5952 (N_5952,N_5306,N_5117);
nand U5953 (N_5953,N_5135,N_5194);
nor U5954 (N_5954,N_5023,N_5117);
nor U5955 (N_5955,N_5374,N_5315);
nor U5956 (N_5956,N_5449,N_5329);
or U5957 (N_5957,N_5068,N_5107);
and U5958 (N_5958,N_5009,N_5158);
nand U5959 (N_5959,N_5001,N_5097);
and U5960 (N_5960,N_5021,N_5316);
or U5961 (N_5961,N_5021,N_5466);
nand U5962 (N_5962,N_5056,N_5223);
xor U5963 (N_5963,N_5052,N_5241);
or U5964 (N_5964,N_5353,N_5361);
nor U5965 (N_5965,N_5060,N_5101);
or U5966 (N_5966,N_5365,N_5122);
or U5967 (N_5967,N_5081,N_5425);
or U5968 (N_5968,N_5481,N_5436);
nor U5969 (N_5969,N_5188,N_5355);
nand U5970 (N_5970,N_5365,N_5007);
and U5971 (N_5971,N_5358,N_5308);
nor U5972 (N_5972,N_5499,N_5436);
nor U5973 (N_5973,N_5461,N_5180);
nand U5974 (N_5974,N_5357,N_5279);
nand U5975 (N_5975,N_5490,N_5191);
nand U5976 (N_5976,N_5464,N_5303);
or U5977 (N_5977,N_5002,N_5106);
nor U5978 (N_5978,N_5020,N_5480);
and U5979 (N_5979,N_5091,N_5258);
xnor U5980 (N_5980,N_5134,N_5354);
and U5981 (N_5981,N_5374,N_5091);
or U5982 (N_5982,N_5134,N_5148);
nand U5983 (N_5983,N_5250,N_5179);
nor U5984 (N_5984,N_5230,N_5049);
or U5985 (N_5985,N_5436,N_5199);
nor U5986 (N_5986,N_5259,N_5191);
and U5987 (N_5987,N_5316,N_5254);
or U5988 (N_5988,N_5131,N_5113);
xnor U5989 (N_5989,N_5328,N_5207);
nand U5990 (N_5990,N_5451,N_5237);
nor U5991 (N_5991,N_5238,N_5210);
and U5992 (N_5992,N_5101,N_5098);
or U5993 (N_5993,N_5477,N_5403);
nor U5994 (N_5994,N_5181,N_5259);
and U5995 (N_5995,N_5092,N_5211);
and U5996 (N_5996,N_5160,N_5048);
or U5997 (N_5997,N_5411,N_5099);
and U5998 (N_5998,N_5181,N_5376);
nand U5999 (N_5999,N_5277,N_5451);
or U6000 (N_6000,N_5690,N_5766);
nand U6001 (N_6001,N_5926,N_5789);
nor U6002 (N_6002,N_5527,N_5964);
or U6003 (N_6003,N_5618,N_5621);
nor U6004 (N_6004,N_5595,N_5764);
xnor U6005 (N_6005,N_5530,N_5542);
or U6006 (N_6006,N_5689,N_5614);
and U6007 (N_6007,N_5773,N_5893);
and U6008 (N_6008,N_5551,N_5899);
nand U6009 (N_6009,N_5914,N_5993);
nand U6010 (N_6010,N_5509,N_5747);
nor U6011 (N_6011,N_5655,N_5695);
xnor U6012 (N_6012,N_5841,N_5897);
xor U6013 (N_6013,N_5732,N_5617);
nor U6014 (N_6014,N_5792,N_5763);
and U6015 (N_6015,N_5734,N_5672);
nand U6016 (N_6016,N_5600,N_5541);
nor U6017 (N_6017,N_5913,N_5996);
xnor U6018 (N_6018,N_5526,N_5584);
or U6019 (N_6019,N_5995,N_5610);
and U6020 (N_6020,N_5649,N_5828);
and U6021 (N_6021,N_5639,N_5795);
nor U6022 (N_6022,N_5794,N_5592);
and U6023 (N_6023,N_5846,N_5825);
nand U6024 (N_6024,N_5706,N_5683);
or U6025 (N_6025,N_5814,N_5659);
and U6026 (N_6026,N_5619,N_5945);
and U6027 (N_6027,N_5924,N_5788);
nand U6028 (N_6028,N_5622,N_5571);
nor U6029 (N_6029,N_5790,N_5912);
or U6030 (N_6030,N_5705,N_5575);
and U6031 (N_6031,N_5546,N_5717);
nand U6032 (N_6032,N_5881,N_5851);
and U6033 (N_6033,N_5770,N_5955);
nand U6034 (N_6034,N_5835,N_5529);
nor U6035 (N_6035,N_5965,N_5975);
nor U6036 (N_6036,N_5808,N_5615);
xor U6037 (N_6037,N_5940,N_5858);
nand U6038 (N_6038,N_5632,N_5875);
or U6039 (N_6039,N_5710,N_5572);
or U6040 (N_6040,N_5979,N_5939);
nand U6041 (N_6041,N_5942,N_5888);
nand U6042 (N_6042,N_5654,N_5820);
nor U6043 (N_6043,N_5671,N_5512);
or U6044 (N_6044,N_5508,N_5601);
nor U6045 (N_6045,N_5757,N_5603);
nor U6046 (N_6046,N_5714,N_5643);
and U6047 (N_6047,N_5535,N_5531);
nand U6048 (N_6048,N_5980,N_5736);
nand U6049 (N_6049,N_5843,N_5831);
or U6050 (N_6050,N_5696,N_5554);
and U6051 (N_6051,N_5597,N_5755);
nand U6052 (N_6052,N_5577,N_5506);
nand U6053 (N_6053,N_5693,N_5974);
nand U6054 (N_6054,N_5886,N_5515);
and U6055 (N_6055,N_5839,N_5768);
nand U6056 (N_6056,N_5877,N_5910);
nor U6057 (N_6057,N_5564,N_5948);
nor U6058 (N_6058,N_5849,N_5907);
nand U6059 (N_6059,N_5803,N_5589);
or U6060 (N_6060,N_5813,N_5549);
nand U6061 (N_6061,N_5887,N_5548);
and U6062 (N_6062,N_5806,N_5981);
or U6063 (N_6063,N_5663,N_5898);
nor U6064 (N_6064,N_5868,N_5743);
nor U6065 (N_6065,N_5605,N_5517);
xor U6066 (N_6066,N_5532,N_5561);
or U6067 (N_6067,N_5552,N_5507);
xnor U6068 (N_6068,N_5657,N_5954);
and U6069 (N_6069,N_5999,N_5781);
nand U6070 (N_6070,N_5751,N_5812);
and U6071 (N_6071,N_5748,N_5973);
nand U6072 (N_6072,N_5982,N_5896);
nor U6073 (N_6073,N_5578,N_5834);
and U6074 (N_6074,N_5867,N_5593);
xor U6075 (N_6075,N_5890,N_5647);
or U6076 (N_6076,N_5819,N_5857);
nand U6077 (N_6077,N_5501,N_5780);
or U6078 (N_6078,N_5923,N_5536);
xor U6079 (N_6079,N_5811,N_5866);
or U6080 (N_6080,N_5873,N_5970);
or U6081 (N_6081,N_5938,N_5514);
nand U6082 (N_6082,N_5756,N_5627);
nor U6083 (N_6083,N_5556,N_5534);
or U6084 (N_6084,N_5775,N_5662);
or U6085 (N_6085,N_5692,N_5626);
or U6086 (N_6086,N_5528,N_5673);
xnor U6087 (N_6087,N_5901,N_5922);
nor U6088 (N_6088,N_5869,N_5956);
and U6089 (N_6089,N_5565,N_5590);
or U6090 (N_6090,N_5967,N_5720);
and U6091 (N_6091,N_5550,N_5563);
and U6092 (N_6092,N_5579,N_5772);
nor U6093 (N_6093,N_5917,N_5567);
nor U6094 (N_6094,N_5951,N_5933);
or U6095 (N_6095,N_5545,N_5539);
or U6096 (N_6096,N_5953,N_5596);
nor U6097 (N_6097,N_5521,N_5966);
or U6098 (N_6098,N_5997,N_5978);
nor U6099 (N_6099,N_5700,N_5816);
xnor U6100 (N_6100,N_5574,N_5651);
xor U6101 (N_6101,N_5568,N_5932);
xnor U6102 (N_6102,N_5730,N_5670);
nand U6103 (N_6103,N_5969,N_5776);
nor U6104 (N_6104,N_5909,N_5629);
or U6105 (N_6105,N_5698,N_5800);
or U6106 (N_6106,N_5959,N_5807);
and U6107 (N_6107,N_5809,N_5707);
nor U6108 (N_6108,N_5859,N_5599);
and U6109 (N_6109,N_5708,N_5797);
or U6110 (N_6110,N_5694,N_5667);
nor U6111 (N_6111,N_5968,N_5798);
or U6112 (N_6112,N_5726,N_5620);
nor U6113 (N_6113,N_5845,N_5885);
xnor U6114 (N_6114,N_5860,N_5746);
xor U6115 (N_6115,N_5523,N_5684);
xor U6116 (N_6116,N_5697,N_5669);
or U6117 (N_6117,N_5598,N_5837);
xor U6118 (N_6118,N_5738,N_5861);
nor U6119 (N_6119,N_5740,N_5796);
nand U6120 (N_6120,N_5986,N_5892);
and U6121 (N_6121,N_5958,N_5678);
nand U6122 (N_6122,N_5555,N_5761);
nor U6123 (N_6123,N_5716,N_5544);
or U6124 (N_6124,N_5641,N_5994);
and U6125 (N_6125,N_5637,N_5645);
xor U6126 (N_6126,N_5821,N_5674);
xnor U6127 (N_6127,N_5602,N_5502);
or U6128 (N_6128,N_5871,N_5636);
and U6129 (N_6129,N_5510,N_5949);
or U6130 (N_6130,N_5937,N_5947);
and U6131 (N_6131,N_5960,N_5739);
nor U6132 (N_6132,N_5988,N_5883);
nand U6133 (N_6133,N_5941,N_5902);
nand U6134 (N_6134,N_5850,N_5876);
nand U6135 (N_6135,N_5553,N_5786);
or U6136 (N_6136,N_5930,N_5987);
nor U6137 (N_6137,N_5744,N_5826);
xnor U6138 (N_6138,N_5658,N_5559);
nor U6139 (N_6139,N_5984,N_5934);
xor U6140 (N_6140,N_5864,N_5853);
or U6141 (N_6141,N_5504,N_5856);
nand U6142 (N_6142,N_5983,N_5870);
nor U6143 (N_6143,N_5903,N_5919);
nand U6144 (N_6144,N_5687,N_5525);
nor U6145 (N_6145,N_5633,N_5865);
nand U6146 (N_6146,N_5900,N_5946);
nand U6147 (N_6147,N_5961,N_5891);
xor U6148 (N_6148,N_5762,N_5712);
xnor U6149 (N_6149,N_5580,N_5591);
xnor U6150 (N_6150,N_5840,N_5962);
xnor U6151 (N_6151,N_5665,N_5588);
xor U6152 (N_6152,N_5827,N_5936);
and U6153 (N_6153,N_5918,N_5802);
xor U6154 (N_6154,N_5518,N_5688);
nor U6155 (N_6155,N_5822,N_5852);
and U6156 (N_6156,N_5884,N_5915);
nor U6157 (N_6157,N_5774,N_5569);
nor U6158 (N_6158,N_5990,N_5685);
and U6159 (N_6159,N_5573,N_5950);
nand U6160 (N_6160,N_5963,N_5511);
xor U6161 (N_6161,N_5681,N_5906);
nor U6162 (N_6162,N_5842,N_5503);
nor U6163 (N_6163,N_5652,N_5725);
or U6164 (N_6164,N_5759,N_5661);
nor U6165 (N_6165,N_5566,N_5880);
xnor U6166 (N_6166,N_5735,N_5711);
xor U6167 (N_6167,N_5513,N_5741);
xor U6168 (N_6168,N_5624,N_5824);
nor U6169 (N_6169,N_5522,N_5646);
or U6170 (N_6170,N_5991,N_5943);
nand U6171 (N_6171,N_5771,N_5728);
nor U6172 (N_6172,N_5648,N_5718);
nor U6173 (N_6173,N_5823,N_5872);
or U6174 (N_6174,N_5804,N_5976);
nand U6175 (N_6175,N_5699,N_5628);
and U6176 (N_6176,N_5754,N_5829);
or U6177 (N_6177,N_5971,N_5640);
or U6178 (N_6178,N_5791,N_5724);
nand U6179 (N_6179,N_5838,N_5989);
or U6180 (N_6180,N_5611,N_5935);
nor U6181 (N_6181,N_5516,N_5682);
nand U6182 (N_6182,N_5815,N_5832);
nand U6183 (N_6183,N_5650,N_5562);
nor U6184 (N_6184,N_5863,N_5929);
or U6185 (N_6185,N_5889,N_5855);
and U6186 (N_6186,N_5904,N_5928);
nand U6187 (N_6187,N_5558,N_5547);
nand U6188 (N_6188,N_5778,N_5810);
and U6189 (N_6189,N_5606,N_5878);
nor U6190 (N_6190,N_5644,N_5931);
and U6191 (N_6191,N_5540,N_5957);
and U6192 (N_6192,N_5557,N_5782);
nor U6193 (N_6193,N_5769,N_5666);
nand U6194 (N_6194,N_5801,N_5701);
xnor U6195 (N_6195,N_5836,N_5727);
and U6196 (N_6196,N_5642,N_5664);
nor U6197 (N_6197,N_5713,N_5653);
or U6198 (N_6198,N_5607,N_5721);
and U6199 (N_6199,N_5952,N_5911);
or U6200 (N_6200,N_5719,N_5635);
nor U6201 (N_6201,N_5533,N_5679);
xor U6202 (N_6202,N_5758,N_5920);
nor U6203 (N_6203,N_5818,N_5704);
and U6204 (N_6204,N_5998,N_5874);
nor U6205 (N_6205,N_5765,N_5630);
nand U6206 (N_6206,N_5703,N_5927);
and U6207 (N_6207,N_5777,N_5753);
nor U6208 (N_6208,N_5537,N_5972);
or U6209 (N_6209,N_5745,N_5844);
xnor U6210 (N_6210,N_5742,N_5582);
and U6211 (N_6211,N_5731,N_5767);
xor U6212 (N_6212,N_5604,N_5894);
xnor U6213 (N_6213,N_5752,N_5660);
nand U6214 (N_6214,N_5560,N_5785);
nand U6215 (N_6215,N_5702,N_5519);
xor U6216 (N_6216,N_5905,N_5847);
nand U6217 (N_6217,N_5992,N_5680);
xor U6218 (N_6218,N_5505,N_5848);
or U6219 (N_6219,N_5921,N_5908);
nand U6220 (N_6220,N_5784,N_5805);
xor U6221 (N_6221,N_5676,N_5691);
nand U6222 (N_6222,N_5587,N_5722);
nand U6223 (N_6223,N_5817,N_5686);
or U6224 (N_6224,N_5916,N_5882);
nor U6225 (N_6225,N_5586,N_5608);
nor U6226 (N_6226,N_5862,N_5977);
or U6227 (N_6227,N_5609,N_5830);
nand U6228 (N_6228,N_5985,N_5500);
nor U6229 (N_6229,N_5616,N_5638);
xnor U6230 (N_6230,N_5799,N_5594);
nand U6231 (N_6231,N_5723,N_5656);
or U6232 (N_6232,N_5709,N_5668);
nor U6233 (N_6233,N_5520,N_5925);
or U6234 (N_6234,N_5625,N_5750);
xnor U6235 (N_6235,N_5715,N_5895);
and U6236 (N_6236,N_5634,N_5787);
and U6237 (N_6237,N_5675,N_5733);
xnor U6238 (N_6238,N_5729,N_5879);
xor U6239 (N_6239,N_5631,N_5783);
xnor U6240 (N_6240,N_5944,N_5538);
xor U6241 (N_6241,N_5623,N_5576);
nor U6242 (N_6242,N_5677,N_5749);
nor U6243 (N_6243,N_5833,N_5524);
xor U6244 (N_6244,N_5570,N_5583);
nor U6245 (N_6245,N_5543,N_5585);
and U6246 (N_6246,N_5737,N_5612);
xnor U6247 (N_6247,N_5581,N_5760);
nand U6248 (N_6248,N_5779,N_5793);
nand U6249 (N_6249,N_5613,N_5854);
or U6250 (N_6250,N_5795,N_5785);
nand U6251 (N_6251,N_5701,N_5604);
xor U6252 (N_6252,N_5972,N_5745);
nor U6253 (N_6253,N_5925,N_5694);
xnor U6254 (N_6254,N_5716,N_5930);
or U6255 (N_6255,N_5909,N_5641);
xor U6256 (N_6256,N_5778,N_5578);
nor U6257 (N_6257,N_5651,N_5972);
or U6258 (N_6258,N_5622,N_5896);
xor U6259 (N_6259,N_5875,N_5572);
or U6260 (N_6260,N_5597,N_5998);
or U6261 (N_6261,N_5778,N_5621);
or U6262 (N_6262,N_5748,N_5913);
nand U6263 (N_6263,N_5973,N_5658);
and U6264 (N_6264,N_5744,N_5963);
nor U6265 (N_6265,N_5725,N_5755);
nor U6266 (N_6266,N_5717,N_5923);
xnor U6267 (N_6267,N_5812,N_5620);
nor U6268 (N_6268,N_5915,N_5924);
and U6269 (N_6269,N_5998,N_5611);
and U6270 (N_6270,N_5554,N_5789);
xor U6271 (N_6271,N_5722,N_5721);
nand U6272 (N_6272,N_5700,N_5969);
xnor U6273 (N_6273,N_5715,N_5729);
or U6274 (N_6274,N_5824,N_5612);
or U6275 (N_6275,N_5969,N_5637);
nor U6276 (N_6276,N_5629,N_5973);
nor U6277 (N_6277,N_5932,N_5756);
nand U6278 (N_6278,N_5636,N_5576);
xnor U6279 (N_6279,N_5636,N_5501);
nor U6280 (N_6280,N_5991,N_5599);
nor U6281 (N_6281,N_5855,N_5831);
nor U6282 (N_6282,N_5827,N_5863);
nand U6283 (N_6283,N_5865,N_5882);
xnor U6284 (N_6284,N_5652,N_5924);
and U6285 (N_6285,N_5706,N_5863);
or U6286 (N_6286,N_5944,N_5523);
or U6287 (N_6287,N_5672,N_5510);
nor U6288 (N_6288,N_5699,N_5576);
or U6289 (N_6289,N_5813,N_5898);
nor U6290 (N_6290,N_5522,N_5573);
and U6291 (N_6291,N_5971,N_5955);
xnor U6292 (N_6292,N_5976,N_5532);
nor U6293 (N_6293,N_5654,N_5925);
and U6294 (N_6294,N_5938,N_5955);
xor U6295 (N_6295,N_5661,N_5629);
and U6296 (N_6296,N_5640,N_5683);
and U6297 (N_6297,N_5995,N_5991);
nor U6298 (N_6298,N_5955,N_5904);
and U6299 (N_6299,N_5977,N_5903);
or U6300 (N_6300,N_5859,N_5754);
or U6301 (N_6301,N_5954,N_5601);
nor U6302 (N_6302,N_5912,N_5781);
or U6303 (N_6303,N_5791,N_5992);
or U6304 (N_6304,N_5593,N_5909);
or U6305 (N_6305,N_5617,N_5738);
xnor U6306 (N_6306,N_5977,N_5609);
nor U6307 (N_6307,N_5700,N_5542);
and U6308 (N_6308,N_5907,N_5605);
and U6309 (N_6309,N_5646,N_5881);
nand U6310 (N_6310,N_5876,N_5838);
and U6311 (N_6311,N_5503,N_5735);
or U6312 (N_6312,N_5853,N_5867);
or U6313 (N_6313,N_5661,N_5951);
or U6314 (N_6314,N_5840,N_5934);
and U6315 (N_6315,N_5564,N_5653);
nor U6316 (N_6316,N_5558,N_5548);
nand U6317 (N_6317,N_5687,N_5539);
and U6318 (N_6318,N_5791,N_5668);
nor U6319 (N_6319,N_5592,N_5654);
and U6320 (N_6320,N_5897,N_5544);
nor U6321 (N_6321,N_5714,N_5953);
nor U6322 (N_6322,N_5969,N_5952);
nand U6323 (N_6323,N_5544,N_5677);
and U6324 (N_6324,N_5568,N_5750);
and U6325 (N_6325,N_5517,N_5803);
nand U6326 (N_6326,N_5562,N_5826);
and U6327 (N_6327,N_5767,N_5738);
nor U6328 (N_6328,N_5579,N_5605);
nand U6329 (N_6329,N_5999,N_5876);
xnor U6330 (N_6330,N_5540,N_5601);
and U6331 (N_6331,N_5863,N_5503);
nand U6332 (N_6332,N_5956,N_5523);
nor U6333 (N_6333,N_5566,N_5638);
xor U6334 (N_6334,N_5962,N_5889);
or U6335 (N_6335,N_5901,N_5672);
and U6336 (N_6336,N_5759,N_5566);
xor U6337 (N_6337,N_5831,N_5750);
nand U6338 (N_6338,N_5752,N_5760);
nand U6339 (N_6339,N_5510,N_5779);
or U6340 (N_6340,N_5862,N_5715);
and U6341 (N_6341,N_5638,N_5619);
nor U6342 (N_6342,N_5669,N_5504);
or U6343 (N_6343,N_5673,N_5743);
and U6344 (N_6344,N_5731,N_5777);
nor U6345 (N_6345,N_5918,N_5528);
nor U6346 (N_6346,N_5932,N_5722);
nand U6347 (N_6347,N_5697,N_5535);
xnor U6348 (N_6348,N_5517,N_5919);
nand U6349 (N_6349,N_5549,N_5994);
nand U6350 (N_6350,N_5805,N_5819);
and U6351 (N_6351,N_5699,N_5849);
nor U6352 (N_6352,N_5588,N_5666);
nor U6353 (N_6353,N_5603,N_5787);
nand U6354 (N_6354,N_5816,N_5508);
nand U6355 (N_6355,N_5552,N_5832);
nor U6356 (N_6356,N_5718,N_5734);
or U6357 (N_6357,N_5916,N_5936);
and U6358 (N_6358,N_5963,N_5998);
and U6359 (N_6359,N_5852,N_5783);
nor U6360 (N_6360,N_5739,N_5803);
nand U6361 (N_6361,N_5571,N_5866);
and U6362 (N_6362,N_5951,N_5919);
xnor U6363 (N_6363,N_5979,N_5695);
or U6364 (N_6364,N_5814,N_5729);
or U6365 (N_6365,N_5628,N_5550);
nor U6366 (N_6366,N_5778,N_5582);
nand U6367 (N_6367,N_5613,N_5583);
xor U6368 (N_6368,N_5901,N_5607);
nand U6369 (N_6369,N_5796,N_5567);
xnor U6370 (N_6370,N_5817,N_5552);
nand U6371 (N_6371,N_5528,N_5845);
nor U6372 (N_6372,N_5820,N_5677);
or U6373 (N_6373,N_5618,N_5739);
xnor U6374 (N_6374,N_5504,N_5960);
or U6375 (N_6375,N_5912,N_5989);
or U6376 (N_6376,N_5995,N_5882);
xor U6377 (N_6377,N_5722,N_5501);
nor U6378 (N_6378,N_5720,N_5961);
nand U6379 (N_6379,N_5824,N_5631);
nor U6380 (N_6380,N_5697,N_5753);
xor U6381 (N_6381,N_5510,N_5581);
xnor U6382 (N_6382,N_5554,N_5674);
and U6383 (N_6383,N_5540,N_5652);
nand U6384 (N_6384,N_5996,N_5915);
and U6385 (N_6385,N_5908,N_5806);
and U6386 (N_6386,N_5969,N_5953);
or U6387 (N_6387,N_5577,N_5984);
nor U6388 (N_6388,N_5680,N_5930);
or U6389 (N_6389,N_5833,N_5543);
xnor U6390 (N_6390,N_5753,N_5960);
nor U6391 (N_6391,N_5678,N_5671);
xnor U6392 (N_6392,N_5660,N_5772);
or U6393 (N_6393,N_5686,N_5842);
and U6394 (N_6394,N_5764,N_5643);
or U6395 (N_6395,N_5570,N_5861);
xor U6396 (N_6396,N_5787,N_5624);
and U6397 (N_6397,N_5664,N_5837);
xnor U6398 (N_6398,N_5993,N_5843);
nand U6399 (N_6399,N_5810,N_5989);
xnor U6400 (N_6400,N_5659,N_5888);
or U6401 (N_6401,N_5632,N_5759);
xor U6402 (N_6402,N_5937,N_5849);
and U6403 (N_6403,N_5841,N_5524);
nor U6404 (N_6404,N_5975,N_5585);
nand U6405 (N_6405,N_5921,N_5822);
xnor U6406 (N_6406,N_5814,N_5534);
nand U6407 (N_6407,N_5600,N_5656);
or U6408 (N_6408,N_5690,N_5618);
nand U6409 (N_6409,N_5719,N_5921);
nand U6410 (N_6410,N_5900,N_5732);
nand U6411 (N_6411,N_5751,N_5647);
nor U6412 (N_6412,N_5836,N_5774);
or U6413 (N_6413,N_5749,N_5581);
nor U6414 (N_6414,N_5697,N_5916);
nand U6415 (N_6415,N_5597,N_5712);
nor U6416 (N_6416,N_5714,N_5505);
and U6417 (N_6417,N_5898,N_5900);
nand U6418 (N_6418,N_5795,N_5659);
and U6419 (N_6419,N_5891,N_5719);
or U6420 (N_6420,N_5990,N_5590);
or U6421 (N_6421,N_5974,N_5743);
nor U6422 (N_6422,N_5522,N_5615);
or U6423 (N_6423,N_5715,N_5694);
or U6424 (N_6424,N_5587,N_5550);
xnor U6425 (N_6425,N_5620,N_5966);
nand U6426 (N_6426,N_5959,N_5896);
nand U6427 (N_6427,N_5638,N_5726);
or U6428 (N_6428,N_5835,N_5594);
xnor U6429 (N_6429,N_5565,N_5504);
nand U6430 (N_6430,N_5564,N_5889);
or U6431 (N_6431,N_5790,N_5953);
and U6432 (N_6432,N_5570,N_5824);
xor U6433 (N_6433,N_5712,N_5973);
or U6434 (N_6434,N_5918,N_5743);
xor U6435 (N_6435,N_5537,N_5545);
or U6436 (N_6436,N_5927,N_5525);
and U6437 (N_6437,N_5553,N_5577);
nor U6438 (N_6438,N_5513,N_5691);
or U6439 (N_6439,N_5587,N_5833);
nand U6440 (N_6440,N_5674,N_5880);
nor U6441 (N_6441,N_5982,N_5837);
xor U6442 (N_6442,N_5598,N_5725);
and U6443 (N_6443,N_5809,N_5683);
nor U6444 (N_6444,N_5833,N_5966);
nor U6445 (N_6445,N_5536,N_5826);
or U6446 (N_6446,N_5627,N_5892);
nand U6447 (N_6447,N_5866,N_5981);
nor U6448 (N_6448,N_5893,N_5671);
xnor U6449 (N_6449,N_5604,N_5583);
or U6450 (N_6450,N_5555,N_5992);
and U6451 (N_6451,N_5825,N_5827);
or U6452 (N_6452,N_5716,N_5714);
xnor U6453 (N_6453,N_5689,N_5912);
and U6454 (N_6454,N_5776,N_5961);
or U6455 (N_6455,N_5969,N_5866);
or U6456 (N_6456,N_5665,N_5981);
xnor U6457 (N_6457,N_5874,N_5948);
xor U6458 (N_6458,N_5826,N_5801);
or U6459 (N_6459,N_5827,N_5549);
xor U6460 (N_6460,N_5711,N_5726);
xnor U6461 (N_6461,N_5919,N_5924);
and U6462 (N_6462,N_5619,N_5887);
and U6463 (N_6463,N_5542,N_5789);
and U6464 (N_6464,N_5706,N_5881);
xnor U6465 (N_6465,N_5786,N_5703);
nand U6466 (N_6466,N_5830,N_5869);
or U6467 (N_6467,N_5531,N_5802);
nand U6468 (N_6468,N_5662,N_5711);
or U6469 (N_6469,N_5890,N_5661);
and U6470 (N_6470,N_5809,N_5697);
nand U6471 (N_6471,N_5638,N_5998);
nor U6472 (N_6472,N_5624,N_5527);
nand U6473 (N_6473,N_5633,N_5882);
nor U6474 (N_6474,N_5676,N_5646);
nor U6475 (N_6475,N_5729,N_5665);
or U6476 (N_6476,N_5999,N_5977);
and U6477 (N_6477,N_5827,N_5996);
nor U6478 (N_6478,N_5762,N_5941);
or U6479 (N_6479,N_5971,N_5699);
or U6480 (N_6480,N_5686,N_5800);
nand U6481 (N_6481,N_5892,N_5898);
nand U6482 (N_6482,N_5580,N_5990);
and U6483 (N_6483,N_5952,N_5899);
or U6484 (N_6484,N_5871,N_5867);
or U6485 (N_6485,N_5822,N_5939);
xnor U6486 (N_6486,N_5897,N_5904);
and U6487 (N_6487,N_5784,N_5760);
nand U6488 (N_6488,N_5807,N_5802);
xnor U6489 (N_6489,N_5850,N_5553);
and U6490 (N_6490,N_5722,N_5677);
and U6491 (N_6491,N_5923,N_5640);
xor U6492 (N_6492,N_5550,N_5707);
and U6493 (N_6493,N_5679,N_5901);
and U6494 (N_6494,N_5881,N_5886);
nor U6495 (N_6495,N_5812,N_5529);
or U6496 (N_6496,N_5813,N_5625);
xor U6497 (N_6497,N_5541,N_5864);
xor U6498 (N_6498,N_5561,N_5509);
and U6499 (N_6499,N_5597,N_5719);
xor U6500 (N_6500,N_6349,N_6466);
xor U6501 (N_6501,N_6153,N_6264);
or U6502 (N_6502,N_6363,N_6198);
and U6503 (N_6503,N_6078,N_6445);
and U6504 (N_6504,N_6008,N_6042);
xor U6505 (N_6505,N_6353,N_6339);
nand U6506 (N_6506,N_6218,N_6086);
and U6507 (N_6507,N_6321,N_6407);
nand U6508 (N_6508,N_6205,N_6290);
and U6509 (N_6509,N_6098,N_6019);
xnor U6510 (N_6510,N_6118,N_6117);
and U6511 (N_6511,N_6389,N_6040);
and U6512 (N_6512,N_6240,N_6108);
and U6513 (N_6513,N_6248,N_6041);
and U6514 (N_6514,N_6159,N_6379);
nor U6515 (N_6515,N_6322,N_6007);
and U6516 (N_6516,N_6273,N_6369);
or U6517 (N_6517,N_6103,N_6491);
nor U6518 (N_6518,N_6224,N_6386);
xor U6519 (N_6519,N_6021,N_6374);
or U6520 (N_6520,N_6012,N_6392);
or U6521 (N_6521,N_6282,N_6469);
xor U6522 (N_6522,N_6383,N_6373);
and U6523 (N_6523,N_6320,N_6256);
or U6524 (N_6524,N_6497,N_6064);
nand U6525 (N_6525,N_6483,N_6201);
or U6526 (N_6526,N_6430,N_6289);
nand U6527 (N_6527,N_6160,N_6452);
or U6528 (N_6528,N_6357,N_6366);
and U6529 (N_6529,N_6095,N_6423);
xnor U6530 (N_6530,N_6332,N_6310);
and U6531 (N_6531,N_6154,N_6152);
nand U6532 (N_6532,N_6482,N_6355);
xor U6533 (N_6533,N_6395,N_6192);
nand U6534 (N_6534,N_6415,N_6306);
nand U6535 (N_6535,N_6125,N_6486);
or U6536 (N_6536,N_6167,N_6227);
xnor U6537 (N_6537,N_6171,N_6314);
and U6538 (N_6538,N_6024,N_6146);
xnor U6539 (N_6539,N_6058,N_6250);
or U6540 (N_6540,N_6473,N_6069);
nor U6541 (N_6541,N_6197,N_6189);
nor U6542 (N_6542,N_6283,N_6063);
or U6543 (N_6543,N_6061,N_6252);
nor U6544 (N_6544,N_6259,N_6182);
and U6545 (N_6545,N_6105,N_6422);
and U6546 (N_6546,N_6472,N_6009);
or U6547 (N_6547,N_6246,N_6362);
or U6548 (N_6548,N_6443,N_6387);
xnor U6549 (N_6549,N_6420,N_6335);
and U6550 (N_6550,N_6367,N_6066);
xor U6551 (N_6551,N_6408,N_6276);
or U6552 (N_6552,N_6270,N_6225);
nand U6553 (N_6553,N_6128,N_6275);
xor U6554 (N_6554,N_6032,N_6404);
xnor U6555 (N_6555,N_6333,N_6114);
or U6556 (N_6556,N_6203,N_6476);
xnor U6557 (N_6557,N_6255,N_6072);
and U6558 (N_6558,N_6375,N_6399);
xnor U6559 (N_6559,N_6220,N_6079);
nand U6560 (N_6560,N_6313,N_6204);
or U6561 (N_6561,N_6456,N_6281);
xnor U6562 (N_6562,N_6429,N_6342);
xor U6563 (N_6563,N_6223,N_6149);
or U6564 (N_6564,N_6142,N_6150);
nand U6565 (N_6565,N_6331,N_6348);
or U6566 (N_6566,N_6442,N_6434);
or U6567 (N_6567,N_6265,N_6002);
nor U6568 (N_6568,N_6376,N_6168);
nand U6569 (N_6569,N_6318,N_6060);
xor U6570 (N_6570,N_6351,N_6485);
nand U6571 (N_6571,N_6065,N_6188);
or U6572 (N_6572,N_6499,N_6120);
nand U6573 (N_6573,N_6412,N_6101);
nand U6574 (N_6574,N_6488,N_6481);
or U6575 (N_6575,N_6294,N_6479);
nand U6576 (N_6576,N_6228,N_6083);
xnor U6577 (N_6577,N_6451,N_6341);
nor U6578 (N_6578,N_6176,N_6001);
nand U6579 (N_6579,N_6358,N_6444);
and U6580 (N_6580,N_6003,N_6496);
nor U6581 (N_6581,N_6277,N_6365);
and U6582 (N_6582,N_6409,N_6028);
nor U6583 (N_6583,N_6298,N_6226);
nand U6584 (N_6584,N_6133,N_6196);
or U6585 (N_6585,N_6242,N_6311);
xnor U6586 (N_6586,N_6081,N_6401);
or U6587 (N_6587,N_6241,N_6454);
nor U6588 (N_6588,N_6006,N_6174);
nand U6589 (N_6589,N_6300,N_6193);
and U6590 (N_6590,N_6080,N_6088);
or U6591 (N_6591,N_6402,N_6087);
or U6592 (N_6592,N_6170,N_6030);
nand U6593 (N_6593,N_6183,N_6364);
and U6594 (N_6594,N_6140,N_6119);
or U6595 (N_6595,N_6112,N_6372);
or U6596 (N_6596,N_6207,N_6417);
or U6597 (N_6597,N_6157,N_6286);
xor U6598 (N_6598,N_6144,N_6410);
nor U6599 (N_6599,N_6102,N_6347);
nand U6600 (N_6600,N_6037,N_6050);
xor U6601 (N_6601,N_6371,N_6464);
and U6602 (N_6602,N_6292,N_6460);
xor U6603 (N_6603,N_6453,N_6474);
or U6604 (N_6604,N_6352,N_6465);
and U6605 (N_6605,N_6129,N_6151);
xnor U6606 (N_6606,N_6293,N_6010);
and U6607 (N_6607,N_6084,N_6155);
and U6608 (N_6608,N_6187,N_6051);
and U6609 (N_6609,N_6428,N_6141);
or U6610 (N_6610,N_6044,N_6249);
and U6611 (N_6611,N_6418,N_6437);
nand U6612 (N_6612,N_6446,N_6082);
nand U6613 (N_6613,N_6092,N_6390);
and U6614 (N_6614,N_6109,N_6014);
and U6615 (N_6615,N_6459,N_6016);
nor U6616 (N_6616,N_6023,N_6394);
and U6617 (N_6617,N_6291,N_6457);
nor U6618 (N_6618,N_6097,N_6219);
nand U6619 (N_6619,N_6115,N_6340);
or U6620 (N_6620,N_6400,N_6123);
and U6621 (N_6621,N_6035,N_6278);
nor U6622 (N_6622,N_6162,N_6234);
xor U6623 (N_6623,N_6380,N_6495);
nor U6624 (N_6624,N_6186,N_6492);
nand U6625 (N_6625,N_6271,N_6135);
nand U6626 (N_6626,N_6238,N_6093);
xor U6627 (N_6627,N_6489,N_6048);
or U6628 (N_6628,N_6326,N_6266);
xnor U6629 (N_6629,N_6074,N_6243);
and U6630 (N_6630,N_6161,N_6011);
nor U6631 (N_6631,N_6107,N_6047);
or U6632 (N_6632,N_6480,N_6137);
and U6633 (N_6633,N_6308,N_6164);
or U6634 (N_6634,N_6431,N_6261);
nand U6635 (N_6635,N_6257,N_6034);
nand U6636 (N_6636,N_6020,N_6113);
or U6637 (N_6637,N_6136,N_6462);
nand U6638 (N_6638,N_6054,N_6253);
xor U6639 (N_6639,N_6381,N_6438);
nor U6640 (N_6640,N_6181,N_6163);
xnor U6641 (N_6641,N_6124,N_6104);
or U6642 (N_6642,N_6022,N_6175);
nand U6643 (N_6643,N_6370,N_6406);
nor U6644 (N_6644,N_6089,N_6467);
nor U6645 (N_6645,N_6450,N_6449);
xor U6646 (N_6646,N_6268,N_6377);
xor U6647 (N_6647,N_6049,N_6411);
nand U6648 (N_6648,N_6075,N_6031);
xor U6649 (N_6649,N_6191,N_6235);
xor U6650 (N_6650,N_6000,N_6303);
nand U6651 (N_6651,N_6209,N_6468);
nor U6652 (N_6652,N_6360,N_6165);
nand U6653 (N_6653,N_6071,N_6039);
nor U6654 (N_6654,N_6070,N_6206);
xnor U6655 (N_6655,N_6356,N_6315);
nor U6656 (N_6656,N_6309,N_6384);
nand U6657 (N_6657,N_6396,N_6319);
or U6658 (N_6658,N_6324,N_6148);
or U6659 (N_6659,N_6327,N_6296);
or U6660 (N_6660,N_6287,N_6251);
or U6661 (N_6661,N_6062,N_6116);
and U6662 (N_6662,N_6328,N_6388);
nand U6663 (N_6663,N_6233,N_6130);
or U6664 (N_6664,N_6121,N_6194);
or U6665 (N_6665,N_6132,N_6447);
or U6666 (N_6666,N_6173,N_6214);
or U6667 (N_6667,N_6413,N_6004);
and U6668 (N_6668,N_6269,N_6245);
and U6669 (N_6669,N_6435,N_6279);
nand U6670 (N_6670,N_6230,N_6427);
nor U6671 (N_6671,N_6096,N_6138);
nor U6672 (N_6672,N_6337,N_6237);
and U6673 (N_6673,N_6302,N_6222);
xor U6674 (N_6674,N_6439,N_6131);
or U6675 (N_6675,N_6398,N_6036);
or U6676 (N_6676,N_6359,N_6471);
or U6677 (N_6677,N_6441,N_6263);
nand U6678 (N_6678,N_6229,N_6301);
nand U6679 (N_6679,N_6448,N_6025);
nor U6680 (N_6680,N_6297,N_6247);
xnor U6681 (N_6681,N_6166,N_6426);
and U6682 (N_6682,N_6493,N_6232);
nor U6683 (N_6683,N_6258,N_6052);
nor U6684 (N_6684,N_6385,N_6091);
nand U6685 (N_6685,N_6077,N_6026);
xor U6686 (N_6686,N_6272,N_6433);
nor U6687 (N_6687,N_6334,N_6178);
and U6688 (N_6688,N_6099,N_6033);
or U6689 (N_6689,N_6354,N_6346);
xor U6690 (N_6690,N_6043,N_6414);
nand U6691 (N_6691,N_6260,N_6147);
nor U6692 (N_6692,N_6216,N_6285);
or U6693 (N_6693,N_6158,N_6419);
nor U6694 (N_6694,N_6038,N_6210);
nor U6695 (N_6695,N_6425,N_6323);
and U6696 (N_6696,N_6169,N_6076);
xnor U6697 (N_6697,N_6073,N_6344);
xnor U6698 (N_6698,N_6202,N_6350);
nand U6699 (N_6699,N_6127,N_6382);
xnor U6700 (N_6700,N_6484,N_6057);
and U6701 (N_6701,N_6288,N_6477);
or U6702 (N_6702,N_6100,N_6325);
nor U6703 (N_6703,N_6046,N_6305);
nor U6704 (N_6704,N_6316,N_6126);
nor U6705 (N_6705,N_6304,N_6068);
nand U6706 (N_6706,N_6461,N_6329);
xor U6707 (N_6707,N_6424,N_6343);
xnor U6708 (N_6708,N_6199,N_6027);
or U6709 (N_6709,N_6338,N_6221);
nor U6710 (N_6710,N_6094,N_6180);
or U6711 (N_6711,N_6184,N_6254);
and U6712 (N_6712,N_6336,N_6330);
nor U6713 (N_6713,N_6017,N_6111);
or U6714 (N_6714,N_6211,N_6045);
nor U6715 (N_6715,N_6085,N_6059);
nor U6716 (N_6716,N_6200,N_6274);
or U6717 (N_6717,N_6280,N_6156);
and U6718 (N_6718,N_6185,N_6056);
nand U6719 (N_6719,N_6478,N_6029);
and U6720 (N_6720,N_6317,N_6244);
nand U6721 (N_6721,N_6145,N_6440);
and U6722 (N_6722,N_6498,N_6416);
xor U6723 (N_6723,N_6110,N_6455);
nand U6724 (N_6724,N_6463,N_6134);
or U6725 (N_6725,N_6018,N_6231);
or U6726 (N_6726,N_6378,N_6458);
xnor U6727 (N_6727,N_6393,N_6307);
nand U6728 (N_6728,N_6179,N_6208);
nand U6729 (N_6729,N_6421,N_6312);
nand U6730 (N_6730,N_6470,N_6195);
or U6731 (N_6731,N_6172,N_6236);
nand U6732 (N_6732,N_6190,N_6436);
and U6733 (N_6733,N_6475,N_6177);
xnor U6734 (N_6734,N_6299,N_6405);
nand U6735 (N_6735,N_6432,N_6215);
or U6736 (N_6736,N_6403,N_6494);
nand U6737 (N_6737,N_6361,N_6212);
and U6738 (N_6738,N_6295,N_6345);
nor U6739 (N_6739,N_6139,N_6055);
xnor U6740 (N_6740,N_6067,N_6122);
nor U6741 (N_6741,N_6397,N_6013);
nand U6742 (N_6742,N_6143,N_6267);
or U6743 (N_6743,N_6284,N_6391);
and U6744 (N_6744,N_6490,N_6106);
or U6745 (N_6745,N_6487,N_6368);
nor U6746 (N_6746,N_6015,N_6090);
nor U6747 (N_6747,N_6217,N_6005);
nand U6748 (N_6748,N_6053,N_6262);
nor U6749 (N_6749,N_6213,N_6239);
and U6750 (N_6750,N_6169,N_6135);
or U6751 (N_6751,N_6208,N_6298);
and U6752 (N_6752,N_6012,N_6124);
and U6753 (N_6753,N_6020,N_6431);
nor U6754 (N_6754,N_6193,N_6093);
nand U6755 (N_6755,N_6472,N_6375);
nor U6756 (N_6756,N_6237,N_6301);
or U6757 (N_6757,N_6033,N_6479);
or U6758 (N_6758,N_6209,N_6273);
nor U6759 (N_6759,N_6216,N_6450);
xor U6760 (N_6760,N_6197,N_6460);
nor U6761 (N_6761,N_6142,N_6157);
nor U6762 (N_6762,N_6305,N_6281);
nor U6763 (N_6763,N_6262,N_6114);
and U6764 (N_6764,N_6375,N_6208);
or U6765 (N_6765,N_6035,N_6130);
or U6766 (N_6766,N_6087,N_6489);
and U6767 (N_6767,N_6429,N_6020);
nand U6768 (N_6768,N_6183,N_6421);
xnor U6769 (N_6769,N_6027,N_6035);
xor U6770 (N_6770,N_6017,N_6296);
nor U6771 (N_6771,N_6325,N_6299);
xor U6772 (N_6772,N_6019,N_6252);
and U6773 (N_6773,N_6286,N_6324);
xnor U6774 (N_6774,N_6477,N_6082);
xor U6775 (N_6775,N_6157,N_6124);
xor U6776 (N_6776,N_6499,N_6436);
and U6777 (N_6777,N_6423,N_6422);
nor U6778 (N_6778,N_6126,N_6425);
nor U6779 (N_6779,N_6227,N_6269);
nor U6780 (N_6780,N_6226,N_6075);
or U6781 (N_6781,N_6427,N_6387);
and U6782 (N_6782,N_6261,N_6380);
xor U6783 (N_6783,N_6415,N_6237);
or U6784 (N_6784,N_6226,N_6208);
or U6785 (N_6785,N_6103,N_6406);
xnor U6786 (N_6786,N_6401,N_6179);
xor U6787 (N_6787,N_6376,N_6179);
nand U6788 (N_6788,N_6228,N_6363);
or U6789 (N_6789,N_6386,N_6230);
or U6790 (N_6790,N_6126,N_6170);
or U6791 (N_6791,N_6438,N_6056);
or U6792 (N_6792,N_6431,N_6184);
and U6793 (N_6793,N_6046,N_6158);
nor U6794 (N_6794,N_6244,N_6465);
or U6795 (N_6795,N_6130,N_6121);
xnor U6796 (N_6796,N_6006,N_6285);
nor U6797 (N_6797,N_6395,N_6466);
or U6798 (N_6798,N_6092,N_6123);
and U6799 (N_6799,N_6202,N_6323);
or U6800 (N_6800,N_6484,N_6355);
and U6801 (N_6801,N_6340,N_6483);
or U6802 (N_6802,N_6190,N_6438);
nand U6803 (N_6803,N_6485,N_6059);
xor U6804 (N_6804,N_6152,N_6465);
nor U6805 (N_6805,N_6094,N_6071);
nand U6806 (N_6806,N_6331,N_6192);
nor U6807 (N_6807,N_6446,N_6119);
xor U6808 (N_6808,N_6128,N_6166);
or U6809 (N_6809,N_6421,N_6484);
or U6810 (N_6810,N_6077,N_6305);
xor U6811 (N_6811,N_6319,N_6371);
nand U6812 (N_6812,N_6027,N_6073);
xor U6813 (N_6813,N_6095,N_6093);
and U6814 (N_6814,N_6115,N_6017);
and U6815 (N_6815,N_6391,N_6277);
and U6816 (N_6816,N_6443,N_6141);
and U6817 (N_6817,N_6256,N_6378);
xor U6818 (N_6818,N_6238,N_6295);
nor U6819 (N_6819,N_6107,N_6006);
and U6820 (N_6820,N_6152,N_6187);
nor U6821 (N_6821,N_6476,N_6262);
xnor U6822 (N_6822,N_6041,N_6485);
or U6823 (N_6823,N_6386,N_6344);
xor U6824 (N_6824,N_6094,N_6372);
or U6825 (N_6825,N_6484,N_6414);
xor U6826 (N_6826,N_6099,N_6111);
nand U6827 (N_6827,N_6437,N_6261);
or U6828 (N_6828,N_6089,N_6057);
nor U6829 (N_6829,N_6183,N_6315);
xor U6830 (N_6830,N_6495,N_6232);
nand U6831 (N_6831,N_6181,N_6351);
nand U6832 (N_6832,N_6107,N_6395);
and U6833 (N_6833,N_6368,N_6211);
nand U6834 (N_6834,N_6304,N_6498);
nand U6835 (N_6835,N_6483,N_6404);
xor U6836 (N_6836,N_6285,N_6206);
xnor U6837 (N_6837,N_6177,N_6146);
nand U6838 (N_6838,N_6436,N_6456);
or U6839 (N_6839,N_6016,N_6197);
nor U6840 (N_6840,N_6063,N_6045);
or U6841 (N_6841,N_6343,N_6274);
or U6842 (N_6842,N_6263,N_6390);
xor U6843 (N_6843,N_6484,N_6192);
or U6844 (N_6844,N_6237,N_6391);
nor U6845 (N_6845,N_6454,N_6410);
nand U6846 (N_6846,N_6174,N_6368);
or U6847 (N_6847,N_6402,N_6436);
nand U6848 (N_6848,N_6229,N_6340);
nand U6849 (N_6849,N_6466,N_6025);
and U6850 (N_6850,N_6271,N_6161);
or U6851 (N_6851,N_6081,N_6432);
nand U6852 (N_6852,N_6065,N_6338);
nand U6853 (N_6853,N_6440,N_6233);
and U6854 (N_6854,N_6108,N_6470);
or U6855 (N_6855,N_6273,N_6491);
nand U6856 (N_6856,N_6338,N_6088);
and U6857 (N_6857,N_6011,N_6466);
nand U6858 (N_6858,N_6193,N_6103);
and U6859 (N_6859,N_6045,N_6259);
or U6860 (N_6860,N_6208,N_6103);
or U6861 (N_6861,N_6059,N_6077);
nor U6862 (N_6862,N_6069,N_6154);
nor U6863 (N_6863,N_6135,N_6150);
xnor U6864 (N_6864,N_6264,N_6353);
nor U6865 (N_6865,N_6411,N_6024);
nand U6866 (N_6866,N_6193,N_6395);
xor U6867 (N_6867,N_6100,N_6203);
nor U6868 (N_6868,N_6410,N_6391);
xor U6869 (N_6869,N_6008,N_6228);
xnor U6870 (N_6870,N_6039,N_6076);
nand U6871 (N_6871,N_6214,N_6467);
and U6872 (N_6872,N_6398,N_6497);
xnor U6873 (N_6873,N_6076,N_6206);
xor U6874 (N_6874,N_6105,N_6294);
nor U6875 (N_6875,N_6010,N_6154);
nand U6876 (N_6876,N_6429,N_6150);
or U6877 (N_6877,N_6039,N_6041);
and U6878 (N_6878,N_6290,N_6249);
nand U6879 (N_6879,N_6168,N_6081);
and U6880 (N_6880,N_6472,N_6314);
and U6881 (N_6881,N_6472,N_6499);
xnor U6882 (N_6882,N_6148,N_6039);
xor U6883 (N_6883,N_6099,N_6055);
nand U6884 (N_6884,N_6080,N_6049);
xnor U6885 (N_6885,N_6397,N_6066);
and U6886 (N_6886,N_6272,N_6414);
nand U6887 (N_6887,N_6105,N_6394);
nor U6888 (N_6888,N_6132,N_6103);
and U6889 (N_6889,N_6322,N_6166);
or U6890 (N_6890,N_6077,N_6067);
or U6891 (N_6891,N_6086,N_6365);
and U6892 (N_6892,N_6397,N_6473);
nor U6893 (N_6893,N_6321,N_6492);
and U6894 (N_6894,N_6011,N_6396);
nand U6895 (N_6895,N_6154,N_6267);
nor U6896 (N_6896,N_6134,N_6026);
nor U6897 (N_6897,N_6425,N_6161);
nor U6898 (N_6898,N_6014,N_6212);
nand U6899 (N_6899,N_6084,N_6391);
nor U6900 (N_6900,N_6230,N_6498);
and U6901 (N_6901,N_6472,N_6240);
or U6902 (N_6902,N_6081,N_6270);
and U6903 (N_6903,N_6172,N_6040);
nor U6904 (N_6904,N_6083,N_6324);
or U6905 (N_6905,N_6318,N_6250);
and U6906 (N_6906,N_6093,N_6023);
nor U6907 (N_6907,N_6108,N_6485);
and U6908 (N_6908,N_6143,N_6013);
nor U6909 (N_6909,N_6257,N_6322);
nor U6910 (N_6910,N_6452,N_6270);
or U6911 (N_6911,N_6072,N_6308);
nor U6912 (N_6912,N_6375,N_6231);
xnor U6913 (N_6913,N_6003,N_6065);
xor U6914 (N_6914,N_6269,N_6063);
nand U6915 (N_6915,N_6288,N_6033);
xor U6916 (N_6916,N_6103,N_6497);
nor U6917 (N_6917,N_6434,N_6026);
or U6918 (N_6918,N_6021,N_6236);
nand U6919 (N_6919,N_6471,N_6397);
or U6920 (N_6920,N_6354,N_6389);
xor U6921 (N_6921,N_6158,N_6359);
xnor U6922 (N_6922,N_6181,N_6221);
nor U6923 (N_6923,N_6476,N_6113);
or U6924 (N_6924,N_6023,N_6063);
nor U6925 (N_6925,N_6162,N_6258);
and U6926 (N_6926,N_6295,N_6050);
and U6927 (N_6927,N_6060,N_6471);
xor U6928 (N_6928,N_6102,N_6324);
and U6929 (N_6929,N_6056,N_6370);
nand U6930 (N_6930,N_6184,N_6093);
nor U6931 (N_6931,N_6149,N_6249);
xor U6932 (N_6932,N_6313,N_6008);
nand U6933 (N_6933,N_6075,N_6024);
and U6934 (N_6934,N_6173,N_6369);
or U6935 (N_6935,N_6300,N_6002);
or U6936 (N_6936,N_6455,N_6434);
or U6937 (N_6937,N_6021,N_6250);
nand U6938 (N_6938,N_6255,N_6049);
nor U6939 (N_6939,N_6153,N_6198);
nor U6940 (N_6940,N_6153,N_6341);
xnor U6941 (N_6941,N_6095,N_6292);
nand U6942 (N_6942,N_6317,N_6125);
xnor U6943 (N_6943,N_6422,N_6171);
nand U6944 (N_6944,N_6122,N_6222);
and U6945 (N_6945,N_6214,N_6065);
and U6946 (N_6946,N_6243,N_6294);
xor U6947 (N_6947,N_6497,N_6104);
or U6948 (N_6948,N_6120,N_6067);
xnor U6949 (N_6949,N_6107,N_6263);
nand U6950 (N_6950,N_6084,N_6072);
xor U6951 (N_6951,N_6475,N_6169);
or U6952 (N_6952,N_6268,N_6009);
nand U6953 (N_6953,N_6175,N_6032);
or U6954 (N_6954,N_6134,N_6129);
nand U6955 (N_6955,N_6384,N_6159);
nand U6956 (N_6956,N_6279,N_6485);
nand U6957 (N_6957,N_6025,N_6255);
nor U6958 (N_6958,N_6096,N_6141);
nor U6959 (N_6959,N_6304,N_6181);
or U6960 (N_6960,N_6178,N_6312);
nand U6961 (N_6961,N_6433,N_6327);
or U6962 (N_6962,N_6145,N_6466);
or U6963 (N_6963,N_6041,N_6286);
xnor U6964 (N_6964,N_6166,N_6360);
nand U6965 (N_6965,N_6335,N_6090);
nor U6966 (N_6966,N_6337,N_6145);
and U6967 (N_6967,N_6365,N_6456);
nand U6968 (N_6968,N_6064,N_6065);
and U6969 (N_6969,N_6222,N_6497);
and U6970 (N_6970,N_6439,N_6323);
xor U6971 (N_6971,N_6122,N_6339);
or U6972 (N_6972,N_6380,N_6351);
nand U6973 (N_6973,N_6283,N_6166);
nor U6974 (N_6974,N_6029,N_6292);
or U6975 (N_6975,N_6427,N_6022);
and U6976 (N_6976,N_6131,N_6435);
or U6977 (N_6977,N_6221,N_6189);
and U6978 (N_6978,N_6431,N_6178);
and U6979 (N_6979,N_6102,N_6068);
xor U6980 (N_6980,N_6475,N_6126);
nor U6981 (N_6981,N_6362,N_6012);
nor U6982 (N_6982,N_6200,N_6146);
nor U6983 (N_6983,N_6201,N_6308);
nor U6984 (N_6984,N_6443,N_6213);
xnor U6985 (N_6985,N_6232,N_6412);
or U6986 (N_6986,N_6344,N_6051);
xor U6987 (N_6987,N_6102,N_6375);
xor U6988 (N_6988,N_6428,N_6412);
xnor U6989 (N_6989,N_6144,N_6380);
nor U6990 (N_6990,N_6138,N_6348);
and U6991 (N_6991,N_6371,N_6021);
xor U6992 (N_6992,N_6093,N_6341);
and U6993 (N_6993,N_6173,N_6223);
nand U6994 (N_6994,N_6468,N_6234);
and U6995 (N_6995,N_6192,N_6054);
xor U6996 (N_6996,N_6008,N_6167);
xnor U6997 (N_6997,N_6393,N_6423);
or U6998 (N_6998,N_6160,N_6457);
and U6999 (N_6999,N_6072,N_6298);
and U7000 (N_7000,N_6891,N_6707);
xor U7001 (N_7001,N_6742,N_6817);
nand U7002 (N_7002,N_6961,N_6989);
nand U7003 (N_7003,N_6938,N_6716);
xnor U7004 (N_7004,N_6741,N_6559);
nand U7005 (N_7005,N_6619,N_6608);
nand U7006 (N_7006,N_6708,N_6797);
or U7007 (N_7007,N_6591,N_6852);
nor U7008 (N_7008,N_6954,N_6916);
xnor U7009 (N_7009,N_6884,N_6600);
nand U7010 (N_7010,N_6779,N_6509);
and U7011 (N_7011,N_6581,N_6740);
or U7012 (N_7012,N_6935,N_6712);
and U7013 (N_7013,N_6860,N_6547);
nand U7014 (N_7014,N_6930,N_6504);
nor U7015 (N_7015,N_6668,N_6861);
nand U7016 (N_7016,N_6620,N_6722);
nand U7017 (N_7017,N_6728,N_6832);
xor U7018 (N_7018,N_6531,N_6900);
or U7019 (N_7019,N_6637,N_6751);
nand U7020 (N_7020,N_6758,N_6720);
and U7021 (N_7021,N_6967,N_6725);
xor U7022 (N_7022,N_6950,N_6840);
nor U7023 (N_7023,N_6634,N_6786);
and U7024 (N_7024,N_6656,N_6703);
or U7025 (N_7025,N_6543,N_6812);
and U7026 (N_7026,N_6567,N_6622);
xnor U7027 (N_7027,N_6664,N_6841);
nand U7028 (N_7028,N_6881,N_6635);
nor U7029 (N_7029,N_6548,N_6919);
nand U7030 (N_7030,N_6941,N_6612);
nand U7031 (N_7031,N_6533,N_6507);
or U7032 (N_7032,N_6746,N_6765);
nand U7033 (N_7033,N_6909,N_6944);
nor U7034 (N_7034,N_6711,N_6523);
nor U7035 (N_7035,N_6987,N_6848);
or U7036 (N_7036,N_6966,N_6690);
nand U7037 (N_7037,N_6697,N_6870);
xnor U7038 (N_7038,N_6988,N_6671);
xnor U7039 (N_7039,N_6638,N_6649);
nand U7040 (N_7040,N_6997,N_6945);
and U7041 (N_7041,N_6560,N_6578);
and U7042 (N_7042,N_6563,N_6974);
xor U7043 (N_7043,N_6971,N_6685);
nand U7044 (N_7044,N_6538,N_6680);
or U7045 (N_7045,N_6541,N_6570);
nor U7046 (N_7046,N_6962,N_6788);
nor U7047 (N_7047,N_6611,N_6598);
xnor U7048 (N_7048,N_6862,N_6748);
nor U7049 (N_7049,N_6757,N_6926);
and U7050 (N_7050,N_6929,N_6546);
or U7051 (N_7051,N_6763,N_6502);
xor U7052 (N_7052,N_6630,N_6605);
and U7053 (N_7053,N_6624,N_6903);
xor U7054 (N_7054,N_6667,N_6921);
nor U7055 (N_7055,N_6760,N_6535);
nor U7056 (N_7056,N_6991,N_6554);
nor U7057 (N_7057,N_6659,N_6985);
and U7058 (N_7058,N_6984,N_6647);
nand U7059 (N_7059,N_6837,N_6815);
xnor U7060 (N_7060,N_6947,N_6830);
nor U7061 (N_7061,N_6596,N_6931);
or U7062 (N_7062,N_6510,N_6617);
or U7063 (N_7063,N_6769,N_6787);
nor U7064 (N_7064,N_6995,N_6529);
and U7065 (N_7065,N_6770,N_6828);
or U7066 (N_7066,N_6928,N_6863);
xnor U7067 (N_7067,N_6642,N_6799);
nand U7068 (N_7068,N_6876,N_6654);
xnor U7069 (N_7069,N_6552,N_6964);
nor U7070 (N_7070,N_6963,N_6606);
or U7071 (N_7071,N_6628,N_6917);
nand U7072 (N_7072,N_6899,N_6705);
nor U7073 (N_7073,N_6805,N_6820);
nor U7074 (N_7074,N_6717,N_6942);
nor U7075 (N_7075,N_6882,N_6579);
or U7076 (N_7076,N_6896,N_6990);
and U7077 (N_7077,N_6802,N_6776);
nand U7078 (N_7078,N_6975,N_6885);
xor U7079 (N_7079,N_6993,N_6747);
or U7080 (N_7080,N_6678,N_6616);
or U7081 (N_7081,N_6661,N_6652);
and U7082 (N_7082,N_6924,N_6726);
or U7083 (N_7083,N_6994,N_6681);
xnor U7084 (N_7084,N_6835,N_6925);
nand U7085 (N_7085,N_6922,N_6519);
nor U7086 (N_7086,N_6851,N_6674);
nor U7087 (N_7087,N_6969,N_6810);
nand U7088 (N_7088,N_6599,N_6887);
or U7089 (N_7089,N_6819,N_6526);
xnor U7090 (N_7090,N_6764,N_6693);
and U7091 (N_7091,N_6845,N_6901);
nor U7092 (N_7092,N_6595,N_6713);
xnor U7093 (N_7093,N_6827,N_6958);
nand U7094 (N_7094,N_6610,N_6539);
nor U7095 (N_7095,N_6673,N_6582);
xnor U7096 (N_7096,N_6934,N_6773);
nor U7097 (N_7097,N_6853,N_6576);
and U7098 (N_7098,N_6771,N_6683);
xor U7099 (N_7099,N_6515,N_6601);
or U7100 (N_7100,N_6687,N_6551);
nand U7101 (N_7101,N_6530,N_6524);
nor U7102 (N_7102,N_6977,N_6998);
xnor U7103 (N_7103,N_6505,N_6886);
nor U7104 (N_7104,N_6645,N_6556);
nor U7105 (N_7105,N_6633,N_6575);
nor U7106 (N_7106,N_6960,N_6933);
nor U7107 (N_7107,N_6749,N_6709);
and U7108 (N_7108,N_6537,N_6972);
and U7109 (N_7109,N_6590,N_6508);
xor U7110 (N_7110,N_6566,N_6883);
nor U7111 (N_7111,N_6544,N_6952);
xor U7112 (N_7112,N_6604,N_6937);
nand U7113 (N_7113,N_6892,N_6676);
nand U7114 (N_7114,N_6784,N_6532);
nand U7115 (N_7115,N_6593,N_6842);
and U7116 (N_7116,N_6948,N_6516);
nor U7117 (N_7117,N_6754,N_6890);
nand U7118 (N_7118,N_6906,N_6733);
nand U7119 (N_7119,N_6923,N_6744);
and U7120 (N_7120,N_6545,N_6694);
and U7121 (N_7121,N_6677,N_6872);
nor U7122 (N_7122,N_6918,N_6970);
nor U7123 (N_7123,N_6996,N_6889);
or U7124 (N_7124,N_6855,N_6833);
xor U7125 (N_7125,N_6636,N_6957);
and U7126 (N_7126,N_6914,N_6809);
xor U7127 (N_7127,N_6528,N_6500);
nand U7128 (N_7128,N_6755,N_6761);
or U7129 (N_7129,N_6806,N_6506);
xnor U7130 (N_7130,N_6540,N_6793);
and U7131 (N_7131,N_6573,N_6568);
nor U7132 (N_7132,N_6874,N_6829);
nand U7133 (N_7133,N_6609,N_6669);
and U7134 (N_7134,N_6702,N_6873);
and U7135 (N_7135,N_6586,N_6785);
and U7136 (N_7136,N_6580,N_6911);
and U7137 (N_7137,N_6557,N_6627);
xor U7138 (N_7138,N_6825,N_6721);
or U7139 (N_7139,N_6912,N_6574);
xnor U7140 (N_7140,N_6865,N_6864);
and U7141 (N_7141,N_6814,N_6572);
or U7142 (N_7142,N_6613,N_6655);
nand U7143 (N_7143,N_6589,N_6796);
or U7144 (N_7144,N_6897,N_6959);
nor U7145 (N_7145,N_6893,N_6846);
nor U7146 (N_7146,N_6880,N_6867);
and U7147 (N_7147,N_6587,N_6768);
or U7148 (N_7148,N_6672,N_6780);
and U7149 (N_7149,N_6907,N_6710);
xnor U7150 (N_7150,N_6759,N_6550);
nand U7151 (N_7151,N_6953,N_6525);
nor U7152 (N_7152,N_6940,N_6982);
nand U7153 (N_7153,N_6735,N_6908);
or U7154 (N_7154,N_6781,N_6653);
nand U7155 (N_7155,N_6752,N_6879);
or U7156 (N_7156,N_6571,N_6729);
or U7157 (N_7157,N_6976,N_6804);
and U7158 (N_7158,N_6738,N_6650);
or U7159 (N_7159,N_6795,N_6807);
and U7160 (N_7160,N_6902,N_6691);
and U7161 (N_7161,N_6818,N_6737);
nor U7162 (N_7162,N_6730,N_6555);
nor U7163 (N_7163,N_6866,N_6648);
and U7164 (N_7164,N_6943,N_6670);
nor U7165 (N_7165,N_6665,N_6868);
or U7166 (N_7166,N_6727,N_6803);
nand U7167 (N_7167,N_6986,N_6715);
nand U7168 (N_7168,N_6839,N_6679);
nor U7169 (N_7169,N_6932,N_6520);
and U7170 (N_7170,N_6626,N_6513);
or U7171 (N_7171,N_6856,N_6564);
and U7172 (N_7172,N_6767,N_6615);
and U7173 (N_7173,N_6542,N_6847);
and U7174 (N_7174,N_6849,N_6791);
nand U7175 (N_7175,N_6501,N_6859);
nand U7176 (N_7176,N_6704,N_6724);
nand U7177 (N_7177,N_6714,N_6651);
nand U7178 (N_7178,N_6898,N_6894);
nand U7179 (N_7179,N_6983,N_6871);
xnor U7180 (N_7180,N_6913,N_6992);
nand U7181 (N_7181,N_6745,N_6657);
or U7182 (N_7182,N_6646,N_6583);
nand U7183 (N_7183,N_6844,N_6731);
nor U7184 (N_7184,N_6965,N_6723);
nor U7185 (N_7185,N_6831,N_6904);
or U7186 (N_7186,N_6558,N_6739);
nor U7187 (N_7187,N_6927,N_6663);
nor U7188 (N_7188,N_6823,N_6623);
or U7189 (N_7189,N_6675,N_6521);
xnor U7190 (N_7190,N_6905,N_6701);
or U7191 (N_7191,N_6684,N_6632);
xnor U7192 (N_7192,N_6843,N_6792);
and U7193 (N_7193,N_6565,N_6584);
nor U7194 (N_7194,N_6621,N_6920);
or U7195 (N_7195,N_6698,N_6949);
nand U7196 (N_7196,N_6790,N_6618);
nor U7197 (N_7197,N_6813,N_6699);
and U7198 (N_7198,N_6700,N_6696);
and U7199 (N_7199,N_6801,N_6999);
and U7200 (N_7200,N_6614,N_6869);
or U7201 (N_7201,N_6895,N_6689);
nand U7202 (N_7202,N_6798,N_6512);
nand U7203 (N_7203,N_6732,N_6518);
nor U7204 (N_7204,N_6822,N_6762);
xnor U7205 (N_7205,N_6602,N_6658);
and U7206 (N_7206,N_6756,N_6750);
and U7207 (N_7207,N_6625,N_6640);
nand U7208 (N_7208,N_6816,N_6777);
nand U7209 (N_7209,N_6607,N_6527);
and U7210 (N_7210,N_6808,N_6838);
and U7211 (N_7211,N_6666,N_6955);
or U7212 (N_7212,N_6973,N_6603);
or U7213 (N_7213,N_6718,N_6644);
nor U7214 (N_7214,N_6800,N_6695);
nor U7215 (N_7215,N_6743,N_6719);
or U7216 (N_7216,N_6734,N_6878);
nand U7217 (N_7217,N_6766,N_6774);
xor U7218 (N_7218,N_6688,N_6951);
nor U7219 (N_7219,N_6794,N_6824);
nand U7220 (N_7220,N_6854,N_6811);
xnor U7221 (N_7221,N_6778,N_6789);
and U7222 (N_7222,N_6775,N_6753);
xor U7223 (N_7223,N_6597,N_6834);
xor U7224 (N_7224,N_6826,N_6686);
and U7225 (N_7225,N_6660,N_6850);
or U7226 (N_7226,N_6875,N_6858);
nand U7227 (N_7227,N_6631,N_6821);
xnor U7228 (N_7228,N_6978,N_6956);
nor U7229 (N_7229,N_6888,N_6592);
nand U7230 (N_7230,N_6594,N_6772);
and U7231 (N_7231,N_6561,N_6736);
nand U7232 (N_7232,N_6836,N_6936);
nand U7233 (N_7233,N_6980,N_6629);
xor U7234 (N_7234,N_6643,N_6511);
nand U7235 (N_7235,N_6522,N_6585);
and U7236 (N_7236,N_6562,N_6692);
and U7237 (N_7237,N_6536,N_6857);
nand U7238 (N_7238,N_6534,N_6939);
and U7239 (N_7239,N_6782,N_6639);
nor U7240 (N_7240,N_6783,N_6514);
xnor U7241 (N_7241,N_6588,N_6662);
and U7242 (N_7242,N_6569,N_6910);
or U7243 (N_7243,N_6979,N_6981);
nor U7244 (N_7244,N_6641,N_6577);
nor U7245 (N_7245,N_6549,N_6553);
and U7246 (N_7246,N_6706,N_6946);
nor U7247 (N_7247,N_6968,N_6915);
xnor U7248 (N_7248,N_6682,N_6503);
or U7249 (N_7249,N_6877,N_6517);
or U7250 (N_7250,N_6533,N_6724);
xnor U7251 (N_7251,N_6748,N_6939);
nor U7252 (N_7252,N_6894,N_6515);
and U7253 (N_7253,N_6707,N_6777);
or U7254 (N_7254,N_6673,N_6523);
nor U7255 (N_7255,N_6576,N_6705);
and U7256 (N_7256,N_6920,N_6827);
nand U7257 (N_7257,N_6596,N_6939);
and U7258 (N_7258,N_6849,N_6718);
nor U7259 (N_7259,N_6860,N_6514);
nand U7260 (N_7260,N_6513,N_6543);
and U7261 (N_7261,N_6791,N_6709);
nor U7262 (N_7262,N_6699,N_6871);
nand U7263 (N_7263,N_6966,N_6994);
and U7264 (N_7264,N_6801,N_6571);
nor U7265 (N_7265,N_6661,N_6881);
nor U7266 (N_7266,N_6611,N_6575);
or U7267 (N_7267,N_6939,N_6862);
nor U7268 (N_7268,N_6842,N_6749);
nand U7269 (N_7269,N_6734,N_6566);
or U7270 (N_7270,N_6849,N_6892);
and U7271 (N_7271,N_6781,N_6675);
or U7272 (N_7272,N_6641,N_6527);
nand U7273 (N_7273,N_6897,N_6863);
nor U7274 (N_7274,N_6685,N_6599);
xnor U7275 (N_7275,N_6599,N_6915);
nand U7276 (N_7276,N_6528,N_6723);
nor U7277 (N_7277,N_6870,N_6782);
nand U7278 (N_7278,N_6850,N_6902);
nand U7279 (N_7279,N_6513,N_6768);
and U7280 (N_7280,N_6970,N_6618);
and U7281 (N_7281,N_6850,N_6508);
or U7282 (N_7282,N_6533,N_6677);
nor U7283 (N_7283,N_6565,N_6882);
or U7284 (N_7284,N_6993,N_6806);
or U7285 (N_7285,N_6789,N_6841);
and U7286 (N_7286,N_6623,N_6951);
and U7287 (N_7287,N_6577,N_6684);
and U7288 (N_7288,N_6980,N_6982);
or U7289 (N_7289,N_6823,N_6896);
and U7290 (N_7290,N_6841,N_6532);
or U7291 (N_7291,N_6794,N_6695);
nor U7292 (N_7292,N_6824,N_6609);
xnor U7293 (N_7293,N_6671,N_6919);
xor U7294 (N_7294,N_6679,N_6584);
and U7295 (N_7295,N_6543,N_6762);
and U7296 (N_7296,N_6598,N_6657);
nor U7297 (N_7297,N_6906,N_6601);
nor U7298 (N_7298,N_6737,N_6642);
nor U7299 (N_7299,N_6622,N_6558);
xor U7300 (N_7300,N_6972,N_6717);
or U7301 (N_7301,N_6932,N_6845);
nand U7302 (N_7302,N_6974,N_6763);
nand U7303 (N_7303,N_6573,N_6566);
nor U7304 (N_7304,N_6647,N_6717);
nand U7305 (N_7305,N_6705,N_6546);
xor U7306 (N_7306,N_6944,N_6923);
nor U7307 (N_7307,N_6858,N_6840);
and U7308 (N_7308,N_6740,N_6922);
xnor U7309 (N_7309,N_6990,N_6508);
nand U7310 (N_7310,N_6981,N_6974);
nor U7311 (N_7311,N_6672,N_6872);
and U7312 (N_7312,N_6809,N_6583);
and U7313 (N_7313,N_6963,N_6629);
or U7314 (N_7314,N_6754,N_6589);
nand U7315 (N_7315,N_6928,N_6895);
nor U7316 (N_7316,N_6531,N_6914);
xnor U7317 (N_7317,N_6830,N_6913);
xor U7318 (N_7318,N_6964,N_6752);
xor U7319 (N_7319,N_6877,N_6711);
nor U7320 (N_7320,N_6772,N_6514);
or U7321 (N_7321,N_6950,N_6812);
and U7322 (N_7322,N_6958,N_6910);
nor U7323 (N_7323,N_6950,N_6737);
nor U7324 (N_7324,N_6791,N_6504);
nor U7325 (N_7325,N_6921,N_6762);
nor U7326 (N_7326,N_6668,N_6603);
nand U7327 (N_7327,N_6565,N_6964);
and U7328 (N_7328,N_6982,N_6952);
and U7329 (N_7329,N_6516,N_6604);
nand U7330 (N_7330,N_6644,N_6812);
nor U7331 (N_7331,N_6805,N_6959);
nand U7332 (N_7332,N_6675,N_6563);
or U7333 (N_7333,N_6773,N_6590);
and U7334 (N_7334,N_6879,N_6676);
or U7335 (N_7335,N_6819,N_6689);
and U7336 (N_7336,N_6627,N_6865);
nor U7337 (N_7337,N_6978,N_6985);
nand U7338 (N_7338,N_6893,N_6955);
xor U7339 (N_7339,N_6669,N_6657);
nand U7340 (N_7340,N_6605,N_6618);
and U7341 (N_7341,N_6666,N_6872);
and U7342 (N_7342,N_6770,N_6929);
nand U7343 (N_7343,N_6563,N_6812);
and U7344 (N_7344,N_6860,N_6504);
nand U7345 (N_7345,N_6868,N_6850);
nand U7346 (N_7346,N_6970,N_6570);
and U7347 (N_7347,N_6995,N_6816);
and U7348 (N_7348,N_6713,N_6579);
nor U7349 (N_7349,N_6552,N_6768);
nor U7350 (N_7350,N_6832,N_6999);
xor U7351 (N_7351,N_6956,N_6591);
or U7352 (N_7352,N_6897,N_6914);
nand U7353 (N_7353,N_6504,N_6983);
and U7354 (N_7354,N_6847,N_6551);
nand U7355 (N_7355,N_6986,N_6574);
xnor U7356 (N_7356,N_6583,N_6584);
nand U7357 (N_7357,N_6854,N_6612);
xor U7358 (N_7358,N_6889,N_6989);
nand U7359 (N_7359,N_6668,N_6606);
nor U7360 (N_7360,N_6759,N_6656);
nand U7361 (N_7361,N_6609,N_6580);
or U7362 (N_7362,N_6670,N_6600);
nand U7363 (N_7363,N_6930,N_6583);
nand U7364 (N_7364,N_6717,N_6846);
nor U7365 (N_7365,N_6840,N_6564);
xor U7366 (N_7366,N_6799,N_6949);
nor U7367 (N_7367,N_6797,N_6842);
nor U7368 (N_7368,N_6618,N_6653);
xnor U7369 (N_7369,N_6509,N_6746);
and U7370 (N_7370,N_6780,N_6800);
and U7371 (N_7371,N_6738,N_6752);
nor U7372 (N_7372,N_6568,N_6724);
or U7373 (N_7373,N_6529,N_6991);
xor U7374 (N_7374,N_6797,N_6696);
or U7375 (N_7375,N_6778,N_6727);
xnor U7376 (N_7376,N_6836,N_6688);
nor U7377 (N_7377,N_6607,N_6504);
xor U7378 (N_7378,N_6884,N_6750);
nand U7379 (N_7379,N_6998,N_6946);
xnor U7380 (N_7380,N_6721,N_6838);
nand U7381 (N_7381,N_6925,N_6882);
nand U7382 (N_7382,N_6940,N_6882);
xnor U7383 (N_7383,N_6753,N_6738);
nor U7384 (N_7384,N_6588,N_6666);
nand U7385 (N_7385,N_6937,N_6606);
nand U7386 (N_7386,N_6893,N_6750);
nand U7387 (N_7387,N_6851,N_6727);
and U7388 (N_7388,N_6814,N_6622);
and U7389 (N_7389,N_6687,N_6714);
nand U7390 (N_7390,N_6559,N_6831);
or U7391 (N_7391,N_6757,N_6738);
nor U7392 (N_7392,N_6727,N_6755);
nor U7393 (N_7393,N_6561,N_6529);
and U7394 (N_7394,N_6858,N_6663);
or U7395 (N_7395,N_6776,N_6504);
or U7396 (N_7396,N_6794,N_6926);
nand U7397 (N_7397,N_6704,N_6931);
and U7398 (N_7398,N_6584,N_6989);
and U7399 (N_7399,N_6607,N_6524);
xnor U7400 (N_7400,N_6983,N_6864);
xor U7401 (N_7401,N_6531,N_6778);
nor U7402 (N_7402,N_6610,N_6698);
and U7403 (N_7403,N_6576,N_6806);
nand U7404 (N_7404,N_6572,N_6748);
xor U7405 (N_7405,N_6842,N_6535);
or U7406 (N_7406,N_6875,N_6782);
or U7407 (N_7407,N_6798,N_6707);
or U7408 (N_7408,N_6944,N_6766);
or U7409 (N_7409,N_6988,N_6670);
nand U7410 (N_7410,N_6634,N_6817);
nand U7411 (N_7411,N_6882,N_6859);
or U7412 (N_7412,N_6620,N_6540);
and U7413 (N_7413,N_6545,N_6514);
or U7414 (N_7414,N_6985,N_6514);
xnor U7415 (N_7415,N_6629,N_6728);
nand U7416 (N_7416,N_6954,N_6919);
nor U7417 (N_7417,N_6661,N_6755);
nand U7418 (N_7418,N_6876,N_6872);
nand U7419 (N_7419,N_6875,N_6953);
nor U7420 (N_7420,N_6508,N_6781);
or U7421 (N_7421,N_6790,N_6871);
xor U7422 (N_7422,N_6895,N_6857);
and U7423 (N_7423,N_6998,N_6886);
or U7424 (N_7424,N_6863,N_6503);
xnor U7425 (N_7425,N_6613,N_6852);
or U7426 (N_7426,N_6747,N_6635);
or U7427 (N_7427,N_6652,N_6590);
and U7428 (N_7428,N_6994,N_6910);
or U7429 (N_7429,N_6928,N_6817);
or U7430 (N_7430,N_6968,N_6501);
or U7431 (N_7431,N_6995,N_6919);
xor U7432 (N_7432,N_6716,N_6879);
nand U7433 (N_7433,N_6791,N_6509);
nand U7434 (N_7434,N_6914,N_6561);
and U7435 (N_7435,N_6766,N_6764);
or U7436 (N_7436,N_6600,N_6936);
nor U7437 (N_7437,N_6703,N_6826);
nor U7438 (N_7438,N_6653,N_6665);
nand U7439 (N_7439,N_6807,N_6508);
nand U7440 (N_7440,N_6743,N_6661);
nor U7441 (N_7441,N_6763,N_6765);
xnor U7442 (N_7442,N_6594,N_6971);
or U7443 (N_7443,N_6516,N_6998);
nor U7444 (N_7444,N_6711,N_6707);
xor U7445 (N_7445,N_6635,N_6680);
or U7446 (N_7446,N_6901,N_6898);
nor U7447 (N_7447,N_6590,N_6780);
nand U7448 (N_7448,N_6784,N_6849);
nor U7449 (N_7449,N_6526,N_6914);
nand U7450 (N_7450,N_6727,N_6949);
nand U7451 (N_7451,N_6829,N_6611);
xnor U7452 (N_7452,N_6552,N_6550);
and U7453 (N_7453,N_6750,N_6789);
xnor U7454 (N_7454,N_6996,N_6830);
and U7455 (N_7455,N_6683,N_6936);
nand U7456 (N_7456,N_6605,N_6504);
or U7457 (N_7457,N_6524,N_6697);
nand U7458 (N_7458,N_6772,N_6848);
or U7459 (N_7459,N_6737,N_6885);
xnor U7460 (N_7460,N_6732,N_6870);
nand U7461 (N_7461,N_6716,N_6516);
xnor U7462 (N_7462,N_6709,N_6661);
or U7463 (N_7463,N_6890,N_6671);
nor U7464 (N_7464,N_6934,N_6929);
or U7465 (N_7465,N_6922,N_6950);
nand U7466 (N_7466,N_6790,N_6890);
or U7467 (N_7467,N_6747,N_6710);
nand U7468 (N_7468,N_6506,N_6550);
or U7469 (N_7469,N_6501,N_6911);
and U7470 (N_7470,N_6522,N_6899);
or U7471 (N_7471,N_6750,N_6699);
xor U7472 (N_7472,N_6820,N_6697);
and U7473 (N_7473,N_6900,N_6547);
xor U7474 (N_7474,N_6613,N_6680);
or U7475 (N_7475,N_6840,N_6893);
xnor U7476 (N_7476,N_6516,N_6992);
or U7477 (N_7477,N_6929,N_6986);
and U7478 (N_7478,N_6555,N_6678);
or U7479 (N_7479,N_6770,N_6784);
nor U7480 (N_7480,N_6619,N_6711);
xnor U7481 (N_7481,N_6784,N_6591);
xnor U7482 (N_7482,N_6923,N_6884);
or U7483 (N_7483,N_6542,N_6796);
xor U7484 (N_7484,N_6861,N_6781);
nor U7485 (N_7485,N_6571,N_6939);
or U7486 (N_7486,N_6920,N_6809);
or U7487 (N_7487,N_6769,N_6682);
or U7488 (N_7488,N_6785,N_6874);
nand U7489 (N_7489,N_6613,N_6973);
nand U7490 (N_7490,N_6840,N_6912);
xor U7491 (N_7491,N_6949,N_6932);
nor U7492 (N_7492,N_6783,N_6887);
or U7493 (N_7493,N_6875,N_6752);
nand U7494 (N_7494,N_6588,N_6553);
or U7495 (N_7495,N_6707,N_6603);
nand U7496 (N_7496,N_6969,N_6513);
nand U7497 (N_7497,N_6753,N_6779);
nand U7498 (N_7498,N_6658,N_6631);
or U7499 (N_7499,N_6791,N_6588);
nand U7500 (N_7500,N_7256,N_7075);
and U7501 (N_7501,N_7045,N_7096);
nor U7502 (N_7502,N_7266,N_7193);
nand U7503 (N_7503,N_7363,N_7206);
nand U7504 (N_7504,N_7413,N_7458);
and U7505 (N_7505,N_7109,N_7497);
nand U7506 (N_7506,N_7235,N_7416);
nor U7507 (N_7507,N_7414,N_7084);
xnor U7508 (N_7508,N_7349,N_7319);
or U7509 (N_7509,N_7032,N_7291);
xor U7510 (N_7510,N_7384,N_7324);
and U7511 (N_7511,N_7415,N_7073);
and U7512 (N_7512,N_7483,N_7473);
or U7513 (N_7513,N_7217,N_7371);
nand U7514 (N_7514,N_7447,N_7432);
nand U7515 (N_7515,N_7167,N_7429);
nand U7516 (N_7516,N_7452,N_7309);
nor U7517 (N_7517,N_7239,N_7000);
nand U7518 (N_7518,N_7488,N_7176);
nand U7519 (N_7519,N_7214,N_7022);
or U7520 (N_7520,N_7436,N_7301);
nand U7521 (N_7521,N_7086,N_7188);
xor U7522 (N_7522,N_7281,N_7372);
xnor U7523 (N_7523,N_7146,N_7407);
nand U7524 (N_7524,N_7278,N_7476);
xor U7525 (N_7525,N_7289,N_7139);
nor U7526 (N_7526,N_7168,N_7249);
nand U7527 (N_7527,N_7016,N_7264);
nor U7528 (N_7528,N_7333,N_7240);
nor U7529 (N_7529,N_7216,N_7008);
xnor U7530 (N_7530,N_7190,N_7156);
and U7531 (N_7531,N_7150,N_7378);
xnor U7532 (N_7532,N_7338,N_7160);
or U7533 (N_7533,N_7445,N_7236);
nand U7534 (N_7534,N_7177,N_7388);
nor U7535 (N_7535,N_7268,N_7002);
xor U7536 (N_7536,N_7035,N_7387);
nand U7537 (N_7537,N_7392,N_7058);
and U7538 (N_7538,N_7263,N_7020);
or U7539 (N_7539,N_7283,N_7007);
or U7540 (N_7540,N_7307,N_7316);
or U7541 (N_7541,N_7197,N_7230);
xnor U7542 (N_7542,N_7358,N_7229);
and U7543 (N_7543,N_7171,N_7438);
xor U7544 (N_7544,N_7039,N_7344);
and U7545 (N_7545,N_7009,N_7061);
and U7546 (N_7546,N_7012,N_7159);
nor U7547 (N_7547,N_7325,N_7332);
nor U7548 (N_7548,N_7042,N_7192);
and U7549 (N_7549,N_7311,N_7290);
or U7550 (N_7550,N_7466,N_7199);
xor U7551 (N_7551,N_7106,N_7318);
xnor U7552 (N_7552,N_7469,N_7345);
or U7553 (N_7553,N_7468,N_7180);
or U7554 (N_7554,N_7437,N_7356);
nand U7555 (N_7555,N_7145,N_7470);
xnor U7556 (N_7556,N_7010,N_7487);
xnor U7557 (N_7557,N_7201,N_7148);
nor U7558 (N_7558,N_7183,N_7011);
or U7559 (N_7559,N_7120,N_7243);
or U7560 (N_7560,N_7433,N_7315);
xnor U7561 (N_7561,N_7082,N_7037);
xnor U7562 (N_7562,N_7444,N_7124);
and U7563 (N_7563,N_7248,N_7280);
xnor U7564 (N_7564,N_7129,N_7089);
nand U7565 (N_7565,N_7398,N_7152);
nor U7566 (N_7566,N_7453,N_7080);
or U7567 (N_7567,N_7153,N_7136);
and U7568 (N_7568,N_7259,N_7285);
and U7569 (N_7569,N_7222,N_7021);
and U7570 (N_7570,N_7361,N_7001);
nand U7571 (N_7571,N_7182,N_7261);
or U7572 (N_7572,N_7454,N_7114);
and U7573 (N_7573,N_7040,N_7006);
or U7574 (N_7574,N_7303,N_7155);
and U7575 (N_7575,N_7127,N_7165);
and U7576 (N_7576,N_7133,N_7421);
and U7577 (N_7577,N_7110,N_7059);
nand U7578 (N_7578,N_7149,N_7360);
and U7579 (N_7579,N_7245,N_7134);
and U7580 (N_7580,N_7386,N_7401);
and U7581 (N_7581,N_7163,N_7296);
and U7582 (N_7582,N_7463,N_7339);
nand U7583 (N_7583,N_7232,N_7379);
nor U7584 (N_7584,N_7317,N_7026);
nand U7585 (N_7585,N_7158,N_7265);
nand U7586 (N_7586,N_7288,N_7352);
nand U7587 (N_7587,N_7081,N_7342);
nand U7588 (N_7588,N_7471,N_7485);
or U7589 (N_7589,N_7383,N_7065);
and U7590 (N_7590,N_7431,N_7277);
or U7591 (N_7591,N_7043,N_7094);
xnor U7592 (N_7592,N_7178,N_7088);
xnor U7593 (N_7593,N_7018,N_7353);
nor U7594 (N_7594,N_7068,N_7169);
nor U7595 (N_7595,N_7375,N_7422);
or U7596 (N_7596,N_7271,N_7287);
nand U7597 (N_7597,N_7166,N_7412);
or U7598 (N_7598,N_7117,N_7226);
and U7599 (N_7599,N_7337,N_7119);
xor U7600 (N_7600,N_7403,N_7064);
or U7601 (N_7601,N_7121,N_7292);
and U7602 (N_7602,N_7434,N_7479);
nor U7603 (N_7603,N_7198,N_7396);
or U7604 (N_7604,N_7126,N_7400);
xor U7605 (N_7605,N_7449,N_7213);
and U7606 (N_7606,N_7099,N_7308);
or U7607 (N_7607,N_7365,N_7448);
nand U7608 (N_7608,N_7368,N_7210);
nor U7609 (N_7609,N_7297,N_7340);
nor U7610 (N_7610,N_7402,N_7184);
and U7611 (N_7611,N_7326,N_7464);
nor U7612 (N_7612,N_7406,N_7204);
xor U7613 (N_7613,N_7175,N_7461);
xnor U7614 (N_7614,N_7279,N_7474);
and U7615 (N_7615,N_7257,N_7147);
xnor U7616 (N_7616,N_7202,N_7393);
nor U7617 (N_7617,N_7275,N_7328);
xor U7618 (N_7618,N_7395,N_7072);
nand U7619 (N_7619,N_7382,N_7131);
xor U7620 (N_7620,N_7046,N_7066);
nand U7621 (N_7621,N_7215,N_7189);
nand U7622 (N_7622,N_7460,N_7252);
xnor U7623 (N_7623,N_7354,N_7496);
or U7624 (N_7624,N_7376,N_7404);
and U7625 (N_7625,N_7334,N_7427);
xor U7626 (N_7626,N_7273,N_7298);
nand U7627 (N_7627,N_7049,N_7357);
nand U7628 (N_7628,N_7013,N_7241);
and U7629 (N_7629,N_7142,N_7377);
and U7630 (N_7630,N_7385,N_7170);
and U7631 (N_7631,N_7036,N_7098);
nor U7632 (N_7632,N_7227,N_7397);
xnor U7633 (N_7633,N_7237,N_7052);
nand U7634 (N_7634,N_7380,N_7472);
and U7635 (N_7635,N_7172,N_7220);
nand U7636 (N_7636,N_7456,N_7137);
nand U7637 (N_7637,N_7212,N_7033);
nand U7638 (N_7638,N_7095,N_7087);
xnor U7639 (N_7639,N_7076,N_7459);
xor U7640 (N_7640,N_7154,N_7442);
nand U7641 (N_7641,N_7242,N_7348);
and U7642 (N_7642,N_7195,N_7313);
or U7643 (N_7643,N_7441,N_7200);
or U7644 (N_7644,N_7304,N_7302);
nor U7645 (N_7645,N_7439,N_7027);
xor U7646 (N_7646,N_7091,N_7105);
nor U7647 (N_7647,N_7462,N_7381);
xor U7648 (N_7648,N_7116,N_7260);
or U7649 (N_7649,N_7102,N_7221);
and U7650 (N_7650,N_7262,N_7209);
xnor U7651 (N_7651,N_7218,N_7330);
or U7652 (N_7652,N_7205,N_7366);
or U7653 (N_7653,N_7113,N_7369);
xor U7654 (N_7654,N_7092,N_7420);
nand U7655 (N_7655,N_7069,N_7362);
xor U7656 (N_7656,N_7100,N_7250);
and U7657 (N_7657,N_7122,N_7132);
nor U7658 (N_7658,N_7219,N_7181);
xnor U7659 (N_7659,N_7062,N_7244);
nor U7660 (N_7660,N_7491,N_7327);
and U7661 (N_7661,N_7054,N_7034);
and U7662 (N_7662,N_7104,N_7017);
xor U7663 (N_7663,N_7482,N_7305);
nor U7664 (N_7664,N_7194,N_7004);
or U7665 (N_7665,N_7295,N_7481);
or U7666 (N_7666,N_7029,N_7467);
or U7667 (N_7667,N_7067,N_7495);
nand U7668 (N_7668,N_7071,N_7079);
and U7669 (N_7669,N_7128,N_7196);
and U7670 (N_7670,N_7424,N_7103);
nor U7671 (N_7671,N_7351,N_7314);
nand U7672 (N_7672,N_7480,N_7329);
xor U7673 (N_7673,N_7428,N_7053);
xor U7674 (N_7674,N_7320,N_7331);
nor U7675 (N_7675,N_7093,N_7486);
nor U7676 (N_7676,N_7499,N_7225);
nor U7677 (N_7677,N_7247,N_7173);
xnor U7678 (N_7678,N_7151,N_7475);
nand U7679 (N_7679,N_7123,N_7030);
and U7680 (N_7680,N_7389,N_7233);
xnor U7681 (N_7681,N_7272,N_7135);
or U7682 (N_7682,N_7055,N_7097);
nor U7683 (N_7683,N_7208,N_7355);
xnor U7684 (N_7684,N_7455,N_7370);
nand U7685 (N_7685,N_7490,N_7423);
nand U7686 (N_7686,N_7115,N_7228);
xor U7687 (N_7687,N_7294,N_7391);
xnor U7688 (N_7688,N_7258,N_7418);
or U7689 (N_7689,N_7083,N_7350);
nor U7690 (N_7690,N_7270,N_7174);
or U7691 (N_7691,N_7161,N_7410);
and U7692 (N_7692,N_7057,N_7435);
nor U7693 (N_7693,N_7457,N_7276);
or U7694 (N_7694,N_7187,N_7077);
xor U7695 (N_7695,N_7364,N_7191);
or U7696 (N_7696,N_7185,N_7108);
nand U7697 (N_7697,N_7028,N_7443);
or U7698 (N_7698,N_7112,N_7025);
and U7699 (N_7699,N_7321,N_7111);
nand U7700 (N_7700,N_7101,N_7269);
and U7701 (N_7701,N_7090,N_7254);
or U7702 (N_7702,N_7143,N_7405);
nand U7703 (N_7703,N_7477,N_7107);
or U7704 (N_7704,N_7478,N_7005);
or U7705 (N_7705,N_7323,N_7019);
or U7706 (N_7706,N_7203,N_7419);
nor U7707 (N_7707,N_7231,N_7041);
xor U7708 (N_7708,N_7425,N_7207);
nand U7709 (N_7709,N_7138,N_7335);
nand U7710 (N_7710,N_7408,N_7446);
nor U7711 (N_7711,N_7223,N_7050);
nand U7712 (N_7712,N_7038,N_7224);
or U7713 (N_7713,N_7253,N_7267);
nor U7714 (N_7714,N_7063,N_7031);
nand U7715 (N_7715,N_7234,N_7312);
nand U7716 (N_7716,N_7238,N_7373);
or U7717 (N_7717,N_7465,N_7056);
nor U7718 (N_7718,N_7003,N_7274);
or U7719 (N_7719,N_7014,N_7394);
or U7720 (N_7720,N_7359,N_7399);
nor U7721 (N_7721,N_7284,N_7024);
nand U7722 (N_7722,N_7440,N_7417);
and U7723 (N_7723,N_7498,N_7282);
and U7724 (N_7724,N_7157,N_7374);
and U7725 (N_7725,N_7306,N_7347);
nand U7726 (N_7726,N_7343,N_7484);
xor U7727 (N_7727,N_7336,N_7078);
nand U7728 (N_7728,N_7450,N_7118);
nand U7729 (N_7729,N_7390,N_7489);
nor U7730 (N_7730,N_7048,N_7051);
and U7731 (N_7731,N_7186,N_7125);
nand U7732 (N_7732,N_7060,N_7411);
nand U7733 (N_7733,N_7140,N_7300);
and U7734 (N_7734,N_7130,N_7144);
and U7735 (N_7735,N_7141,N_7310);
xor U7736 (N_7736,N_7246,N_7070);
or U7737 (N_7737,N_7492,N_7015);
or U7738 (N_7738,N_7251,N_7179);
nand U7739 (N_7739,N_7085,N_7023);
or U7740 (N_7740,N_7164,N_7255);
or U7741 (N_7741,N_7430,N_7367);
nor U7742 (N_7742,N_7346,N_7286);
nor U7743 (N_7743,N_7293,N_7494);
nand U7744 (N_7744,N_7299,N_7322);
xnor U7745 (N_7745,N_7044,N_7341);
and U7746 (N_7746,N_7074,N_7162);
or U7747 (N_7747,N_7451,N_7211);
nor U7748 (N_7748,N_7047,N_7493);
nor U7749 (N_7749,N_7409,N_7426);
xnor U7750 (N_7750,N_7171,N_7457);
or U7751 (N_7751,N_7040,N_7167);
nand U7752 (N_7752,N_7353,N_7111);
nor U7753 (N_7753,N_7170,N_7359);
or U7754 (N_7754,N_7483,N_7439);
xor U7755 (N_7755,N_7463,N_7486);
and U7756 (N_7756,N_7173,N_7123);
and U7757 (N_7757,N_7154,N_7033);
or U7758 (N_7758,N_7194,N_7360);
nand U7759 (N_7759,N_7369,N_7463);
nor U7760 (N_7760,N_7352,N_7280);
and U7761 (N_7761,N_7174,N_7139);
or U7762 (N_7762,N_7334,N_7330);
nor U7763 (N_7763,N_7031,N_7042);
nor U7764 (N_7764,N_7248,N_7330);
nand U7765 (N_7765,N_7046,N_7383);
nand U7766 (N_7766,N_7341,N_7017);
xor U7767 (N_7767,N_7219,N_7104);
nor U7768 (N_7768,N_7315,N_7047);
xnor U7769 (N_7769,N_7222,N_7085);
or U7770 (N_7770,N_7084,N_7357);
or U7771 (N_7771,N_7411,N_7267);
xnor U7772 (N_7772,N_7223,N_7376);
xor U7773 (N_7773,N_7407,N_7436);
nand U7774 (N_7774,N_7409,N_7154);
nor U7775 (N_7775,N_7135,N_7379);
xnor U7776 (N_7776,N_7467,N_7219);
and U7777 (N_7777,N_7290,N_7335);
nand U7778 (N_7778,N_7216,N_7274);
nor U7779 (N_7779,N_7031,N_7361);
nor U7780 (N_7780,N_7290,N_7432);
or U7781 (N_7781,N_7356,N_7237);
or U7782 (N_7782,N_7178,N_7297);
nor U7783 (N_7783,N_7151,N_7072);
and U7784 (N_7784,N_7246,N_7243);
nor U7785 (N_7785,N_7094,N_7134);
and U7786 (N_7786,N_7040,N_7003);
xor U7787 (N_7787,N_7115,N_7014);
or U7788 (N_7788,N_7461,N_7056);
and U7789 (N_7789,N_7179,N_7379);
or U7790 (N_7790,N_7428,N_7160);
xnor U7791 (N_7791,N_7298,N_7047);
xnor U7792 (N_7792,N_7078,N_7077);
xor U7793 (N_7793,N_7149,N_7306);
or U7794 (N_7794,N_7248,N_7290);
nor U7795 (N_7795,N_7149,N_7300);
nand U7796 (N_7796,N_7027,N_7332);
nor U7797 (N_7797,N_7404,N_7153);
or U7798 (N_7798,N_7211,N_7181);
nor U7799 (N_7799,N_7198,N_7061);
nor U7800 (N_7800,N_7458,N_7465);
xor U7801 (N_7801,N_7465,N_7382);
and U7802 (N_7802,N_7208,N_7146);
xnor U7803 (N_7803,N_7352,N_7125);
nand U7804 (N_7804,N_7415,N_7262);
xor U7805 (N_7805,N_7467,N_7194);
nand U7806 (N_7806,N_7404,N_7493);
nor U7807 (N_7807,N_7029,N_7119);
xor U7808 (N_7808,N_7472,N_7170);
or U7809 (N_7809,N_7247,N_7419);
nand U7810 (N_7810,N_7001,N_7393);
nand U7811 (N_7811,N_7404,N_7256);
nand U7812 (N_7812,N_7240,N_7103);
and U7813 (N_7813,N_7303,N_7080);
xor U7814 (N_7814,N_7177,N_7009);
or U7815 (N_7815,N_7338,N_7387);
nor U7816 (N_7816,N_7229,N_7055);
nor U7817 (N_7817,N_7093,N_7362);
or U7818 (N_7818,N_7363,N_7484);
nor U7819 (N_7819,N_7328,N_7087);
nor U7820 (N_7820,N_7257,N_7093);
xnor U7821 (N_7821,N_7204,N_7461);
or U7822 (N_7822,N_7146,N_7401);
or U7823 (N_7823,N_7013,N_7243);
nand U7824 (N_7824,N_7077,N_7004);
or U7825 (N_7825,N_7185,N_7222);
nor U7826 (N_7826,N_7281,N_7472);
nor U7827 (N_7827,N_7491,N_7042);
and U7828 (N_7828,N_7262,N_7347);
xnor U7829 (N_7829,N_7282,N_7095);
or U7830 (N_7830,N_7213,N_7079);
xor U7831 (N_7831,N_7094,N_7300);
nand U7832 (N_7832,N_7315,N_7497);
xnor U7833 (N_7833,N_7264,N_7174);
and U7834 (N_7834,N_7118,N_7339);
or U7835 (N_7835,N_7359,N_7224);
nor U7836 (N_7836,N_7415,N_7356);
xnor U7837 (N_7837,N_7238,N_7363);
xor U7838 (N_7838,N_7026,N_7453);
xor U7839 (N_7839,N_7254,N_7374);
nand U7840 (N_7840,N_7096,N_7496);
or U7841 (N_7841,N_7113,N_7168);
nor U7842 (N_7842,N_7252,N_7220);
xor U7843 (N_7843,N_7223,N_7153);
nor U7844 (N_7844,N_7375,N_7142);
nor U7845 (N_7845,N_7417,N_7353);
or U7846 (N_7846,N_7416,N_7378);
and U7847 (N_7847,N_7445,N_7299);
nor U7848 (N_7848,N_7206,N_7117);
nor U7849 (N_7849,N_7494,N_7459);
nand U7850 (N_7850,N_7281,N_7336);
nor U7851 (N_7851,N_7192,N_7096);
nand U7852 (N_7852,N_7130,N_7042);
nor U7853 (N_7853,N_7300,N_7368);
nand U7854 (N_7854,N_7093,N_7467);
xor U7855 (N_7855,N_7480,N_7149);
or U7856 (N_7856,N_7365,N_7236);
nand U7857 (N_7857,N_7097,N_7436);
and U7858 (N_7858,N_7282,N_7397);
xor U7859 (N_7859,N_7114,N_7369);
xnor U7860 (N_7860,N_7490,N_7112);
or U7861 (N_7861,N_7088,N_7280);
nor U7862 (N_7862,N_7293,N_7300);
or U7863 (N_7863,N_7018,N_7001);
nand U7864 (N_7864,N_7075,N_7096);
nand U7865 (N_7865,N_7158,N_7134);
nor U7866 (N_7866,N_7476,N_7472);
or U7867 (N_7867,N_7024,N_7414);
nor U7868 (N_7868,N_7260,N_7466);
xor U7869 (N_7869,N_7267,N_7287);
and U7870 (N_7870,N_7445,N_7149);
nand U7871 (N_7871,N_7353,N_7044);
and U7872 (N_7872,N_7256,N_7154);
nand U7873 (N_7873,N_7163,N_7337);
and U7874 (N_7874,N_7162,N_7032);
or U7875 (N_7875,N_7380,N_7335);
and U7876 (N_7876,N_7144,N_7367);
or U7877 (N_7877,N_7387,N_7256);
nand U7878 (N_7878,N_7435,N_7007);
or U7879 (N_7879,N_7110,N_7116);
or U7880 (N_7880,N_7301,N_7273);
nor U7881 (N_7881,N_7267,N_7449);
nand U7882 (N_7882,N_7439,N_7063);
and U7883 (N_7883,N_7208,N_7248);
or U7884 (N_7884,N_7354,N_7468);
nand U7885 (N_7885,N_7361,N_7343);
xnor U7886 (N_7886,N_7032,N_7180);
nand U7887 (N_7887,N_7236,N_7414);
nand U7888 (N_7888,N_7170,N_7167);
or U7889 (N_7889,N_7138,N_7041);
and U7890 (N_7890,N_7239,N_7220);
or U7891 (N_7891,N_7253,N_7488);
xor U7892 (N_7892,N_7207,N_7276);
xnor U7893 (N_7893,N_7479,N_7318);
and U7894 (N_7894,N_7124,N_7295);
and U7895 (N_7895,N_7382,N_7393);
and U7896 (N_7896,N_7400,N_7183);
and U7897 (N_7897,N_7381,N_7077);
nand U7898 (N_7898,N_7270,N_7177);
or U7899 (N_7899,N_7074,N_7043);
and U7900 (N_7900,N_7306,N_7160);
nor U7901 (N_7901,N_7421,N_7187);
or U7902 (N_7902,N_7005,N_7053);
nor U7903 (N_7903,N_7054,N_7330);
and U7904 (N_7904,N_7235,N_7253);
nand U7905 (N_7905,N_7491,N_7351);
xor U7906 (N_7906,N_7348,N_7317);
and U7907 (N_7907,N_7340,N_7022);
nand U7908 (N_7908,N_7023,N_7479);
nor U7909 (N_7909,N_7449,N_7375);
and U7910 (N_7910,N_7069,N_7461);
and U7911 (N_7911,N_7381,N_7100);
and U7912 (N_7912,N_7316,N_7198);
or U7913 (N_7913,N_7188,N_7121);
nor U7914 (N_7914,N_7457,N_7095);
nor U7915 (N_7915,N_7091,N_7073);
and U7916 (N_7916,N_7113,N_7193);
and U7917 (N_7917,N_7496,N_7083);
or U7918 (N_7918,N_7019,N_7132);
and U7919 (N_7919,N_7154,N_7101);
nor U7920 (N_7920,N_7421,N_7449);
xor U7921 (N_7921,N_7488,N_7425);
nand U7922 (N_7922,N_7348,N_7332);
or U7923 (N_7923,N_7234,N_7268);
nor U7924 (N_7924,N_7386,N_7240);
nand U7925 (N_7925,N_7434,N_7180);
and U7926 (N_7926,N_7118,N_7180);
and U7927 (N_7927,N_7284,N_7217);
xnor U7928 (N_7928,N_7329,N_7372);
nand U7929 (N_7929,N_7390,N_7404);
and U7930 (N_7930,N_7196,N_7428);
or U7931 (N_7931,N_7060,N_7330);
xnor U7932 (N_7932,N_7043,N_7068);
xnor U7933 (N_7933,N_7437,N_7477);
or U7934 (N_7934,N_7100,N_7384);
nand U7935 (N_7935,N_7228,N_7397);
or U7936 (N_7936,N_7466,N_7247);
xnor U7937 (N_7937,N_7324,N_7200);
or U7938 (N_7938,N_7241,N_7065);
nand U7939 (N_7939,N_7261,N_7101);
and U7940 (N_7940,N_7276,N_7113);
xor U7941 (N_7941,N_7351,N_7040);
nand U7942 (N_7942,N_7233,N_7194);
xor U7943 (N_7943,N_7472,N_7272);
nand U7944 (N_7944,N_7071,N_7349);
nor U7945 (N_7945,N_7007,N_7213);
nand U7946 (N_7946,N_7468,N_7250);
and U7947 (N_7947,N_7274,N_7201);
xnor U7948 (N_7948,N_7129,N_7316);
and U7949 (N_7949,N_7133,N_7327);
or U7950 (N_7950,N_7170,N_7412);
nor U7951 (N_7951,N_7077,N_7136);
and U7952 (N_7952,N_7030,N_7237);
or U7953 (N_7953,N_7237,N_7207);
nor U7954 (N_7954,N_7302,N_7309);
or U7955 (N_7955,N_7407,N_7011);
nor U7956 (N_7956,N_7164,N_7251);
xor U7957 (N_7957,N_7075,N_7232);
nor U7958 (N_7958,N_7476,N_7432);
nor U7959 (N_7959,N_7278,N_7489);
and U7960 (N_7960,N_7025,N_7323);
or U7961 (N_7961,N_7024,N_7207);
and U7962 (N_7962,N_7355,N_7220);
or U7963 (N_7963,N_7139,N_7381);
or U7964 (N_7964,N_7279,N_7310);
or U7965 (N_7965,N_7466,N_7325);
or U7966 (N_7966,N_7026,N_7248);
nand U7967 (N_7967,N_7223,N_7363);
xnor U7968 (N_7968,N_7234,N_7226);
nand U7969 (N_7969,N_7279,N_7086);
nor U7970 (N_7970,N_7005,N_7101);
nand U7971 (N_7971,N_7230,N_7354);
nor U7972 (N_7972,N_7017,N_7235);
xnor U7973 (N_7973,N_7371,N_7399);
or U7974 (N_7974,N_7306,N_7243);
nor U7975 (N_7975,N_7467,N_7113);
and U7976 (N_7976,N_7282,N_7046);
and U7977 (N_7977,N_7031,N_7032);
xor U7978 (N_7978,N_7198,N_7019);
nand U7979 (N_7979,N_7181,N_7054);
nor U7980 (N_7980,N_7446,N_7121);
and U7981 (N_7981,N_7209,N_7210);
and U7982 (N_7982,N_7111,N_7286);
nor U7983 (N_7983,N_7367,N_7129);
nor U7984 (N_7984,N_7027,N_7414);
or U7985 (N_7985,N_7411,N_7263);
nand U7986 (N_7986,N_7306,N_7020);
and U7987 (N_7987,N_7177,N_7122);
nor U7988 (N_7988,N_7175,N_7128);
and U7989 (N_7989,N_7079,N_7416);
xor U7990 (N_7990,N_7352,N_7247);
xnor U7991 (N_7991,N_7463,N_7014);
nor U7992 (N_7992,N_7383,N_7025);
nor U7993 (N_7993,N_7343,N_7280);
nand U7994 (N_7994,N_7386,N_7031);
xnor U7995 (N_7995,N_7423,N_7127);
xor U7996 (N_7996,N_7344,N_7402);
nand U7997 (N_7997,N_7150,N_7230);
or U7998 (N_7998,N_7068,N_7150);
nor U7999 (N_7999,N_7157,N_7492);
nor U8000 (N_8000,N_7908,N_7795);
xnor U8001 (N_8001,N_7827,N_7800);
nand U8002 (N_8002,N_7713,N_7724);
and U8003 (N_8003,N_7929,N_7890);
and U8004 (N_8004,N_7869,N_7938);
nor U8005 (N_8005,N_7695,N_7544);
or U8006 (N_8006,N_7793,N_7792);
nand U8007 (N_8007,N_7794,N_7801);
nor U8008 (N_8008,N_7732,N_7741);
xor U8009 (N_8009,N_7930,N_7865);
or U8010 (N_8010,N_7567,N_7956);
or U8011 (N_8011,N_7615,N_7691);
or U8012 (N_8012,N_7555,N_7513);
nor U8013 (N_8013,N_7876,N_7642);
and U8014 (N_8014,N_7599,N_7603);
xor U8015 (N_8015,N_7650,N_7970);
xnor U8016 (N_8016,N_7996,N_7565);
or U8017 (N_8017,N_7980,N_7592);
nand U8018 (N_8018,N_7822,N_7504);
xor U8019 (N_8019,N_7804,N_7781);
nor U8020 (N_8020,N_7645,N_7813);
nor U8021 (N_8021,N_7805,N_7569);
xnor U8022 (N_8022,N_7632,N_7553);
nor U8023 (N_8023,N_7923,N_7641);
xnor U8024 (N_8024,N_7944,N_7806);
or U8025 (N_8025,N_7959,N_7653);
and U8026 (N_8026,N_7867,N_7767);
or U8027 (N_8027,N_7943,N_7772);
nor U8028 (N_8028,N_7681,N_7643);
nand U8029 (N_8029,N_7976,N_7882);
nor U8030 (N_8030,N_7937,N_7647);
xor U8031 (N_8031,N_7639,N_7593);
or U8032 (N_8032,N_7849,N_7658);
xnor U8033 (N_8033,N_7942,N_7935);
xor U8034 (N_8034,N_7954,N_7836);
xor U8035 (N_8035,N_7963,N_7936);
and U8036 (N_8036,N_7987,N_7564);
nand U8037 (N_8037,N_7534,N_7861);
xnor U8038 (N_8038,N_7674,N_7893);
xnor U8039 (N_8039,N_7973,N_7608);
and U8040 (N_8040,N_7939,N_7558);
nand U8041 (N_8041,N_7560,N_7711);
or U8042 (N_8042,N_7840,N_7699);
nor U8043 (N_8043,N_7521,N_7562);
nand U8044 (N_8044,N_7576,N_7831);
or U8045 (N_8045,N_7633,N_7759);
and U8046 (N_8046,N_7843,N_7702);
nor U8047 (N_8047,N_7978,N_7766);
xnor U8048 (N_8048,N_7610,N_7878);
nand U8049 (N_8049,N_7541,N_7587);
or U8050 (N_8050,N_7539,N_7689);
nor U8051 (N_8051,N_7517,N_7907);
nand U8052 (N_8052,N_7900,N_7966);
and U8053 (N_8053,N_7991,N_7749);
xor U8054 (N_8054,N_7515,N_7850);
or U8055 (N_8055,N_7789,N_7500);
or U8056 (N_8056,N_7809,N_7946);
or U8057 (N_8057,N_7656,N_7915);
or U8058 (N_8058,N_7769,N_7510);
and U8059 (N_8059,N_7928,N_7543);
xnor U8060 (N_8060,N_7685,N_7715);
xnor U8061 (N_8061,N_7596,N_7780);
nor U8062 (N_8062,N_7718,N_7514);
and U8063 (N_8063,N_7950,N_7965);
nand U8064 (N_8064,N_7802,N_7547);
and U8065 (N_8065,N_7888,N_7590);
xnor U8066 (N_8066,N_7579,N_7649);
and U8067 (N_8067,N_7858,N_7644);
or U8068 (N_8068,N_7824,N_7548);
nand U8069 (N_8069,N_7927,N_7670);
xor U8070 (N_8070,N_7984,N_7595);
nor U8071 (N_8071,N_7648,N_7771);
or U8072 (N_8072,N_7652,N_7982);
xor U8073 (N_8073,N_7763,N_7953);
and U8074 (N_8074,N_7873,N_7785);
and U8075 (N_8075,N_7667,N_7631);
xnor U8076 (N_8076,N_7559,N_7744);
nor U8077 (N_8077,N_7725,N_7941);
or U8078 (N_8078,N_7584,N_7975);
xnor U8079 (N_8079,N_7846,N_7743);
nor U8080 (N_8080,N_7518,N_7512);
or U8081 (N_8081,N_7669,N_7556);
or U8082 (N_8082,N_7527,N_7625);
nor U8083 (N_8083,N_7952,N_7971);
xor U8084 (N_8084,N_7524,N_7997);
nand U8085 (N_8085,N_7550,N_7851);
nor U8086 (N_8086,N_7756,N_7619);
or U8087 (N_8087,N_7845,N_7630);
nor U8088 (N_8088,N_7945,N_7676);
xor U8089 (N_8089,N_7828,N_7777);
nor U8090 (N_8090,N_7529,N_7750);
nand U8091 (N_8091,N_7602,N_7583);
and U8092 (N_8092,N_7716,N_7852);
nor U8093 (N_8093,N_7951,N_7784);
xor U8094 (N_8094,N_7796,N_7662);
nor U8095 (N_8095,N_7621,N_7617);
and U8096 (N_8096,N_7572,N_7705);
xor U8097 (N_8097,N_7968,N_7707);
or U8098 (N_8098,N_7932,N_7825);
and U8099 (N_8099,N_7889,N_7549);
xor U8100 (N_8100,N_7773,N_7540);
nand U8101 (N_8101,N_7783,N_7764);
nor U8102 (N_8102,N_7819,N_7877);
and U8103 (N_8103,N_7508,N_7934);
or U8104 (N_8104,N_7838,N_7886);
and U8105 (N_8105,N_7812,N_7629);
and U8106 (N_8106,N_7910,N_7790);
nor U8107 (N_8107,N_7628,N_7995);
or U8108 (N_8108,N_7964,N_7989);
and U8109 (N_8109,N_7906,N_7501);
nor U8110 (N_8110,N_7606,N_7916);
xor U8111 (N_8111,N_7891,N_7526);
nor U8112 (N_8112,N_7791,N_7779);
nand U8113 (N_8113,N_7918,N_7671);
xnor U8114 (N_8114,N_7727,N_7992);
or U8115 (N_8115,N_7651,N_7519);
nor U8116 (N_8116,N_7697,N_7881);
and U8117 (N_8117,N_7775,N_7638);
nor U8118 (N_8118,N_7757,N_7884);
and U8119 (N_8119,N_7589,N_7672);
nand U8120 (N_8120,N_7655,N_7530);
and U8121 (N_8121,N_7532,N_7566);
or U8122 (N_8122,N_7815,N_7646);
nor U8123 (N_8123,N_7575,N_7879);
and U8124 (N_8124,N_7611,N_7730);
nand U8125 (N_8125,N_7974,N_7626);
xnor U8126 (N_8126,N_7758,N_7588);
and U8127 (N_8127,N_7640,N_7538);
nand U8128 (N_8128,N_7620,N_7854);
nand U8129 (N_8129,N_7803,N_7578);
nor U8130 (N_8130,N_7753,N_7859);
or U8131 (N_8131,N_7925,N_7533);
nor U8132 (N_8132,N_7511,N_7998);
xnor U8133 (N_8133,N_7823,N_7622);
or U8134 (N_8134,N_7736,N_7692);
xor U8135 (N_8135,N_7690,N_7969);
or U8136 (N_8136,N_7726,N_7598);
xnor U8137 (N_8137,N_7913,N_7684);
and U8138 (N_8138,N_7693,N_7563);
xor U8139 (N_8139,N_7537,N_7568);
or U8140 (N_8140,N_7922,N_7931);
or U8141 (N_8141,N_7712,N_7687);
nand U8142 (N_8142,N_7990,N_7573);
or U8143 (N_8143,N_7847,N_7797);
xor U8144 (N_8144,N_7799,N_7940);
nand U8145 (N_8145,N_7614,N_7503);
nand U8146 (N_8146,N_7604,N_7731);
nand U8147 (N_8147,N_7830,N_7546);
xnor U8148 (N_8148,N_7832,N_7875);
or U8149 (N_8149,N_7751,N_7844);
xor U8150 (N_8150,N_7542,N_7708);
nor U8151 (N_8151,N_7586,N_7755);
nor U8152 (N_8152,N_7600,N_7871);
or U8153 (N_8153,N_7580,N_7762);
xor U8154 (N_8154,N_7505,N_7597);
and U8155 (N_8155,N_7577,N_7798);
xor U8156 (N_8156,N_7682,N_7735);
nand U8157 (N_8157,N_7901,N_7894);
or U8158 (N_8158,N_7680,N_7778);
nand U8159 (N_8159,N_7960,N_7709);
and U8160 (N_8160,N_7788,N_7782);
nor U8161 (N_8161,N_7627,N_7921);
or U8162 (N_8162,N_7665,N_7637);
nor U8163 (N_8163,N_7862,N_7898);
or U8164 (N_8164,N_7745,N_7748);
nor U8165 (N_8165,N_7892,N_7752);
nand U8166 (N_8166,N_7839,N_7666);
nor U8167 (N_8167,N_7818,N_7754);
nand U8168 (N_8168,N_7591,N_7912);
nor U8169 (N_8169,N_7686,N_7520);
xor U8170 (N_8170,N_7833,N_7863);
and U8171 (N_8171,N_7961,N_7919);
or U8172 (N_8172,N_7636,N_7986);
xor U8173 (N_8173,N_7856,N_7948);
nor U8174 (N_8174,N_7955,N_7739);
or U8175 (N_8175,N_7820,N_7988);
or U8176 (N_8176,N_7904,N_7634);
nand U8177 (N_8177,N_7826,N_7897);
and U8178 (N_8178,N_7874,N_7623);
and U8179 (N_8179,N_7612,N_7883);
nor U8180 (N_8180,N_7765,N_7723);
xor U8181 (N_8181,N_7994,N_7594);
and U8182 (N_8182,N_7853,N_7770);
and U8183 (N_8183,N_7981,N_7917);
nor U8184 (N_8184,N_7761,N_7535);
xnor U8185 (N_8185,N_7677,N_7860);
nand U8186 (N_8186,N_7554,N_7857);
or U8187 (N_8187,N_7842,N_7525);
nor U8188 (N_8188,N_7523,N_7841);
nand U8189 (N_8189,N_7509,N_7866);
nand U8190 (N_8190,N_7909,N_7679);
and U8191 (N_8191,N_7581,N_7811);
nor U8192 (N_8192,N_7816,N_7659);
nor U8193 (N_8193,N_7962,N_7872);
and U8194 (N_8194,N_7885,N_7507);
xnor U8195 (N_8195,N_7911,N_7786);
xor U8196 (N_8196,N_7657,N_7660);
nand U8197 (N_8197,N_7920,N_7949);
and U8198 (N_8198,N_7678,N_7808);
xnor U8199 (N_8199,N_7516,N_7821);
nor U8200 (N_8200,N_7895,N_7701);
or U8201 (N_8201,N_7582,N_7902);
nand U8202 (N_8202,N_7967,N_7561);
and U8203 (N_8203,N_7664,N_7574);
or U8204 (N_8204,N_7545,N_7896);
xor U8205 (N_8205,N_7663,N_7933);
xor U8206 (N_8206,N_7720,N_7864);
xnor U8207 (N_8207,N_7710,N_7722);
and U8208 (N_8208,N_7635,N_7835);
xor U8209 (N_8209,N_7719,N_7585);
nand U8210 (N_8210,N_7848,N_7760);
and U8211 (N_8211,N_7729,N_7536);
nor U8212 (N_8212,N_7887,N_7570);
and U8213 (N_8213,N_7528,N_7605);
and U8214 (N_8214,N_7924,N_7829);
nand U8215 (N_8215,N_7675,N_7870);
nor U8216 (N_8216,N_7698,N_7721);
nand U8217 (N_8217,N_7926,N_7977);
nor U8218 (N_8218,N_7601,N_7683);
and U8219 (N_8219,N_7714,N_7983);
nand U8220 (N_8220,N_7696,N_7899);
xnor U8221 (N_8221,N_7737,N_7993);
xnor U8222 (N_8222,N_7740,N_7837);
nor U8223 (N_8223,N_7807,N_7728);
nand U8224 (N_8224,N_7768,N_7673);
xor U8225 (N_8225,N_7742,N_7903);
xor U8226 (N_8226,N_7502,N_7914);
xor U8227 (N_8227,N_7506,N_7624);
and U8228 (N_8228,N_7834,N_7787);
nor U8229 (N_8229,N_7817,N_7814);
and U8230 (N_8230,N_7703,N_7571);
and U8231 (N_8231,N_7957,N_7979);
xnor U8232 (N_8232,N_7947,N_7958);
nor U8233 (N_8233,N_7738,N_7616);
nor U8234 (N_8234,N_7717,N_7880);
or U8235 (N_8235,N_7905,N_7747);
and U8236 (N_8236,N_7734,N_7774);
nor U8237 (N_8237,N_7618,N_7694);
and U8238 (N_8238,N_7704,N_7522);
and U8239 (N_8239,N_7706,N_7552);
xnor U8240 (N_8240,N_7700,N_7668);
nand U8241 (N_8241,N_7607,N_7531);
xor U8242 (N_8242,N_7661,N_7999);
nand U8243 (N_8243,N_7985,N_7654);
xor U8244 (N_8244,N_7613,N_7972);
or U8245 (N_8245,N_7733,N_7688);
xnor U8246 (N_8246,N_7551,N_7776);
and U8247 (N_8247,N_7557,N_7868);
nor U8248 (N_8248,N_7810,N_7609);
nor U8249 (N_8249,N_7746,N_7855);
xor U8250 (N_8250,N_7839,N_7837);
and U8251 (N_8251,N_7503,N_7630);
nor U8252 (N_8252,N_7885,N_7963);
and U8253 (N_8253,N_7536,N_7760);
and U8254 (N_8254,N_7953,N_7761);
nand U8255 (N_8255,N_7672,N_7899);
nand U8256 (N_8256,N_7980,N_7959);
nor U8257 (N_8257,N_7898,N_7995);
nand U8258 (N_8258,N_7737,N_7710);
nand U8259 (N_8259,N_7717,N_7538);
xor U8260 (N_8260,N_7718,N_7662);
nand U8261 (N_8261,N_7715,N_7578);
and U8262 (N_8262,N_7823,N_7870);
nor U8263 (N_8263,N_7779,N_7928);
or U8264 (N_8264,N_7940,N_7670);
nor U8265 (N_8265,N_7577,N_7837);
nor U8266 (N_8266,N_7858,N_7786);
nor U8267 (N_8267,N_7991,N_7563);
or U8268 (N_8268,N_7977,N_7746);
or U8269 (N_8269,N_7827,N_7859);
nand U8270 (N_8270,N_7746,N_7729);
or U8271 (N_8271,N_7576,N_7690);
or U8272 (N_8272,N_7802,N_7973);
or U8273 (N_8273,N_7680,N_7660);
or U8274 (N_8274,N_7749,N_7691);
nand U8275 (N_8275,N_7560,N_7659);
nand U8276 (N_8276,N_7970,N_7850);
xnor U8277 (N_8277,N_7514,N_7592);
nor U8278 (N_8278,N_7625,N_7958);
and U8279 (N_8279,N_7845,N_7949);
and U8280 (N_8280,N_7911,N_7631);
xor U8281 (N_8281,N_7549,N_7864);
xor U8282 (N_8282,N_7956,N_7731);
nor U8283 (N_8283,N_7696,N_7637);
nor U8284 (N_8284,N_7547,N_7521);
or U8285 (N_8285,N_7528,N_7832);
or U8286 (N_8286,N_7947,N_7900);
and U8287 (N_8287,N_7651,N_7971);
xor U8288 (N_8288,N_7896,N_7919);
nand U8289 (N_8289,N_7656,N_7798);
nor U8290 (N_8290,N_7637,N_7921);
xor U8291 (N_8291,N_7746,N_7878);
xnor U8292 (N_8292,N_7532,N_7715);
and U8293 (N_8293,N_7613,N_7814);
nand U8294 (N_8294,N_7882,N_7662);
nor U8295 (N_8295,N_7608,N_7744);
nor U8296 (N_8296,N_7744,N_7999);
nor U8297 (N_8297,N_7812,N_7840);
nand U8298 (N_8298,N_7992,N_7851);
or U8299 (N_8299,N_7804,N_7671);
and U8300 (N_8300,N_7753,N_7622);
or U8301 (N_8301,N_7900,N_7773);
or U8302 (N_8302,N_7716,N_7547);
nand U8303 (N_8303,N_7712,N_7895);
nor U8304 (N_8304,N_7851,N_7560);
and U8305 (N_8305,N_7592,N_7656);
nor U8306 (N_8306,N_7806,N_7991);
or U8307 (N_8307,N_7716,N_7984);
nand U8308 (N_8308,N_7522,N_7504);
nor U8309 (N_8309,N_7981,N_7998);
nand U8310 (N_8310,N_7936,N_7508);
xor U8311 (N_8311,N_7768,N_7860);
and U8312 (N_8312,N_7846,N_7695);
nand U8313 (N_8313,N_7638,N_7724);
nor U8314 (N_8314,N_7725,N_7571);
nand U8315 (N_8315,N_7880,N_7714);
nand U8316 (N_8316,N_7621,N_7985);
xor U8317 (N_8317,N_7882,N_7733);
xnor U8318 (N_8318,N_7863,N_7634);
xnor U8319 (N_8319,N_7923,N_7824);
nor U8320 (N_8320,N_7723,N_7857);
nand U8321 (N_8321,N_7519,N_7578);
nor U8322 (N_8322,N_7753,N_7930);
nand U8323 (N_8323,N_7934,N_7797);
and U8324 (N_8324,N_7918,N_7503);
nor U8325 (N_8325,N_7765,N_7960);
nand U8326 (N_8326,N_7545,N_7723);
nor U8327 (N_8327,N_7928,N_7569);
and U8328 (N_8328,N_7679,N_7880);
nor U8329 (N_8329,N_7885,N_7606);
nand U8330 (N_8330,N_7994,N_7811);
or U8331 (N_8331,N_7964,N_7559);
nor U8332 (N_8332,N_7787,N_7892);
nor U8333 (N_8333,N_7942,N_7883);
and U8334 (N_8334,N_7763,N_7792);
xor U8335 (N_8335,N_7504,N_7858);
or U8336 (N_8336,N_7756,N_7835);
nor U8337 (N_8337,N_7761,N_7693);
or U8338 (N_8338,N_7694,N_7561);
and U8339 (N_8339,N_7647,N_7983);
and U8340 (N_8340,N_7608,N_7511);
nand U8341 (N_8341,N_7967,N_7983);
nor U8342 (N_8342,N_7878,N_7603);
or U8343 (N_8343,N_7770,N_7817);
nand U8344 (N_8344,N_7998,N_7930);
or U8345 (N_8345,N_7655,N_7940);
nand U8346 (N_8346,N_7630,N_7678);
and U8347 (N_8347,N_7661,N_7829);
nor U8348 (N_8348,N_7903,N_7730);
and U8349 (N_8349,N_7504,N_7502);
xnor U8350 (N_8350,N_7760,N_7922);
nand U8351 (N_8351,N_7911,N_7611);
nor U8352 (N_8352,N_7743,N_7515);
xor U8353 (N_8353,N_7685,N_7560);
xor U8354 (N_8354,N_7834,N_7747);
or U8355 (N_8355,N_7518,N_7997);
nor U8356 (N_8356,N_7645,N_7573);
or U8357 (N_8357,N_7871,N_7960);
nor U8358 (N_8358,N_7815,N_7505);
xnor U8359 (N_8359,N_7990,N_7661);
nor U8360 (N_8360,N_7742,N_7731);
and U8361 (N_8361,N_7855,N_7625);
xnor U8362 (N_8362,N_7515,N_7583);
nor U8363 (N_8363,N_7752,N_7999);
xor U8364 (N_8364,N_7606,N_7730);
nor U8365 (N_8365,N_7776,N_7665);
xnor U8366 (N_8366,N_7882,N_7910);
or U8367 (N_8367,N_7989,N_7864);
nand U8368 (N_8368,N_7634,N_7746);
or U8369 (N_8369,N_7622,N_7695);
nand U8370 (N_8370,N_7702,N_7740);
or U8371 (N_8371,N_7652,N_7740);
nand U8372 (N_8372,N_7765,N_7833);
nor U8373 (N_8373,N_7919,N_7528);
or U8374 (N_8374,N_7629,N_7914);
nor U8375 (N_8375,N_7913,N_7509);
or U8376 (N_8376,N_7538,N_7819);
nand U8377 (N_8377,N_7843,N_7846);
or U8378 (N_8378,N_7964,N_7978);
and U8379 (N_8379,N_7783,N_7711);
nor U8380 (N_8380,N_7686,N_7811);
nand U8381 (N_8381,N_7749,N_7686);
nor U8382 (N_8382,N_7914,N_7950);
and U8383 (N_8383,N_7514,N_7614);
and U8384 (N_8384,N_7739,N_7576);
or U8385 (N_8385,N_7940,N_7745);
and U8386 (N_8386,N_7760,N_7836);
and U8387 (N_8387,N_7722,N_7977);
and U8388 (N_8388,N_7622,N_7541);
or U8389 (N_8389,N_7789,N_7677);
nand U8390 (N_8390,N_7838,N_7992);
nand U8391 (N_8391,N_7928,N_7636);
nor U8392 (N_8392,N_7891,N_7694);
nand U8393 (N_8393,N_7834,N_7611);
nor U8394 (N_8394,N_7937,N_7684);
nand U8395 (N_8395,N_7945,N_7703);
nor U8396 (N_8396,N_7591,N_7851);
nor U8397 (N_8397,N_7592,N_7864);
and U8398 (N_8398,N_7647,N_7569);
and U8399 (N_8399,N_7752,N_7539);
or U8400 (N_8400,N_7718,N_7767);
nand U8401 (N_8401,N_7613,N_7668);
nor U8402 (N_8402,N_7689,N_7525);
xor U8403 (N_8403,N_7709,N_7690);
and U8404 (N_8404,N_7977,N_7984);
or U8405 (N_8405,N_7527,N_7573);
or U8406 (N_8406,N_7948,N_7852);
xor U8407 (N_8407,N_7655,N_7944);
nor U8408 (N_8408,N_7541,N_7955);
and U8409 (N_8409,N_7741,N_7669);
nor U8410 (N_8410,N_7581,N_7850);
and U8411 (N_8411,N_7760,N_7893);
xor U8412 (N_8412,N_7910,N_7661);
or U8413 (N_8413,N_7647,N_7939);
or U8414 (N_8414,N_7768,N_7839);
xor U8415 (N_8415,N_7802,N_7858);
nor U8416 (N_8416,N_7576,N_7634);
nand U8417 (N_8417,N_7840,N_7684);
or U8418 (N_8418,N_7931,N_7514);
or U8419 (N_8419,N_7534,N_7902);
xor U8420 (N_8420,N_7760,N_7607);
or U8421 (N_8421,N_7820,N_7558);
xor U8422 (N_8422,N_7914,N_7983);
and U8423 (N_8423,N_7594,N_7702);
and U8424 (N_8424,N_7913,N_7916);
nand U8425 (N_8425,N_7735,N_7815);
nor U8426 (N_8426,N_7741,N_7918);
or U8427 (N_8427,N_7925,N_7941);
nor U8428 (N_8428,N_7706,N_7609);
or U8429 (N_8429,N_7804,N_7703);
and U8430 (N_8430,N_7705,N_7563);
xnor U8431 (N_8431,N_7522,N_7761);
nand U8432 (N_8432,N_7939,N_7731);
nand U8433 (N_8433,N_7685,N_7546);
xor U8434 (N_8434,N_7844,N_7813);
xor U8435 (N_8435,N_7623,N_7890);
xor U8436 (N_8436,N_7616,N_7756);
or U8437 (N_8437,N_7905,N_7863);
and U8438 (N_8438,N_7605,N_7663);
nand U8439 (N_8439,N_7931,N_7864);
nor U8440 (N_8440,N_7881,N_7795);
nand U8441 (N_8441,N_7693,N_7696);
and U8442 (N_8442,N_7773,N_7851);
nor U8443 (N_8443,N_7734,N_7723);
or U8444 (N_8444,N_7570,N_7609);
or U8445 (N_8445,N_7920,N_7829);
or U8446 (N_8446,N_7799,N_7587);
xor U8447 (N_8447,N_7605,N_7863);
xor U8448 (N_8448,N_7703,N_7573);
nor U8449 (N_8449,N_7816,N_7817);
nor U8450 (N_8450,N_7531,N_7650);
nand U8451 (N_8451,N_7667,N_7500);
xnor U8452 (N_8452,N_7939,N_7769);
or U8453 (N_8453,N_7724,N_7895);
xnor U8454 (N_8454,N_7648,N_7518);
and U8455 (N_8455,N_7568,N_7579);
or U8456 (N_8456,N_7707,N_7949);
nor U8457 (N_8457,N_7960,N_7828);
nor U8458 (N_8458,N_7592,N_7651);
nand U8459 (N_8459,N_7918,N_7912);
nand U8460 (N_8460,N_7899,N_7940);
and U8461 (N_8461,N_7833,N_7826);
nand U8462 (N_8462,N_7640,N_7559);
or U8463 (N_8463,N_7730,N_7904);
nor U8464 (N_8464,N_7610,N_7834);
and U8465 (N_8465,N_7971,N_7655);
and U8466 (N_8466,N_7988,N_7545);
nor U8467 (N_8467,N_7750,N_7691);
xor U8468 (N_8468,N_7638,N_7680);
nand U8469 (N_8469,N_7735,N_7616);
or U8470 (N_8470,N_7959,N_7902);
and U8471 (N_8471,N_7848,N_7799);
and U8472 (N_8472,N_7661,N_7916);
xor U8473 (N_8473,N_7620,N_7954);
and U8474 (N_8474,N_7659,N_7577);
and U8475 (N_8475,N_7580,N_7749);
nor U8476 (N_8476,N_7755,N_7772);
xor U8477 (N_8477,N_7859,N_7734);
nand U8478 (N_8478,N_7850,N_7810);
xnor U8479 (N_8479,N_7874,N_7551);
or U8480 (N_8480,N_7705,N_7596);
or U8481 (N_8481,N_7903,N_7698);
and U8482 (N_8482,N_7871,N_7799);
and U8483 (N_8483,N_7805,N_7688);
and U8484 (N_8484,N_7874,N_7628);
and U8485 (N_8485,N_7942,N_7714);
or U8486 (N_8486,N_7993,N_7578);
xnor U8487 (N_8487,N_7662,N_7675);
nand U8488 (N_8488,N_7587,N_7770);
nor U8489 (N_8489,N_7805,N_7684);
xnor U8490 (N_8490,N_7621,N_7642);
and U8491 (N_8491,N_7702,N_7672);
xnor U8492 (N_8492,N_7789,N_7824);
nand U8493 (N_8493,N_7539,N_7680);
xor U8494 (N_8494,N_7898,N_7882);
or U8495 (N_8495,N_7977,N_7713);
nand U8496 (N_8496,N_7525,N_7879);
and U8497 (N_8497,N_7810,N_7746);
or U8498 (N_8498,N_7525,N_7931);
nor U8499 (N_8499,N_7606,N_7984);
or U8500 (N_8500,N_8454,N_8393);
or U8501 (N_8501,N_8182,N_8145);
or U8502 (N_8502,N_8401,N_8423);
nor U8503 (N_8503,N_8297,N_8239);
or U8504 (N_8504,N_8242,N_8064);
or U8505 (N_8505,N_8309,N_8281);
or U8506 (N_8506,N_8057,N_8267);
and U8507 (N_8507,N_8303,N_8439);
nand U8508 (N_8508,N_8336,N_8089);
xnor U8509 (N_8509,N_8348,N_8105);
xor U8510 (N_8510,N_8042,N_8301);
nor U8511 (N_8511,N_8080,N_8453);
nor U8512 (N_8512,N_8160,N_8295);
and U8513 (N_8513,N_8065,N_8441);
and U8514 (N_8514,N_8021,N_8358);
nand U8515 (N_8515,N_8285,N_8005);
or U8516 (N_8516,N_8070,N_8487);
and U8517 (N_8517,N_8258,N_8485);
or U8518 (N_8518,N_8055,N_8433);
xnor U8519 (N_8519,N_8354,N_8186);
xor U8520 (N_8520,N_8168,N_8227);
nor U8521 (N_8521,N_8253,N_8394);
nor U8522 (N_8522,N_8015,N_8233);
or U8523 (N_8523,N_8202,N_8130);
and U8524 (N_8524,N_8096,N_8094);
and U8525 (N_8525,N_8032,N_8197);
nor U8526 (N_8526,N_8151,N_8254);
nand U8527 (N_8527,N_8109,N_8405);
nand U8528 (N_8528,N_8238,N_8156);
and U8529 (N_8529,N_8184,N_8035);
nor U8530 (N_8530,N_8463,N_8283);
xnor U8531 (N_8531,N_8178,N_8325);
nand U8532 (N_8532,N_8058,N_8273);
nor U8533 (N_8533,N_8322,N_8078);
xor U8534 (N_8534,N_8472,N_8249);
nand U8535 (N_8535,N_8025,N_8210);
nor U8536 (N_8536,N_8189,N_8101);
and U8537 (N_8537,N_8396,N_8050);
xnor U8538 (N_8538,N_8061,N_8246);
nand U8539 (N_8539,N_8215,N_8469);
xnor U8540 (N_8540,N_8222,N_8046);
or U8541 (N_8541,N_8365,N_8428);
nor U8542 (N_8542,N_8279,N_8288);
nand U8543 (N_8543,N_8087,N_8123);
nor U8544 (N_8544,N_8430,N_8024);
or U8545 (N_8545,N_8033,N_8257);
nor U8546 (N_8546,N_8172,N_8136);
nor U8547 (N_8547,N_8334,N_8196);
or U8548 (N_8548,N_8415,N_8079);
nor U8549 (N_8549,N_8175,N_8290);
or U8550 (N_8550,N_8038,N_8434);
xor U8551 (N_8551,N_8417,N_8459);
nor U8552 (N_8552,N_8116,N_8241);
xor U8553 (N_8553,N_8011,N_8438);
nand U8554 (N_8554,N_8170,N_8216);
nor U8555 (N_8555,N_8308,N_8353);
nor U8556 (N_8556,N_8131,N_8384);
nand U8557 (N_8557,N_8444,N_8041);
and U8558 (N_8558,N_8107,N_8187);
and U8559 (N_8559,N_8134,N_8474);
and U8560 (N_8560,N_8299,N_8022);
nor U8561 (N_8561,N_8263,N_8104);
nand U8562 (N_8562,N_8318,N_8012);
or U8563 (N_8563,N_8014,N_8375);
nand U8564 (N_8564,N_8352,N_8237);
xnor U8565 (N_8565,N_8490,N_8207);
and U8566 (N_8566,N_8044,N_8199);
and U8567 (N_8567,N_8436,N_8460);
xnor U8568 (N_8568,N_8223,N_8408);
nor U8569 (N_8569,N_8464,N_8016);
nand U8570 (N_8570,N_8007,N_8244);
xnor U8571 (N_8571,N_8225,N_8208);
or U8572 (N_8572,N_8129,N_8133);
nor U8573 (N_8573,N_8072,N_8378);
and U8574 (N_8574,N_8009,N_8001);
xor U8575 (N_8575,N_8086,N_8496);
or U8576 (N_8576,N_8114,N_8435);
nand U8577 (N_8577,N_8037,N_8473);
nand U8578 (N_8578,N_8491,N_8478);
nand U8579 (N_8579,N_8219,N_8306);
nand U8580 (N_8580,N_8211,N_8240);
and U8581 (N_8581,N_8218,N_8363);
and U8582 (N_8582,N_8250,N_8406);
xor U8583 (N_8583,N_8482,N_8135);
or U8584 (N_8584,N_8385,N_8204);
xnor U8585 (N_8585,N_8390,N_8316);
xnor U8586 (N_8586,N_8402,N_8403);
or U8587 (N_8587,N_8088,N_8243);
nand U8588 (N_8588,N_8339,N_8071);
xnor U8589 (N_8589,N_8304,N_8040);
nand U8590 (N_8590,N_8455,N_8000);
nand U8591 (N_8591,N_8117,N_8426);
and U8592 (N_8592,N_8023,N_8361);
xnor U8593 (N_8593,N_8293,N_8280);
or U8594 (N_8594,N_8359,N_8262);
nand U8595 (N_8595,N_8122,N_8251);
nand U8596 (N_8596,N_8127,N_8150);
nand U8597 (N_8597,N_8261,N_8128);
nor U8598 (N_8598,N_8180,N_8458);
and U8599 (N_8599,N_8447,N_8412);
nand U8600 (N_8600,N_8108,N_8201);
and U8601 (N_8601,N_8260,N_8326);
nor U8602 (N_8602,N_8320,N_8450);
nor U8603 (N_8603,N_8143,N_8422);
xor U8604 (N_8604,N_8315,N_8159);
and U8605 (N_8605,N_8154,N_8291);
or U8606 (N_8606,N_8067,N_8062);
or U8607 (N_8607,N_8083,N_8468);
xnor U8608 (N_8608,N_8307,N_8333);
nor U8609 (N_8609,N_8418,N_8093);
nand U8610 (N_8610,N_8410,N_8097);
xor U8611 (N_8611,N_8051,N_8031);
nor U8612 (N_8612,N_8486,N_8395);
and U8613 (N_8613,N_8466,N_8442);
nand U8614 (N_8614,N_8355,N_8125);
nand U8615 (N_8615,N_8179,N_8224);
nor U8616 (N_8616,N_8347,N_8443);
xor U8617 (N_8617,N_8121,N_8462);
nor U8618 (N_8618,N_8092,N_8386);
or U8619 (N_8619,N_8248,N_8198);
xor U8620 (N_8620,N_8158,N_8006);
xor U8621 (N_8621,N_8142,N_8271);
or U8622 (N_8622,N_8028,N_8029);
and U8623 (N_8623,N_8467,N_8185);
nand U8624 (N_8624,N_8076,N_8327);
or U8625 (N_8625,N_8205,N_8282);
or U8626 (N_8626,N_8465,N_8372);
nor U8627 (N_8627,N_8494,N_8177);
nor U8628 (N_8628,N_8157,N_8342);
and U8629 (N_8629,N_8409,N_8118);
or U8630 (N_8630,N_8445,N_8312);
nor U8631 (N_8631,N_8212,N_8321);
xnor U8632 (N_8632,N_8077,N_8099);
and U8633 (N_8633,N_8167,N_8457);
or U8634 (N_8634,N_8337,N_8477);
nor U8635 (N_8635,N_8300,N_8027);
nand U8636 (N_8636,N_8475,N_8499);
xor U8637 (N_8637,N_8020,N_8330);
nor U8638 (N_8638,N_8095,N_8146);
nand U8639 (N_8639,N_8343,N_8139);
or U8640 (N_8640,N_8416,N_8119);
xor U8641 (N_8641,N_8338,N_8424);
nand U8642 (N_8642,N_8013,N_8010);
or U8643 (N_8643,N_8106,N_8328);
or U8644 (N_8644,N_8045,N_8413);
and U8645 (N_8645,N_8068,N_8404);
nor U8646 (N_8646,N_8421,N_8100);
xnor U8647 (N_8647,N_8230,N_8302);
or U8648 (N_8648,N_8069,N_8234);
xor U8649 (N_8649,N_8272,N_8429);
xor U8650 (N_8650,N_8488,N_8340);
nor U8651 (N_8651,N_8148,N_8493);
nor U8652 (N_8652,N_8190,N_8399);
nor U8653 (N_8653,N_8305,N_8245);
nand U8654 (N_8654,N_8018,N_8275);
xor U8655 (N_8655,N_8411,N_8432);
nand U8656 (N_8656,N_8141,N_8059);
and U8657 (N_8657,N_8296,N_8317);
nand U8658 (N_8658,N_8235,N_8360);
and U8659 (N_8659,N_8414,N_8171);
xnor U8660 (N_8660,N_8349,N_8173);
and U8661 (N_8661,N_8448,N_8252);
or U8662 (N_8662,N_8495,N_8377);
or U8663 (N_8663,N_8379,N_8226);
or U8664 (N_8664,N_8091,N_8110);
nor U8665 (N_8665,N_8373,N_8111);
and U8666 (N_8666,N_8229,N_8200);
or U8667 (N_8667,N_8098,N_8357);
nand U8668 (N_8668,N_8188,N_8102);
and U8669 (N_8669,N_8484,N_8313);
nor U8670 (N_8670,N_8419,N_8112);
or U8671 (N_8671,N_8269,N_8049);
nor U8672 (N_8672,N_8264,N_8155);
nor U8673 (N_8673,N_8203,N_8481);
nor U8674 (N_8674,N_8278,N_8228);
and U8675 (N_8675,N_8370,N_8276);
or U8676 (N_8676,N_8374,N_8060);
xnor U8677 (N_8677,N_8075,N_8169);
nand U8678 (N_8678,N_8287,N_8369);
or U8679 (N_8679,N_8480,N_8341);
or U8680 (N_8680,N_8174,N_8476);
nand U8681 (N_8681,N_8026,N_8247);
or U8682 (N_8682,N_8380,N_8124);
xnor U8683 (N_8683,N_8319,N_8213);
xor U8684 (N_8684,N_8400,N_8452);
xor U8685 (N_8685,N_8266,N_8479);
nor U8686 (N_8686,N_8073,N_8389);
nand U8687 (N_8687,N_8113,N_8449);
and U8688 (N_8688,N_8367,N_8074);
xor U8689 (N_8689,N_8346,N_8376);
or U8690 (N_8690,N_8483,N_8066);
and U8691 (N_8691,N_8497,N_8163);
and U8692 (N_8692,N_8289,N_8397);
nor U8693 (N_8693,N_8420,N_8331);
or U8694 (N_8694,N_8456,N_8206);
nand U8695 (N_8695,N_8470,N_8492);
xor U8696 (N_8696,N_8388,N_8149);
nor U8697 (N_8697,N_8221,N_8191);
nand U8698 (N_8698,N_8392,N_8161);
nand U8699 (N_8699,N_8383,N_8003);
xor U8700 (N_8700,N_8350,N_8084);
xor U8701 (N_8701,N_8398,N_8082);
xnor U8702 (N_8702,N_8183,N_8194);
and U8703 (N_8703,N_8366,N_8039);
and U8704 (N_8704,N_8209,N_8162);
nor U8705 (N_8705,N_8364,N_8220);
and U8706 (N_8706,N_8054,N_8371);
or U8707 (N_8707,N_8451,N_8292);
and U8708 (N_8708,N_8407,N_8166);
nor U8709 (N_8709,N_8498,N_8165);
nand U8710 (N_8710,N_8427,N_8034);
or U8711 (N_8711,N_8043,N_8126);
nor U8712 (N_8712,N_8085,N_8132);
and U8713 (N_8713,N_8489,N_8277);
nand U8714 (N_8714,N_8255,N_8090);
xor U8715 (N_8715,N_8298,N_8310);
nand U8716 (N_8716,N_8425,N_8138);
nor U8717 (N_8717,N_8344,N_8345);
nor U8718 (N_8718,N_8446,N_8387);
nor U8719 (N_8719,N_8368,N_8284);
and U8720 (N_8720,N_8256,N_8471);
and U8721 (N_8721,N_8053,N_8181);
xor U8722 (N_8722,N_8461,N_8236);
or U8723 (N_8723,N_8382,N_8286);
nor U8724 (N_8724,N_8314,N_8019);
xnor U8725 (N_8725,N_8120,N_8176);
and U8726 (N_8726,N_8004,N_8232);
nor U8727 (N_8727,N_8329,N_8008);
nor U8728 (N_8728,N_8324,N_8017);
xnor U8729 (N_8729,N_8323,N_8047);
and U8730 (N_8730,N_8311,N_8431);
nand U8731 (N_8731,N_8274,N_8391);
nand U8732 (N_8732,N_8192,N_8362);
or U8733 (N_8733,N_8103,N_8440);
and U8734 (N_8734,N_8048,N_8356);
xnor U8735 (N_8735,N_8115,N_8351);
or U8736 (N_8736,N_8144,N_8270);
nand U8737 (N_8737,N_8195,N_8217);
or U8738 (N_8738,N_8381,N_8164);
xor U8739 (N_8739,N_8231,N_8437);
xnor U8740 (N_8740,N_8052,N_8153);
nand U8741 (N_8741,N_8036,N_8259);
and U8742 (N_8742,N_8268,N_8193);
xor U8743 (N_8743,N_8140,N_8152);
or U8744 (N_8744,N_8214,N_8063);
or U8745 (N_8745,N_8335,N_8265);
and U8746 (N_8746,N_8081,N_8056);
nand U8747 (N_8747,N_8030,N_8294);
nor U8748 (N_8748,N_8332,N_8002);
or U8749 (N_8749,N_8147,N_8137);
nand U8750 (N_8750,N_8106,N_8274);
nand U8751 (N_8751,N_8249,N_8418);
or U8752 (N_8752,N_8331,N_8395);
nor U8753 (N_8753,N_8026,N_8235);
nor U8754 (N_8754,N_8237,N_8103);
xnor U8755 (N_8755,N_8314,N_8481);
nor U8756 (N_8756,N_8466,N_8437);
nor U8757 (N_8757,N_8206,N_8087);
xor U8758 (N_8758,N_8378,N_8011);
and U8759 (N_8759,N_8296,N_8226);
or U8760 (N_8760,N_8342,N_8203);
or U8761 (N_8761,N_8229,N_8133);
nor U8762 (N_8762,N_8420,N_8419);
nand U8763 (N_8763,N_8289,N_8490);
nor U8764 (N_8764,N_8072,N_8270);
xnor U8765 (N_8765,N_8060,N_8188);
or U8766 (N_8766,N_8157,N_8073);
and U8767 (N_8767,N_8164,N_8465);
nor U8768 (N_8768,N_8083,N_8050);
nor U8769 (N_8769,N_8358,N_8108);
xnor U8770 (N_8770,N_8087,N_8241);
nor U8771 (N_8771,N_8225,N_8041);
xnor U8772 (N_8772,N_8371,N_8009);
nor U8773 (N_8773,N_8420,N_8362);
or U8774 (N_8774,N_8338,N_8146);
nor U8775 (N_8775,N_8397,N_8052);
and U8776 (N_8776,N_8186,N_8236);
nand U8777 (N_8777,N_8320,N_8204);
or U8778 (N_8778,N_8150,N_8259);
nor U8779 (N_8779,N_8406,N_8178);
or U8780 (N_8780,N_8350,N_8473);
nand U8781 (N_8781,N_8153,N_8192);
nand U8782 (N_8782,N_8331,N_8280);
nor U8783 (N_8783,N_8322,N_8489);
xor U8784 (N_8784,N_8002,N_8210);
nor U8785 (N_8785,N_8347,N_8287);
nor U8786 (N_8786,N_8384,N_8443);
or U8787 (N_8787,N_8021,N_8363);
and U8788 (N_8788,N_8059,N_8045);
and U8789 (N_8789,N_8157,N_8055);
xnor U8790 (N_8790,N_8390,N_8194);
nor U8791 (N_8791,N_8438,N_8036);
xor U8792 (N_8792,N_8277,N_8212);
nand U8793 (N_8793,N_8275,N_8205);
nand U8794 (N_8794,N_8085,N_8260);
xnor U8795 (N_8795,N_8052,N_8310);
nand U8796 (N_8796,N_8203,N_8286);
or U8797 (N_8797,N_8486,N_8400);
nor U8798 (N_8798,N_8160,N_8251);
nand U8799 (N_8799,N_8191,N_8117);
nand U8800 (N_8800,N_8016,N_8048);
and U8801 (N_8801,N_8053,N_8442);
nor U8802 (N_8802,N_8061,N_8320);
or U8803 (N_8803,N_8324,N_8105);
nor U8804 (N_8804,N_8435,N_8471);
nand U8805 (N_8805,N_8114,N_8087);
nand U8806 (N_8806,N_8360,N_8401);
nand U8807 (N_8807,N_8324,N_8499);
or U8808 (N_8808,N_8265,N_8206);
nor U8809 (N_8809,N_8280,N_8168);
and U8810 (N_8810,N_8023,N_8475);
xor U8811 (N_8811,N_8168,N_8030);
nand U8812 (N_8812,N_8247,N_8437);
nor U8813 (N_8813,N_8114,N_8130);
nand U8814 (N_8814,N_8013,N_8451);
nor U8815 (N_8815,N_8051,N_8384);
nand U8816 (N_8816,N_8187,N_8238);
and U8817 (N_8817,N_8123,N_8259);
xnor U8818 (N_8818,N_8189,N_8148);
or U8819 (N_8819,N_8000,N_8422);
and U8820 (N_8820,N_8365,N_8278);
or U8821 (N_8821,N_8350,N_8076);
or U8822 (N_8822,N_8417,N_8082);
and U8823 (N_8823,N_8203,N_8086);
or U8824 (N_8824,N_8437,N_8107);
nand U8825 (N_8825,N_8125,N_8086);
or U8826 (N_8826,N_8455,N_8247);
and U8827 (N_8827,N_8052,N_8043);
nor U8828 (N_8828,N_8410,N_8079);
nor U8829 (N_8829,N_8206,N_8225);
xnor U8830 (N_8830,N_8479,N_8260);
nand U8831 (N_8831,N_8060,N_8224);
or U8832 (N_8832,N_8349,N_8430);
nand U8833 (N_8833,N_8000,N_8419);
xor U8834 (N_8834,N_8467,N_8144);
and U8835 (N_8835,N_8339,N_8017);
and U8836 (N_8836,N_8045,N_8471);
nand U8837 (N_8837,N_8252,N_8426);
nand U8838 (N_8838,N_8140,N_8044);
nand U8839 (N_8839,N_8275,N_8080);
or U8840 (N_8840,N_8019,N_8113);
and U8841 (N_8841,N_8027,N_8069);
and U8842 (N_8842,N_8042,N_8013);
or U8843 (N_8843,N_8145,N_8430);
and U8844 (N_8844,N_8030,N_8109);
nor U8845 (N_8845,N_8006,N_8339);
and U8846 (N_8846,N_8487,N_8444);
xor U8847 (N_8847,N_8267,N_8080);
nand U8848 (N_8848,N_8351,N_8000);
nand U8849 (N_8849,N_8108,N_8027);
and U8850 (N_8850,N_8148,N_8033);
nor U8851 (N_8851,N_8314,N_8154);
or U8852 (N_8852,N_8059,N_8239);
and U8853 (N_8853,N_8413,N_8240);
nand U8854 (N_8854,N_8021,N_8297);
and U8855 (N_8855,N_8113,N_8475);
nand U8856 (N_8856,N_8021,N_8459);
nand U8857 (N_8857,N_8044,N_8098);
nand U8858 (N_8858,N_8366,N_8350);
nor U8859 (N_8859,N_8202,N_8209);
nor U8860 (N_8860,N_8335,N_8268);
nor U8861 (N_8861,N_8070,N_8188);
xnor U8862 (N_8862,N_8307,N_8488);
nor U8863 (N_8863,N_8279,N_8417);
nor U8864 (N_8864,N_8063,N_8403);
xor U8865 (N_8865,N_8340,N_8234);
or U8866 (N_8866,N_8381,N_8455);
nor U8867 (N_8867,N_8259,N_8486);
or U8868 (N_8868,N_8162,N_8000);
nand U8869 (N_8869,N_8224,N_8448);
and U8870 (N_8870,N_8413,N_8303);
nor U8871 (N_8871,N_8486,N_8143);
nand U8872 (N_8872,N_8432,N_8122);
xor U8873 (N_8873,N_8224,N_8343);
nand U8874 (N_8874,N_8250,N_8354);
nand U8875 (N_8875,N_8052,N_8245);
nand U8876 (N_8876,N_8389,N_8109);
xnor U8877 (N_8877,N_8152,N_8046);
and U8878 (N_8878,N_8253,N_8454);
or U8879 (N_8879,N_8489,N_8324);
xnor U8880 (N_8880,N_8097,N_8400);
nand U8881 (N_8881,N_8034,N_8254);
nor U8882 (N_8882,N_8489,N_8022);
xnor U8883 (N_8883,N_8070,N_8109);
or U8884 (N_8884,N_8129,N_8075);
or U8885 (N_8885,N_8412,N_8416);
nand U8886 (N_8886,N_8128,N_8166);
xnor U8887 (N_8887,N_8191,N_8133);
and U8888 (N_8888,N_8392,N_8046);
nor U8889 (N_8889,N_8033,N_8171);
xnor U8890 (N_8890,N_8139,N_8449);
nor U8891 (N_8891,N_8357,N_8493);
nand U8892 (N_8892,N_8460,N_8388);
nand U8893 (N_8893,N_8202,N_8080);
nor U8894 (N_8894,N_8171,N_8258);
nor U8895 (N_8895,N_8455,N_8355);
and U8896 (N_8896,N_8408,N_8005);
xor U8897 (N_8897,N_8200,N_8081);
and U8898 (N_8898,N_8123,N_8346);
nand U8899 (N_8899,N_8194,N_8476);
or U8900 (N_8900,N_8430,N_8427);
and U8901 (N_8901,N_8132,N_8448);
nand U8902 (N_8902,N_8076,N_8055);
and U8903 (N_8903,N_8375,N_8445);
nor U8904 (N_8904,N_8052,N_8007);
and U8905 (N_8905,N_8080,N_8239);
xor U8906 (N_8906,N_8378,N_8410);
nand U8907 (N_8907,N_8414,N_8158);
nor U8908 (N_8908,N_8149,N_8140);
nor U8909 (N_8909,N_8170,N_8108);
nand U8910 (N_8910,N_8333,N_8131);
nor U8911 (N_8911,N_8106,N_8370);
nor U8912 (N_8912,N_8451,N_8299);
and U8913 (N_8913,N_8196,N_8467);
nor U8914 (N_8914,N_8388,N_8338);
xor U8915 (N_8915,N_8295,N_8372);
or U8916 (N_8916,N_8180,N_8452);
and U8917 (N_8917,N_8188,N_8050);
nor U8918 (N_8918,N_8427,N_8212);
or U8919 (N_8919,N_8226,N_8334);
or U8920 (N_8920,N_8215,N_8399);
and U8921 (N_8921,N_8481,N_8081);
nor U8922 (N_8922,N_8253,N_8465);
or U8923 (N_8923,N_8352,N_8437);
or U8924 (N_8924,N_8251,N_8227);
nand U8925 (N_8925,N_8083,N_8209);
nand U8926 (N_8926,N_8119,N_8180);
nor U8927 (N_8927,N_8335,N_8310);
nor U8928 (N_8928,N_8172,N_8374);
nand U8929 (N_8929,N_8484,N_8447);
or U8930 (N_8930,N_8355,N_8389);
nand U8931 (N_8931,N_8421,N_8210);
nor U8932 (N_8932,N_8321,N_8063);
and U8933 (N_8933,N_8463,N_8233);
or U8934 (N_8934,N_8344,N_8129);
xor U8935 (N_8935,N_8407,N_8187);
nor U8936 (N_8936,N_8409,N_8066);
nand U8937 (N_8937,N_8350,N_8169);
nor U8938 (N_8938,N_8219,N_8361);
xnor U8939 (N_8939,N_8022,N_8264);
or U8940 (N_8940,N_8351,N_8206);
nand U8941 (N_8941,N_8463,N_8183);
xnor U8942 (N_8942,N_8116,N_8453);
or U8943 (N_8943,N_8429,N_8238);
or U8944 (N_8944,N_8337,N_8275);
and U8945 (N_8945,N_8460,N_8148);
or U8946 (N_8946,N_8028,N_8235);
nor U8947 (N_8947,N_8211,N_8066);
nor U8948 (N_8948,N_8218,N_8000);
and U8949 (N_8949,N_8315,N_8415);
xor U8950 (N_8950,N_8075,N_8321);
or U8951 (N_8951,N_8425,N_8182);
nor U8952 (N_8952,N_8259,N_8371);
nor U8953 (N_8953,N_8162,N_8481);
xor U8954 (N_8954,N_8354,N_8024);
nor U8955 (N_8955,N_8186,N_8329);
or U8956 (N_8956,N_8480,N_8029);
or U8957 (N_8957,N_8431,N_8333);
nand U8958 (N_8958,N_8228,N_8329);
nand U8959 (N_8959,N_8108,N_8364);
nor U8960 (N_8960,N_8365,N_8147);
nand U8961 (N_8961,N_8352,N_8307);
nor U8962 (N_8962,N_8387,N_8381);
or U8963 (N_8963,N_8326,N_8389);
or U8964 (N_8964,N_8130,N_8399);
nor U8965 (N_8965,N_8109,N_8034);
nand U8966 (N_8966,N_8233,N_8433);
nor U8967 (N_8967,N_8433,N_8472);
nand U8968 (N_8968,N_8077,N_8287);
nor U8969 (N_8969,N_8031,N_8029);
nor U8970 (N_8970,N_8020,N_8445);
or U8971 (N_8971,N_8465,N_8083);
or U8972 (N_8972,N_8025,N_8196);
or U8973 (N_8973,N_8475,N_8392);
or U8974 (N_8974,N_8430,N_8120);
nand U8975 (N_8975,N_8237,N_8434);
nand U8976 (N_8976,N_8206,N_8353);
nor U8977 (N_8977,N_8427,N_8069);
xnor U8978 (N_8978,N_8243,N_8248);
nand U8979 (N_8979,N_8176,N_8156);
xor U8980 (N_8980,N_8179,N_8045);
nand U8981 (N_8981,N_8165,N_8288);
and U8982 (N_8982,N_8409,N_8117);
xnor U8983 (N_8983,N_8446,N_8328);
nor U8984 (N_8984,N_8435,N_8196);
nand U8985 (N_8985,N_8140,N_8372);
xor U8986 (N_8986,N_8082,N_8187);
and U8987 (N_8987,N_8213,N_8154);
nand U8988 (N_8988,N_8237,N_8215);
or U8989 (N_8989,N_8110,N_8054);
xor U8990 (N_8990,N_8424,N_8373);
and U8991 (N_8991,N_8489,N_8294);
nand U8992 (N_8992,N_8450,N_8267);
nand U8993 (N_8993,N_8007,N_8316);
nand U8994 (N_8994,N_8198,N_8379);
xnor U8995 (N_8995,N_8399,N_8488);
nor U8996 (N_8996,N_8280,N_8292);
nor U8997 (N_8997,N_8213,N_8395);
and U8998 (N_8998,N_8461,N_8262);
xor U8999 (N_8999,N_8291,N_8139);
and U9000 (N_9000,N_8546,N_8744);
and U9001 (N_9001,N_8808,N_8692);
xor U9002 (N_9002,N_8694,N_8535);
and U9003 (N_9003,N_8759,N_8776);
nand U9004 (N_9004,N_8953,N_8840);
nand U9005 (N_9005,N_8570,N_8997);
xor U9006 (N_9006,N_8859,N_8856);
and U9007 (N_9007,N_8940,N_8871);
nor U9008 (N_9008,N_8565,N_8966);
nand U9009 (N_9009,N_8676,N_8879);
or U9010 (N_9010,N_8616,N_8561);
or U9011 (N_9011,N_8778,N_8833);
nor U9012 (N_9012,N_8573,N_8643);
or U9013 (N_9013,N_8900,N_8787);
or U9014 (N_9014,N_8615,N_8960);
and U9015 (N_9015,N_8948,N_8606);
nand U9016 (N_9016,N_8685,N_8766);
nor U9017 (N_9017,N_8996,N_8598);
xor U9018 (N_9018,N_8939,N_8608);
nand U9019 (N_9019,N_8563,N_8624);
nor U9020 (N_9020,N_8684,N_8709);
xnor U9021 (N_9021,N_8890,N_8741);
xnor U9022 (N_9022,N_8930,N_8534);
nor U9023 (N_9023,N_8989,N_8523);
and U9024 (N_9024,N_8805,N_8780);
xnor U9025 (N_9025,N_8530,N_8500);
or U9026 (N_9026,N_8589,N_8680);
xor U9027 (N_9027,N_8786,N_8994);
or U9028 (N_9028,N_8797,N_8799);
nor U9029 (N_9029,N_8774,N_8854);
or U9030 (N_9030,N_8678,N_8739);
nand U9031 (N_9031,N_8751,N_8999);
or U9032 (N_9032,N_8941,N_8647);
or U9033 (N_9033,N_8949,N_8702);
nand U9034 (N_9034,N_8920,N_8782);
nand U9035 (N_9035,N_8807,N_8593);
or U9036 (N_9036,N_8911,N_8526);
nor U9037 (N_9037,N_8512,N_8555);
xnor U9038 (N_9038,N_8663,N_8517);
or U9039 (N_9039,N_8798,N_8897);
nand U9040 (N_9040,N_8902,N_8945);
nand U9041 (N_9041,N_8888,N_8728);
or U9042 (N_9042,N_8541,N_8677);
xor U9043 (N_9043,N_8601,N_8746);
xor U9044 (N_9044,N_8910,N_8907);
and U9045 (N_9045,N_8612,N_8794);
or U9046 (N_9046,N_8800,N_8891);
xor U9047 (N_9047,N_8659,N_8986);
or U9048 (N_9048,N_8803,N_8571);
xor U9049 (N_9049,N_8923,N_8763);
nand U9050 (N_9050,N_8642,N_8586);
xnor U9051 (N_9051,N_8935,N_8717);
or U9052 (N_9052,N_8718,N_8884);
and U9053 (N_9053,N_8864,N_8506);
nor U9054 (N_9054,N_8858,N_8756);
and U9055 (N_9055,N_8587,N_8784);
or U9056 (N_9056,N_8696,N_8823);
nor U9057 (N_9057,N_8533,N_8922);
and U9058 (N_9058,N_8625,N_8795);
or U9059 (N_9059,N_8550,N_8824);
and U9060 (N_9060,N_8671,N_8686);
nor U9061 (N_9061,N_8557,N_8826);
nand U9062 (N_9062,N_8574,N_8576);
and U9063 (N_9063,N_8820,N_8635);
or U9064 (N_9064,N_8572,N_8552);
xnor U9065 (N_9065,N_8946,N_8944);
and U9066 (N_9066,N_8981,N_8855);
or U9067 (N_9067,N_8832,N_8626);
xnor U9068 (N_9068,N_8725,N_8765);
or U9069 (N_9069,N_8841,N_8704);
nor U9070 (N_9070,N_8628,N_8700);
nand U9071 (N_9071,N_8619,N_8658);
nand U9072 (N_9072,N_8812,N_8657);
nand U9073 (N_9073,N_8967,N_8731);
or U9074 (N_9074,N_8781,N_8896);
xnor U9075 (N_9075,N_8998,N_8973);
xor U9076 (N_9076,N_8750,N_8977);
xor U9077 (N_9077,N_8822,N_8964);
and U9078 (N_9078,N_8687,N_8577);
nor U9079 (N_9079,N_8880,N_8584);
and U9080 (N_9080,N_8970,N_8847);
and U9081 (N_9081,N_8792,N_8938);
xor U9082 (N_9082,N_8919,N_8697);
xnor U9083 (N_9083,N_8852,N_8749);
xor U9084 (N_9084,N_8887,N_8633);
nor U9085 (N_9085,N_8991,N_8758);
nand U9086 (N_9086,N_8585,N_8664);
and U9087 (N_9087,N_8547,N_8599);
or U9088 (N_9088,N_8828,N_8582);
or U9089 (N_9089,N_8931,N_8761);
nand U9090 (N_9090,N_8544,N_8690);
and U9091 (N_9091,N_8992,N_8844);
and U9092 (N_9092,N_8965,N_8505);
or U9093 (N_9093,N_8933,N_8834);
and U9094 (N_9094,N_8623,N_8914);
and U9095 (N_9095,N_8532,N_8747);
nor U9096 (N_9096,N_8513,N_8733);
or U9097 (N_9097,N_8508,N_8893);
xnor U9098 (N_9098,N_8839,N_8843);
and U9099 (N_9099,N_8760,N_8915);
xnor U9100 (N_9100,N_8525,N_8668);
or U9101 (N_9101,N_8768,N_8644);
nand U9102 (N_9102,N_8894,N_8816);
xor U9103 (N_9103,N_8724,N_8762);
and U9104 (N_9104,N_8609,N_8610);
or U9105 (N_9105,N_8729,N_8982);
or U9106 (N_9106,N_8957,N_8602);
or U9107 (N_9107,N_8595,N_8885);
nand U9108 (N_9108,N_8874,N_8722);
and U9109 (N_9109,N_8522,N_8934);
nor U9110 (N_9110,N_8556,N_8681);
xor U9111 (N_9111,N_8575,N_8521);
nor U9112 (N_9112,N_8516,N_8578);
and U9113 (N_9113,N_8951,N_8695);
xor U9114 (N_9114,N_8591,N_8912);
xor U9115 (N_9115,N_8764,N_8883);
nor U9116 (N_9116,N_8861,N_8735);
xor U9117 (N_9117,N_8503,N_8712);
and U9118 (N_9118,N_8959,N_8706);
xnor U9119 (N_9119,N_8985,N_8904);
and U9120 (N_9120,N_8929,N_8501);
xnor U9121 (N_9121,N_8566,N_8708);
or U9122 (N_9122,N_8707,N_8614);
nor U9123 (N_9123,N_8638,N_8531);
nor U9124 (N_9124,N_8675,N_8838);
nand U9125 (N_9125,N_8537,N_8845);
nand U9126 (N_9126,N_8754,N_8688);
nor U9127 (N_9127,N_8846,N_8952);
or U9128 (N_9128,N_8850,N_8790);
xnor U9129 (N_9129,N_8588,N_8925);
and U9130 (N_9130,N_8881,N_8889);
xnor U9131 (N_9131,N_8813,N_8752);
nand U9132 (N_9132,N_8811,N_8634);
or U9133 (N_9133,N_8716,N_8711);
nor U9134 (N_9134,N_8650,N_8667);
nand U9135 (N_9135,N_8757,N_8867);
nand U9136 (N_9136,N_8720,N_8672);
nor U9137 (N_9137,N_8723,N_8617);
nor U9138 (N_9138,N_8748,N_8662);
xnor U9139 (N_9139,N_8983,N_8962);
nor U9140 (N_9140,N_8769,N_8990);
or U9141 (N_9141,N_8549,N_8528);
and U9142 (N_9142,N_8630,N_8520);
nor U9143 (N_9143,N_8654,N_8569);
nand U9144 (N_9144,N_8639,N_8683);
nand U9145 (N_9145,N_8559,N_8969);
or U9146 (N_9146,N_8527,N_8974);
and U9147 (N_9147,N_8580,N_8771);
or U9148 (N_9148,N_8652,N_8627);
nand U9149 (N_9149,N_8987,N_8507);
or U9150 (N_9150,N_8538,N_8950);
nor U9151 (N_9151,N_8873,N_8866);
nor U9152 (N_9152,N_8705,N_8567);
xor U9153 (N_9153,N_8937,N_8594);
and U9154 (N_9154,N_8581,N_8726);
or U9155 (N_9155,N_8851,N_8600);
nor U9156 (N_9156,N_8562,N_8783);
nand U9157 (N_9157,N_8976,N_8835);
xor U9158 (N_9158,N_8509,N_8791);
nor U9159 (N_9159,N_8956,N_8514);
or U9160 (N_9160,N_8876,N_8984);
nor U9161 (N_9161,N_8958,N_8814);
and U9162 (N_9162,N_8877,N_8645);
xnor U9163 (N_9163,N_8656,N_8740);
or U9164 (N_9164,N_8917,N_8742);
and U9165 (N_9165,N_8560,N_8857);
nand U9166 (N_9166,N_8903,N_8540);
or U9167 (N_9167,N_8863,N_8796);
nor U9168 (N_9168,N_8511,N_8921);
nand U9169 (N_9169,N_8699,N_8653);
nor U9170 (N_9170,N_8777,N_8730);
and U9171 (N_9171,N_8849,N_8603);
xnor U9172 (N_9172,N_8770,N_8568);
and U9173 (N_9173,N_8518,N_8755);
and U9174 (N_9174,N_8862,N_8721);
nor U9175 (N_9175,N_8669,N_8955);
nand U9176 (N_9176,N_8703,N_8637);
xor U9177 (N_9177,N_8636,N_8607);
and U9178 (N_9178,N_8789,N_8916);
or U9179 (N_9179,N_8745,N_8551);
nor U9180 (N_9180,N_8753,N_8853);
nor U9181 (N_9181,N_8943,N_8827);
xnor U9182 (N_9182,N_8670,N_8682);
xnor U9183 (N_9183,N_8882,N_8908);
nor U9184 (N_9184,N_8646,N_8817);
and U9185 (N_9185,N_8772,N_8622);
or U9186 (N_9186,N_8860,N_8927);
nand U9187 (N_9187,N_8515,N_8775);
nand U9188 (N_9188,N_8979,N_8815);
or U9189 (N_9189,N_8579,N_8674);
or U9190 (N_9190,N_8714,N_8596);
and U9191 (N_9191,N_8504,N_8802);
nand U9192 (N_9192,N_8913,N_8963);
and U9193 (N_9193,N_8631,N_8804);
xor U9194 (N_9194,N_8819,N_8701);
or U9195 (N_9195,N_8736,N_8836);
xor U9196 (N_9196,N_8661,N_8558);
nand U9197 (N_9197,N_8810,N_8691);
nand U9198 (N_9198,N_8924,N_8629);
and U9199 (N_9199,N_8932,N_8665);
and U9200 (N_9200,N_8821,N_8524);
and U9201 (N_9201,N_8830,N_8710);
and U9202 (N_9202,N_8898,N_8954);
and U9203 (N_9203,N_8868,N_8928);
and U9204 (N_9204,N_8564,N_8978);
and U9205 (N_9205,N_8734,N_8611);
or U9206 (N_9206,N_8536,N_8870);
nor U9207 (N_9207,N_8620,N_8583);
nor U9208 (N_9208,N_8679,N_8901);
or U9209 (N_9209,N_8738,N_8743);
nor U9210 (N_9210,N_8942,N_8666);
nand U9211 (N_9211,N_8875,N_8906);
xnor U9212 (N_9212,N_8886,N_8737);
and U9213 (N_9213,N_8993,N_8773);
xnor U9214 (N_9214,N_8892,N_8825);
or U9215 (N_9215,N_8632,N_8878);
xnor U9216 (N_9216,N_8947,N_8673);
nor U9217 (N_9217,N_8988,N_8529);
nor U9218 (N_9218,N_8895,N_8848);
xor U9219 (N_9219,N_8592,N_8837);
nand U9220 (N_9220,N_8732,N_8649);
or U9221 (N_9221,N_8621,N_8809);
or U9222 (N_9222,N_8767,N_8548);
nor U9223 (N_9223,N_8539,N_8613);
and U9224 (N_9224,N_8554,N_8590);
and U9225 (N_9225,N_8788,N_8648);
and U9226 (N_9226,N_8727,N_8829);
xnor U9227 (N_9227,N_8693,N_8713);
nor U9228 (N_9228,N_8689,N_8779);
and U9229 (N_9229,N_8698,N_8553);
or U9230 (N_9230,N_8909,N_8543);
nor U9231 (N_9231,N_8818,N_8519);
nor U9232 (N_9232,N_8968,N_8899);
nand U9233 (N_9233,N_8926,N_8971);
nand U9234 (N_9234,N_8660,N_8785);
xor U9235 (N_9235,N_8806,N_8502);
nand U9236 (N_9236,N_8640,N_8831);
and U9237 (N_9237,N_8597,N_8542);
nor U9238 (N_9238,N_8905,N_8842);
nor U9239 (N_9239,N_8872,N_8975);
xor U9240 (N_9240,N_8604,N_8605);
nand U9241 (N_9241,N_8641,N_8655);
xnor U9242 (N_9242,N_8801,N_8793);
nor U9243 (N_9243,N_8961,N_8715);
nor U9244 (N_9244,N_8651,N_8719);
nand U9245 (N_9245,N_8972,N_8545);
and U9246 (N_9246,N_8865,N_8936);
nor U9247 (N_9247,N_8618,N_8918);
and U9248 (N_9248,N_8869,N_8995);
nand U9249 (N_9249,N_8510,N_8980);
xnor U9250 (N_9250,N_8930,N_8553);
nor U9251 (N_9251,N_8797,N_8921);
or U9252 (N_9252,N_8694,N_8920);
xor U9253 (N_9253,N_8744,N_8964);
nor U9254 (N_9254,N_8865,N_8537);
nand U9255 (N_9255,N_8511,N_8819);
xnor U9256 (N_9256,N_8637,N_8604);
nor U9257 (N_9257,N_8612,N_8684);
and U9258 (N_9258,N_8646,N_8728);
xor U9259 (N_9259,N_8991,N_8872);
and U9260 (N_9260,N_8959,N_8514);
and U9261 (N_9261,N_8620,N_8997);
and U9262 (N_9262,N_8808,N_8508);
xnor U9263 (N_9263,N_8630,N_8724);
xor U9264 (N_9264,N_8568,N_8791);
xnor U9265 (N_9265,N_8641,N_8575);
nor U9266 (N_9266,N_8823,N_8508);
nor U9267 (N_9267,N_8776,N_8883);
xnor U9268 (N_9268,N_8675,N_8855);
nor U9269 (N_9269,N_8608,N_8741);
and U9270 (N_9270,N_8795,N_8563);
xor U9271 (N_9271,N_8623,N_8763);
nand U9272 (N_9272,N_8856,N_8882);
or U9273 (N_9273,N_8732,N_8509);
nor U9274 (N_9274,N_8685,N_8979);
and U9275 (N_9275,N_8997,N_8667);
nor U9276 (N_9276,N_8592,N_8540);
nand U9277 (N_9277,N_8753,N_8977);
or U9278 (N_9278,N_8940,N_8647);
xor U9279 (N_9279,N_8769,N_8741);
nand U9280 (N_9280,N_8603,N_8758);
xnor U9281 (N_9281,N_8615,N_8838);
nor U9282 (N_9282,N_8927,N_8544);
or U9283 (N_9283,N_8534,N_8712);
xnor U9284 (N_9284,N_8577,N_8591);
and U9285 (N_9285,N_8724,N_8864);
xnor U9286 (N_9286,N_8979,N_8948);
and U9287 (N_9287,N_8500,N_8763);
nand U9288 (N_9288,N_8621,N_8595);
xnor U9289 (N_9289,N_8562,N_8688);
nand U9290 (N_9290,N_8905,N_8966);
or U9291 (N_9291,N_8945,N_8816);
nand U9292 (N_9292,N_8866,N_8728);
nand U9293 (N_9293,N_8540,N_8714);
and U9294 (N_9294,N_8586,N_8538);
and U9295 (N_9295,N_8822,N_8747);
or U9296 (N_9296,N_8786,N_8917);
or U9297 (N_9297,N_8610,N_8795);
or U9298 (N_9298,N_8898,N_8972);
nor U9299 (N_9299,N_8946,N_8632);
or U9300 (N_9300,N_8716,N_8975);
nor U9301 (N_9301,N_8625,N_8735);
xnor U9302 (N_9302,N_8663,N_8832);
nand U9303 (N_9303,N_8784,N_8656);
nand U9304 (N_9304,N_8531,N_8622);
nor U9305 (N_9305,N_8674,N_8886);
nor U9306 (N_9306,N_8921,N_8851);
or U9307 (N_9307,N_8903,N_8860);
nand U9308 (N_9308,N_8698,N_8603);
xnor U9309 (N_9309,N_8577,N_8617);
nand U9310 (N_9310,N_8838,N_8823);
xor U9311 (N_9311,N_8676,N_8563);
nand U9312 (N_9312,N_8895,N_8723);
and U9313 (N_9313,N_8535,N_8748);
or U9314 (N_9314,N_8556,N_8851);
nand U9315 (N_9315,N_8707,N_8598);
or U9316 (N_9316,N_8745,N_8722);
nand U9317 (N_9317,N_8712,N_8664);
xor U9318 (N_9318,N_8645,N_8620);
and U9319 (N_9319,N_8502,N_8855);
xnor U9320 (N_9320,N_8894,N_8920);
nand U9321 (N_9321,N_8970,N_8961);
nand U9322 (N_9322,N_8807,N_8949);
and U9323 (N_9323,N_8851,N_8615);
xnor U9324 (N_9324,N_8570,N_8709);
nor U9325 (N_9325,N_8543,N_8922);
and U9326 (N_9326,N_8533,N_8625);
nand U9327 (N_9327,N_8587,N_8771);
xnor U9328 (N_9328,N_8999,N_8824);
nand U9329 (N_9329,N_8660,N_8688);
nor U9330 (N_9330,N_8558,N_8507);
nor U9331 (N_9331,N_8541,N_8845);
nand U9332 (N_9332,N_8690,N_8836);
xor U9333 (N_9333,N_8511,N_8717);
nor U9334 (N_9334,N_8618,N_8901);
or U9335 (N_9335,N_8657,N_8546);
nand U9336 (N_9336,N_8500,N_8621);
nor U9337 (N_9337,N_8947,N_8816);
nand U9338 (N_9338,N_8781,N_8667);
xnor U9339 (N_9339,N_8689,N_8667);
nor U9340 (N_9340,N_8510,N_8534);
and U9341 (N_9341,N_8793,N_8876);
nor U9342 (N_9342,N_8920,N_8816);
or U9343 (N_9343,N_8970,N_8753);
or U9344 (N_9344,N_8563,N_8883);
xor U9345 (N_9345,N_8619,N_8636);
nor U9346 (N_9346,N_8957,N_8566);
or U9347 (N_9347,N_8551,N_8579);
and U9348 (N_9348,N_8841,N_8570);
nor U9349 (N_9349,N_8931,N_8560);
nand U9350 (N_9350,N_8691,N_8942);
xor U9351 (N_9351,N_8731,N_8876);
nor U9352 (N_9352,N_8809,N_8514);
or U9353 (N_9353,N_8905,N_8702);
and U9354 (N_9354,N_8648,N_8645);
nor U9355 (N_9355,N_8627,N_8651);
and U9356 (N_9356,N_8963,N_8655);
and U9357 (N_9357,N_8589,N_8728);
nand U9358 (N_9358,N_8916,N_8787);
xor U9359 (N_9359,N_8673,N_8990);
xnor U9360 (N_9360,N_8674,N_8572);
xnor U9361 (N_9361,N_8685,N_8975);
xor U9362 (N_9362,N_8848,N_8779);
nand U9363 (N_9363,N_8821,N_8981);
or U9364 (N_9364,N_8635,N_8836);
and U9365 (N_9365,N_8904,N_8816);
and U9366 (N_9366,N_8767,N_8664);
nand U9367 (N_9367,N_8832,N_8919);
nand U9368 (N_9368,N_8538,N_8655);
and U9369 (N_9369,N_8905,N_8990);
nor U9370 (N_9370,N_8519,N_8684);
or U9371 (N_9371,N_8968,N_8737);
xnor U9372 (N_9372,N_8591,N_8998);
nand U9373 (N_9373,N_8935,N_8933);
or U9374 (N_9374,N_8608,N_8916);
and U9375 (N_9375,N_8857,N_8582);
nand U9376 (N_9376,N_8763,N_8942);
nor U9377 (N_9377,N_8645,N_8883);
nor U9378 (N_9378,N_8714,N_8622);
nand U9379 (N_9379,N_8810,N_8757);
nand U9380 (N_9380,N_8818,N_8812);
nor U9381 (N_9381,N_8959,N_8881);
nand U9382 (N_9382,N_8694,N_8735);
xor U9383 (N_9383,N_8577,N_8550);
nor U9384 (N_9384,N_8597,N_8630);
or U9385 (N_9385,N_8552,N_8660);
nand U9386 (N_9386,N_8881,N_8636);
and U9387 (N_9387,N_8556,N_8775);
nand U9388 (N_9388,N_8528,N_8601);
or U9389 (N_9389,N_8945,N_8601);
nand U9390 (N_9390,N_8967,N_8615);
and U9391 (N_9391,N_8767,N_8959);
nor U9392 (N_9392,N_8979,N_8535);
and U9393 (N_9393,N_8907,N_8641);
or U9394 (N_9394,N_8839,N_8748);
and U9395 (N_9395,N_8891,N_8540);
nor U9396 (N_9396,N_8665,N_8578);
nor U9397 (N_9397,N_8965,N_8862);
nor U9398 (N_9398,N_8617,N_8555);
or U9399 (N_9399,N_8546,N_8979);
nand U9400 (N_9400,N_8725,N_8551);
xor U9401 (N_9401,N_8831,N_8902);
or U9402 (N_9402,N_8875,N_8670);
nor U9403 (N_9403,N_8611,N_8833);
xor U9404 (N_9404,N_8864,N_8853);
xnor U9405 (N_9405,N_8507,N_8585);
nand U9406 (N_9406,N_8613,N_8611);
xor U9407 (N_9407,N_8907,N_8521);
nand U9408 (N_9408,N_8959,N_8701);
and U9409 (N_9409,N_8701,N_8743);
nor U9410 (N_9410,N_8647,N_8689);
xnor U9411 (N_9411,N_8578,N_8742);
nand U9412 (N_9412,N_8862,N_8593);
and U9413 (N_9413,N_8588,N_8915);
nand U9414 (N_9414,N_8811,N_8504);
xor U9415 (N_9415,N_8507,N_8736);
nand U9416 (N_9416,N_8869,N_8689);
and U9417 (N_9417,N_8899,N_8825);
nand U9418 (N_9418,N_8694,N_8764);
nand U9419 (N_9419,N_8808,N_8750);
nand U9420 (N_9420,N_8942,N_8644);
nor U9421 (N_9421,N_8856,N_8771);
xor U9422 (N_9422,N_8594,N_8902);
nor U9423 (N_9423,N_8758,N_8685);
xnor U9424 (N_9424,N_8712,N_8873);
or U9425 (N_9425,N_8832,N_8837);
xnor U9426 (N_9426,N_8560,N_8584);
xnor U9427 (N_9427,N_8566,N_8960);
or U9428 (N_9428,N_8661,N_8897);
or U9429 (N_9429,N_8861,N_8536);
and U9430 (N_9430,N_8732,N_8739);
or U9431 (N_9431,N_8789,N_8585);
xnor U9432 (N_9432,N_8667,N_8564);
nor U9433 (N_9433,N_8880,N_8616);
nor U9434 (N_9434,N_8877,N_8758);
and U9435 (N_9435,N_8929,N_8989);
and U9436 (N_9436,N_8869,N_8755);
nand U9437 (N_9437,N_8994,N_8703);
xnor U9438 (N_9438,N_8599,N_8643);
nand U9439 (N_9439,N_8503,N_8697);
and U9440 (N_9440,N_8809,N_8958);
or U9441 (N_9441,N_8501,N_8727);
or U9442 (N_9442,N_8809,N_8703);
or U9443 (N_9443,N_8982,N_8601);
and U9444 (N_9444,N_8983,N_8706);
or U9445 (N_9445,N_8794,N_8600);
and U9446 (N_9446,N_8542,N_8956);
or U9447 (N_9447,N_8929,N_8857);
nand U9448 (N_9448,N_8572,N_8511);
nor U9449 (N_9449,N_8943,N_8779);
nand U9450 (N_9450,N_8662,N_8881);
xnor U9451 (N_9451,N_8729,N_8845);
nor U9452 (N_9452,N_8696,N_8876);
nand U9453 (N_9453,N_8936,N_8904);
or U9454 (N_9454,N_8781,N_8595);
nand U9455 (N_9455,N_8807,N_8758);
and U9456 (N_9456,N_8927,N_8762);
nor U9457 (N_9457,N_8747,N_8873);
or U9458 (N_9458,N_8802,N_8924);
or U9459 (N_9459,N_8557,N_8867);
nor U9460 (N_9460,N_8535,N_8864);
nand U9461 (N_9461,N_8600,N_8943);
nor U9462 (N_9462,N_8767,N_8807);
or U9463 (N_9463,N_8747,N_8686);
nand U9464 (N_9464,N_8938,N_8949);
and U9465 (N_9465,N_8996,N_8673);
or U9466 (N_9466,N_8633,N_8578);
or U9467 (N_9467,N_8529,N_8722);
and U9468 (N_9468,N_8519,N_8975);
nand U9469 (N_9469,N_8501,N_8933);
xnor U9470 (N_9470,N_8981,N_8760);
and U9471 (N_9471,N_8924,N_8509);
nand U9472 (N_9472,N_8714,N_8796);
xnor U9473 (N_9473,N_8796,N_8527);
and U9474 (N_9474,N_8864,N_8741);
and U9475 (N_9475,N_8594,N_8528);
and U9476 (N_9476,N_8572,N_8995);
or U9477 (N_9477,N_8789,N_8669);
xor U9478 (N_9478,N_8925,N_8641);
and U9479 (N_9479,N_8781,N_8577);
and U9480 (N_9480,N_8914,N_8775);
nand U9481 (N_9481,N_8754,N_8681);
and U9482 (N_9482,N_8667,N_8646);
nand U9483 (N_9483,N_8884,N_8692);
nor U9484 (N_9484,N_8643,N_8882);
nor U9485 (N_9485,N_8533,N_8857);
and U9486 (N_9486,N_8631,N_8829);
and U9487 (N_9487,N_8734,N_8952);
or U9488 (N_9488,N_8689,N_8614);
xnor U9489 (N_9489,N_8555,N_8525);
and U9490 (N_9490,N_8957,N_8664);
xnor U9491 (N_9491,N_8573,N_8835);
nor U9492 (N_9492,N_8717,N_8631);
xnor U9493 (N_9493,N_8893,N_8775);
xor U9494 (N_9494,N_8683,N_8679);
xnor U9495 (N_9495,N_8518,N_8564);
and U9496 (N_9496,N_8811,N_8676);
or U9497 (N_9497,N_8746,N_8983);
xnor U9498 (N_9498,N_8652,N_8590);
nor U9499 (N_9499,N_8904,N_8879);
xnor U9500 (N_9500,N_9077,N_9052);
nand U9501 (N_9501,N_9314,N_9169);
xor U9502 (N_9502,N_9000,N_9460);
xnor U9503 (N_9503,N_9458,N_9206);
or U9504 (N_9504,N_9049,N_9115);
xnor U9505 (N_9505,N_9465,N_9236);
and U9506 (N_9506,N_9081,N_9132);
xor U9507 (N_9507,N_9209,N_9357);
and U9508 (N_9508,N_9348,N_9406);
and U9509 (N_9509,N_9280,N_9420);
and U9510 (N_9510,N_9198,N_9494);
xnor U9511 (N_9511,N_9144,N_9341);
or U9512 (N_9512,N_9190,N_9479);
nand U9513 (N_9513,N_9445,N_9367);
and U9514 (N_9514,N_9120,N_9374);
or U9515 (N_9515,N_9402,N_9204);
xor U9516 (N_9516,N_9271,N_9355);
and U9517 (N_9517,N_9097,N_9295);
xnor U9518 (N_9518,N_9189,N_9369);
or U9519 (N_9519,N_9118,N_9105);
nand U9520 (N_9520,N_9281,N_9087);
nor U9521 (N_9521,N_9304,N_9139);
nor U9522 (N_9522,N_9387,N_9110);
or U9523 (N_9523,N_9074,N_9421);
nand U9524 (N_9524,N_9359,N_9409);
or U9525 (N_9525,N_9286,N_9478);
and U9526 (N_9526,N_9142,N_9436);
nor U9527 (N_9527,N_9243,N_9317);
and U9528 (N_9528,N_9426,N_9256);
or U9529 (N_9529,N_9145,N_9037);
and U9530 (N_9530,N_9311,N_9340);
and U9531 (N_9531,N_9213,N_9193);
or U9532 (N_9532,N_9123,N_9318);
xor U9533 (N_9533,N_9017,N_9122);
and U9534 (N_9534,N_9399,N_9060);
and U9535 (N_9535,N_9214,N_9151);
or U9536 (N_9536,N_9331,N_9245);
and U9537 (N_9537,N_9362,N_9027);
or U9538 (N_9538,N_9287,N_9444);
or U9539 (N_9539,N_9156,N_9497);
and U9540 (N_9540,N_9099,N_9158);
xnor U9541 (N_9541,N_9411,N_9002);
and U9542 (N_9542,N_9024,N_9152);
and U9543 (N_9543,N_9408,N_9289);
or U9544 (N_9544,N_9384,N_9454);
nand U9545 (N_9545,N_9372,N_9263);
nor U9546 (N_9546,N_9136,N_9038);
xnor U9547 (N_9547,N_9045,N_9053);
nor U9548 (N_9548,N_9373,N_9016);
and U9549 (N_9549,N_9013,N_9095);
and U9550 (N_9550,N_9473,N_9019);
nor U9551 (N_9551,N_9004,N_9199);
or U9552 (N_9552,N_9468,N_9201);
xnor U9553 (N_9553,N_9227,N_9325);
nand U9554 (N_9554,N_9288,N_9031);
or U9555 (N_9555,N_9065,N_9160);
nand U9556 (N_9556,N_9101,N_9447);
nor U9557 (N_9557,N_9219,N_9350);
nand U9558 (N_9558,N_9187,N_9223);
and U9559 (N_9559,N_9055,N_9003);
nor U9560 (N_9560,N_9252,N_9010);
nor U9561 (N_9561,N_9018,N_9246);
xor U9562 (N_9562,N_9107,N_9057);
xor U9563 (N_9563,N_9435,N_9329);
nand U9564 (N_9564,N_9062,N_9481);
nor U9565 (N_9565,N_9143,N_9486);
or U9566 (N_9566,N_9240,N_9459);
xor U9567 (N_9567,N_9165,N_9407);
nor U9568 (N_9568,N_9381,N_9197);
nand U9569 (N_9569,N_9174,N_9114);
and U9570 (N_9570,N_9309,N_9100);
nor U9571 (N_9571,N_9021,N_9098);
nor U9572 (N_9572,N_9302,N_9225);
nand U9573 (N_9573,N_9112,N_9360);
nor U9574 (N_9574,N_9490,N_9443);
nand U9575 (N_9575,N_9092,N_9231);
xor U9576 (N_9576,N_9424,N_9290);
nand U9577 (N_9577,N_9033,N_9358);
xnor U9578 (N_9578,N_9433,N_9398);
or U9579 (N_9579,N_9361,N_9244);
or U9580 (N_9580,N_9255,N_9432);
nand U9581 (N_9581,N_9242,N_9086);
xor U9582 (N_9582,N_9161,N_9438);
and U9583 (N_9583,N_9078,N_9119);
nand U9584 (N_9584,N_9025,N_9232);
xor U9585 (N_9585,N_9430,N_9066);
and U9586 (N_9586,N_9036,N_9182);
and U9587 (N_9587,N_9382,N_9059);
nor U9588 (N_9588,N_9186,N_9166);
and U9589 (N_9589,N_9267,N_9346);
xor U9590 (N_9590,N_9032,N_9293);
and U9591 (N_9591,N_9285,N_9393);
xor U9592 (N_9592,N_9268,N_9073);
nor U9593 (N_9593,N_9154,N_9009);
nand U9594 (N_9594,N_9487,N_9451);
nand U9595 (N_9595,N_9212,N_9303);
nand U9596 (N_9596,N_9217,N_9224);
or U9597 (N_9597,N_9334,N_9397);
xnor U9598 (N_9598,N_9104,N_9416);
xor U9599 (N_9599,N_9046,N_9134);
xor U9600 (N_9600,N_9040,N_9183);
nor U9601 (N_9601,N_9493,N_9264);
nor U9602 (N_9602,N_9258,N_9185);
or U9603 (N_9603,N_9248,N_9272);
and U9604 (N_9604,N_9047,N_9167);
nand U9605 (N_9605,N_9457,N_9129);
xor U9606 (N_9606,N_9425,N_9137);
and U9607 (N_9607,N_9423,N_9043);
xor U9608 (N_9608,N_9323,N_9389);
or U9609 (N_9609,N_9277,N_9220);
nand U9610 (N_9610,N_9403,N_9450);
xnor U9611 (N_9611,N_9306,N_9313);
nor U9612 (N_9612,N_9237,N_9241);
or U9613 (N_9613,N_9216,N_9273);
and U9614 (N_9614,N_9181,N_9064);
nor U9615 (N_9615,N_9157,N_9483);
xnor U9616 (N_9616,N_9184,N_9117);
xor U9617 (N_9617,N_9370,N_9482);
xor U9618 (N_9618,N_9188,N_9298);
or U9619 (N_9619,N_9054,N_9067);
and U9620 (N_9620,N_9251,N_9279);
xnor U9621 (N_9621,N_9068,N_9449);
or U9622 (N_9622,N_9001,N_9475);
nor U9623 (N_9623,N_9322,N_9442);
and U9624 (N_9624,N_9324,N_9395);
nor U9625 (N_9625,N_9363,N_9096);
xor U9626 (N_9626,N_9210,N_9337);
or U9627 (N_9627,N_9491,N_9386);
and U9628 (N_9628,N_9388,N_9326);
or U9629 (N_9629,N_9401,N_9297);
and U9630 (N_9630,N_9283,N_9422);
xnor U9631 (N_9631,N_9321,N_9146);
nand U9632 (N_9632,N_9495,N_9261);
xnor U9633 (N_9633,N_9332,N_9180);
nand U9634 (N_9634,N_9392,N_9028);
nand U9635 (N_9635,N_9130,N_9070);
and U9636 (N_9636,N_9274,N_9441);
xnor U9637 (N_9637,N_9396,N_9138);
xnor U9638 (N_9638,N_9415,N_9315);
or U9639 (N_9639,N_9404,N_9368);
and U9640 (N_9640,N_9075,N_9345);
or U9641 (N_9641,N_9434,N_9480);
nand U9642 (N_9642,N_9365,N_9235);
and U9643 (N_9643,N_9414,N_9194);
or U9644 (N_9644,N_9125,N_9464);
nor U9645 (N_9645,N_9470,N_9039);
nor U9646 (N_9646,N_9292,N_9347);
nand U9647 (N_9647,N_9353,N_9485);
nand U9648 (N_9648,N_9191,N_9305);
or U9649 (N_9649,N_9342,N_9394);
or U9650 (N_9650,N_9147,N_9429);
or U9651 (N_9651,N_9207,N_9333);
and U9652 (N_9652,N_9462,N_9192);
and U9653 (N_9653,N_9455,N_9140);
xor U9654 (N_9654,N_9354,N_9291);
nor U9655 (N_9655,N_9103,N_9083);
nand U9656 (N_9656,N_9308,N_9312);
nand U9657 (N_9657,N_9093,N_9205);
nand U9658 (N_9658,N_9089,N_9133);
and U9659 (N_9659,N_9418,N_9344);
nand U9660 (N_9660,N_9044,N_9176);
and U9661 (N_9661,N_9048,N_9319);
and U9662 (N_9662,N_9106,N_9006);
xor U9663 (N_9663,N_9484,N_9200);
and U9664 (N_9664,N_9474,N_9400);
nor U9665 (N_9665,N_9034,N_9278);
xnor U9666 (N_9666,N_9330,N_9069);
and U9667 (N_9667,N_9247,N_9061);
xor U9668 (N_9668,N_9159,N_9179);
or U9669 (N_9669,N_9467,N_9379);
or U9670 (N_9670,N_9296,N_9164);
and U9671 (N_9671,N_9440,N_9020);
nand U9672 (N_9672,N_9356,N_9488);
nor U9673 (N_9673,N_9076,N_9383);
or U9674 (N_9674,N_9352,N_9111);
nand U9675 (N_9675,N_9471,N_9090);
xnor U9676 (N_9676,N_9253,N_9472);
xor U9677 (N_9677,N_9489,N_9014);
and U9678 (N_9678,N_9327,N_9377);
nor U9679 (N_9679,N_9022,N_9109);
nand U9680 (N_9680,N_9476,N_9371);
xnor U9681 (N_9681,N_9222,N_9349);
xor U9682 (N_9682,N_9084,N_9072);
and U9683 (N_9683,N_9127,N_9128);
xnor U9684 (N_9684,N_9265,N_9226);
nor U9685 (N_9685,N_9300,N_9203);
xnor U9686 (N_9686,N_9177,N_9051);
and U9687 (N_9687,N_9294,N_9148);
xor U9688 (N_9688,N_9269,N_9262);
xnor U9689 (N_9689,N_9239,N_9376);
or U9690 (N_9690,N_9266,N_9080);
nor U9691 (N_9691,N_9439,N_9260);
and U9692 (N_9692,N_9116,N_9390);
xnor U9693 (N_9693,N_9463,N_9230);
and U9694 (N_9694,N_9050,N_9058);
xnor U9695 (N_9695,N_9088,N_9108);
nor U9696 (N_9696,N_9015,N_9008);
and U9697 (N_9697,N_9320,N_9082);
nand U9698 (N_9698,N_9419,N_9316);
nor U9699 (N_9699,N_9063,N_9113);
nand U9700 (N_9700,N_9035,N_9446);
xor U9701 (N_9701,N_9466,N_9498);
nor U9702 (N_9702,N_9085,N_9155);
or U9703 (N_9703,N_9171,N_9131);
nand U9704 (N_9704,N_9417,N_9456);
and U9705 (N_9705,N_9173,N_9041);
nor U9706 (N_9706,N_9307,N_9238);
xnor U9707 (N_9707,N_9150,N_9195);
nand U9708 (N_9708,N_9276,N_9405);
or U9709 (N_9709,N_9079,N_9135);
or U9710 (N_9710,N_9328,N_9410);
and U9711 (N_9711,N_9221,N_9228);
or U9712 (N_9712,N_9141,N_9094);
nor U9713 (N_9713,N_9366,N_9124);
xnor U9714 (N_9714,N_9452,N_9023);
nor U9715 (N_9715,N_9208,N_9499);
xor U9716 (N_9716,N_9437,N_9153);
and U9717 (N_9717,N_9310,N_9102);
xnor U9718 (N_9718,N_9428,N_9121);
xor U9719 (N_9719,N_9364,N_9071);
nor U9720 (N_9720,N_9351,N_9202);
and U9721 (N_9721,N_9229,N_9233);
nor U9722 (N_9722,N_9492,N_9335);
xor U9723 (N_9723,N_9211,N_9427);
xor U9724 (N_9724,N_9282,N_9042);
or U9725 (N_9725,N_9234,N_9284);
and U9726 (N_9726,N_9336,N_9343);
nor U9727 (N_9727,N_9030,N_9196);
or U9728 (N_9728,N_9162,N_9380);
or U9729 (N_9729,N_9218,N_9496);
nand U9730 (N_9730,N_9375,N_9170);
nand U9731 (N_9731,N_9215,N_9453);
xnor U9732 (N_9732,N_9178,N_9026);
nor U9733 (N_9733,N_9338,N_9012);
xnor U9734 (N_9734,N_9275,N_9469);
nor U9735 (N_9735,N_9011,N_9029);
nor U9736 (N_9736,N_9091,N_9259);
xor U9737 (N_9737,N_9299,N_9448);
nand U9738 (N_9738,N_9257,N_9301);
nand U9739 (N_9739,N_9413,N_9126);
nor U9740 (N_9740,N_9391,N_9149);
and U9741 (N_9741,N_9385,N_9378);
or U9742 (N_9742,N_9168,N_9412);
nand U9743 (N_9743,N_9007,N_9172);
or U9744 (N_9744,N_9163,N_9477);
nor U9745 (N_9745,N_9431,N_9339);
xnor U9746 (N_9746,N_9461,N_9056);
and U9747 (N_9747,N_9250,N_9249);
and U9748 (N_9748,N_9005,N_9270);
or U9749 (N_9749,N_9175,N_9254);
or U9750 (N_9750,N_9419,N_9052);
xor U9751 (N_9751,N_9111,N_9118);
or U9752 (N_9752,N_9106,N_9157);
nand U9753 (N_9753,N_9422,N_9159);
and U9754 (N_9754,N_9203,N_9162);
and U9755 (N_9755,N_9416,N_9209);
and U9756 (N_9756,N_9408,N_9001);
nand U9757 (N_9757,N_9210,N_9412);
or U9758 (N_9758,N_9109,N_9488);
xnor U9759 (N_9759,N_9181,N_9213);
xnor U9760 (N_9760,N_9077,N_9178);
nand U9761 (N_9761,N_9060,N_9214);
xnor U9762 (N_9762,N_9413,N_9081);
and U9763 (N_9763,N_9205,N_9005);
nor U9764 (N_9764,N_9385,N_9402);
xor U9765 (N_9765,N_9023,N_9052);
or U9766 (N_9766,N_9322,N_9427);
nand U9767 (N_9767,N_9277,N_9299);
xor U9768 (N_9768,N_9008,N_9101);
nor U9769 (N_9769,N_9315,N_9459);
nand U9770 (N_9770,N_9372,N_9115);
nor U9771 (N_9771,N_9287,N_9183);
nand U9772 (N_9772,N_9296,N_9150);
and U9773 (N_9773,N_9445,N_9063);
nor U9774 (N_9774,N_9108,N_9466);
nor U9775 (N_9775,N_9326,N_9176);
and U9776 (N_9776,N_9484,N_9298);
and U9777 (N_9777,N_9347,N_9221);
xor U9778 (N_9778,N_9141,N_9309);
nand U9779 (N_9779,N_9434,N_9181);
and U9780 (N_9780,N_9222,N_9480);
or U9781 (N_9781,N_9319,N_9328);
and U9782 (N_9782,N_9269,N_9226);
nor U9783 (N_9783,N_9125,N_9018);
or U9784 (N_9784,N_9459,N_9231);
nand U9785 (N_9785,N_9131,N_9070);
and U9786 (N_9786,N_9160,N_9207);
nand U9787 (N_9787,N_9116,N_9144);
and U9788 (N_9788,N_9101,N_9286);
or U9789 (N_9789,N_9193,N_9055);
nor U9790 (N_9790,N_9003,N_9238);
or U9791 (N_9791,N_9029,N_9019);
or U9792 (N_9792,N_9130,N_9076);
nor U9793 (N_9793,N_9028,N_9197);
nor U9794 (N_9794,N_9335,N_9029);
nand U9795 (N_9795,N_9106,N_9306);
nor U9796 (N_9796,N_9200,N_9079);
and U9797 (N_9797,N_9349,N_9327);
or U9798 (N_9798,N_9247,N_9187);
nand U9799 (N_9799,N_9087,N_9304);
xor U9800 (N_9800,N_9186,N_9323);
and U9801 (N_9801,N_9491,N_9314);
nand U9802 (N_9802,N_9043,N_9421);
nor U9803 (N_9803,N_9008,N_9007);
nand U9804 (N_9804,N_9443,N_9242);
or U9805 (N_9805,N_9109,N_9025);
and U9806 (N_9806,N_9306,N_9022);
nor U9807 (N_9807,N_9365,N_9273);
nor U9808 (N_9808,N_9263,N_9254);
xnor U9809 (N_9809,N_9235,N_9155);
xnor U9810 (N_9810,N_9128,N_9324);
or U9811 (N_9811,N_9465,N_9401);
xor U9812 (N_9812,N_9483,N_9289);
nor U9813 (N_9813,N_9449,N_9431);
xnor U9814 (N_9814,N_9209,N_9220);
or U9815 (N_9815,N_9110,N_9389);
and U9816 (N_9816,N_9472,N_9343);
nand U9817 (N_9817,N_9421,N_9231);
nor U9818 (N_9818,N_9157,N_9320);
and U9819 (N_9819,N_9441,N_9352);
nor U9820 (N_9820,N_9440,N_9327);
or U9821 (N_9821,N_9293,N_9406);
xor U9822 (N_9822,N_9360,N_9319);
nand U9823 (N_9823,N_9392,N_9147);
nor U9824 (N_9824,N_9395,N_9106);
and U9825 (N_9825,N_9135,N_9455);
or U9826 (N_9826,N_9059,N_9435);
nor U9827 (N_9827,N_9035,N_9168);
nor U9828 (N_9828,N_9200,N_9227);
and U9829 (N_9829,N_9037,N_9245);
nand U9830 (N_9830,N_9218,N_9008);
nor U9831 (N_9831,N_9163,N_9440);
nor U9832 (N_9832,N_9090,N_9302);
nand U9833 (N_9833,N_9421,N_9405);
nor U9834 (N_9834,N_9092,N_9371);
or U9835 (N_9835,N_9340,N_9076);
or U9836 (N_9836,N_9110,N_9014);
nor U9837 (N_9837,N_9126,N_9216);
nand U9838 (N_9838,N_9134,N_9463);
xor U9839 (N_9839,N_9242,N_9121);
and U9840 (N_9840,N_9024,N_9253);
nand U9841 (N_9841,N_9302,N_9411);
xor U9842 (N_9842,N_9148,N_9494);
nor U9843 (N_9843,N_9308,N_9007);
nand U9844 (N_9844,N_9003,N_9464);
nor U9845 (N_9845,N_9137,N_9405);
xnor U9846 (N_9846,N_9326,N_9158);
nand U9847 (N_9847,N_9490,N_9060);
nand U9848 (N_9848,N_9183,N_9293);
xnor U9849 (N_9849,N_9339,N_9372);
xor U9850 (N_9850,N_9375,N_9162);
nand U9851 (N_9851,N_9455,N_9214);
nor U9852 (N_9852,N_9003,N_9186);
xnor U9853 (N_9853,N_9464,N_9067);
nand U9854 (N_9854,N_9181,N_9406);
or U9855 (N_9855,N_9140,N_9227);
nand U9856 (N_9856,N_9401,N_9014);
and U9857 (N_9857,N_9116,N_9457);
nor U9858 (N_9858,N_9265,N_9051);
or U9859 (N_9859,N_9345,N_9338);
nand U9860 (N_9860,N_9079,N_9112);
xor U9861 (N_9861,N_9282,N_9219);
nand U9862 (N_9862,N_9206,N_9343);
xor U9863 (N_9863,N_9135,N_9289);
nand U9864 (N_9864,N_9391,N_9089);
or U9865 (N_9865,N_9285,N_9127);
and U9866 (N_9866,N_9386,N_9107);
nand U9867 (N_9867,N_9037,N_9271);
or U9868 (N_9868,N_9111,N_9309);
nor U9869 (N_9869,N_9091,N_9097);
nand U9870 (N_9870,N_9102,N_9034);
and U9871 (N_9871,N_9481,N_9101);
and U9872 (N_9872,N_9203,N_9158);
xor U9873 (N_9873,N_9228,N_9337);
nand U9874 (N_9874,N_9470,N_9418);
nand U9875 (N_9875,N_9216,N_9240);
xor U9876 (N_9876,N_9483,N_9478);
or U9877 (N_9877,N_9024,N_9317);
xor U9878 (N_9878,N_9177,N_9013);
nand U9879 (N_9879,N_9282,N_9487);
xnor U9880 (N_9880,N_9420,N_9410);
or U9881 (N_9881,N_9498,N_9419);
xnor U9882 (N_9882,N_9134,N_9036);
xor U9883 (N_9883,N_9033,N_9318);
and U9884 (N_9884,N_9295,N_9223);
or U9885 (N_9885,N_9474,N_9154);
and U9886 (N_9886,N_9464,N_9045);
xnor U9887 (N_9887,N_9060,N_9165);
nor U9888 (N_9888,N_9493,N_9077);
xor U9889 (N_9889,N_9473,N_9305);
nand U9890 (N_9890,N_9126,N_9335);
or U9891 (N_9891,N_9084,N_9479);
or U9892 (N_9892,N_9122,N_9205);
nor U9893 (N_9893,N_9117,N_9211);
and U9894 (N_9894,N_9195,N_9146);
nor U9895 (N_9895,N_9227,N_9275);
and U9896 (N_9896,N_9308,N_9327);
or U9897 (N_9897,N_9412,N_9131);
nor U9898 (N_9898,N_9290,N_9054);
or U9899 (N_9899,N_9120,N_9329);
nand U9900 (N_9900,N_9322,N_9104);
nand U9901 (N_9901,N_9299,N_9357);
nor U9902 (N_9902,N_9120,N_9311);
or U9903 (N_9903,N_9200,N_9289);
nand U9904 (N_9904,N_9026,N_9261);
nand U9905 (N_9905,N_9128,N_9100);
or U9906 (N_9906,N_9019,N_9011);
xnor U9907 (N_9907,N_9025,N_9304);
and U9908 (N_9908,N_9011,N_9170);
nor U9909 (N_9909,N_9241,N_9142);
or U9910 (N_9910,N_9260,N_9157);
and U9911 (N_9911,N_9418,N_9446);
or U9912 (N_9912,N_9105,N_9023);
and U9913 (N_9913,N_9148,N_9345);
nor U9914 (N_9914,N_9238,N_9250);
nor U9915 (N_9915,N_9133,N_9401);
nand U9916 (N_9916,N_9438,N_9203);
nand U9917 (N_9917,N_9424,N_9327);
or U9918 (N_9918,N_9297,N_9268);
nor U9919 (N_9919,N_9269,N_9270);
nor U9920 (N_9920,N_9021,N_9346);
or U9921 (N_9921,N_9356,N_9010);
xnor U9922 (N_9922,N_9189,N_9284);
nand U9923 (N_9923,N_9407,N_9071);
xor U9924 (N_9924,N_9356,N_9048);
nor U9925 (N_9925,N_9059,N_9429);
nor U9926 (N_9926,N_9308,N_9204);
nand U9927 (N_9927,N_9257,N_9009);
or U9928 (N_9928,N_9064,N_9008);
or U9929 (N_9929,N_9322,N_9083);
or U9930 (N_9930,N_9343,N_9451);
nor U9931 (N_9931,N_9140,N_9232);
xnor U9932 (N_9932,N_9038,N_9145);
xnor U9933 (N_9933,N_9338,N_9184);
nand U9934 (N_9934,N_9204,N_9022);
or U9935 (N_9935,N_9206,N_9270);
or U9936 (N_9936,N_9463,N_9051);
nand U9937 (N_9937,N_9263,N_9258);
and U9938 (N_9938,N_9175,N_9304);
or U9939 (N_9939,N_9209,N_9397);
and U9940 (N_9940,N_9479,N_9159);
nor U9941 (N_9941,N_9056,N_9270);
nor U9942 (N_9942,N_9384,N_9277);
nand U9943 (N_9943,N_9015,N_9207);
xor U9944 (N_9944,N_9431,N_9195);
or U9945 (N_9945,N_9042,N_9247);
nand U9946 (N_9946,N_9054,N_9090);
or U9947 (N_9947,N_9239,N_9290);
nand U9948 (N_9948,N_9040,N_9212);
nand U9949 (N_9949,N_9355,N_9291);
and U9950 (N_9950,N_9309,N_9162);
nor U9951 (N_9951,N_9355,N_9174);
xnor U9952 (N_9952,N_9067,N_9111);
or U9953 (N_9953,N_9040,N_9267);
xor U9954 (N_9954,N_9330,N_9162);
and U9955 (N_9955,N_9404,N_9426);
nand U9956 (N_9956,N_9184,N_9189);
nor U9957 (N_9957,N_9113,N_9122);
or U9958 (N_9958,N_9304,N_9431);
nor U9959 (N_9959,N_9139,N_9101);
nand U9960 (N_9960,N_9434,N_9324);
nand U9961 (N_9961,N_9182,N_9460);
nor U9962 (N_9962,N_9340,N_9446);
or U9963 (N_9963,N_9015,N_9329);
nand U9964 (N_9964,N_9419,N_9173);
and U9965 (N_9965,N_9204,N_9383);
nand U9966 (N_9966,N_9185,N_9111);
nand U9967 (N_9967,N_9376,N_9079);
and U9968 (N_9968,N_9370,N_9081);
and U9969 (N_9969,N_9064,N_9172);
nor U9970 (N_9970,N_9154,N_9425);
and U9971 (N_9971,N_9424,N_9174);
or U9972 (N_9972,N_9480,N_9197);
and U9973 (N_9973,N_9292,N_9060);
nor U9974 (N_9974,N_9103,N_9340);
or U9975 (N_9975,N_9207,N_9145);
xnor U9976 (N_9976,N_9104,N_9109);
nor U9977 (N_9977,N_9332,N_9024);
xor U9978 (N_9978,N_9066,N_9484);
xnor U9979 (N_9979,N_9002,N_9176);
or U9980 (N_9980,N_9435,N_9354);
xor U9981 (N_9981,N_9343,N_9094);
or U9982 (N_9982,N_9267,N_9018);
and U9983 (N_9983,N_9109,N_9064);
xor U9984 (N_9984,N_9140,N_9120);
and U9985 (N_9985,N_9252,N_9489);
or U9986 (N_9986,N_9040,N_9123);
nor U9987 (N_9987,N_9088,N_9375);
or U9988 (N_9988,N_9311,N_9454);
and U9989 (N_9989,N_9008,N_9407);
or U9990 (N_9990,N_9021,N_9256);
nor U9991 (N_9991,N_9067,N_9154);
nand U9992 (N_9992,N_9344,N_9347);
nor U9993 (N_9993,N_9194,N_9195);
xor U9994 (N_9994,N_9133,N_9202);
or U9995 (N_9995,N_9292,N_9221);
nor U9996 (N_9996,N_9398,N_9132);
and U9997 (N_9997,N_9485,N_9031);
and U9998 (N_9998,N_9320,N_9432);
nand U9999 (N_9999,N_9040,N_9195);
xnor U10000 (N_10000,N_9953,N_9521);
nor U10001 (N_10001,N_9894,N_9872);
xor U10002 (N_10002,N_9536,N_9566);
and U10003 (N_10003,N_9622,N_9795);
and U10004 (N_10004,N_9721,N_9895);
or U10005 (N_10005,N_9513,N_9746);
and U10006 (N_10006,N_9708,N_9585);
and U10007 (N_10007,N_9524,N_9979);
nand U10008 (N_10008,N_9621,N_9542);
xnor U10009 (N_10009,N_9885,N_9763);
nor U10010 (N_10010,N_9933,N_9645);
nand U10011 (N_10011,N_9984,N_9541);
xnor U10012 (N_10012,N_9792,N_9606);
xor U10013 (N_10013,N_9549,N_9725);
and U10014 (N_10014,N_9829,N_9640);
nand U10015 (N_10015,N_9976,N_9773);
xnor U10016 (N_10016,N_9660,N_9589);
or U10017 (N_10017,N_9540,N_9579);
nor U10018 (N_10018,N_9952,N_9887);
or U10019 (N_10019,N_9701,N_9569);
and U10020 (N_10020,N_9962,N_9989);
xor U10021 (N_10021,N_9946,N_9571);
xnor U10022 (N_10022,N_9652,N_9698);
and U10023 (N_10023,N_9884,N_9926);
nand U10024 (N_10024,N_9662,N_9882);
nand U10025 (N_10025,N_9557,N_9915);
or U10026 (N_10026,N_9604,N_9747);
xnor U10027 (N_10027,N_9696,N_9768);
nand U10028 (N_10028,N_9883,N_9972);
xnor U10029 (N_10029,N_9734,N_9617);
xnor U10030 (N_10030,N_9689,N_9899);
nor U10031 (N_10031,N_9871,N_9517);
and U10032 (N_10032,N_9879,N_9668);
or U10033 (N_10033,N_9749,N_9685);
nor U10034 (N_10034,N_9826,N_9651);
and U10035 (N_10035,N_9803,N_9527);
xnor U10036 (N_10036,N_9612,N_9788);
nand U10037 (N_10037,N_9684,N_9729);
nand U10038 (N_10038,N_9702,N_9922);
xor U10039 (N_10039,N_9714,N_9675);
nor U10040 (N_10040,N_9634,N_9906);
nor U10041 (N_10041,N_9947,N_9995);
xnor U10042 (N_10042,N_9780,N_9587);
and U10043 (N_10043,N_9761,N_9841);
and U10044 (N_10044,N_9713,N_9740);
xnor U10045 (N_10045,N_9608,N_9968);
or U10046 (N_10046,N_9808,N_9655);
and U10047 (N_10047,N_9874,N_9560);
and U10048 (N_10048,N_9593,N_9727);
xnor U10049 (N_10049,N_9902,N_9985);
nand U10050 (N_10050,N_9633,N_9870);
or U10051 (N_10051,N_9813,N_9515);
nand U10052 (N_10052,N_9750,N_9590);
nand U10053 (N_10053,N_9762,N_9562);
or U10054 (N_10054,N_9663,N_9938);
nand U10055 (N_10055,N_9558,N_9733);
nor U10056 (N_10056,N_9584,N_9856);
or U10057 (N_10057,N_9635,N_9983);
or U10058 (N_10058,N_9807,N_9583);
nor U10059 (N_10059,N_9508,N_9657);
and U10060 (N_10060,N_9965,N_9751);
nor U10061 (N_10061,N_9567,N_9719);
or U10062 (N_10062,N_9935,N_9741);
xnor U10063 (N_10063,N_9799,N_9615);
or U10064 (N_10064,N_9511,N_9950);
or U10065 (N_10065,N_9838,N_9930);
xor U10066 (N_10066,N_9544,N_9552);
xor U10067 (N_10067,N_9502,N_9978);
and U10068 (N_10068,N_9876,N_9865);
xor U10069 (N_10069,N_9743,N_9994);
or U10070 (N_10070,N_9691,N_9949);
or U10071 (N_10071,N_9681,N_9987);
and U10072 (N_10072,N_9538,N_9921);
nand U10073 (N_10073,N_9526,N_9969);
nor U10074 (N_10074,N_9832,N_9873);
nand U10075 (N_10075,N_9863,N_9929);
and U10076 (N_10076,N_9754,N_9744);
nand U10077 (N_10077,N_9755,N_9613);
or U10078 (N_10078,N_9506,N_9955);
nor U10079 (N_10079,N_9957,N_9996);
xor U10080 (N_10080,N_9945,N_9582);
and U10081 (N_10081,N_9827,N_9644);
and U10082 (N_10082,N_9893,N_9777);
nand U10083 (N_10083,N_9618,N_9507);
nand U10084 (N_10084,N_9784,N_9686);
nor U10085 (N_10085,N_9673,N_9975);
and U10086 (N_10086,N_9697,N_9992);
nand U10087 (N_10087,N_9948,N_9594);
and U10088 (N_10088,N_9501,N_9973);
nand U10089 (N_10089,N_9804,N_9716);
nor U10090 (N_10090,N_9522,N_9928);
nand U10091 (N_10091,N_9722,N_9598);
nor U10092 (N_10092,N_9852,N_9533);
xor U10093 (N_10093,N_9703,N_9658);
nor U10094 (N_10094,N_9636,N_9610);
nor U10095 (N_10095,N_9539,N_9659);
nor U10096 (N_10096,N_9596,N_9919);
and U10097 (N_10097,N_9869,N_9556);
or U10098 (N_10098,N_9866,N_9855);
nor U10099 (N_10099,N_9731,N_9738);
nand U10100 (N_10100,N_9981,N_9927);
nand U10101 (N_10101,N_9626,N_9599);
and U10102 (N_10102,N_9525,N_9537);
xor U10103 (N_10103,N_9553,N_9988);
xor U10104 (N_10104,N_9580,N_9806);
and U10105 (N_10105,N_9670,N_9790);
and U10106 (N_10106,N_9889,N_9509);
nand U10107 (N_10107,N_9920,N_9656);
or U10108 (N_10108,N_9817,N_9966);
nor U10109 (N_10109,N_9529,N_9816);
nand U10110 (N_10110,N_9682,N_9842);
nand U10111 (N_10111,N_9564,N_9646);
nor U10112 (N_10112,N_9774,N_9575);
and U10113 (N_10113,N_9900,N_9923);
nor U10114 (N_10114,N_9964,N_9998);
nor U10115 (N_10115,N_9530,N_9959);
and U10116 (N_10116,N_9665,N_9849);
or U10117 (N_10117,N_9783,N_9862);
and U10118 (N_10118,N_9867,N_9916);
nor U10119 (N_10119,N_9624,N_9531);
xnor U10120 (N_10120,N_9548,N_9999);
and U10121 (N_10121,N_9910,N_9875);
and U10122 (N_10122,N_9825,N_9909);
nor U10123 (N_10123,N_9631,N_9643);
and U10124 (N_10124,N_9718,N_9595);
and U10125 (N_10125,N_9504,N_9831);
xnor U10126 (N_10126,N_9601,N_9756);
xnor U10127 (N_10127,N_9528,N_9822);
xnor U10128 (N_10128,N_9925,N_9737);
or U10129 (N_10129,N_9888,N_9735);
xor U10130 (N_10130,N_9648,N_9778);
and U10131 (N_10131,N_9937,N_9514);
or U10132 (N_10132,N_9802,N_9694);
nand U10133 (N_10133,N_9674,N_9934);
or U10134 (N_10134,N_9758,N_9791);
or U10135 (N_10135,N_9914,N_9629);
nor U10136 (N_10136,N_9667,N_9864);
and U10137 (N_10137,N_9980,N_9620);
nand U10138 (N_10138,N_9877,N_9551);
xnor U10139 (N_10139,N_9690,N_9903);
xor U10140 (N_10140,N_9990,N_9638);
and U10141 (N_10141,N_9739,N_9971);
xnor U10142 (N_10142,N_9611,N_9745);
and U10143 (N_10143,N_9858,N_9772);
nand U10144 (N_10144,N_9770,N_9878);
or U10145 (N_10145,N_9680,N_9677);
xor U10146 (N_10146,N_9700,N_9545);
xnor U10147 (N_10147,N_9821,N_9664);
nor U10148 (N_10148,N_9845,N_9764);
nand U10149 (N_10149,N_9880,N_9688);
nand U10150 (N_10150,N_9786,N_9518);
nand U10151 (N_10151,N_9912,N_9785);
and U10152 (N_10152,N_9707,N_9809);
or U10153 (N_10153,N_9661,N_9759);
xnor U10154 (N_10154,N_9890,N_9717);
or U10155 (N_10155,N_9844,N_9710);
and U10156 (N_10156,N_9840,N_9534);
xnor U10157 (N_10157,N_9997,N_9881);
nand U10158 (N_10158,N_9850,N_9641);
nor U10159 (N_10159,N_9603,N_9535);
and U10160 (N_10160,N_9924,N_9766);
nor U10161 (N_10161,N_9628,N_9779);
nor U10162 (N_10162,N_9810,N_9576);
or U10163 (N_10163,N_9723,N_9720);
or U10164 (N_10164,N_9848,N_9588);
or U10165 (N_10165,N_9781,N_9847);
nand U10166 (N_10166,N_9752,N_9715);
or U10167 (N_10167,N_9577,N_9555);
or U10168 (N_10168,N_9861,N_9753);
or U10169 (N_10169,N_9907,N_9547);
or U10170 (N_10170,N_9854,N_9695);
and U10171 (N_10171,N_9836,N_9775);
and U10172 (N_10172,N_9820,N_9500);
nand U10173 (N_10173,N_9730,N_9616);
or U10174 (N_10174,N_9614,N_9835);
nor U10175 (N_10175,N_9956,N_9597);
nand U10176 (N_10176,N_9570,N_9742);
or U10177 (N_10177,N_9932,N_9812);
or U10178 (N_10178,N_9591,N_9666);
and U10179 (N_10179,N_9982,N_9503);
and U10180 (N_10180,N_9819,N_9600);
xnor U10181 (N_10181,N_9574,N_9853);
xnor U10182 (N_10182,N_9942,N_9523);
xor U10183 (N_10183,N_9961,N_9732);
xor U10184 (N_10184,N_9602,N_9805);
nand U10185 (N_10185,N_9728,N_9970);
xor U10186 (N_10186,N_9512,N_9532);
xnor U10187 (N_10187,N_9823,N_9798);
nor U10188 (N_10188,N_9771,N_9828);
and U10189 (N_10189,N_9619,N_9625);
or U10190 (N_10190,N_9510,N_9904);
and U10191 (N_10191,N_9650,N_9649);
nand U10192 (N_10192,N_9519,N_9931);
and U10193 (N_10193,N_9572,N_9859);
nand U10194 (N_10194,N_9669,N_9793);
nor U10195 (N_10195,N_9627,N_9706);
nand U10196 (N_10196,N_9672,N_9679);
nor U10197 (N_10197,N_9676,N_9986);
nor U10198 (N_10198,N_9561,N_9958);
or U10199 (N_10199,N_9693,N_9712);
nor U10200 (N_10200,N_9559,N_9767);
and U10201 (N_10201,N_9839,N_9917);
and U10202 (N_10202,N_9607,N_9898);
or U10203 (N_10203,N_9578,N_9776);
xnor U10204 (N_10204,N_9581,N_9757);
or U10205 (N_10205,N_9760,N_9833);
nand U10206 (N_10206,N_9568,N_9726);
nand U10207 (N_10207,N_9837,N_9609);
or U10208 (N_10208,N_9991,N_9993);
nand U10209 (N_10209,N_9846,N_9683);
nor U10210 (N_10210,N_9769,N_9797);
xor U10211 (N_10211,N_9505,N_9811);
and U10212 (N_10212,N_9520,N_9851);
or U10213 (N_10213,N_9642,N_9913);
and U10214 (N_10214,N_9671,N_9789);
xor U10215 (N_10215,N_9905,N_9605);
and U10216 (N_10216,N_9834,N_9748);
and U10217 (N_10217,N_9765,N_9939);
xor U10218 (N_10218,N_9573,N_9974);
and U10219 (N_10219,N_9830,N_9711);
xnor U10220 (N_10220,N_9516,N_9586);
nand U10221 (N_10221,N_9891,N_9654);
xnor U10222 (N_10222,N_9901,N_9857);
nor U10223 (N_10223,N_9886,N_9843);
xnor U10224 (N_10224,N_9796,N_9554);
and U10225 (N_10225,N_9687,N_9941);
or U10226 (N_10226,N_9782,N_9709);
or U10227 (N_10227,N_9892,N_9692);
and U10228 (N_10228,N_9860,N_9818);
and U10229 (N_10229,N_9736,N_9936);
xor U10230 (N_10230,N_9951,N_9546);
nor U10231 (N_10231,N_9960,N_9550);
and U10232 (N_10232,N_9815,N_9940);
and U10233 (N_10233,N_9699,N_9897);
nor U10234 (N_10234,N_9647,N_9896);
or U10235 (N_10235,N_9678,N_9705);
and U10236 (N_10236,N_9977,N_9632);
nor U10237 (N_10237,N_9943,N_9814);
nand U10238 (N_10238,N_9653,N_9800);
or U10239 (N_10239,N_9637,N_9954);
nand U10240 (N_10240,N_9543,N_9787);
xor U10241 (N_10241,N_9967,N_9824);
xor U10242 (N_10242,N_9724,N_9963);
nand U10243 (N_10243,N_9592,N_9801);
xor U10244 (N_10244,N_9630,N_9868);
xor U10245 (N_10245,N_9918,N_9639);
or U10246 (N_10246,N_9623,N_9944);
or U10247 (N_10247,N_9794,N_9565);
nor U10248 (N_10248,N_9563,N_9704);
xnor U10249 (N_10249,N_9908,N_9911);
nor U10250 (N_10250,N_9940,N_9619);
and U10251 (N_10251,N_9770,N_9630);
nand U10252 (N_10252,N_9990,N_9984);
nand U10253 (N_10253,N_9991,N_9795);
xnor U10254 (N_10254,N_9898,N_9905);
nand U10255 (N_10255,N_9669,N_9519);
and U10256 (N_10256,N_9892,N_9644);
or U10257 (N_10257,N_9699,N_9857);
and U10258 (N_10258,N_9775,N_9801);
or U10259 (N_10259,N_9611,N_9502);
xnor U10260 (N_10260,N_9856,N_9805);
xnor U10261 (N_10261,N_9505,N_9551);
and U10262 (N_10262,N_9818,N_9945);
xnor U10263 (N_10263,N_9973,N_9730);
and U10264 (N_10264,N_9948,N_9977);
and U10265 (N_10265,N_9510,N_9692);
xor U10266 (N_10266,N_9920,N_9966);
or U10267 (N_10267,N_9835,N_9738);
or U10268 (N_10268,N_9629,N_9604);
nand U10269 (N_10269,N_9837,N_9993);
xor U10270 (N_10270,N_9861,N_9905);
xor U10271 (N_10271,N_9643,N_9790);
nand U10272 (N_10272,N_9579,N_9718);
or U10273 (N_10273,N_9852,N_9859);
nand U10274 (N_10274,N_9589,N_9900);
nor U10275 (N_10275,N_9777,N_9665);
nor U10276 (N_10276,N_9772,N_9954);
xor U10277 (N_10277,N_9796,N_9563);
and U10278 (N_10278,N_9775,N_9671);
nor U10279 (N_10279,N_9618,N_9679);
xor U10280 (N_10280,N_9899,N_9606);
nor U10281 (N_10281,N_9862,N_9976);
and U10282 (N_10282,N_9656,N_9716);
xnor U10283 (N_10283,N_9683,N_9832);
nor U10284 (N_10284,N_9569,N_9972);
nor U10285 (N_10285,N_9504,N_9625);
or U10286 (N_10286,N_9957,N_9723);
nor U10287 (N_10287,N_9503,N_9692);
xor U10288 (N_10288,N_9745,N_9893);
or U10289 (N_10289,N_9535,N_9752);
and U10290 (N_10290,N_9551,N_9788);
and U10291 (N_10291,N_9542,N_9989);
nand U10292 (N_10292,N_9946,N_9996);
or U10293 (N_10293,N_9632,N_9724);
and U10294 (N_10294,N_9818,N_9623);
xnor U10295 (N_10295,N_9719,N_9659);
and U10296 (N_10296,N_9790,N_9782);
nand U10297 (N_10297,N_9725,N_9783);
nor U10298 (N_10298,N_9503,N_9867);
xnor U10299 (N_10299,N_9645,N_9532);
nor U10300 (N_10300,N_9643,N_9530);
nand U10301 (N_10301,N_9798,N_9588);
nor U10302 (N_10302,N_9571,N_9747);
nand U10303 (N_10303,N_9978,N_9600);
or U10304 (N_10304,N_9762,N_9523);
or U10305 (N_10305,N_9669,N_9837);
nand U10306 (N_10306,N_9836,N_9571);
or U10307 (N_10307,N_9932,N_9826);
nor U10308 (N_10308,N_9726,N_9789);
nor U10309 (N_10309,N_9612,N_9514);
nor U10310 (N_10310,N_9763,N_9716);
or U10311 (N_10311,N_9871,N_9576);
nor U10312 (N_10312,N_9501,N_9649);
and U10313 (N_10313,N_9734,N_9758);
nor U10314 (N_10314,N_9708,N_9917);
xor U10315 (N_10315,N_9843,N_9776);
or U10316 (N_10316,N_9551,N_9817);
or U10317 (N_10317,N_9673,N_9575);
nor U10318 (N_10318,N_9635,N_9708);
and U10319 (N_10319,N_9901,N_9884);
nand U10320 (N_10320,N_9558,N_9627);
or U10321 (N_10321,N_9994,N_9910);
nand U10322 (N_10322,N_9615,N_9776);
nor U10323 (N_10323,N_9964,N_9526);
nand U10324 (N_10324,N_9851,N_9691);
nor U10325 (N_10325,N_9519,N_9935);
nor U10326 (N_10326,N_9615,N_9866);
xor U10327 (N_10327,N_9713,N_9863);
or U10328 (N_10328,N_9947,N_9502);
nand U10329 (N_10329,N_9609,N_9702);
and U10330 (N_10330,N_9698,N_9961);
xor U10331 (N_10331,N_9888,N_9938);
or U10332 (N_10332,N_9748,N_9540);
nor U10333 (N_10333,N_9825,N_9841);
and U10334 (N_10334,N_9984,N_9971);
xor U10335 (N_10335,N_9668,N_9636);
nor U10336 (N_10336,N_9764,N_9934);
or U10337 (N_10337,N_9886,N_9796);
xor U10338 (N_10338,N_9991,N_9727);
xnor U10339 (N_10339,N_9556,N_9884);
nand U10340 (N_10340,N_9601,N_9863);
or U10341 (N_10341,N_9659,N_9880);
xnor U10342 (N_10342,N_9599,N_9828);
nor U10343 (N_10343,N_9532,N_9803);
nor U10344 (N_10344,N_9551,N_9924);
nor U10345 (N_10345,N_9864,N_9772);
or U10346 (N_10346,N_9637,N_9640);
and U10347 (N_10347,N_9975,N_9537);
and U10348 (N_10348,N_9867,N_9505);
xor U10349 (N_10349,N_9861,N_9826);
nand U10350 (N_10350,N_9900,N_9634);
nand U10351 (N_10351,N_9856,N_9783);
and U10352 (N_10352,N_9666,N_9533);
and U10353 (N_10353,N_9778,N_9866);
nand U10354 (N_10354,N_9724,N_9542);
xnor U10355 (N_10355,N_9791,N_9927);
xnor U10356 (N_10356,N_9715,N_9829);
nand U10357 (N_10357,N_9522,N_9523);
and U10358 (N_10358,N_9581,N_9692);
or U10359 (N_10359,N_9857,N_9568);
and U10360 (N_10360,N_9653,N_9581);
nand U10361 (N_10361,N_9827,N_9564);
or U10362 (N_10362,N_9554,N_9736);
nor U10363 (N_10363,N_9937,N_9539);
nand U10364 (N_10364,N_9873,N_9561);
nand U10365 (N_10365,N_9562,N_9722);
and U10366 (N_10366,N_9600,N_9602);
or U10367 (N_10367,N_9528,N_9553);
nand U10368 (N_10368,N_9808,N_9721);
or U10369 (N_10369,N_9736,N_9846);
nor U10370 (N_10370,N_9926,N_9971);
and U10371 (N_10371,N_9577,N_9792);
nand U10372 (N_10372,N_9605,N_9674);
and U10373 (N_10373,N_9641,N_9926);
nor U10374 (N_10374,N_9695,N_9662);
nand U10375 (N_10375,N_9763,N_9874);
or U10376 (N_10376,N_9536,N_9662);
nand U10377 (N_10377,N_9833,N_9585);
nand U10378 (N_10378,N_9537,N_9879);
or U10379 (N_10379,N_9897,N_9772);
nor U10380 (N_10380,N_9609,N_9955);
and U10381 (N_10381,N_9566,N_9580);
and U10382 (N_10382,N_9821,N_9592);
xnor U10383 (N_10383,N_9913,N_9833);
and U10384 (N_10384,N_9916,N_9983);
xor U10385 (N_10385,N_9680,N_9767);
xor U10386 (N_10386,N_9956,N_9831);
nand U10387 (N_10387,N_9608,N_9997);
xnor U10388 (N_10388,N_9676,N_9750);
and U10389 (N_10389,N_9557,N_9930);
nor U10390 (N_10390,N_9669,N_9711);
and U10391 (N_10391,N_9647,N_9537);
nand U10392 (N_10392,N_9902,N_9892);
nand U10393 (N_10393,N_9629,N_9552);
nand U10394 (N_10394,N_9757,N_9732);
nor U10395 (N_10395,N_9508,N_9831);
or U10396 (N_10396,N_9917,N_9504);
or U10397 (N_10397,N_9707,N_9680);
and U10398 (N_10398,N_9781,N_9700);
nand U10399 (N_10399,N_9738,N_9718);
or U10400 (N_10400,N_9896,N_9871);
and U10401 (N_10401,N_9507,N_9795);
xnor U10402 (N_10402,N_9761,N_9642);
nor U10403 (N_10403,N_9541,N_9759);
nand U10404 (N_10404,N_9995,N_9683);
and U10405 (N_10405,N_9833,N_9714);
nand U10406 (N_10406,N_9783,N_9641);
nand U10407 (N_10407,N_9961,N_9733);
nand U10408 (N_10408,N_9714,N_9711);
and U10409 (N_10409,N_9796,N_9618);
nor U10410 (N_10410,N_9583,N_9715);
or U10411 (N_10411,N_9736,N_9614);
or U10412 (N_10412,N_9779,N_9676);
and U10413 (N_10413,N_9521,N_9731);
nor U10414 (N_10414,N_9706,N_9658);
and U10415 (N_10415,N_9625,N_9532);
nor U10416 (N_10416,N_9512,N_9928);
nand U10417 (N_10417,N_9640,N_9709);
nor U10418 (N_10418,N_9958,N_9575);
and U10419 (N_10419,N_9936,N_9915);
nand U10420 (N_10420,N_9526,N_9931);
nor U10421 (N_10421,N_9550,N_9696);
or U10422 (N_10422,N_9656,N_9721);
xor U10423 (N_10423,N_9905,N_9779);
or U10424 (N_10424,N_9838,N_9559);
or U10425 (N_10425,N_9761,N_9970);
xor U10426 (N_10426,N_9973,N_9883);
and U10427 (N_10427,N_9636,N_9509);
and U10428 (N_10428,N_9627,N_9628);
or U10429 (N_10429,N_9796,N_9809);
nand U10430 (N_10430,N_9522,N_9965);
nor U10431 (N_10431,N_9635,N_9966);
and U10432 (N_10432,N_9947,N_9994);
or U10433 (N_10433,N_9701,N_9550);
nand U10434 (N_10434,N_9612,N_9973);
nand U10435 (N_10435,N_9505,N_9868);
nor U10436 (N_10436,N_9595,N_9955);
and U10437 (N_10437,N_9503,N_9650);
nor U10438 (N_10438,N_9706,N_9906);
xnor U10439 (N_10439,N_9636,N_9517);
and U10440 (N_10440,N_9980,N_9806);
and U10441 (N_10441,N_9967,N_9819);
and U10442 (N_10442,N_9757,N_9896);
nand U10443 (N_10443,N_9562,N_9569);
xor U10444 (N_10444,N_9846,N_9605);
and U10445 (N_10445,N_9889,N_9863);
or U10446 (N_10446,N_9732,N_9872);
or U10447 (N_10447,N_9567,N_9535);
or U10448 (N_10448,N_9958,N_9960);
nor U10449 (N_10449,N_9675,N_9915);
and U10450 (N_10450,N_9916,N_9627);
xnor U10451 (N_10451,N_9782,N_9830);
xor U10452 (N_10452,N_9960,N_9671);
and U10453 (N_10453,N_9615,N_9958);
or U10454 (N_10454,N_9528,N_9612);
nand U10455 (N_10455,N_9953,N_9879);
xnor U10456 (N_10456,N_9749,N_9755);
and U10457 (N_10457,N_9552,N_9770);
nand U10458 (N_10458,N_9974,N_9945);
or U10459 (N_10459,N_9810,N_9596);
nand U10460 (N_10460,N_9580,N_9915);
or U10461 (N_10461,N_9608,N_9599);
xor U10462 (N_10462,N_9510,N_9650);
and U10463 (N_10463,N_9748,N_9931);
xor U10464 (N_10464,N_9644,N_9932);
or U10465 (N_10465,N_9756,N_9503);
or U10466 (N_10466,N_9916,N_9502);
or U10467 (N_10467,N_9984,N_9615);
xnor U10468 (N_10468,N_9611,N_9715);
or U10469 (N_10469,N_9915,N_9853);
xnor U10470 (N_10470,N_9616,N_9853);
or U10471 (N_10471,N_9555,N_9613);
and U10472 (N_10472,N_9512,N_9597);
nor U10473 (N_10473,N_9916,N_9941);
nor U10474 (N_10474,N_9552,N_9570);
nor U10475 (N_10475,N_9716,N_9973);
xor U10476 (N_10476,N_9647,N_9787);
and U10477 (N_10477,N_9852,N_9523);
nand U10478 (N_10478,N_9771,N_9759);
nand U10479 (N_10479,N_9686,N_9917);
xnor U10480 (N_10480,N_9907,N_9725);
nand U10481 (N_10481,N_9915,N_9584);
nand U10482 (N_10482,N_9509,N_9873);
nand U10483 (N_10483,N_9983,N_9853);
or U10484 (N_10484,N_9594,N_9945);
nor U10485 (N_10485,N_9628,N_9993);
or U10486 (N_10486,N_9517,N_9723);
and U10487 (N_10487,N_9791,N_9600);
nand U10488 (N_10488,N_9902,N_9955);
nand U10489 (N_10489,N_9899,N_9887);
or U10490 (N_10490,N_9582,N_9779);
nor U10491 (N_10491,N_9894,N_9805);
and U10492 (N_10492,N_9560,N_9653);
or U10493 (N_10493,N_9559,N_9734);
and U10494 (N_10494,N_9862,N_9781);
xnor U10495 (N_10495,N_9502,N_9623);
xnor U10496 (N_10496,N_9691,N_9521);
nand U10497 (N_10497,N_9754,N_9848);
nor U10498 (N_10498,N_9913,N_9914);
or U10499 (N_10499,N_9850,N_9824);
and U10500 (N_10500,N_10207,N_10486);
xor U10501 (N_10501,N_10396,N_10475);
nor U10502 (N_10502,N_10218,N_10476);
or U10503 (N_10503,N_10230,N_10042);
or U10504 (N_10504,N_10110,N_10141);
and U10505 (N_10505,N_10283,N_10293);
and U10506 (N_10506,N_10397,N_10077);
and U10507 (N_10507,N_10348,N_10213);
and U10508 (N_10508,N_10172,N_10227);
xor U10509 (N_10509,N_10105,N_10342);
nand U10510 (N_10510,N_10058,N_10177);
nand U10511 (N_10511,N_10387,N_10037);
or U10512 (N_10512,N_10125,N_10067);
xnor U10513 (N_10513,N_10115,N_10246);
nand U10514 (N_10514,N_10338,N_10161);
or U10515 (N_10515,N_10118,N_10367);
xor U10516 (N_10516,N_10210,N_10461);
nand U10517 (N_10517,N_10312,N_10109);
nand U10518 (N_10518,N_10340,N_10262);
and U10519 (N_10519,N_10386,N_10143);
xor U10520 (N_10520,N_10473,N_10052);
nor U10521 (N_10521,N_10045,N_10343);
or U10522 (N_10522,N_10019,N_10256);
nand U10523 (N_10523,N_10026,N_10147);
nor U10524 (N_10524,N_10378,N_10003);
nor U10525 (N_10525,N_10316,N_10390);
nor U10526 (N_10526,N_10201,N_10306);
nand U10527 (N_10527,N_10490,N_10251);
or U10528 (N_10528,N_10453,N_10439);
nand U10529 (N_10529,N_10322,N_10195);
and U10530 (N_10530,N_10469,N_10139);
nand U10531 (N_10531,N_10173,N_10225);
xor U10532 (N_10532,N_10265,N_10267);
xnor U10533 (N_10533,N_10122,N_10468);
xor U10534 (N_10534,N_10126,N_10063);
nor U10535 (N_10535,N_10268,N_10248);
or U10536 (N_10536,N_10442,N_10382);
and U10537 (N_10537,N_10361,N_10385);
nor U10538 (N_10538,N_10437,N_10011);
and U10539 (N_10539,N_10409,N_10184);
or U10540 (N_10540,N_10325,N_10178);
nor U10541 (N_10541,N_10354,N_10159);
and U10542 (N_10542,N_10229,N_10169);
or U10543 (N_10543,N_10328,N_10440);
and U10544 (N_10544,N_10100,N_10152);
xnor U10545 (N_10545,N_10443,N_10188);
nand U10546 (N_10546,N_10456,N_10404);
or U10547 (N_10547,N_10001,N_10131);
xnor U10548 (N_10548,N_10451,N_10164);
and U10549 (N_10549,N_10311,N_10355);
nor U10550 (N_10550,N_10029,N_10344);
and U10551 (N_10551,N_10465,N_10000);
nand U10552 (N_10552,N_10193,N_10155);
and U10553 (N_10553,N_10481,N_10447);
nor U10554 (N_10554,N_10096,N_10472);
nand U10555 (N_10555,N_10309,N_10085);
nor U10556 (N_10556,N_10408,N_10036);
xor U10557 (N_10557,N_10179,N_10013);
and U10558 (N_10558,N_10324,N_10016);
and U10559 (N_10559,N_10307,N_10452);
and U10560 (N_10560,N_10030,N_10339);
nor U10561 (N_10561,N_10388,N_10427);
nor U10562 (N_10562,N_10241,N_10223);
nor U10563 (N_10563,N_10253,N_10182);
and U10564 (N_10564,N_10133,N_10369);
and U10565 (N_10565,N_10148,N_10445);
nor U10566 (N_10566,N_10090,N_10236);
xor U10567 (N_10567,N_10022,N_10235);
nand U10568 (N_10568,N_10429,N_10033);
or U10569 (N_10569,N_10093,N_10135);
nand U10570 (N_10570,N_10480,N_10413);
xnor U10571 (N_10571,N_10217,N_10204);
nand U10572 (N_10572,N_10402,N_10086);
xor U10573 (N_10573,N_10154,N_10292);
or U10574 (N_10574,N_10424,N_10051);
or U10575 (N_10575,N_10166,N_10124);
or U10576 (N_10576,N_10203,N_10289);
and U10577 (N_10577,N_10286,N_10057);
or U10578 (N_10578,N_10291,N_10336);
and U10579 (N_10579,N_10112,N_10081);
and U10580 (N_10580,N_10346,N_10394);
xor U10581 (N_10581,N_10260,N_10295);
xor U10582 (N_10582,N_10103,N_10047);
xor U10583 (N_10583,N_10384,N_10138);
nor U10584 (N_10584,N_10220,N_10238);
and U10585 (N_10585,N_10454,N_10027);
nor U10586 (N_10586,N_10314,N_10215);
or U10587 (N_10587,N_10175,N_10243);
xnor U10588 (N_10588,N_10163,N_10315);
nor U10589 (N_10589,N_10471,N_10463);
and U10590 (N_10590,N_10351,N_10145);
or U10591 (N_10591,N_10299,N_10279);
and U10592 (N_10592,N_10405,N_10107);
and U10593 (N_10593,N_10054,N_10353);
nor U10594 (N_10594,N_10214,N_10282);
xnor U10595 (N_10595,N_10134,N_10298);
and U10596 (N_10596,N_10320,N_10167);
and U10597 (N_10597,N_10383,N_10464);
and U10598 (N_10598,N_10233,N_10467);
nor U10599 (N_10599,N_10357,N_10259);
xnor U10600 (N_10600,N_10209,N_10035);
or U10601 (N_10601,N_10423,N_10417);
nand U10602 (N_10602,N_10375,N_10428);
and U10603 (N_10603,N_10121,N_10261);
or U10604 (N_10604,N_10129,N_10313);
and U10605 (N_10605,N_10123,N_10478);
xor U10606 (N_10606,N_10113,N_10263);
nand U10607 (N_10607,N_10075,N_10380);
and U10608 (N_10608,N_10335,N_10174);
and U10609 (N_10609,N_10162,N_10015);
and U10610 (N_10610,N_10171,N_10021);
or U10611 (N_10611,N_10458,N_10247);
nor U10612 (N_10612,N_10140,N_10410);
nand U10613 (N_10613,N_10494,N_10258);
nor U10614 (N_10614,N_10434,N_10421);
nor U10615 (N_10615,N_10412,N_10466);
and U10616 (N_10616,N_10190,N_10366);
nor U10617 (N_10617,N_10219,N_10297);
nand U10618 (N_10618,N_10108,N_10395);
and U10619 (N_10619,N_10005,N_10270);
nor U10620 (N_10620,N_10371,N_10091);
xor U10621 (N_10621,N_10128,N_10043);
nor U10622 (N_10622,N_10023,N_10255);
or U10623 (N_10623,N_10450,N_10012);
xnor U10624 (N_10624,N_10492,N_10422);
and U10625 (N_10625,N_10448,N_10381);
nand U10626 (N_10626,N_10474,N_10333);
nand U10627 (N_10627,N_10205,N_10137);
or U10628 (N_10628,N_10431,N_10222);
nand U10629 (N_10629,N_10416,N_10127);
nand U10630 (N_10630,N_10020,N_10226);
xor U10631 (N_10631,N_10053,N_10014);
nor U10632 (N_10632,N_10358,N_10379);
or U10633 (N_10633,N_10323,N_10294);
nand U10634 (N_10634,N_10455,N_10157);
xnor U10635 (N_10635,N_10069,N_10132);
xnor U10636 (N_10636,N_10274,N_10362);
nand U10637 (N_10637,N_10094,N_10496);
or U10638 (N_10638,N_10040,N_10497);
xor U10639 (N_10639,N_10277,N_10136);
nand U10640 (N_10640,N_10116,N_10304);
nand U10641 (N_10641,N_10071,N_10446);
and U10642 (N_10642,N_10106,N_10482);
and U10643 (N_10643,N_10060,N_10046);
xor U10644 (N_10644,N_10004,N_10089);
xnor U10645 (N_10645,N_10206,N_10250);
xor U10646 (N_10646,N_10444,N_10317);
xnor U10647 (N_10647,N_10006,N_10048);
nor U10648 (N_10648,N_10153,N_10158);
xor U10649 (N_10649,N_10165,N_10460);
and U10650 (N_10650,N_10080,N_10007);
and U10651 (N_10651,N_10326,N_10280);
nand U10652 (N_10652,N_10187,N_10038);
nand U10653 (N_10653,N_10308,N_10287);
xor U10654 (N_10654,N_10170,N_10319);
or U10655 (N_10655,N_10156,N_10407);
nor U10656 (N_10656,N_10079,N_10149);
and U10657 (N_10657,N_10401,N_10373);
nand U10658 (N_10658,N_10426,N_10266);
xor U10659 (N_10659,N_10087,N_10252);
or U10660 (N_10660,N_10088,N_10073);
nor U10661 (N_10661,N_10400,N_10078);
xnor U10662 (N_10662,N_10403,N_10150);
nor U10663 (N_10663,N_10025,N_10321);
or U10664 (N_10664,N_10199,N_10430);
or U10665 (N_10665,N_10024,N_10111);
nor U10666 (N_10666,N_10151,N_10099);
and U10667 (N_10667,N_10420,N_10212);
nand U10668 (N_10668,N_10031,N_10245);
nand U10669 (N_10669,N_10232,N_10216);
nor U10670 (N_10670,N_10425,N_10327);
and U10671 (N_10671,N_10377,N_10041);
nand U10672 (N_10672,N_10269,N_10296);
xnor U10673 (N_10673,N_10484,N_10104);
xor U10674 (N_10674,N_10363,N_10228);
xnor U10675 (N_10675,N_10186,N_10406);
nor U10676 (N_10676,N_10275,N_10376);
nor U10677 (N_10677,N_10114,N_10374);
nor U10678 (N_10678,N_10084,N_10176);
and U10679 (N_10679,N_10415,N_10370);
xor U10680 (N_10680,N_10160,N_10345);
nand U10681 (N_10681,N_10364,N_10144);
nor U10682 (N_10682,N_10393,N_10208);
xor U10683 (N_10683,N_10183,N_10389);
nor U10684 (N_10684,N_10337,N_10462);
xor U10685 (N_10685,N_10008,N_10264);
nor U10686 (N_10686,N_10276,N_10350);
nand U10687 (N_10687,N_10441,N_10146);
xor U10688 (N_10688,N_10498,N_10168);
nor U10689 (N_10689,N_10002,N_10330);
nand U10690 (N_10690,N_10049,N_10244);
or U10691 (N_10691,N_10194,N_10300);
xor U10692 (N_10692,N_10301,N_10050);
and U10693 (N_10693,N_10055,N_10302);
nor U10694 (N_10694,N_10198,N_10368);
nand U10695 (N_10695,N_10284,N_10281);
and U10696 (N_10696,N_10010,N_10449);
and U10697 (N_10697,N_10399,N_10189);
xor U10698 (N_10698,N_10365,N_10117);
nor U10699 (N_10699,N_10436,N_10334);
and U10700 (N_10700,N_10082,N_10142);
xor U10701 (N_10701,N_10391,N_10477);
or U10702 (N_10702,N_10331,N_10039);
or U10703 (N_10703,N_10418,N_10392);
xnor U10704 (N_10704,N_10211,N_10181);
nand U10705 (N_10705,N_10196,N_10095);
nand U10706 (N_10706,N_10076,N_10242);
nor U10707 (N_10707,N_10062,N_10070);
or U10708 (N_10708,N_10254,N_10059);
and U10709 (N_10709,N_10098,N_10290);
and U10710 (N_10710,N_10192,N_10285);
and U10711 (N_10711,N_10221,N_10349);
and U10712 (N_10712,N_10332,N_10288);
nand U10713 (N_10713,N_10028,N_10119);
nor U10714 (N_10714,N_10257,N_10065);
and U10715 (N_10715,N_10032,N_10278);
xor U10716 (N_10716,N_10074,N_10329);
and U10717 (N_10717,N_10224,N_10191);
xor U10718 (N_10718,N_10120,N_10249);
nor U10719 (N_10719,N_10352,N_10347);
nor U10720 (N_10720,N_10305,N_10061);
xor U10721 (N_10721,N_10239,N_10034);
xnor U10722 (N_10722,N_10068,N_10341);
nor U10723 (N_10723,N_10491,N_10470);
nand U10724 (N_10724,N_10372,N_10438);
nand U10725 (N_10725,N_10495,N_10064);
nor U10726 (N_10726,N_10493,N_10414);
and U10727 (N_10727,N_10411,N_10487);
xor U10728 (N_10728,N_10130,N_10310);
nand U10729 (N_10729,N_10092,N_10083);
or U10730 (N_10730,N_10419,N_10272);
or U10731 (N_10731,N_10435,N_10483);
and U10732 (N_10732,N_10101,N_10432);
xnor U10733 (N_10733,N_10185,N_10433);
and U10734 (N_10734,N_10240,N_10489);
nor U10735 (N_10735,N_10018,N_10271);
and U10736 (N_10736,N_10197,N_10273);
or U10737 (N_10737,N_10359,N_10237);
or U10738 (N_10738,N_10200,N_10231);
and U10739 (N_10739,N_10066,N_10485);
or U10740 (N_10740,N_10009,N_10488);
or U10741 (N_10741,N_10097,N_10056);
nor U10742 (N_10742,N_10356,N_10457);
nor U10743 (N_10743,N_10303,N_10044);
or U10744 (N_10744,N_10318,N_10202);
and U10745 (N_10745,N_10360,N_10102);
or U10746 (N_10746,N_10459,N_10234);
or U10747 (N_10747,N_10180,N_10499);
nand U10748 (N_10748,N_10479,N_10017);
nand U10749 (N_10749,N_10398,N_10072);
xnor U10750 (N_10750,N_10019,N_10315);
and U10751 (N_10751,N_10464,N_10257);
nand U10752 (N_10752,N_10003,N_10147);
and U10753 (N_10753,N_10474,N_10053);
nor U10754 (N_10754,N_10338,N_10296);
nor U10755 (N_10755,N_10356,N_10209);
nor U10756 (N_10756,N_10014,N_10418);
xnor U10757 (N_10757,N_10051,N_10035);
nand U10758 (N_10758,N_10320,N_10037);
nor U10759 (N_10759,N_10228,N_10065);
or U10760 (N_10760,N_10198,N_10104);
or U10761 (N_10761,N_10198,N_10355);
xnor U10762 (N_10762,N_10157,N_10467);
or U10763 (N_10763,N_10304,N_10228);
nand U10764 (N_10764,N_10121,N_10097);
and U10765 (N_10765,N_10091,N_10408);
nand U10766 (N_10766,N_10281,N_10407);
xor U10767 (N_10767,N_10465,N_10285);
or U10768 (N_10768,N_10495,N_10353);
xnor U10769 (N_10769,N_10412,N_10029);
nor U10770 (N_10770,N_10202,N_10422);
and U10771 (N_10771,N_10049,N_10234);
xnor U10772 (N_10772,N_10388,N_10128);
and U10773 (N_10773,N_10466,N_10097);
or U10774 (N_10774,N_10187,N_10012);
xnor U10775 (N_10775,N_10422,N_10069);
nor U10776 (N_10776,N_10385,N_10437);
and U10777 (N_10777,N_10125,N_10197);
and U10778 (N_10778,N_10373,N_10056);
xnor U10779 (N_10779,N_10181,N_10462);
or U10780 (N_10780,N_10083,N_10065);
or U10781 (N_10781,N_10113,N_10435);
nand U10782 (N_10782,N_10414,N_10148);
and U10783 (N_10783,N_10458,N_10182);
nand U10784 (N_10784,N_10024,N_10263);
nand U10785 (N_10785,N_10118,N_10340);
and U10786 (N_10786,N_10177,N_10092);
or U10787 (N_10787,N_10441,N_10052);
and U10788 (N_10788,N_10352,N_10329);
or U10789 (N_10789,N_10279,N_10475);
or U10790 (N_10790,N_10438,N_10288);
nor U10791 (N_10791,N_10070,N_10491);
nor U10792 (N_10792,N_10348,N_10177);
xor U10793 (N_10793,N_10411,N_10461);
or U10794 (N_10794,N_10369,N_10270);
and U10795 (N_10795,N_10229,N_10210);
xnor U10796 (N_10796,N_10204,N_10363);
or U10797 (N_10797,N_10129,N_10294);
xor U10798 (N_10798,N_10352,N_10358);
and U10799 (N_10799,N_10434,N_10428);
nor U10800 (N_10800,N_10391,N_10119);
nor U10801 (N_10801,N_10267,N_10272);
nor U10802 (N_10802,N_10062,N_10331);
xnor U10803 (N_10803,N_10060,N_10146);
and U10804 (N_10804,N_10008,N_10199);
xor U10805 (N_10805,N_10383,N_10466);
nor U10806 (N_10806,N_10341,N_10029);
nor U10807 (N_10807,N_10397,N_10073);
xor U10808 (N_10808,N_10164,N_10025);
or U10809 (N_10809,N_10172,N_10350);
and U10810 (N_10810,N_10395,N_10387);
nand U10811 (N_10811,N_10156,N_10131);
or U10812 (N_10812,N_10202,N_10150);
and U10813 (N_10813,N_10221,N_10302);
nand U10814 (N_10814,N_10142,N_10485);
nor U10815 (N_10815,N_10109,N_10292);
or U10816 (N_10816,N_10490,N_10129);
xor U10817 (N_10817,N_10465,N_10250);
nor U10818 (N_10818,N_10222,N_10046);
and U10819 (N_10819,N_10286,N_10444);
nand U10820 (N_10820,N_10458,N_10253);
xor U10821 (N_10821,N_10218,N_10207);
xnor U10822 (N_10822,N_10071,N_10275);
or U10823 (N_10823,N_10059,N_10199);
and U10824 (N_10824,N_10091,N_10005);
and U10825 (N_10825,N_10354,N_10395);
nor U10826 (N_10826,N_10192,N_10388);
or U10827 (N_10827,N_10424,N_10290);
xor U10828 (N_10828,N_10026,N_10374);
nand U10829 (N_10829,N_10203,N_10227);
nand U10830 (N_10830,N_10148,N_10081);
nor U10831 (N_10831,N_10377,N_10131);
or U10832 (N_10832,N_10436,N_10208);
and U10833 (N_10833,N_10475,N_10282);
nand U10834 (N_10834,N_10347,N_10257);
nand U10835 (N_10835,N_10243,N_10480);
nor U10836 (N_10836,N_10084,N_10091);
and U10837 (N_10837,N_10301,N_10091);
and U10838 (N_10838,N_10369,N_10338);
xor U10839 (N_10839,N_10086,N_10017);
nor U10840 (N_10840,N_10467,N_10002);
nand U10841 (N_10841,N_10461,N_10153);
xor U10842 (N_10842,N_10456,N_10365);
or U10843 (N_10843,N_10453,N_10353);
or U10844 (N_10844,N_10293,N_10247);
or U10845 (N_10845,N_10395,N_10432);
and U10846 (N_10846,N_10196,N_10375);
xor U10847 (N_10847,N_10166,N_10144);
or U10848 (N_10848,N_10210,N_10089);
nand U10849 (N_10849,N_10087,N_10224);
or U10850 (N_10850,N_10317,N_10418);
xor U10851 (N_10851,N_10106,N_10183);
nor U10852 (N_10852,N_10129,N_10092);
or U10853 (N_10853,N_10166,N_10460);
nor U10854 (N_10854,N_10329,N_10094);
xnor U10855 (N_10855,N_10475,N_10074);
nand U10856 (N_10856,N_10151,N_10336);
nor U10857 (N_10857,N_10007,N_10018);
nor U10858 (N_10858,N_10357,N_10197);
and U10859 (N_10859,N_10265,N_10217);
nor U10860 (N_10860,N_10084,N_10156);
nor U10861 (N_10861,N_10045,N_10001);
nor U10862 (N_10862,N_10158,N_10164);
nand U10863 (N_10863,N_10073,N_10223);
or U10864 (N_10864,N_10449,N_10485);
xor U10865 (N_10865,N_10306,N_10490);
or U10866 (N_10866,N_10183,N_10004);
and U10867 (N_10867,N_10426,N_10420);
and U10868 (N_10868,N_10449,N_10308);
nand U10869 (N_10869,N_10013,N_10386);
nand U10870 (N_10870,N_10007,N_10030);
nor U10871 (N_10871,N_10268,N_10304);
or U10872 (N_10872,N_10327,N_10034);
or U10873 (N_10873,N_10481,N_10125);
or U10874 (N_10874,N_10466,N_10149);
and U10875 (N_10875,N_10332,N_10491);
and U10876 (N_10876,N_10002,N_10373);
or U10877 (N_10877,N_10127,N_10093);
nand U10878 (N_10878,N_10234,N_10120);
or U10879 (N_10879,N_10222,N_10204);
nor U10880 (N_10880,N_10105,N_10134);
or U10881 (N_10881,N_10215,N_10451);
or U10882 (N_10882,N_10477,N_10403);
nand U10883 (N_10883,N_10453,N_10280);
or U10884 (N_10884,N_10415,N_10270);
and U10885 (N_10885,N_10271,N_10443);
or U10886 (N_10886,N_10146,N_10244);
and U10887 (N_10887,N_10139,N_10441);
xnor U10888 (N_10888,N_10112,N_10299);
xor U10889 (N_10889,N_10164,N_10206);
xor U10890 (N_10890,N_10041,N_10238);
nand U10891 (N_10891,N_10364,N_10162);
nand U10892 (N_10892,N_10100,N_10403);
xor U10893 (N_10893,N_10395,N_10377);
nand U10894 (N_10894,N_10287,N_10186);
or U10895 (N_10895,N_10494,N_10300);
nor U10896 (N_10896,N_10297,N_10277);
nand U10897 (N_10897,N_10271,N_10051);
and U10898 (N_10898,N_10176,N_10051);
or U10899 (N_10899,N_10244,N_10070);
nor U10900 (N_10900,N_10107,N_10430);
nand U10901 (N_10901,N_10067,N_10378);
nand U10902 (N_10902,N_10277,N_10133);
nand U10903 (N_10903,N_10129,N_10467);
nor U10904 (N_10904,N_10433,N_10274);
nand U10905 (N_10905,N_10238,N_10177);
and U10906 (N_10906,N_10499,N_10335);
or U10907 (N_10907,N_10257,N_10365);
nor U10908 (N_10908,N_10092,N_10104);
nor U10909 (N_10909,N_10284,N_10017);
nand U10910 (N_10910,N_10122,N_10104);
xor U10911 (N_10911,N_10273,N_10128);
or U10912 (N_10912,N_10436,N_10090);
and U10913 (N_10913,N_10247,N_10190);
or U10914 (N_10914,N_10117,N_10025);
xnor U10915 (N_10915,N_10101,N_10496);
nor U10916 (N_10916,N_10082,N_10179);
xnor U10917 (N_10917,N_10361,N_10256);
nand U10918 (N_10918,N_10006,N_10269);
or U10919 (N_10919,N_10192,N_10290);
nor U10920 (N_10920,N_10156,N_10394);
nor U10921 (N_10921,N_10049,N_10073);
nor U10922 (N_10922,N_10492,N_10472);
nand U10923 (N_10923,N_10343,N_10344);
nand U10924 (N_10924,N_10137,N_10152);
or U10925 (N_10925,N_10062,N_10384);
nor U10926 (N_10926,N_10286,N_10431);
nand U10927 (N_10927,N_10295,N_10388);
and U10928 (N_10928,N_10111,N_10312);
nand U10929 (N_10929,N_10115,N_10052);
and U10930 (N_10930,N_10172,N_10417);
xnor U10931 (N_10931,N_10020,N_10087);
xnor U10932 (N_10932,N_10104,N_10460);
nor U10933 (N_10933,N_10313,N_10449);
and U10934 (N_10934,N_10445,N_10451);
or U10935 (N_10935,N_10357,N_10330);
nor U10936 (N_10936,N_10161,N_10198);
and U10937 (N_10937,N_10181,N_10025);
nand U10938 (N_10938,N_10293,N_10213);
nand U10939 (N_10939,N_10002,N_10391);
and U10940 (N_10940,N_10328,N_10019);
and U10941 (N_10941,N_10294,N_10186);
nand U10942 (N_10942,N_10203,N_10398);
or U10943 (N_10943,N_10452,N_10489);
nand U10944 (N_10944,N_10030,N_10298);
xor U10945 (N_10945,N_10237,N_10376);
xor U10946 (N_10946,N_10335,N_10320);
nand U10947 (N_10947,N_10065,N_10396);
nand U10948 (N_10948,N_10315,N_10056);
xnor U10949 (N_10949,N_10260,N_10189);
or U10950 (N_10950,N_10309,N_10048);
nor U10951 (N_10951,N_10024,N_10002);
nand U10952 (N_10952,N_10242,N_10182);
or U10953 (N_10953,N_10019,N_10246);
nand U10954 (N_10954,N_10249,N_10388);
nand U10955 (N_10955,N_10151,N_10243);
xor U10956 (N_10956,N_10065,N_10070);
nor U10957 (N_10957,N_10255,N_10008);
or U10958 (N_10958,N_10041,N_10202);
or U10959 (N_10959,N_10189,N_10326);
xnor U10960 (N_10960,N_10497,N_10474);
or U10961 (N_10961,N_10239,N_10412);
and U10962 (N_10962,N_10060,N_10110);
nor U10963 (N_10963,N_10268,N_10360);
nand U10964 (N_10964,N_10074,N_10126);
and U10965 (N_10965,N_10296,N_10382);
nand U10966 (N_10966,N_10261,N_10253);
xor U10967 (N_10967,N_10339,N_10372);
or U10968 (N_10968,N_10207,N_10301);
and U10969 (N_10969,N_10054,N_10228);
nand U10970 (N_10970,N_10224,N_10480);
nand U10971 (N_10971,N_10390,N_10353);
nor U10972 (N_10972,N_10054,N_10367);
nand U10973 (N_10973,N_10460,N_10144);
and U10974 (N_10974,N_10124,N_10323);
xnor U10975 (N_10975,N_10322,N_10415);
nand U10976 (N_10976,N_10491,N_10182);
xnor U10977 (N_10977,N_10496,N_10459);
and U10978 (N_10978,N_10491,N_10163);
xor U10979 (N_10979,N_10131,N_10175);
nand U10980 (N_10980,N_10201,N_10211);
and U10981 (N_10981,N_10246,N_10159);
nor U10982 (N_10982,N_10239,N_10083);
nand U10983 (N_10983,N_10002,N_10275);
or U10984 (N_10984,N_10399,N_10110);
or U10985 (N_10985,N_10138,N_10492);
xnor U10986 (N_10986,N_10173,N_10494);
or U10987 (N_10987,N_10116,N_10141);
nor U10988 (N_10988,N_10234,N_10153);
xnor U10989 (N_10989,N_10484,N_10167);
nand U10990 (N_10990,N_10288,N_10358);
nand U10991 (N_10991,N_10378,N_10055);
nand U10992 (N_10992,N_10136,N_10368);
and U10993 (N_10993,N_10080,N_10059);
and U10994 (N_10994,N_10270,N_10155);
or U10995 (N_10995,N_10222,N_10244);
and U10996 (N_10996,N_10168,N_10124);
or U10997 (N_10997,N_10034,N_10019);
xor U10998 (N_10998,N_10235,N_10464);
nor U10999 (N_10999,N_10414,N_10486);
nand U11000 (N_11000,N_10963,N_10567);
xor U11001 (N_11001,N_10537,N_10545);
nor U11002 (N_11002,N_10588,N_10548);
nand U11003 (N_11003,N_10500,N_10968);
nand U11004 (N_11004,N_10656,N_10584);
nor U11005 (N_11005,N_10531,N_10877);
nor U11006 (N_11006,N_10648,N_10789);
xor U11007 (N_11007,N_10654,N_10939);
nand U11008 (N_11008,N_10842,N_10521);
and U11009 (N_11009,N_10884,N_10989);
nand U11010 (N_11010,N_10611,N_10909);
nand U11011 (N_11011,N_10976,N_10730);
nor U11012 (N_11012,N_10686,N_10755);
or U11013 (N_11013,N_10946,N_10724);
or U11014 (N_11014,N_10979,N_10625);
xnor U11015 (N_11015,N_10536,N_10514);
or U11016 (N_11016,N_10661,N_10636);
nand U11017 (N_11017,N_10763,N_10922);
xor U11018 (N_11018,N_10704,N_10703);
nor U11019 (N_11019,N_10809,N_10746);
nand U11020 (N_11020,N_10830,N_10882);
and U11021 (N_11021,N_10549,N_10699);
or U11022 (N_11022,N_10762,N_10639);
and U11023 (N_11023,N_10702,N_10624);
nor U11024 (N_11024,N_10538,N_10794);
nand U11025 (N_11025,N_10660,N_10953);
nand U11026 (N_11026,N_10838,N_10714);
xnor U11027 (N_11027,N_10700,N_10541);
or U11028 (N_11028,N_10655,N_10859);
xor U11029 (N_11029,N_10834,N_10621);
nand U11030 (N_11030,N_10959,N_10994);
or U11031 (N_11031,N_10582,N_10825);
and U11032 (N_11032,N_10677,N_10863);
nand U11033 (N_11033,N_10592,N_10681);
or U11034 (N_11034,N_10561,N_10965);
xnor U11035 (N_11035,N_10650,N_10964);
or U11036 (N_11036,N_10568,N_10733);
xor U11037 (N_11037,N_10982,N_10504);
nor U11038 (N_11038,N_10908,N_10605);
or U11039 (N_11039,N_10669,N_10855);
and U11040 (N_11040,N_10555,N_10969);
nand U11041 (N_11041,N_10898,N_10716);
nor U11042 (N_11042,N_10958,N_10515);
xnor U11043 (N_11043,N_10607,N_10528);
nand U11044 (N_11044,N_10552,N_10786);
xor U11045 (N_11045,N_10623,N_10657);
or U11046 (N_11046,N_10576,N_10543);
and U11047 (N_11047,N_10807,N_10742);
nor U11048 (N_11048,N_10617,N_10516);
xnor U11049 (N_11049,N_10858,N_10803);
nand U11050 (N_11050,N_10868,N_10950);
nand U11051 (N_11051,N_10764,N_10943);
and U11052 (N_11052,N_10851,N_10894);
or U11053 (N_11053,N_10634,N_10784);
nor U11054 (N_11054,N_10826,N_10823);
nand U11055 (N_11055,N_10659,N_10772);
nand U11056 (N_11056,N_10542,N_10673);
or U11057 (N_11057,N_10983,N_10525);
xnor U11058 (N_11058,N_10577,N_10523);
nand U11059 (N_11059,N_10881,N_10684);
nand U11060 (N_11060,N_10885,N_10915);
nand U11061 (N_11061,N_10988,N_10749);
nand U11062 (N_11062,N_10539,N_10866);
nor U11063 (N_11063,N_10613,N_10864);
and U11064 (N_11064,N_10569,N_10619);
or U11065 (N_11065,N_10741,N_10903);
xnor U11066 (N_11066,N_10596,N_10805);
nand U11067 (N_11067,N_10574,N_10916);
xor U11068 (N_11068,N_10604,N_10771);
nor U11069 (N_11069,N_10731,N_10853);
or U11070 (N_11070,N_10783,N_10776);
xor U11071 (N_11071,N_10532,N_10601);
nor U11072 (N_11072,N_10902,N_10770);
and U11073 (N_11073,N_10573,N_10978);
and U11074 (N_11074,N_10759,N_10986);
and U11075 (N_11075,N_10641,N_10896);
or U11076 (N_11076,N_10630,N_10706);
or U11077 (N_11077,N_10768,N_10682);
xor U11078 (N_11078,N_10737,N_10757);
nand U11079 (N_11079,N_10558,N_10690);
nor U11080 (N_11080,N_10937,N_10527);
and U11081 (N_11081,N_10705,N_10678);
xor U11082 (N_11082,N_10869,N_10729);
and U11083 (N_11083,N_10519,N_10529);
nor U11084 (N_11084,N_10696,N_10880);
nor U11085 (N_11085,N_10980,N_10775);
nor U11086 (N_11086,N_10725,N_10886);
or U11087 (N_11087,N_10591,N_10740);
and U11088 (N_11088,N_10874,N_10565);
and U11089 (N_11089,N_10754,N_10698);
or U11090 (N_11090,N_10791,N_10919);
nor U11091 (N_11091,N_10649,N_10918);
xor U11092 (N_11092,N_10629,N_10945);
nand U11093 (N_11093,N_10839,N_10872);
xor U11094 (N_11094,N_10887,N_10815);
nor U11095 (N_11095,N_10998,N_10674);
or U11096 (N_11096,N_10713,N_10895);
nand U11097 (N_11097,N_10665,N_10511);
or U11098 (N_11098,N_10793,N_10712);
xor U11099 (N_11099,N_10873,N_10972);
and U11100 (N_11100,N_10942,N_10966);
and U11101 (N_11101,N_10501,N_10824);
nand U11102 (N_11102,N_10897,N_10813);
or U11103 (N_11103,N_10828,N_10888);
nand U11104 (N_11104,N_10981,N_10554);
nor U11105 (N_11105,N_10638,N_10721);
xnor U11106 (N_11106,N_10645,N_10810);
or U11107 (N_11107,N_10556,N_10910);
xnor U11108 (N_11108,N_10688,N_10760);
nor U11109 (N_11109,N_10540,N_10782);
nor U11110 (N_11110,N_10871,N_10914);
nand U11111 (N_11111,N_10883,N_10564);
nor U11112 (N_11112,N_10879,N_10788);
or U11113 (N_11113,N_10583,N_10854);
xnor U11114 (N_11114,N_10701,N_10522);
and U11115 (N_11115,N_10827,N_10820);
nand U11116 (N_11116,N_10751,N_10808);
or U11117 (N_11117,N_10557,N_10736);
xnor U11118 (N_11118,N_10819,N_10923);
and U11119 (N_11119,N_10683,N_10679);
xnor U11120 (N_11120,N_10753,N_10550);
nand U11121 (N_11121,N_10995,N_10610);
or U11122 (N_11122,N_10961,N_10628);
xnor U11123 (N_11123,N_10812,N_10637);
and U11124 (N_11124,N_10547,N_10503);
and U11125 (N_11125,N_10920,N_10814);
or U11126 (N_11126,N_10671,N_10818);
and U11127 (N_11127,N_10856,N_10780);
and U11128 (N_11128,N_10925,N_10620);
nand U11129 (N_11129,N_10921,N_10798);
nor U11130 (N_11130,N_10892,N_10672);
nand U11131 (N_11131,N_10860,N_10773);
or U11132 (N_11132,N_10640,N_10750);
and U11133 (N_11133,N_10734,N_10710);
nor U11134 (N_11134,N_10692,N_10912);
nor U11135 (N_11135,N_10546,N_10840);
or U11136 (N_11136,N_10662,N_10935);
or U11137 (N_11137,N_10796,N_10951);
or U11138 (N_11138,N_10695,N_10831);
xor U11139 (N_11139,N_10586,N_10534);
nand U11140 (N_11140,N_10580,N_10572);
or U11141 (N_11141,N_10829,N_10956);
nand U11142 (N_11142,N_10551,N_10571);
nand U11143 (N_11143,N_10595,N_10520);
or U11144 (N_11144,N_10934,N_10930);
nand U11145 (N_11145,N_10594,N_10949);
nand U11146 (N_11146,N_10837,N_10985);
or U11147 (N_11147,N_10779,N_10926);
xor U11148 (N_11148,N_10924,N_10901);
and U11149 (N_11149,N_10728,N_10835);
or U11150 (N_11150,N_10990,N_10893);
nor U11151 (N_11151,N_10857,N_10785);
xor U11152 (N_11152,N_10526,N_10590);
nor U11153 (N_11153,N_10752,N_10954);
nand U11154 (N_11154,N_10744,N_10570);
or U11155 (N_11155,N_10867,N_10875);
and U11156 (N_11156,N_10562,N_10761);
and U11157 (N_11157,N_10606,N_10566);
xor U11158 (N_11158,N_10797,N_10693);
or U11159 (N_11159,N_10502,N_10651);
nor U11160 (N_11160,N_10599,N_10900);
xnor U11161 (N_11161,N_10533,N_10646);
or U11162 (N_11162,N_10781,N_10685);
nand U11163 (N_11163,N_10579,N_10553);
xor U11164 (N_11164,N_10518,N_10747);
and U11165 (N_11165,N_10609,N_10585);
and U11166 (N_11166,N_10849,N_10563);
or U11167 (N_11167,N_10769,N_10913);
and U11168 (N_11168,N_10974,N_10932);
xor U11169 (N_11169,N_10598,N_10627);
or U11170 (N_11170,N_10722,N_10844);
nor U11171 (N_11171,N_10952,N_10984);
and U11172 (N_11172,N_10633,N_10929);
xor U11173 (N_11173,N_10689,N_10708);
nor U11174 (N_11174,N_10711,N_10664);
or U11175 (N_11175,N_10847,N_10836);
nand U11176 (N_11176,N_10970,N_10512);
xor U11177 (N_11177,N_10524,N_10719);
and U11178 (N_11178,N_10559,N_10967);
nand U11179 (N_11179,N_10732,N_10774);
nand U11180 (N_11180,N_10643,N_10944);
nor U11181 (N_11181,N_10632,N_10928);
and U11182 (N_11182,N_10991,N_10992);
nand U11183 (N_11183,N_10756,N_10668);
or U11184 (N_11184,N_10635,N_10841);
or U11185 (N_11185,N_10581,N_10971);
and U11186 (N_11186,N_10631,N_10941);
and U11187 (N_11187,N_10707,N_10890);
or U11188 (N_11188,N_10626,N_10603);
xnor U11189 (N_11189,N_10911,N_10653);
nor U11190 (N_11190,N_10999,N_10962);
or U11191 (N_11191,N_10777,N_10906);
and U11192 (N_11192,N_10765,N_10767);
and U11193 (N_11193,N_10938,N_10720);
nand U11194 (N_11194,N_10622,N_10723);
and U11195 (N_11195,N_10589,N_10667);
and U11196 (N_11196,N_10670,N_10506);
nor U11197 (N_11197,N_10821,N_10933);
xor U11198 (N_11198,N_10587,N_10865);
xnor U11199 (N_11199,N_10878,N_10644);
or U11200 (N_11200,N_10709,N_10993);
nand U11201 (N_11201,N_10832,N_10870);
xnor U11202 (N_11202,N_10848,N_10697);
and U11203 (N_11203,N_10616,N_10578);
nand U11204 (N_11204,N_10694,N_10822);
xor U11205 (N_11205,N_10852,N_10955);
or U11206 (N_11206,N_10597,N_10801);
and U11207 (N_11207,N_10904,N_10530);
nor U11208 (N_11208,N_10975,N_10680);
nor U11209 (N_11209,N_10715,N_10739);
and U11210 (N_11210,N_10743,N_10735);
and U11211 (N_11211,N_10927,N_10996);
nor U11212 (N_11212,N_10766,N_10726);
or U11213 (N_11213,N_10727,N_10917);
nand U11214 (N_11214,N_10799,N_10899);
nand U11215 (N_11215,N_10987,N_10652);
nand U11216 (N_11216,N_10560,N_10618);
xor U11217 (N_11217,N_10612,N_10608);
nor U11218 (N_11218,N_10843,N_10931);
and U11219 (N_11219,N_10748,N_10505);
and U11220 (N_11220,N_10507,N_10907);
nand U11221 (N_11221,N_10948,N_10997);
nand U11222 (N_11222,N_10614,N_10675);
nand U11223 (N_11223,N_10745,N_10889);
nand U11224 (N_11224,N_10802,N_10936);
and U11225 (N_11225,N_10508,N_10891);
and U11226 (N_11226,N_10787,N_10658);
nor U11227 (N_11227,N_10666,N_10811);
nor U11228 (N_11228,N_10544,N_10513);
or U11229 (N_11229,N_10816,N_10861);
nand U11230 (N_11230,N_10977,N_10800);
or U11231 (N_11231,N_10804,N_10509);
or U11232 (N_11232,N_10676,N_10510);
nor U11233 (N_11233,N_10602,N_10973);
or U11234 (N_11234,N_10517,N_10758);
nand U11235 (N_11235,N_10940,N_10600);
xnor U11236 (N_11236,N_10905,N_10642);
and U11237 (N_11237,N_10833,N_10960);
nor U11238 (N_11238,N_10663,N_10738);
xor U11239 (N_11239,N_10795,N_10615);
nor U11240 (N_11240,N_10957,N_10862);
nand U11241 (N_11241,N_10778,N_10718);
or U11242 (N_11242,N_10876,N_10806);
and U11243 (N_11243,N_10792,N_10717);
nand U11244 (N_11244,N_10535,N_10687);
nor U11245 (N_11245,N_10845,N_10846);
or U11246 (N_11246,N_10850,N_10790);
nand U11247 (N_11247,N_10593,N_10575);
or U11248 (N_11248,N_10691,N_10947);
nand U11249 (N_11249,N_10647,N_10817);
nand U11250 (N_11250,N_10554,N_10809);
or U11251 (N_11251,N_10515,N_10890);
nand U11252 (N_11252,N_10847,N_10700);
xnor U11253 (N_11253,N_10961,N_10957);
nor U11254 (N_11254,N_10742,N_10736);
nand U11255 (N_11255,N_10690,N_10932);
nor U11256 (N_11256,N_10757,N_10744);
nand U11257 (N_11257,N_10841,N_10784);
and U11258 (N_11258,N_10692,N_10744);
or U11259 (N_11259,N_10530,N_10865);
nand U11260 (N_11260,N_10761,N_10753);
or U11261 (N_11261,N_10985,N_10894);
nand U11262 (N_11262,N_10834,N_10753);
xor U11263 (N_11263,N_10711,N_10667);
xnor U11264 (N_11264,N_10821,N_10785);
or U11265 (N_11265,N_10968,N_10733);
and U11266 (N_11266,N_10891,N_10573);
nor U11267 (N_11267,N_10527,N_10758);
nor U11268 (N_11268,N_10837,N_10594);
and U11269 (N_11269,N_10502,N_10943);
nor U11270 (N_11270,N_10566,N_10841);
nor U11271 (N_11271,N_10730,N_10582);
nand U11272 (N_11272,N_10525,N_10779);
nor U11273 (N_11273,N_10730,N_10984);
or U11274 (N_11274,N_10742,N_10952);
xor U11275 (N_11275,N_10919,N_10611);
nand U11276 (N_11276,N_10723,N_10801);
or U11277 (N_11277,N_10576,N_10636);
nand U11278 (N_11278,N_10760,N_10894);
and U11279 (N_11279,N_10566,N_10993);
and U11280 (N_11280,N_10731,N_10855);
and U11281 (N_11281,N_10780,N_10582);
xor U11282 (N_11282,N_10667,N_10892);
and U11283 (N_11283,N_10950,N_10569);
nor U11284 (N_11284,N_10800,N_10638);
or U11285 (N_11285,N_10924,N_10915);
and U11286 (N_11286,N_10509,N_10891);
or U11287 (N_11287,N_10787,N_10596);
xnor U11288 (N_11288,N_10783,N_10561);
nand U11289 (N_11289,N_10738,N_10513);
nor U11290 (N_11290,N_10782,N_10545);
xor U11291 (N_11291,N_10612,N_10710);
and U11292 (N_11292,N_10776,N_10739);
or U11293 (N_11293,N_10548,N_10975);
and U11294 (N_11294,N_10849,N_10896);
nand U11295 (N_11295,N_10913,N_10603);
xnor U11296 (N_11296,N_10978,N_10734);
and U11297 (N_11297,N_10838,N_10810);
or U11298 (N_11298,N_10691,N_10924);
and U11299 (N_11299,N_10939,N_10971);
nor U11300 (N_11300,N_10748,N_10953);
nor U11301 (N_11301,N_10781,N_10655);
nand U11302 (N_11302,N_10773,N_10840);
and U11303 (N_11303,N_10728,N_10556);
and U11304 (N_11304,N_10544,N_10965);
nand U11305 (N_11305,N_10747,N_10618);
nor U11306 (N_11306,N_10873,N_10516);
nand U11307 (N_11307,N_10918,N_10809);
or U11308 (N_11308,N_10608,N_10645);
xor U11309 (N_11309,N_10741,N_10558);
nor U11310 (N_11310,N_10524,N_10666);
xnor U11311 (N_11311,N_10779,N_10825);
nand U11312 (N_11312,N_10950,N_10775);
nor U11313 (N_11313,N_10648,N_10821);
or U11314 (N_11314,N_10619,N_10895);
nor U11315 (N_11315,N_10613,N_10909);
xnor U11316 (N_11316,N_10980,N_10581);
nor U11317 (N_11317,N_10630,N_10850);
or U11318 (N_11318,N_10756,N_10859);
nor U11319 (N_11319,N_10575,N_10917);
nand U11320 (N_11320,N_10522,N_10705);
nand U11321 (N_11321,N_10672,N_10792);
and U11322 (N_11322,N_10510,N_10937);
xnor U11323 (N_11323,N_10588,N_10580);
xnor U11324 (N_11324,N_10624,N_10812);
nor U11325 (N_11325,N_10601,N_10763);
nor U11326 (N_11326,N_10743,N_10546);
xnor U11327 (N_11327,N_10828,N_10865);
and U11328 (N_11328,N_10967,N_10982);
or U11329 (N_11329,N_10819,N_10869);
nand U11330 (N_11330,N_10970,N_10722);
nand U11331 (N_11331,N_10517,N_10514);
or U11332 (N_11332,N_10743,N_10941);
or U11333 (N_11333,N_10855,N_10576);
and U11334 (N_11334,N_10955,N_10778);
nor U11335 (N_11335,N_10635,N_10616);
or U11336 (N_11336,N_10690,N_10731);
nor U11337 (N_11337,N_10509,N_10731);
or U11338 (N_11338,N_10758,N_10685);
or U11339 (N_11339,N_10652,N_10828);
or U11340 (N_11340,N_10703,N_10707);
xor U11341 (N_11341,N_10763,N_10895);
or U11342 (N_11342,N_10638,N_10576);
and U11343 (N_11343,N_10982,N_10706);
xor U11344 (N_11344,N_10580,N_10917);
nor U11345 (N_11345,N_10720,N_10755);
xor U11346 (N_11346,N_10950,N_10587);
nand U11347 (N_11347,N_10748,N_10586);
nand U11348 (N_11348,N_10589,N_10982);
and U11349 (N_11349,N_10820,N_10822);
or U11350 (N_11350,N_10622,N_10867);
or U11351 (N_11351,N_10518,N_10658);
and U11352 (N_11352,N_10638,N_10665);
and U11353 (N_11353,N_10846,N_10557);
nor U11354 (N_11354,N_10677,N_10659);
nand U11355 (N_11355,N_10606,N_10946);
and U11356 (N_11356,N_10767,N_10894);
xor U11357 (N_11357,N_10623,N_10567);
and U11358 (N_11358,N_10955,N_10602);
or U11359 (N_11359,N_10801,N_10839);
and U11360 (N_11360,N_10735,N_10935);
and U11361 (N_11361,N_10976,N_10969);
and U11362 (N_11362,N_10508,N_10611);
xor U11363 (N_11363,N_10953,N_10872);
or U11364 (N_11364,N_10597,N_10769);
and U11365 (N_11365,N_10549,N_10653);
xnor U11366 (N_11366,N_10612,N_10992);
and U11367 (N_11367,N_10727,N_10843);
nand U11368 (N_11368,N_10988,N_10936);
nand U11369 (N_11369,N_10936,N_10947);
and U11370 (N_11370,N_10907,N_10541);
nand U11371 (N_11371,N_10887,N_10657);
and U11372 (N_11372,N_10652,N_10628);
xnor U11373 (N_11373,N_10925,N_10795);
nor U11374 (N_11374,N_10625,N_10505);
xor U11375 (N_11375,N_10611,N_10968);
xor U11376 (N_11376,N_10529,N_10637);
nor U11377 (N_11377,N_10628,N_10849);
or U11378 (N_11378,N_10599,N_10929);
and U11379 (N_11379,N_10887,N_10709);
or U11380 (N_11380,N_10916,N_10983);
xnor U11381 (N_11381,N_10543,N_10661);
or U11382 (N_11382,N_10691,N_10610);
nor U11383 (N_11383,N_10766,N_10684);
xor U11384 (N_11384,N_10584,N_10984);
nor U11385 (N_11385,N_10738,N_10512);
xnor U11386 (N_11386,N_10569,N_10599);
nor U11387 (N_11387,N_10822,N_10505);
nor U11388 (N_11388,N_10903,N_10935);
xor U11389 (N_11389,N_10503,N_10880);
nand U11390 (N_11390,N_10813,N_10792);
and U11391 (N_11391,N_10670,N_10631);
nor U11392 (N_11392,N_10504,N_10797);
nand U11393 (N_11393,N_10899,N_10734);
nor U11394 (N_11394,N_10733,N_10898);
xnor U11395 (N_11395,N_10768,N_10870);
or U11396 (N_11396,N_10648,N_10658);
nor U11397 (N_11397,N_10983,N_10633);
nand U11398 (N_11398,N_10510,N_10609);
or U11399 (N_11399,N_10726,N_10903);
and U11400 (N_11400,N_10678,N_10632);
xor U11401 (N_11401,N_10938,N_10644);
nor U11402 (N_11402,N_10725,N_10998);
nand U11403 (N_11403,N_10641,N_10597);
nand U11404 (N_11404,N_10991,N_10692);
and U11405 (N_11405,N_10727,N_10756);
nand U11406 (N_11406,N_10505,N_10717);
nand U11407 (N_11407,N_10683,N_10871);
and U11408 (N_11408,N_10620,N_10537);
or U11409 (N_11409,N_10831,N_10871);
or U11410 (N_11410,N_10621,N_10620);
xor U11411 (N_11411,N_10692,N_10769);
and U11412 (N_11412,N_10530,N_10564);
or U11413 (N_11413,N_10551,N_10960);
nand U11414 (N_11414,N_10811,N_10950);
nand U11415 (N_11415,N_10900,N_10720);
or U11416 (N_11416,N_10530,N_10607);
or U11417 (N_11417,N_10554,N_10836);
and U11418 (N_11418,N_10791,N_10644);
nor U11419 (N_11419,N_10889,N_10540);
xor U11420 (N_11420,N_10533,N_10603);
nor U11421 (N_11421,N_10751,N_10973);
xnor U11422 (N_11422,N_10516,N_10653);
nor U11423 (N_11423,N_10908,N_10699);
nand U11424 (N_11424,N_10988,N_10657);
xnor U11425 (N_11425,N_10772,N_10971);
nand U11426 (N_11426,N_10759,N_10990);
or U11427 (N_11427,N_10919,N_10713);
xnor U11428 (N_11428,N_10773,N_10624);
nor U11429 (N_11429,N_10761,N_10905);
and U11430 (N_11430,N_10707,N_10962);
nor U11431 (N_11431,N_10893,N_10607);
xnor U11432 (N_11432,N_10983,N_10893);
nand U11433 (N_11433,N_10956,N_10578);
xnor U11434 (N_11434,N_10811,N_10897);
and U11435 (N_11435,N_10796,N_10741);
or U11436 (N_11436,N_10799,N_10947);
nor U11437 (N_11437,N_10638,N_10814);
xnor U11438 (N_11438,N_10940,N_10617);
nor U11439 (N_11439,N_10666,N_10828);
and U11440 (N_11440,N_10606,N_10696);
and U11441 (N_11441,N_10678,N_10520);
nand U11442 (N_11442,N_10735,N_10981);
and U11443 (N_11443,N_10873,N_10632);
nand U11444 (N_11444,N_10553,N_10969);
or U11445 (N_11445,N_10506,N_10843);
xnor U11446 (N_11446,N_10889,N_10797);
nor U11447 (N_11447,N_10640,N_10769);
xor U11448 (N_11448,N_10905,N_10552);
or U11449 (N_11449,N_10692,N_10609);
xor U11450 (N_11450,N_10987,N_10953);
xnor U11451 (N_11451,N_10999,N_10565);
and U11452 (N_11452,N_10839,N_10754);
xnor U11453 (N_11453,N_10821,N_10670);
xor U11454 (N_11454,N_10586,N_10892);
or U11455 (N_11455,N_10867,N_10523);
nand U11456 (N_11456,N_10909,N_10648);
nor U11457 (N_11457,N_10712,N_10675);
and U11458 (N_11458,N_10952,N_10547);
nand U11459 (N_11459,N_10527,N_10860);
or U11460 (N_11460,N_10574,N_10972);
and U11461 (N_11461,N_10891,N_10533);
and U11462 (N_11462,N_10681,N_10585);
xor U11463 (N_11463,N_10631,N_10503);
and U11464 (N_11464,N_10857,N_10964);
nor U11465 (N_11465,N_10942,N_10731);
nor U11466 (N_11466,N_10905,N_10823);
or U11467 (N_11467,N_10627,N_10951);
nor U11468 (N_11468,N_10541,N_10790);
xor U11469 (N_11469,N_10812,N_10941);
nand U11470 (N_11470,N_10602,N_10816);
and U11471 (N_11471,N_10755,N_10862);
or U11472 (N_11472,N_10928,N_10660);
or U11473 (N_11473,N_10840,N_10921);
nand U11474 (N_11474,N_10712,N_10936);
and U11475 (N_11475,N_10691,N_10871);
or U11476 (N_11476,N_10707,N_10807);
or U11477 (N_11477,N_10870,N_10978);
nor U11478 (N_11478,N_10783,N_10653);
nor U11479 (N_11479,N_10987,N_10672);
and U11480 (N_11480,N_10704,N_10599);
or U11481 (N_11481,N_10592,N_10851);
or U11482 (N_11482,N_10629,N_10714);
nor U11483 (N_11483,N_10674,N_10793);
and U11484 (N_11484,N_10888,N_10565);
xor U11485 (N_11485,N_10667,N_10871);
nor U11486 (N_11486,N_10581,N_10703);
or U11487 (N_11487,N_10833,N_10558);
xnor U11488 (N_11488,N_10704,N_10789);
and U11489 (N_11489,N_10983,N_10905);
nand U11490 (N_11490,N_10685,N_10811);
and U11491 (N_11491,N_10723,N_10833);
nand U11492 (N_11492,N_10765,N_10738);
or U11493 (N_11493,N_10693,N_10853);
nand U11494 (N_11494,N_10789,N_10773);
nand U11495 (N_11495,N_10814,N_10970);
nor U11496 (N_11496,N_10889,N_10545);
nand U11497 (N_11497,N_10997,N_10593);
or U11498 (N_11498,N_10909,N_10878);
nand U11499 (N_11499,N_10707,N_10671);
nor U11500 (N_11500,N_11436,N_11143);
or U11501 (N_11501,N_11356,N_11403);
xnor U11502 (N_11502,N_11429,N_11337);
nor U11503 (N_11503,N_11102,N_11407);
nand U11504 (N_11504,N_11409,N_11112);
nand U11505 (N_11505,N_11258,N_11274);
nor U11506 (N_11506,N_11267,N_11304);
xor U11507 (N_11507,N_11485,N_11362);
nand U11508 (N_11508,N_11192,N_11217);
xnor U11509 (N_11509,N_11423,N_11248);
or U11510 (N_11510,N_11284,N_11059);
and U11511 (N_11511,N_11153,N_11052);
or U11512 (N_11512,N_11493,N_11074);
xor U11513 (N_11513,N_11213,N_11032);
or U11514 (N_11514,N_11378,N_11061);
nand U11515 (N_11515,N_11463,N_11397);
and U11516 (N_11516,N_11374,N_11176);
and U11517 (N_11517,N_11308,N_11431);
nand U11518 (N_11518,N_11370,N_11168);
and U11519 (N_11519,N_11413,N_11218);
and U11520 (N_11520,N_11044,N_11490);
nor U11521 (N_11521,N_11132,N_11279);
and U11522 (N_11522,N_11442,N_11247);
or U11523 (N_11523,N_11263,N_11345);
nor U11524 (N_11524,N_11329,N_11161);
nor U11525 (N_11525,N_11088,N_11380);
xor U11526 (N_11526,N_11177,N_11483);
nand U11527 (N_11527,N_11474,N_11203);
nor U11528 (N_11528,N_11195,N_11300);
or U11529 (N_11529,N_11410,N_11243);
nor U11530 (N_11530,N_11198,N_11072);
or U11531 (N_11531,N_11441,N_11317);
nand U11532 (N_11532,N_11424,N_11487);
xor U11533 (N_11533,N_11219,N_11053);
nor U11534 (N_11534,N_11259,N_11125);
nand U11535 (N_11535,N_11037,N_11376);
xnor U11536 (N_11536,N_11012,N_11349);
and U11537 (N_11537,N_11173,N_11361);
nor U11538 (N_11538,N_11149,N_11309);
nor U11539 (N_11539,N_11253,N_11164);
and U11540 (N_11540,N_11470,N_11367);
and U11541 (N_11541,N_11294,N_11202);
or U11542 (N_11542,N_11138,N_11034);
or U11543 (N_11543,N_11462,N_11426);
or U11544 (N_11544,N_11447,N_11341);
xnor U11545 (N_11545,N_11301,N_11001);
or U11546 (N_11546,N_11049,N_11150);
or U11547 (N_11547,N_11172,N_11136);
nand U11548 (N_11548,N_11127,N_11122);
nand U11549 (N_11549,N_11120,N_11295);
xor U11550 (N_11550,N_11414,N_11231);
xnor U11551 (N_11551,N_11326,N_11481);
or U11552 (N_11552,N_11244,N_11098);
and U11553 (N_11553,N_11291,N_11196);
or U11554 (N_11554,N_11316,N_11346);
nand U11555 (N_11555,N_11009,N_11446);
or U11556 (N_11556,N_11359,N_11338);
or U11557 (N_11557,N_11273,N_11265);
and U11558 (N_11558,N_11392,N_11223);
nand U11559 (N_11559,N_11352,N_11070);
or U11560 (N_11560,N_11420,N_11113);
or U11561 (N_11561,N_11031,N_11347);
and U11562 (N_11562,N_11369,N_11178);
xnor U11563 (N_11563,N_11323,N_11236);
and U11564 (N_11564,N_11353,N_11108);
nor U11565 (N_11565,N_11110,N_11327);
nor U11566 (N_11566,N_11118,N_11254);
nor U11567 (N_11567,N_11461,N_11030);
nand U11568 (N_11568,N_11180,N_11473);
and U11569 (N_11569,N_11408,N_11303);
nand U11570 (N_11570,N_11205,N_11241);
nor U11571 (N_11571,N_11038,N_11078);
or U11572 (N_11572,N_11068,N_11250);
or U11573 (N_11573,N_11277,N_11114);
nand U11574 (N_11574,N_11499,N_11107);
nor U11575 (N_11575,N_11008,N_11175);
and U11576 (N_11576,N_11307,N_11228);
and U11577 (N_11577,N_11421,N_11268);
nor U11578 (N_11578,N_11073,N_11024);
and U11579 (N_11579,N_11233,N_11046);
and U11580 (N_11580,N_11182,N_11451);
nor U11581 (N_11581,N_11146,N_11290);
nand U11582 (N_11582,N_11390,N_11297);
or U11583 (N_11583,N_11375,N_11283);
xnor U11584 (N_11584,N_11459,N_11453);
and U11585 (N_11585,N_11472,N_11324);
and U11586 (N_11586,N_11210,N_11251);
xor U11587 (N_11587,N_11235,N_11054);
nor U11588 (N_11588,N_11045,N_11402);
and U11589 (N_11589,N_11147,N_11366);
nand U11590 (N_11590,N_11092,N_11340);
nor U11591 (N_11591,N_11204,N_11377);
xnor U11592 (N_11592,N_11400,N_11129);
xor U11593 (N_11593,N_11165,N_11325);
nor U11594 (N_11594,N_11494,N_11296);
or U11595 (N_11595,N_11497,N_11220);
nor U11596 (N_11596,N_11057,N_11492);
nand U11597 (N_11597,N_11062,N_11200);
nor U11598 (N_11598,N_11055,N_11170);
xor U11599 (N_11599,N_11444,N_11124);
and U11600 (N_11600,N_11428,N_11276);
nand U11601 (N_11601,N_11238,N_11117);
or U11602 (N_11602,N_11027,N_11401);
xor U11603 (N_11603,N_11006,N_11355);
xnor U11604 (N_11604,N_11368,N_11159);
nor U11605 (N_11605,N_11019,N_11386);
nand U11606 (N_11606,N_11100,N_11091);
nor U11607 (N_11607,N_11293,N_11270);
or U11608 (N_11608,N_11358,N_11306);
nor U11609 (N_11609,N_11373,N_11448);
nor U11610 (N_11610,N_11333,N_11162);
xor U11611 (N_11611,N_11004,N_11021);
xor U11612 (N_11612,N_11186,N_11281);
xnor U11613 (N_11613,N_11260,N_11257);
xnor U11614 (N_11614,N_11111,N_11464);
or U11615 (N_11615,N_11140,N_11311);
nand U11616 (N_11616,N_11320,N_11422);
nor U11617 (N_11617,N_11232,N_11419);
or U11618 (N_11618,N_11363,N_11015);
xor U11619 (N_11619,N_11264,N_11237);
or U11620 (N_11620,N_11496,N_11443);
nor U11621 (N_11621,N_11454,N_11191);
and U11622 (N_11622,N_11000,N_11332);
nand U11623 (N_11623,N_11187,N_11066);
nand U11624 (N_11624,N_11084,N_11142);
nor U11625 (N_11625,N_11221,N_11134);
nand U11626 (N_11626,N_11269,N_11216);
nor U11627 (N_11627,N_11109,N_11089);
xor U11628 (N_11628,N_11394,N_11212);
nor U11629 (N_11629,N_11016,N_11152);
or U11630 (N_11630,N_11230,N_11155);
nand U11631 (N_11631,N_11416,N_11387);
nor U11632 (N_11632,N_11002,N_11069);
nand U11633 (N_11633,N_11188,N_11239);
nor U11634 (N_11634,N_11227,N_11047);
nand U11635 (N_11635,N_11335,N_11145);
or U11636 (N_11636,N_11133,N_11123);
and U11637 (N_11637,N_11224,N_11096);
nand U11638 (N_11638,N_11183,N_11388);
nand U11639 (N_11639,N_11194,N_11287);
and U11640 (N_11640,N_11406,N_11495);
nor U11641 (N_11641,N_11384,N_11417);
nor U11642 (N_11642,N_11071,N_11121);
or U11643 (N_11643,N_11382,N_11225);
and U11644 (N_11644,N_11206,N_11005);
nor U11645 (N_11645,N_11344,N_11399);
or U11646 (N_11646,N_11476,N_11104);
nor U11647 (N_11647,N_11090,N_11299);
nor U11648 (N_11648,N_11302,N_11130);
nor U11649 (N_11649,N_11101,N_11292);
or U11650 (N_11650,N_11036,N_11106);
nor U11651 (N_11651,N_11395,N_11181);
nor U11652 (N_11652,N_11151,N_11432);
nand U11653 (N_11653,N_11023,N_11215);
and U11654 (N_11654,N_11010,N_11240);
or U11655 (N_11655,N_11467,N_11094);
xor U11656 (N_11656,N_11086,N_11014);
or U11657 (N_11657,N_11262,N_11482);
xor U11658 (N_11658,N_11007,N_11314);
or U11659 (N_11659,N_11275,N_11116);
and U11660 (N_11660,N_11449,N_11312);
nor U11661 (N_11661,N_11411,N_11026);
xnor U11662 (N_11662,N_11020,N_11163);
and U11663 (N_11663,N_11029,N_11011);
and U11664 (N_11664,N_11360,N_11280);
nor U11665 (N_11665,N_11339,N_11455);
xnor U11666 (N_11666,N_11135,N_11418);
and U11667 (N_11667,N_11425,N_11271);
nand U11668 (N_11668,N_11435,N_11322);
xor U11669 (N_11669,N_11105,N_11081);
nor U11670 (N_11670,N_11310,N_11077);
and U11671 (N_11671,N_11427,N_11357);
and U11672 (N_11672,N_11365,N_11013);
nor U11673 (N_11673,N_11087,N_11393);
nor U11674 (N_11674,N_11348,N_11396);
xnor U11675 (N_11675,N_11063,N_11331);
or U11676 (N_11676,N_11160,N_11298);
xor U11677 (N_11677,N_11043,N_11255);
or U11678 (N_11678,N_11336,N_11246);
nor U11679 (N_11679,N_11128,N_11478);
xnor U11680 (N_11680,N_11452,N_11157);
nor U11681 (N_11681,N_11214,N_11389);
xnor U11682 (N_11682,N_11041,N_11434);
and U11683 (N_11683,N_11226,N_11199);
nand U11684 (N_11684,N_11430,N_11285);
nand U11685 (N_11685,N_11437,N_11018);
nor U11686 (N_11686,N_11252,N_11450);
xnor U11687 (N_11687,N_11315,N_11334);
xnor U11688 (N_11688,N_11412,N_11371);
xor U11689 (N_11689,N_11342,N_11471);
nor U11690 (N_11690,N_11184,N_11085);
or U11691 (N_11691,N_11131,N_11119);
xor U11692 (N_11692,N_11035,N_11156);
nand U11693 (N_11693,N_11003,N_11040);
and U11694 (N_11694,N_11234,N_11475);
and U11695 (N_11695,N_11477,N_11189);
nand U11696 (N_11696,N_11479,N_11115);
nor U11697 (N_11697,N_11433,N_11439);
nor U11698 (N_11698,N_11017,N_11351);
and U11699 (N_11699,N_11289,N_11385);
xor U11700 (N_11700,N_11458,N_11174);
and U11701 (N_11701,N_11209,N_11381);
nand U11702 (N_11702,N_11354,N_11060);
and U11703 (N_11703,N_11148,N_11093);
nand U11704 (N_11704,N_11169,N_11158);
or U11705 (N_11705,N_11033,N_11404);
or U11706 (N_11706,N_11288,N_11190);
xnor U11707 (N_11707,N_11082,N_11440);
nand U11708 (N_11708,N_11445,N_11343);
nand U11709 (N_11709,N_11318,N_11064);
and U11710 (N_11710,N_11065,N_11211);
and U11711 (N_11711,N_11405,N_11488);
xnor U11712 (N_11712,N_11166,N_11330);
and U11713 (N_11713,N_11067,N_11039);
nand U11714 (N_11714,N_11469,N_11185);
xnor U11715 (N_11715,N_11095,N_11075);
and U11716 (N_11716,N_11028,N_11079);
and U11717 (N_11717,N_11468,N_11364);
nand U11718 (N_11718,N_11025,N_11466);
or U11719 (N_11719,N_11076,N_11048);
or U11720 (N_11720,N_11144,N_11460);
or U11721 (N_11721,N_11207,N_11179);
nand U11722 (N_11722,N_11498,N_11167);
nand U11723 (N_11723,N_11465,N_11056);
xnor U11724 (N_11724,N_11282,N_11141);
xnor U11725 (N_11725,N_11080,N_11201);
nor U11726 (N_11726,N_11126,N_11261);
or U11727 (N_11727,N_11222,N_11083);
xnor U11728 (N_11728,N_11321,N_11438);
and U11729 (N_11729,N_11486,N_11272);
or U11730 (N_11730,N_11154,N_11099);
nand U11731 (N_11731,N_11042,N_11286);
nor U11732 (N_11732,N_11319,N_11197);
or U11733 (N_11733,N_11328,N_11266);
and U11734 (N_11734,N_11139,N_11256);
nor U11735 (N_11735,N_11229,N_11391);
and U11736 (N_11736,N_11278,N_11103);
xnor U11737 (N_11737,N_11245,N_11456);
nand U11738 (N_11738,N_11313,N_11137);
and U11739 (N_11739,N_11491,N_11350);
nand U11740 (N_11740,N_11249,N_11372);
nor U11741 (N_11741,N_11171,N_11383);
or U11742 (N_11742,N_11022,N_11379);
xnor U11743 (N_11743,N_11242,N_11208);
nor U11744 (N_11744,N_11193,N_11058);
or U11745 (N_11745,N_11415,N_11484);
nand U11746 (N_11746,N_11305,N_11398);
nor U11747 (N_11747,N_11489,N_11050);
and U11748 (N_11748,N_11051,N_11480);
nand U11749 (N_11749,N_11097,N_11457);
xnor U11750 (N_11750,N_11166,N_11371);
xor U11751 (N_11751,N_11029,N_11064);
nand U11752 (N_11752,N_11490,N_11064);
or U11753 (N_11753,N_11018,N_11424);
or U11754 (N_11754,N_11107,N_11326);
or U11755 (N_11755,N_11355,N_11077);
and U11756 (N_11756,N_11261,N_11449);
or U11757 (N_11757,N_11169,N_11467);
nand U11758 (N_11758,N_11470,N_11140);
xnor U11759 (N_11759,N_11229,N_11280);
nand U11760 (N_11760,N_11318,N_11018);
and U11761 (N_11761,N_11221,N_11422);
nor U11762 (N_11762,N_11403,N_11442);
nor U11763 (N_11763,N_11076,N_11459);
xor U11764 (N_11764,N_11074,N_11369);
nand U11765 (N_11765,N_11335,N_11469);
and U11766 (N_11766,N_11380,N_11272);
or U11767 (N_11767,N_11437,N_11397);
nand U11768 (N_11768,N_11035,N_11248);
and U11769 (N_11769,N_11015,N_11040);
nor U11770 (N_11770,N_11088,N_11176);
and U11771 (N_11771,N_11386,N_11285);
and U11772 (N_11772,N_11359,N_11227);
and U11773 (N_11773,N_11333,N_11457);
or U11774 (N_11774,N_11043,N_11475);
xor U11775 (N_11775,N_11272,N_11439);
nor U11776 (N_11776,N_11143,N_11384);
or U11777 (N_11777,N_11481,N_11290);
nor U11778 (N_11778,N_11127,N_11297);
nand U11779 (N_11779,N_11452,N_11138);
xor U11780 (N_11780,N_11000,N_11006);
nor U11781 (N_11781,N_11477,N_11335);
xor U11782 (N_11782,N_11257,N_11105);
and U11783 (N_11783,N_11240,N_11244);
xor U11784 (N_11784,N_11329,N_11370);
nand U11785 (N_11785,N_11361,N_11194);
or U11786 (N_11786,N_11078,N_11430);
nand U11787 (N_11787,N_11148,N_11463);
xnor U11788 (N_11788,N_11044,N_11325);
nand U11789 (N_11789,N_11270,N_11306);
xor U11790 (N_11790,N_11367,N_11288);
and U11791 (N_11791,N_11413,N_11049);
nand U11792 (N_11792,N_11481,N_11206);
or U11793 (N_11793,N_11465,N_11034);
and U11794 (N_11794,N_11182,N_11322);
xnor U11795 (N_11795,N_11335,N_11443);
nor U11796 (N_11796,N_11286,N_11311);
nand U11797 (N_11797,N_11290,N_11463);
and U11798 (N_11798,N_11307,N_11086);
xor U11799 (N_11799,N_11487,N_11396);
nand U11800 (N_11800,N_11327,N_11214);
or U11801 (N_11801,N_11443,N_11064);
nand U11802 (N_11802,N_11461,N_11453);
or U11803 (N_11803,N_11228,N_11326);
or U11804 (N_11804,N_11282,N_11053);
and U11805 (N_11805,N_11397,N_11427);
nor U11806 (N_11806,N_11393,N_11207);
and U11807 (N_11807,N_11499,N_11488);
nor U11808 (N_11808,N_11365,N_11179);
and U11809 (N_11809,N_11139,N_11035);
or U11810 (N_11810,N_11128,N_11480);
nand U11811 (N_11811,N_11410,N_11044);
nand U11812 (N_11812,N_11160,N_11442);
xnor U11813 (N_11813,N_11245,N_11474);
nor U11814 (N_11814,N_11129,N_11038);
or U11815 (N_11815,N_11444,N_11174);
xnor U11816 (N_11816,N_11238,N_11379);
nor U11817 (N_11817,N_11338,N_11121);
nand U11818 (N_11818,N_11422,N_11456);
or U11819 (N_11819,N_11007,N_11102);
or U11820 (N_11820,N_11476,N_11363);
xnor U11821 (N_11821,N_11376,N_11282);
and U11822 (N_11822,N_11131,N_11137);
xor U11823 (N_11823,N_11295,N_11240);
nor U11824 (N_11824,N_11020,N_11070);
and U11825 (N_11825,N_11398,N_11480);
nand U11826 (N_11826,N_11104,N_11364);
or U11827 (N_11827,N_11165,N_11244);
and U11828 (N_11828,N_11403,N_11389);
xnor U11829 (N_11829,N_11048,N_11292);
xor U11830 (N_11830,N_11139,N_11198);
nor U11831 (N_11831,N_11202,N_11489);
nor U11832 (N_11832,N_11432,N_11143);
and U11833 (N_11833,N_11118,N_11415);
nand U11834 (N_11834,N_11233,N_11002);
and U11835 (N_11835,N_11217,N_11332);
nor U11836 (N_11836,N_11450,N_11110);
nor U11837 (N_11837,N_11047,N_11347);
and U11838 (N_11838,N_11254,N_11231);
or U11839 (N_11839,N_11135,N_11335);
nand U11840 (N_11840,N_11024,N_11256);
nand U11841 (N_11841,N_11432,N_11435);
nand U11842 (N_11842,N_11021,N_11399);
and U11843 (N_11843,N_11116,N_11022);
or U11844 (N_11844,N_11037,N_11336);
and U11845 (N_11845,N_11410,N_11139);
nand U11846 (N_11846,N_11215,N_11476);
xor U11847 (N_11847,N_11223,N_11245);
nor U11848 (N_11848,N_11486,N_11264);
nor U11849 (N_11849,N_11174,N_11218);
nand U11850 (N_11850,N_11305,N_11480);
or U11851 (N_11851,N_11405,N_11298);
and U11852 (N_11852,N_11072,N_11334);
nand U11853 (N_11853,N_11346,N_11212);
and U11854 (N_11854,N_11350,N_11441);
nand U11855 (N_11855,N_11138,N_11148);
and U11856 (N_11856,N_11276,N_11430);
xnor U11857 (N_11857,N_11497,N_11196);
or U11858 (N_11858,N_11469,N_11117);
xnor U11859 (N_11859,N_11495,N_11398);
or U11860 (N_11860,N_11164,N_11396);
nor U11861 (N_11861,N_11023,N_11287);
xor U11862 (N_11862,N_11224,N_11431);
and U11863 (N_11863,N_11493,N_11131);
and U11864 (N_11864,N_11392,N_11401);
nand U11865 (N_11865,N_11431,N_11111);
or U11866 (N_11866,N_11095,N_11014);
xor U11867 (N_11867,N_11211,N_11042);
and U11868 (N_11868,N_11460,N_11336);
nand U11869 (N_11869,N_11193,N_11402);
and U11870 (N_11870,N_11050,N_11042);
and U11871 (N_11871,N_11440,N_11024);
nor U11872 (N_11872,N_11440,N_11436);
or U11873 (N_11873,N_11198,N_11024);
xor U11874 (N_11874,N_11404,N_11181);
and U11875 (N_11875,N_11152,N_11207);
and U11876 (N_11876,N_11178,N_11337);
nor U11877 (N_11877,N_11038,N_11051);
nand U11878 (N_11878,N_11167,N_11073);
nor U11879 (N_11879,N_11158,N_11460);
nor U11880 (N_11880,N_11436,N_11223);
or U11881 (N_11881,N_11321,N_11121);
nand U11882 (N_11882,N_11013,N_11425);
or U11883 (N_11883,N_11226,N_11009);
or U11884 (N_11884,N_11263,N_11125);
nand U11885 (N_11885,N_11157,N_11077);
and U11886 (N_11886,N_11133,N_11329);
or U11887 (N_11887,N_11194,N_11456);
or U11888 (N_11888,N_11483,N_11444);
nor U11889 (N_11889,N_11412,N_11114);
nand U11890 (N_11890,N_11264,N_11137);
and U11891 (N_11891,N_11312,N_11303);
or U11892 (N_11892,N_11086,N_11336);
nor U11893 (N_11893,N_11255,N_11204);
or U11894 (N_11894,N_11435,N_11014);
and U11895 (N_11895,N_11149,N_11107);
nand U11896 (N_11896,N_11102,N_11079);
xnor U11897 (N_11897,N_11010,N_11431);
or U11898 (N_11898,N_11265,N_11274);
nand U11899 (N_11899,N_11412,N_11399);
nor U11900 (N_11900,N_11302,N_11033);
or U11901 (N_11901,N_11171,N_11214);
nor U11902 (N_11902,N_11087,N_11305);
or U11903 (N_11903,N_11355,N_11123);
and U11904 (N_11904,N_11232,N_11438);
xor U11905 (N_11905,N_11273,N_11311);
xnor U11906 (N_11906,N_11129,N_11391);
or U11907 (N_11907,N_11397,N_11440);
and U11908 (N_11908,N_11103,N_11071);
and U11909 (N_11909,N_11297,N_11489);
nand U11910 (N_11910,N_11081,N_11310);
xnor U11911 (N_11911,N_11423,N_11250);
and U11912 (N_11912,N_11190,N_11107);
or U11913 (N_11913,N_11237,N_11388);
and U11914 (N_11914,N_11390,N_11052);
xnor U11915 (N_11915,N_11305,N_11377);
or U11916 (N_11916,N_11204,N_11463);
nor U11917 (N_11917,N_11013,N_11165);
and U11918 (N_11918,N_11007,N_11201);
or U11919 (N_11919,N_11037,N_11174);
nor U11920 (N_11920,N_11283,N_11234);
xor U11921 (N_11921,N_11366,N_11370);
xor U11922 (N_11922,N_11456,N_11413);
or U11923 (N_11923,N_11218,N_11248);
xnor U11924 (N_11924,N_11181,N_11477);
or U11925 (N_11925,N_11376,N_11284);
nand U11926 (N_11926,N_11041,N_11348);
nor U11927 (N_11927,N_11049,N_11420);
xnor U11928 (N_11928,N_11232,N_11305);
or U11929 (N_11929,N_11135,N_11155);
nor U11930 (N_11930,N_11414,N_11144);
xnor U11931 (N_11931,N_11472,N_11120);
nand U11932 (N_11932,N_11096,N_11034);
nand U11933 (N_11933,N_11232,N_11076);
xnor U11934 (N_11934,N_11155,N_11092);
and U11935 (N_11935,N_11169,N_11460);
and U11936 (N_11936,N_11063,N_11153);
nand U11937 (N_11937,N_11391,N_11235);
nand U11938 (N_11938,N_11294,N_11258);
and U11939 (N_11939,N_11378,N_11156);
and U11940 (N_11940,N_11185,N_11104);
or U11941 (N_11941,N_11259,N_11043);
nor U11942 (N_11942,N_11012,N_11192);
or U11943 (N_11943,N_11063,N_11299);
or U11944 (N_11944,N_11440,N_11001);
xnor U11945 (N_11945,N_11280,N_11422);
nand U11946 (N_11946,N_11293,N_11215);
nand U11947 (N_11947,N_11137,N_11101);
nor U11948 (N_11948,N_11433,N_11427);
nor U11949 (N_11949,N_11267,N_11023);
xnor U11950 (N_11950,N_11400,N_11053);
xnor U11951 (N_11951,N_11142,N_11499);
and U11952 (N_11952,N_11495,N_11016);
xor U11953 (N_11953,N_11299,N_11250);
or U11954 (N_11954,N_11136,N_11286);
xor U11955 (N_11955,N_11158,N_11206);
or U11956 (N_11956,N_11202,N_11090);
and U11957 (N_11957,N_11478,N_11030);
or U11958 (N_11958,N_11069,N_11453);
and U11959 (N_11959,N_11166,N_11226);
xnor U11960 (N_11960,N_11005,N_11166);
and U11961 (N_11961,N_11059,N_11283);
nor U11962 (N_11962,N_11131,N_11048);
or U11963 (N_11963,N_11099,N_11190);
xnor U11964 (N_11964,N_11245,N_11287);
nor U11965 (N_11965,N_11367,N_11018);
xnor U11966 (N_11966,N_11199,N_11238);
xnor U11967 (N_11967,N_11233,N_11396);
and U11968 (N_11968,N_11109,N_11420);
and U11969 (N_11969,N_11232,N_11110);
xor U11970 (N_11970,N_11341,N_11423);
nand U11971 (N_11971,N_11241,N_11117);
xnor U11972 (N_11972,N_11066,N_11380);
xnor U11973 (N_11973,N_11267,N_11182);
nand U11974 (N_11974,N_11392,N_11201);
nor U11975 (N_11975,N_11057,N_11270);
and U11976 (N_11976,N_11007,N_11172);
nor U11977 (N_11977,N_11265,N_11458);
xor U11978 (N_11978,N_11388,N_11363);
xor U11979 (N_11979,N_11030,N_11394);
nand U11980 (N_11980,N_11003,N_11282);
or U11981 (N_11981,N_11104,N_11139);
or U11982 (N_11982,N_11365,N_11325);
nor U11983 (N_11983,N_11259,N_11483);
nand U11984 (N_11984,N_11141,N_11313);
and U11985 (N_11985,N_11088,N_11183);
xnor U11986 (N_11986,N_11091,N_11369);
and U11987 (N_11987,N_11045,N_11360);
xor U11988 (N_11988,N_11235,N_11093);
nand U11989 (N_11989,N_11215,N_11258);
and U11990 (N_11990,N_11214,N_11492);
nand U11991 (N_11991,N_11066,N_11346);
nand U11992 (N_11992,N_11039,N_11138);
and U11993 (N_11993,N_11051,N_11194);
nand U11994 (N_11994,N_11229,N_11352);
nand U11995 (N_11995,N_11434,N_11068);
or U11996 (N_11996,N_11185,N_11236);
and U11997 (N_11997,N_11255,N_11453);
or U11998 (N_11998,N_11141,N_11409);
nand U11999 (N_11999,N_11123,N_11397);
nor U12000 (N_12000,N_11988,N_11847);
nor U12001 (N_12001,N_11773,N_11739);
or U12002 (N_12002,N_11743,N_11570);
nor U12003 (N_12003,N_11961,N_11909);
and U12004 (N_12004,N_11529,N_11654);
or U12005 (N_12005,N_11955,N_11874);
nor U12006 (N_12006,N_11919,N_11602);
xor U12007 (N_12007,N_11515,N_11780);
and U12008 (N_12008,N_11678,N_11823);
nor U12009 (N_12009,N_11781,N_11645);
nor U12010 (N_12010,N_11849,N_11718);
or U12011 (N_12011,N_11982,N_11558);
and U12012 (N_12012,N_11600,N_11628);
and U12013 (N_12013,N_11956,N_11524);
nor U12014 (N_12014,N_11998,N_11798);
and U12015 (N_12015,N_11688,N_11794);
nor U12016 (N_12016,N_11980,N_11997);
or U12017 (N_12017,N_11624,N_11971);
nand U12018 (N_12018,N_11670,N_11875);
xor U12019 (N_12019,N_11603,N_11972);
xor U12020 (N_12020,N_11950,N_11711);
or U12021 (N_12021,N_11845,N_11785);
or U12022 (N_12022,N_11712,N_11755);
or U12023 (N_12023,N_11817,N_11698);
nand U12024 (N_12024,N_11680,N_11585);
xor U12025 (N_12025,N_11837,N_11729);
and U12026 (N_12026,N_11935,N_11533);
xor U12027 (N_12027,N_11793,N_11520);
and U12028 (N_12028,N_11860,N_11967);
nor U12029 (N_12029,N_11801,N_11888);
nand U12030 (N_12030,N_11735,N_11588);
or U12031 (N_12031,N_11548,N_11502);
xnor U12032 (N_12032,N_11852,N_11775);
or U12033 (N_12033,N_11836,N_11746);
and U12034 (N_12034,N_11942,N_11815);
nand U12035 (N_12035,N_11606,N_11699);
xor U12036 (N_12036,N_11983,N_11995);
or U12037 (N_12037,N_11800,N_11807);
and U12038 (N_12038,N_11648,N_11541);
xor U12039 (N_12039,N_11557,N_11978);
or U12040 (N_12040,N_11578,N_11723);
or U12041 (N_12041,N_11841,N_11689);
nor U12042 (N_12042,N_11776,N_11632);
nor U12043 (N_12043,N_11973,N_11898);
or U12044 (N_12044,N_11531,N_11677);
xor U12045 (N_12045,N_11864,N_11911);
nor U12046 (N_12046,N_11709,N_11617);
nand U12047 (N_12047,N_11681,N_11822);
xnor U12048 (N_12048,N_11749,N_11625);
nand U12049 (N_12049,N_11762,N_11834);
and U12050 (N_12050,N_11721,N_11519);
or U12051 (N_12051,N_11902,N_11503);
nand U12052 (N_12052,N_11716,N_11663);
nand U12053 (N_12053,N_11782,N_11991);
and U12054 (N_12054,N_11806,N_11564);
and U12055 (N_12055,N_11959,N_11952);
nand U12056 (N_12056,N_11906,N_11535);
and U12057 (N_12057,N_11510,N_11863);
nand U12058 (N_12058,N_11941,N_11897);
and U12059 (N_12059,N_11777,N_11984);
or U12060 (N_12060,N_11544,N_11958);
xnor U12061 (N_12061,N_11752,N_11674);
or U12062 (N_12062,N_11797,N_11910);
xnor U12063 (N_12063,N_11804,N_11900);
nor U12064 (N_12064,N_11808,N_11646);
xor U12065 (N_12065,N_11504,N_11827);
or U12066 (N_12066,N_11922,N_11741);
and U12067 (N_12067,N_11597,N_11856);
nor U12068 (N_12068,N_11715,N_11946);
or U12069 (N_12069,N_11891,N_11756);
and U12070 (N_12070,N_11599,N_11929);
nand U12071 (N_12071,N_11682,N_11728);
and U12072 (N_12072,N_11870,N_11561);
and U12073 (N_12073,N_11620,N_11990);
nor U12074 (N_12074,N_11788,N_11799);
nor U12075 (N_12075,N_11894,N_11885);
xnor U12076 (N_12076,N_11904,N_11934);
xor U12077 (N_12077,N_11812,N_11517);
nor U12078 (N_12078,N_11905,N_11683);
nor U12079 (N_12079,N_11744,N_11613);
nor U12080 (N_12080,N_11994,N_11887);
nand U12081 (N_12081,N_11965,N_11501);
and U12082 (N_12082,N_11884,N_11825);
nor U12083 (N_12083,N_11824,N_11719);
nor U12084 (N_12084,N_11697,N_11577);
xor U12085 (N_12085,N_11987,N_11700);
xnor U12086 (N_12086,N_11704,N_11920);
nor U12087 (N_12087,N_11575,N_11754);
and U12088 (N_12088,N_11572,N_11805);
or U12089 (N_12089,N_11895,N_11758);
nand U12090 (N_12090,N_11552,N_11516);
nand U12091 (N_12091,N_11886,N_11616);
nor U12092 (N_12092,N_11927,N_11556);
or U12093 (N_12093,N_11720,N_11615);
xor U12094 (N_12094,N_11926,N_11634);
and U12095 (N_12095,N_11896,N_11742);
nor U12096 (N_12096,N_11644,N_11623);
and U12097 (N_12097,N_11566,N_11550);
and U12098 (N_12098,N_11530,N_11523);
or U12099 (N_12099,N_11907,N_11859);
nand U12100 (N_12100,N_11977,N_11810);
and U12101 (N_12101,N_11707,N_11921);
and U12102 (N_12102,N_11702,N_11507);
or U12103 (N_12103,N_11727,N_11667);
or U12104 (N_12104,N_11976,N_11944);
xor U12105 (N_12105,N_11713,N_11893);
or U12106 (N_12106,N_11771,N_11732);
nor U12107 (N_12107,N_11768,N_11914);
xnor U12108 (N_12108,N_11916,N_11511);
or U12109 (N_12109,N_11586,N_11760);
and U12110 (N_12110,N_11803,N_11652);
xor U12111 (N_12111,N_11855,N_11751);
xor U12112 (N_12112,N_11953,N_11555);
and U12113 (N_12113,N_11937,N_11779);
or U12114 (N_12114,N_11705,N_11611);
nand U12115 (N_12115,N_11876,N_11996);
nand U12116 (N_12116,N_11506,N_11649);
nand U12117 (N_12117,N_11607,N_11598);
xor U12118 (N_12118,N_11641,N_11505);
nand U12119 (N_12119,N_11701,N_11753);
and U12120 (N_12120,N_11818,N_11672);
nor U12121 (N_12121,N_11786,N_11629);
xnor U12122 (N_12122,N_11925,N_11609);
and U12123 (N_12123,N_11717,N_11656);
nand U12124 (N_12124,N_11665,N_11745);
and U12125 (N_12125,N_11630,N_11936);
nor U12126 (N_12126,N_11542,N_11589);
nor U12127 (N_12127,N_11733,N_11576);
nand U12128 (N_12128,N_11584,N_11545);
nor U12129 (N_12129,N_11591,N_11869);
and U12130 (N_12130,N_11872,N_11608);
or U12131 (N_12131,N_11787,N_11693);
and U12132 (N_12132,N_11651,N_11692);
or U12133 (N_12133,N_11748,N_11833);
nand U12134 (N_12134,N_11842,N_11547);
xnor U12135 (N_12135,N_11851,N_11695);
nand U12136 (N_12136,N_11974,N_11830);
nand U12137 (N_12137,N_11708,N_11571);
xnor U12138 (N_12138,N_11500,N_11846);
and U12139 (N_12139,N_11525,N_11881);
or U12140 (N_12140,N_11553,N_11923);
nand U12141 (N_12141,N_11819,N_11738);
nand U12142 (N_12142,N_11573,N_11590);
and U12143 (N_12143,N_11828,N_11594);
nand U12144 (N_12144,N_11759,N_11774);
nand U12145 (N_12145,N_11631,N_11789);
nand U12146 (N_12146,N_11538,N_11690);
nor U12147 (N_12147,N_11962,N_11612);
nand U12148 (N_12148,N_11899,N_11873);
or U12149 (N_12149,N_11867,N_11696);
xnor U12150 (N_12150,N_11521,N_11622);
or U12151 (N_12151,N_11795,N_11981);
and U12152 (N_12152,N_11853,N_11924);
xnor U12153 (N_12153,N_11635,N_11737);
and U12154 (N_12154,N_11569,N_11838);
and U12155 (N_12155,N_11731,N_11858);
xnor U12156 (N_12156,N_11559,N_11862);
or U12157 (N_12157,N_11673,N_11587);
or U12158 (N_12158,N_11889,N_11540);
or U12159 (N_12159,N_11593,N_11664);
nand U12160 (N_12160,N_11660,N_11595);
nand U12161 (N_12161,N_11592,N_11618);
and U12162 (N_12162,N_11657,N_11669);
xor U12163 (N_12163,N_11835,N_11975);
nor U12164 (N_12164,N_11912,N_11596);
nand U12165 (N_12165,N_11957,N_11843);
and U12166 (N_12166,N_11605,N_11802);
xnor U12167 (N_12167,N_11883,N_11676);
or U12168 (N_12168,N_11943,N_11796);
and U12169 (N_12169,N_11903,N_11966);
xnor U12170 (N_12170,N_11765,N_11901);
nand U12171 (N_12171,N_11850,N_11546);
or U12172 (N_12172,N_11933,N_11642);
xnor U12173 (N_12173,N_11757,N_11964);
xnor U12174 (N_12174,N_11979,N_11528);
xor U12175 (N_12175,N_11627,N_11908);
or U12176 (N_12176,N_11948,N_11890);
or U12177 (N_12177,N_11614,N_11650);
nand U12178 (N_12178,N_11960,N_11684);
nand U12179 (N_12179,N_11522,N_11999);
nor U12180 (N_12180,N_11767,N_11949);
nand U12181 (N_12181,N_11565,N_11579);
nor U12182 (N_12182,N_11954,N_11826);
nor U12183 (N_12183,N_11604,N_11724);
nor U12184 (N_12184,N_11537,N_11963);
xor U12185 (N_12185,N_11857,N_11951);
nand U12186 (N_12186,N_11580,N_11915);
nand U12187 (N_12187,N_11726,N_11918);
nor U12188 (N_12188,N_11568,N_11633);
xnor U12189 (N_12189,N_11985,N_11534);
nand U12190 (N_12190,N_11626,N_11583);
xor U12191 (N_12191,N_11513,N_11947);
nand U12192 (N_12192,N_11551,N_11878);
or U12193 (N_12193,N_11784,N_11560);
nand U12194 (N_12194,N_11725,N_11582);
or U12195 (N_12195,N_11816,N_11791);
nor U12196 (N_12196,N_11621,N_11706);
or U12197 (N_12197,N_11829,N_11740);
or U12198 (N_12198,N_11871,N_11854);
or U12199 (N_12199,N_11832,N_11730);
and U12200 (N_12200,N_11714,N_11750);
or U12201 (N_12201,N_11666,N_11970);
and U12202 (N_12202,N_11993,N_11992);
nand U12203 (N_12203,N_11882,N_11679);
xor U12204 (N_12204,N_11518,N_11928);
xnor U12205 (N_12205,N_11769,N_11989);
xnor U12206 (N_12206,N_11831,N_11747);
and U12207 (N_12207,N_11763,N_11968);
nor U12208 (N_12208,N_11514,N_11655);
xnor U12209 (N_12209,N_11809,N_11839);
nor U12210 (N_12210,N_11581,N_11844);
nand U12211 (N_12211,N_11880,N_11790);
or U12212 (N_12212,N_11686,N_11938);
or U12213 (N_12213,N_11821,N_11526);
nor U12214 (N_12214,N_11930,N_11764);
nor U12215 (N_12215,N_11868,N_11512);
nand U12216 (N_12216,N_11866,N_11865);
or U12217 (N_12217,N_11574,N_11668);
nor U12218 (N_12218,N_11601,N_11662);
and U12219 (N_12219,N_11772,N_11792);
nor U12220 (N_12220,N_11913,N_11685);
nor U12221 (N_12221,N_11527,N_11734);
nor U12222 (N_12222,N_11820,N_11761);
xnor U12223 (N_12223,N_11539,N_11932);
nor U12224 (N_12224,N_11637,N_11653);
nand U12225 (N_12225,N_11687,N_11879);
or U12226 (N_12226,N_11770,N_11940);
nand U12227 (N_12227,N_11783,N_11619);
or U12228 (N_12228,N_11532,N_11563);
nor U12229 (N_12229,N_11636,N_11694);
or U12230 (N_12230,N_11917,N_11861);
xnor U12231 (N_12231,N_11877,N_11508);
and U12232 (N_12232,N_11945,N_11610);
nand U12233 (N_12233,N_11736,N_11778);
or U12234 (N_12234,N_11536,N_11643);
nand U12235 (N_12235,N_11661,N_11811);
and U12236 (N_12236,N_11691,N_11722);
nor U12237 (N_12237,N_11840,N_11813);
or U12238 (N_12238,N_11671,N_11658);
and U12239 (N_12239,N_11640,N_11814);
xor U12240 (N_12240,N_11647,N_11710);
xnor U12241 (N_12241,N_11986,N_11969);
or U12242 (N_12242,N_11567,N_11543);
nand U12243 (N_12243,N_11939,N_11892);
xnor U12244 (N_12244,N_11766,N_11509);
nand U12245 (N_12245,N_11639,N_11931);
nor U12246 (N_12246,N_11549,N_11554);
xnor U12247 (N_12247,N_11675,N_11659);
and U12248 (N_12248,N_11703,N_11848);
xnor U12249 (N_12249,N_11562,N_11638);
and U12250 (N_12250,N_11593,N_11571);
nand U12251 (N_12251,N_11540,N_11526);
and U12252 (N_12252,N_11945,N_11847);
and U12253 (N_12253,N_11571,N_11917);
xnor U12254 (N_12254,N_11761,N_11828);
and U12255 (N_12255,N_11521,N_11660);
and U12256 (N_12256,N_11784,N_11968);
and U12257 (N_12257,N_11646,N_11595);
nor U12258 (N_12258,N_11515,N_11718);
nor U12259 (N_12259,N_11632,N_11921);
or U12260 (N_12260,N_11876,N_11668);
xnor U12261 (N_12261,N_11567,N_11772);
nand U12262 (N_12262,N_11597,N_11864);
xnor U12263 (N_12263,N_11891,N_11994);
and U12264 (N_12264,N_11575,N_11560);
and U12265 (N_12265,N_11644,N_11656);
nor U12266 (N_12266,N_11843,N_11833);
or U12267 (N_12267,N_11946,N_11759);
or U12268 (N_12268,N_11922,N_11543);
xor U12269 (N_12269,N_11566,N_11548);
and U12270 (N_12270,N_11782,N_11791);
or U12271 (N_12271,N_11515,N_11503);
nand U12272 (N_12272,N_11993,N_11719);
nand U12273 (N_12273,N_11724,N_11646);
and U12274 (N_12274,N_11536,N_11746);
nand U12275 (N_12275,N_11639,N_11673);
xnor U12276 (N_12276,N_11702,N_11550);
nor U12277 (N_12277,N_11543,N_11628);
or U12278 (N_12278,N_11876,N_11643);
or U12279 (N_12279,N_11676,N_11550);
nand U12280 (N_12280,N_11537,N_11940);
and U12281 (N_12281,N_11670,N_11584);
nand U12282 (N_12282,N_11518,N_11685);
xor U12283 (N_12283,N_11943,N_11509);
nand U12284 (N_12284,N_11860,N_11583);
xor U12285 (N_12285,N_11705,N_11648);
nor U12286 (N_12286,N_11890,N_11512);
nor U12287 (N_12287,N_11943,N_11827);
or U12288 (N_12288,N_11874,N_11836);
or U12289 (N_12289,N_11996,N_11922);
nand U12290 (N_12290,N_11594,N_11575);
and U12291 (N_12291,N_11694,N_11695);
and U12292 (N_12292,N_11758,N_11996);
or U12293 (N_12293,N_11575,N_11807);
nand U12294 (N_12294,N_11877,N_11800);
nor U12295 (N_12295,N_11730,N_11654);
nor U12296 (N_12296,N_11941,N_11639);
or U12297 (N_12297,N_11707,N_11764);
and U12298 (N_12298,N_11868,N_11976);
nand U12299 (N_12299,N_11947,N_11730);
and U12300 (N_12300,N_11891,N_11775);
nor U12301 (N_12301,N_11816,N_11945);
and U12302 (N_12302,N_11551,N_11740);
xnor U12303 (N_12303,N_11937,N_11741);
xnor U12304 (N_12304,N_11909,N_11932);
nand U12305 (N_12305,N_11550,N_11932);
xor U12306 (N_12306,N_11874,N_11919);
xor U12307 (N_12307,N_11704,N_11598);
xnor U12308 (N_12308,N_11786,N_11780);
nand U12309 (N_12309,N_11786,N_11728);
and U12310 (N_12310,N_11552,N_11671);
xnor U12311 (N_12311,N_11903,N_11620);
and U12312 (N_12312,N_11963,N_11806);
xnor U12313 (N_12313,N_11961,N_11566);
and U12314 (N_12314,N_11523,N_11611);
xor U12315 (N_12315,N_11554,N_11715);
nor U12316 (N_12316,N_11853,N_11640);
or U12317 (N_12317,N_11935,N_11668);
and U12318 (N_12318,N_11691,N_11596);
nand U12319 (N_12319,N_11781,N_11507);
nand U12320 (N_12320,N_11511,N_11690);
and U12321 (N_12321,N_11995,N_11905);
nand U12322 (N_12322,N_11687,N_11781);
and U12323 (N_12323,N_11710,N_11840);
xnor U12324 (N_12324,N_11870,N_11690);
or U12325 (N_12325,N_11756,N_11652);
nor U12326 (N_12326,N_11911,N_11705);
xnor U12327 (N_12327,N_11814,N_11660);
and U12328 (N_12328,N_11865,N_11841);
nor U12329 (N_12329,N_11585,N_11743);
nand U12330 (N_12330,N_11810,N_11995);
nand U12331 (N_12331,N_11561,N_11695);
xnor U12332 (N_12332,N_11551,N_11757);
or U12333 (N_12333,N_11655,N_11622);
nand U12334 (N_12334,N_11745,N_11793);
nor U12335 (N_12335,N_11768,N_11542);
nor U12336 (N_12336,N_11510,N_11958);
nor U12337 (N_12337,N_11691,N_11666);
nor U12338 (N_12338,N_11916,N_11594);
xnor U12339 (N_12339,N_11672,N_11529);
xor U12340 (N_12340,N_11891,N_11512);
or U12341 (N_12341,N_11701,N_11704);
nand U12342 (N_12342,N_11726,N_11968);
and U12343 (N_12343,N_11914,N_11588);
xnor U12344 (N_12344,N_11795,N_11794);
xor U12345 (N_12345,N_11834,N_11840);
and U12346 (N_12346,N_11941,N_11577);
and U12347 (N_12347,N_11510,N_11783);
nand U12348 (N_12348,N_11918,N_11718);
nor U12349 (N_12349,N_11709,N_11751);
and U12350 (N_12350,N_11948,N_11968);
or U12351 (N_12351,N_11612,N_11516);
nor U12352 (N_12352,N_11843,N_11887);
nand U12353 (N_12353,N_11634,N_11749);
nor U12354 (N_12354,N_11530,N_11895);
nand U12355 (N_12355,N_11548,N_11618);
or U12356 (N_12356,N_11550,N_11565);
nand U12357 (N_12357,N_11833,N_11708);
nand U12358 (N_12358,N_11844,N_11867);
nor U12359 (N_12359,N_11947,N_11965);
and U12360 (N_12360,N_11572,N_11561);
xnor U12361 (N_12361,N_11827,N_11749);
xor U12362 (N_12362,N_11973,N_11904);
or U12363 (N_12363,N_11583,N_11853);
nor U12364 (N_12364,N_11652,N_11865);
nor U12365 (N_12365,N_11842,N_11863);
nor U12366 (N_12366,N_11905,N_11562);
and U12367 (N_12367,N_11508,N_11892);
nor U12368 (N_12368,N_11612,N_11995);
and U12369 (N_12369,N_11640,N_11977);
and U12370 (N_12370,N_11946,N_11890);
xor U12371 (N_12371,N_11827,N_11679);
and U12372 (N_12372,N_11710,N_11963);
or U12373 (N_12373,N_11809,N_11782);
or U12374 (N_12374,N_11925,N_11750);
nand U12375 (N_12375,N_11870,N_11862);
nor U12376 (N_12376,N_11737,N_11636);
nor U12377 (N_12377,N_11943,N_11803);
or U12378 (N_12378,N_11508,N_11857);
nand U12379 (N_12379,N_11666,N_11594);
nand U12380 (N_12380,N_11864,N_11764);
nor U12381 (N_12381,N_11929,N_11570);
nand U12382 (N_12382,N_11680,N_11582);
or U12383 (N_12383,N_11660,N_11534);
nor U12384 (N_12384,N_11503,N_11542);
and U12385 (N_12385,N_11507,N_11704);
xnor U12386 (N_12386,N_11611,N_11707);
nor U12387 (N_12387,N_11656,N_11688);
xnor U12388 (N_12388,N_11887,N_11981);
and U12389 (N_12389,N_11517,N_11959);
and U12390 (N_12390,N_11996,N_11957);
or U12391 (N_12391,N_11679,N_11618);
or U12392 (N_12392,N_11708,N_11840);
or U12393 (N_12393,N_11952,N_11591);
or U12394 (N_12394,N_11924,N_11964);
nand U12395 (N_12395,N_11954,N_11968);
nand U12396 (N_12396,N_11579,N_11832);
or U12397 (N_12397,N_11784,N_11617);
nor U12398 (N_12398,N_11797,N_11716);
and U12399 (N_12399,N_11574,N_11536);
xor U12400 (N_12400,N_11744,N_11838);
xnor U12401 (N_12401,N_11801,N_11889);
nor U12402 (N_12402,N_11693,N_11753);
nor U12403 (N_12403,N_11715,N_11568);
nand U12404 (N_12404,N_11624,N_11748);
xor U12405 (N_12405,N_11842,N_11520);
and U12406 (N_12406,N_11778,N_11883);
xnor U12407 (N_12407,N_11550,N_11694);
or U12408 (N_12408,N_11901,N_11611);
nor U12409 (N_12409,N_11593,N_11659);
and U12410 (N_12410,N_11691,N_11778);
and U12411 (N_12411,N_11888,N_11626);
and U12412 (N_12412,N_11783,N_11694);
xor U12413 (N_12413,N_11658,N_11833);
xor U12414 (N_12414,N_11802,N_11660);
or U12415 (N_12415,N_11910,N_11841);
and U12416 (N_12416,N_11929,N_11624);
or U12417 (N_12417,N_11692,N_11919);
or U12418 (N_12418,N_11988,N_11944);
nor U12419 (N_12419,N_11946,N_11665);
nand U12420 (N_12420,N_11691,N_11587);
nand U12421 (N_12421,N_11722,N_11527);
and U12422 (N_12422,N_11818,N_11970);
or U12423 (N_12423,N_11520,N_11855);
nand U12424 (N_12424,N_11761,N_11524);
or U12425 (N_12425,N_11550,N_11531);
and U12426 (N_12426,N_11747,N_11784);
and U12427 (N_12427,N_11628,N_11705);
nor U12428 (N_12428,N_11758,N_11765);
nor U12429 (N_12429,N_11925,N_11747);
nand U12430 (N_12430,N_11858,N_11802);
or U12431 (N_12431,N_11626,N_11947);
xor U12432 (N_12432,N_11945,N_11543);
nor U12433 (N_12433,N_11897,N_11547);
nand U12434 (N_12434,N_11599,N_11585);
nor U12435 (N_12435,N_11924,N_11830);
or U12436 (N_12436,N_11803,N_11749);
nor U12437 (N_12437,N_11715,N_11518);
and U12438 (N_12438,N_11529,N_11710);
xnor U12439 (N_12439,N_11729,N_11957);
xnor U12440 (N_12440,N_11984,N_11989);
nor U12441 (N_12441,N_11949,N_11775);
or U12442 (N_12442,N_11512,N_11810);
nor U12443 (N_12443,N_11595,N_11928);
and U12444 (N_12444,N_11685,N_11553);
xor U12445 (N_12445,N_11508,N_11505);
nand U12446 (N_12446,N_11604,N_11960);
or U12447 (N_12447,N_11724,N_11888);
nor U12448 (N_12448,N_11502,N_11535);
nand U12449 (N_12449,N_11844,N_11547);
or U12450 (N_12450,N_11949,N_11560);
and U12451 (N_12451,N_11734,N_11926);
nor U12452 (N_12452,N_11814,N_11925);
xor U12453 (N_12453,N_11809,N_11868);
and U12454 (N_12454,N_11929,N_11596);
nand U12455 (N_12455,N_11563,N_11720);
or U12456 (N_12456,N_11543,N_11767);
nand U12457 (N_12457,N_11776,N_11719);
xnor U12458 (N_12458,N_11970,N_11882);
and U12459 (N_12459,N_11735,N_11666);
xnor U12460 (N_12460,N_11900,N_11743);
or U12461 (N_12461,N_11911,N_11599);
xnor U12462 (N_12462,N_11806,N_11591);
and U12463 (N_12463,N_11745,N_11734);
nand U12464 (N_12464,N_11682,N_11991);
and U12465 (N_12465,N_11681,N_11554);
and U12466 (N_12466,N_11778,N_11677);
xor U12467 (N_12467,N_11658,N_11801);
nor U12468 (N_12468,N_11810,N_11877);
or U12469 (N_12469,N_11533,N_11799);
xor U12470 (N_12470,N_11890,N_11867);
xor U12471 (N_12471,N_11514,N_11658);
nand U12472 (N_12472,N_11997,N_11676);
or U12473 (N_12473,N_11512,N_11729);
nor U12474 (N_12474,N_11975,N_11831);
nor U12475 (N_12475,N_11591,N_11989);
xnor U12476 (N_12476,N_11943,N_11564);
or U12477 (N_12477,N_11691,N_11972);
nand U12478 (N_12478,N_11708,N_11815);
nor U12479 (N_12479,N_11928,N_11657);
nand U12480 (N_12480,N_11769,N_11720);
and U12481 (N_12481,N_11603,N_11535);
xor U12482 (N_12482,N_11853,N_11801);
xnor U12483 (N_12483,N_11524,N_11726);
nor U12484 (N_12484,N_11724,N_11721);
or U12485 (N_12485,N_11917,N_11559);
or U12486 (N_12486,N_11608,N_11946);
nand U12487 (N_12487,N_11546,N_11674);
nor U12488 (N_12488,N_11723,N_11636);
or U12489 (N_12489,N_11913,N_11544);
nand U12490 (N_12490,N_11562,N_11762);
and U12491 (N_12491,N_11628,N_11760);
and U12492 (N_12492,N_11832,N_11819);
nand U12493 (N_12493,N_11824,N_11975);
nor U12494 (N_12494,N_11601,N_11881);
and U12495 (N_12495,N_11741,N_11784);
or U12496 (N_12496,N_11810,N_11768);
nor U12497 (N_12497,N_11681,N_11585);
xnor U12498 (N_12498,N_11592,N_11977);
and U12499 (N_12499,N_11526,N_11645);
or U12500 (N_12500,N_12368,N_12005);
nor U12501 (N_12501,N_12215,N_12362);
nor U12502 (N_12502,N_12477,N_12141);
or U12503 (N_12503,N_12355,N_12148);
nor U12504 (N_12504,N_12070,N_12492);
nor U12505 (N_12505,N_12069,N_12346);
nor U12506 (N_12506,N_12391,N_12003);
and U12507 (N_12507,N_12016,N_12091);
or U12508 (N_12508,N_12295,N_12390);
or U12509 (N_12509,N_12487,N_12190);
nor U12510 (N_12510,N_12094,N_12344);
or U12511 (N_12511,N_12235,N_12058);
nand U12512 (N_12512,N_12345,N_12481);
nand U12513 (N_12513,N_12373,N_12065);
or U12514 (N_12514,N_12145,N_12030);
xnor U12515 (N_12515,N_12157,N_12056);
and U12516 (N_12516,N_12227,N_12146);
xnor U12517 (N_12517,N_12417,N_12310);
xnor U12518 (N_12518,N_12000,N_12316);
nor U12519 (N_12519,N_12176,N_12133);
nor U12520 (N_12520,N_12137,N_12024);
nand U12521 (N_12521,N_12040,N_12049);
and U12522 (N_12522,N_12407,N_12131);
nand U12523 (N_12523,N_12472,N_12102);
nand U12524 (N_12524,N_12122,N_12011);
and U12525 (N_12525,N_12413,N_12339);
and U12526 (N_12526,N_12020,N_12113);
nand U12527 (N_12527,N_12135,N_12100);
or U12528 (N_12528,N_12367,N_12464);
nor U12529 (N_12529,N_12357,N_12231);
xnor U12530 (N_12530,N_12175,N_12479);
nand U12531 (N_12531,N_12258,N_12107);
and U12532 (N_12532,N_12441,N_12035);
and U12533 (N_12533,N_12151,N_12170);
xnor U12534 (N_12534,N_12178,N_12382);
xnor U12535 (N_12535,N_12017,N_12395);
or U12536 (N_12536,N_12437,N_12315);
and U12537 (N_12537,N_12116,N_12248);
xnor U12538 (N_12538,N_12433,N_12436);
and U12539 (N_12539,N_12121,N_12105);
and U12540 (N_12540,N_12473,N_12338);
nor U12541 (N_12541,N_12155,N_12266);
xnor U12542 (N_12542,N_12241,N_12474);
xor U12543 (N_12543,N_12160,N_12370);
xor U12544 (N_12544,N_12119,N_12244);
nand U12545 (N_12545,N_12335,N_12279);
and U12546 (N_12546,N_12312,N_12114);
xnor U12547 (N_12547,N_12064,N_12221);
and U12548 (N_12548,N_12055,N_12467);
nor U12549 (N_12549,N_12053,N_12340);
or U12550 (N_12550,N_12080,N_12410);
nor U12551 (N_12551,N_12220,N_12015);
or U12552 (N_12552,N_12277,N_12354);
nor U12553 (N_12553,N_12229,N_12036);
and U12554 (N_12554,N_12478,N_12249);
xnor U12555 (N_12555,N_12179,N_12187);
nor U12556 (N_12556,N_12047,N_12198);
and U12557 (N_12557,N_12171,N_12404);
nor U12558 (N_12558,N_12378,N_12434);
nor U12559 (N_12559,N_12439,N_12324);
and U12560 (N_12560,N_12387,N_12485);
nand U12561 (N_12561,N_12325,N_12350);
or U12562 (N_12562,N_12161,N_12250);
nand U12563 (N_12563,N_12284,N_12242);
xor U12564 (N_12564,N_12012,N_12351);
and U12565 (N_12565,N_12348,N_12044);
and U12566 (N_12566,N_12411,N_12383);
nor U12567 (N_12567,N_12123,N_12446);
nand U12568 (N_12568,N_12431,N_12112);
xor U12569 (N_12569,N_12128,N_12422);
xnor U12570 (N_12570,N_12063,N_12163);
nor U12571 (N_12571,N_12453,N_12222);
nand U12572 (N_12572,N_12104,N_12469);
nor U12573 (N_12573,N_12247,N_12461);
or U12574 (N_12574,N_12330,N_12271);
or U12575 (N_12575,N_12255,N_12214);
nand U12576 (N_12576,N_12369,N_12318);
and U12577 (N_12577,N_12033,N_12239);
nand U12578 (N_12578,N_12207,N_12319);
nand U12579 (N_12579,N_12287,N_12209);
and U12580 (N_12580,N_12167,N_12072);
xor U12581 (N_12581,N_12275,N_12412);
nor U12582 (N_12582,N_12392,N_12211);
nor U12583 (N_12583,N_12313,N_12193);
and U12584 (N_12584,N_12272,N_12142);
or U12585 (N_12585,N_12010,N_12085);
xnor U12586 (N_12586,N_12483,N_12257);
nand U12587 (N_12587,N_12356,N_12071);
and U12588 (N_12588,N_12043,N_12019);
nor U12589 (N_12589,N_12031,N_12343);
or U12590 (N_12590,N_12371,N_12219);
and U12591 (N_12591,N_12217,N_12365);
and U12592 (N_12592,N_12195,N_12223);
or U12593 (N_12593,N_12398,N_12432);
nand U12594 (N_12594,N_12048,N_12199);
or U12595 (N_12595,N_12327,N_12182);
or U12596 (N_12596,N_12092,N_12078);
or U12597 (N_12597,N_12471,N_12082);
nor U12598 (N_12598,N_12083,N_12259);
or U12599 (N_12599,N_12401,N_12321);
nand U12600 (N_12600,N_12165,N_12352);
or U12601 (N_12601,N_12061,N_12136);
nand U12602 (N_12602,N_12347,N_12129);
nand U12603 (N_12603,N_12006,N_12212);
nor U12604 (N_12604,N_12008,N_12329);
or U12605 (N_12605,N_12173,N_12416);
nand U12606 (N_12606,N_12311,N_12408);
nand U12607 (N_12607,N_12110,N_12465);
or U12608 (N_12608,N_12445,N_12029);
nor U12609 (N_12609,N_12451,N_12463);
xnor U12610 (N_12610,N_12200,N_12290);
nand U12611 (N_12611,N_12045,N_12337);
and U12612 (N_12612,N_12309,N_12460);
or U12613 (N_12613,N_12188,N_12034);
xnor U12614 (N_12614,N_12147,N_12066);
or U12615 (N_12615,N_12489,N_12323);
nor U12616 (N_12616,N_12456,N_12307);
nor U12617 (N_12617,N_12495,N_12426);
or U12618 (N_12618,N_12095,N_12134);
nand U12619 (N_12619,N_12184,N_12084);
or U12620 (N_12620,N_12256,N_12096);
nor U12621 (N_12621,N_12196,N_12238);
or U12622 (N_12622,N_12269,N_12482);
xor U12623 (N_12623,N_12442,N_12225);
nor U12624 (N_12624,N_12208,N_12490);
or U12625 (N_12625,N_12399,N_12427);
or U12626 (N_12626,N_12414,N_12067);
nor U12627 (N_12627,N_12380,N_12430);
and U12628 (N_12628,N_12077,N_12218);
or U12629 (N_12629,N_12042,N_12332);
nand U12630 (N_12630,N_12353,N_12059);
nand U12631 (N_12631,N_12039,N_12375);
and U12632 (N_12632,N_12341,N_12156);
or U12633 (N_12633,N_12449,N_12201);
nand U12634 (N_12634,N_12496,N_12491);
and U12635 (N_12635,N_12298,N_12180);
and U12636 (N_12636,N_12192,N_12484);
and U12637 (N_12637,N_12237,N_12475);
and U12638 (N_12638,N_12118,N_12013);
or U12639 (N_12639,N_12224,N_12216);
or U12640 (N_12640,N_12308,N_12153);
xor U12641 (N_12641,N_12018,N_12359);
or U12642 (N_12642,N_12021,N_12028);
xnor U12643 (N_12643,N_12488,N_12458);
nor U12644 (N_12644,N_12289,N_12124);
or U12645 (N_12645,N_12400,N_12304);
nor U12646 (N_12646,N_12074,N_12087);
and U12647 (N_12647,N_12470,N_12418);
or U12648 (N_12648,N_12009,N_12455);
nor U12649 (N_12649,N_12204,N_12361);
xnor U12650 (N_12650,N_12385,N_12405);
or U12651 (N_12651,N_12301,N_12486);
and U12652 (N_12652,N_12425,N_12299);
nor U12653 (N_12653,N_12403,N_12297);
xnor U12654 (N_12654,N_12164,N_12079);
and U12655 (N_12655,N_12393,N_12389);
nand U12656 (N_12656,N_12169,N_12366);
or U12657 (N_12657,N_12253,N_12194);
and U12658 (N_12658,N_12415,N_12384);
nand U12659 (N_12659,N_12240,N_12245);
nor U12660 (N_12660,N_12260,N_12440);
nand U12661 (N_12661,N_12191,N_12144);
and U12662 (N_12662,N_12448,N_12333);
nand U12663 (N_12663,N_12314,N_12203);
and U12664 (N_12664,N_12420,N_12127);
nand U12665 (N_12665,N_12158,N_12268);
nand U12666 (N_12666,N_12197,N_12435);
and U12667 (N_12667,N_12172,N_12076);
nor U12668 (N_12668,N_12181,N_12462);
nand U12669 (N_12669,N_12305,N_12109);
and U12670 (N_12670,N_12139,N_12183);
xor U12671 (N_12671,N_12334,N_12364);
xor U12672 (N_12672,N_12326,N_12428);
nor U12673 (N_12673,N_12494,N_12050);
or U12674 (N_12674,N_12014,N_12454);
xor U12675 (N_12675,N_12177,N_12001);
xor U12676 (N_12676,N_12376,N_12349);
or U12677 (N_12677,N_12377,N_12261);
and U12678 (N_12678,N_12336,N_12281);
or U12679 (N_12679,N_12394,N_12073);
and U12680 (N_12680,N_12358,N_12103);
nand U12681 (N_12681,N_12468,N_12154);
and U12682 (N_12682,N_12372,N_12062);
or U12683 (N_12683,N_12007,N_12497);
or U12684 (N_12684,N_12093,N_12111);
or U12685 (N_12685,N_12189,N_12379);
nand U12686 (N_12686,N_12186,N_12120);
xor U12687 (N_12687,N_12360,N_12152);
and U12688 (N_12688,N_12002,N_12283);
nand U12689 (N_12689,N_12088,N_12317);
or U12690 (N_12690,N_12168,N_12037);
or U12691 (N_12691,N_12230,N_12125);
or U12692 (N_12692,N_12233,N_12081);
or U12693 (N_12693,N_12130,N_12243);
nor U12694 (N_12694,N_12331,N_12264);
nand U12695 (N_12695,N_12068,N_12457);
nand U12696 (N_12696,N_12252,N_12251);
nor U12697 (N_12697,N_12138,N_12274);
nand U12698 (N_12698,N_12174,N_12388);
and U12699 (N_12699,N_12402,N_12086);
or U12700 (N_12700,N_12342,N_12150);
nor U12701 (N_12701,N_12444,N_12228);
and U12702 (N_12702,N_12278,N_12262);
and U12703 (N_12703,N_12480,N_12089);
nor U12704 (N_12704,N_12106,N_12406);
or U12705 (N_12705,N_12117,N_12386);
and U12706 (N_12706,N_12263,N_12026);
nor U12707 (N_12707,N_12108,N_12149);
and U12708 (N_12708,N_12051,N_12159);
nand U12709 (N_12709,N_12057,N_12226);
and U12710 (N_12710,N_12285,N_12363);
or U12711 (N_12711,N_12097,N_12499);
or U12712 (N_12712,N_12032,N_12374);
nor U12713 (N_12713,N_12320,N_12202);
nor U12714 (N_12714,N_12276,N_12267);
nand U12715 (N_12715,N_12166,N_12126);
and U12716 (N_12716,N_12476,N_12419);
nand U12717 (N_12717,N_12041,N_12273);
nand U12718 (N_12718,N_12234,N_12075);
xor U12719 (N_12719,N_12322,N_12421);
or U12720 (N_12720,N_12265,N_12296);
nor U12721 (N_12721,N_12288,N_12022);
nor U12722 (N_12722,N_12452,N_12246);
and U12723 (N_12723,N_12302,N_12381);
nor U12724 (N_12724,N_12099,N_12293);
nor U12725 (N_12725,N_12396,N_12450);
nor U12726 (N_12726,N_12397,N_12424);
nand U12727 (N_12727,N_12027,N_12038);
xor U12728 (N_12728,N_12286,N_12115);
xnor U12729 (N_12729,N_12306,N_12025);
xor U12730 (N_12730,N_12023,N_12162);
nand U12731 (N_12731,N_12206,N_12185);
or U12732 (N_12732,N_12438,N_12328);
nand U12733 (N_12733,N_12132,N_12140);
nor U12734 (N_12734,N_12300,N_12292);
nand U12735 (N_12735,N_12210,N_12052);
nand U12736 (N_12736,N_12493,N_12060);
xnor U12737 (N_12737,N_12498,N_12004);
xor U12738 (N_12738,N_12447,N_12232);
and U12739 (N_12739,N_12213,N_12423);
nand U12740 (N_12740,N_12429,N_12054);
or U12741 (N_12741,N_12143,N_12409);
xnor U12742 (N_12742,N_12270,N_12466);
xnor U12743 (N_12743,N_12294,N_12101);
and U12744 (N_12744,N_12291,N_12254);
xor U12745 (N_12745,N_12443,N_12090);
and U12746 (N_12746,N_12282,N_12046);
nor U12747 (N_12747,N_12098,N_12205);
or U12748 (N_12748,N_12303,N_12236);
or U12749 (N_12749,N_12280,N_12459);
xnor U12750 (N_12750,N_12261,N_12155);
or U12751 (N_12751,N_12046,N_12017);
or U12752 (N_12752,N_12166,N_12379);
and U12753 (N_12753,N_12000,N_12107);
and U12754 (N_12754,N_12005,N_12484);
nand U12755 (N_12755,N_12290,N_12149);
and U12756 (N_12756,N_12352,N_12093);
and U12757 (N_12757,N_12158,N_12480);
nor U12758 (N_12758,N_12120,N_12414);
nor U12759 (N_12759,N_12442,N_12317);
nor U12760 (N_12760,N_12200,N_12381);
xnor U12761 (N_12761,N_12366,N_12053);
or U12762 (N_12762,N_12042,N_12218);
nand U12763 (N_12763,N_12071,N_12331);
nand U12764 (N_12764,N_12222,N_12290);
and U12765 (N_12765,N_12349,N_12388);
nor U12766 (N_12766,N_12439,N_12321);
xnor U12767 (N_12767,N_12121,N_12357);
xnor U12768 (N_12768,N_12368,N_12064);
and U12769 (N_12769,N_12391,N_12166);
xnor U12770 (N_12770,N_12024,N_12266);
or U12771 (N_12771,N_12433,N_12000);
nor U12772 (N_12772,N_12314,N_12180);
nand U12773 (N_12773,N_12041,N_12244);
or U12774 (N_12774,N_12211,N_12275);
or U12775 (N_12775,N_12266,N_12351);
xor U12776 (N_12776,N_12380,N_12006);
and U12777 (N_12777,N_12288,N_12283);
nor U12778 (N_12778,N_12339,N_12189);
and U12779 (N_12779,N_12409,N_12181);
or U12780 (N_12780,N_12008,N_12254);
nand U12781 (N_12781,N_12097,N_12218);
and U12782 (N_12782,N_12451,N_12371);
xor U12783 (N_12783,N_12049,N_12012);
nand U12784 (N_12784,N_12002,N_12480);
nand U12785 (N_12785,N_12474,N_12401);
or U12786 (N_12786,N_12163,N_12459);
nand U12787 (N_12787,N_12455,N_12151);
xnor U12788 (N_12788,N_12219,N_12476);
and U12789 (N_12789,N_12122,N_12056);
and U12790 (N_12790,N_12163,N_12265);
and U12791 (N_12791,N_12424,N_12245);
or U12792 (N_12792,N_12123,N_12146);
nor U12793 (N_12793,N_12020,N_12382);
and U12794 (N_12794,N_12036,N_12429);
or U12795 (N_12795,N_12375,N_12385);
nand U12796 (N_12796,N_12164,N_12136);
and U12797 (N_12797,N_12491,N_12071);
or U12798 (N_12798,N_12328,N_12107);
and U12799 (N_12799,N_12057,N_12259);
nor U12800 (N_12800,N_12382,N_12479);
xnor U12801 (N_12801,N_12117,N_12002);
nand U12802 (N_12802,N_12253,N_12293);
nand U12803 (N_12803,N_12164,N_12261);
and U12804 (N_12804,N_12011,N_12140);
or U12805 (N_12805,N_12152,N_12370);
nor U12806 (N_12806,N_12242,N_12318);
xor U12807 (N_12807,N_12352,N_12062);
nor U12808 (N_12808,N_12475,N_12236);
nor U12809 (N_12809,N_12181,N_12177);
nand U12810 (N_12810,N_12389,N_12117);
nand U12811 (N_12811,N_12020,N_12362);
nand U12812 (N_12812,N_12161,N_12312);
and U12813 (N_12813,N_12212,N_12093);
and U12814 (N_12814,N_12341,N_12489);
nand U12815 (N_12815,N_12247,N_12019);
or U12816 (N_12816,N_12266,N_12227);
nand U12817 (N_12817,N_12093,N_12008);
or U12818 (N_12818,N_12087,N_12475);
and U12819 (N_12819,N_12305,N_12296);
nand U12820 (N_12820,N_12366,N_12061);
nand U12821 (N_12821,N_12391,N_12440);
nor U12822 (N_12822,N_12223,N_12198);
or U12823 (N_12823,N_12358,N_12373);
nand U12824 (N_12824,N_12397,N_12343);
or U12825 (N_12825,N_12220,N_12127);
nand U12826 (N_12826,N_12314,N_12292);
nand U12827 (N_12827,N_12362,N_12237);
and U12828 (N_12828,N_12249,N_12427);
or U12829 (N_12829,N_12422,N_12201);
nand U12830 (N_12830,N_12403,N_12150);
xor U12831 (N_12831,N_12330,N_12474);
xor U12832 (N_12832,N_12435,N_12182);
or U12833 (N_12833,N_12090,N_12284);
and U12834 (N_12834,N_12328,N_12026);
xor U12835 (N_12835,N_12406,N_12024);
and U12836 (N_12836,N_12145,N_12462);
or U12837 (N_12837,N_12047,N_12134);
or U12838 (N_12838,N_12446,N_12085);
nand U12839 (N_12839,N_12324,N_12288);
nand U12840 (N_12840,N_12270,N_12027);
or U12841 (N_12841,N_12083,N_12135);
xor U12842 (N_12842,N_12180,N_12329);
or U12843 (N_12843,N_12111,N_12230);
and U12844 (N_12844,N_12075,N_12374);
or U12845 (N_12845,N_12290,N_12257);
nor U12846 (N_12846,N_12174,N_12010);
xor U12847 (N_12847,N_12370,N_12341);
nand U12848 (N_12848,N_12381,N_12030);
or U12849 (N_12849,N_12095,N_12455);
nor U12850 (N_12850,N_12043,N_12374);
nand U12851 (N_12851,N_12319,N_12060);
nand U12852 (N_12852,N_12473,N_12000);
xor U12853 (N_12853,N_12165,N_12108);
xnor U12854 (N_12854,N_12066,N_12269);
or U12855 (N_12855,N_12404,N_12418);
nor U12856 (N_12856,N_12334,N_12232);
xor U12857 (N_12857,N_12224,N_12110);
xnor U12858 (N_12858,N_12383,N_12153);
or U12859 (N_12859,N_12282,N_12171);
xor U12860 (N_12860,N_12129,N_12457);
and U12861 (N_12861,N_12198,N_12002);
or U12862 (N_12862,N_12219,N_12101);
nor U12863 (N_12863,N_12308,N_12290);
or U12864 (N_12864,N_12368,N_12425);
nor U12865 (N_12865,N_12349,N_12273);
nor U12866 (N_12866,N_12452,N_12359);
xnor U12867 (N_12867,N_12273,N_12042);
or U12868 (N_12868,N_12398,N_12191);
nand U12869 (N_12869,N_12134,N_12023);
xor U12870 (N_12870,N_12011,N_12166);
xnor U12871 (N_12871,N_12354,N_12420);
nor U12872 (N_12872,N_12367,N_12301);
nand U12873 (N_12873,N_12147,N_12262);
nand U12874 (N_12874,N_12015,N_12427);
and U12875 (N_12875,N_12477,N_12374);
nor U12876 (N_12876,N_12438,N_12167);
or U12877 (N_12877,N_12405,N_12382);
and U12878 (N_12878,N_12058,N_12420);
xor U12879 (N_12879,N_12335,N_12223);
xor U12880 (N_12880,N_12059,N_12174);
xnor U12881 (N_12881,N_12057,N_12134);
nor U12882 (N_12882,N_12062,N_12357);
or U12883 (N_12883,N_12279,N_12447);
and U12884 (N_12884,N_12227,N_12265);
xor U12885 (N_12885,N_12229,N_12374);
or U12886 (N_12886,N_12006,N_12443);
or U12887 (N_12887,N_12236,N_12330);
and U12888 (N_12888,N_12365,N_12401);
nor U12889 (N_12889,N_12453,N_12410);
or U12890 (N_12890,N_12223,N_12468);
or U12891 (N_12891,N_12473,N_12449);
nor U12892 (N_12892,N_12182,N_12024);
or U12893 (N_12893,N_12250,N_12009);
xor U12894 (N_12894,N_12178,N_12003);
xnor U12895 (N_12895,N_12485,N_12201);
or U12896 (N_12896,N_12497,N_12439);
nor U12897 (N_12897,N_12131,N_12322);
xnor U12898 (N_12898,N_12265,N_12340);
and U12899 (N_12899,N_12469,N_12427);
or U12900 (N_12900,N_12027,N_12126);
nor U12901 (N_12901,N_12295,N_12456);
nor U12902 (N_12902,N_12254,N_12463);
nor U12903 (N_12903,N_12301,N_12072);
nand U12904 (N_12904,N_12004,N_12362);
nand U12905 (N_12905,N_12216,N_12330);
and U12906 (N_12906,N_12410,N_12070);
xor U12907 (N_12907,N_12473,N_12210);
xnor U12908 (N_12908,N_12235,N_12011);
xor U12909 (N_12909,N_12440,N_12426);
xnor U12910 (N_12910,N_12018,N_12120);
or U12911 (N_12911,N_12095,N_12053);
and U12912 (N_12912,N_12242,N_12285);
and U12913 (N_12913,N_12297,N_12319);
nand U12914 (N_12914,N_12224,N_12009);
xnor U12915 (N_12915,N_12319,N_12392);
nand U12916 (N_12916,N_12351,N_12422);
or U12917 (N_12917,N_12113,N_12107);
or U12918 (N_12918,N_12295,N_12318);
nor U12919 (N_12919,N_12165,N_12422);
xnor U12920 (N_12920,N_12145,N_12033);
nand U12921 (N_12921,N_12034,N_12189);
or U12922 (N_12922,N_12127,N_12184);
nor U12923 (N_12923,N_12340,N_12475);
nor U12924 (N_12924,N_12243,N_12044);
nand U12925 (N_12925,N_12274,N_12259);
xor U12926 (N_12926,N_12428,N_12131);
nand U12927 (N_12927,N_12185,N_12404);
nand U12928 (N_12928,N_12306,N_12117);
and U12929 (N_12929,N_12163,N_12039);
or U12930 (N_12930,N_12384,N_12478);
nor U12931 (N_12931,N_12416,N_12337);
or U12932 (N_12932,N_12277,N_12413);
or U12933 (N_12933,N_12083,N_12188);
and U12934 (N_12934,N_12053,N_12198);
nand U12935 (N_12935,N_12418,N_12308);
nor U12936 (N_12936,N_12271,N_12149);
xor U12937 (N_12937,N_12217,N_12260);
nor U12938 (N_12938,N_12174,N_12233);
nor U12939 (N_12939,N_12280,N_12335);
and U12940 (N_12940,N_12261,N_12179);
and U12941 (N_12941,N_12254,N_12104);
and U12942 (N_12942,N_12090,N_12039);
nand U12943 (N_12943,N_12120,N_12173);
xnor U12944 (N_12944,N_12453,N_12496);
and U12945 (N_12945,N_12037,N_12009);
and U12946 (N_12946,N_12427,N_12342);
nor U12947 (N_12947,N_12431,N_12275);
and U12948 (N_12948,N_12325,N_12166);
xor U12949 (N_12949,N_12258,N_12324);
or U12950 (N_12950,N_12255,N_12160);
xor U12951 (N_12951,N_12223,N_12349);
nand U12952 (N_12952,N_12399,N_12030);
or U12953 (N_12953,N_12382,N_12374);
xnor U12954 (N_12954,N_12458,N_12150);
xnor U12955 (N_12955,N_12068,N_12474);
xor U12956 (N_12956,N_12188,N_12236);
nand U12957 (N_12957,N_12363,N_12069);
or U12958 (N_12958,N_12354,N_12103);
xor U12959 (N_12959,N_12206,N_12410);
or U12960 (N_12960,N_12397,N_12483);
or U12961 (N_12961,N_12421,N_12295);
nand U12962 (N_12962,N_12454,N_12389);
xor U12963 (N_12963,N_12444,N_12047);
nor U12964 (N_12964,N_12036,N_12475);
nand U12965 (N_12965,N_12227,N_12018);
or U12966 (N_12966,N_12316,N_12045);
or U12967 (N_12967,N_12340,N_12351);
nand U12968 (N_12968,N_12481,N_12065);
and U12969 (N_12969,N_12086,N_12423);
and U12970 (N_12970,N_12236,N_12309);
nor U12971 (N_12971,N_12466,N_12261);
nor U12972 (N_12972,N_12350,N_12216);
and U12973 (N_12973,N_12428,N_12034);
nor U12974 (N_12974,N_12442,N_12345);
nor U12975 (N_12975,N_12448,N_12217);
nand U12976 (N_12976,N_12370,N_12018);
nor U12977 (N_12977,N_12132,N_12279);
or U12978 (N_12978,N_12495,N_12014);
or U12979 (N_12979,N_12230,N_12112);
or U12980 (N_12980,N_12210,N_12434);
nand U12981 (N_12981,N_12447,N_12223);
nor U12982 (N_12982,N_12453,N_12268);
nand U12983 (N_12983,N_12383,N_12299);
xor U12984 (N_12984,N_12417,N_12205);
nand U12985 (N_12985,N_12018,N_12471);
nor U12986 (N_12986,N_12211,N_12340);
nand U12987 (N_12987,N_12205,N_12185);
xnor U12988 (N_12988,N_12393,N_12171);
nor U12989 (N_12989,N_12258,N_12078);
and U12990 (N_12990,N_12192,N_12401);
and U12991 (N_12991,N_12014,N_12222);
and U12992 (N_12992,N_12403,N_12375);
or U12993 (N_12993,N_12410,N_12098);
and U12994 (N_12994,N_12420,N_12474);
and U12995 (N_12995,N_12447,N_12347);
or U12996 (N_12996,N_12045,N_12225);
nand U12997 (N_12997,N_12012,N_12110);
and U12998 (N_12998,N_12458,N_12307);
xor U12999 (N_12999,N_12159,N_12464);
and U13000 (N_13000,N_12966,N_12786);
xor U13001 (N_13001,N_12736,N_12514);
xnor U13002 (N_13002,N_12944,N_12856);
or U13003 (N_13003,N_12679,N_12564);
nor U13004 (N_13004,N_12763,N_12882);
nor U13005 (N_13005,N_12577,N_12951);
nand U13006 (N_13006,N_12542,N_12698);
xor U13007 (N_13007,N_12629,N_12847);
nor U13008 (N_13008,N_12541,N_12999);
nor U13009 (N_13009,N_12625,N_12669);
nor U13010 (N_13010,N_12920,N_12568);
or U13011 (N_13011,N_12503,N_12653);
or U13012 (N_13012,N_12533,N_12605);
or U13013 (N_13013,N_12659,N_12774);
xnor U13014 (N_13014,N_12798,N_12628);
and U13015 (N_13015,N_12502,N_12796);
and U13016 (N_13016,N_12905,N_12612);
or U13017 (N_13017,N_12917,N_12753);
xnor U13018 (N_13018,N_12545,N_12543);
and U13019 (N_13019,N_12616,N_12525);
nor U13020 (N_13020,N_12903,N_12715);
nor U13021 (N_13021,N_12692,N_12797);
nor U13022 (N_13022,N_12752,N_12948);
nor U13023 (N_13023,N_12734,N_12892);
or U13024 (N_13024,N_12881,N_12800);
and U13025 (N_13025,N_12650,N_12821);
xor U13026 (N_13026,N_12932,N_12997);
nor U13027 (N_13027,N_12654,N_12695);
nand U13028 (N_13028,N_12936,N_12744);
and U13029 (N_13029,N_12524,N_12619);
or U13030 (N_13030,N_12947,N_12730);
xor U13031 (N_13031,N_12704,N_12805);
or U13032 (N_13032,N_12647,N_12762);
nand U13033 (N_13033,N_12773,N_12964);
or U13034 (N_13034,N_12998,N_12842);
and U13035 (N_13035,N_12615,N_12671);
or U13036 (N_13036,N_12632,N_12924);
or U13037 (N_13037,N_12833,N_12517);
and U13038 (N_13038,N_12575,N_12723);
nand U13039 (N_13039,N_12927,N_12759);
xor U13040 (N_13040,N_12790,N_12553);
nor U13041 (N_13041,N_12521,N_12626);
and U13042 (N_13042,N_12957,N_12931);
xnor U13043 (N_13043,N_12620,N_12583);
xor U13044 (N_13044,N_12703,N_12571);
and U13045 (N_13045,N_12883,N_12858);
xor U13046 (N_13046,N_12781,N_12635);
xor U13047 (N_13047,N_12642,N_12665);
xnor U13048 (N_13048,N_12634,N_12572);
xnor U13049 (N_13049,N_12649,N_12540);
and U13050 (N_13050,N_12535,N_12828);
and U13051 (N_13051,N_12561,N_12707);
and U13052 (N_13052,N_12587,N_12676);
xor U13053 (N_13053,N_12900,N_12868);
or U13054 (N_13054,N_12969,N_12600);
and U13055 (N_13055,N_12806,N_12861);
and U13056 (N_13056,N_12559,N_12501);
nor U13057 (N_13057,N_12973,N_12611);
nand U13058 (N_13058,N_12511,N_12689);
nor U13059 (N_13059,N_12850,N_12808);
nor U13060 (N_13060,N_12918,N_12618);
and U13061 (N_13061,N_12954,N_12563);
or U13062 (N_13062,N_12739,N_12764);
nand U13063 (N_13063,N_12767,N_12547);
xor U13064 (N_13064,N_12636,N_12557);
xor U13065 (N_13065,N_12896,N_12777);
xor U13066 (N_13066,N_12562,N_12934);
or U13067 (N_13067,N_12990,N_12826);
nand U13068 (N_13068,N_12757,N_12804);
and U13069 (N_13069,N_12522,N_12725);
or U13070 (N_13070,N_12724,N_12694);
xor U13071 (N_13071,N_12652,N_12586);
xor U13072 (N_13072,N_12803,N_12980);
and U13073 (N_13073,N_12766,N_12565);
and U13074 (N_13074,N_12686,N_12729);
and U13075 (N_13075,N_12728,N_12656);
xnor U13076 (N_13076,N_12749,N_12841);
nand U13077 (N_13077,N_12961,N_12529);
nor U13078 (N_13078,N_12959,N_12640);
nand U13079 (N_13079,N_12809,N_12621);
nand U13080 (N_13080,N_12945,N_12670);
nand U13081 (N_13081,N_12641,N_12672);
nand U13082 (N_13082,N_12580,N_12899);
nand U13083 (N_13083,N_12791,N_12995);
nand U13084 (N_13084,N_12885,N_12817);
nor U13085 (N_13085,N_12977,N_12911);
or U13086 (N_13086,N_12538,N_12741);
nand U13087 (N_13087,N_12705,N_12507);
or U13088 (N_13088,N_12779,N_12527);
and U13089 (N_13089,N_12732,N_12960);
and U13090 (N_13090,N_12550,N_12633);
and U13091 (N_13091,N_12500,N_12607);
or U13092 (N_13092,N_12875,N_12992);
nand U13093 (N_13093,N_12539,N_12727);
xnor U13094 (N_13094,N_12836,N_12567);
xnor U13095 (N_13095,N_12520,N_12528);
xnor U13096 (N_13096,N_12716,N_12878);
or U13097 (N_13097,N_12589,N_12512);
nor U13098 (N_13098,N_12776,N_12747);
xnor U13099 (N_13099,N_12737,N_12505);
and U13100 (N_13100,N_12504,N_12816);
nor U13101 (N_13101,N_12590,N_12854);
xor U13102 (N_13102,N_12802,N_12637);
xor U13103 (N_13103,N_12735,N_12606);
xor U13104 (N_13104,N_12518,N_12989);
nor U13105 (N_13105,N_12601,N_12687);
nand U13106 (N_13106,N_12846,N_12921);
or U13107 (N_13107,N_12617,N_12596);
nand U13108 (N_13108,N_12783,N_12784);
xnor U13109 (N_13109,N_12799,N_12748);
and U13110 (N_13110,N_12860,N_12987);
xnor U13111 (N_13111,N_12793,N_12866);
nand U13112 (N_13112,N_12840,N_12971);
nor U13113 (N_13113,N_12982,N_12949);
and U13114 (N_13114,N_12834,N_12699);
nor U13115 (N_13115,N_12985,N_12785);
or U13116 (N_13116,N_12714,N_12674);
nor U13117 (N_13117,N_12581,N_12720);
xnor U13118 (N_13118,N_12801,N_12693);
and U13119 (N_13119,N_12942,N_12579);
xnor U13120 (N_13120,N_12662,N_12886);
and U13121 (N_13121,N_12974,N_12782);
and U13122 (N_13122,N_12991,N_12677);
and U13123 (N_13123,N_12682,N_12754);
and U13124 (N_13124,N_12691,N_12509);
or U13125 (N_13125,N_12609,N_12895);
nor U13126 (N_13126,N_12893,N_12830);
nor U13127 (N_13127,N_12913,N_12852);
xor U13128 (N_13128,N_12717,N_12986);
nor U13129 (N_13129,N_12638,N_12839);
nor U13130 (N_13130,N_12688,N_12523);
nand U13131 (N_13131,N_12645,N_12660);
xor U13132 (N_13132,N_12554,N_12814);
and U13133 (N_13133,N_12743,N_12862);
and U13134 (N_13134,N_12979,N_12812);
nand U13135 (N_13135,N_12576,N_12871);
and U13136 (N_13136,N_12630,N_12941);
nor U13137 (N_13137,N_12702,N_12758);
xnor U13138 (N_13138,N_12769,N_12851);
and U13139 (N_13139,N_12667,N_12938);
xnor U13140 (N_13140,N_12552,N_12910);
xnor U13141 (N_13141,N_12972,N_12962);
and U13142 (N_13142,N_12597,N_12929);
nand U13143 (N_13143,N_12788,N_12914);
nand U13144 (N_13144,N_12558,N_12531);
nor U13145 (N_13145,N_12810,N_12978);
or U13146 (N_13146,N_12516,N_12815);
and U13147 (N_13147,N_12879,N_12746);
and U13148 (N_13148,N_12683,N_12916);
or U13149 (N_13149,N_12891,N_12582);
or U13150 (N_13150,N_12578,N_12646);
nand U13151 (N_13151,N_12874,N_12768);
and U13152 (N_13152,N_12639,N_12820);
xnor U13153 (N_13153,N_12726,N_12819);
nand U13154 (N_13154,N_12952,N_12666);
nor U13155 (N_13155,N_12988,N_12608);
xnor U13156 (N_13156,N_12919,N_12889);
nor U13157 (N_13157,N_12549,N_12775);
nor U13158 (N_13158,N_12718,N_12537);
nand U13159 (N_13159,N_12673,N_12643);
and U13160 (N_13160,N_12937,N_12984);
and U13161 (N_13161,N_12923,N_12623);
xor U13162 (N_13162,N_12664,N_12661);
or U13163 (N_13163,N_12950,N_12551);
nor U13164 (N_13164,N_12844,N_12731);
xor U13165 (N_13165,N_12867,N_12668);
nor U13166 (N_13166,N_12684,N_12901);
and U13167 (N_13167,N_12696,N_12849);
xor U13168 (N_13168,N_12902,N_12701);
nor U13169 (N_13169,N_12711,N_12955);
nor U13170 (N_13170,N_12631,N_12928);
or U13171 (N_13171,N_12888,N_12544);
nor U13172 (N_13172,N_12823,N_12560);
and U13173 (N_13173,N_12930,N_12708);
xnor U13174 (N_13174,N_12872,N_12663);
nand U13175 (N_13175,N_12678,N_12807);
nor U13176 (N_13176,N_12613,N_12648);
and U13177 (N_13177,N_12738,N_12824);
or U13178 (N_13178,N_12644,N_12588);
and U13179 (N_13179,N_12765,N_12651);
or U13180 (N_13180,N_12778,N_12894);
and U13181 (N_13181,N_12865,N_12794);
xnor U13182 (N_13182,N_12943,N_12967);
and U13183 (N_13183,N_12831,N_12710);
and U13184 (N_13184,N_12877,N_12935);
and U13185 (N_13185,N_12602,N_12829);
xnor U13186 (N_13186,N_12904,N_12761);
and U13187 (N_13187,N_12598,N_12864);
or U13188 (N_13188,N_12981,N_12968);
or U13189 (N_13189,N_12870,N_12570);
nand U13190 (N_13190,N_12548,N_12566);
or U13191 (N_13191,N_12912,N_12787);
xor U13192 (N_13192,N_12832,N_12884);
xnor U13193 (N_13193,N_12573,N_12908);
or U13194 (N_13194,N_12515,N_12835);
nand U13195 (N_13195,N_12976,N_12593);
or U13196 (N_13196,N_12965,N_12709);
nand U13197 (N_13197,N_12770,N_12880);
nand U13198 (N_13198,N_12939,N_12780);
nand U13199 (N_13199,N_12855,N_12536);
and U13200 (N_13200,N_12657,N_12771);
nor U13201 (N_13201,N_12933,N_12845);
nor U13202 (N_13202,N_12822,N_12733);
xor U13203 (N_13203,N_12700,N_12772);
xnor U13204 (N_13204,N_12706,N_12655);
nand U13205 (N_13205,N_12690,N_12721);
nand U13206 (N_13206,N_12713,N_12591);
nor U13207 (N_13207,N_12993,N_12750);
nand U13208 (N_13208,N_12996,N_12556);
and U13209 (N_13209,N_12843,N_12745);
or U13210 (N_13210,N_12604,N_12946);
and U13211 (N_13211,N_12574,N_12915);
nand U13212 (N_13212,N_12890,N_12795);
nor U13213 (N_13213,N_12859,N_12624);
xor U13214 (N_13214,N_12584,N_12958);
and U13215 (N_13215,N_12681,N_12756);
nor U13216 (N_13216,N_12680,N_12983);
nor U13217 (N_13217,N_12508,N_12526);
or U13218 (N_13218,N_12848,N_12599);
and U13219 (N_13219,N_12970,N_12789);
nor U13220 (N_13220,N_12585,N_12863);
xnor U13221 (N_13221,N_12658,N_12751);
or U13222 (N_13222,N_12685,N_12837);
or U13223 (N_13223,N_12534,N_12675);
nand U13224 (N_13224,N_12740,N_12510);
or U13225 (N_13225,N_12712,N_12760);
nand U13226 (N_13226,N_12603,N_12627);
nand U13227 (N_13227,N_12742,N_12869);
and U13228 (N_13228,N_12922,N_12594);
nand U13229 (N_13229,N_12595,N_12838);
and U13230 (N_13230,N_12697,N_12506);
or U13231 (N_13231,N_12876,N_12898);
and U13232 (N_13232,N_12906,N_12825);
and U13233 (N_13233,N_12755,N_12975);
and U13234 (N_13234,N_12792,N_12907);
nor U13235 (N_13235,N_12956,N_12530);
nand U13236 (N_13236,N_12963,N_12513);
nor U13237 (N_13237,N_12813,N_12897);
nand U13238 (N_13238,N_12909,N_12622);
nand U13239 (N_13239,N_12953,N_12546);
nor U13240 (N_13240,N_12610,N_12555);
nor U13241 (N_13241,N_12926,N_12592);
and U13242 (N_13242,N_12887,N_12569);
or U13243 (N_13243,N_12827,N_12853);
nand U13244 (N_13244,N_12722,N_12873);
and U13245 (N_13245,N_12857,N_12994);
nor U13246 (N_13246,N_12811,N_12719);
nor U13247 (N_13247,N_12925,N_12532);
nor U13248 (N_13248,N_12614,N_12818);
or U13249 (N_13249,N_12940,N_12519);
nand U13250 (N_13250,N_12767,N_12842);
nor U13251 (N_13251,N_12661,N_12968);
nand U13252 (N_13252,N_12587,N_12554);
or U13253 (N_13253,N_12734,N_12605);
nor U13254 (N_13254,N_12775,N_12607);
and U13255 (N_13255,N_12701,N_12658);
xnor U13256 (N_13256,N_12538,N_12588);
xnor U13257 (N_13257,N_12992,N_12642);
nor U13258 (N_13258,N_12990,N_12748);
nand U13259 (N_13259,N_12569,N_12760);
nor U13260 (N_13260,N_12568,N_12889);
nor U13261 (N_13261,N_12737,N_12886);
nand U13262 (N_13262,N_12854,N_12618);
or U13263 (N_13263,N_12723,N_12869);
or U13264 (N_13264,N_12584,N_12622);
nor U13265 (N_13265,N_12566,N_12612);
or U13266 (N_13266,N_12856,N_12756);
xor U13267 (N_13267,N_12624,N_12881);
or U13268 (N_13268,N_12629,N_12535);
xnor U13269 (N_13269,N_12894,N_12582);
and U13270 (N_13270,N_12686,N_12596);
xnor U13271 (N_13271,N_12727,N_12902);
or U13272 (N_13272,N_12952,N_12625);
nand U13273 (N_13273,N_12909,N_12968);
or U13274 (N_13274,N_12551,N_12558);
and U13275 (N_13275,N_12613,N_12617);
and U13276 (N_13276,N_12857,N_12860);
or U13277 (N_13277,N_12974,N_12964);
xor U13278 (N_13278,N_12759,N_12795);
and U13279 (N_13279,N_12576,N_12910);
xor U13280 (N_13280,N_12715,N_12521);
and U13281 (N_13281,N_12832,N_12757);
nor U13282 (N_13282,N_12645,N_12610);
or U13283 (N_13283,N_12515,N_12657);
xor U13284 (N_13284,N_12678,N_12675);
or U13285 (N_13285,N_12860,N_12780);
nor U13286 (N_13286,N_12931,N_12544);
or U13287 (N_13287,N_12955,N_12813);
xor U13288 (N_13288,N_12975,N_12756);
xor U13289 (N_13289,N_12677,N_12713);
nand U13290 (N_13290,N_12965,N_12755);
nand U13291 (N_13291,N_12762,N_12725);
nor U13292 (N_13292,N_12825,N_12927);
nand U13293 (N_13293,N_12935,N_12944);
and U13294 (N_13294,N_12558,N_12556);
nor U13295 (N_13295,N_12858,N_12561);
xnor U13296 (N_13296,N_12686,N_12955);
nand U13297 (N_13297,N_12624,N_12988);
or U13298 (N_13298,N_12593,N_12599);
xnor U13299 (N_13299,N_12722,N_12984);
xor U13300 (N_13300,N_12703,N_12762);
xor U13301 (N_13301,N_12828,N_12721);
or U13302 (N_13302,N_12970,N_12965);
nor U13303 (N_13303,N_12704,N_12744);
or U13304 (N_13304,N_12829,N_12948);
nor U13305 (N_13305,N_12783,N_12726);
or U13306 (N_13306,N_12646,N_12693);
or U13307 (N_13307,N_12776,N_12570);
xnor U13308 (N_13308,N_12929,N_12656);
xor U13309 (N_13309,N_12755,N_12646);
nor U13310 (N_13310,N_12549,N_12856);
nand U13311 (N_13311,N_12666,N_12675);
xor U13312 (N_13312,N_12693,N_12992);
nor U13313 (N_13313,N_12964,N_12806);
and U13314 (N_13314,N_12611,N_12722);
nand U13315 (N_13315,N_12847,N_12538);
xor U13316 (N_13316,N_12722,N_12529);
xor U13317 (N_13317,N_12832,N_12969);
xor U13318 (N_13318,N_12837,N_12934);
and U13319 (N_13319,N_12964,N_12634);
xnor U13320 (N_13320,N_12778,N_12826);
nand U13321 (N_13321,N_12937,N_12956);
and U13322 (N_13322,N_12973,N_12801);
or U13323 (N_13323,N_12566,N_12795);
xor U13324 (N_13324,N_12895,N_12602);
nor U13325 (N_13325,N_12913,N_12833);
nand U13326 (N_13326,N_12778,N_12814);
or U13327 (N_13327,N_12643,N_12916);
or U13328 (N_13328,N_12950,N_12655);
nand U13329 (N_13329,N_12885,N_12609);
xor U13330 (N_13330,N_12513,N_12798);
nand U13331 (N_13331,N_12721,N_12754);
and U13332 (N_13332,N_12924,N_12567);
xnor U13333 (N_13333,N_12953,N_12843);
nor U13334 (N_13334,N_12690,N_12523);
xor U13335 (N_13335,N_12515,N_12894);
or U13336 (N_13336,N_12570,N_12716);
nor U13337 (N_13337,N_12525,N_12929);
nand U13338 (N_13338,N_12768,N_12567);
or U13339 (N_13339,N_12975,N_12972);
nor U13340 (N_13340,N_12713,N_12887);
and U13341 (N_13341,N_12566,N_12768);
or U13342 (N_13342,N_12551,N_12884);
nor U13343 (N_13343,N_12591,N_12874);
xnor U13344 (N_13344,N_12934,N_12526);
and U13345 (N_13345,N_12770,N_12866);
or U13346 (N_13346,N_12773,N_12553);
nor U13347 (N_13347,N_12661,N_12604);
xnor U13348 (N_13348,N_12870,N_12896);
or U13349 (N_13349,N_12575,N_12708);
nor U13350 (N_13350,N_12533,N_12637);
or U13351 (N_13351,N_12799,N_12640);
xor U13352 (N_13352,N_12649,N_12959);
nor U13353 (N_13353,N_12617,N_12586);
nor U13354 (N_13354,N_12944,N_12747);
nand U13355 (N_13355,N_12977,N_12913);
xnor U13356 (N_13356,N_12945,N_12842);
or U13357 (N_13357,N_12651,N_12976);
nor U13358 (N_13358,N_12870,N_12923);
and U13359 (N_13359,N_12567,N_12812);
or U13360 (N_13360,N_12612,N_12912);
xor U13361 (N_13361,N_12848,N_12681);
nor U13362 (N_13362,N_12684,N_12827);
nor U13363 (N_13363,N_12873,N_12934);
or U13364 (N_13364,N_12642,N_12673);
and U13365 (N_13365,N_12912,N_12934);
xor U13366 (N_13366,N_12534,N_12777);
and U13367 (N_13367,N_12844,N_12728);
or U13368 (N_13368,N_12541,N_12954);
or U13369 (N_13369,N_12851,N_12723);
xor U13370 (N_13370,N_12949,N_12935);
nand U13371 (N_13371,N_12869,N_12841);
or U13372 (N_13372,N_12735,N_12763);
nand U13373 (N_13373,N_12695,N_12836);
nor U13374 (N_13374,N_12965,N_12895);
and U13375 (N_13375,N_12965,N_12825);
xor U13376 (N_13376,N_12923,N_12757);
nor U13377 (N_13377,N_12682,N_12880);
or U13378 (N_13378,N_12600,N_12865);
nor U13379 (N_13379,N_12750,N_12567);
nor U13380 (N_13380,N_12505,N_12509);
nor U13381 (N_13381,N_12686,N_12932);
xnor U13382 (N_13382,N_12522,N_12979);
and U13383 (N_13383,N_12684,N_12599);
xnor U13384 (N_13384,N_12666,N_12997);
nand U13385 (N_13385,N_12588,N_12843);
xor U13386 (N_13386,N_12702,N_12945);
nand U13387 (N_13387,N_12962,N_12873);
and U13388 (N_13388,N_12683,N_12694);
or U13389 (N_13389,N_12600,N_12803);
nand U13390 (N_13390,N_12759,N_12772);
or U13391 (N_13391,N_12659,N_12688);
or U13392 (N_13392,N_12709,N_12585);
xor U13393 (N_13393,N_12712,N_12555);
or U13394 (N_13394,N_12552,N_12647);
xor U13395 (N_13395,N_12626,N_12766);
or U13396 (N_13396,N_12824,N_12744);
nand U13397 (N_13397,N_12809,N_12725);
and U13398 (N_13398,N_12746,N_12515);
or U13399 (N_13399,N_12505,N_12759);
nand U13400 (N_13400,N_12695,N_12807);
xnor U13401 (N_13401,N_12930,N_12911);
and U13402 (N_13402,N_12943,N_12792);
xnor U13403 (N_13403,N_12992,N_12650);
xnor U13404 (N_13404,N_12962,N_12510);
or U13405 (N_13405,N_12576,N_12880);
nor U13406 (N_13406,N_12910,N_12709);
xor U13407 (N_13407,N_12721,N_12854);
and U13408 (N_13408,N_12948,N_12868);
nor U13409 (N_13409,N_12828,N_12776);
nor U13410 (N_13410,N_12706,N_12563);
or U13411 (N_13411,N_12855,N_12520);
nand U13412 (N_13412,N_12810,N_12797);
nor U13413 (N_13413,N_12943,N_12634);
nor U13414 (N_13414,N_12699,N_12609);
and U13415 (N_13415,N_12557,N_12988);
nor U13416 (N_13416,N_12765,N_12865);
nor U13417 (N_13417,N_12959,N_12604);
or U13418 (N_13418,N_12570,N_12999);
or U13419 (N_13419,N_12659,N_12611);
nor U13420 (N_13420,N_12654,N_12503);
and U13421 (N_13421,N_12672,N_12620);
xor U13422 (N_13422,N_12944,N_12673);
and U13423 (N_13423,N_12910,N_12638);
nand U13424 (N_13424,N_12683,N_12887);
xnor U13425 (N_13425,N_12532,N_12542);
nor U13426 (N_13426,N_12587,N_12671);
xor U13427 (N_13427,N_12640,N_12901);
xnor U13428 (N_13428,N_12715,N_12581);
nand U13429 (N_13429,N_12523,N_12528);
and U13430 (N_13430,N_12872,N_12990);
nand U13431 (N_13431,N_12755,N_12503);
nand U13432 (N_13432,N_12721,N_12934);
nand U13433 (N_13433,N_12671,N_12644);
nand U13434 (N_13434,N_12855,N_12807);
and U13435 (N_13435,N_12865,N_12617);
or U13436 (N_13436,N_12535,N_12891);
or U13437 (N_13437,N_12882,N_12612);
or U13438 (N_13438,N_12626,N_12859);
and U13439 (N_13439,N_12516,N_12629);
or U13440 (N_13440,N_12852,N_12939);
xnor U13441 (N_13441,N_12966,N_12971);
and U13442 (N_13442,N_12845,N_12741);
nor U13443 (N_13443,N_12991,N_12535);
nor U13444 (N_13444,N_12830,N_12602);
and U13445 (N_13445,N_12579,N_12673);
or U13446 (N_13446,N_12729,N_12867);
xor U13447 (N_13447,N_12699,N_12882);
nor U13448 (N_13448,N_12547,N_12813);
nand U13449 (N_13449,N_12978,N_12829);
and U13450 (N_13450,N_12905,N_12676);
or U13451 (N_13451,N_12808,N_12654);
and U13452 (N_13452,N_12885,N_12759);
nand U13453 (N_13453,N_12688,N_12630);
or U13454 (N_13454,N_12551,N_12912);
nor U13455 (N_13455,N_12883,N_12932);
and U13456 (N_13456,N_12582,N_12602);
or U13457 (N_13457,N_12778,N_12514);
xor U13458 (N_13458,N_12864,N_12840);
or U13459 (N_13459,N_12573,N_12748);
and U13460 (N_13460,N_12838,N_12565);
and U13461 (N_13461,N_12786,N_12618);
or U13462 (N_13462,N_12694,N_12964);
or U13463 (N_13463,N_12801,N_12798);
xnor U13464 (N_13464,N_12646,N_12893);
xor U13465 (N_13465,N_12968,N_12758);
and U13466 (N_13466,N_12556,N_12956);
and U13467 (N_13467,N_12893,N_12680);
or U13468 (N_13468,N_12647,N_12539);
xor U13469 (N_13469,N_12983,N_12807);
xor U13470 (N_13470,N_12628,N_12817);
or U13471 (N_13471,N_12793,N_12680);
and U13472 (N_13472,N_12879,N_12582);
or U13473 (N_13473,N_12981,N_12620);
and U13474 (N_13474,N_12795,N_12589);
and U13475 (N_13475,N_12988,N_12741);
or U13476 (N_13476,N_12659,N_12835);
and U13477 (N_13477,N_12531,N_12908);
or U13478 (N_13478,N_12791,N_12879);
nor U13479 (N_13479,N_12943,N_12794);
nand U13480 (N_13480,N_12731,N_12635);
or U13481 (N_13481,N_12811,N_12677);
nand U13482 (N_13482,N_12598,N_12641);
nor U13483 (N_13483,N_12922,N_12997);
and U13484 (N_13484,N_12965,N_12772);
or U13485 (N_13485,N_12938,N_12895);
nand U13486 (N_13486,N_12572,N_12954);
or U13487 (N_13487,N_12822,N_12926);
xor U13488 (N_13488,N_12744,N_12974);
nand U13489 (N_13489,N_12836,N_12514);
nand U13490 (N_13490,N_12997,N_12558);
or U13491 (N_13491,N_12564,N_12991);
and U13492 (N_13492,N_12831,N_12626);
nand U13493 (N_13493,N_12986,N_12596);
nor U13494 (N_13494,N_12581,N_12605);
xor U13495 (N_13495,N_12931,N_12968);
nor U13496 (N_13496,N_12905,N_12672);
nand U13497 (N_13497,N_12900,N_12632);
nand U13498 (N_13498,N_12869,N_12904);
nor U13499 (N_13499,N_12819,N_12610);
and U13500 (N_13500,N_13351,N_13409);
and U13501 (N_13501,N_13034,N_13115);
nor U13502 (N_13502,N_13094,N_13460);
nand U13503 (N_13503,N_13314,N_13370);
or U13504 (N_13504,N_13044,N_13407);
nor U13505 (N_13505,N_13096,N_13257);
or U13506 (N_13506,N_13199,N_13219);
nor U13507 (N_13507,N_13089,N_13304);
or U13508 (N_13508,N_13059,N_13374);
or U13509 (N_13509,N_13395,N_13254);
or U13510 (N_13510,N_13321,N_13237);
xor U13511 (N_13511,N_13246,N_13424);
nand U13512 (N_13512,N_13359,N_13426);
nand U13513 (N_13513,N_13099,N_13003);
nor U13514 (N_13514,N_13435,N_13140);
nor U13515 (N_13515,N_13156,N_13436);
or U13516 (N_13516,N_13307,N_13255);
nor U13517 (N_13517,N_13090,N_13129);
xor U13518 (N_13518,N_13079,N_13421);
or U13519 (N_13519,N_13072,N_13406);
or U13520 (N_13520,N_13442,N_13174);
or U13521 (N_13521,N_13142,N_13434);
nand U13522 (N_13522,N_13158,N_13268);
nand U13523 (N_13523,N_13104,N_13371);
xor U13524 (N_13524,N_13009,N_13160);
nor U13525 (N_13525,N_13367,N_13390);
nor U13526 (N_13526,N_13214,N_13282);
and U13527 (N_13527,N_13098,N_13049);
nor U13528 (N_13528,N_13473,N_13499);
nor U13529 (N_13529,N_13283,N_13352);
xnor U13530 (N_13530,N_13339,N_13067);
or U13531 (N_13531,N_13029,N_13083);
or U13532 (N_13532,N_13037,N_13317);
and U13533 (N_13533,N_13392,N_13184);
and U13534 (N_13534,N_13462,N_13244);
nand U13535 (N_13535,N_13335,N_13487);
nand U13536 (N_13536,N_13366,N_13126);
or U13537 (N_13537,N_13386,N_13124);
and U13538 (N_13538,N_13217,N_13313);
nor U13539 (N_13539,N_13302,N_13380);
or U13540 (N_13540,N_13058,N_13311);
nand U13541 (N_13541,N_13060,N_13100);
and U13542 (N_13542,N_13064,N_13391);
nand U13543 (N_13543,N_13484,N_13438);
and U13544 (N_13544,N_13143,N_13312);
or U13545 (N_13545,N_13210,N_13422);
xor U13546 (N_13546,N_13343,N_13284);
nand U13547 (N_13547,N_13485,N_13154);
or U13548 (N_13548,N_13087,N_13136);
or U13549 (N_13549,N_13019,N_13239);
xor U13550 (N_13550,N_13266,N_13014);
or U13551 (N_13551,N_13465,N_13084);
nand U13552 (N_13552,N_13474,N_13057);
nor U13553 (N_13553,N_13111,N_13250);
and U13554 (N_13554,N_13137,N_13112);
nand U13555 (N_13555,N_13103,N_13375);
and U13556 (N_13556,N_13287,N_13444);
xor U13557 (N_13557,N_13320,N_13167);
xor U13558 (N_13558,N_13147,N_13364);
nand U13559 (N_13559,N_13439,N_13001);
nor U13560 (N_13560,N_13027,N_13213);
nand U13561 (N_13561,N_13316,N_13150);
nor U13562 (N_13562,N_13293,N_13216);
and U13563 (N_13563,N_13202,N_13128);
xor U13564 (N_13564,N_13035,N_13412);
or U13565 (N_13565,N_13116,N_13269);
or U13566 (N_13566,N_13233,N_13068);
or U13567 (N_13567,N_13480,N_13220);
xnor U13568 (N_13568,N_13388,N_13069);
and U13569 (N_13569,N_13379,N_13288);
nand U13570 (N_13570,N_13413,N_13030);
and U13571 (N_13571,N_13417,N_13496);
nand U13572 (N_13572,N_13159,N_13240);
nor U13573 (N_13573,N_13145,N_13344);
and U13574 (N_13574,N_13226,N_13455);
or U13575 (N_13575,N_13248,N_13117);
nor U13576 (N_13576,N_13397,N_13222);
xnor U13577 (N_13577,N_13075,N_13324);
or U13578 (N_13578,N_13290,N_13182);
and U13579 (N_13579,N_13401,N_13491);
xor U13580 (N_13580,N_13171,N_13144);
nor U13581 (N_13581,N_13373,N_13251);
and U13582 (N_13582,N_13400,N_13095);
and U13583 (N_13583,N_13356,N_13055);
or U13584 (N_13584,N_13448,N_13038);
or U13585 (N_13585,N_13173,N_13039);
nand U13586 (N_13586,N_13186,N_13082);
xnor U13587 (N_13587,N_13394,N_13271);
or U13588 (N_13588,N_13056,N_13120);
and U13589 (N_13589,N_13309,N_13420);
nor U13590 (N_13590,N_13423,N_13085);
nand U13591 (N_13591,N_13489,N_13497);
xnor U13592 (N_13592,N_13461,N_13478);
nand U13593 (N_13593,N_13361,N_13076);
xor U13594 (N_13594,N_13315,N_13146);
or U13595 (N_13595,N_13358,N_13326);
or U13596 (N_13596,N_13481,N_13322);
nand U13597 (N_13597,N_13236,N_13040);
nand U13598 (N_13598,N_13265,N_13353);
nor U13599 (N_13599,N_13264,N_13050);
or U13600 (N_13600,N_13225,N_13490);
or U13601 (N_13601,N_13139,N_13006);
xor U13602 (N_13602,N_13195,N_13270);
and U13603 (N_13603,N_13091,N_13482);
nand U13604 (N_13604,N_13172,N_13350);
xor U13605 (N_13605,N_13048,N_13041);
and U13606 (N_13606,N_13121,N_13303);
nand U13607 (N_13607,N_13340,N_13242);
nand U13608 (N_13608,N_13215,N_13188);
and U13609 (N_13609,N_13292,N_13410);
or U13610 (N_13610,N_13025,N_13403);
nand U13611 (N_13611,N_13325,N_13336);
and U13612 (N_13612,N_13110,N_13175);
and U13613 (N_13613,N_13308,N_13252);
and U13614 (N_13614,N_13261,N_13472);
nand U13615 (N_13615,N_13052,N_13232);
xor U13616 (N_13616,N_13263,N_13004);
nand U13617 (N_13617,N_13437,N_13164);
nand U13618 (N_13618,N_13342,N_13300);
or U13619 (N_13619,N_13123,N_13127);
or U13620 (N_13620,N_13241,N_13238);
or U13621 (N_13621,N_13152,N_13245);
nand U13622 (N_13622,N_13023,N_13476);
and U13623 (N_13623,N_13278,N_13260);
or U13624 (N_13624,N_13221,N_13341);
and U13625 (N_13625,N_13365,N_13190);
and U13626 (N_13626,N_13494,N_13493);
and U13627 (N_13627,N_13377,N_13185);
xor U13628 (N_13628,N_13405,N_13495);
or U13629 (N_13629,N_13071,N_13475);
and U13630 (N_13630,N_13141,N_13022);
nor U13631 (N_13631,N_13450,N_13196);
or U13632 (N_13632,N_13431,N_13328);
nor U13633 (N_13633,N_13243,N_13452);
or U13634 (N_13634,N_13223,N_13101);
and U13635 (N_13635,N_13181,N_13306);
nor U13636 (N_13636,N_13253,N_13451);
nor U13637 (N_13637,N_13492,N_13433);
nor U13638 (N_13638,N_13273,N_13020);
nor U13639 (N_13639,N_13212,N_13047);
or U13640 (N_13640,N_13053,N_13256);
and U13641 (N_13641,N_13258,N_13446);
nor U13642 (N_13642,N_13227,N_13183);
xnor U13643 (N_13643,N_13419,N_13398);
and U13644 (N_13644,N_13454,N_13418);
nand U13645 (N_13645,N_13319,N_13387);
and U13646 (N_13646,N_13180,N_13017);
or U13647 (N_13647,N_13205,N_13193);
or U13648 (N_13648,N_13203,N_13468);
nand U13649 (N_13649,N_13201,N_13078);
and U13650 (N_13650,N_13280,N_13042);
nand U13651 (N_13651,N_13402,N_13272);
nor U13652 (N_13652,N_13192,N_13362);
or U13653 (N_13653,N_13088,N_13289);
nor U13654 (N_13654,N_13396,N_13153);
and U13655 (N_13655,N_13323,N_13063);
nand U13656 (N_13656,N_13228,N_13330);
xor U13657 (N_13657,N_13125,N_13376);
and U13658 (N_13658,N_13080,N_13310);
or U13659 (N_13659,N_13331,N_13207);
xor U13660 (N_13660,N_13119,N_13333);
xnor U13661 (N_13661,N_13295,N_13337);
nor U13662 (N_13662,N_13285,N_13011);
nand U13663 (N_13663,N_13198,N_13021);
nor U13664 (N_13664,N_13399,N_13262);
or U13665 (N_13665,N_13428,N_13384);
nor U13666 (N_13666,N_13276,N_13133);
nand U13667 (N_13667,N_13334,N_13045);
and U13668 (N_13668,N_13345,N_13447);
and U13669 (N_13669,N_13230,N_13179);
and U13670 (N_13670,N_13176,N_13408);
and U13671 (N_13671,N_13346,N_13281);
and U13672 (N_13672,N_13274,N_13109);
xor U13673 (N_13673,N_13355,N_13389);
or U13674 (N_13674,N_13443,N_13073);
xor U13675 (N_13675,N_13372,N_13368);
xor U13676 (N_13676,N_13329,N_13224);
nand U13677 (N_13677,N_13015,N_13369);
and U13678 (N_13678,N_13032,N_13187);
nor U13679 (N_13679,N_13235,N_13211);
nor U13680 (N_13680,N_13065,N_13477);
and U13681 (N_13681,N_13297,N_13046);
or U13682 (N_13682,N_13024,N_13122);
nand U13683 (N_13683,N_13130,N_13054);
and U13684 (N_13684,N_13275,N_13018);
xor U13685 (N_13685,N_13231,N_13208);
nand U13686 (N_13686,N_13469,N_13301);
xor U13687 (N_13687,N_13005,N_13381);
xnor U13688 (N_13688,N_13411,N_13393);
nor U13689 (N_13689,N_13151,N_13498);
or U13690 (N_13690,N_13028,N_13013);
and U13691 (N_13691,N_13166,N_13385);
xnor U13692 (N_13692,N_13163,N_13070);
nor U13693 (N_13693,N_13286,N_13204);
nand U13694 (N_13694,N_13445,N_13294);
xor U13695 (N_13695,N_13327,N_13108);
xnor U13696 (N_13696,N_13177,N_13354);
nand U13697 (N_13697,N_13197,N_13458);
and U13698 (N_13698,N_13170,N_13031);
and U13699 (N_13699,N_13234,N_13348);
xnor U13700 (N_13700,N_13161,N_13105);
xor U13701 (N_13701,N_13404,N_13149);
and U13702 (N_13702,N_13007,N_13206);
or U13703 (N_13703,N_13277,N_13081);
nor U13704 (N_13704,N_13414,N_13036);
nor U13705 (N_13705,N_13165,N_13459);
nor U13706 (N_13706,N_13092,N_13033);
nand U13707 (N_13707,N_13016,N_13086);
nand U13708 (N_13708,N_13157,N_13132);
and U13709 (N_13709,N_13299,N_13093);
nor U13710 (N_13710,N_13349,N_13382);
or U13711 (N_13711,N_13113,N_13114);
nand U13712 (N_13712,N_13191,N_13415);
nor U13713 (N_13713,N_13357,N_13118);
xor U13714 (N_13714,N_13051,N_13194);
or U13715 (N_13715,N_13135,N_13010);
and U13716 (N_13716,N_13363,N_13077);
nor U13717 (N_13717,N_13483,N_13247);
or U13718 (N_13718,N_13427,N_13026);
and U13719 (N_13719,N_13148,N_13259);
nand U13720 (N_13720,N_13464,N_13457);
nand U13721 (N_13721,N_13162,N_13209);
xnor U13722 (N_13722,N_13383,N_13338);
xnor U13723 (N_13723,N_13066,N_13298);
and U13724 (N_13724,N_13318,N_13043);
and U13725 (N_13725,N_13138,N_13378);
nand U13726 (N_13726,N_13218,N_13467);
and U13727 (N_13727,N_13430,N_13296);
nand U13728 (N_13728,N_13471,N_13168);
nor U13729 (N_13729,N_13305,N_13200);
xnor U13730 (N_13730,N_13347,N_13106);
nand U13731 (N_13731,N_13012,N_13449);
or U13732 (N_13732,N_13102,N_13429);
and U13733 (N_13733,N_13189,N_13008);
nand U13734 (N_13734,N_13061,N_13178);
or U13735 (N_13735,N_13479,N_13229);
xnor U13736 (N_13736,N_13279,N_13002);
and U13737 (N_13737,N_13425,N_13134);
nand U13738 (N_13738,N_13131,N_13267);
xor U13739 (N_13739,N_13456,N_13441);
nand U13740 (N_13740,N_13360,N_13416);
nor U13741 (N_13741,N_13486,N_13097);
nor U13742 (N_13742,N_13155,N_13000);
and U13743 (N_13743,N_13488,N_13249);
xor U13744 (N_13744,N_13453,N_13107);
nand U13745 (N_13745,N_13074,N_13169);
xnor U13746 (N_13746,N_13062,N_13463);
xor U13747 (N_13747,N_13432,N_13440);
nor U13748 (N_13748,N_13332,N_13470);
nor U13749 (N_13749,N_13466,N_13291);
or U13750 (N_13750,N_13189,N_13176);
nand U13751 (N_13751,N_13281,N_13334);
or U13752 (N_13752,N_13358,N_13037);
nand U13753 (N_13753,N_13073,N_13427);
or U13754 (N_13754,N_13314,N_13491);
and U13755 (N_13755,N_13086,N_13164);
nor U13756 (N_13756,N_13357,N_13256);
nor U13757 (N_13757,N_13161,N_13129);
or U13758 (N_13758,N_13353,N_13359);
nand U13759 (N_13759,N_13113,N_13487);
nand U13760 (N_13760,N_13207,N_13220);
nand U13761 (N_13761,N_13016,N_13047);
xnor U13762 (N_13762,N_13487,N_13246);
or U13763 (N_13763,N_13445,N_13158);
nor U13764 (N_13764,N_13388,N_13128);
xnor U13765 (N_13765,N_13293,N_13108);
nand U13766 (N_13766,N_13044,N_13359);
xor U13767 (N_13767,N_13173,N_13018);
nand U13768 (N_13768,N_13090,N_13323);
or U13769 (N_13769,N_13372,N_13130);
or U13770 (N_13770,N_13356,N_13455);
and U13771 (N_13771,N_13006,N_13086);
xor U13772 (N_13772,N_13054,N_13497);
nand U13773 (N_13773,N_13048,N_13180);
nor U13774 (N_13774,N_13214,N_13308);
nand U13775 (N_13775,N_13095,N_13301);
nor U13776 (N_13776,N_13275,N_13444);
nand U13777 (N_13777,N_13348,N_13005);
nor U13778 (N_13778,N_13213,N_13143);
and U13779 (N_13779,N_13272,N_13410);
nor U13780 (N_13780,N_13224,N_13014);
or U13781 (N_13781,N_13091,N_13334);
or U13782 (N_13782,N_13185,N_13301);
and U13783 (N_13783,N_13169,N_13222);
nor U13784 (N_13784,N_13207,N_13349);
nand U13785 (N_13785,N_13276,N_13181);
xor U13786 (N_13786,N_13204,N_13197);
xor U13787 (N_13787,N_13290,N_13070);
xnor U13788 (N_13788,N_13230,N_13409);
xnor U13789 (N_13789,N_13230,N_13259);
xor U13790 (N_13790,N_13439,N_13112);
nor U13791 (N_13791,N_13182,N_13072);
or U13792 (N_13792,N_13041,N_13153);
xnor U13793 (N_13793,N_13217,N_13452);
and U13794 (N_13794,N_13179,N_13384);
or U13795 (N_13795,N_13264,N_13130);
and U13796 (N_13796,N_13136,N_13190);
xnor U13797 (N_13797,N_13105,N_13281);
nor U13798 (N_13798,N_13008,N_13222);
nand U13799 (N_13799,N_13289,N_13198);
nand U13800 (N_13800,N_13474,N_13101);
xor U13801 (N_13801,N_13078,N_13249);
nand U13802 (N_13802,N_13162,N_13319);
and U13803 (N_13803,N_13253,N_13391);
xnor U13804 (N_13804,N_13117,N_13158);
nor U13805 (N_13805,N_13411,N_13206);
or U13806 (N_13806,N_13212,N_13354);
xnor U13807 (N_13807,N_13303,N_13042);
and U13808 (N_13808,N_13212,N_13264);
and U13809 (N_13809,N_13305,N_13443);
nor U13810 (N_13810,N_13235,N_13065);
and U13811 (N_13811,N_13265,N_13083);
xnor U13812 (N_13812,N_13133,N_13270);
and U13813 (N_13813,N_13137,N_13182);
or U13814 (N_13814,N_13409,N_13488);
nand U13815 (N_13815,N_13081,N_13017);
and U13816 (N_13816,N_13125,N_13244);
nor U13817 (N_13817,N_13361,N_13434);
xnor U13818 (N_13818,N_13257,N_13199);
nand U13819 (N_13819,N_13353,N_13101);
or U13820 (N_13820,N_13460,N_13219);
nand U13821 (N_13821,N_13057,N_13361);
nand U13822 (N_13822,N_13493,N_13323);
nor U13823 (N_13823,N_13080,N_13396);
and U13824 (N_13824,N_13241,N_13151);
xor U13825 (N_13825,N_13039,N_13413);
and U13826 (N_13826,N_13482,N_13421);
xor U13827 (N_13827,N_13352,N_13072);
nor U13828 (N_13828,N_13178,N_13040);
or U13829 (N_13829,N_13196,N_13312);
nand U13830 (N_13830,N_13074,N_13381);
nand U13831 (N_13831,N_13039,N_13480);
and U13832 (N_13832,N_13144,N_13417);
and U13833 (N_13833,N_13003,N_13468);
and U13834 (N_13834,N_13107,N_13290);
nor U13835 (N_13835,N_13492,N_13126);
nor U13836 (N_13836,N_13088,N_13453);
xor U13837 (N_13837,N_13472,N_13061);
xor U13838 (N_13838,N_13311,N_13232);
and U13839 (N_13839,N_13184,N_13213);
nand U13840 (N_13840,N_13278,N_13232);
or U13841 (N_13841,N_13068,N_13408);
nor U13842 (N_13842,N_13075,N_13110);
nand U13843 (N_13843,N_13165,N_13132);
xor U13844 (N_13844,N_13423,N_13139);
nand U13845 (N_13845,N_13161,N_13118);
nor U13846 (N_13846,N_13227,N_13198);
nor U13847 (N_13847,N_13313,N_13112);
nand U13848 (N_13848,N_13417,N_13162);
nand U13849 (N_13849,N_13466,N_13214);
and U13850 (N_13850,N_13490,N_13173);
nand U13851 (N_13851,N_13364,N_13009);
nand U13852 (N_13852,N_13375,N_13278);
xor U13853 (N_13853,N_13265,N_13458);
nor U13854 (N_13854,N_13345,N_13250);
nor U13855 (N_13855,N_13052,N_13442);
and U13856 (N_13856,N_13149,N_13027);
xor U13857 (N_13857,N_13430,N_13028);
nor U13858 (N_13858,N_13128,N_13156);
xnor U13859 (N_13859,N_13236,N_13496);
or U13860 (N_13860,N_13222,N_13167);
and U13861 (N_13861,N_13401,N_13404);
or U13862 (N_13862,N_13216,N_13271);
xor U13863 (N_13863,N_13315,N_13387);
or U13864 (N_13864,N_13299,N_13374);
or U13865 (N_13865,N_13393,N_13023);
or U13866 (N_13866,N_13479,N_13006);
xnor U13867 (N_13867,N_13343,N_13451);
and U13868 (N_13868,N_13216,N_13172);
nand U13869 (N_13869,N_13497,N_13121);
xnor U13870 (N_13870,N_13114,N_13366);
and U13871 (N_13871,N_13275,N_13157);
and U13872 (N_13872,N_13284,N_13311);
and U13873 (N_13873,N_13434,N_13263);
or U13874 (N_13874,N_13111,N_13099);
or U13875 (N_13875,N_13428,N_13174);
and U13876 (N_13876,N_13070,N_13059);
nand U13877 (N_13877,N_13359,N_13028);
nand U13878 (N_13878,N_13445,N_13130);
or U13879 (N_13879,N_13294,N_13131);
xnor U13880 (N_13880,N_13296,N_13095);
xor U13881 (N_13881,N_13004,N_13336);
or U13882 (N_13882,N_13127,N_13185);
or U13883 (N_13883,N_13468,N_13201);
nand U13884 (N_13884,N_13392,N_13234);
nor U13885 (N_13885,N_13012,N_13153);
xnor U13886 (N_13886,N_13043,N_13082);
nor U13887 (N_13887,N_13190,N_13355);
or U13888 (N_13888,N_13342,N_13440);
or U13889 (N_13889,N_13427,N_13488);
and U13890 (N_13890,N_13005,N_13344);
nor U13891 (N_13891,N_13350,N_13114);
or U13892 (N_13892,N_13446,N_13127);
and U13893 (N_13893,N_13370,N_13137);
nor U13894 (N_13894,N_13078,N_13348);
xor U13895 (N_13895,N_13354,N_13227);
xnor U13896 (N_13896,N_13243,N_13446);
or U13897 (N_13897,N_13430,N_13155);
or U13898 (N_13898,N_13363,N_13486);
and U13899 (N_13899,N_13381,N_13000);
or U13900 (N_13900,N_13304,N_13003);
nor U13901 (N_13901,N_13199,N_13288);
xnor U13902 (N_13902,N_13254,N_13477);
and U13903 (N_13903,N_13366,N_13454);
xnor U13904 (N_13904,N_13089,N_13213);
nor U13905 (N_13905,N_13168,N_13483);
or U13906 (N_13906,N_13344,N_13135);
nand U13907 (N_13907,N_13391,N_13442);
and U13908 (N_13908,N_13220,N_13414);
or U13909 (N_13909,N_13353,N_13111);
nand U13910 (N_13910,N_13436,N_13055);
nand U13911 (N_13911,N_13148,N_13217);
xnor U13912 (N_13912,N_13438,N_13205);
nor U13913 (N_13913,N_13356,N_13338);
and U13914 (N_13914,N_13091,N_13050);
or U13915 (N_13915,N_13253,N_13031);
and U13916 (N_13916,N_13012,N_13135);
xnor U13917 (N_13917,N_13455,N_13367);
nor U13918 (N_13918,N_13371,N_13328);
nor U13919 (N_13919,N_13069,N_13214);
or U13920 (N_13920,N_13478,N_13496);
xor U13921 (N_13921,N_13058,N_13216);
or U13922 (N_13922,N_13102,N_13239);
nor U13923 (N_13923,N_13151,N_13239);
nand U13924 (N_13924,N_13251,N_13104);
and U13925 (N_13925,N_13112,N_13437);
xor U13926 (N_13926,N_13361,N_13019);
xnor U13927 (N_13927,N_13082,N_13211);
nor U13928 (N_13928,N_13063,N_13377);
nor U13929 (N_13929,N_13066,N_13156);
or U13930 (N_13930,N_13069,N_13321);
and U13931 (N_13931,N_13059,N_13395);
nor U13932 (N_13932,N_13184,N_13180);
nand U13933 (N_13933,N_13222,N_13067);
nor U13934 (N_13934,N_13302,N_13259);
or U13935 (N_13935,N_13414,N_13325);
xor U13936 (N_13936,N_13167,N_13136);
xor U13937 (N_13937,N_13007,N_13249);
nor U13938 (N_13938,N_13443,N_13031);
nand U13939 (N_13939,N_13279,N_13340);
nor U13940 (N_13940,N_13247,N_13280);
nand U13941 (N_13941,N_13343,N_13230);
xnor U13942 (N_13942,N_13251,N_13449);
nand U13943 (N_13943,N_13336,N_13096);
nor U13944 (N_13944,N_13006,N_13374);
xor U13945 (N_13945,N_13462,N_13341);
and U13946 (N_13946,N_13117,N_13019);
nor U13947 (N_13947,N_13064,N_13382);
xnor U13948 (N_13948,N_13344,N_13126);
nand U13949 (N_13949,N_13264,N_13346);
or U13950 (N_13950,N_13359,N_13208);
nor U13951 (N_13951,N_13459,N_13054);
nand U13952 (N_13952,N_13455,N_13340);
and U13953 (N_13953,N_13478,N_13370);
xnor U13954 (N_13954,N_13465,N_13450);
nor U13955 (N_13955,N_13056,N_13469);
and U13956 (N_13956,N_13245,N_13221);
nor U13957 (N_13957,N_13179,N_13074);
nor U13958 (N_13958,N_13219,N_13390);
xnor U13959 (N_13959,N_13091,N_13077);
and U13960 (N_13960,N_13249,N_13064);
nand U13961 (N_13961,N_13475,N_13021);
or U13962 (N_13962,N_13039,N_13479);
and U13963 (N_13963,N_13497,N_13411);
xnor U13964 (N_13964,N_13154,N_13037);
or U13965 (N_13965,N_13421,N_13407);
and U13966 (N_13966,N_13186,N_13137);
nand U13967 (N_13967,N_13318,N_13499);
and U13968 (N_13968,N_13203,N_13317);
nor U13969 (N_13969,N_13403,N_13206);
or U13970 (N_13970,N_13267,N_13321);
xor U13971 (N_13971,N_13215,N_13107);
nand U13972 (N_13972,N_13374,N_13163);
and U13973 (N_13973,N_13414,N_13093);
nand U13974 (N_13974,N_13007,N_13434);
or U13975 (N_13975,N_13353,N_13321);
nor U13976 (N_13976,N_13076,N_13392);
and U13977 (N_13977,N_13055,N_13149);
and U13978 (N_13978,N_13047,N_13221);
and U13979 (N_13979,N_13291,N_13393);
and U13980 (N_13980,N_13080,N_13388);
xor U13981 (N_13981,N_13463,N_13497);
xor U13982 (N_13982,N_13182,N_13335);
and U13983 (N_13983,N_13138,N_13497);
or U13984 (N_13984,N_13240,N_13304);
xor U13985 (N_13985,N_13056,N_13090);
nand U13986 (N_13986,N_13417,N_13437);
nand U13987 (N_13987,N_13366,N_13265);
and U13988 (N_13988,N_13447,N_13257);
and U13989 (N_13989,N_13284,N_13306);
and U13990 (N_13990,N_13221,N_13373);
xor U13991 (N_13991,N_13180,N_13374);
xor U13992 (N_13992,N_13402,N_13216);
or U13993 (N_13993,N_13453,N_13379);
nor U13994 (N_13994,N_13111,N_13134);
nand U13995 (N_13995,N_13064,N_13143);
xnor U13996 (N_13996,N_13361,N_13436);
xor U13997 (N_13997,N_13353,N_13474);
or U13998 (N_13998,N_13436,N_13184);
and U13999 (N_13999,N_13156,N_13121);
nor U14000 (N_14000,N_13742,N_13670);
xor U14001 (N_14001,N_13513,N_13602);
xnor U14002 (N_14002,N_13960,N_13887);
nor U14003 (N_14003,N_13992,N_13973);
nor U14004 (N_14004,N_13942,N_13669);
nor U14005 (N_14005,N_13537,N_13959);
nand U14006 (N_14006,N_13784,N_13638);
nor U14007 (N_14007,N_13934,N_13896);
xnor U14008 (N_14008,N_13587,N_13706);
and U14009 (N_14009,N_13585,N_13768);
or U14010 (N_14010,N_13528,N_13953);
or U14011 (N_14011,N_13857,N_13508);
or U14012 (N_14012,N_13990,N_13552);
xnor U14013 (N_14013,N_13788,N_13958);
xnor U14014 (N_14014,N_13851,N_13580);
nor U14015 (N_14015,N_13627,N_13662);
nand U14016 (N_14016,N_13910,N_13625);
or U14017 (N_14017,N_13522,N_13805);
nand U14018 (N_14018,N_13916,N_13858);
and U14019 (N_14019,N_13545,N_13898);
nor U14020 (N_14020,N_13699,N_13765);
nor U14021 (N_14021,N_13658,N_13976);
nor U14022 (N_14022,N_13751,N_13752);
nor U14023 (N_14023,N_13901,N_13754);
xor U14024 (N_14024,N_13503,N_13512);
xnor U14025 (N_14025,N_13883,N_13578);
nand U14026 (N_14026,N_13935,N_13519);
or U14027 (N_14027,N_13741,N_13886);
nor U14028 (N_14028,N_13649,N_13715);
xnor U14029 (N_14029,N_13782,N_13590);
xnor U14030 (N_14030,N_13581,N_13971);
nand U14031 (N_14031,N_13837,N_13774);
nor U14032 (N_14032,N_13829,N_13530);
and U14033 (N_14033,N_13536,N_13769);
and U14034 (N_14034,N_13588,N_13997);
or U14035 (N_14035,N_13703,N_13605);
nand U14036 (N_14036,N_13659,N_13770);
and U14037 (N_14037,N_13761,N_13616);
and U14038 (N_14038,N_13702,N_13654);
and U14039 (N_14039,N_13760,N_13750);
nor U14040 (N_14040,N_13965,N_13977);
xor U14041 (N_14041,N_13560,N_13607);
xnor U14042 (N_14042,N_13758,N_13817);
xnor U14043 (N_14043,N_13866,N_13833);
and U14044 (N_14044,N_13665,N_13984);
nor U14045 (N_14045,N_13611,N_13591);
nor U14046 (N_14046,N_13505,N_13907);
and U14047 (N_14047,N_13961,N_13593);
nand U14048 (N_14048,N_13860,N_13839);
or U14049 (N_14049,N_13773,N_13720);
nor U14050 (N_14050,N_13957,N_13775);
or U14051 (N_14051,N_13853,N_13810);
nor U14052 (N_14052,N_13629,N_13917);
xor U14053 (N_14053,N_13951,N_13708);
and U14054 (N_14054,N_13739,N_13885);
or U14055 (N_14055,N_13852,N_13834);
and U14056 (N_14056,N_13707,N_13712);
or U14057 (N_14057,N_13546,N_13812);
or U14058 (N_14058,N_13640,N_13936);
nor U14059 (N_14059,N_13680,N_13811);
or U14060 (N_14060,N_13541,N_13677);
xnor U14061 (N_14061,N_13574,N_13798);
or U14062 (N_14062,N_13873,N_13912);
nand U14063 (N_14063,N_13986,N_13717);
nand U14064 (N_14064,N_13978,N_13766);
or U14065 (N_14065,N_13763,N_13818);
nor U14066 (N_14066,N_13617,N_13909);
nand U14067 (N_14067,N_13930,N_13737);
nand U14068 (N_14068,N_13686,N_13759);
or U14069 (N_14069,N_13989,N_13569);
xnor U14070 (N_14070,N_13937,N_13690);
or U14071 (N_14071,N_13727,N_13913);
nor U14072 (N_14072,N_13779,N_13848);
nor U14073 (N_14073,N_13663,N_13675);
or U14074 (N_14074,N_13781,N_13696);
nand U14075 (N_14075,N_13501,N_13988);
or U14076 (N_14076,N_13711,N_13946);
and U14077 (N_14077,N_13882,N_13791);
xor U14078 (N_14078,N_13684,N_13600);
and U14079 (N_14079,N_13732,N_13846);
and U14080 (N_14080,N_13550,N_13604);
nand U14081 (N_14081,N_13830,N_13943);
xor U14082 (N_14082,N_13985,N_13735);
xnor U14083 (N_14083,N_13914,N_13724);
nor U14084 (N_14084,N_13728,N_13840);
or U14085 (N_14085,N_13744,N_13504);
xor U14086 (N_14086,N_13999,N_13994);
and U14087 (N_14087,N_13924,N_13859);
xor U14088 (N_14088,N_13679,N_13911);
nand U14089 (N_14089,N_13667,N_13705);
and U14090 (N_14090,N_13874,N_13921);
or U14091 (N_14091,N_13844,N_13621);
and U14092 (N_14092,N_13870,N_13648);
xor U14093 (N_14093,N_13693,N_13804);
and U14094 (N_14094,N_13624,N_13687);
or U14095 (N_14095,N_13630,N_13568);
or U14096 (N_14096,N_13955,N_13738);
or U14097 (N_14097,N_13968,N_13966);
nor U14098 (N_14098,N_13842,N_13656);
and U14099 (N_14099,N_13736,N_13967);
or U14100 (N_14100,N_13856,N_13918);
xor U14101 (N_14101,N_13540,N_13704);
and U14102 (N_14102,N_13877,N_13601);
and U14103 (N_14103,N_13824,N_13963);
and U14104 (N_14104,N_13716,N_13645);
nand U14105 (N_14105,N_13867,N_13944);
nand U14106 (N_14106,N_13940,N_13511);
and U14107 (N_14107,N_13542,N_13729);
nand U14108 (N_14108,N_13962,N_13655);
nand U14109 (N_14109,N_13836,N_13772);
and U14110 (N_14110,N_13531,N_13553);
or U14111 (N_14111,N_13776,N_13905);
nand U14112 (N_14112,N_13664,N_13778);
or U14113 (N_14113,N_13923,N_13691);
nand U14114 (N_14114,N_13628,N_13660);
or U14115 (N_14115,N_13878,N_13785);
or U14116 (N_14116,N_13895,N_13740);
or U14117 (N_14117,N_13948,N_13900);
xor U14118 (N_14118,N_13719,N_13863);
nand U14119 (N_14119,N_13599,N_13606);
or U14120 (N_14120,N_13734,N_13821);
nor U14121 (N_14121,N_13796,N_13579);
or U14122 (N_14122,N_13730,N_13845);
or U14123 (N_14123,N_13523,N_13695);
and U14124 (N_14124,N_13748,N_13676);
nand U14125 (N_14125,N_13800,N_13619);
and U14126 (N_14126,N_13925,N_13570);
xnor U14127 (N_14127,N_13661,N_13783);
nand U14128 (N_14128,N_13577,N_13718);
nand U14129 (N_14129,N_13762,N_13673);
nor U14130 (N_14130,N_13562,N_13652);
nor U14131 (N_14131,N_13743,N_13982);
nand U14132 (N_14132,N_13635,N_13755);
or U14133 (N_14133,N_13710,N_13603);
nand U14134 (N_14134,N_13548,N_13543);
xor U14135 (N_14135,N_13820,N_13803);
nor U14136 (N_14136,N_13731,N_13701);
nand U14137 (N_14137,N_13615,N_13509);
nor U14138 (N_14138,N_13771,N_13709);
xor U14139 (N_14139,N_13933,N_13674);
xnor U14140 (N_14140,N_13612,N_13538);
xor U14141 (N_14141,N_13854,N_13979);
or U14142 (N_14142,N_13980,N_13631);
nor U14143 (N_14143,N_13726,N_13903);
and U14144 (N_14144,N_13610,N_13808);
nor U14145 (N_14145,N_13714,N_13534);
nand U14146 (N_14146,N_13525,N_13746);
xor U14147 (N_14147,N_13517,N_13794);
nand U14148 (N_14148,N_13609,N_13972);
nor U14149 (N_14149,N_13597,N_13700);
nor U14150 (N_14150,N_13747,N_13725);
xnor U14151 (N_14151,N_13713,N_13556);
nand U14152 (N_14152,N_13950,N_13850);
or U14153 (N_14153,N_13801,N_13897);
and U14154 (N_14154,N_13890,N_13894);
or U14155 (N_14155,N_13582,N_13780);
nor U14156 (N_14156,N_13634,N_13567);
or U14157 (N_14157,N_13643,N_13906);
and U14158 (N_14158,N_13757,N_13688);
nor U14159 (N_14159,N_13613,N_13952);
nand U14160 (N_14160,N_13849,N_13639);
nand U14161 (N_14161,N_13892,N_13641);
xnor U14162 (N_14162,N_13520,N_13539);
or U14163 (N_14163,N_13814,N_13880);
nor U14164 (N_14164,N_13875,N_13847);
nor U14165 (N_14165,N_13931,N_13576);
xor U14166 (N_14166,N_13516,N_13721);
nor U14167 (N_14167,N_13626,N_13749);
xor U14168 (N_14168,N_13502,N_13823);
xnor U14169 (N_14169,N_13793,N_13644);
nand U14170 (N_14170,N_13789,N_13983);
and U14171 (N_14171,N_13767,N_13908);
nand U14172 (N_14172,N_13826,N_13583);
or U14173 (N_14173,N_13993,N_13682);
xnor U14174 (N_14174,N_13533,N_13668);
or U14175 (N_14175,N_13904,N_13529);
nand U14176 (N_14176,N_13685,N_13919);
xor U14177 (N_14177,N_13799,N_13868);
nand U14178 (N_14178,N_13650,N_13756);
xor U14179 (N_14179,N_13975,N_13722);
and U14180 (N_14180,N_13608,N_13862);
and U14181 (N_14181,N_13532,N_13970);
or U14182 (N_14182,N_13618,N_13753);
nor U14183 (N_14183,N_13872,N_13506);
and U14184 (N_14184,N_13865,N_13807);
nand U14185 (N_14185,N_13592,N_13828);
or U14186 (N_14186,N_13786,N_13518);
and U14187 (N_14187,N_13555,N_13795);
or U14188 (N_14188,N_13777,N_13584);
xnor U14189 (N_14189,N_13838,N_13558);
nand U14190 (N_14190,N_13792,N_13598);
nor U14191 (N_14191,N_13816,N_13893);
or U14192 (N_14192,N_13764,N_13871);
and U14193 (N_14193,N_13802,N_13787);
nand U14194 (N_14194,N_13864,N_13733);
nand U14195 (N_14195,N_13987,N_13813);
nand U14196 (N_14196,N_13678,N_13595);
xnor U14197 (N_14197,N_13891,N_13938);
xor U14198 (N_14198,N_13510,N_13694);
nor U14199 (N_14199,N_13745,N_13651);
nand U14200 (N_14200,N_13527,N_13881);
nor U14201 (N_14201,N_13825,N_13790);
and U14202 (N_14202,N_13949,N_13827);
or U14203 (N_14203,N_13974,N_13797);
xor U14204 (N_14204,N_13551,N_13926);
or U14205 (N_14205,N_13697,N_13637);
nand U14206 (N_14206,N_13647,N_13941);
nor U14207 (N_14207,N_13969,N_13932);
or U14208 (N_14208,N_13559,N_13832);
or U14209 (N_14209,N_13594,N_13561);
or U14210 (N_14210,N_13572,N_13500);
xor U14211 (N_14211,N_13671,N_13689);
xor U14212 (N_14212,N_13922,N_13899);
or U14213 (N_14213,N_13831,N_13683);
nor U14214 (N_14214,N_13571,N_13956);
and U14215 (N_14215,N_13636,N_13589);
or U14216 (N_14216,N_13819,N_13642);
nand U14217 (N_14217,N_13575,N_13586);
nor U14218 (N_14218,N_13928,N_13563);
nor U14219 (N_14219,N_13547,N_13623);
xor U14220 (N_14220,N_13902,N_13939);
nor U14221 (N_14221,N_13981,N_13526);
and U14222 (N_14222,N_13672,N_13573);
and U14223 (N_14223,N_13549,N_13666);
nor U14224 (N_14224,N_13622,N_13879);
and U14225 (N_14225,N_13998,N_13927);
xnor U14226 (N_14226,N_13915,N_13947);
xnor U14227 (N_14227,N_13557,N_13535);
xnor U14228 (N_14228,N_13514,N_13809);
and U14229 (N_14229,N_13995,N_13632);
xnor U14230 (N_14230,N_13876,N_13657);
xnor U14231 (N_14231,N_13692,N_13815);
nand U14232 (N_14232,N_13554,N_13806);
or U14233 (N_14233,N_13954,N_13566);
xnor U14234 (N_14234,N_13544,N_13822);
or U14235 (N_14235,N_13681,N_13884);
nand U14236 (N_14236,N_13507,N_13920);
xor U14237 (N_14237,N_13596,N_13861);
nand U14238 (N_14238,N_13515,N_13565);
nand U14239 (N_14239,N_13633,N_13698);
and U14240 (N_14240,N_13964,N_13843);
nor U14241 (N_14241,N_13614,N_13888);
nand U14242 (N_14242,N_13889,N_13945);
or U14243 (N_14243,N_13524,N_13620);
nor U14244 (N_14244,N_13653,N_13929);
nor U14245 (N_14245,N_13855,N_13991);
nand U14246 (N_14246,N_13996,N_13869);
and U14247 (N_14247,N_13646,N_13841);
nand U14248 (N_14248,N_13564,N_13723);
nand U14249 (N_14249,N_13835,N_13521);
and U14250 (N_14250,N_13611,N_13757);
xor U14251 (N_14251,N_13888,N_13947);
or U14252 (N_14252,N_13821,N_13506);
nor U14253 (N_14253,N_13813,N_13776);
nand U14254 (N_14254,N_13512,N_13936);
or U14255 (N_14255,N_13693,N_13647);
or U14256 (N_14256,N_13702,N_13984);
or U14257 (N_14257,N_13954,N_13667);
or U14258 (N_14258,N_13750,N_13991);
nand U14259 (N_14259,N_13703,N_13993);
nor U14260 (N_14260,N_13530,N_13835);
xor U14261 (N_14261,N_13928,N_13518);
nor U14262 (N_14262,N_13825,N_13717);
or U14263 (N_14263,N_13741,N_13534);
nor U14264 (N_14264,N_13955,N_13858);
or U14265 (N_14265,N_13740,N_13970);
nand U14266 (N_14266,N_13868,N_13814);
or U14267 (N_14267,N_13735,N_13566);
nand U14268 (N_14268,N_13694,N_13896);
xor U14269 (N_14269,N_13532,N_13802);
xor U14270 (N_14270,N_13564,N_13611);
or U14271 (N_14271,N_13699,N_13638);
xor U14272 (N_14272,N_13885,N_13888);
and U14273 (N_14273,N_13944,N_13761);
and U14274 (N_14274,N_13998,N_13568);
nand U14275 (N_14275,N_13643,N_13876);
and U14276 (N_14276,N_13617,N_13953);
and U14277 (N_14277,N_13819,N_13840);
xnor U14278 (N_14278,N_13952,N_13923);
or U14279 (N_14279,N_13666,N_13880);
or U14280 (N_14280,N_13670,N_13576);
or U14281 (N_14281,N_13966,N_13846);
xnor U14282 (N_14282,N_13764,N_13812);
nor U14283 (N_14283,N_13528,N_13929);
nand U14284 (N_14284,N_13911,N_13792);
xnor U14285 (N_14285,N_13537,N_13778);
or U14286 (N_14286,N_13589,N_13751);
or U14287 (N_14287,N_13523,N_13947);
nand U14288 (N_14288,N_13942,N_13863);
nor U14289 (N_14289,N_13874,N_13650);
nand U14290 (N_14290,N_13521,N_13800);
and U14291 (N_14291,N_13898,N_13591);
or U14292 (N_14292,N_13942,N_13831);
and U14293 (N_14293,N_13684,N_13998);
nand U14294 (N_14294,N_13807,N_13673);
or U14295 (N_14295,N_13649,N_13592);
nand U14296 (N_14296,N_13700,N_13567);
and U14297 (N_14297,N_13861,N_13519);
and U14298 (N_14298,N_13927,N_13993);
nor U14299 (N_14299,N_13566,N_13870);
nor U14300 (N_14300,N_13512,N_13831);
and U14301 (N_14301,N_13818,N_13715);
nand U14302 (N_14302,N_13503,N_13550);
nand U14303 (N_14303,N_13752,N_13623);
and U14304 (N_14304,N_13845,N_13825);
xnor U14305 (N_14305,N_13764,N_13785);
xnor U14306 (N_14306,N_13509,N_13744);
xor U14307 (N_14307,N_13557,N_13590);
and U14308 (N_14308,N_13928,N_13533);
or U14309 (N_14309,N_13569,N_13579);
or U14310 (N_14310,N_13581,N_13662);
and U14311 (N_14311,N_13658,N_13507);
or U14312 (N_14312,N_13943,N_13761);
xnor U14313 (N_14313,N_13880,N_13961);
nor U14314 (N_14314,N_13742,N_13578);
or U14315 (N_14315,N_13888,N_13953);
nand U14316 (N_14316,N_13715,N_13902);
or U14317 (N_14317,N_13572,N_13651);
nor U14318 (N_14318,N_13532,N_13708);
nand U14319 (N_14319,N_13735,N_13776);
and U14320 (N_14320,N_13506,N_13707);
and U14321 (N_14321,N_13933,N_13661);
nand U14322 (N_14322,N_13504,N_13999);
xor U14323 (N_14323,N_13692,N_13653);
xor U14324 (N_14324,N_13647,N_13969);
xnor U14325 (N_14325,N_13766,N_13545);
xnor U14326 (N_14326,N_13968,N_13687);
nand U14327 (N_14327,N_13579,N_13827);
nand U14328 (N_14328,N_13536,N_13710);
nor U14329 (N_14329,N_13698,N_13547);
or U14330 (N_14330,N_13668,N_13662);
nor U14331 (N_14331,N_13649,N_13808);
or U14332 (N_14332,N_13930,N_13526);
and U14333 (N_14333,N_13507,N_13533);
and U14334 (N_14334,N_13658,N_13797);
nand U14335 (N_14335,N_13767,N_13744);
nor U14336 (N_14336,N_13908,N_13733);
nor U14337 (N_14337,N_13566,N_13952);
nand U14338 (N_14338,N_13947,N_13869);
xnor U14339 (N_14339,N_13811,N_13699);
or U14340 (N_14340,N_13537,N_13775);
nand U14341 (N_14341,N_13655,N_13651);
nor U14342 (N_14342,N_13594,N_13589);
xnor U14343 (N_14343,N_13854,N_13623);
or U14344 (N_14344,N_13802,N_13511);
and U14345 (N_14345,N_13653,N_13804);
or U14346 (N_14346,N_13674,N_13700);
or U14347 (N_14347,N_13938,N_13526);
nand U14348 (N_14348,N_13806,N_13762);
and U14349 (N_14349,N_13538,N_13521);
or U14350 (N_14350,N_13713,N_13961);
or U14351 (N_14351,N_13801,N_13966);
xor U14352 (N_14352,N_13854,N_13727);
nand U14353 (N_14353,N_13966,N_13512);
xnor U14354 (N_14354,N_13505,N_13810);
nand U14355 (N_14355,N_13654,N_13703);
nor U14356 (N_14356,N_13673,N_13759);
or U14357 (N_14357,N_13803,N_13893);
nor U14358 (N_14358,N_13878,N_13873);
nand U14359 (N_14359,N_13717,N_13936);
and U14360 (N_14360,N_13817,N_13833);
xor U14361 (N_14361,N_13603,N_13890);
or U14362 (N_14362,N_13740,N_13759);
xnor U14363 (N_14363,N_13574,N_13658);
xor U14364 (N_14364,N_13646,N_13979);
xnor U14365 (N_14365,N_13541,N_13619);
nor U14366 (N_14366,N_13546,N_13526);
nand U14367 (N_14367,N_13866,N_13536);
nand U14368 (N_14368,N_13901,N_13899);
nand U14369 (N_14369,N_13564,N_13785);
nand U14370 (N_14370,N_13991,N_13788);
nor U14371 (N_14371,N_13763,N_13501);
xor U14372 (N_14372,N_13791,N_13768);
xnor U14373 (N_14373,N_13824,N_13603);
and U14374 (N_14374,N_13598,N_13995);
and U14375 (N_14375,N_13621,N_13865);
xnor U14376 (N_14376,N_13982,N_13749);
or U14377 (N_14377,N_13592,N_13692);
nand U14378 (N_14378,N_13976,N_13524);
nor U14379 (N_14379,N_13861,N_13642);
or U14380 (N_14380,N_13773,N_13694);
xor U14381 (N_14381,N_13618,N_13626);
nor U14382 (N_14382,N_13873,N_13984);
nor U14383 (N_14383,N_13816,N_13923);
nand U14384 (N_14384,N_13843,N_13977);
and U14385 (N_14385,N_13515,N_13591);
or U14386 (N_14386,N_13896,N_13595);
nand U14387 (N_14387,N_13807,N_13827);
and U14388 (N_14388,N_13633,N_13737);
xnor U14389 (N_14389,N_13958,N_13986);
or U14390 (N_14390,N_13731,N_13904);
and U14391 (N_14391,N_13948,N_13504);
and U14392 (N_14392,N_13862,N_13683);
or U14393 (N_14393,N_13698,N_13996);
nor U14394 (N_14394,N_13643,N_13728);
and U14395 (N_14395,N_13765,N_13871);
xnor U14396 (N_14396,N_13969,N_13771);
and U14397 (N_14397,N_13903,N_13781);
nand U14398 (N_14398,N_13683,N_13645);
nand U14399 (N_14399,N_13716,N_13735);
xnor U14400 (N_14400,N_13735,N_13523);
xnor U14401 (N_14401,N_13840,N_13805);
or U14402 (N_14402,N_13590,N_13833);
and U14403 (N_14403,N_13613,N_13738);
nor U14404 (N_14404,N_13683,N_13585);
xnor U14405 (N_14405,N_13943,N_13551);
nor U14406 (N_14406,N_13769,N_13856);
nand U14407 (N_14407,N_13764,N_13575);
or U14408 (N_14408,N_13929,N_13734);
nand U14409 (N_14409,N_13983,N_13719);
nand U14410 (N_14410,N_13750,N_13500);
and U14411 (N_14411,N_13843,N_13989);
and U14412 (N_14412,N_13675,N_13722);
nor U14413 (N_14413,N_13935,N_13598);
nor U14414 (N_14414,N_13890,N_13994);
and U14415 (N_14415,N_13743,N_13591);
nand U14416 (N_14416,N_13632,N_13732);
nand U14417 (N_14417,N_13670,N_13528);
xnor U14418 (N_14418,N_13930,N_13902);
xnor U14419 (N_14419,N_13734,N_13535);
and U14420 (N_14420,N_13786,N_13687);
nand U14421 (N_14421,N_13568,N_13840);
nor U14422 (N_14422,N_13788,N_13710);
nand U14423 (N_14423,N_13602,N_13711);
xor U14424 (N_14424,N_13974,N_13681);
xor U14425 (N_14425,N_13530,N_13565);
nand U14426 (N_14426,N_13609,N_13760);
and U14427 (N_14427,N_13965,N_13846);
nor U14428 (N_14428,N_13769,N_13853);
and U14429 (N_14429,N_13727,N_13608);
nand U14430 (N_14430,N_13740,N_13774);
nand U14431 (N_14431,N_13607,N_13697);
or U14432 (N_14432,N_13645,N_13671);
nand U14433 (N_14433,N_13666,N_13581);
and U14434 (N_14434,N_13748,N_13792);
xor U14435 (N_14435,N_13893,N_13567);
nand U14436 (N_14436,N_13713,N_13862);
nor U14437 (N_14437,N_13949,N_13785);
xnor U14438 (N_14438,N_13591,N_13783);
nor U14439 (N_14439,N_13880,N_13527);
xnor U14440 (N_14440,N_13711,N_13781);
nand U14441 (N_14441,N_13653,N_13847);
nand U14442 (N_14442,N_13790,N_13902);
or U14443 (N_14443,N_13552,N_13705);
nand U14444 (N_14444,N_13788,N_13817);
nand U14445 (N_14445,N_13919,N_13615);
nor U14446 (N_14446,N_13821,N_13980);
xor U14447 (N_14447,N_13808,N_13752);
nand U14448 (N_14448,N_13990,N_13962);
and U14449 (N_14449,N_13624,N_13571);
xnor U14450 (N_14450,N_13963,N_13703);
nor U14451 (N_14451,N_13729,N_13760);
and U14452 (N_14452,N_13938,N_13584);
xnor U14453 (N_14453,N_13835,N_13503);
and U14454 (N_14454,N_13671,N_13639);
or U14455 (N_14455,N_13972,N_13665);
nand U14456 (N_14456,N_13555,N_13709);
xnor U14457 (N_14457,N_13875,N_13804);
xnor U14458 (N_14458,N_13685,N_13567);
nor U14459 (N_14459,N_13580,N_13704);
nand U14460 (N_14460,N_13664,N_13516);
nand U14461 (N_14461,N_13548,N_13811);
xor U14462 (N_14462,N_13896,N_13815);
nand U14463 (N_14463,N_13538,N_13907);
or U14464 (N_14464,N_13631,N_13807);
nor U14465 (N_14465,N_13992,N_13570);
nand U14466 (N_14466,N_13899,N_13537);
xor U14467 (N_14467,N_13595,N_13958);
or U14468 (N_14468,N_13516,N_13520);
nand U14469 (N_14469,N_13788,N_13835);
or U14470 (N_14470,N_13842,N_13765);
nand U14471 (N_14471,N_13871,N_13710);
or U14472 (N_14472,N_13925,N_13736);
nand U14473 (N_14473,N_13983,N_13909);
nand U14474 (N_14474,N_13528,N_13507);
or U14475 (N_14475,N_13868,N_13524);
and U14476 (N_14476,N_13501,N_13692);
nand U14477 (N_14477,N_13640,N_13808);
nor U14478 (N_14478,N_13658,N_13986);
xor U14479 (N_14479,N_13938,N_13836);
or U14480 (N_14480,N_13968,N_13951);
and U14481 (N_14481,N_13591,N_13734);
xnor U14482 (N_14482,N_13844,N_13523);
xor U14483 (N_14483,N_13720,N_13837);
xor U14484 (N_14484,N_13626,N_13789);
nor U14485 (N_14485,N_13886,N_13622);
nor U14486 (N_14486,N_13831,N_13523);
xnor U14487 (N_14487,N_13828,N_13990);
xnor U14488 (N_14488,N_13506,N_13552);
or U14489 (N_14489,N_13748,N_13914);
xnor U14490 (N_14490,N_13958,N_13577);
nand U14491 (N_14491,N_13958,N_13625);
and U14492 (N_14492,N_13963,N_13666);
and U14493 (N_14493,N_13555,N_13968);
nand U14494 (N_14494,N_13901,N_13922);
or U14495 (N_14495,N_13669,N_13897);
or U14496 (N_14496,N_13657,N_13555);
nor U14497 (N_14497,N_13795,N_13569);
nand U14498 (N_14498,N_13889,N_13664);
or U14499 (N_14499,N_13635,N_13761);
nand U14500 (N_14500,N_14341,N_14472);
nand U14501 (N_14501,N_14252,N_14033);
xor U14502 (N_14502,N_14339,N_14350);
nor U14503 (N_14503,N_14156,N_14176);
and U14504 (N_14504,N_14145,N_14439);
nor U14505 (N_14505,N_14440,N_14105);
and U14506 (N_14506,N_14427,N_14488);
and U14507 (N_14507,N_14046,N_14400);
or U14508 (N_14508,N_14358,N_14122);
and U14509 (N_14509,N_14493,N_14024);
and U14510 (N_14510,N_14376,N_14343);
and U14511 (N_14511,N_14482,N_14269);
nor U14512 (N_14512,N_14014,N_14178);
xnor U14513 (N_14513,N_14090,N_14115);
or U14514 (N_14514,N_14282,N_14037);
nand U14515 (N_14515,N_14352,N_14408);
and U14516 (N_14516,N_14007,N_14331);
nor U14517 (N_14517,N_14457,N_14095);
xnor U14518 (N_14518,N_14478,N_14034);
nand U14519 (N_14519,N_14491,N_14107);
nand U14520 (N_14520,N_14398,N_14255);
or U14521 (N_14521,N_14464,N_14008);
or U14522 (N_14522,N_14078,N_14066);
xnor U14523 (N_14523,N_14285,N_14371);
or U14524 (N_14524,N_14299,N_14264);
or U14525 (N_14525,N_14366,N_14053);
xnor U14526 (N_14526,N_14195,N_14075);
or U14527 (N_14527,N_14238,N_14311);
and U14528 (N_14528,N_14042,N_14498);
xnor U14529 (N_14529,N_14169,N_14184);
and U14530 (N_14530,N_14128,N_14197);
nor U14531 (N_14531,N_14302,N_14487);
and U14532 (N_14532,N_14304,N_14324);
or U14533 (N_14533,N_14079,N_14104);
or U14534 (N_14534,N_14381,N_14340);
xnor U14535 (N_14535,N_14388,N_14308);
xnor U14536 (N_14536,N_14136,N_14306);
nor U14537 (N_14537,N_14097,N_14330);
xnor U14538 (N_14538,N_14142,N_14461);
and U14539 (N_14539,N_14447,N_14060);
or U14540 (N_14540,N_14173,N_14077);
xnor U14541 (N_14541,N_14384,N_14023);
or U14542 (N_14542,N_14061,N_14259);
xor U14543 (N_14543,N_14470,N_14154);
and U14544 (N_14544,N_14120,N_14429);
or U14545 (N_14545,N_14260,N_14207);
and U14546 (N_14546,N_14146,N_14329);
or U14547 (N_14547,N_14283,N_14138);
xnor U14548 (N_14548,N_14214,N_14017);
nor U14549 (N_14549,N_14396,N_14319);
or U14550 (N_14550,N_14127,N_14148);
nand U14551 (N_14551,N_14425,N_14293);
nor U14552 (N_14552,N_14256,N_14266);
nor U14553 (N_14553,N_14399,N_14222);
xnor U14554 (N_14554,N_14415,N_14432);
and U14555 (N_14555,N_14094,N_14475);
and U14556 (N_14556,N_14118,N_14333);
or U14557 (N_14557,N_14010,N_14224);
nand U14558 (N_14558,N_14239,N_14430);
xor U14559 (N_14559,N_14141,N_14393);
and U14560 (N_14560,N_14402,N_14389);
nor U14561 (N_14561,N_14454,N_14431);
and U14562 (N_14562,N_14158,N_14392);
nand U14563 (N_14563,N_14211,N_14407);
xnor U14564 (N_14564,N_14323,N_14290);
nor U14565 (N_14565,N_14316,N_14117);
nor U14566 (N_14566,N_14191,N_14228);
nor U14567 (N_14567,N_14110,N_14446);
nand U14568 (N_14568,N_14433,N_14153);
and U14569 (N_14569,N_14313,N_14423);
and U14570 (N_14570,N_14111,N_14139);
nand U14571 (N_14571,N_14058,N_14021);
nand U14572 (N_14572,N_14353,N_14373);
nor U14573 (N_14573,N_14474,N_14100);
and U14574 (N_14574,N_14159,N_14043);
nor U14575 (N_14575,N_14426,N_14337);
nand U14576 (N_14576,N_14403,N_14436);
or U14577 (N_14577,N_14057,N_14377);
xnor U14578 (N_14578,N_14074,N_14121);
xor U14579 (N_14579,N_14204,N_14418);
and U14580 (N_14580,N_14096,N_14404);
nor U14581 (N_14581,N_14036,N_14480);
xnor U14582 (N_14582,N_14244,N_14296);
or U14583 (N_14583,N_14278,N_14087);
xnor U14584 (N_14584,N_14364,N_14417);
nor U14585 (N_14585,N_14182,N_14124);
xor U14586 (N_14586,N_14062,N_14137);
nand U14587 (N_14587,N_14442,N_14167);
or U14588 (N_14588,N_14450,N_14466);
or U14589 (N_14589,N_14005,N_14428);
nor U14590 (N_14590,N_14391,N_14355);
nor U14591 (N_14591,N_14463,N_14233);
nand U14592 (N_14592,N_14254,N_14183);
xor U14593 (N_14593,N_14044,N_14499);
nand U14594 (N_14594,N_14106,N_14280);
and U14595 (N_14595,N_14144,N_14274);
xor U14596 (N_14596,N_14190,N_14130);
and U14597 (N_14597,N_14284,N_14245);
nand U14598 (N_14598,N_14114,N_14237);
or U14599 (N_14599,N_14199,N_14370);
xor U14600 (N_14600,N_14483,N_14192);
or U14601 (N_14601,N_14451,N_14019);
xnor U14602 (N_14602,N_14015,N_14441);
nand U14603 (N_14603,N_14273,N_14312);
or U14604 (N_14604,N_14288,N_14026);
nand U14605 (N_14605,N_14289,N_14368);
or U14606 (N_14606,N_14149,N_14452);
nor U14607 (N_14607,N_14286,N_14372);
nand U14608 (N_14608,N_14342,N_14098);
nor U14609 (N_14609,N_14049,N_14011);
nand U14610 (N_14610,N_14242,N_14134);
xnor U14611 (N_14611,N_14301,N_14367);
or U14612 (N_14612,N_14481,N_14484);
and U14613 (N_14613,N_14344,N_14420);
nor U14614 (N_14614,N_14186,N_14453);
or U14615 (N_14615,N_14068,N_14133);
or U14616 (N_14616,N_14116,N_14486);
xnor U14617 (N_14617,N_14150,N_14129);
or U14618 (N_14618,N_14421,N_14218);
xnor U14619 (N_14619,N_14022,N_14047);
and U14620 (N_14620,N_14201,N_14152);
or U14621 (N_14621,N_14492,N_14262);
nand U14622 (N_14622,N_14385,N_14101);
nor U14623 (N_14623,N_14071,N_14243);
nand U14624 (N_14624,N_14067,N_14202);
or U14625 (N_14625,N_14084,N_14170);
or U14626 (N_14626,N_14161,N_14485);
and U14627 (N_14627,N_14336,N_14162);
nor U14628 (N_14628,N_14276,N_14261);
and U14629 (N_14629,N_14303,N_14348);
or U14630 (N_14630,N_14210,N_14444);
nand U14631 (N_14631,N_14497,N_14268);
xor U14632 (N_14632,N_14048,N_14291);
or U14633 (N_14633,N_14328,N_14179);
or U14634 (N_14634,N_14458,N_14012);
nor U14635 (N_14635,N_14018,N_14369);
nand U14636 (N_14636,N_14305,N_14409);
xnor U14637 (N_14637,N_14471,N_14424);
nand U14638 (N_14638,N_14379,N_14467);
or U14639 (N_14639,N_14132,N_14295);
and U14640 (N_14640,N_14172,N_14346);
nor U14641 (N_14641,N_14332,N_14270);
nand U14642 (N_14642,N_14247,N_14265);
or U14643 (N_14643,N_14263,N_14397);
nor U14644 (N_14644,N_14249,N_14227);
nand U14645 (N_14645,N_14160,N_14135);
nand U14646 (N_14646,N_14318,N_14089);
or U14647 (N_14647,N_14401,N_14166);
nand U14648 (N_14648,N_14193,N_14052);
nand U14649 (N_14649,N_14006,N_14416);
or U14650 (N_14650,N_14310,N_14411);
xor U14651 (N_14651,N_14203,N_14275);
and U14652 (N_14652,N_14382,N_14035);
xor U14653 (N_14653,N_14443,N_14272);
or U14654 (N_14654,N_14347,N_14473);
nand U14655 (N_14655,N_14386,N_14032);
nor U14656 (N_14656,N_14085,N_14212);
or U14657 (N_14657,N_14220,N_14147);
nor U14658 (N_14658,N_14025,N_14004);
or U14659 (N_14659,N_14279,N_14248);
nor U14660 (N_14660,N_14020,N_14000);
xnor U14661 (N_14661,N_14083,N_14315);
xor U14662 (N_14662,N_14476,N_14394);
nor U14663 (N_14663,N_14174,N_14165);
xnor U14664 (N_14664,N_14200,N_14143);
or U14665 (N_14665,N_14216,N_14390);
and U14666 (N_14666,N_14039,N_14215);
nand U14667 (N_14667,N_14002,N_14406);
nor U14668 (N_14668,N_14297,N_14236);
or U14669 (N_14669,N_14040,N_14405);
nand U14670 (N_14670,N_14065,N_14414);
nand U14671 (N_14671,N_14119,N_14157);
xor U14672 (N_14672,N_14327,N_14365);
nand U14673 (N_14673,N_14086,N_14459);
nor U14674 (N_14674,N_14300,N_14437);
and U14675 (N_14675,N_14335,N_14155);
nor U14676 (N_14676,N_14448,N_14378);
nand U14677 (N_14677,N_14325,N_14320);
nor U14678 (N_14678,N_14038,N_14309);
nand U14679 (N_14679,N_14091,N_14226);
or U14680 (N_14680,N_14395,N_14027);
or U14681 (N_14681,N_14455,N_14281);
and U14682 (N_14682,N_14064,N_14462);
and U14683 (N_14683,N_14349,N_14240);
nand U14684 (N_14684,N_14208,N_14001);
xor U14685 (N_14685,N_14168,N_14334);
xnor U14686 (N_14686,N_14338,N_14198);
xor U14687 (N_14687,N_14465,N_14003);
and U14688 (N_14688,N_14232,N_14050);
xor U14689 (N_14689,N_14082,N_14359);
or U14690 (N_14690,N_14449,N_14189);
nor U14691 (N_14691,N_14073,N_14460);
nor U14692 (N_14692,N_14292,N_14185);
and U14693 (N_14693,N_14051,N_14194);
and U14694 (N_14694,N_14271,N_14181);
nand U14695 (N_14695,N_14250,N_14307);
and U14696 (N_14696,N_14231,N_14469);
or U14697 (N_14697,N_14219,N_14028);
nand U14698 (N_14698,N_14380,N_14317);
and U14699 (N_14699,N_14112,N_14054);
nand U14700 (N_14700,N_14030,N_14434);
or U14701 (N_14701,N_14056,N_14321);
xor U14702 (N_14702,N_14477,N_14093);
and U14703 (N_14703,N_14251,N_14069);
or U14704 (N_14704,N_14375,N_14221);
nand U14705 (N_14705,N_14357,N_14209);
nor U14706 (N_14706,N_14205,N_14387);
and U14707 (N_14707,N_14246,N_14383);
nor U14708 (N_14708,N_14125,N_14140);
nor U14709 (N_14709,N_14081,N_14171);
and U14710 (N_14710,N_14496,N_14229);
xor U14711 (N_14711,N_14351,N_14412);
or U14712 (N_14712,N_14102,N_14187);
xnor U14713 (N_14713,N_14468,N_14277);
nor U14714 (N_14714,N_14479,N_14490);
or U14715 (N_14715,N_14445,N_14230);
nor U14716 (N_14716,N_14410,N_14287);
or U14717 (N_14717,N_14126,N_14435);
nand U14718 (N_14718,N_14206,N_14267);
xnor U14719 (N_14719,N_14456,N_14180);
xnor U14720 (N_14720,N_14163,N_14055);
nor U14721 (N_14721,N_14298,N_14361);
nand U14722 (N_14722,N_14109,N_14177);
or U14723 (N_14723,N_14294,N_14131);
and U14724 (N_14724,N_14164,N_14151);
nor U14725 (N_14725,N_14072,N_14494);
or U14726 (N_14726,N_14059,N_14345);
or U14727 (N_14727,N_14175,N_14360);
nor U14728 (N_14728,N_14253,N_14213);
nand U14729 (N_14729,N_14217,N_14223);
or U14730 (N_14730,N_14354,N_14031);
nand U14731 (N_14731,N_14103,N_14092);
nand U14732 (N_14732,N_14489,N_14009);
xnor U14733 (N_14733,N_14495,N_14123);
xnor U14734 (N_14734,N_14419,N_14322);
xnor U14735 (N_14735,N_14045,N_14029);
xnor U14736 (N_14736,N_14076,N_14356);
nand U14737 (N_14737,N_14099,N_14258);
xnor U14738 (N_14738,N_14196,N_14013);
nand U14739 (N_14739,N_14063,N_14235);
or U14740 (N_14740,N_14241,N_14016);
nand U14741 (N_14741,N_14374,N_14108);
and U14742 (N_14742,N_14188,N_14088);
or U14743 (N_14743,N_14080,N_14113);
and U14744 (N_14744,N_14070,N_14326);
and U14745 (N_14745,N_14363,N_14225);
or U14746 (N_14746,N_14234,N_14362);
and U14747 (N_14747,N_14413,N_14314);
nor U14748 (N_14748,N_14041,N_14422);
nand U14749 (N_14749,N_14257,N_14438);
nor U14750 (N_14750,N_14335,N_14059);
nand U14751 (N_14751,N_14298,N_14410);
nand U14752 (N_14752,N_14316,N_14317);
or U14753 (N_14753,N_14059,N_14203);
or U14754 (N_14754,N_14154,N_14391);
or U14755 (N_14755,N_14254,N_14441);
or U14756 (N_14756,N_14165,N_14333);
nand U14757 (N_14757,N_14317,N_14131);
nand U14758 (N_14758,N_14061,N_14400);
or U14759 (N_14759,N_14216,N_14491);
xnor U14760 (N_14760,N_14211,N_14493);
nand U14761 (N_14761,N_14106,N_14036);
xnor U14762 (N_14762,N_14489,N_14087);
or U14763 (N_14763,N_14050,N_14151);
nand U14764 (N_14764,N_14009,N_14377);
nand U14765 (N_14765,N_14201,N_14310);
nand U14766 (N_14766,N_14412,N_14421);
or U14767 (N_14767,N_14133,N_14348);
nand U14768 (N_14768,N_14061,N_14114);
nor U14769 (N_14769,N_14375,N_14396);
or U14770 (N_14770,N_14137,N_14494);
or U14771 (N_14771,N_14333,N_14457);
xnor U14772 (N_14772,N_14342,N_14043);
nor U14773 (N_14773,N_14465,N_14290);
and U14774 (N_14774,N_14393,N_14444);
and U14775 (N_14775,N_14386,N_14394);
xor U14776 (N_14776,N_14130,N_14302);
nor U14777 (N_14777,N_14239,N_14250);
and U14778 (N_14778,N_14489,N_14115);
nor U14779 (N_14779,N_14475,N_14048);
or U14780 (N_14780,N_14335,N_14290);
and U14781 (N_14781,N_14136,N_14053);
xor U14782 (N_14782,N_14433,N_14151);
and U14783 (N_14783,N_14269,N_14337);
or U14784 (N_14784,N_14453,N_14175);
or U14785 (N_14785,N_14353,N_14179);
nand U14786 (N_14786,N_14421,N_14450);
nand U14787 (N_14787,N_14081,N_14176);
nor U14788 (N_14788,N_14076,N_14365);
nor U14789 (N_14789,N_14248,N_14072);
and U14790 (N_14790,N_14039,N_14353);
and U14791 (N_14791,N_14234,N_14014);
or U14792 (N_14792,N_14121,N_14216);
and U14793 (N_14793,N_14237,N_14165);
or U14794 (N_14794,N_14125,N_14330);
nor U14795 (N_14795,N_14099,N_14059);
nor U14796 (N_14796,N_14362,N_14447);
nor U14797 (N_14797,N_14174,N_14436);
and U14798 (N_14798,N_14220,N_14213);
nor U14799 (N_14799,N_14074,N_14452);
nor U14800 (N_14800,N_14327,N_14128);
nand U14801 (N_14801,N_14400,N_14251);
xor U14802 (N_14802,N_14106,N_14040);
nor U14803 (N_14803,N_14419,N_14017);
nor U14804 (N_14804,N_14055,N_14135);
nor U14805 (N_14805,N_14109,N_14324);
nand U14806 (N_14806,N_14402,N_14317);
nand U14807 (N_14807,N_14145,N_14429);
xnor U14808 (N_14808,N_14004,N_14479);
nand U14809 (N_14809,N_14454,N_14219);
nor U14810 (N_14810,N_14346,N_14395);
and U14811 (N_14811,N_14056,N_14211);
nand U14812 (N_14812,N_14244,N_14203);
and U14813 (N_14813,N_14285,N_14010);
and U14814 (N_14814,N_14126,N_14219);
nand U14815 (N_14815,N_14189,N_14459);
xor U14816 (N_14816,N_14428,N_14293);
xor U14817 (N_14817,N_14034,N_14089);
and U14818 (N_14818,N_14447,N_14282);
nand U14819 (N_14819,N_14466,N_14496);
xor U14820 (N_14820,N_14200,N_14449);
and U14821 (N_14821,N_14147,N_14403);
xor U14822 (N_14822,N_14437,N_14242);
nand U14823 (N_14823,N_14390,N_14130);
nor U14824 (N_14824,N_14392,N_14310);
nor U14825 (N_14825,N_14187,N_14132);
nor U14826 (N_14826,N_14227,N_14361);
and U14827 (N_14827,N_14306,N_14156);
or U14828 (N_14828,N_14252,N_14008);
or U14829 (N_14829,N_14491,N_14413);
or U14830 (N_14830,N_14152,N_14393);
nand U14831 (N_14831,N_14048,N_14295);
and U14832 (N_14832,N_14451,N_14459);
nand U14833 (N_14833,N_14250,N_14066);
nor U14834 (N_14834,N_14240,N_14286);
and U14835 (N_14835,N_14043,N_14194);
and U14836 (N_14836,N_14231,N_14325);
nor U14837 (N_14837,N_14360,N_14398);
nor U14838 (N_14838,N_14228,N_14083);
nand U14839 (N_14839,N_14337,N_14315);
nor U14840 (N_14840,N_14300,N_14259);
xor U14841 (N_14841,N_14432,N_14194);
and U14842 (N_14842,N_14122,N_14364);
xnor U14843 (N_14843,N_14050,N_14057);
nand U14844 (N_14844,N_14249,N_14008);
or U14845 (N_14845,N_14147,N_14170);
nand U14846 (N_14846,N_14027,N_14463);
xnor U14847 (N_14847,N_14304,N_14080);
nand U14848 (N_14848,N_14127,N_14246);
or U14849 (N_14849,N_14147,N_14156);
or U14850 (N_14850,N_14196,N_14447);
or U14851 (N_14851,N_14206,N_14278);
or U14852 (N_14852,N_14388,N_14450);
xnor U14853 (N_14853,N_14041,N_14285);
and U14854 (N_14854,N_14436,N_14467);
nand U14855 (N_14855,N_14406,N_14036);
nor U14856 (N_14856,N_14440,N_14131);
and U14857 (N_14857,N_14038,N_14346);
and U14858 (N_14858,N_14061,N_14292);
nand U14859 (N_14859,N_14385,N_14282);
xnor U14860 (N_14860,N_14047,N_14313);
nand U14861 (N_14861,N_14412,N_14214);
nor U14862 (N_14862,N_14208,N_14260);
and U14863 (N_14863,N_14141,N_14135);
or U14864 (N_14864,N_14243,N_14073);
nor U14865 (N_14865,N_14079,N_14210);
nand U14866 (N_14866,N_14331,N_14230);
xnor U14867 (N_14867,N_14050,N_14177);
nand U14868 (N_14868,N_14053,N_14025);
nand U14869 (N_14869,N_14021,N_14086);
nand U14870 (N_14870,N_14479,N_14108);
xor U14871 (N_14871,N_14159,N_14382);
nor U14872 (N_14872,N_14432,N_14109);
or U14873 (N_14873,N_14340,N_14058);
nand U14874 (N_14874,N_14192,N_14384);
and U14875 (N_14875,N_14449,N_14184);
nand U14876 (N_14876,N_14373,N_14460);
and U14877 (N_14877,N_14012,N_14288);
nand U14878 (N_14878,N_14344,N_14261);
nor U14879 (N_14879,N_14121,N_14405);
nand U14880 (N_14880,N_14107,N_14385);
and U14881 (N_14881,N_14209,N_14014);
or U14882 (N_14882,N_14067,N_14161);
xnor U14883 (N_14883,N_14215,N_14368);
nand U14884 (N_14884,N_14300,N_14475);
nand U14885 (N_14885,N_14358,N_14455);
or U14886 (N_14886,N_14297,N_14483);
xor U14887 (N_14887,N_14306,N_14265);
xnor U14888 (N_14888,N_14261,N_14145);
xor U14889 (N_14889,N_14492,N_14460);
and U14890 (N_14890,N_14281,N_14216);
xnor U14891 (N_14891,N_14375,N_14476);
and U14892 (N_14892,N_14025,N_14060);
and U14893 (N_14893,N_14404,N_14088);
or U14894 (N_14894,N_14384,N_14401);
nand U14895 (N_14895,N_14468,N_14404);
or U14896 (N_14896,N_14470,N_14108);
nand U14897 (N_14897,N_14490,N_14218);
nand U14898 (N_14898,N_14347,N_14253);
or U14899 (N_14899,N_14474,N_14062);
and U14900 (N_14900,N_14222,N_14367);
xor U14901 (N_14901,N_14048,N_14415);
or U14902 (N_14902,N_14066,N_14135);
or U14903 (N_14903,N_14196,N_14060);
or U14904 (N_14904,N_14110,N_14109);
and U14905 (N_14905,N_14452,N_14106);
nor U14906 (N_14906,N_14464,N_14014);
nand U14907 (N_14907,N_14145,N_14050);
nand U14908 (N_14908,N_14300,N_14026);
xnor U14909 (N_14909,N_14445,N_14103);
nand U14910 (N_14910,N_14396,N_14019);
nand U14911 (N_14911,N_14343,N_14036);
xor U14912 (N_14912,N_14360,N_14041);
and U14913 (N_14913,N_14321,N_14061);
nand U14914 (N_14914,N_14393,N_14385);
nor U14915 (N_14915,N_14249,N_14340);
xor U14916 (N_14916,N_14363,N_14102);
or U14917 (N_14917,N_14387,N_14326);
nand U14918 (N_14918,N_14114,N_14247);
xor U14919 (N_14919,N_14438,N_14266);
xor U14920 (N_14920,N_14243,N_14330);
nor U14921 (N_14921,N_14037,N_14006);
nand U14922 (N_14922,N_14042,N_14054);
xnor U14923 (N_14923,N_14178,N_14496);
nand U14924 (N_14924,N_14114,N_14262);
xor U14925 (N_14925,N_14266,N_14237);
nand U14926 (N_14926,N_14311,N_14169);
nor U14927 (N_14927,N_14212,N_14458);
nand U14928 (N_14928,N_14332,N_14044);
nand U14929 (N_14929,N_14386,N_14332);
or U14930 (N_14930,N_14024,N_14375);
nand U14931 (N_14931,N_14447,N_14179);
nor U14932 (N_14932,N_14451,N_14315);
and U14933 (N_14933,N_14389,N_14275);
or U14934 (N_14934,N_14416,N_14015);
or U14935 (N_14935,N_14489,N_14088);
xor U14936 (N_14936,N_14153,N_14207);
nand U14937 (N_14937,N_14073,N_14215);
and U14938 (N_14938,N_14184,N_14358);
or U14939 (N_14939,N_14208,N_14099);
xnor U14940 (N_14940,N_14297,N_14199);
or U14941 (N_14941,N_14196,N_14419);
and U14942 (N_14942,N_14323,N_14247);
nor U14943 (N_14943,N_14165,N_14287);
nand U14944 (N_14944,N_14303,N_14129);
xnor U14945 (N_14945,N_14437,N_14245);
and U14946 (N_14946,N_14213,N_14131);
nor U14947 (N_14947,N_14392,N_14495);
or U14948 (N_14948,N_14032,N_14188);
and U14949 (N_14949,N_14378,N_14427);
or U14950 (N_14950,N_14365,N_14332);
xnor U14951 (N_14951,N_14201,N_14336);
or U14952 (N_14952,N_14220,N_14166);
nor U14953 (N_14953,N_14258,N_14352);
nor U14954 (N_14954,N_14319,N_14446);
nor U14955 (N_14955,N_14300,N_14463);
or U14956 (N_14956,N_14281,N_14457);
nand U14957 (N_14957,N_14402,N_14059);
nor U14958 (N_14958,N_14392,N_14250);
xnor U14959 (N_14959,N_14397,N_14238);
nand U14960 (N_14960,N_14085,N_14267);
and U14961 (N_14961,N_14122,N_14262);
nor U14962 (N_14962,N_14384,N_14138);
or U14963 (N_14963,N_14107,N_14118);
nand U14964 (N_14964,N_14393,N_14322);
nor U14965 (N_14965,N_14305,N_14294);
nand U14966 (N_14966,N_14361,N_14100);
or U14967 (N_14967,N_14277,N_14208);
nor U14968 (N_14968,N_14308,N_14070);
or U14969 (N_14969,N_14169,N_14411);
nor U14970 (N_14970,N_14381,N_14276);
xnor U14971 (N_14971,N_14418,N_14281);
and U14972 (N_14972,N_14030,N_14154);
nand U14973 (N_14973,N_14261,N_14339);
nor U14974 (N_14974,N_14417,N_14031);
nand U14975 (N_14975,N_14204,N_14423);
nor U14976 (N_14976,N_14115,N_14212);
nand U14977 (N_14977,N_14320,N_14459);
xor U14978 (N_14978,N_14423,N_14272);
or U14979 (N_14979,N_14466,N_14311);
nand U14980 (N_14980,N_14012,N_14004);
xor U14981 (N_14981,N_14216,N_14395);
nand U14982 (N_14982,N_14184,N_14257);
xor U14983 (N_14983,N_14017,N_14329);
nor U14984 (N_14984,N_14376,N_14448);
nand U14985 (N_14985,N_14166,N_14067);
xnor U14986 (N_14986,N_14084,N_14487);
and U14987 (N_14987,N_14386,N_14218);
nand U14988 (N_14988,N_14095,N_14327);
nand U14989 (N_14989,N_14451,N_14393);
or U14990 (N_14990,N_14228,N_14265);
and U14991 (N_14991,N_14457,N_14421);
nand U14992 (N_14992,N_14042,N_14466);
nand U14993 (N_14993,N_14076,N_14499);
nand U14994 (N_14994,N_14488,N_14476);
and U14995 (N_14995,N_14286,N_14032);
nor U14996 (N_14996,N_14347,N_14222);
xnor U14997 (N_14997,N_14281,N_14116);
xnor U14998 (N_14998,N_14152,N_14121);
and U14999 (N_14999,N_14359,N_14030);
and UO_0 (O_0,N_14654,N_14664);
and UO_1 (O_1,N_14560,N_14824);
xor UO_2 (O_2,N_14571,N_14954);
xnor UO_3 (O_3,N_14676,N_14886);
nand UO_4 (O_4,N_14967,N_14862);
nand UO_5 (O_5,N_14830,N_14696);
or UO_6 (O_6,N_14625,N_14586);
xor UO_7 (O_7,N_14906,N_14840);
xor UO_8 (O_8,N_14945,N_14507);
nor UO_9 (O_9,N_14551,N_14624);
nor UO_10 (O_10,N_14899,N_14759);
or UO_11 (O_11,N_14666,N_14803);
xor UO_12 (O_12,N_14546,N_14744);
or UO_13 (O_13,N_14538,N_14526);
nor UO_14 (O_14,N_14589,N_14822);
nand UO_15 (O_15,N_14993,N_14806);
and UO_16 (O_16,N_14575,N_14962);
nand UO_17 (O_17,N_14860,N_14504);
and UO_18 (O_18,N_14807,N_14880);
xor UO_19 (O_19,N_14535,N_14980);
or UO_20 (O_20,N_14726,N_14528);
and UO_21 (O_21,N_14653,N_14606);
and UO_22 (O_22,N_14952,N_14835);
nand UO_23 (O_23,N_14969,N_14739);
or UO_24 (O_24,N_14770,N_14976);
and UO_25 (O_25,N_14693,N_14553);
xnor UO_26 (O_26,N_14940,N_14794);
nand UO_27 (O_27,N_14821,N_14787);
xor UO_28 (O_28,N_14673,N_14556);
nand UO_29 (O_29,N_14772,N_14585);
xnor UO_30 (O_30,N_14718,N_14631);
or UO_31 (O_31,N_14518,N_14508);
nand UO_32 (O_32,N_14709,N_14514);
and UO_33 (O_33,N_14800,N_14846);
xnor UO_34 (O_34,N_14655,N_14557);
or UO_35 (O_35,N_14513,N_14876);
xor UO_36 (O_36,N_14939,N_14684);
or UO_37 (O_37,N_14836,N_14501);
or UO_38 (O_38,N_14647,N_14651);
nand UO_39 (O_39,N_14865,N_14619);
nand UO_40 (O_40,N_14713,N_14905);
nor UO_41 (O_41,N_14533,N_14930);
nand UO_42 (O_42,N_14725,N_14804);
nor UO_43 (O_43,N_14764,N_14755);
nor UO_44 (O_44,N_14889,N_14790);
or UO_45 (O_45,N_14628,N_14791);
and UO_46 (O_46,N_14861,N_14638);
nor UO_47 (O_47,N_14616,N_14925);
or UO_48 (O_48,N_14531,N_14555);
xor UO_49 (O_49,N_14918,N_14736);
or UO_50 (O_50,N_14750,N_14866);
and UO_51 (O_51,N_14611,N_14885);
xnor UO_52 (O_52,N_14541,N_14809);
nand UO_53 (O_53,N_14982,N_14833);
and UO_54 (O_54,N_14748,N_14639);
or UO_55 (O_55,N_14687,N_14933);
or UO_56 (O_56,N_14977,N_14956);
nor UO_57 (O_57,N_14763,N_14966);
xor UO_58 (O_58,N_14715,N_14594);
nor UO_59 (O_59,N_14892,N_14608);
xor UO_60 (O_60,N_14743,N_14714);
and UO_61 (O_61,N_14922,N_14949);
nor UO_62 (O_62,N_14900,N_14968);
nand UO_63 (O_63,N_14587,N_14641);
or UO_64 (O_64,N_14574,N_14988);
nand UO_65 (O_65,N_14847,N_14838);
nor UO_66 (O_66,N_14622,N_14707);
or UO_67 (O_67,N_14563,N_14771);
or UO_68 (O_68,N_14853,N_14576);
nand UO_69 (O_69,N_14991,N_14815);
and UO_70 (O_70,N_14500,N_14592);
nor UO_71 (O_71,N_14682,N_14566);
nand UO_72 (O_72,N_14706,N_14694);
xnor UO_73 (O_73,N_14524,N_14916);
nand UO_74 (O_74,N_14510,N_14747);
or UO_75 (O_75,N_14786,N_14637);
xor UO_76 (O_76,N_14642,N_14699);
or UO_77 (O_77,N_14947,N_14797);
or UO_78 (O_78,N_14636,N_14702);
nand UO_79 (O_79,N_14875,N_14506);
and UO_80 (O_80,N_14908,N_14970);
xor UO_81 (O_81,N_14542,N_14537);
nand UO_82 (O_82,N_14893,N_14527);
xnor UO_83 (O_83,N_14891,N_14859);
xnor UO_84 (O_84,N_14521,N_14643);
or UO_85 (O_85,N_14850,N_14897);
nand UO_86 (O_86,N_14870,N_14722);
xnor UO_87 (O_87,N_14887,N_14584);
or UO_88 (O_88,N_14590,N_14998);
xnor UO_89 (O_89,N_14517,N_14877);
nor UO_90 (O_90,N_14519,N_14627);
nand UO_91 (O_91,N_14832,N_14857);
xor UO_92 (O_92,N_14564,N_14728);
nor UO_93 (O_93,N_14766,N_14650);
xnor UO_94 (O_94,N_14935,N_14516);
nand UO_95 (O_95,N_14737,N_14547);
or UO_96 (O_96,N_14769,N_14668);
nand UO_97 (O_97,N_14931,N_14689);
xnor UO_98 (O_98,N_14754,N_14963);
or UO_99 (O_99,N_14663,N_14974);
nor UO_100 (O_100,N_14789,N_14792);
nor UO_101 (O_101,N_14995,N_14680);
or UO_102 (O_102,N_14843,N_14649);
xor UO_103 (O_103,N_14529,N_14894);
or UO_104 (O_104,N_14544,N_14734);
or UO_105 (O_105,N_14831,N_14983);
or UO_106 (O_106,N_14955,N_14674);
and UO_107 (O_107,N_14697,N_14598);
nor UO_108 (O_108,N_14614,N_14730);
nand UO_109 (O_109,N_14914,N_14757);
xor UO_110 (O_110,N_14758,N_14852);
nand UO_111 (O_111,N_14999,N_14536);
and UO_112 (O_112,N_14996,N_14779);
or UO_113 (O_113,N_14767,N_14733);
or UO_114 (O_114,N_14872,N_14826);
nand UO_115 (O_115,N_14841,N_14973);
nor UO_116 (O_116,N_14583,N_14796);
nand UO_117 (O_117,N_14640,N_14581);
nor UO_118 (O_118,N_14670,N_14912);
nor UO_119 (O_119,N_14749,N_14633);
or UO_120 (O_120,N_14515,N_14570);
or UO_121 (O_121,N_14957,N_14958);
nor UO_122 (O_122,N_14927,N_14868);
and UO_123 (O_123,N_14879,N_14992);
and UO_124 (O_124,N_14823,N_14729);
nand UO_125 (O_125,N_14740,N_14910);
or UO_126 (O_126,N_14632,N_14812);
and UO_127 (O_127,N_14675,N_14793);
nor UO_128 (O_128,N_14985,N_14530);
nand UO_129 (O_129,N_14903,N_14782);
and UO_130 (O_130,N_14657,N_14591);
or UO_131 (O_131,N_14677,N_14617);
and UO_132 (O_132,N_14741,N_14950);
xor UO_133 (O_133,N_14781,N_14981);
nor UO_134 (O_134,N_14686,N_14817);
and UO_135 (O_135,N_14856,N_14562);
or UO_136 (O_136,N_14871,N_14610);
nor UO_137 (O_137,N_14929,N_14944);
nand UO_138 (O_138,N_14540,N_14788);
or UO_139 (O_139,N_14690,N_14735);
xor UO_140 (O_140,N_14844,N_14780);
nand UO_141 (O_141,N_14795,N_14760);
nor UO_142 (O_142,N_14612,N_14921);
and UO_143 (O_143,N_14678,N_14774);
and UO_144 (O_144,N_14805,N_14669);
xnor UO_145 (O_145,N_14705,N_14503);
xnor UO_146 (O_146,N_14660,N_14762);
or UO_147 (O_147,N_14913,N_14723);
nand UO_148 (O_148,N_14549,N_14652);
nor UO_149 (O_149,N_14882,N_14842);
xor UO_150 (O_150,N_14602,N_14588);
nand UO_151 (O_151,N_14601,N_14813);
and UO_152 (O_152,N_14942,N_14811);
or UO_153 (O_153,N_14600,N_14828);
nand UO_154 (O_154,N_14634,N_14580);
and UO_155 (O_155,N_14646,N_14569);
or UO_156 (O_156,N_14665,N_14845);
or UO_157 (O_157,N_14911,N_14878);
and UO_158 (O_158,N_14511,N_14727);
and UO_159 (O_159,N_14672,N_14884);
and UO_160 (O_160,N_14520,N_14621);
nor UO_161 (O_161,N_14512,N_14599);
nand UO_162 (O_162,N_14827,N_14953);
nand UO_163 (O_163,N_14658,N_14579);
nand UO_164 (O_164,N_14979,N_14773);
or UO_165 (O_165,N_14550,N_14742);
and UO_166 (O_166,N_14543,N_14907);
and UO_167 (O_167,N_14717,N_14946);
nor UO_168 (O_168,N_14923,N_14909);
or UO_169 (O_169,N_14752,N_14685);
xnor UO_170 (O_170,N_14799,N_14902);
nand UO_171 (O_171,N_14924,N_14895);
and UO_172 (O_172,N_14716,N_14618);
nor UO_173 (O_173,N_14644,N_14656);
and UO_174 (O_174,N_14607,N_14597);
or UO_175 (O_175,N_14578,N_14552);
xnor UO_176 (O_176,N_14888,N_14839);
or UO_177 (O_177,N_14701,N_14765);
nand UO_178 (O_178,N_14561,N_14761);
xnor UO_179 (O_179,N_14623,N_14881);
nand UO_180 (O_180,N_14573,N_14681);
nand UO_181 (O_181,N_14959,N_14784);
nor UO_182 (O_182,N_14820,N_14915);
or UO_183 (O_183,N_14802,N_14932);
or UO_184 (O_184,N_14509,N_14997);
nand UO_185 (O_185,N_14648,N_14943);
nor UO_186 (O_186,N_14712,N_14937);
and UO_187 (O_187,N_14753,N_14635);
or UO_188 (O_188,N_14626,N_14534);
or UO_189 (O_189,N_14818,N_14711);
nor UO_190 (O_190,N_14990,N_14559);
xor UO_191 (O_191,N_14720,N_14928);
nand UO_192 (O_192,N_14603,N_14890);
nor UO_193 (O_193,N_14719,N_14816);
or UO_194 (O_194,N_14691,N_14898);
nand UO_195 (O_195,N_14941,N_14863);
and UO_196 (O_196,N_14938,N_14874);
xor UO_197 (O_197,N_14746,N_14873);
nand UO_198 (O_198,N_14775,N_14867);
or UO_199 (O_199,N_14810,N_14698);
xor UO_200 (O_200,N_14572,N_14819);
and UO_201 (O_201,N_14778,N_14522);
nand UO_202 (O_202,N_14776,N_14978);
xor UO_203 (O_203,N_14936,N_14994);
nor UO_204 (O_204,N_14703,N_14904);
xor UO_205 (O_205,N_14629,N_14724);
nand UO_206 (O_206,N_14984,N_14738);
xnor UO_207 (O_207,N_14849,N_14613);
xnor UO_208 (O_208,N_14987,N_14808);
xor UO_209 (O_209,N_14539,N_14645);
nor UO_210 (O_210,N_14934,N_14558);
nor UO_211 (O_211,N_14986,N_14692);
or UO_212 (O_212,N_14731,N_14783);
xor UO_213 (O_213,N_14896,N_14568);
nor UO_214 (O_214,N_14864,N_14751);
or UO_215 (O_215,N_14554,N_14700);
nand UO_216 (O_216,N_14567,N_14960);
or UO_217 (O_217,N_14834,N_14683);
and UO_218 (O_218,N_14785,N_14756);
nor UO_219 (O_219,N_14695,N_14883);
xor UO_220 (O_220,N_14964,N_14667);
nor UO_221 (O_221,N_14525,N_14801);
nand UO_222 (O_222,N_14661,N_14565);
or UO_223 (O_223,N_14965,N_14721);
xnor UO_224 (O_224,N_14605,N_14659);
or UO_225 (O_225,N_14951,N_14502);
nand UO_226 (O_226,N_14975,N_14829);
nor UO_227 (O_227,N_14593,N_14577);
nand UO_228 (O_228,N_14768,N_14825);
or UO_229 (O_229,N_14596,N_14777);
nor UO_230 (O_230,N_14523,N_14798);
and UO_231 (O_231,N_14545,N_14837);
nand UO_232 (O_232,N_14869,N_14620);
nor UO_233 (O_233,N_14630,N_14971);
nor UO_234 (O_234,N_14732,N_14604);
xnor UO_235 (O_235,N_14972,N_14505);
xnor UO_236 (O_236,N_14595,N_14609);
nand UO_237 (O_237,N_14919,N_14855);
nand UO_238 (O_238,N_14532,N_14615);
xnor UO_239 (O_239,N_14745,N_14548);
and UO_240 (O_240,N_14961,N_14688);
xor UO_241 (O_241,N_14671,N_14858);
and UO_242 (O_242,N_14848,N_14920);
xor UO_243 (O_243,N_14851,N_14901);
nor UO_244 (O_244,N_14662,N_14704);
xor UO_245 (O_245,N_14708,N_14854);
and UO_246 (O_246,N_14582,N_14948);
nor UO_247 (O_247,N_14989,N_14710);
and UO_248 (O_248,N_14917,N_14926);
or UO_249 (O_249,N_14679,N_14814);
xor UO_250 (O_250,N_14953,N_14666);
or UO_251 (O_251,N_14724,N_14951);
nand UO_252 (O_252,N_14810,N_14876);
and UO_253 (O_253,N_14716,N_14980);
and UO_254 (O_254,N_14687,N_14952);
nor UO_255 (O_255,N_14921,N_14557);
xnor UO_256 (O_256,N_14673,N_14719);
nand UO_257 (O_257,N_14591,N_14669);
nor UO_258 (O_258,N_14561,N_14662);
xor UO_259 (O_259,N_14850,N_14924);
and UO_260 (O_260,N_14547,N_14767);
xor UO_261 (O_261,N_14952,N_14523);
or UO_262 (O_262,N_14537,N_14644);
nand UO_263 (O_263,N_14609,N_14837);
or UO_264 (O_264,N_14716,N_14604);
nor UO_265 (O_265,N_14948,N_14937);
nand UO_266 (O_266,N_14650,N_14613);
nor UO_267 (O_267,N_14943,N_14999);
xor UO_268 (O_268,N_14701,N_14936);
nor UO_269 (O_269,N_14984,N_14788);
nand UO_270 (O_270,N_14518,N_14616);
xor UO_271 (O_271,N_14607,N_14923);
nor UO_272 (O_272,N_14956,N_14528);
and UO_273 (O_273,N_14792,N_14755);
xor UO_274 (O_274,N_14965,N_14839);
xor UO_275 (O_275,N_14782,N_14943);
nand UO_276 (O_276,N_14849,N_14600);
and UO_277 (O_277,N_14622,N_14936);
and UO_278 (O_278,N_14900,N_14918);
nand UO_279 (O_279,N_14857,N_14531);
nor UO_280 (O_280,N_14837,N_14546);
and UO_281 (O_281,N_14786,N_14729);
and UO_282 (O_282,N_14824,N_14648);
xnor UO_283 (O_283,N_14663,N_14500);
nor UO_284 (O_284,N_14911,N_14988);
nand UO_285 (O_285,N_14906,N_14773);
or UO_286 (O_286,N_14806,N_14930);
nand UO_287 (O_287,N_14899,N_14878);
xnor UO_288 (O_288,N_14511,N_14792);
and UO_289 (O_289,N_14715,N_14861);
and UO_290 (O_290,N_14913,N_14717);
xor UO_291 (O_291,N_14735,N_14874);
and UO_292 (O_292,N_14740,N_14845);
and UO_293 (O_293,N_14514,N_14752);
and UO_294 (O_294,N_14605,N_14619);
xnor UO_295 (O_295,N_14510,N_14643);
and UO_296 (O_296,N_14650,N_14674);
xor UO_297 (O_297,N_14520,N_14997);
or UO_298 (O_298,N_14976,N_14714);
nand UO_299 (O_299,N_14911,N_14541);
and UO_300 (O_300,N_14624,N_14642);
or UO_301 (O_301,N_14875,N_14933);
nor UO_302 (O_302,N_14728,N_14885);
xnor UO_303 (O_303,N_14643,N_14981);
or UO_304 (O_304,N_14714,N_14610);
and UO_305 (O_305,N_14634,N_14617);
nand UO_306 (O_306,N_14858,N_14755);
nor UO_307 (O_307,N_14719,N_14712);
nor UO_308 (O_308,N_14521,N_14759);
nand UO_309 (O_309,N_14567,N_14592);
nor UO_310 (O_310,N_14861,N_14947);
nor UO_311 (O_311,N_14812,N_14702);
nor UO_312 (O_312,N_14656,N_14567);
and UO_313 (O_313,N_14606,N_14502);
and UO_314 (O_314,N_14664,N_14775);
nor UO_315 (O_315,N_14677,N_14788);
and UO_316 (O_316,N_14614,N_14644);
nand UO_317 (O_317,N_14989,N_14988);
nand UO_318 (O_318,N_14698,N_14543);
xnor UO_319 (O_319,N_14526,N_14768);
and UO_320 (O_320,N_14820,N_14860);
nor UO_321 (O_321,N_14816,N_14916);
nor UO_322 (O_322,N_14802,N_14642);
nand UO_323 (O_323,N_14509,N_14752);
xnor UO_324 (O_324,N_14850,N_14974);
and UO_325 (O_325,N_14994,N_14975);
and UO_326 (O_326,N_14817,N_14616);
nand UO_327 (O_327,N_14968,N_14827);
nor UO_328 (O_328,N_14758,N_14769);
or UO_329 (O_329,N_14993,N_14882);
or UO_330 (O_330,N_14671,N_14552);
nand UO_331 (O_331,N_14694,N_14959);
nor UO_332 (O_332,N_14720,N_14995);
xor UO_333 (O_333,N_14576,N_14633);
or UO_334 (O_334,N_14943,N_14696);
and UO_335 (O_335,N_14728,N_14961);
xnor UO_336 (O_336,N_14844,N_14779);
and UO_337 (O_337,N_14821,N_14833);
or UO_338 (O_338,N_14726,N_14907);
and UO_339 (O_339,N_14904,N_14548);
and UO_340 (O_340,N_14553,N_14840);
and UO_341 (O_341,N_14913,N_14882);
or UO_342 (O_342,N_14585,N_14780);
xor UO_343 (O_343,N_14673,N_14574);
nor UO_344 (O_344,N_14556,N_14762);
xor UO_345 (O_345,N_14892,N_14837);
nor UO_346 (O_346,N_14867,N_14642);
xnor UO_347 (O_347,N_14594,N_14941);
and UO_348 (O_348,N_14549,N_14726);
nor UO_349 (O_349,N_14985,N_14986);
xor UO_350 (O_350,N_14864,N_14546);
xor UO_351 (O_351,N_14629,N_14803);
and UO_352 (O_352,N_14742,N_14673);
or UO_353 (O_353,N_14805,N_14715);
nor UO_354 (O_354,N_14557,N_14514);
nor UO_355 (O_355,N_14679,N_14905);
and UO_356 (O_356,N_14927,N_14504);
or UO_357 (O_357,N_14926,N_14523);
nand UO_358 (O_358,N_14930,N_14609);
or UO_359 (O_359,N_14554,N_14935);
xnor UO_360 (O_360,N_14986,N_14577);
nand UO_361 (O_361,N_14760,N_14990);
and UO_362 (O_362,N_14666,N_14667);
or UO_363 (O_363,N_14948,N_14844);
nand UO_364 (O_364,N_14574,N_14709);
nand UO_365 (O_365,N_14785,N_14919);
xor UO_366 (O_366,N_14704,N_14913);
nand UO_367 (O_367,N_14917,N_14558);
nand UO_368 (O_368,N_14987,N_14891);
nand UO_369 (O_369,N_14945,N_14797);
nor UO_370 (O_370,N_14697,N_14768);
or UO_371 (O_371,N_14740,N_14514);
nor UO_372 (O_372,N_14770,N_14551);
nand UO_373 (O_373,N_14683,N_14861);
and UO_374 (O_374,N_14848,N_14734);
or UO_375 (O_375,N_14778,N_14715);
and UO_376 (O_376,N_14748,N_14587);
or UO_377 (O_377,N_14520,N_14818);
nor UO_378 (O_378,N_14922,N_14682);
xor UO_379 (O_379,N_14544,N_14802);
nor UO_380 (O_380,N_14574,N_14677);
xnor UO_381 (O_381,N_14989,N_14849);
xor UO_382 (O_382,N_14935,N_14923);
and UO_383 (O_383,N_14600,N_14715);
nor UO_384 (O_384,N_14779,N_14648);
xnor UO_385 (O_385,N_14540,N_14823);
and UO_386 (O_386,N_14954,N_14758);
and UO_387 (O_387,N_14679,N_14987);
or UO_388 (O_388,N_14687,N_14968);
xor UO_389 (O_389,N_14688,N_14686);
or UO_390 (O_390,N_14619,N_14695);
nor UO_391 (O_391,N_14887,N_14938);
and UO_392 (O_392,N_14836,N_14582);
and UO_393 (O_393,N_14625,N_14536);
xor UO_394 (O_394,N_14930,N_14532);
and UO_395 (O_395,N_14621,N_14688);
nor UO_396 (O_396,N_14847,N_14745);
nand UO_397 (O_397,N_14880,N_14840);
nand UO_398 (O_398,N_14723,N_14684);
xor UO_399 (O_399,N_14668,N_14891);
or UO_400 (O_400,N_14802,N_14950);
and UO_401 (O_401,N_14627,N_14652);
nor UO_402 (O_402,N_14952,N_14859);
and UO_403 (O_403,N_14640,N_14773);
and UO_404 (O_404,N_14577,N_14709);
and UO_405 (O_405,N_14869,N_14981);
nand UO_406 (O_406,N_14785,N_14933);
and UO_407 (O_407,N_14567,N_14843);
xor UO_408 (O_408,N_14596,N_14618);
nand UO_409 (O_409,N_14630,N_14799);
nand UO_410 (O_410,N_14794,N_14933);
nor UO_411 (O_411,N_14857,N_14787);
nor UO_412 (O_412,N_14608,N_14911);
xnor UO_413 (O_413,N_14840,N_14846);
xor UO_414 (O_414,N_14760,N_14978);
nand UO_415 (O_415,N_14711,N_14649);
or UO_416 (O_416,N_14618,N_14930);
or UO_417 (O_417,N_14946,N_14745);
or UO_418 (O_418,N_14809,N_14691);
xnor UO_419 (O_419,N_14885,N_14896);
nor UO_420 (O_420,N_14612,N_14732);
or UO_421 (O_421,N_14894,N_14575);
xnor UO_422 (O_422,N_14980,N_14784);
nand UO_423 (O_423,N_14787,N_14941);
xnor UO_424 (O_424,N_14931,N_14610);
xnor UO_425 (O_425,N_14547,N_14916);
xnor UO_426 (O_426,N_14521,N_14932);
nand UO_427 (O_427,N_14838,N_14986);
nor UO_428 (O_428,N_14668,N_14600);
or UO_429 (O_429,N_14656,N_14858);
nor UO_430 (O_430,N_14800,N_14535);
or UO_431 (O_431,N_14863,N_14653);
nor UO_432 (O_432,N_14582,N_14914);
nor UO_433 (O_433,N_14604,N_14582);
xor UO_434 (O_434,N_14601,N_14919);
or UO_435 (O_435,N_14760,N_14606);
nor UO_436 (O_436,N_14737,N_14643);
nand UO_437 (O_437,N_14547,N_14743);
xnor UO_438 (O_438,N_14765,N_14884);
xor UO_439 (O_439,N_14704,N_14842);
nor UO_440 (O_440,N_14549,N_14933);
xor UO_441 (O_441,N_14998,N_14871);
xnor UO_442 (O_442,N_14602,N_14988);
nand UO_443 (O_443,N_14801,N_14500);
nand UO_444 (O_444,N_14779,N_14786);
or UO_445 (O_445,N_14788,N_14639);
nand UO_446 (O_446,N_14693,N_14695);
and UO_447 (O_447,N_14716,N_14886);
nand UO_448 (O_448,N_14927,N_14737);
nand UO_449 (O_449,N_14653,N_14611);
or UO_450 (O_450,N_14714,N_14843);
or UO_451 (O_451,N_14904,N_14829);
nand UO_452 (O_452,N_14817,N_14691);
nor UO_453 (O_453,N_14583,N_14979);
nor UO_454 (O_454,N_14514,N_14561);
or UO_455 (O_455,N_14749,N_14594);
nand UO_456 (O_456,N_14660,N_14920);
xnor UO_457 (O_457,N_14881,N_14723);
nor UO_458 (O_458,N_14593,N_14695);
and UO_459 (O_459,N_14956,N_14721);
nand UO_460 (O_460,N_14922,N_14751);
or UO_461 (O_461,N_14526,N_14658);
nor UO_462 (O_462,N_14801,N_14967);
and UO_463 (O_463,N_14863,N_14637);
and UO_464 (O_464,N_14600,N_14573);
xnor UO_465 (O_465,N_14678,N_14727);
xor UO_466 (O_466,N_14729,N_14572);
nand UO_467 (O_467,N_14626,N_14704);
nor UO_468 (O_468,N_14979,N_14525);
xor UO_469 (O_469,N_14784,N_14750);
or UO_470 (O_470,N_14912,N_14624);
and UO_471 (O_471,N_14948,N_14727);
or UO_472 (O_472,N_14709,N_14809);
nand UO_473 (O_473,N_14693,N_14670);
xnor UO_474 (O_474,N_14821,N_14928);
or UO_475 (O_475,N_14655,N_14616);
or UO_476 (O_476,N_14546,N_14960);
nor UO_477 (O_477,N_14899,N_14502);
nor UO_478 (O_478,N_14810,N_14945);
nand UO_479 (O_479,N_14957,N_14551);
xnor UO_480 (O_480,N_14785,N_14975);
nor UO_481 (O_481,N_14524,N_14898);
nor UO_482 (O_482,N_14522,N_14951);
and UO_483 (O_483,N_14793,N_14875);
nor UO_484 (O_484,N_14667,N_14739);
nor UO_485 (O_485,N_14635,N_14683);
nand UO_486 (O_486,N_14751,N_14789);
and UO_487 (O_487,N_14830,N_14952);
nor UO_488 (O_488,N_14717,N_14568);
nor UO_489 (O_489,N_14684,N_14670);
xnor UO_490 (O_490,N_14526,N_14751);
or UO_491 (O_491,N_14683,N_14652);
or UO_492 (O_492,N_14989,N_14929);
xor UO_493 (O_493,N_14629,N_14812);
and UO_494 (O_494,N_14862,N_14812);
nand UO_495 (O_495,N_14977,N_14830);
xnor UO_496 (O_496,N_14979,N_14554);
nand UO_497 (O_497,N_14837,N_14905);
and UO_498 (O_498,N_14991,N_14651);
xor UO_499 (O_499,N_14843,N_14638);
nand UO_500 (O_500,N_14708,N_14845);
nor UO_501 (O_501,N_14971,N_14870);
and UO_502 (O_502,N_14558,N_14849);
or UO_503 (O_503,N_14939,N_14680);
xor UO_504 (O_504,N_14902,N_14966);
and UO_505 (O_505,N_14969,N_14545);
nor UO_506 (O_506,N_14968,N_14787);
nor UO_507 (O_507,N_14892,N_14590);
or UO_508 (O_508,N_14617,N_14882);
xor UO_509 (O_509,N_14904,N_14516);
and UO_510 (O_510,N_14638,N_14817);
nor UO_511 (O_511,N_14545,N_14916);
xor UO_512 (O_512,N_14585,N_14706);
nand UO_513 (O_513,N_14633,N_14856);
and UO_514 (O_514,N_14644,N_14910);
nand UO_515 (O_515,N_14822,N_14755);
nor UO_516 (O_516,N_14808,N_14984);
or UO_517 (O_517,N_14917,N_14891);
and UO_518 (O_518,N_14568,N_14579);
xnor UO_519 (O_519,N_14655,N_14856);
or UO_520 (O_520,N_14754,N_14504);
nor UO_521 (O_521,N_14723,N_14780);
nor UO_522 (O_522,N_14877,N_14888);
nand UO_523 (O_523,N_14785,N_14518);
and UO_524 (O_524,N_14900,N_14578);
xor UO_525 (O_525,N_14680,N_14736);
xor UO_526 (O_526,N_14987,N_14558);
and UO_527 (O_527,N_14683,N_14629);
nor UO_528 (O_528,N_14594,N_14797);
xnor UO_529 (O_529,N_14538,N_14723);
nor UO_530 (O_530,N_14697,N_14658);
or UO_531 (O_531,N_14724,N_14829);
nand UO_532 (O_532,N_14750,N_14831);
or UO_533 (O_533,N_14819,N_14674);
or UO_534 (O_534,N_14937,N_14573);
nor UO_535 (O_535,N_14670,N_14519);
nand UO_536 (O_536,N_14941,N_14687);
xor UO_537 (O_537,N_14828,N_14981);
nand UO_538 (O_538,N_14783,N_14509);
xor UO_539 (O_539,N_14859,N_14847);
or UO_540 (O_540,N_14654,N_14515);
nor UO_541 (O_541,N_14687,N_14819);
xor UO_542 (O_542,N_14772,N_14965);
nor UO_543 (O_543,N_14995,N_14674);
nand UO_544 (O_544,N_14866,N_14624);
or UO_545 (O_545,N_14863,N_14792);
nor UO_546 (O_546,N_14584,N_14752);
xnor UO_547 (O_547,N_14554,N_14645);
nand UO_548 (O_548,N_14998,N_14894);
and UO_549 (O_549,N_14814,N_14720);
or UO_550 (O_550,N_14907,N_14692);
nand UO_551 (O_551,N_14644,N_14691);
or UO_552 (O_552,N_14993,N_14622);
or UO_553 (O_553,N_14949,N_14565);
or UO_554 (O_554,N_14848,N_14789);
xor UO_555 (O_555,N_14511,N_14573);
nor UO_556 (O_556,N_14994,N_14804);
nor UO_557 (O_557,N_14820,N_14638);
nor UO_558 (O_558,N_14824,N_14606);
nand UO_559 (O_559,N_14663,N_14655);
nand UO_560 (O_560,N_14856,N_14682);
nand UO_561 (O_561,N_14945,N_14596);
nand UO_562 (O_562,N_14945,N_14629);
nor UO_563 (O_563,N_14714,N_14865);
and UO_564 (O_564,N_14902,N_14739);
and UO_565 (O_565,N_14554,N_14668);
or UO_566 (O_566,N_14538,N_14567);
and UO_567 (O_567,N_14747,N_14611);
or UO_568 (O_568,N_14622,N_14732);
xnor UO_569 (O_569,N_14933,N_14878);
or UO_570 (O_570,N_14723,N_14787);
and UO_571 (O_571,N_14656,N_14801);
xor UO_572 (O_572,N_14785,N_14574);
and UO_573 (O_573,N_14634,N_14652);
and UO_574 (O_574,N_14996,N_14807);
xor UO_575 (O_575,N_14514,N_14963);
nor UO_576 (O_576,N_14702,N_14907);
and UO_577 (O_577,N_14759,N_14952);
and UO_578 (O_578,N_14895,N_14897);
xnor UO_579 (O_579,N_14986,N_14814);
nand UO_580 (O_580,N_14525,N_14804);
or UO_581 (O_581,N_14840,N_14883);
nand UO_582 (O_582,N_14892,N_14749);
nand UO_583 (O_583,N_14743,N_14695);
or UO_584 (O_584,N_14651,N_14951);
nand UO_585 (O_585,N_14624,N_14900);
xor UO_586 (O_586,N_14880,N_14612);
xnor UO_587 (O_587,N_14782,N_14537);
and UO_588 (O_588,N_14844,N_14724);
xnor UO_589 (O_589,N_14961,N_14754);
nand UO_590 (O_590,N_14687,N_14746);
nor UO_591 (O_591,N_14655,N_14984);
xor UO_592 (O_592,N_14727,N_14990);
xor UO_593 (O_593,N_14996,N_14687);
nor UO_594 (O_594,N_14688,N_14902);
nor UO_595 (O_595,N_14603,N_14959);
and UO_596 (O_596,N_14680,N_14948);
or UO_597 (O_597,N_14560,N_14943);
and UO_598 (O_598,N_14744,N_14717);
and UO_599 (O_599,N_14931,N_14786);
or UO_600 (O_600,N_14589,N_14543);
and UO_601 (O_601,N_14636,N_14645);
or UO_602 (O_602,N_14925,N_14672);
xor UO_603 (O_603,N_14766,N_14978);
and UO_604 (O_604,N_14528,N_14842);
xnor UO_605 (O_605,N_14789,N_14928);
or UO_606 (O_606,N_14792,N_14799);
xnor UO_607 (O_607,N_14765,N_14907);
and UO_608 (O_608,N_14657,N_14554);
nand UO_609 (O_609,N_14705,N_14923);
xor UO_610 (O_610,N_14952,N_14515);
xnor UO_611 (O_611,N_14856,N_14935);
xnor UO_612 (O_612,N_14935,N_14934);
nor UO_613 (O_613,N_14533,N_14544);
and UO_614 (O_614,N_14766,N_14615);
nand UO_615 (O_615,N_14806,N_14605);
nand UO_616 (O_616,N_14796,N_14699);
xnor UO_617 (O_617,N_14939,N_14898);
or UO_618 (O_618,N_14761,N_14949);
or UO_619 (O_619,N_14826,N_14801);
or UO_620 (O_620,N_14857,N_14721);
xor UO_621 (O_621,N_14778,N_14842);
and UO_622 (O_622,N_14699,N_14912);
or UO_623 (O_623,N_14768,N_14974);
and UO_624 (O_624,N_14771,N_14846);
xnor UO_625 (O_625,N_14913,N_14881);
nor UO_626 (O_626,N_14877,N_14823);
nor UO_627 (O_627,N_14931,N_14914);
nor UO_628 (O_628,N_14655,N_14650);
or UO_629 (O_629,N_14729,N_14754);
nor UO_630 (O_630,N_14866,N_14899);
nor UO_631 (O_631,N_14704,N_14694);
or UO_632 (O_632,N_14766,N_14635);
or UO_633 (O_633,N_14885,N_14998);
nor UO_634 (O_634,N_14714,N_14746);
or UO_635 (O_635,N_14534,N_14840);
nand UO_636 (O_636,N_14813,N_14609);
and UO_637 (O_637,N_14562,N_14568);
xor UO_638 (O_638,N_14558,N_14678);
nor UO_639 (O_639,N_14547,N_14802);
nand UO_640 (O_640,N_14535,N_14705);
nand UO_641 (O_641,N_14801,N_14975);
xor UO_642 (O_642,N_14925,N_14637);
xnor UO_643 (O_643,N_14699,N_14557);
nor UO_644 (O_644,N_14715,N_14571);
xnor UO_645 (O_645,N_14710,N_14952);
nand UO_646 (O_646,N_14830,N_14886);
or UO_647 (O_647,N_14885,N_14868);
and UO_648 (O_648,N_14941,N_14599);
and UO_649 (O_649,N_14737,N_14881);
nand UO_650 (O_650,N_14818,N_14977);
xnor UO_651 (O_651,N_14777,N_14977);
xnor UO_652 (O_652,N_14930,N_14933);
and UO_653 (O_653,N_14884,N_14999);
nor UO_654 (O_654,N_14804,N_14645);
xor UO_655 (O_655,N_14868,N_14589);
xnor UO_656 (O_656,N_14943,N_14776);
xnor UO_657 (O_657,N_14890,N_14722);
or UO_658 (O_658,N_14964,N_14780);
nor UO_659 (O_659,N_14964,N_14713);
xnor UO_660 (O_660,N_14612,N_14764);
nor UO_661 (O_661,N_14809,N_14735);
or UO_662 (O_662,N_14861,N_14913);
or UO_663 (O_663,N_14823,N_14549);
xnor UO_664 (O_664,N_14661,N_14793);
or UO_665 (O_665,N_14717,N_14929);
nand UO_666 (O_666,N_14537,N_14877);
nand UO_667 (O_667,N_14572,N_14741);
or UO_668 (O_668,N_14799,N_14514);
and UO_669 (O_669,N_14852,N_14505);
or UO_670 (O_670,N_14921,N_14912);
xnor UO_671 (O_671,N_14565,N_14741);
xor UO_672 (O_672,N_14518,N_14834);
or UO_673 (O_673,N_14656,N_14550);
nor UO_674 (O_674,N_14759,N_14716);
or UO_675 (O_675,N_14773,N_14581);
and UO_676 (O_676,N_14725,N_14726);
nor UO_677 (O_677,N_14696,N_14642);
xor UO_678 (O_678,N_14830,N_14778);
or UO_679 (O_679,N_14788,N_14645);
nor UO_680 (O_680,N_14578,N_14949);
nor UO_681 (O_681,N_14904,N_14867);
xor UO_682 (O_682,N_14543,N_14560);
nor UO_683 (O_683,N_14577,N_14961);
or UO_684 (O_684,N_14547,N_14572);
nand UO_685 (O_685,N_14829,N_14687);
nand UO_686 (O_686,N_14921,N_14886);
and UO_687 (O_687,N_14592,N_14744);
or UO_688 (O_688,N_14827,N_14900);
and UO_689 (O_689,N_14526,N_14785);
xor UO_690 (O_690,N_14582,N_14832);
or UO_691 (O_691,N_14896,N_14549);
nor UO_692 (O_692,N_14776,N_14722);
xnor UO_693 (O_693,N_14521,N_14703);
xnor UO_694 (O_694,N_14805,N_14533);
xor UO_695 (O_695,N_14743,N_14907);
and UO_696 (O_696,N_14780,N_14744);
xor UO_697 (O_697,N_14724,N_14860);
nor UO_698 (O_698,N_14963,N_14699);
xnor UO_699 (O_699,N_14974,N_14861);
nand UO_700 (O_700,N_14860,N_14858);
xnor UO_701 (O_701,N_14652,N_14553);
nor UO_702 (O_702,N_14899,N_14804);
nand UO_703 (O_703,N_14856,N_14541);
nor UO_704 (O_704,N_14681,N_14632);
and UO_705 (O_705,N_14927,N_14813);
xnor UO_706 (O_706,N_14878,N_14905);
xor UO_707 (O_707,N_14683,N_14622);
nand UO_708 (O_708,N_14748,N_14528);
nor UO_709 (O_709,N_14685,N_14708);
xor UO_710 (O_710,N_14885,N_14971);
and UO_711 (O_711,N_14943,N_14811);
and UO_712 (O_712,N_14946,N_14768);
or UO_713 (O_713,N_14717,N_14846);
nand UO_714 (O_714,N_14717,N_14813);
nor UO_715 (O_715,N_14830,N_14906);
and UO_716 (O_716,N_14907,N_14682);
nor UO_717 (O_717,N_14657,N_14547);
xor UO_718 (O_718,N_14590,N_14954);
and UO_719 (O_719,N_14515,N_14895);
or UO_720 (O_720,N_14692,N_14619);
xnor UO_721 (O_721,N_14513,N_14548);
nand UO_722 (O_722,N_14663,N_14863);
xor UO_723 (O_723,N_14511,N_14655);
xor UO_724 (O_724,N_14912,N_14534);
nand UO_725 (O_725,N_14687,N_14672);
nor UO_726 (O_726,N_14544,N_14940);
xnor UO_727 (O_727,N_14550,N_14873);
and UO_728 (O_728,N_14739,N_14547);
xor UO_729 (O_729,N_14743,N_14610);
nand UO_730 (O_730,N_14569,N_14521);
or UO_731 (O_731,N_14637,N_14761);
and UO_732 (O_732,N_14918,N_14667);
or UO_733 (O_733,N_14843,N_14641);
and UO_734 (O_734,N_14692,N_14501);
nor UO_735 (O_735,N_14907,N_14569);
or UO_736 (O_736,N_14988,N_14666);
nand UO_737 (O_737,N_14888,N_14613);
nand UO_738 (O_738,N_14678,N_14753);
nand UO_739 (O_739,N_14591,N_14696);
or UO_740 (O_740,N_14544,N_14587);
or UO_741 (O_741,N_14822,N_14663);
nand UO_742 (O_742,N_14806,N_14650);
xnor UO_743 (O_743,N_14660,N_14545);
nand UO_744 (O_744,N_14842,N_14652);
or UO_745 (O_745,N_14718,N_14674);
xnor UO_746 (O_746,N_14573,N_14554);
xnor UO_747 (O_747,N_14638,N_14511);
nor UO_748 (O_748,N_14661,N_14866);
xnor UO_749 (O_749,N_14724,N_14599);
or UO_750 (O_750,N_14573,N_14712);
and UO_751 (O_751,N_14681,N_14548);
nor UO_752 (O_752,N_14673,N_14937);
and UO_753 (O_753,N_14725,N_14706);
and UO_754 (O_754,N_14928,N_14620);
nand UO_755 (O_755,N_14586,N_14753);
or UO_756 (O_756,N_14852,N_14695);
and UO_757 (O_757,N_14630,N_14672);
nand UO_758 (O_758,N_14721,N_14812);
nand UO_759 (O_759,N_14723,N_14747);
nor UO_760 (O_760,N_14749,N_14776);
and UO_761 (O_761,N_14755,N_14892);
nor UO_762 (O_762,N_14651,N_14666);
nor UO_763 (O_763,N_14605,N_14778);
xor UO_764 (O_764,N_14869,N_14673);
nand UO_765 (O_765,N_14724,N_14659);
nand UO_766 (O_766,N_14805,N_14643);
or UO_767 (O_767,N_14656,N_14705);
nor UO_768 (O_768,N_14540,N_14772);
xnor UO_769 (O_769,N_14764,N_14679);
and UO_770 (O_770,N_14860,N_14536);
nor UO_771 (O_771,N_14650,N_14550);
or UO_772 (O_772,N_14720,N_14733);
nand UO_773 (O_773,N_14501,N_14760);
nand UO_774 (O_774,N_14876,N_14595);
or UO_775 (O_775,N_14912,N_14785);
nor UO_776 (O_776,N_14865,N_14686);
nand UO_777 (O_777,N_14552,N_14779);
and UO_778 (O_778,N_14579,N_14819);
or UO_779 (O_779,N_14549,N_14564);
nor UO_780 (O_780,N_14721,N_14683);
nor UO_781 (O_781,N_14827,N_14903);
nor UO_782 (O_782,N_14637,N_14817);
nor UO_783 (O_783,N_14927,N_14662);
nand UO_784 (O_784,N_14727,N_14559);
xor UO_785 (O_785,N_14953,N_14740);
nor UO_786 (O_786,N_14918,N_14709);
xor UO_787 (O_787,N_14853,N_14868);
nor UO_788 (O_788,N_14819,N_14633);
xnor UO_789 (O_789,N_14585,N_14531);
and UO_790 (O_790,N_14935,N_14547);
or UO_791 (O_791,N_14850,N_14675);
xor UO_792 (O_792,N_14827,N_14517);
xor UO_793 (O_793,N_14593,N_14745);
nand UO_794 (O_794,N_14829,N_14783);
nor UO_795 (O_795,N_14971,N_14650);
nand UO_796 (O_796,N_14567,N_14618);
nor UO_797 (O_797,N_14761,N_14990);
or UO_798 (O_798,N_14949,N_14529);
nand UO_799 (O_799,N_14820,N_14895);
or UO_800 (O_800,N_14786,N_14608);
and UO_801 (O_801,N_14565,N_14826);
and UO_802 (O_802,N_14676,N_14707);
nand UO_803 (O_803,N_14702,N_14650);
nor UO_804 (O_804,N_14522,N_14502);
or UO_805 (O_805,N_14734,N_14653);
nor UO_806 (O_806,N_14564,N_14570);
and UO_807 (O_807,N_14580,N_14716);
and UO_808 (O_808,N_14657,N_14723);
and UO_809 (O_809,N_14706,N_14792);
and UO_810 (O_810,N_14574,N_14624);
nand UO_811 (O_811,N_14813,N_14552);
and UO_812 (O_812,N_14686,N_14878);
or UO_813 (O_813,N_14683,N_14596);
xnor UO_814 (O_814,N_14935,N_14860);
and UO_815 (O_815,N_14839,N_14926);
and UO_816 (O_816,N_14664,N_14607);
and UO_817 (O_817,N_14669,N_14851);
nand UO_818 (O_818,N_14997,N_14978);
nand UO_819 (O_819,N_14658,N_14946);
and UO_820 (O_820,N_14774,N_14664);
or UO_821 (O_821,N_14912,N_14705);
and UO_822 (O_822,N_14959,N_14976);
xor UO_823 (O_823,N_14515,N_14666);
or UO_824 (O_824,N_14846,N_14836);
nand UO_825 (O_825,N_14951,N_14999);
nor UO_826 (O_826,N_14855,N_14550);
xor UO_827 (O_827,N_14783,N_14894);
or UO_828 (O_828,N_14842,N_14659);
and UO_829 (O_829,N_14970,N_14872);
xnor UO_830 (O_830,N_14623,N_14817);
nand UO_831 (O_831,N_14601,N_14941);
nand UO_832 (O_832,N_14529,N_14527);
or UO_833 (O_833,N_14695,N_14796);
and UO_834 (O_834,N_14942,N_14762);
nand UO_835 (O_835,N_14865,N_14991);
xnor UO_836 (O_836,N_14513,N_14578);
and UO_837 (O_837,N_14632,N_14996);
and UO_838 (O_838,N_14769,N_14555);
and UO_839 (O_839,N_14831,N_14934);
nor UO_840 (O_840,N_14571,N_14522);
nor UO_841 (O_841,N_14849,N_14575);
or UO_842 (O_842,N_14867,N_14724);
xor UO_843 (O_843,N_14599,N_14665);
or UO_844 (O_844,N_14899,N_14998);
and UO_845 (O_845,N_14615,N_14935);
nand UO_846 (O_846,N_14860,N_14567);
nand UO_847 (O_847,N_14553,N_14802);
xor UO_848 (O_848,N_14802,N_14849);
nand UO_849 (O_849,N_14609,N_14614);
or UO_850 (O_850,N_14632,N_14825);
nand UO_851 (O_851,N_14885,N_14693);
or UO_852 (O_852,N_14940,N_14945);
or UO_853 (O_853,N_14864,N_14951);
xnor UO_854 (O_854,N_14869,N_14748);
nor UO_855 (O_855,N_14789,N_14582);
or UO_856 (O_856,N_14697,N_14873);
nand UO_857 (O_857,N_14691,N_14927);
xnor UO_858 (O_858,N_14596,N_14981);
or UO_859 (O_859,N_14620,N_14965);
xnor UO_860 (O_860,N_14794,N_14778);
nor UO_861 (O_861,N_14576,N_14520);
and UO_862 (O_862,N_14769,N_14551);
nand UO_863 (O_863,N_14712,N_14513);
xor UO_864 (O_864,N_14728,N_14858);
xor UO_865 (O_865,N_14894,N_14542);
xnor UO_866 (O_866,N_14771,N_14777);
xor UO_867 (O_867,N_14676,N_14922);
nand UO_868 (O_868,N_14798,N_14528);
and UO_869 (O_869,N_14896,N_14869);
and UO_870 (O_870,N_14850,N_14552);
and UO_871 (O_871,N_14797,N_14502);
nand UO_872 (O_872,N_14605,N_14552);
nor UO_873 (O_873,N_14657,N_14557);
xor UO_874 (O_874,N_14637,N_14810);
and UO_875 (O_875,N_14704,N_14906);
nor UO_876 (O_876,N_14557,N_14712);
or UO_877 (O_877,N_14838,N_14906);
and UO_878 (O_878,N_14947,N_14948);
nor UO_879 (O_879,N_14731,N_14897);
nor UO_880 (O_880,N_14868,N_14718);
nor UO_881 (O_881,N_14894,N_14744);
xor UO_882 (O_882,N_14907,N_14664);
nor UO_883 (O_883,N_14972,N_14561);
xor UO_884 (O_884,N_14916,N_14782);
nand UO_885 (O_885,N_14645,N_14889);
or UO_886 (O_886,N_14849,N_14783);
and UO_887 (O_887,N_14547,N_14653);
nor UO_888 (O_888,N_14783,N_14991);
and UO_889 (O_889,N_14961,N_14600);
or UO_890 (O_890,N_14790,N_14576);
xor UO_891 (O_891,N_14506,N_14613);
nand UO_892 (O_892,N_14902,N_14750);
nor UO_893 (O_893,N_14518,N_14815);
nor UO_894 (O_894,N_14932,N_14661);
nand UO_895 (O_895,N_14540,N_14796);
xnor UO_896 (O_896,N_14880,N_14986);
or UO_897 (O_897,N_14799,N_14836);
or UO_898 (O_898,N_14867,N_14770);
xnor UO_899 (O_899,N_14947,N_14698);
and UO_900 (O_900,N_14734,N_14607);
xor UO_901 (O_901,N_14909,N_14882);
xor UO_902 (O_902,N_14910,N_14713);
nor UO_903 (O_903,N_14511,N_14826);
or UO_904 (O_904,N_14827,N_14657);
and UO_905 (O_905,N_14570,N_14679);
nor UO_906 (O_906,N_14820,N_14617);
nand UO_907 (O_907,N_14572,N_14933);
nand UO_908 (O_908,N_14694,N_14874);
xor UO_909 (O_909,N_14997,N_14789);
nand UO_910 (O_910,N_14725,N_14937);
nor UO_911 (O_911,N_14579,N_14886);
or UO_912 (O_912,N_14566,N_14752);
nand UO_913 (O_913,N_14871,N_14813);
or UO_914 (O_914,N_14508,N_14847);
and UO_915 (O_915,N_14511,N_14813);
or UO_916 (O_916,N_14550,N_14540);
nand UO_917 (O_917,N_14574,N_14968);
or UO_918 (O_918,N_14599,N_14728);
nand UO_919 (O_919,N_14800,N_14576);
or UO_920 (O_920,N_14595,N_14852);
and UO_921 (O_921,N_14613,N_14611);
nor UO_922 (O_922,N_14567,N_14665);
nand UO_923 (O_923,N_14963,N_14665);
xnor UO_924 (O_924,N_14643,N_14747);
nor UO_925 (O_925,N_14544,N_14737);
and UO_926 (O_926,N_14679,N_14836);
xnor UO_927 (O_927,N_14532,N_14790);
xor UO_928 (O_928,N_14750,N_14687);
or UO_929 (O_929,N_14957,N_14862);
xor UO_930 (O_930,N_14621,N_14937);
or UO_931 (O_931,N_14762,N_14781);
xor UO_932 (O_932,N_14742,N_14797);
nand UO_933 (O_933,N_14664,N_14649);
or UO_934 (O_934,N_14892,N_14668);
nor UO_935 (O_935,N_14677,N_14947);
nand UO_936 (O_936,N_14867,N_14559);
or UO_937 (O_937,N_14790,N_14787);
and UO_938 (O_938,N_14974,N_14784);
or UO_939 (O_939,N_14757,N_14592);
and UO_940 (O_940,N_14621,N_14786);
nor UO_941 (O_941,N_14768,N_14605);
and UO_942 (O_942,N_14904,N_14679);
xnor UO_943 (O_943,N_14779,N_14814);
nand UO_944 (O_944,N_14769,N_14755);
nor UO_945 (O_945,N_14625,N_14635);
xor UO_946 (O_946,N_14704,N_14572);
nor UO_947 (O_947,N_14638,N_14939);
nor UO_948 (O_948,N_14897,N_14523);
xnor UO_949 (O_949,N_14766,N_14914);
or UO_950 (O_950,N_14817,N_14654);
xor UO_951 (O_951,N_14615,N_14928);
and UO_952 (O_952,N_14815,N_14600);
nand UO_953 (O_953,N_14871,N_14883);
xor UO_954 (O_954,N_14986,N_14564);
xnor UO_955 (O_955,N_14641,N_14584);
xnor UO_956 (O_956,N_14632,N_14664);
nand UO_957 (O_957,N_14694,N_14973);
and UO_958 (O_958,N_14745,N_14591);
and UO_959 (O_959,N_14585,N_14600);
and UO_960 (O_960,N_14786,N_14689);
nor UO_961 (O_961,N_14545,N_14979);
nand UO_962 (O_962,N_14788,N_14554);
nand UO_963 (O_963,N_14912,N_14569);
nand UO_964 (O_964,N_14580,N_14506);
nand UO_965 (O_965,N_14961,N_14727);
nand UO_966 (O_966,N_14571,N_14897);
and UO_967 (O_967,N_14865,N_14814);
and UO_968 (O_968,N_14878,N_14708);
nand UO_969 (O_969,N_14582,N_14641);
xnor UO_970 (O_970,N_14911,N_14511);
nand UO_971 (O_971,N_14925,N_14683);
xnor UO_972 (O_972,N_14907,N_14737);
and UO_973 (O_973,N_14934,N_14989);
nor UO_974 (O_974,N_14538,N_14714);
nor UO_975 (O_975,N_14578,N_14693);
and UO_976 (O_976,N_14575,N_14818);
nor UO_977 (O_977,N_14952,N_14903);
nor UO_978 (O_978,N_14762,N_14592);
xnor UO_979 (O_979,N_14767,N_14921);
nor UO_980 (O_980,N_14769,N_14810);
nand UO_981 (O_981,N_14974,N_14585);
nand UO_982 (O_982,N_14937,N_14601);
nor UO_983 (O_983,N_14514,N_14678);
or UO_984 (O_984,N_14934,N_14508);
nor UO_985 (O_985,N_14692,N_14939);
nor UO_986 (O_986,N_14738,N_14671);
xor UO_987 (O_987,N_14607,N_14667);
nor UO_988 (O_988,N_14962,N_14596);
xor UO_989 (O_989,N_14949,N_14589);
nor UO_990 (O_990,N_14603,N_14857);
nand UO_991 (O_991,N_14623,N_14511);
nor UO_992 (O_992,N_14510,N_14956);
xor UO_993 (O_993,N_14726,N_14682);
and UO_994 (O_994,N_14760,N_14851);
nand UO_995 (O_995,N_14623,N_14828);
nor UO_996 (O_996,N_14898,N_14690);
nor UO_997 (O_997,N_14558,N_14960);
nor UO_998 (O_998,N_14983,N_14764);
and UO_999 (O_999,N_14722,N_14826);
xor UO_1000 (O_1000,N_14854,N_14739);
nand UO_1001 (O_1001,N_14768,N_14818);
and UO_1002 (O_1002,N_14801,N_14536);
nor UO_1003 (O_1003,N_14773,N_14745);
xor UO_1004 (O_1004,N_14657,N_14869);
or UO_1005 (O_1005,N_14945,N_14704);
and UO_1006 (O_1006,N_14685,N_14611);
or UO_1007 (O_1007,N_14522,N_14505);
xor UO_1008 (O_1008,N_14674,N_14925);
or UO_1009 (O_1009,N_14652,N_14513);
xor UO_1010 (O_1010,N_14537,N_14844);
xor UO_1011 (O_1011,N_14660,N_14785);
and UO_1012 (O_1012,N_14849,N_14612);
nand UO_1013 (O_1013,N_14964,N_14909);
xnor UO_1014 (O_1014,N_14780,N_14661);
xor UO_1015 (O_1015,N_14873,N_14965);
or UO_1016 (O_1016,N_14814,N_14610);
and UO_1017 (O_1017,N_14919,N_14827);
nand UO_1018 (O_1018,N_14842,N_14711);
xnor UO_1019 (O_1019,N_14825,N_14659);
and UO_1020 (O_1020,N_14530,N_14743);
and UO_1021 (O_1021,N_14779,N_14600);
nand UO_1022 (O_1022,N_14950,N_14663);
xor UO_1023 (O_1023,N_14681,N_14536);
xor UO_1024 (O_1024,N_14768,N_14637);
xnor UO_1025 (O_1025,N_14644,N_14505);
and UO_1026 (O_1026,N_14547,N_14748);
or UO_1027 (O_1027,N_14885,N_14822);
or UO_1028 (O_1028,N_14776,N_14780);
xor UO_1029 (O_1029,N_14527,N_14646);
nor UO_1030 (O_1030,N_14708,N_14523);
or UO_1031 (O_1031,N_14607,N_14699);
nand UO_1032 (O_1032,N_14877,N_14967);
xor UO_1033 (O_1033,N_14909,N_14918);
nor UO_1034 (O_1034,N_14624,N_14567);
or UO_1035 (O_1035,N_14564,N_14796);
xor UO_1036 (O_1036,N_14661,N_14904);
nand UO_1037 (O_1037,N_14862,N_14566);
or UO_1038 (O_1038,N_14965,N_14563);
or UO_1039 (O_1039,N_14644,N_14786);
and UO_1040 (O_1040,N_14833,N_14750);
or UO_1041 (O_1041,N_14623,N_14947);
nor UO_1042 (O_1042,N_14845,N_14940);
nor UO_1043 (O_1043,N_14685,N_14698);
or UO_1044 (O_1044,N_14503,N_14505);
and UO_1045 (O_1045,N_14507,N_14649);
nor UO_1046 (O_1046,N_14589,N_14763);
nand UO_1047 (O_1047,N_14957,N_14632);
and UO_1048 (O_1048,N_14564,N_14787);
or UO_1049 (O_1049,N_14640,N_14796);
and UO_1050 (O_1050,N_14501,N_14505);
or UO_1051 (O_1051,N_14558,N_14696);
and UO_1052 (O_1052,N_14759,N_14974);
xnor UO_1053 (O_1053,N_14918,N_14883);
nor UO_1054 (O_1054,N_14803,N_14725);
xnor UO_1055 (O_1055,N_14707,N_14873);
nand UO_1056 (O_1056,N_14729,N_14780);
nor UO_1057 (O_1057,N_14930,N_14920);
or UO_1058 (O_1058,N_14772,N_14779);
nor UO_1059 (O_1059,N_14678,N_14663);
xor UO_1060 (O_1060,N_14611,N_14684);
xnor UO_1061 (O_1061,N_14808,N_14516);
xnor UO_1062 (O_1062,N_14721,N_14626);
nand UO_1063 (O_1063,N_14642,N_14712);
and UO_1064 (O_1064,N_14537,N_14772);
nor UO_1065 (O_1065,N_14630,N_14581);
or UO_1066 (O_1066,N_14976,N_14787);
and UO_1067 (O_1067,N_14851,N_14535);
and UO_1068 (O_1068,N_14745,N_14935);
xor UO_1069 (O_1069,N_14954,N_14597);
nand UO_1070 (O_1070,N_14967,N_14592);
xnor UO_1071 (O_1071,N_14994,N_14726);
nand UO_1072 (O_1072,N_14779,N_14972);
nor UO_1073 (O_1073,N_14737,N_14993);
and UO_1074 (O_1074,N_14727,N_14801);
and UO_1075 (O_1075,N_14986,N_14534);
nand UO_1076 (O_1076,N_14633,N_14618);
or UO_1077 (O_1077,N_14547,N_14934);
xnor UO_1078 (O_1078,N_14910,N_14760);
nor UO_1079 (O_1079,N_14617,N_14761);
xnor UO_1080 (O_1080,N_14982,N_14641);
xnor UO_1081 (O_1081,N_14684,N_14834);
nand UO_1082 (O_1082,N_14811,N_14725);
or UO_1083 (O_1083,N_14744,N_14760);
nor UO_1084 (O_1084,N_14500,N_14518);
or UO_1085 (O_1085,N_14682,N_14501);
or UO_1086 (O_1086,N_14538,N_14622);
xnor UO_1087 (O_1087,N_14772,N_14909);
xor UO_1088 (O_1088,N_14967,N_14879);
nor UO_1089 (O_1089,N_14972,N_14689);
xor UO_1090 (O_1090,N_14559,N_14836);
or UO_1091 (O_1091,N_14848,N_14989);
nor UO_1092 (O_1092,N_14725,N_14734);
xnor UO_1093 (O_1093,N_14836,N_14761);
or UO_1094 (O_1094,N_14925,N_14570);
and UO_1095 (O_1095,N_14955,N_14671);
xor UO_1096 (O_1096,N_14788,N_14766);
xnor UO_1097 (O_1097,N_14937,N_14516);
and UO_1098 (O_1098,N_14857,N_14898);
xnor UO_1099 (O_1099,N_14725,N_14652);
nor UO_1100 (O_1100,N_14627,N_14855);
xor UO_1101 (O_1101,N_14730,N_14971);
and UO_1102 (O_1102,N_14647,N_14654);
and UO_1103 (O_1103,N_14647,N_14630);
nand UO_1104 (O_1104,N_14507,N_14789);
nor UO_1105 (O_1105,N_14950,N_14871);
or UO_1106 (O_1106,N_14637,N_14892);
and UO_1107 (O_1107,N_14974,N_14833);
and UO_1108 (O_1108,N_14597,N_14536);
or UO_1109 (O_1109,N_14786,N_14835);
and UO_1110 (O_1110,N_14804,N_14529);
nand UO_1111 (O_1111,N_14964,N_14864);
nand UO_1112 (O_1112,N_14991,N_14589);
xnor UO_1113 (O_1113,N_14546,N_14961);
and UO_1114 (O_1114,N_14510,N_14903);
xor UO_1115 (O_1115,N_14793,N_14912);
xor UO_1116 (O_1116,N_14899,N_14600);
or UO_1117 (O_1117,N_14700,N_14821);
nand UO_1118 (O_1118,N_14775,N_14746);
or UO_1119 (O_1119,N_14508,N_14781);
or UO_1120 (O_1120,N_14988,N_14705);
xnor UO_1121 (O_1121,N_14796,N_14707);
or UO_1122 (O_1122,N_14717,N_14934);
nand UO_1123 (O_1123,N_14704,N_14802);
xor UO_1124 (O_1124,N_14718,N_14658);
nor UO_1125 (O_1125,N_14709,N_14995);
and UO_1126 (O_1126,N_14978,N_14979);
xnor UO_1127 (O_1127,N_14513,N_14740);
nand UO_1128 (O_1128,N_14539,N_14861);
nand UO_1129 (O_1129,N_14669,N_14543);
xor UO_1130 (O_1130,N_14819,N_14822);
xnor UO_1131 (O_1131,N_14706,N_14693);
or UO_1132 (O_1132,N_14969,N_14749);
xor UO_1133 (O_1133,N_14783,N_14979);
nand UO_1134 (O_1134,N_14516,N_14973);
and UO_1135 (O_1135,N_14583,N_14735);
nor UO_1136 (O_1136,N_14866,N_14660);
nor UO_1137 (O_1137,N_14826,N_14639);
xor UO_1138 (O_1138,N_14608,N_14517);
nor UO_1139 (O_1139,N_14868,N_14971);
and UO_1140 (O_1140,N_14575,N_14714);
and UO_1141 (O_1141,N_14539,N_14639);
xor UO_1142 (O_1142,N_14693,N_14546);
xnor UO_1143 (O_1143,N_14680,N_14560);
and UO_1144 (O_1144,N_14979,N_14528);
nor UO_1145 (O_1145,N_14907,N_14695);
or UO_1146 (O_1146,N_14873,N_14674);
nor UO_1147 (O_1147,N_14599,N_14894);
nand UO_1148 (O_1148,N_14993,N_14772);
and UO_1149 (O_1149,N_14952,N_14818);
and UO_1150 (O_1150,N_14697,N_14776);
xor UO_1151 (O_1151,N_14924,N_14911);
or UO_1152 (O_1152,N_14880,N_14658);
or UO_1153 (O_1153,N_14936,N_14644);
nor UO_1154 (O_1154,N_14849,N_14795);
or UO_1155 (O_1155,N_14518,N_14977);
or UO_1156 (O_1156,N_14694,N_14648);
xor UO_1157 (O_1157,N_14522,N_14849);
nor UO_1158 (O_1158,N_14930,N_14749);
or UO_1159 (O_1159,N_14988,N_14902);
nor UO_1160 (O_1160,N_14826,N_14663);
and UO_1161 (O_1161,N_14896,N_14755);
nor UO_1162 (O_1162,N_14632,N_14509);
xnor UO_1163 (O_1163,N_14500,N_14784);
xnor UO_1164 (O_1164,N_14923,N_14600);
or UO_1165 (O_1165,N_14594,N_14666);
xor UO_1166 (O_1166,N_14656,N_14552);
or UO_1167 (O_1167,N_14708,N_14727);
nand UO_1168 (O_1168,N_14678,N_14542);
xnor UO_1169 (O_1169,N_14892,N_14595);
xor UO_1170 (O_1170,N_14531,N_14879);
or UO_1171 (O_1171,N_14532,N_14751);
nand UO_1172 (O_1172,N_14524,N_14507);
or UO_1173 (O_1173,N_14544,N_14668);
and UO_1174 (O_1174,N_14964,N_14918);
or UO_1175 (O_1175,N_14729,N_14978);
nand UO_1176 (O_1176,N_14605,N_14666);
nand UO_1177 (O_1177,N_14762,N_14822);
and UO_1178 (O_1178,N_14796,N_14794);
nand UO_1179 (O_1179,N_14590,N_14928);
nor UO_1180 (O_1180,N_14808,N_14600);
nand UO_1181 (O_1181,N_14938,N_14916);
and UO_1182 (O_1182,N_14848,N_14608);
xnor UO_1183 (O_1183,N_14877,N_14714);
and UO_1184 (O_1184,N_14745,N_14641);
nor UO_1185 (O_1185,N_14607,N_14516);
xnor UO_1186 (O_1186,N_14577,N_14977);
nand UO_1187 (O_1187,N_14578,N_14883);
or UO_1188 (O_1188,N_14881,N_14960);
or UO_1189 (O_1189,N_14650,N_14609);
nor UO_1190 (O_1190,N_14864,N_14551);
xor UO_1191 (O_1191,N_14557,N_14893);
nand UO_1192 (O_1192,N_14869,N_14611);
or UO_1193 (O_1193,N_14999,N_14922);
nand UO_1194 (O_1194,N_14645,N_14778);
xor UO_1195 (O_1195,N_14599,N_14882);
nand UO_1196 (O_1196,N_14663,N_14869);
and UO_1197 (O_1197,N_14912,N_14770);
nor UO_1198 (O_1198,N_14533,N_14705);
xnor UO_1199 (O_1199,N_14929,N_14595);
nor UO_1200 (O_1200,N_14791,N_14549);
xor UO_1201 (O_1201,N_14717,N_14628);
nand UO_1202 (O_1202,N_14837,N_14993);
or UO_1203 (O_1203,N_14942,N_14603);
and UO_1204 (O_1204,N_14912,N_14874);
and UO_1205 (O_1205,N_14628,N_14735);
and UO_1206 (O_1206,N_14880,N_14739);
nand UO_1207 (O_1207,N_14531,N_14596);
nor UO_1208 (O_1208,N_14559,N_14902);
nor UO_1209 (O_1209,N_14592,N_14770);
nor UO_1210 (O_1210,N_14984,N_14986);
nor UO_1211 (O_1211,N_14570,N_14651);
and UO_1212 (O_1212,N_14732,N_14667);
and UO_1213 (O_1213,N_14729,N_14894);
xor UO_1214 (O_1214,N_14609,N_14710);
xor UO_1215 (O_1215,N_14691,N_14696);
nand UO_1216 (O_1216,N_14895,N_14970);
nor UO_1217 (O_1217,N_14966,N_14588);
and UO_1218 (O_1218,N_14866,N_14699);
and UO_1219 (O_1219,N_14964,N_14947);
xor UO_1220 (O_1220,N_14935,N_14861);
xor UO_1221 (O_1221,N_14847,N_14639);
nand UO_1222 (O_1222,N_14677,N_14749);
or UO_1223 (O_1223,N_14591,N_14908);
or UO_1224 (O_1224,N_14755,N_14926);
xor UO_1225 (O_1225,N_14607,N_14836);
xor UO_1226 (O_1226,N_14940,N_14787);
nand UO_1227 (O_1227,N_14794,N_14755);
xor UO_1228 (O_1228,N_14746,N_14783);
and UO_1229 (O_1229,N_14824,N_14898);
and UO_1230 (O_1230,N_14638,N_14803);
and UO_1231 (O_1231,N_14560,N_14988);
nor UO_1232 (O_1232,N_14962,N_14831);
and UO_1233 (O_1233,N_14814,N_14529);
nor UO_1234 (O_1234,N_14776,N_14827);
or UO_1235 (O_1235,N_14707,N_14880);
nand UO_1236 (O_1236,N_14742,N_14926);
nand UO_1237 (O_1237,N_14763,N_14674);
nor UO_1238 (O_1238,N_14948,N_14940);
nand UO_1239 (O_1239,N_14738,N_14974);
nand UO_1240 (O_1240,N_14874,N_14867);
xnor UO_1241 (O_1241,N_14934,N_14775);
and UO_1242 (O_1242,N_14637,N_14781);
nand UO_1243 (O_1243,N_14531,N_14530);
xor UO_1244 (O_1244,N_14679,N_14692);
nand UO_1245 (O_1245,N_14566,N_14573);
or UO_1246 (O_1246,N_14666,N_14976);
nor UO_1247 (O_1247,N_14635,N_14743);
nand UO_1248 (O_1248,N_14506,N_14996);
nand UO_1249 (O_1249,N_14618,N_14865);
nand UO_1250 (O_1250,N_14617,N_14626);
xnor UO_1251 (O_1251,N_14800,N_14679);
nor UO_1252 (O_1252,N_14755,N_14580);
and UO_1253 (O_1253,N_14596,N_14757);
or UO_1254 (O_1254,N_14862,N_14525);
nor UO_1255 (O_1255,N_14720,N_14749);
nand UO_1256 (O_1256,N_14741,N_14923);
or UO_1257 (O_1257,N_14733,N_14611);
nand UO_1258 (O_1258,N_14548,N_14957);
or UO_1259 (O_1259,N_14696,N_14571);
and UO_1260 (O_1260,N_14583,N_14819);
xnor UO_1261 (O_1261,N_14539,N_14563);
nor UO_1262 (O_1262,N_14537,N_14648);
and UO_1263 (O_1263,N_14823,N_14607);
nor UO_1264 (O_1264,N_14789,N_14636);
xnor UO_1265 (O_1265,N_14611,N_14887);
nand UO_1266 (O_1266,N_14852,N_14836);
and UO_1267 (O_1267,N_14843,N_14903);
nor UO_1268 (O_1268,N_14989,N_14576);
nor UO_1269 (O_1269,N_14725,N_14801);
or UO_1270 (O_1270,N_14837,N_14819);
or UO_1271 (O_1271,N_14510,N_14695);
and UO_1272 (O_1272,N_14929,N_14860);
nor UO_1273 (O_1273,N_14589,N_14686);
nand UO_1274 (O_1274,N_14546,N_14536);
xor UO_1275 (O_1275,N_14626,N_14858);
nor UO_1276 (O_1276,N_14821,N_14763);
nand UO_1277 (O_1277,N_14627,N_14962);
nor UO_1278 (O_1278,N_14706,N_14697);
xor UO_1279 (O_1279,N_14954,N_14603);
and UO_1280 (O_1280,N_14625,N_14751);
xor UO_1281 (O_1281,N_14533,N_14854);
and UO_1282 (O_1282,N_14880,N_14909);
nor UO_1283 (O_1283,N_14697,N_14699);
nor UO_1284 (O_1284,N_14703,N_14723);
or UO_1285 (O_1285,N_14568,N_14614);
xor UO_1286 (O_1286,N_14640,N_14762);
xor UO_1287 (O_1287,N_14550,N_14707);
nor UO_1288 (O_1288,N_14961,N_14942);
or UO_1289 (O_1289,N_14754,N_14887);
xor UO_1290 (O_1290,N_14745,N_14687);
nor UO_1291 (O_1291,N_14547,N_14758);
nor UO_1292 (O_1292,N_14548,N_14628);
or UO_1293 (O_1293,N_14664,N_14668);
nand UO_1294 (O_1294,N_14998,N_14952);
xor UO_1295 (O_1295,N_14617,N_14665);
and UO_1296 (O_1296,N_14702,N_14794);
and UO_1297 (O_1297,N_14835,N_14555);
xor UO_1298 (O_1298,N_14866,N_14590);
or UO_1299 (O_1299,N_14650,N_14552);
nand UO_1300 (O_1300,N_14838,N_14900);
nor UO_1301 (O_1301,N_14847,N_14821);
xor UO_1302 (O_1302,N_14578,N_14728);
xor UO_1303 (O_1303,N_14834,N_14825);
and UO_1304 (O_1304,N_14884,N_14904);
and UO_1305 (O_1305,N_14718,N_14919);
xor UO_1306 (O_1306,N_14954,N_14859);
xor UO_1307 (O_1307,N_14772,N_14676);
and UO_1308 (O_1308,N_14520,N_14806);
or UO_1309 (O_1309,N_14810,N_14563);
nor UO_1310 (O_1310,N_14853,N_14832);
nand UO_1311 (O_1311,N_14936,N_14579);
or UO_1312 (O_1312,N_14767,N_14862);
nand UO_1313 (O_1313,N_14905,N_14503);
and UO_1314 (O_1314,N_14752,N_14913);
nor UO_1315 (O_1315,N_14896,N_14763);
and UO_1316 (O_1316,N_14825,N_14974);
xor UO_1317 (O_1317,N_14993,N_14834);
xnor UO_1318 (O_1318,N_14782,N_14977);
xor UO_1319 (O_1319,N_14777,N_14801);
nor UO_1320 (O_1320,N_14792,N_14669);
nand UO_1321 (O_1321,N_14655,N_14633);
or UO_1322 (O_1322,N_14666,N_14664);
nor UO_1323 (O_1323,N_14556,N_14662);
and UO_1324 (O_1324,N_14690,N_14864);
nor UO_1325 (O_1325,N_14603,N_14811);
nor UO_1326 (O_1326,N_14857,N_14694);
nand UO_1327 (O_1327,N_14626,N_14533);
nor UO_1328 (O_1328,N_14730,N_14853);
nand UO_1329 (O_1329,N_14839,N_14853);
nand UO_1330 (O_1330,N_14903,N_14568);
nand UO_1331 (O_1331,N_14606,N_14971);
xnor UO_1332 (O_1332,N_14944,N_14815);
or UO_1333 (O_1333,N_14693,N_14927);
xor UO_1334 (O_1334,N_14649,N_14968);
xor UO_1335 (O_1335,N_14678,N_14988);
nor UO_1336 (O_1336,N_14556,N_14574);
or UO_1337 (O_1337,N_14728,N_14662);
nor UO_1338 (O_1338,N_14949,N_14504);
and UO_1339 (O_1339,N_14557,N_14925);
xor UO_1340 (O_1340,N_14817,N_14627);
and UO_1341 (O_1341,N_14684,N_14773);
nor UO_1342 (O_1342,N_14948,N_14944);
nor UO_1343 (O_1343,N_14527,N_14726);
or UO_1344 (O_1344,N_14851,N_14882);
or UO_1345 (O_1345,N_14851,N_14593);
or UO_1346 (O_1346,N_14928,N_14903);
xnor UO_1347 (O_1347,N_14915,N_14739);
nor UO_1348 (O_1348,N_14539,N_14677);
or UO_1349 (O_1349,N_14891,N_14709);
xor UO_1350 (O_1350,N_14965,N_14829);
xor UO_1351 (O_1351,N_14745,N_14713);
or UO_1352 (O_1352,N_14679,N_14838);
nor UO_1353 (O_1353,N_14877,N_14652);
xor UO_1354 (O_1354,N_14992,N_14978);
or UO_1355 (O_1355,N_14706,N_14677);
nor UO_1356 (O_1356,N_14698,N_14538);
nor UO_1357 (O_1357,N_14550,N_14826);
or UO_1358 (O_1358,N_14718,N_14520);
xor UO_1359 (O_1359,N_14634,N_14892);
or UO_1360 (O_1360,N_14567,N_14692);
nor UO_1361 (O_1361,N_14671,N_14506);
nand UO_1362 (O_1362,N_14904,N_14922);
and UO_1363 (O_1363,N_14859,N_14616);
nand UO_1364 (O_1364,N_14735,N_14986);
nand UO_1365 (O_1365,N_14832,N_14882);
xnor UO_1366 (O_1366,N_14593,N_14949);
or UO_1367 (O_1367,N_14975,N_14909);
xnor UO_1368 (O_1368,N_14770,N_14517);
nand UO_1369 (O_1369,N_14798,N_14835);
or UO_1370 (O_1370,N_14787,N_14671);
nor UO_1371 (O_1371,N_14706,N_14676);
xor UO_1372 (O_1372,N_14653,N_14801);
xnor UO_1373 (O_1373,N_14861,N_14809);
nor UO_1374 (O_1374,N_14632,N_14521);
nor UO_1375 (O_1375,N_14623,N_14850);
nor UO_1376 (O_1376,N_14676,N_14542);
nand UO_1377 (O_1377,N_14758,N_14649);
and UO_1378 (O_1378,N_14809,N_14647);
nand UO_1379 (O_1379,N_14519,N_14991);
nor UO_1380 (O_1380,N_14944,N_14548);
or UO_1381 (O_1381,N_14536,N_14947);
or UO_1382 (O_1382,N_14873,N_14878);
nor UO_1383 (O_1383,N_14584,N_14629);
nand UO_1384 (O_1384,N_14624,N_14758);
nand UO_1385 (O_1385,N_14515,N_14930);
or UO_1386 (O_1386,N_14994,N_14968);
or UO_1387 (O_1387,N_14542,N_14556);
and UO_1388 (O_1388,N_14514,N_14831);
or UO_1389 (O_1389,N_14808,N_14964);
xor UO_1390 (O_1390,N_14540,N_14927);
xor UO_1391 (O_1391,N_14574,N_14750);
nand UO_1392 (O_1392,N_14585,N_14845);
nand UO_1393 (O_1393,N_14977,N_14630);
xor UO_1394 (O_1394,N_14881,N_14569);
xor UO_1395 (O_1395,N_14983,N_14839);
and UO_1396 (O_1396,N_14724,N_14541);
and UO_1397 (O_1397,N_14820,N_14806);
nor UO_1398 (O_1398,N_14515,N_14607);
and UO_1399 (O_1399,N_14846,N_14651);
nor UO_1400 (O_1400,N_14712,N_14791);
or UO_1401 (O_1401,N_14716,N_14625);
nand UO_1402 (O_1402,N_14914,N_14922);
nand UO_1403 (O_1403,N_14566,N_14744);
and UO_1404 (O_1404,N_14605,N_14882);
nor UO_1405 (O_1405,N_14609,N_14719);
or UO_1406 (O_1406,N_14705,N_14584);
nand UO_1407 (O_1407,N_14885,N_14833);
nor UO_1408 (O_1408,N_14532,N_14850);
or UO_1409 (O_1409,N_14952,N_14890);
nor UO_1410 (O_1410,N_14996,N_14655);
nor UO_1411 (O_1411,N_14614,N_14941);
nand UO_1412 (O_1412,N_14998,N_14902);
and UO_1413 (O_1413,N_14683,N_14633);
xor UO_1414 (O_1414,N_14578,N_14803);
xnor UO_1415 (O_1415,N_14575,N_14960);
and UO_1416 (O_1416,N_14964,N_14651);
or UO_1417 (O_1417,N_14542,N_14715);
or UO_1418 (O_1418,N_14655,N_14691);
or UO_1419 (O_1419,N_14734,N_14880);
or UO_1420 (O_1420,N_14607,N_14631);
nor UO_1421 (O_1421,N_14830,N_14766);
and UO_1422 (O_1422,N_14520,N_14823);
nand UO_1423 (O_1423,N_14920,N_14733);
xnor UO_1424 (O_1424,N_14692,N_14728);
or UO_1425 (O_1425,N_14733,N_14863);
or UO_1426 (O_1426,N_14877,N_14827);
nor UO_1427 (O_1427,N_14505,N_14938);
or UO_1428 (O_1428,N_14504,N_14636);
xnor UO_1429 (O_1429,N_14737,N_14947);
nand UO_1430 (O_1430,N_14688,N_14575);
nor UO_1431 (O_1431,N_14655,N_14853);
or UO_1432 (O_1432,N_14875,N_14741);
nor UO_1433 (O_1433,N_14672,N_14938);
xor UO_1434 (O_1434,N_14893,N_14762);
nor UO_1435 (O_1435,N_14592,N_14746);
nor UO_1436 (O_1436,N_14909,N_14755);
nand UO_1437 (O_1437,N_14841,N_14926);
nand UO_1438 (O_1438,N_14845,N_14719);
and UO_1439 (O_1439,N_14800,N_14649);
nor UO_1440 (O_1440,N_14652,N_14761);
nand UO_1441 (O_1441,N_14766,N_14509);
or UO_1442 (O_1442,N_14851,N_14735);
or UO_1443 (O_1443,N_14687,N_14787);
and UO_1444 (O_1444,N_14518,N_14916);
nor UO_1445 (O_1445,N_14766,N_14746);
nor UO_1446 (O_1446,N_14529,N_14750);
or UO_1447 (O_1447,N_14557,N_14711);
nand UO_1448 (O_1448,N_14529,N_14799);
xor UO_1449 (O_1449,N_14531,N_14868);
and UO_1450 (O_1450,N_14873,N_14682);
xnor UO_1451 (O_1451,N_14880,N_14802);
and UO_1452 (O_1452,N_14856,N_14880);
xor UO_1453 (O_1453,N_14890,N_14659);
nand UO_1454 (O_1454,N_14828,N_14990);
nor UO_1455 (O_1455,N_14884,N_14774);
nand UO_1456 (O_1456,N_14952,N_14689);
xor UO_1457 (O_1457,N_14672,N_14778);
nor UO_1458 (O_1458,N_14606,N_14615);
and UO_1459 (O_1459,N_14873,N_14625);
and UO_1460 (O_1460,N_14953,N_14608);
xor UO_1461 (O_1461,N_14992,N_14751);
nor UO_1462 (O_1462,N_14795,N_14685);
nand UO_1463 (O_1463,N_14793,N_14722);
nand UO_1464 (O_1464,N_14534,N_14982);
nor UO_1465 (O_1465,N_14664,N_14540);
and UO_1466 (O_1466,N_14982,N_14950);
nand UO_1467 (O_1467,N_14647,N_14680);
nor UO_1468 (O_1468,N_14790,N_14896);
xor UO_1469 (O_1469,N_14956,N_14886);
xor UO_1470 (O_1470,N_14571,N_14744);
nor UO_1471 (O_1471,N_14660,N_14786);
nand UO_1472 (O_1472,N_14728,N_14852);
xor UO_1473 (O_1473,N_14606,N_14625);
nand UO_1474 (O_1474,N_14727,N_14772);
nor UO_1475 (O_1475,N_14508,N_14551);
nand UO_1476 (O_1476,N_14677,N_14615);
or UO_1477 (O_1477,N_14949,N_14716);
or UO_1478 (O_1478,N_14514,N_14722);
and UO_1479 (O_1479,N_14537,N_14840);
or UO_1480 (O_1480,N_14623,N_14790);
xor UO_1481 (O_1481,N_14691,N_14904);
xor UO_1482 (O_1482,N_14719,N_14738);
and UO_1483 (O_1483,N_14954,N_14915);
nor UO_1484 (O_1484,N_14576,N_14620);
and UO_1485 (O_1485,N_14651,N_14626);
nor UO_1486 (O_1486,N_14781,N_14666);
nand UO_1487 (O_1487,N_14564,N_14596);
nor UO_1488 (O_1488,N_14944,N_14709);
xnor UO_1489 (O_1489,N_14902,N_14518);
or UO_1490 (O_1490,N_14579,N_14670);
nor UO_1491 (O_1491,N_14998,N_14873);
xnor UO_1492 (O_1492,N_14520,N_14559);
nor UO_1493 (O_1493,N_14502,N_14791);
and UO_1494 (O_1494,N_14799,N_14730);
and UO_1495 (O_1495,N_14807,N_14911);
or UO_1496 (O_1496,N_14649,N_14939);
nor UO_1497 (O_1497,N_14915,N_14704);
and UO_1498 (O_1498,N_14736,N_14582);
nand UO_1499 (O_1499,N_14554,N_14606);
and UO_1500 (O_1500,N_14554,N_14960);
xnor UO_1501 (O_1501,N_14771,N_14877);
xnor UO_1502 (O_1502,N_14811,N_14572);
or UO_1503 (O_1503,N_14649,N_14655);
xor UO_1504 (O_1504,N_14867,N_14791);
or UO_1505 (O_1505,N_14840,N_14812);
nand UO_1506 (O_1506,N_14576,N_14637);
and UO_1507 (O_1507,N_14551,N_14667);
nor UO_1508 (O_1508,N_14607,N_14878);
and UO_1509 (O_1509,N_14603,N_14934);
xnor UO_1510 (O_1510,N_14950,N_14592);
or UO_1511 (O_1511,N_14815,N_14701);
or UO_1512 (O_1512,N_14762,N_14800);
or UO_1513 (O_1513,N_14891,N_14719);
nor UO_1514 (O_1514,N_14578,N_14817);
nand UO_1515 (O_1515,N_14962,N_14850);
or UO_1516 (O_1516,N_14850,N_14781);
xor UO_1517 (O_1517,N_14575,N_14614);
nor UO_1518 (O_1518,N_14718,N_14677);
or UO_1519 (O_1519,N_14641,N_14865);
xor UO_1520 (O_1520,N_14527,N_14985);
or UO_1521 (O_1521,N_14567,N_14632);
xnor UO_1522 (O_1522,N_14656,N_14951);
nor UO_1523 (O_1523,N_14784,N_14782);
xor UO_1524 (O_1524,N_14688,N_14787);
nor UO_1525 (O_1525,N_14887,N_14840);
xor UO_1526 (O_1526,N_14662,N_14782);
or UO_1527 (O_1527,N_14969,N_14904);
xnor UO_1528 (O_1528,N_14991,N_14906);
and UO_1529 (O_1529,N_14966,N_14781);
or UO_1530 (O_1530,N_14746,N_14638);
nand UO_1531 (O_1531,N_14967,N_14544);
nand UO_1532 (O_1532,N_14636,N_14805);
xor UO_1533 (O_1533,N_14828,N_14505);
nand UO_1534 (O_1534,N_14901,N_14711);
xor UO_1535 (O_1535,N_14748,N_14855);
nor UO_1536 (O_1536,N_14684,N_14928);
or UO_1537 (O_1537,N_14863,N_14901);
nand UO_1538 (O_1538,N_14964,N_14756);
nor UO_1539 (O_1539,N_14549,N_14732);
xnor UO_1540 (O_1540,N_14668,N_14941);
xnor UO_1541 (O_1541,N_14847,N_14980);
and UO_1542 (O_1542,N_14908,N_14798);
nor UO_1543 (O_1543,N_14818,N_14577);
or UO_1544 (O_1544,N_14502,N_14731);
or UO_1545 (O_1545,N_14762,N_14519);
nor UO_1546 (O_1546,N_14862,N_14868);
xor UO_1547 (O_1547,N_14832,N_14891);
and UO_1548 (O_1548,N_14553,N_14687);
or UO_1549 (O_1549,N_14543,N_14943);
or UO_1550 (O_1550,N_14847,N_14931);
xor UO_1551 (O_1551,N_14752,N_14633);
and UO_1552 (O_1552,N_14782,N_14728);
and UO_1553 (O_1553,N_14772,N_14912);
or UO_1554 (O_1554,N_14631,N_14597);
or UO_1555 (O_1555,N_14539,N_14702);
nand UO_1556 (O_1556,N_14820,N_14894);
xor UO_1557 (O_1557,N_14782,N_14791);
nor UO_1558 (O_1558,N_14842,N_14667);
nand UO_1559 (O_1559,N_14847,N_14892);
and UO_1560 (O_1560,N_14697,N_14527);
or UO_1561 (O_1561,N_14728,N_14573);
nand UO_1562 (O_1562,N_14531,N_14508);
nor UO_1563 (O_1563,N_14586,N_14820);
nand UO_1564 (O_1564,N_14510,N_14525);
or UO_1565 (O_1565,N_14819,N_14787);
xnor UO_1566 (O_1566,N_14875,N_14661);
or UO_1567 (O_1567,N_14975,N_14930);
xor UO_1568 (O_1568,N_14721,N_14762);
nand UO_1569 (O_1569,N_14511,N_14534);
xnor UO_1570 (O_1570,N_14506,N_14624);
nand UO_1571 (O_1571,N_14654,N_14593);
nor UO_1572 (O_1572,N_14853,N_14598);
xnor UO_1573 (O_1573,N_14634,N_14780);
xnor UO_1574 (O_1574,N_14838,N_14715);
and UO_1575 (O_1575,N_14911,N_14667);
nand UO_1576 (O_1576,N_14552,N_14763);
nand UO_1577 (O_1577,N_14611,N_14823);
nor UO_1578 (O_1578,N_14525,N_14645);
nor UO_1579 (O_1579,N_14817,N_14653);
and UO_1580 (O_1580,N_14705,N_14566);
and UO_1581 (O_1581,N_14747,N_14727);
nor UO_1582 (O_1582,N_14915,N_14561);
nor UO_1583 (O_1583,N_14640,N_14845);
or UO_1584 (O_1584,N_14514,N_14515);
and UO_1585 (O_1585,N_14639,N_14857);
nand UO_1586 (O_1586,N_14818,N_14981);
nand UO_1587 (O_1587,N_14944,N_14504);
nor UO_1588 (O_1588,N_14773,N_14959);
xnor UO_1589 (O_1589,N_14594,N_14625);
nor UO_1590 (O_1590,N_14569,N_14958);
nand UO_1591 (O_1591,N_14847,N_14907);
and UO_1592 (O_1592,N_14666,N_14941);
xnor UO_1593 (O_1593,N_14939,N_14507);
xnor UO_1594 (O_1594,N_14747,N_14985);
or UO_1595 (O_1595,N_14822,N_14868);
xnor UO_1596 (O_1596,N_14790,N_14702);
or UO_1597 (O_1597,N_14696,N_14598);
nor UO_1598 (O_1598,N_14841,N_14717);
nor UO_1599 (O_1599,N_14795,N_14938);
xor UO_1600 (O_1600,N_14745,N_14976);
nand UO_1601 (O_1601,N_14904,N_14540);
nor UO_1602 (O_1602,N_14879,N_14599);
nand UO_1603 (O_1603,N_14934,N_14589);
nor UO_1604 (O_1604,N_14597,N_14772);
xor UO_1605 (O_1605,N_14852,N_14739);
nor UO_1606 (O_1606,N_14823,N_14927);
and UO_1607 (O_1607,N_14766,N_14941);
xor UO_1608 (O_1608,N_14646,N_14683);
or UO_1609 (O_1609,N_14597,N_14842);
nor UO_1610 (O_1610,N_14848,N_14733);
or UO_1611 (O_1611,N_14942,N_14559);
or UO_1612 (O_1612,N_14598,N_14562);
or UO_1613 (O_1613,N_14598,N_14763);
xor UO_1614 (O_1614,N_14848,N_14627);
nor UO_1615 (O_1615,N_14561,N_14884);
and UO_1616 (O_1616,N_14909,N_14634);
or UO_1617 (O_1617,N_14840,N_14843);
or UO_1618 (O_1618,N_14630,N_14659);
nor UO_1619 (O_1619,N_14934,N_14632);
nand UO_1620 (O_1620,N_14689,N_14753);
nand UO_1621 (O_1621,N_14992,N_14526);
or UO_1622 (O_1622,N_14820,N_14775);
and UO_1623 (O_1623,N_14539,N_14511);
nand UO_1624 (O_1624,N_14885,N_14637);
nand UO_1625 (O_1625,N_14824,N_14908);
xor UO_1626 (O_1626,N_14542,N_14804);
and UO_1627 (O_1627,N_14659,N_14646);
or UO_1628 (O_1628,N_14524,N_14714);
nand UO_1629 (O_1629,N_14859,N_14719);
nand UO_1630 (O_1630,N_14849,N_14599);
or UO_1631 (O_1631,N_14817,N_14804);
nand UO_1632 (O_1632,N_14694,N_14637);
or UO_1633 (O_1633,N_14719,N_14716);
nor UO_1634 (O_1634,N_14968,N_14929);
nor UO_1635 (O_1635,N_14838,N_14558);
nor UO_1636 (O_1636,N_14591,N_14813);
or UO_1637 (O_1637,N_14627,N_14877);
xnor UO_1638 (O_1638,N_14600,N_14959);
nor UO_1639 (O_1639,N_14799,N_14862);
xnor UO_1640 (O_1640,N_14836,N_14878);
or UO_1641 (O_1641,N_14885,N_14751);
nand UO_1642 (O_1642,N_14829,N_14960);
nor UO_1643 (O_1643,N_14759,N_14571);
nand UO_1644 (O_1644,N_14511,N_14814);
nand UO_1645 (O_1645,N_14719,N_14523);
and UO_1646 (O_1646,N_14616,N_14660);
xnor UO_1647 (O_1647,N_14861,N_14966);
nor UO_1648 (O_1648,N_14557,N_14598);
nand UO_1649 (O_1649,N_14726,N_14605);
or UO_1650 (O_1650,N_14784,N_14828);
or UO_1651 (O_1651,N_14801,N_14881);
nor UO_1652 (O_1652,N_14528,N_14522);
nor UO_1653 (O_1653,N_14930,N_14518);
nor UO_1654 (O_1654,N_14880,N_14710);
xor UO_1655 (O_1655,N_14622,N_14709);
nand UO_1656 (O_1656,N_14869,N_14521);
nor UO_1657 (O_1657,N_14592,N_14918);
and UO_1658 (O_1658,N_14739,N_14960);
nand UO_1659 (O_1659,N_14591,N_14744);
and UO_1660 (O_1660,N_14692,N_14526);
xor UO_1661 (O_1661,N_14583,N_14560);
nand UO_1662 (O_1662,N_14993,N_14952);
and UO_1663 (O_1663,N_14743,N_14812);
xnor UO_1664 (O_1664,N_14670,N_14501);
nand UO_1665 (O_1665,N_14912,N_14924);
and UO_1666 (O_1666,N_14741,N_14779);
and UO_1667 (O_1667,N_14620,N_14814);
nor UO_1668 (O_1668,N_14722,N_14512);
or UO_1669 (O_1669,N_14577,N_14533);
nand UO_1670 (O_1670,N_14579,N_14978);
xor UO_1671 (O_1671,N_14654,N_14543);
and UO_1672 (O_1672,N_14703,N_14596);
xor UO_1673 (O_1673,N_14750,N_14807);
nand UO_1674 (O_1674,N_14834,N_14836);
or UO_1675 (O_1675,N_14539,N_14623);
and UO_1676 (O_1676,N_14620,N_14843);
nor UO_1677 (O_1677,N_14796,N_14827);
nor UO_1678 (O_1678,N_14607,N_14569);
xor UO_1679 (O_1679,N_14524,N_14882);
or UO_1680 (O_1680,N_14958,N_14612);
xnor UO_1681 (O_1681,N_14551,N_14879);
and UO_1682 (O_1682,N_14779,N_14701);
nor UO_1683 (O_1683,N_14688,N_14649);
nand UO_1684 (O_1684,N_14617,N_14895);
or UO_1685 (O_1685,N_14835,N_14714);
and UO_1686 (O_1686,N_14993,N_14514);
nor UO_1687 (O_1687,N_14957,N_14878);
and UO_1688 (O_1688,N_14521,N_14916);
xnor UO_1689 (O_1689,N_14637,N_14697);
and UO_1690 (O_1690,N_14667,N_14617);
xor UO_1691 (O_1691,N_14815,N_14999);
or UO_1692 (O_1692,N_14503,N_14923);
and UO_1693 (O_1693,N_14786,N_14809);
or UO_1694 (O_1694,N_14997,N_14925);
nor UO_1695 (O_1695,N_14555,N_14887);
nor UO_1696 (O_1696,N_14574,N_14680);
or UO_1697 (O_1697,N_14971,N_14735);
nor UO_1698 (O_1698,N_14598,N_14545);
xnor UO_1699 (O_1699,N_14937,N_14935);
and UO_1700 (O_1700,N_14789,N_14828);
nand UO_1701 (O_1701,N_14955,N_14870);
xor UO_1702 (O_1702,N_14760,N_14663);
xor UO_1703 (O_1703,N_14584,N_14625);
or UO_1704 (O_1704,N_14734,N_14599);
nor UO_1705 (O_1705,N_14959,N_14532);
nor UO_1706 (O_1706,N_14933,N_14510);
and UO_1707 (O_1707,N_14917,N_14928);
nor UO_1708 (O_1708,N_14916,N_14864);
xor UO_1709 (O_1709,N_14801,N_14876);
nor UO_1710 (O_1710,N_14652,N_14708);
or UO_1711 (O_1711,N_14935,N_14521);
xnor UO_1712 (O_1712,N_14859,N_14883);
nor UO_1713 (O_1713,N_14774,N_14941);
nor UO_1714 (O_1714,N_14630,N_14683);
or UO_1715 (O_1715,N_14871,N_14932);
nor UO_1716 (O_1716,N_14503,N_14979);
or UO_1717 (O_1717,N_14654,N_14813);
nand UO_1718 (O_1718,N_14837,N_14760);
and UO_1719 (O_1719,N_14641,N_14921);
and UO_1720 (O_1720,N_14663,N_14570);
and UO_1721 (O_1721,N_14760,N_14714);
or UO_1722 (O_1722,N_14669,N_14940);
and UO_1723 (O_1723,N_14933,N_14601);
or UO_1724 (O_1724,N_14885,N_14895);
or UO_1725 (O_1725,N_14690,N_14612);
nand UO_1726 (O_1726,N_14979,N_14717);
nand UO_1727 (O_1727,N_14658,N_14568);
nand UO_1728 (O_1728,N_14978,N_14991);
nor UO_1729 (O_1729,N_14764,N_14704);
xor UO_1730 (O_1730,N_14821,N_14557);
xnor UO_1731 (O_1731,N_14597,N_14887);
or UO_1732 (O_1732,N_14979,N_14739);
nand UO_1733 (O_1733,N_14785,N_14836);
nand UO_1734 (O_1734,N_14553,N_14849);
xor UO_1735 (O_1735,N_14528,N_14686);
xnor UO_1736 (O_1736,N_14767,N_14919);
or UO_1737 (O_1737,N_14729,N_14603);
xor UO_1738 (O_1738,N_14646,N_14716);
nand UO_1739 (O_1739,N_14766,N_14911);
and UO_1740 (O_1740,N_14546,N_14876);
xnor UO_1741 (O_1741,N_14607,N_14862);
or UO_1742 (O_1742,N_14555,N_14500);
or UO_1743 (O_1743,N_14907,N_14886);
nand UO_1744 (O_1744,N_14784,N_14736);
xnor UO_1745 (O_1745,N_14771,N_14919);
xnor UO_1746 (O_1746,N_14915,N_14759);
or UO_1747 (O_1747,N_14957,N_14748);
or UO_1748 (O_1748,N_14979,N_14829);
xnor UO_1749 (O_1749,N_14744,N_14582);
and UO_1750 (O_1750,N_14622,N_14514);
or UO_1751 (O_1751,N_14604,N_14642);
and UO_1752 (O_1752,N_14721,N_14598);
xor UO_1753 (O_1753,N_14659,N_14506);
or UO_1754 (O_1754,N_14916,N_14625);
nand UO_1755 (O_1755,N_14965,N_14544);
nor UO_1756 (O_1756,N_14792,N_14816);
nor UO_1757 (O_1757,N_14897,N_14890);
and UO_1758 (O_1758,N_14674,N_14977);
nor UO_1759 (O_1759,N_14620,N_14736);
and UO_1760 (O_1760,N_14886,N_14963);
or UO_1761 (O_1761,N_14818,N_14926);
or UO_1762 (O_1762,N_14670,N_14934);
nand UO_1763 (O_1763,N_14868,N_14626);
nor UO_1764 (O_1764,N_14807,N_14708);
nand UO_1765 (O_1765,N_14663,N_14550);
nand UO_1766 (O_1766,N_14915,N_14600);
xor UO_1767 (O_1767,N_14627,N_14508);
nor UO_1768 (O_1768,N_14695,N_14781);
and UO_1769 (O_1769,N_14950,N_14573);
nor UO_1770 (O_1770,N_14893,N_14806);
nor UO_1771 (O_1771,N_14766,N_14887);
and UO_1772 (O_1772,N_14983,N_14781);
or UO_1773 (O_1773,N_14873,N_14916);
nor UO_1774 (O_1774,N_14554,N_14783);
xor UO_1775 (O_1775,N_14691,N_14568);
nor UO_1776 (O_1776,N_14580,N_14800);
nor UO_1777 (O_1777,N_14986,N_14608);
nor UO_1778 (O_1778,N_14666,N_14510);
nand UO_1779 (O_1779,N_14962,N_14662);
xor UO_1780 (O_1780,N_14545,N_14912);
xor UO_1781 (O_1781,N_14682,N_14556);
and UO_1782 (O_1782,N_14720,N_14807);
or UO_1783 (O_1783,N_14910,N_14857);
xor UO_1784 (O_1784,N_14710,N_14563);
and UO_1785 (O_1785,N_14861,N_14757);
nor UO_1786 (O_1786,N_14500,N_14596);
and UO_1787 (O_1787,N_14958,N_14711);
nor UO_1788 (O_1788,N_14916,N_14503);
xnor UO_1789 (O_1789,N_14568,N_14650);
and UO_1790 (O_1790,N_14538,N_14643);
and UO_1791 (O_1791,N_14788,N_14671);
nand UO_1792 (O_1792,N_14969,N_14678);
xor UO_1793 (O_1793,N_14750,N_14644);
nand UO_1794 (O_1794,N_14618,N_14706);
xor UO_1795 (O_1795,N_14577,N_14570);
or UO_1796 (O_1796,N_14649,N_14531);
nand UO_1797 (O_1797,N_14526,N_14731);
and UO_1798 (O_1798,N_14979,N_14948);
nor UO_1799 (O_1799,N_14698,N_14856);
or UO_1800 (O_1800,N_14503,N_14696);
xor UO_1801 (O_1801,N_14679,N_14716);
nor UO_1802 (O_1802,N_14789,N_14570);
and UO_1803 (O_1803,N_14728,N_14581);
nor UO_1804 (O_1804,N_14722,N_14993);
nand UO_1805 (O_1805,N_14569,N_14925);
nor UO_1806 (O_1806,N_14674,N_14881);
nor UO_1807 (O_1807,N_14789,N_14847);
nand UO_1808 (O_1808,N_14970,N_14935);
xor UO_1809 (O_1809,N_14550,N_14516);
and UO_1810 (O_1810,N_14951,N_14532);
nor UO_1811 (O_1811,N_14517,N_14994);
xor UO_1812 (O_1812,N_14528,N_14773);
xnor UO_1813 (O_1813,N_14558,N_14979);
or UO_1814 (O_1814,N_14811,N_14685);
nor UO_1815 (O_1815,N_14543,N_14791);
nand UO_1816 (O_1816,N_14537,N_14821);
and UO_1817 (O_1817,N_14544,N_14634);
nor UO_1818 (O_1818,N_14521,N_14774);
xor UO_1819 (O_1819,N_14965,N_14688);
and UO_1820 (O_1820,N_14684,N_14835);
xnor UO_1821 (O_1821,N_14711,N_14607);
and UO_1822 (O_1822,N_14942,N_14555);
nor UO_1823 (O_1823,N_14726,N_14644);
and UO_1824 (O_1824,N_14697,N_14927);
nor UO_1825 (O_1825,N_14896,N_14842);
or UO_1826 (O_1826,N_14929,N_14804);
and UO_1827 (O_1827,N_14998,N_14712);
nor UO_1828 (O_1828,N_14822,N_14860);
nand UO_1829 (O_1829,N_14686,N_14941);
nor UO_1830 (O_1830,N_14532,N_14931);
nor UO_1831 (O_1831,N_14532,N_14576);
and UO_1832 (O_1832,N_14553,N_14871);
or UO_1833 (O_1833,N_14631,N_14771);
nor UO_1834 (O_1834,N_14861,N_14815);
xnor UO_1835 (O_1835,N_14789,N_14610);
xnor UO_1836 (O_1836,N_14858,N_14855);
nor UO_1837 (O_1837,N_14542,N_14723);
and UO_1838 (O_1838,N_14944,N_14720);
nand UO_1839 (O_1839,N_14687,N_14868);
and UO_1840 (O_1840,N_14698,N_14780);
nor UO_1841 (O_1841,N_14846,N_14885);
and UO_1842 (O_1842,N_14946,N_14701);
nand UO_1843 (O_1843,N_14746,N_14859);
nor UO_1844 (O_1844,N_14651,N_14587);
nor UO_1845 (O_1845,N_14886,N_14895);
nand UO_1846 (O_1846,N_14874,N_14987);
or UO_1847 (O_1847,N_14654,N_14503);
and UO_1848 (O_1848,N_14537,N_14903);
nor UO_1849 (O_1849,N_14668,N_14847);
nand UO_1850 (O_1850,N_14994,N_14836);
nor UO_1851 (O_1851,N_14681,N_14652);
nand UO_1852 (O_1852,N_14732,N_14981);
nor UO_1853 (O_1853,N_14574,N_14522);
or UO_1854 (O_1854,N_14656,N_14760);
or UO_1855 (O_1855,N_14994,N_14773);
nand UO_1856 (O_1856,N_14886,N_14888);
or UO_1857 (O_1857,N_14759,N_14809);
nand UO_1858 (O_1858,N_14611,N_14681);
and UO_1859 (O_1859,N_14785,N_14951);
and UO_1860 (O_1860,N_14738,N_14540);
or UO_1861 (O_1861,N_14819,N_14663);
nand UO_1862 (O_1862,N_14828,N_14527);
nor UO_1863 (O_1863,N_14632,N_14941);
xor UO_1864 (O_1864,N_14901,N_14645);
or UO_1865 (O_1865,N_14954,N_14500);
and UO_1866 (O_1866,N_14788,N_14833);
or UO_1867 (O_1867,N_14724,N_14556);
nor UO_1868 (O_1868,N_14812,N_14841);
xor UO_1869 (O_1869,N_14979,N_14542);
or UO_1870 (O_1870,N_14709,N_14691);
nand UO_1871 (O_1871,N_14673,N_14841);
nor UO_1872 (O_1872,N_14798,N_14991);
nor UO_1873 (O_1873,N_14946,N_14541);
nand UO_1874 (O_1874,N_14741,N_14983);
xor UO_1875 (O_1875,N_14565,N_14977);
and UO_1876 (O_1876,N_14666,N_14868);
or UO_1877 (O_1877,N_14735,N_14575);
nor UO_1878 (O_1878,N_14698,N_14694);
and UO_1879 (O_1879,N_14867,N_14796);
and UO_1880 (O_1880,N_14744,N_14779);
nand UO_1881 (O_1881,N_14911,N_14516);
nand UO_1882 (O_1882,N_14817,N_14669);
or UO_1883 (O_1883,N_14931,N_14860);
and UO_1884 (O_1884,N_14815,N_14667);
nor UO_1885 (O_1885,N_14663,N_14647);
xor UO_1886 (O_1886,N_14867,N_14635);
nor UO_1887 (O_1887,N_14608,N_14729);
xor UO_1888 (O_1888,N_14957,N_14754);
nor UO_1889 (O_1889,N_14792,N_14657);
and UO_1890 (O_1890,N_14904,N_14694);
xnor UO_1891 (O_1891,N_14870,N_14595);
and UO_1892 (O_1892,N_14614,N_14781);
nand UO_1893 (O_1893,N_14954,N_14609);
nand UO_1894 (O_1894,N_14580,N_14641);
and UO_1895 (O_1895,N_14638,N_14726);
or UO_1896 (O_1896,N_14915,N_14984);
nand UO_1897 (O_1897,N_14890,N_14938);
and UO_1898 (O_1898,N_14998,N_14690);
and UO_1899 (O_1899,N_14603,N_14680);
or UO_1900 (O_1900,N_14739,N_14843);
nand UO_1901 (O_1901,N_14592,N_14653);
nand UO_1902 (O_1902,N_14934,N_14765);
nand UO_1903 (O_1903,N_14868,N_14591);
xnor UO_1904 (O_1904,N_14747,N_14821);
and UO_1905 (O_1905,N_14609,N_14716);
and UO_1906 (O_1906,N_14959,N_14515);
or UO_1907 (O_1907,N_14509,N_14946);
nand UO_1908 (O_1908,N_14575,N_14662);
nand UO_1909 (O_1909,N_14666,N_14783);
or UO_1910 (O_1910,N_14724,N_14901);
xnor UO_1911 (O_1911,N_14564,N_14828);
xor UO_1912 (O_1912,N_14570,N_14860);
nand UO_1913 (O_1913,N_14714,N_14520);
nand UO_1914 (O_1914,N_14834,N_14843);
or UO_1915 (O_1915,N_14912,N_14720);
nor UO_1916 (O_1916,N_14563,N_14757);
or UO_1917 (O_1917,N_14601,N_14578);
and UO_1918 (O_1918,N_14544,N_14627);
xnor UO_1919 (O_1919,N_14737,N_14575);
nand UO_1920 (O_1920,N_14893,N_14896);
or UO_1921 (O_1921,N_14764,N_14878);
xnor UO_1922 (O_1922,N_14617,N_14945);
nor UO_1923 (O_1923,N_14513,N_14777);
and UO_1924 (O_1924,N_14958,N_14932);
and UO_1925 (O_1925,N_14757,N_14976);
nor UO_1926 (O_1926,N_14714,N_14909);
nand UO_1927 (O_1927,N_14989,N_14951);
nor UO_1928 (O_1928,N_14638,N_14612);
nand UO_1929 (O_1929,N_14672,N_14541);
or UO_1930 (O_1930,N_14974,N_14577);
and UO_1931 (O_1931,N_14500,N_14974);
nor UO_1932 (O_1932,N_14955,N_14597);
and UO_1933 (O_1933,N_14617,N_14774);
and UO_1934 (O_1934,N_14758,N_14578);
or UO_1935 (O_1935,N_14990,N_14712);
and UO_1936 (O_1936,N_14924,N_14972);
nor UO_1937 (O_1937,N_14530,N_14950);
xnor UO_1938 (O_1938,N_14517,N_14533);
or UO_1939 (O_1939,N_14969,N_14523);
and UO_1940 (O_1940,N_14652,N_14695);
xnor UO_1941 (O_1941,N_14940,N_14922);
nand UO_1942 (O_1942,N_14974,N_14641);
nand UO_1943 (O_1943,N_14969,N_14973);
nand UO_1944 (O_1944,N_14607,N_14554);
and UO_1945 (O_1945,N_14695,N_14559);
or UO_1946 (O_1946,N_14672,N_14506);
nor UO_1947 (O_1947,N_14564,N_14765);
nand UO_1948 (O_1948,N_14580,N_14764);
nand UO_1949 (O_1949,N_14517,N_14581);
and UO_1950 (O_1950,N_14653,N_14604);
xor UO_1951 (O_1951,N_14555,N_14944);
and UO_1952 (O_1952,N_14708,N_14697);
or UO_1953 (O_1953,N_14951,N_14851);
nand UO_1954 (O_1954,N_14711,N_14907);
and UO_1955 (O_1955,N_14534,N_14999);
nand UO_1956 (O_1956,N_14695,N_14806);
or UO_1957 (O_1957,N_14845,N_14951);
nor UO_1958 (O_1958,N_14990,N_14552);
and UO_1959 (O_1959,N_14955,N_14850);
nor UO_1960 (O_1960,N_14686,N_14536);
or UO_1961 (O_1961,N_14520,N_14750);
xnor UO_1962 (O_1962,N_14799,N_14698);
nor UO_1963 (O_1963,N_14990,N_14574);
or UO_1964 (O_1964,N_14973,N_14509);
or UO_1965 (O_1965,N_14582,N_14597);
xor UO_1966 (O_1966,N_14863,N_14568);
nand UO_1967 (O_1967,N_14734,N_14686);
nand UO_1968 (O_1968,N_14933,N_14848);
xnor UO_1969 (O_1969,N_14745,N_14774);
or UO_1970 (O_1970,N_14524,N_14880);
or UO_1971 (O_1971,N_14990,N_14861);
xor UO_1972 (O_1972,N_14785,N_14551);
nor UO_1973 (O_1973,N_14920,N_14863);
nand UO_1974 (O_1974,N_14828,N_14824);
nor UO_1975 (O_1975,N_14624,N_14812);
or UO_1976 (O_1976,N_14794,N_14841);
or UO_1977 (O_1977,N_14936,N_14500);
nand UO_1978 (O_1978,N_14755,N_14639);
or UO_1979 (O_1979,N_14673,N_14531);
nand UO_1980 (O_1980,N_14705,N_14649);
or UO_1981 (O_1981,N_14590,N_14791);
xor UO_1982 (O_1982,N_14915,N_14758);
nand UO_1983 (O_1983,N_14754,N_14931);
and UO_1984 (O_1984,N_14840,N_14992);
and UO_1985 (O_1985,N_14569,N_14573);
xnor UO_1986 (O_1986,N_14832,N_14706);
nor UO_1987 (O_1987,N_14904,N_14597);
or UO_1988 (O_1988,N_14801,N_14999);
nor UO_1989 (O_1989,N_14654,N_14546);
xor UO_1990 (O_1990,N_14759,N_14930);
nand UO_1991 (O_1991,N_14890,N_14858);
or UO_1992 (O_1992,N_14973,N_14644);
and UO_1993 (O_1993,N_14547,N_14516);
nor UO_1994 (O_1994,N_14767,N_14732);
nand UO_1995 (O_1995,N_14860,N_14682);
nor UO_1996 (O_1996,N_14592,N_14747);
or UO_1997 (O_1997,N_14585,N_14599);
or UO_1998 (O_1998,N_14870,N_14505);
nor UO_1999 (O_1999,N_14821,N_14879);
endmodule