module basic_2500_25000_3000_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_913,In_2035);
or U1 (N_1,In_900,In_1914);
and U2 (N_2,In_322,In_1308);
xor U3 (N_3,In_1038,In_2172);
and U4 (N_4,In_1042,In_1260);
nor U5 (N_5,In_1328,In_1591);
xor U6 (N_6,In_418,In_2375);
xnor U7 (N_7,In_129,In_241);
and U8 (N_8,In_1726,In_1334);
xnor U9 (N_9,In_396,In_640);
and U10 (N_10,In_1539,In_748);
nand U11 (N_11,In_113,In_684);
and U12 (N_12,In_1882,In_1001);
xnor U13 (N_13,In_2395,In_553);
nand U14 (N_14,In_679,In_1122);
xnor U15 (N_15,In_1926,In_7);
xnor U16 (N_16,In_472,In_1300);
or U17 (N_17,In_116,In_1250);
xnor U18 (N_18,In_2236,In_284);
xnor U19 (N_19,In_2162,In_2198);
nand U20 (N_20,In_1477,In_2000);
nand U21 (N_21,In_1292,In_1521);
nor U22 (N_22,In_221,In_2224);
nor U23 (N_23,In_1320,In_1850);
and U24 (N_24,In_428,In_40);
nor U25 (N_25,In_192,In_2194);
nand U26 (N_26,In_2452,In_257);
nand U27 (N_27,In_514,In_471);
and U28 (N_28,In_1186,In_1262);
or U29 (N_29,In_2130,In_2079);
nor U30 (N_30,In_924,In_1963);
nor U31 (N_31,In_2281,In_1945);
and U32 (N_32,In_1612,In_321);
and U33 (N_33,In_82,In_1708);
nor U34 (N_34,In_2317,In_1062);
xor U35 (N_35,In_711,In_64);
nor U36 (N_36,In_1993,In_1840);
and U37 (N_37,In_1131,In_21);
xor U38 (N_38,In_1699,In_1057);
nand U39 (N_39,In_1273,In_1854);
nand U40 (N_40,In_2013,In_1112);
nor U41 (N_41,In_857,In_829);
nand U42 (N_42,In_448,In_254);
or U43 (N_43,In_2409,In_1104);
and U44 (N_44,In_1567,In_2476);
nand U45 (N_45,In_2125,In_1382);
and U46 (N_46,In_56,In_1698);
nor U47 (N_47,In_2093,In_2420);
nor U48 (N_48,In_981,In_1798);
and U49 (N_49,In_654,In_2331);
xnor U50 (N_50,In_740,In_1748);
xor U51 (N_51,In_653,In_736);
nand U52 (N_52,In_1818,In_706);
nor U53 (N_53,In_60,In_1747);
xor U54 (N_54,In_1330,In_52);
xnor U55 (N_55,In_443,In_1126);
xnor U56 (N_56,In_2306,In_2199);
and U57 (N_57,In_2488,In_1618);
and U58 (N_58,In_390,In_224);
xnor U59 (N_59,In_1461,In_1499);
nor U60 (N_60,In_1865,In_1658);
xnor U61 (N_61,In_1381,In_144);
nor U62 (N_62,In_128,In_1588);
or U63 (N_63,In_1428,In_1366);
xor U64 (N_64,In_1243,In_2201);
nand U65 (N_65,In_1210,In_1206);
and U66 (N_66,In_1183,In_747);
and U67 (N_67,In_1220,In_1981);
nor U68 (N_68,In_1507,In_37);
nor U69 (N_69,In_1103,In_2474);
or U70 (N_70,In_1304,In_1741);
nand U71 (N_71,In_2134,In_2086);
xnor U72 (N_72,In_1140,In_1930);
or U73 (N_73,In_489,In_1019);
or U74 (N_74,In_1291,In_1271);
or U75 (N_75,In_518,In_2104);
nand U76 (N_76,In_1080,In_734);
nand U77 (N_77,In_1830,In_1111);
and U78 (N_78,In_571,In_267);
and U79 (N_79,In_2167,In_138);
or U80 (N_80,In_1848,In_2124);
or U81 (N_81,In_344,In_2370);
or U82 (N_82,In_1996,In_2227);
or U83 (N_83,In_1666,In_2373);
xor U84 (N_84,In_2112,In_122);
nor U85 (N_85,In_843,In_1991);
and U86 (N_86,In_1011,In_1418);
nor U87 (N_87,In_1437,In_1749);
or U88 (N_88,In_2444,In_1227);
nand U89 (N_89,In_877,In_2491);
nand U90 (N_90,In_520,In_1797);
nor U91 (N_91,In_1376,In_1462);
xor U92 (N_92,In_1731,In_2011);
and U93 (N_93,In_146,In_2100);
nor U94 (N_94,In_1026,In_1359);
xnor U95 (N_95,In_865,In_2269);
or U96 (N_96,In_1694,In_899);
xnor U97 (N_97,In_11,In_2188);
and U98 (N_98,In_824,In_2412);
and U99 (N_99,In_278,In_339);
xnor U100 (N_100,In_2047,In_1412);
or U101 (N_101,In_2320,In_1609);
or U102 (N_102,In_2132,In_889);
nor U103 (N_103,In_1225,In_986);
nor U104 (N_104,In_1237,In_746);
and U105 (N_105,In_1447,In_440);
nand U106 (N_106,In_605,In_570);
and U107 (N_107,In_1795,In_1817);
and U108 (N_108,In_326,In_2020);
or U109 (N_109,In_1143,In_1617);
nand U110 (N_110,In_346,In_946);
or U111 (N_111,In_1894,In_1097);
xor U112 (N_112,In_2063,In_1701);
nor U113 (N_113,In_1843,In_2092);
and U114 (N_114,In_2360,In_473);
xnor U115 (N_115,In_2021,In_2085);
or U116 (N_116,In_768,In_407);
nor U117 (N_117,In_1657,In_338);
nor U118 (N_118,In_1254,In_2296);
xor U119 (N_119,In_1472,In_2492);
nor U120 (N_120,In_1092,In_875);
or U121 (N_121,In_6,In_1460);
or U122 (N_122,In_2155,In_356);
and U123 (N_123,In_389,In_94);
or U124 (N_124,In_766,In_2447);
and U125 (N_125,In_1885,In_2329);
and U126 (N_126,In_1547,In_2258);
xnor U127 (N_127,In_1685,In_1009);
nand U128 (N_128,In_1425,In_751);
xnor U129 (N_129,In_667,In_232);
and U130 (N_130,In_234,In_1501);
and U131 (N_131,In_2245,In_1051);
xnor U132 (N_132,In_646,In_531);
nor U133 (N_133,In_225,In_2486);
xnor U134 (N_134,In_853,In_2299);
or U135 (N_135,In_1296,In_806);
and U136 (N_136,In_1934,In_1989);
xor U137 (N_137,In_1692,In_1691);
nand U138 (N_138,In_2267,In_850);
xnor U139 (N_139,In_1956,In_1649);
and U140 (N_140,In_2138,In_598);
nand U141 (N_141,In_1377,In_1994);
and U142 (N_142,In_1369,In_2300);
xnor U143 (N_143,In_468,In_2025);
and U144 (N_144,In_950,In_770);
nand U145 (N_145,In_231,In_625);
nand U146 (N_146,In_1804,In_687);
and U147 (N_147,In_1864,In_1238);
nor U148 (N_148,In_1975,In_2131);
or U149 (N_149,In_233,In_228);
or U150 (N_150,In_891,In_24);
nor U151 (N_151,In_2323,In_1556);
or U152 (N_152,In_1253,In_1760);
nor U153 (N_153,In_554,In_1397);
nor U154 (N_154,In_584,In_272);
and U155 (N_155,In_543,In_483);
and U156 (N_156,In_682,In_1141);
or U157 (N_157,In_894,In_1125);
and U158 (N_158,In_1577,In_1811);
nand U159 (N_159,In_1889,In_2365);
xor U160 (N_160,In_317,In_504);
nor U161 (N_161,In_561,In_2284);
nand U162 (N_162,In_1442,In_1786);
nor U163 (N_163,In_1927,In_1343);
or U164 (N_164,In_941,In_1039);
nand U165 (N_165,In_2228,In_719);
nand U166 (N_166,In_2352,In_179);
nand U167 (N_167,In_1219,In_2128);
nand U168 (N_168,In_691,In_935);
xor U169 (N_169,In_2213,In_1118);
nor U170 (N_170,In_147,In_1587);
nor U171 (N_171,In_2393,In_488);
nor U172 (N_172,In_2127,In_2216);
and U173 (N_173,In_1791,In_1076);
nor U174 (N_174,In_1826,In_2206);
nor U175 (N_175,In_1720,In_217);
nor U176 (N_176,In_929,In_970);
or U177 (N_177,In_1813,In_1498);
xor U178 (N_178,In_1710,In_972);
and U179 (N_179,In_2405,In_817);
and U180 (N_180,In_329,In_1548);
nor U181 (N_181,In_2295,In_1959);
and U182 (N_182,In_919,In_1347);
xnor U183 (N_183,In_481,In_2310);
and U184 (N_184,In_874,In_2432);
and U185 (N_185,In_1435,In_2460);
or U186 (N_186,In_1806,In_1652);
and U187 (N_187,In_505,In_693);
or U188 (N_188,In_1890,In_1695);
and U189 (N_189,In_593,In_14);
xnor U190 (N_190,In_1054,In_189);
and U191 (N_191,In_1871,In_1490);
and U192 (N_192,In_2034,In_1302);
nor U193 (N_193,In_340,In_1506);
nor U194 (N_194,In_2232,In_1439);
or U195 (N_195,In_676,In_771);
xor U196 (N_196,In_1,In_2303);
and U197 (N_197,In_292,In_487);
nor U198 (N_198,In_1241,In_1069);
nor U199 (N_199,In_500,In_1383);
nor U200 (N_200,In_1642,In_1113);
or U201 (N_201,In_1318,In_1966);
and U202 (N_202,In_136,In_2146);
nand U203 (N_203,In_1458,In_883);
and U204 (N_204,In_2218,In_989);
or U205 (N_205,In_2166,In_1646);
or U206 (N_206,In_484,In_1230);
or U207 (N_207,In_2390,In_1083);
and U208 (N_208,In_810,In_290);
nor U209 (N_209,In_669,In_2164);
nor U210 (N_210,In_410,In_635);
nand U211 (N_211,In_738,In_2380);
nand U212 (N_212,In_2304,In_218);
nand U213 (N_213,In_1732,In_261);
nand U214 (N_214,In_2297,In_967);
or U215 (N_215,In_195,In_1488);
nand U216 (N_216,In_1492,In_955);
nor U217 (N_217,In_1373,In_403);
and U218 (N_218,In_1182,In_2436);
xnor U219 (N_219,In_162,In_25);
xor U220 (N_220,In_2046,In_2001);
xor U221 (N_221,In_1638,In_2429);
or U222 (N_222,In_1820,In_1772);
xor U223 (N_223,In_2066,In_1423);
and U224 (N_224,In_1473,In_475);
and U225 (N_225,In_2345,In_2276);
or U226 (N_226,In_69,In_1440);
or U227 (N_227,In_909,In_1457);
nand U228 (N_228,In_1936,In_840);
nor U229 (N_229,In_2457,In_809);
or U230 (N_230,In_651,In_2038);
nor U231 (N_231,In_72,In_1689);
and U232 (N_232,In_2449,In_681);
and U233 (N_233,In_1625,In_786);
nor U234 (N_234,In_1297,In_2424);
nand U235 (N_235,In_1082,In_1718);
or U236 (N_236,In_616,In_490);
nand U237 (N_237,In_1816,In_1604);
and U238 (N_238,In_452,In_1846);
nand U239 (N_239,In_931,In_1041);
xnor U240 (N_240,In_541,In_1315);
or U241 (N_241,In_2059,In_515);
nand U242 (N_242,In_708,In_145);
or U243 (N_243,In_2248,In_1399);
nand U244 (N_244,In_818,In_1116);
xor U245 (N_245,In_96,In_2110);
nand U246 (N_246,In_414,In_4);
nand U247 (N_247,In_1419,In_188);
nor U248 (N_248,In_1724,In_2207);
or U249 (N_249,In_3,In_1348);
and U250 (N_250,In_633,In_271);
and U251 (N_251,In_2448,In_2142);
xnor U252 (N_252,In_943,In_243);
nand U253 (N_253,In_2455,In_1615);
xor U254 (N_254,In_49,In_103);
nor U255 (N_255,In_2347,In_1660);
or U256 (N_256,In_1124,In_1520);
xnor U257 (N_257,In_1757,In_334);
or U258 (N_258,In_1775,In_212);
nand U259 (N_259,In_1332,In_2439);
nor U260 (N_260,In_1810,In_2179);
nand U261 (N_261,In_201,In_976);
xnor U262 (N_262,In_2010,In_2438);
nor U263 (N_263,In_2264,In_19);
and U264 (N_264,In_199,In_1246);
nor U265 (N_265,In_741,In_2386);
nand U266 (N_266,In_978,In_626);
xnor U267 (N_267,In_577,In_1187);
xnor U268 (N_268,In_269,In_1168);
nand U269 (N_269,In_1481,In_2009);
xor U270 (N_270,In_2261,In_1663);
nor U271 (N_271,In_1362,In_1607);
nand U272 (N_272,In_2048,In_672);
xor U273 (N_273,In_363,In_1029);
nand U274 (N_274,In_2374,In_265);
or U275 (N_275,In_2073,In_545);
xnor U276 (N_276,In_1845,In_730);
xnor U277 (N_277,In_1368,In_157);
nand U278 (N_278,In_957,In_130);
nand U279 (N_279,In_932,In_841);
or U280 (N_280,In_132,In_790);
and U281 (N_281,In_1783,In_222);
nor U282 (N_282,In_1782,In_1570);
xor U283 (N_283,In_1110,In_1193);
nand U284 (N_284,In_1217,In_610);
or U285 (N_285,In_433,In_1768);
nand U286 (N_286,In_470,In_1231);
or U287 (N_287,In_629,In_108);
or U288 (N_288,In_1537,In_1478);
or U289 (N_289,In_1221,In_839);
and U290 (N_290,In_259,In_1849);
nor U291 (N_291,In_1878,In_670);
or U292 (N_292,In_235,In_1269);
xnor U293 (N_293,In_1668,In_1678);
xor U294 (N_294,In_798,In_2381);
nand U295 (N_295,In_2174,In_9);
and U296 (N_296,In_1593,In_2200);
or U297 (N_297,In_2487,In_83);
and U298 (N_298,In_675,In_2400);
xor U299 (N_299,In_1319,In_851);
or U300 (N_300,In_1831,In_2406);
xor U301 (N_301,In_954,In_213);
or U302 (N_302,In_1151,In_2181);
nor U303 (N_303,In_1215,In_1050);
or U304 (N_304,In_1228,In_365);
and U305 (N_305,In_358,In_1700);
xnor U306 (N_306,In_1165,In_886);
nand U307 (N_307,In_523,In_1900);
nand U308 (N_308,In_247,In_1340);
nor U309 (N_309,In_2493,In_1552);
nand U310 (N_310,In_1713,In_193);
or U311 (N_311,In_1821,In_830);
and U312 (N_312,In_1863,In_1200);
or U313 (N_313,In_975,In_623);
xor U314 (N_314,In_1239,In_2252);
and U315 (N_315,In_1654,In_266);
and U316 (N_316,In_1115,In_1363);
and U317 (N_317,In_1367,In_239);
or U318 (N_318,In_996,In_141);
and U319 (N_319,In_1469,In_1190);
or U320 (N_320,In_35,In_1489);
nor U321 (N_321,In_2017,In_30);
nand U322 (N_322,In_174,In_1542);
nor U323 (N_323,In_1261,In_121);
nand U324 (N_324,In_697,In_808);
nor U325 (N_325,In_1455,In_78);
and U326 (N_326,In_778,In_2120);
or U327 (N_327,In_592,In_1941);
and U328 (N_328,In_926,In_2369);
nand U329 (N_329,In_2050,In_1555);
and U330 (N_330,In_1661,In_1703);
nor U331 (N_331,In_1647,In_1378);
nor U332 (N_332,In_148,In_295);
and U333 (N_333,In_630,In_614);
or U334 (N_334,In_200,In_958);
xnor U335 (N_335,In_2278,In_2082);
nand U336 (N_336,In_2437,In_683);
nor U337 (N_337,In_2163,In_1780);
and U338 (N_338,In_1331,In_720);
and U339 (N_339,In_2154,In_793);
xnor U340 (N_340,In_2483,In_1847);
xnor U341 (N_341,In_463,In_1773);
or U342 (N_342,In_451,In_781);
or U343 (N_343,In_2084,In_1453);
and U344 (N_344,In_774,In_952);
nand U345 (N_345,In_462,In_449);
nand U346 (N_346,In_210,In_624);
xor U347 (N_347,In_726,In_392);
nand U348 (N_348,In_1549,In_767);
xnor U349 (N_349,In_53,In_1532);
or U350 (N_350,In_123,In_999);
nand U351 (N_351,In_1248,In_1424);
or U352 (N_352,In_2143,In_2496);
xor U353 (N_353,In_1842,In_1895);
and U354 (N_354,In_2402,In_859);
nor U355 (N_355,In_2006,In_533);
xor U356 (N_356,In_1023,In_2379);
nand U357 (N_357,In_1513,In_236);
nor U358 (N_358,In_1450,In_1166);
or U359 (N_359,In_1997,In_1267);
nor U360 (N_360,In_934,In_2121);
xnor U361 (N_361,In_801,In_1987);
xor U362 (N_362,In_79,In_1526);
or U363 (N_363,In_838,In_2069);
nand U364 (N_364,In_2337,In_167);
nor U365 (N_365,In_2454,In_119);
nor U366 (N_366,In_1733,In_208);
or U367 (N_367,In_1071,In_1280);
or U368 (N_368,In_456,In_1259);
and U369 (N_369,In_2027,In_775);
xnor U370 (N_370,In_495,In_1005);
and U371 (N_371,In_2425,In_700);
nand U372 (N_372,In_2222,In_832);
or U373 (N_373,In_2355,In_301);
nor U374 (N_374,In_1535,In_532);
nor U375 (N_375,In_42,In_1065);
or U376 (N_376,In_1992,In_2328);
xnor U377 (N_377,In_821,In_1942);
or U378 (N_378,In_501,In_1179);
nand U379 (N_379,In_895,In_1946);
or U380 (N_380,In_2256,In_716);
and U381 (N_381,In_1306,In_155);
and U382 (N_382,In_546,In_2356);
nor U383 (N_383,In_1568,In_2113);
or U384 (N_384,In_815,In_2499);
nand U385 (N_385,In_203,In_105);
nor U386 (N_386,In_1497,In_901);
nor U387 (N_387,In_2415,In_283);
or U388 (N_388,In_382,In_2036);
xnor U389 (N_389,In_612,In_1345);
and U390 (N_390,In_2140,In_355);
and U391 (N_391,In_288,In_1040);
or U392 (N_392,In_498,In_848);
or U393 (N_393,In_2145,In_563);
or U394 (N_394,In_707,In_376);
or U395 (N_395,In_1270,In_1986);
nor U396 (N_396,In_1707,In_2141);
and U397 (N_397,In_125,In_1600);
and U398 (N_398,In_548,In_962);
nand U399 (N_399,In_602,In_2288);
nor U400 (N_400,In_2235,In_750);
nand U401 (N_401,In_2335,In_2292);
or U402 (N_402,In_2109,In_198);
nand U403 (N_403,In_384,In_1008);
or U404 (N_404,In_1767,In_1686);
or U405 (N_405,In_1333,In_386);
nand U406 (N_406,In_1309,In_1199);
and U407 (N_407,In_1645,In_1258);
and U408 (N_408,In_914,In_149);
or U409 (N_409,In_2332,In_2456);
xor U410 (N_410,In_1411,In_844);
and U411 (N_411,In_1807,In_114);
nor U412 (N_412,In_1195,In_1432);
xor U413 (N_413,In_1616,In_1740);
nand U414 (N_414,In_1349,In_1105);
nor U415 (N_415,In_357,In_411);
xnor U416 (N_416,In_2185,In_1756);
xnor U417 (N_417,In_536,In_661);
or U418 (N_418,In_1171,In_1024);
nor U419 (N_419,In_2270,In_1211);
and U420 (N_420,In_1873,In_1576);
and U421 (N_421,In_993,In_1393);
xor U422 (N_422,In_1833,In_1913);
nand U423 (N_423,In_1384,In_2391);
xor U424 (N_424,In_2338,In_1192);
or U425 (N_425,In_2171,In_517);
or U426 (N_426,In_1907,In_647);
xor U427 (N_427,In_1142,In_1569);
nand U428 (N_428,In_575,In_1629);
xor U429 (N_429,In_2253,In_606);
nor U430 (N_430,In_1176,In_1705);
or U431 (N_431,In_184,In_760);
xor U432 (N_432,In_1264,In_1013);
nor U433 (N_433,In_1665,In_307);
nand U434 (N_434,In_1173,In_985);
and U435 (N_435,In_2178,In_1504);
nor U436 (N_436,In_1474,In_1117);
nand U437 (N_437,In_1856,In_374);
nand U438 (N_438,In_537,In_1396);
or U439 (N_439,In_2067,In_2250);
nor U440 (N_440,In_542,In_2150);
or U441 (N_441,In_337,In_1620);
xnor U442 (N_442,In_2397,In_1961);
nand U443 (N_443,In_220,In_1870);
nor U444 (N_444,In_1364,In_1788);
nand U445 (N_445,In_1483,In_309);
nand U446 (N_446,In_1020,In_1471);
or U447 (N_447,In_1293,In_2377);
or U448 (N_448,In_923,In_1480);
and U449 (N_449,In_2214,In_1937);
and U450 (N_450,In_702,In_1979);
nor U451 (N_451,In_782,In_1978);
or U452 (N_452,In_480,In_80);
nand U453 (N_453,In_2289,In_215);
and U454 (N_454,In_353,In_1903);
xnor U455 (N_455,In_1633,In_1148);
xnor U456 (N_456,In_104,In_422);
nand U457 (N_457,In_494,In_1880);
xnor U458 (N_458,In_658,In_2419);
or U459 (N_459,In_115,In_1690);
and U460 (N_460,In_1635,In_319);
xor U461 (N_461,In_942,In_2417);
xor U462 (N_462,In_1263,In_1169);
nand U463 (N_463,In_1272,In_732);
nor U464 (N_464,In_1876,In_1375);
and U465 (N_465,In_1759,In_2101);
xor U466 (N_466,In_1582,In_375);
and U467 (N_467,In_512,In_250);
and U468 (N_468,In_1702,In_312);
nand U469 (N_469,In_530,In_974);
nand U470 (N_470,In_727,In_2280);
and U471 (N_471,In_600,In_294);
and U472 (N_472,In_1465,In_2072);
nand U473 (N_473,In_1892,In_85);
or U474 (N_474,In_550,In_2014);
nand U475 (N_475,In_2414,In_1524);
and U476 (N_476,In_302,In_2097);
and U477 (N_477,In_1799,In_1745);
or U478 (N_478,In_2325,In_182);
nand U479 (N_479,In_1960,In_153);
nand U480 (N_480,In_791,In_524);
nand U481 (N_481,In_688,In_749);
and U482 (N_482,In_2485,In_229);
or U483 (N_483,In_1681,In_648);
or U484 (N_484,In_756,In_1282);
and U485 (N_485,In_1409,In_15);
or U486 (N_486,In_1803,In_2293);
and U487 (N_487,In_2008,In_718);
nor U488 (N_488,In_1746,In_1405);
nand U489 (N_489,In_117,In_2398);
nor U490 (N_490,In_1610,In_1912);
xnor U491 (N_491,In_997,In_2411);
or U492 (N_492,In_673,In_1965);
nand U493 (N_493,In_641,In_1257);
nand U494 (N_494,In_432,In_1794);
nand U495 (N_495,In_2182,In_39);
nand U496 (N_496,In_194,In_2045);
xor U497 (N_497,In_219,In_728);
xnor U498 (N_498,In_240,In_982);
or U499 (N_499,In_1717,In_1284);
xor U500 (N_500,In_1922,N_371);
xnor U501 (N_501,N_53,In_1421);
nor U502 (N_502,N_463,In_2040);
and U503 (N_503,In_1044,In_920);
nor U504 (N_504,N_373,In_439);
nor U505 (N_505,In_861,In_1712);
nor U506 (N_506,N_251,N_8);
xnor U507 (N_507,In_2413,In_1824);
or U508 (N_508,In_1413,In_1326);
xnor U509 (N_509,In_163,In_1778);
and U510 (N_510,In_1575,N_174);
or U511 (N_511,In_1518,N_277);
and U512 (N_512,N_260,In_2223);
and U513 (N_513,In_1603,N_398);
xor U514 (N_514,In_120,In_694);
nand U515 (N_515,N_397,In_1360);
or U516 (N_516,In_1559,In_230);
or U517 (N_517,In_1750,In_1920);
or U518 (N_518,In_1444,In_2327);
nor U519 (N_519,In_466,N_129);
nand U520 (N_520,In_1063,In_2404);
or U521 (N_521,In_2220,In_1792);
nand U522 (N_522,In_1601,In_1651);
xor U523 (N_523,In_555,N_380);
or U524 (N_524,In_205,In_634);
xor U525 (N_525,N_135,In_1590);
nand U526 (N_526,In_1312,N_482);
xor U527 (N_527,In_2285,In_1921);
and U528 (N_528,In_1516,In_2431);
or U529 (N_529,N_175,In_351);
nor U530 (N_530,In_1037,In_1055);
nand U531 (N_531,In_1735,N_168);
and U532 (N_532,N_163,In_1990);
xnor U533 (N_533,In_253,In_892);
xnor U534 (N_534,In_1505,In_1408);
and U535 (N_535,N_75,In_2464);
nand U536 (N_536,In_1307,In_1014);
nand U537 (N_537,In_1704,In_17);
or U538 (N_538,N_451,In_1022);
xnor U539 (N_539,In_2031,In_2032);
xor U540 (N_540,In_1077,In_583);
nor U541 (N_541,In_1147,In_2147);
nor U542 (N_542,In_2459,N_471);
and U543 (N_543,N_423,In_1288);
and U544 (N_544,N_248,In_2122);
nor U545 (N_545,N_4,In_1027);
nand U546 (N_546,N_3,In_628);
and U547 (N_547,In_737,In_983);
xor U548 (N_548,In_836,N_491);
nor U549 (N_549,In_1047,In_2230);
nor U550 (N_550,N_191,In_1317);
or U551 (N_551,In_1589,N_70);
xor U552 (N_552,In_722,In_1101);
nand U553 (N_553,In_175,N_125);
nor U554 (N_554,In_1180,In_1006);
nor U555 (N_555,In_933,In_1538);
and U556 (N_556,In_632,N_473);
xor U557 (N_557,In_870,N_254);
or U558 (N_558,In_2168,In_1121);
or U559 (N_559,In_619,N_94);
and U560 (N_560,In_61,In_945);
and U561 (N_561,N_276,In_1881);
nor U562 (N_562,N_73,In_1917);
xor U563 (N_563,In_1925,In_388);
or U564 (N_564,In_1739,N_450);
xnor U565 (N_565,In_1763,In_50);
nand U566 (N_566,In_1018,In_368);
xnor U567 (N_567,N_384,N_332);
or U568 (N_568,In_1725,In_2202);
nor U569 (N_569,In_1943,In_2002);
nor U570 (N_570,In_879,In_316);
or U571 (N_571,In_2161,In_1175);
or U572 (N_572,In_1459,In_887);
and U573 (N_573,In_522,In_2482);
nand U574 (N_574,N_330,In_137);
xnor U575 (N_575,In_1177,In_342);
xor U576 (N_576,N_429,In_2169);
or U577 (N_577,In_2246,In_464);
nor U578 (N_578,In_1886,In_255);
or U579 (N_579,In_1028,In_674);
and U580 (N_580,In_690,In_1358);
xnor U581 (N_581,In_426,N_309);
nor U582 (N_582,In_493,In_2254);
and U583 (N_583,In_963,In_2180);
nand U584 (N_584,In_723,In_124);
nor U585 (N_585,N_15,In_1454);
xnor U586 (N_586,In_710,In_1999);
and U587 (N_587,In_1256,In_2311);
or U588 (N_588,In_2357,N_33);
and U589 (N_589,In_2077,In_618);
and U590 (N_590,In_1536,In_1529);
xnor U591 (N_591,In_1869,In_2382);
xor U592 (N_592,In_51,In_1201);
and U593 (N_593,N_123,N_498);
or U594 (N_594,N_150,In_959);
nor U595 (N_595,In_588,N_171);
nand U596 (N_596,In_1774,N_105);
and U597 (N_597,N_403,In_1722);
nor U598 (N_598,In_343,In_764);
nor U599 (N_599,N_472,In_1858);
and U600 (N_600,In_1410,In_590);
and U601 (N_601,In_313,In_99);
nand U602 (N_602,N_71,N_147);
nor U603 (N_603,In_1170,In_2215);
xor U604 (N_604,In_1525,In_558);
xnor U605 (N_605,In_965,In_1204);
nor U606 (N_606,In_1232,N_95);
xor U607 (N_607,N_385,In_2251);
xnor U608 (N_608,In_140,In_1052);
nor U609 (N_609,In_331,In_416);
nand U610 (N_610,N_149,N_300);
nor U611 (N_611,In_2361,In_805);
and U612 (N_612,In_88,In_93);
xor U613 (N_613,In_2389,In_562);
nor U614 (N_614,In_604,In_1508);
xor U615 (N_615,In_86,In_245);
or U616 (N_616,In_921,N_18);
nand U617 (N_617,In_831,In_421);
nand U618 (N_618,In_349,N_193);
and U619 (N_619,In_1479,In_2037);
and U620 (N_620,In_29,N_183);
and U621 (N_621,In_1094,In_90);
nor U622 (N_622,N_22,In_544);
nand U623 (N_623,In_1790,N_157);
nand U624 (N_624,N_418,N_112);
or U625 (N_625,N_90,In_1000);
nor U626 (N_626,In_896,N_389);
nor U627 (N_627,In_1064,In_2294);
nand U628 (N_628,In_944,In_1463);
and U629 (N_629,N_14,In_405);
nor U630 (N_630,In_2316,In_1470);
nand U631 (N_631,N_323,In_1808);
xor U632 (N_632,In_1887,N_424);
and U633 (N_633,N_360,In_172);
or U634 (N_634,In_2277,N_216);
nand U635 (N_635,In_2392,N_233);
and U636 (N_636,N_173,In_897);
xnor U637 (N_637,In_735,N_374);
nand U638 (N_638,In_2187,In_1036);
nand U639 (N_639,In_1510,In_2153);
nand U640 (N_640,N_227,In_1954);
nor U641 (N_641,N_228,N_270);
and U642 (N_642,In_2209,In_379);
nand U643 (N_643,In_2458,In_1163);
nor U644 (N_644,In_22,In_1819);
nor U645 (N_645,In_1738,N_203);
xnor U646 (N_646,In_325,N_92);
and U647 (N_647,In_2314,N_211);
nor U648 (N_648,N_42,In_564);
nand U649 (N_649,N_465,N_289);
nand U650 (N_650,In_2394,In_401);
nand U651 (N_651,In_565,In_482);
nor U652 (N_652,In_1955,In_1511);
xor U653 (N_653,In_1209,N_0);
and U654 (N_654,In_305,In_2176);
and U655 (N_655,In_378,In_1404);
nor U656 (N_656,In_1233,In_1025);
xor U657 (N_657,In_1391,In_1053);
nand U658 (N_658,In_1935,In_251);
nand U659 (N_659,In_360,In_1229);
nor U660 (N_660,N_292,N_479);
or U661 (N_661,N_232,N_43);
nand U662 (N_662,In_227,In_2081);
nor U663 (N_663,N_62,In_1972);
xnor U664 (N_664,In_1534,N_490);
or U665 (N_665,In_31,N_217);
nor U666 (N_666,In_2403,N_213);
nand U667 (N_667,In_1502,In_1153);
and U668 (N_668,In_486,In_2315);
xnor U669 (N_669,In_847,In_2324);
or U670 (N_670,N_151,In_2430);
or U671 (N_671,In_1560,N_31);
and U672 (N_672,In_1533,In_1433);
nor U673 (N_673,In_1491,In_2044);
nor U674 (N_674,In_763,N_148);
nor U675 (N_675,In_885,In_1485);
nor U676 (N_676,In_1109,N_422);
and U677 (N_677,In_925,In_1553);
or U678 (N_678,N_342,N_72);
nor U679 (N_679,In_1674,N_59);
or U680 (N_680,In_1944,In_2117);
xor U681 (N_681,In_1838,N_107);
nand U682 (N_682,In_394,In_2434);
or U683 (N_683,In_1985,In_2074);
nand U684 (N_684,In_603,In_911);
xor U685 (N_685,In_1904,In_2175);
or U686 (N_686,In_2263,In_873);
or U687 (N_687,In_601,In_845);
nand U688 (N_688,In_32,In_1058);
xnor U689 (N_689,N_468,N_156);
and U690 (N_690,N_29,In_1236);
nor U691 (N_691,In_2481,In_754);
nand U692 (N_692,In_2165,N_268);
or U693 (N_693,In_2156,In_1563);
or U694 (N_694,N_453,In_1087);
and U695 (N_695,N_396,In_677);
xnor U696 (N_696,In_1578,N_154);
and U697 (N_697,In_1303,In_1420);
and U698 (N_698,In_1068,In_668);
or U699 (N_699,In_2385,N_136);
xor U700 (N_700,In_527,In_366);
or U701 (N_701,In_1120,In_1350);
nand U702 (N_702,N_290,In_18);
xor U703 (N_703,In_1464,N_200);
xnor U704 (N_704,In_1968,N_339);
or U705 (N_705,In_1468,In_1766);
and U706 (N_706,In_1801,In_783);
or U707 (N_707,In_1714,N_426);
xnor U708 (N_708,In_1390,In_1519);
nand U709 (N_709,In_2271,In_2433);
nor U710 (N_710,In_1812,In_256);
or U711 (N_711,In_453,In_1947);
or U712 (N_712,In_1606,In_905);
and U713 (N_713,N_476,N_229);
nor U714 (N_714,In_1729,In_1133);
and U715 (N_715,In_1872,In_1496);
or U716 (N_716,In_1755,N_57);
nor U717 (N_717,N_131,N_340);
or U718 (N_718,N_40,N_264);
or U719 (N_719,In_1980,In_743);
xnor U720 (N_720,In_701,N_34);
nand U721 (N_721,N_88,In_731);
nand U722 (N_722,In_2115,N_307);
nand U723 (N_723,In_2016,In_1030);
nor U724 (N_724,In_1728,N_122);
or U725 (N_725,In_2095,N_399);
nor U726 (N_726,N_314,In_1495);
nor U727 (N_727,N_431,N_357);
and U728 (N_728,In_587,In_287);
xor U729 (N_729,In_1098,N_395);
or U730 (N_730,In_1313,In_2058);
nor U731 (N_731,In_1641,In_2358);
nand U732 (N_732,In_2078,In_2435);
xnor U733 (N_733,In_2019,In_1793);
or U734 (N_734,In_2205,In_521);
or U735 (N_735,N_402,In_936);
and U736 (N_736,N_142,In_1060);
nand U737 (N_737,In_373,In_169);
and U738 (N_738,In_36,In_1048);
nor U739 (N_739,In_1977,In_649);
nor U740 (N_740,In_1135,In_2418);
or U741 (N_741,In_627,In_171);
and U742 (N_742,In_797,N_116);
and U743 (N_743,In_928,N_444);
and U744 (N_744,In_1918,N_81);
or U745 (N_745,In_2075,N_89);
nand U746 (N_746,In_1566,In_469);
nor U747 (N_747,In_717,In_576);
xnor U748 (N_748,In_1145,N_298);
nand U749 (N_749,N_492,In_2313);
xnor U750 (N_750,N_489,In_1066);
xnor U751 (N_751,In_57,In_643);
or U752 (N_752,In_1295,N_114);
nand U753 (N_753,In_903,In_400);
nor U754 (N_754,In_1351,In_2062);
xor U755 (N_755,In_2305,In_2054);
xnor U756 (N_756,N_419,In_1298);
xor U757 (N_757,In_1785,In_784);
nor U758 (N_758,In_1181,In_940);
xor U759 (N_759,N_182,In_777);
and U760 (N_760,N_82,In_2090);
xnor U761 (N_761,In_476,In_1178);
xnor U762 (N_762,In_2204,In_1314);
nand U763 (N_763,In_2494,In_2445);
nand U764 (N_764,N_359,In_956);
and U765 (N_765,In_2440,In_2279);
or U766 (N_766,N_153,In_856);
xor U767 (N_767,In_769,In_556);
nand U768 (N_768,In_1128,N_198);
nor U769 (N_769,In_2307,In_1855);
xnor U770 (N_770,In_506,N_2);
or U771 (N_771,In_582,In_1572);
nor U772 (N_772,In_580,N_10);
nor U773 (N_773,N_325,In_1655);
nand U774 (N_774,In_881,In_1896);
and U775 (N_775,In_381,In_615);
nand U776 (N_776,In_1218,N_145);
and U777 (N_777,In_1189,N_108);
and U778 (N_778,In_2136,In_1034);
or U779 (N_779,In_2387,N_212);
xnor U780 (N_780,In_2333,In_922);
and U781 (N_781,In_2410,In_2272);
and U782 (N_782,In_2334,In_2056);
nor U783 (N_783,In_1835,N_343);
or U784 (N_784,N_361,In_491);
nand U785 (N_785,N_138,In_1754);
nand U786 (N_786,In_1860,In_1662);
xor U787 (N_787,In_2238,In_383);
or U788 (N_788,In_118,In_721);
nor U789 (N_789,In_161,N_341);
nand U790 (N_790,N_446,In_1266);
nor U791 (N_791,N_192,In_371);
or U792 (N_792,In_1073,In_2472);
nand U793 (N_793,N_141,N_127);
nor U794 (N_794,In_1096,In_631);
nor U795 (N_795,In_698,N_364);
xnor U796 (N_796,In_1129,In_296);
or U797 (N_797,In_758,In_20);
nand U798 (N_798,In_581,In_1764);
xor U799 (N_799,In_1286,In_1866);
nor U800 (N_800,In_291,In_1049);
or U801 (N_801,In_882,N_274);
or U802 (N_802,N_261,N_181);
or U803 (N_803,N_35,In_455);
nor U804 (N_804,In_97,In_1203);
and U805 (N_805,In_300,N_180);
and U806 (N_806,N_285,N_409);
nor U807 (N_807,In_1446,In_650);
nor U808 (N_808,N_76,In_868);
nand U809 (N_809,In_1346,N_86);
or U810 (N_810,N_199,In_1650);
xnor U811 (N_811,In_237,In_1597);
xnor U812 (N_812,N_293,N_144);
nand U813 (N_813,In_1342,In_1624);
nand U814 (N_814,In_2336,N_338);
or U815 (N_815,In_181,In_912);
nor U816 (N_816,In_511,In_2342);
nand U817 (N_817,In_2119,In_1561);
nor U818 (N_818,N_470,In_1752);
or U819 (N_819,N_235,In_1777);
or U820 (N_820,N_414,In_1299);
xnor U821 (N_821,In_1152,N_126);
xnor U822 (N_822,In_289,In_2170);
nand U823 (N_823,N_449,N_39);
nor U824 (N_824,In_855,N_170);
or U825 (N_825,In_2479,N_80);
xor U826 (N_826,In_2226,In_1730);
and U827 (N_827,In_1216,In_92);
and U828 (N_828,In_1234,N_255);
xor U829 (N_829,N_115,N_495);
nand U830 (N_830,In_1619,In_2051);
nor U831 (N_831,N_178,In_2368);
nand U832 (N_832,In_759,In_336);
and U833 (N_833,N_282,N_47);
nor U834 (N_834,N_329,N_258);
or U835 (N_835,In_1614,In_776);
nor U836 (N_836,N_321,In_77);
xor U837 (N_837,N_45,In_538);
nand U838 (N_838,N_425,In_1235);
nor U839 (N_839,In_1796,N_30);
and U840 (N_840,In_960,In_744);
or U841 (N_841,In_2426,In_2229);
nand U842 (N_842,N_334,In_2018);
xnor U843 (N_843,In_2441,N_328);
nor U844 (N_844,N_372,N_382);
xor U845 (N_845,In_2453,In_1249);
and U846 (N_846,In_1677,N_64);
and U847 (N_847,In_398,In_1632);
or U848 (N_848,In_2064,In_151);
xor U849 (N_849,In_1623,In_509);
xor U850 (N_850,In_1543,In_404);
nand U851 (N_851,In_927,In_415);
nand U852 (N_852,N_185,In_1928);
nor U853 (N_853,N_46,In_893);
or U854 (N_854,In_703,In_223);
nand U855 (N_855,In_2498,In_1431);
xor U856 (N_856,In_1311,In_102);
xnor U857 (N_857,In_2468,In_1430);
or U858 (N_858,In_516,In_264);
or U859 (N_859,In_876,N_120);
nor U860 (N_860,In_459,N_331);
or U861 (N_861,In_293,N_317);
nor U862 (N_862,N_177,N_462);
or U863 (N_863,In_621,N_240);
nor U864 (N_864,In_1119,In_406);
nand U865 (N_865,In_2087,In_1456);
nor U866 (N_866,In_1452,N_100);
or U867 (N_867,N_326,N_480);
and U868 (N_868,N_99,In_742);
xor U869 (N_869,In_1281,In_54);
xor U870 (N_870,In_441,In_1771);
nand U871 (N_871,In_1841,In_1970);
and U872 (N_872,N_188,In_1252);
or U873 (N_873,N_390,In_2203);
xnor U874 (N_874,In_794,In_1998);
or U875 (N_875,In_1207,In_595);
or U876 (N_876,In_596,In_724);
nand U877 (N_877,N_190,In_1213);
nor U878 (N_878,In_1164,In_2319);
xnor U879 (N_879,In_1613,In_431);
nand U880 (N_880,In_1924,In_350);
and U881 (N_881,N_124,In_2290);
xnor U882 (N_882,N_351,In_2340);
xnor U883 (N_883,In_814,In_1275);
xor U884 (N_884,In_1933,In_2341);
xor U885 (N_885,In_2378,In_1584);
nor U886 (N_886,In_1902,In_2042);
nor U887 (N_887,In_825,N_486);
xor U888 (N_888,N_101,In_1734);
or U889 (N_889,In_318,In_1874);
xor U890 (N_890,In_1744,In_1622);
xor U891 (N_891,In_1697,In_1184);
or U892 (N_892,In_1374,In_559);
nand U893 (N_893,In_204,In_1809);
and U894 (N_894,In_799,In_1085);
nand U895 (N_895,In_551,In_910);
nand U896 (N_896,N_222,In_242);
or U897 (N_897,N_244,In_761);
nand U898 (N_898,In_1825,In_1546);
or U899 (N_899,In_1644,In_2135);
xor U900 (N_900,In_833,In_1676);
and U901 (N_901,N_162,In_637);
nor U902 (N_902,In_315,In_579);
and U903 (N_903,N_455,In_1571);
nor U904 (N_904,N_60,In_1208);
nor U905 (N_905,In_938,In_980);
nor U906 (N_906,N_379,In_1915);
xnor U907 (N_907,N_369,In_2012);
nor U908 (N_908,N_9,In_1828);
xnor U909 (N_909,In_973,In_858);
or U910 (N_910,N_301,In_2354);
nor U911 (N_911,N_25,In_1401);
xnor U912 (N_912,N_78,In_816);
and U913 (N_913,N_243,In_1155);
xor U914 (N_914,In_2363,In_884);
nor U915 (N_915,In_1517,In_686);
nor U916 (N_916,In_1325,N_494);
nor U917 (N_917,N_54,In_310);
xnor U918 (N_918,N_336,N_237);
and U919 (N_919,N_269,In_152);
or U920 (N_920,N_437,In_2302);
xnor U921 (N_921,In_2192,In_2071);
nor U922 (N_922,In_569,In_1161);
xnor U923 (N_923,N_85,In_1982);
or U924 (N_924,N_275,In_460);
or U925 (N_925,In_273,In_2396);
or U926 (N_926,In_1910,N_291);
or U927 (N_927,In_333,N_103);
xnor U928 (N_928,N_302,N_420);
xor U929 (N_929,N_165,In_2451);
nand U930 (N_930,N_224,In_2149);
nand U931 (N_931,N_111,In_1279);
or U932 (N_932,In_1605,N_348);
or U933 (N_933,In_2026,In_359);
and U934 (N_934,In_1737,In_2219);
xor U935 (N_935,In_187,In_1742);
and U936 (N_936,In_275,In_1557);
or U937 (N_937,In_1908,In_578);
nor U938 (N_938,N_195,In_191);
xor U939 (N_939,In_1244,N_172);
nand U940 (N_940,In_311,In_1648);
nor U941 (N_941,In_10,In_765);
xor U942 (N_942,In_367,N_404);
nor U943 (N_943,N_353,In_238);
xor U944 (N_944,In_755,N_27);
or U945 (N_945,In_285,In_1196);
nand U946 (N_946,In_585,In_2422);
or U947 (N_947,N_143,In_1223);
nor U948 (N_948,In_395,In_689);
or U949 (N_949,In_663,In_695);
xnor U950 (N_950,In_733,In_1512);
xor U951 (N_951,In_434,N_355);
and U952 (N_952,In_369,N_169);
xor U953 (N_953,In_1072,In_1156);
and U954 (N_954,In_2183,In_2099);
nand U955 (N_955,In_2106,In_1157);
xnor U956 (N_956,In_729,In_1929);
or U957 (N_957,N_393,In_47);
nor U958 (N_958,In_409,N_466);
or U959 (N_959,In_65,In_620);
or U960 (N_960,In_638,In_2105);
xor U961 (N_961,In_2123,In_2301);
nor U962 (N_962,N_335,In_1089);
and U963 (N_963,In_1132,In_1687);
and U964 (N_964,In_852,In_1940);
nor U965 (N_965,In_419,In_1467);
or U966 (N_966,N_412,In_802);
nor U967 (N_967,N_405,In_1079);
and U968 (N_968,N_324,In_2291);
nor U969 (N_969,In_1268,In_2473);
or U970 (N_970,N_7,N_262);
xnor U971 (N_971,N_263,In_1523);
nor U972 (N_972,In_1673,N_21);
nor U973 (N_973,In_1611,In_2461);
and U974 (N_974,N_249,In_2242);
nor U975 (N_975,N_102,In_2094);
nor U976 (N_976,N_176,In_1438);
xor U977 (N_977,In_109,In_2343);
or U978 (N_978,In_860,In_1365);
nand U979 (N_979,N_223,N_134);
nor U980 (N_980,In_1251,In_2349);
and U981 (N_981,N_375,In_260);
xor U982 (N_982,N_84,In_1224);
xor U983 (N_983,In_826,In_2241);
or U984 (N_984,N_474,In_1357);
xnor U985 (N_985,In_671,In_513);
or U986 (N_986,In_499,In_1017);
xnor U987 (N_987,In_1528,In_226);
and U988 (N_988,In_828,In_1906);
nor U989 (N_989,In_1137,N_488);
nand U990 (N_990,In_279,N_297);
and U991 (N_991,N_306,N_58);
or U992 (N_992,In_827,N_295);
or U993 (N_993,N_443,N_284);
nor U994 (N_994,N_352,In_1829);
nand U995 (N_995,N_97,In_2211);
xor U996 (N_996,N_256,In_282);
xor U997 (N_997,In_2350,In_1090);
nor U998 (N_998,In_244,In_2286);
or U999 (N_999,In_1277,In_804);
nand U1000 (N_1000,N_347,In_566);
nand U1001 (N_1001,In_1436,In_110);
nor U1002 (N_1002,N_823,In_1032);
xor U1003 (N_1003,N_726,N_522);
and U1004 (N_1004,In_345,N_536);
nor U1005 (N_1005,N_904,In_450);
nor U1006 (N_1006,N_572,In_1675);
and U1007 (N_1007,In_1445,N_775);
nand U1008 (N_1008,N_531,In_437);
xor U1009 (N_1009,In_98,N_847);
nor U1010 (N_1010,In_2225,N_744);
or U1011 (N_1011,N_721,In_540);
or U1012 (N_1012,In_1822,N_960);
or U1013 (N_1013,In_2239,N_320);
nand U1014 (N_1014,N_219,N_500);
xnor U1015 (N_1015,N_499,N_570);
nor U1016 (N_1016,In_2114,N_523);
xor U1017 (N_1017,In_1573,N_786);
nor U1018 (N_1018,In_2466,In_535);
xor U1019 (N_1019,In_1056,N_152);
or U1020 (N_1020,In_1919,In_1016);
xnor U1021 (N_1021,N_906,N_954);
and U1022 (N_1022,N_825,In_773);
nor U1023 (N_1023,N_247,In_1836);
or U1024 (N_1024,N_601,In_84);
and U1025 (N_1025,N_857,In_1283);
nor U1026 (N_1026,In_154,In_1530);
nor U1027 (N_1027,N_615,In_214);
nand U1028 (N_1028,N_848,In_397);
nand U1029 (N_1029,N_879,N_680);
nand U1030 (N_1030,In_1494,In_2060);
and U1031 (N_1031,N_484,N_666);
or U1032 (N_1032,In_1594,N_877);
nor U1033 (N_1033,N_581,In_2007);
nand U1034 (N_1034,In_1883,N_106);
and U1035 (N_1035,In_2348,In_526);
or U1036 (N_1036,In_2070,In_2091);
nor U1037 (N_1037,In_636,N_635);
nand U1038 (N_1038,N_901,N_349);
and U1039 (N_1039,N_436,In_1743);
and U1040 (N_1040,In_745,In_2061);
or U1041 (N_1041,N_984,In_1679);
nand U1042 (N_1042,In_573,In_902);
and U1043 (N_1043,In_613,In_1033);
nor U1044 (N_1044,N_435,In_1909);
nand U1045 (N_1045,In_387,In_753);
and U1046 (N_1046,In_1212,In_2133);
nand U1047 (N_1047,N_731,N_515);
or U1048 (N_1048,In_685,N_132);
or U1049 (N_1049,N_741,In_297);
nand U1050 (N_1050,N_752,N_505);
nand U1051 (N_1051,In_639,N_571);
and U1052 (N_1052,In_1150,N_83);
and U1053 (N_1053,N_678,N_839);
nand U1054 (N_1054,N_445,N_316);
nand U1055 (N_1055,In_2221,N_808);
nor U1056 (N_1056,N_66,N_591);
nor U1057 (N_1057,N_118,N_638);
or U1058 (N_1058,In_467,In_1706);
xnor U1059 (N_1059,In_101,N_713);
or U1060 (N_1060,In_915,In_2383);
and U1061 (N_1061,In_75,In_1932);
nand U1062 (N_1062,In_158,N_345);
nand U1063 (N_1063,In_796,N_773);
and U1064 (N_1064,In_725,N_861);
nand U1065 (N_1065,N_506,In_772);
or U1066 (N_1066,In_445,N_947);
and U1067 (N_1067,N_207,N_159);
nand U1068 (N_1068,N_642,In_1643);
nor U1069 (N_1069,N_133,In_1242);
xnor U1070 (N_1070,N_485,N_995);
nand U1071 (N_1071,N_179,N_986);
nor U1072 (N_1072,N_377,N_831);
nor U1073 (N_1073,In_341,In_880);
or U1074 (N_1074,N_599,In_1827);
nand U1075 (N_1075,N_777,In_966);
nor U1076 (N_1076,N_951,In_2053);
xor U1077 (N_1077,N_612,N_434);
and U1078 (N_1078,N_755,N_551);
nor U1079 (N_1079,N_630,In_423);
xor U1080 (N_1080,N_356,N_860);
or U1081 (N_1081,N_734,N_559);
xor U1082 (N_1082,N_502,In_611);
xnor U1083 (N_1083,N_368,In_1088);
or U1084 (N_1084,N_23,In_1877);
xnor U1085 (N_1085,In_837,N_793);
nor U1086 (N_1086,N_366,In_2463);
nand U1087 (N_1087,In_2052,N_272);
or U1088 (N_1088,N_584,N_613);
nand U1089 (N_1089,In_2049,In_1897);
and U1090 (N_1090,N_664,In_1716);
and U1091 (N_1091,In_1693,In_2158);
xor U1092 (N_1092,N_703,N_924);
nand U1093 (N_1093,N_641,In_918);
nand U1094 (N_1094,In_820,N_487);
nand U1095 (N_1095,In_2353,N_707);
and U1096 (N_1096,N_273,N_433);
and U1097 (N_1097,In_1514,In_785);
and U1098 (N_1098,N_299,In_168);
nand U1099 (N_1099,N_442,N_759);
and U1100 (N_1100,N_563,N_130);
or U1101 (N_1101,N_819,In_1621);
nand U1102 (N_1102,In_2484,N_892);
or U1103 (N_1103,N_668,N_381);
xor U1104 (N_1104,In_2407,In_2401);
and U1105 (N_1105,N_952,N_874);
or U1106 (N_1106,In_1075,In_2287);
or U1107 (N_1107,N_626,In_1130);
nand U1108 (N_1108,N_113,In_2098);
nand U1109 (N_1109,N_929,In_435);
nor U1110 (N_1110,N_996,N_253);
xor U1111 (N_1111,N_187,N_729);
nand U1112 (N_1112,In_160,N_985);
and U1113 (N_1113,In_1762,In_2351);
nor U1114 (N_1114,In_48,N_911);
and U1115 (N_1115,N_700,In_552);
nor U1116 (N_1116,In_1787,In_1352);
nand U1117 (N_1117,In_1839,In_800);
nand U1118 (N_1118,In_2096,In_447);
nor U1119 (N_1119,N_849,N_236);
nor U1120 (N_1120,N_779,N_870);
xnor U1121 (N_1121,In_979,In_1289);
and U1122 (N_1122,In_206,In_1751);
nand U1123 (N_1123,N_587,N_413);
xor U1124 (N_1124,In_1574,N_257);
xor U1125 (N_1125,In_1627,In_1012);
and U1126 (N_1126,N_851,In_990);
nor U1127 (N_1127,N_955,N_979);
nand U1128 (N_1128,In_1736,In_705);
or U1129 (N_1129,N_681,In_1422);
nor U1130 (N_1130,In_812,N_971);
nand U1131 (N_1131,In_248,N_313);
nand U1132 (N_1132,In_139,In_1637);
or U1133 (N_1133,N_166,N_578);
xnor U1134 (N_1134,N_844,In_715);
nand U1135 (N_1135,N_765,In_202);
or U1136 (N_1136,In_1138,In_1197);
or U1137 (N_1137,N_394,In_1136);
nor U1138 (N_1138,In_916,N_427);
nor U1139 (N_1139,In_16,In_298);
or U1140 (N_1140,In_1031,N_811);
or U1141 (N_1141,N_600,In_1853);
nor U1142 (N_1142,N_525,N_990);
nand U1143 (N_1143,In_1002,In_1386);
nor U1144 (N_1144,In_878,In_534);
xor U1145 (N_1145,N_890,In_2367);
or U1146 (N_1146,In_258,N_876);
nor U1147 (N_1147,N_575,In_2129);
nand U1148 (N_1148,N_843,In_811);
and U1149 (N_1149,N_961,N_628);
or U1150 (N_1150,N_197,In_1434);
xnor U1151 (N_1151,In_1466,In_1580);
xnor U1152 (N_1152,N_68,N_866);
and U1153 (N_1153,In_557,N_467);
nand U1154 (N_1154,N_5,N_854);
or U1155 (N_1155,N_754,In_757);
nor U1156 (N_1156,In_186,In_871);
nand U1157 (N_1157,N_576,N_458);
and U1158 (N_1158,N_496,N_746);
nand U1159 (N_1159,In_2312,N_712);
and U1160 (N_1160,In_1010,N_319);
and U1161 (N_1161,In_2318,N_205);
nand U1162 (N_1162,N_519,N_383);
xor U1163 (N_1163,In_961,In_1952);
xnor U1164 (N_1164,N_999,N_362);
nand U1165 (N_1165,N_546,N_736);
nor U1166 (N_1166,N_288,In_779);
nand U1167 (N_1167,N_764,N_12);
nor U1168 (N_1168,In_2283,In_1400);
nand U1169 (N_1169,N_931,In_823);
nor U1170 (N_1170,N_430,N_271);
and U1171 (N_1171,N_421,In_1815);
nand U1172 (N_1172,N_659,In_2111);
or U1173 (N_1173,In_2208,In_1837);
and U1174 (N_1174,In_971,In_2366);
xnor U1175 (N_1175,In_207,In_2191);
nor U1176 (N_1176,In_503,In_1134);
or U1177 (N_1177,In_2446,In_1361);
or U1178 (N_1178,In_1581,N_675);
nand U1179 (N_1179,N_747,N_894);
nor U1180 (N_1180,N_944,In_1779);
nand U1181 (N_1181,N_883,In_74);
xor U1182 (N_1182,N_927,In_1719);
or U1183 (N_1183,N_327,In_1154);
or U1184 (N_1184,N_805,N_303);
or U1185 (N_1185,In_1247,N_189);
or U1186 (N_1186,N_246,In_1338);
nor U1187 (N_1187,N_975,In_1294);
and U1188 (N_1188,N_834,In_1389);
nand U1189 (N_1189,N_508,In_2443);
or U1190 (N_1190,N_11,In_1784);
nand U1191 (N_1191,N_1,N_702);
nand U1192 (N_1192,In_2495,In_987);
and U1193 (N_1193,N_616,In_209);
nor U1194 (N_1194,In_71,N_521);
xor U1195 (N_1195,In_1631,N_650);
nand U1196 (N_1196,N_676,N_912);
xor U1197 (N_1197,In_1948,In_1395);
xnor U1198 (N_1198,In_1634,N_687);
or U1199 (N_1199,N_619,In_2116);
or U1200 (N_1200,N_459,In_1387);
and U1201 (N_1201,N_921,N_852);
nand U1202 (N_1202,In_1958,N_724);
nor U1203 (N_1203,In_1107,In_2030);
nand U1204 (N_1204,N_534,In_142);
xnor U1205 (N_1205,N_908,In_854);
nor U1206 (N_1206,In_906,N_810);
xor U1207 (N_1207,N_873,In_709);
or U1208 (N_1208,In_1931,N_509);
and U1209 (N_1209,In_2489,In_1851);
nand U1210 (N_1210,N_225,In_2196);
or U1211 (N_1211,In_2197,In_106);
nand U1212 (N_1212,N_517,In_385);
xor U1213 (N_1213,In_2231,In_170);
and U1214 (N_1214,N_477,N_943);
nor U1215 (N_1215,N_202,In_1683);
or U1216 (N_1216,N_310,N_717);
xor U1217 (N_1217,In_2450,In_1905);
nand U1218 (N_1218,N_527,N_750);
and U1219 (N_1219,N_915,In_2029);
nand U1220 (N_1220,In_91,N_620);
and U1221 (N_1221,In_1290,N_910);
nand U1222 (N_1222,N_751,N_41);
nand U1223 (N_1223,N_829,In_178);
nor U1224 (N_1224,N_830,In_55);
or U1225 (N_1225,In_609,N_855);
nand U1226 (N_1226,In_1585,In_133);
and U1227 (N_1227,N_514,In_413);
nor U1228 (N_1228,In_1639,N_816);
xnor U1229 (N_1229,In_2362,N_417);
nor U1230 (N_1230,N_428,In_680);
nand U1231 (N_1231,N_914,In_370);
nor U1232 (N_1232,N_19,N_65);
and U1233 (N_1233,N_588,N_631);
and U1234 (N_1234,In_964,N_464);
nand U1235 (N_1235,N_761,In_1823);
nor U1236 (N_1236,In_2372,N_63);
nor U1237 (N_1237,In_591,In_1372);
and U1238 (N_1238,N_590,In_1123);
xor U1239 (N_1239,In_888,In_1500);
xnor U1240 (N_1240,In_1515,N_441);
xor U1241 (N_1241,N_37,In_1891);
or U1242 (N_1242,N_714,N_561);
xor U1243 (N_1243,N_573,In_324);
nor U1244 (N_1244,N_940,N_722);
and U1245 (N_1245,N_812,In_2083);
nor U1246 (N_1246,In_1964,In_1070);
or U1247 (N_1247,In_2249,N_26);
nor U1248 (N_1248,In_1356,In_1640);
and U1249 (N_1249,In_529,N_137);
nand U1250 (N_1250,N_732,In_1301);
or U1251 (N_1251,In_2212,N_611);
and U1252 (N_1252,N_555,In_655);
xnor U1253 (N_1253,N_391,N_842);
xnor U1254 (N_1254,In_2339,N_448);
or U1255 (N_1255,In_1531,In_572);
nor U1256 (N_1256,In_427,In_1074);
and U1257 (N_1257,N_524,In_2416);
nor U1258 (N_1258,In_519,N_735);
xnor U1259 (N_1259,In_34,N_828);
nor U1260 (N_1260,N_949,N_540);
or U1261 (N_1261,In_1852,N_32);
xnor U1262 (N_1262,In_1167,In_1323);
or U1263 (N_1263,In_1680,N_778);
nand U1264 (N_1264,N_608,N_685);
nor U1265 (N_1265,N_574,In_1086);
nor U1266 (N_1266,In_1857,In_44);
or U1267 (N_1267,In_2193,N_920);
xnor U1268 (N_1268,N_926,N_406);
nand U1269 (N_1269,N_96,N_556);
xor U1270 (N_1270,N_880,In_1776);
nand U1271 (N_1271,In_1305,N_817);
xor U1272 (N_1272,N_392,In_665);
and U1273 (N_1273,In_539,In_43);
or U1274 (N_1274,N_91,N_932);
nand U1275 (N_1275,In_1667,N_942);
nor U1276 (N_1276,N_386,In_953);
xnor U1277 (N_1277,N_796,In_951);
and U1278 (N_1278,N_800,In_1938);
nand U1279 (N_1279,In_594,In_1608);
nand U1280 (N_1280,In_1127,N_684);
or U1281 (N_1281,N_739,In_320);
xnor U1282 (N_1282,In_408,In_574);
nor U1283 (N_1283,N_543,In_787);
and U1284 (N_1284,In_2043,In_713);
nand U1285 (N_1285,In_2442,N_312);
nand U1286 (N_1286,N_79,N_740);
and U1287 (N_1287,N_806,In_692);
xor U1288 (N_1288,In_835,In_1043);
xnor U1289 (N_1289,In_362,In_1800);
and U1290 (N_1290,In_159,N_48);
and U1291 (N_1291,N_452,N_715);
and U1292 (N_1292,N_51,N_503);
xnor U1293 (N_1293,N_585,N_267);
xor U1294 (N_1294,In_59,N_801);
nor U1295 (N_1295,In_492,N_973);
and U1296 (N_1296,In_33,N_28);
xor U1297 (N_1297,In_666,In_1656);
nand U1298 (N_1298,N_965,In_303);
and U1299 (N_1299,N_938,In_2423);
or U1300 (N_1300,In_1522,In_948);
nand U1301 (N_1301,N_286,N_322);
xnor U1302 (N_1302,In_872,N_989);
nor U1303 (N_1303,In_270,In_46);
xor U1304 (N_1304,N_758,In_2266);
or U1305 (N_1305,N_544,N_586);
xnor U1306 (N_1306,N_461,In_949);
or U1307 (N_1307,N_841,In_1769);
and U1308 (N_1308,In_1899,In_2243);
or U1309 (N_1309,In_1670,N_896);
and U1310 (N_1310,In_2041,In_347);
xnor U1311 (N_1311,In_70,In_1160);
nand U1312 (N_1312,N_533,N_835);
or U1313 (N_1313,N_520,N_696);
and U1314 (N_1314,In_1353,N_913);
nand U1315 (N_1315,N_69,N_776);
or U1316 (N_1316,N_743,In_485);
or U1317 (N_1317,In_1185,In_1443);
nand U1318 (N_1318,N_250,In_696);
or U1319 (N_1319,N_532,N_408);
xor U1320 (N_1320,N_770,In_2275);
nor U1321 (N_1321,In_1596,In_438);
xnor U1322 (N_1322,In_2344,N_958);
nand U1323 (N_1323,In_1310,N_206);
nand U1324 (N_1324,N_992,N_560);
and U1325 (N_1325,In_2321,In_2262);
xnor U1326 (N_1326,N_218,N_538);
and U1327 (N_1327,In_1551,N_226);
or U1328 (N_1328,N_121,N_569);
and U1329 (N_1329,In_659,N_558);
xnor U1330 (N_1330,In_998,In_930);
nand U1331 (N_1331,N_662,In_1957);
nand U1332 (N_1332,N_160,In_1371);
nor U1333 (N_1333,In_586,In_478);
and U1334 (N_1334,In_262,N_695);
and U1335 (N_1335,In_1427,N_826);
or U1336 (N_1336,N_647,N_606);
and U1337 (N_1337,N_833,In_984);
xnor U1338 (N_1338,In_1035,N_629);
nand U1339 (N_1339,N_541,In_2477);
nand U1340 (N_1340,In_402,In_2282);
xor U1341 (N_1341,In_2421,In_442);
and U1342 (N_1342,In_2033,N_748);
nand U1343 (N_1343,In_216,N_67);
nor U1344 (N_1344,In_1329,N_867);
nand U1345 (N_1345,In_176,In_867);
xor U1346 (N_1346,In_2359,N_771);
or U1347 (N_1347,N_279,N_974);
nor U1348 (N_1348,In_211,N_354);
and U1349 (N_1349,N_832,N_858);
and U1350 (N_1350,N_194,In_1370);
or U1351 (N_1351,In_2265,In_354);
nand U1352 (N_1352,In_1174,In_111);
nand U1353 (N_1353,In_1916,In_869);
nand U1354 (N_1354,N_644,N_956);
nor U1355 (N_1355,N_311,In_1765);
nand U1356 (N_1356,N_201,N_692);
nor U1357 (N_1357,In_1671,N_557);
xnor U1358 (N_1358,In_1893,N_481);
or U1359 (N_1359,In_274,N_110);
nor U1360 (N_1360,In_165,N_234);
nand U1361 (N_1361,N_643,N_663);
or U1362 (N_1362,In_1558,N_850);
or U1363 (N_1363,N_547,In_1599);
nand U1364 (N_1364,N_737,In_2003);
nand U1365 (N_1365,N_497,In_474);
and U1366 (N_1366,In_8,N_807);
nand U1367 (N_1367,N_987,N_566);
xor U1368 (N_1368,In_1045,In_2184);
xor U1369 (N_1369,N_769,In_2210);
nor U1370 (N_1370,N_836,N_649);
or U1371 (N_1371,In_1715,In_1962);
or U1372 (N_1372,N_780,N_457);
nand U1373 (N_1373,N_903,N_792);
or U1374 (N_1374,In_657,In_2462);
nor U1375 (N_1375,N_885,In_1449);
and U1376 (N_1376,In_263,N_526);
nand U1377 (N_1377,In_461,In_41);
and U1378 (N_1378,In_2055,In_1911);
nand U1379 (N_1379,In_1727,In_567);
or U1380 (N_1380,In_2428,In_813);
or U1381 (N_1381,N_607,In_150);
and U1382 (N_1382,N_797,In_803);
xor U1383 (N_1383,In_1222,In_1355);
xnor U1384 (N_1384,In_2257,In_1598);
nor U1385 (N_1385,In_100,In_2480);
and U1386 (N_1386,In_2024,N_672);
or U1387 (N_1387,In_2126,N_241);
nand U1388 (N_1388,In_304,In_1226);
nor U1389 (N_1389,In_2384,In_1814);
and U1390 (N_1390,In_197,N_953);
xnor U1391 (N_1391,N_919,N_632);
or U1392 (N_1392,N_596,In_1682);
nand U1393 (N_1393,N_475,In_299);
or U1394 (N_1394,In_1761,N_674);
or U1395 (N_1395,In_252,In_1276);
or U1396 (N_1396,In_45,N_598);
xnor U1397 (N_1397,N_853,In_497);
and U1398 (N_1398,N_710,N_483);
nor U1399 (N_1399,N_711,In_1448);
xor U1400 (N_1400,In_28,In_1723);
or U1401 (N_1401,In_712,In_1015);
xnor U1402 (N_1402,N_625,N_787);
nor U1403 (N_1403,N_287,N_969);
and U1404 (N_1404,N_837,In_2152);
nor U1405 (N_1405,N_636,N_998);
and U1406 (N_1406,N_550,N_167);
nor U1407 (N_1407,In_1950,N_582);
or U1408 (N_1408,In_1867,In_1415);
nor U1409 (N_1409,N_977,In_1636);
or U1410 (N_1410,N_597,In_112);
nor U1411 (N_1411,In_762,In_1628);
nand U1412 (N_1412,In_352,In_458);
nor U1413 (N_1413,N_934,N_946);
and U1414 (N_1414,N_304,In_1406);
nand U1415 (N_1415,In_2148,In_937);
nor U1416 (N_1416,In_560,N_553);
xnor U1417 (N_1417,N_993,N_749);
nand U1418 (N_1418,N_959,N_708);
nand U1419 (N_1419,In_23,N_604);
or U1420 (N_1420,In_1198,In_2308);
or U1421 (N_1421,In_134,In_660);
nand U1422 (N_1422,N_296,N_17);
nand U1423 (N_1423,N_609,In_608);
xnor U1424 (N_1424,N_693,N_337);
nand U1425 (N_1425,N_358,N_895);
nor U1426 (N_1426,N_772,In_1709);
xor U1427 (N_1427,In_1484,In_1995);
and U1428 (N_1428,In_1144,In_907);
or U1429 (N_1429,In_1265,N_923);
and U1430 (N_1430,In_2322,N_56);
and U1431 (N_1431,In_2469,In_1684);
nand U1432 (N_1432,N_469,N_738);
nor U1433 (N_1433,N_230,In_862);
or U1434 (N_1434,N_548,In_1159);
xnor U1435 (N_1435,N_627,In_1102);
and U1436 (N_1436,In_2195,In_131);
nor U1437 (N_1437,N_242,In_645);
nand U1438 (N_1438,N_733,N_589);
xor U1439 (N_1439,In_1441,N_438);
or U1440 (N_1440,In_164,N_864);
and U1441 (N_1441,In_1984,In_1316);
nor U1442 (N_1442,N_98,In_2408);
xor U1443 (N_1443,In_1659,In_2255);
nor U1444 (N_1444,N_869,N_939);
nor U1445 (N_1445,In_977,N_603);
nor U1446 (N_1446,N_315,N_614);
nor U1447 (N_1447,N_768,N_865);
nor U1448 (N_1448,In_822,N_117);
and U1449 (N_1449,N_55,In_890);
or U1450 (N_1450,In_377,In_412);
nor U1451 (N_1451,In_917,N_882);
xor U1452 (N_1452,In_1194,In_190);
and U1453 (N_1453,N_705,In_444);
and U1454 (N_1454,N_682,In_465);
or U1455 (N_1455,N_501,N_432);
or U1456 (N_1456,N_539,N_978);
nand U1457 (N_1457,In_1669,N_701);
or U1458 (N_1458,In_525,In_2108);
nand U1459 (N_1459,N_184,N_579);
and U1460 (N_1460,In_1106,N_204);
xnor U1461 (N_1461,In_1146,In_1394);
xnor U1462 (N_1462,N_20,N_623);
and U1463 (N_1463,In_1162,In_2068);
and U1464 (N_1464,In_95,In_1403);
or U1465 (N_1465,N_781,N_6);
or U1466 (N_1466,In_898,N_964);
and U1467 (N_1467,In_1172,In_2326);
nor U1468 (N_1468,In_1949,N_294);
and U1469 (N_1469,In_1398,N_52);
nand U1470 (N_1470,N_694,In_126);
or U1471 (N_1471,In_2260,In_1407);
or U1472 (N_1472,In_2240,N_863);
xnor U1473 (N_1473,N_822,In_1245);
xnor U1474 (N_1474,In_1753,N_706);
nand U1475 (N_1475,N_605,In_992);
nand U1476 (N_1476,In_1493,N_593);
or U1477 (N_1477,N_660,In_2089);
xor U1478 (N_1478,N_937,N_624);
or U1479 (N_1479,In_2259,In_348);
and U1480 (N_1480,In_849,In_1527);
xnor U1481 (N_1481,N_936,In_795);
nor U1482 (N_1482,N_610,In_1475);
nor U1483 (N_1483,In_1095,N_580);
xor U1484 (N_1484,In_1789,In_864);
nand U1485 (N_1485,In_2102,In_589);
and U1486 (N_1486,In_2233,In_380);
and U1487 (N_1487,In_1379,N_49);
or U1488 (N_1488,In_66,N_824);
nand U1489 (N_1489,In_177,N_907);
and U1490 (N_1490,In_2237,In_1592);
xnor U1491 (N_1491,N_266,In_1004);
xor U1492 (N_1492,N_791,In_2080);
and U1493 (N_1493,In_1626,N_367);
or U1494 (N_1494,N_902,N_909);
nand U1495 (N_1495,N_530,In_678);
nor U1496 (N_1496,In_2274,N_119);
xor U1497 (N_1497,N_646,N_220);
and U1498 (N_1498,N_545,In_2);
and U1499 (N_1499,N_378,In_2057);
xor U1500 (N_1500,N_1030,N_699);
and U1501 (N_1501,In_1898,N_1060);
and U1502 (N_1502,N_1435,N_1065);
or U1503 (N_1503,N_1485,N_1450);
xor U1504 (N_1504,N_1044,In_1003);
xnor U1505 (N_1505,In_173,In_2144);
and U1506 (N_1506,N_1163,In_446);
xnor U1507 (N_1507,N_654,N_1169);
nor U1508 (N_1508,N_1199,N_1071);
nand U1509 (N_1509,N_456,In_430);
nand U1510 (N_1510,In_1426,N_898);
and U1511 (N_1511,N_1005,In_939);
nand U1512 (N_1512,N_1360,In_507);
xnor U1513 (N_1513,N_1113,In_1844);
and U1514 (N_1514,In_2427,N_1309);
nand U1515 (N_1515,N_1325,In_1802);
nor U1516 (N_1516,In_607,N_1253);
and U1517 (N_1517,N_1330,In_1579);
nand U1518 (N_1518,N_528,In_1380);
nand U1519 (N_1519,N_602,N_1241);
xor U1520 (N_1520,N_1348,In_699);
nor U1521 (N_1521,N_1024,N_789);
or U1522 (N_1522,In_1078,In_1278);
nand U1523 (N_1523,N_1138,N_730);
nand U1524 (N_1524,N_1463,N_1088);
or U1525 (N_1525,N_77,N_1181);
and U1526 (N_1526,N_618,N_997);
or U1527 (N_1527,N_1135,N_411);
nand U1528 (N_1528,N_1101,N_1176);
nand U1529 (N_1529,In_1046,In_968);
nor U1530 (N_1530,N_1331,N_74);
nand U1531 (N_1531,N_1258,N_1074);
nor U1532 (N_1532,N_209,In_739);
and U1533 (N_1533,N_945,In_2478);
and U1534 (N_1534,N_1032,In_2005);
nand U1535 (N_1535,N_1341,N_1404);
xnor U1536 (N_1536,N_1197,N_196);
nor U1537 (N_1537,N_1312,N_1214);
and U1538 (N_1538,In_792,In_127);
and U1539 (N_1539,N_1180,N_594);
xor U1540 (N_1540,N_1458,In_597);
or U1541 (N_1541,In_547,N_1232);
and U1542 (N_1542,N_818,N_1277);
and U1543 (N_1543,N_656,N_1112);
xor U1544 (N_1544,N_510,N_529);
and U1545 (N_1545,N_1382,N_1063);
or U1546 (N_1546,N_155,N_1082);
nor U1547 (N_1547,N_1087,In_1429);
and U1548 (N_1548,N_1185,N_1303);
or U1549 (N_1549,In_947,N_1263);
or U1550 (N_1550,N_595,In_38);
or U1551 (N_1551,N_862,N_1286);
and U1552 (N_1552,N_871,In_1711);
xnor U1553 (N_1553,In_1287,N_1014);
or U1554 (N_1554,N_1216,N_1218);
nand U1555 (N_1555,In_332,N_1379);
nor U1556 (N_1556,N_1217,N_1480);
nand U1557 (N_1557,N_1049,In_479);
xor U1558 (N_1558,N_794,In_1672);
nand U1559 (N_1559,In_2076,N_704);
xnor U1560 (N_1560,N_1172,In_327);
or U1561 (N_1561,In_2004,N_673);
nor U1562 (N_1562,N_1431,In_1967);
and U1563 (N_1563,N_1254,N_1410);
nor U1564 (N_1564,N_1007,In_1770);
nor U1565 (N_1565,N_1339,N_803);
xnor U1566 (N_1566,N_1323,N_1124);
and U1567 (N_1567,N_1171,N_799);
nor U1568 (N_1568,N_756,N_846);
xor U1569 (N_1569,N_1021,N_1461);
nand U1570 (N_1570,In_1487,N_1354);
and U1571 (N_1571,N_415,N_1015);
nand U1572 (N_1572,N_215,In_1321);
nor U1573 (N_1573,N_1186,N_146);
nor U1574 (N_1574,N_698,N_1483);
nor U1575 (N_1575,N_1342,N_410);
nand U1576 (N_1576,In_393,N_1002);
nor U1577 (N_1577,In_662,In_335);
and U1578 (N_1578,In_1108,N_281);
nand U1579 (N_1579,In_281,N_1152);
nor U1580 (N_1580,N_925,In_1214);
nand U1581 (N_1581,N_401,In_2497);
nor U1582 (N_1582,N_1078,In_425);
and U1583 (N_1583,N_1419,N_1384);
nand U1584 (N_1584,In_1653,N_1104);
and U1585 (N_1585,In_12,N_1210);
nor U1586 (N_1586,In_2015,N_24);
and U1587 (N_1587,N_670,N_669);
and U1588 (N_1588,N_344,In_399);
nand U1589 (N_1589,N_1196,N_1280);
and U1590 (N_1590,N_1444,N_1434);
and U1591 (N_1591,N_333,In_1664);
or U1592 (N_1592,In_1202,N_567);
or U1593 (N_1593,In_1901,N_727);
xor U1594 (N_1594,In_1951,In_1583);
xor U1595 (N_1595,In_846,In_27);
nand U1596 (N_1596,N_265,In_664);
nand U1597 (N_1597,N_888,N_1205);
or U1598 (N_1598,N_1261,N_1440);
or U1599 (N_1599,N_1122,N_1156);
nand U1600 (N_1600,N_1316,N_1110);
and U1601 (N_1601,N_1433,In_89);
xnor U1602 (N_1602,In_2330,N_1275);
or U1603 (N_1603,N_1357,N_1383);
nand U1604 (N_1604,N_1359,N_820);
nor U1605 (N_1605,N_1420,N_905);
nand U1606 (N_1606,In_306,In_863);
or U1607 (N_1607,N_633,N_1034);
or U1608 (N_1608,N_1498,N_1321);
nand U1609 (N_1609,N_1374,In_1486);
nor U1610 (N_1610,In_1344,In_1240);
nand U1611 (N_1611,N_1157,N_813);
xor U1612 (N_1612,N_1429,In_268);
or U1613 (N_1613,In_5,N_158);
nor U1614 (N_1614,N_1243,N_1084);
nand U1615 (N_1615,N_1430,N_1066);
or U1616 (N_1616,In_528,N_1120);
and U1617 (N_1617,N_1329,N_1234);
or U1618 (N_1618,In_617,In_2039);
nand U1619 (N_1619,N_972,N_1402);
nor U1620 (N_1620,N_1067,N_513);
nor U1621 (N_1621,N_981,N_1438);
xnor U1622 (N_1622,In_2107,N_1028);
and U1623 (N_1623,N_1479,N_1064);
or U1624 (N_1624,N_1153,N_1260);
nand U1625 (N_1625,N_439,N_1370);
or U1626 (N_1626,N_1418,N_891);
and U1627 (N_1627,N_679,N_899);
and U1628 (N_1628,N_983,In_1630);
xnor U1629 (N_1629,N_1222,N_1136);
nor U1630 (N_1630,N_688,In_1339);
and U1631 (N_1631,In_2470,In_1336);
nand U1632 (N_1632,N_1226,N_1307);
nor U1633 (N_1633,N_1406,N_941);
xnor U1634 (N_1634,N_1454,N_1393);
xor U1635 (N_1635,N_1011,N_1022);
xor U1636 (N_1636,N_1193,N_1095);
xnor U1637 (N_1637,N_283,N_622);
nand U1638 (N_1638,N_1413,In_1545);
xor U1639 (N_1639,N_1000,In_1191);
xnor U1640 (N_1640,N_1472,N_1236);
nor U1641 (N_1641,N_1211,In_994);
or U1642 (N_1642,N_1392,N_1389);
nand U1643 (N_1643,N_1373,N_930);
xnor U1644 (N_1644,N_691,N_1492);
or U1645 (N_1645,N_87,N_1225);
nor U1646 (N_1646,In_1859,N_164);
xor U1647 (N_1647,In_1884,N_1107);
or U1648 (N_1648,N_1130,N_1097);
or U1649 (N_1649,N_887,In_819);
nand U1650 (N_1650,N_742,N_645);
and U1651 (N_1651,N_1310,N_16);
or U1652 (N_1652,N_1167,N_1414);
or U1653 (N_1653,N_1381,N_1499);
xor U1654 (N_1654,N_1358,N_239);
xnor U1655 (N_1655,N_933,N_592);
and U1656 (N_1656,N_881,N_583);
xnor U1657 (N_1657,N_1183,N_872);
nor U1658 (N_1658,N_1350,N_840);
or U1659 (N_1659,N_104,N_1302);
nor U1660 (N_1660,N_1338,N_416);
nand U1661 (N_1661,In_1602,N_1108);
nor U1662 (N_1662,N_1315,N_1308);
nor U1663 (N_1663,N_1109,N_1201);
and U1664 (N_1664,In_1832,N_661);
nand U1665 (N_1665,N_875,N_1224);
and U1666 (N_1666,In_1021,In_107);
nor U1667 (N_1667,In_1939,In_1540);
and U1668 (N_1668,N_1409,N_1029);
nand U1669 (N_1669,N_1327,N_1056);
xor U1670 (N_1670,N_1213,N_1367);
and U1671 (N_1671,N_1127,N_1070);
nor U1672 (N_1672,N_1343,N_1407);
or U1673 (N_1673,N_1026,N_1004);
or U1674 (N_1674,N_957,In_508);
xor U1675 (N_1675,N_1421,N_1347);
and U1676 (N_1676,N_1198,N_1209);
xnor U1677 (N_1677,N_1207,N_1313);
or U1678 (N_1678,N_963,N_1491);
nand U1679 (N_1679,N_1265,N_1257);
xnor U1680 (N_1680,N_1246,N_454);
nand U1681 (N_1681,N_346,N_1481);
nand U1682 (N_1682,N_1062,In_2490);
nor U1683 (N_1683,In_1416,N_1072);
or U1684 (N_1684,N_1053,N_50);
or U1685 (N_1685,In_477,In_364);
and U1686 (N_1686,In_26,N_1179);
or U1687 (N_1687,N_1158,N_1497);
nand U1688 (N_1688,N_93,N_1304);
and U1689 (N_1689,N_1055,In_63);
and U1690 (N_1690,N_537,N_1114);
or U1691 (N_1691,In_1354,N_900);
or U1692 (N_1692,In_704,N_1284);
nor U1693 (N_1693,N_1092,N_1090);
nand U1694 (N_1694,N_935,N_686);
and U1695 (N_1695,In_2273,In_1971);
xor U1696 (N_1696,N_1194,In_1564);
nand U1697 (N_1697,N_1182,N_1105);
nor U1698 (N_1698,N_1189,N_1267);
nor U1699 (N_1699,In_995,In_417);
and U1700 (N_1700,N_1317,N_1351);
xor U1701 (N_1701,N_1047,N_1437);
nand U1702 (N_1702,N_1477,N_549);
xor U1703 (N_1703,In_135,In_87);
nand U1704 (N_1704,In_1923,N_677);
nor U1705 (N_1705,In_549,N_1045);
xor U1706 (N_1706,N_1355,In_420);
and U1707 (N_1707,N_1314,N_210);
nor U1708 (N_1708,In_1565,N_1239);
and U1709 (N_1709,N_1018,In_789);
xor U1710 (N_1710,N_709,N_1178);
or U1711 (N_1711,N_785,N_1161);
nor U1712 (N_1712,N_1459,N_1126);
nand U1713 (N_1713,In_2186,N_719);
nor U1714 (N_1714,In_991,In_788);
nor U1715 (N_1715,In_502,N_1285);
xor U1716 (N_1716,In_1721,In_2065);
xnor U1717 (N_1717,N_1424,N_1340);
nor U1718 (N_1718,N_308,N_1428);
nand U1719 (N_1719,N_1009,N_1488);
xor U1720 (N_1720,In_391,N_1013);
and U1721 (N_1721,N_1174,N_1150);
or U1722 (N_1722,N_1098,N_542);
and U1723 (N_1723,N_1474,N_1050);
nand U1724 (N_1724,N_1443,N_1371);
and U1725 (N_1725,In_1139,N_1439);
and U1726 (N_1726,N_1332,In_13);
or U1727 (N_1727,N_1447,N_1137);
xnor U1728 (N_1728,N_565,N_1290);
nor U1729 (N_1729,N_1442,N_518);
and U1730 (N_1730,In_1550,N_802);
or U1731 (N_1731,N_1111,N_1173);
and U1732 (N_1732,N_884,In_1337);
xnor U1733 (N_1733,N_1334,In_457);
nand U1734 (N_1734,In_496,N_252);
or U1735 (N_1735,N_1322,In_361);
nor U1736 (N_1736,N_1306,N_966);
and U1737 (N_1737,In_2467,N_1394);
and U1738 (N_1738,In_2189,N_238);
xnor U1739 (N_1739,N_1349,N_350);
nand U1740 (N_1740,N_1276,N_1368);
and U1741 (N_1741,N_980,N_1403);
xor U1742 (N_1742,In_1081,N_1289);
nand U1743 (N_1743,In_1888,N_1395);
xor U1744 (N_1744,N_1490,In_2234);
or U1745 (N_1745,In_1285,N_648);
xor U1746 (N_1746,N_1311,In_1586);
xor U1747 (N_1747,In_568,N_1445);
nand U1748 (N_1748,N_535,N_1282);
nor U1749 (N_1749,N_1085,In_429);
or U1750 (N_1750,N_655,N_1148);
and U1751 (N_1751,In_622,In_2190);
xnor U1752 (N_1752,N_1143,N_1377);
nor U1753 (N_1753,N_61,In_1149);
or U1754 (N_1754,In_62,N_1346);
or U1755 (N_1755,N_1455,N_1345);
nand U1756 (N_1756,N_1184,N_387);
and U1757 (N_1757,N_856,N_1432);
and U1758 (N_1758,N_1077,N_1252);
or U1759 (N_1759,In_1503,N_1344);
or U1760 (N_1760,N_1417,In_1451);
xor U1761 (N_1761,N_1027,In_2159);
and U1762 (N_1762,In_2022,N_1361);
nand U1763 (N_1763,N_1235,N_1423);
xnor U1764 (N_1764,N_1190,N_1133);
xor U1765 (N_1765,N_1221,N_1249);
nor U1766 (N_1766,In_2157,N_1369);
or U1767 (N_1767,In_156,In_2475);
nor U1768 (N_1768,N_1248,N_1228);
xnor U1769 (N_1769,N_1141,N_1264);
nand U1770 (N_1770,In_2465,N_221);
and U1771 (N_1771,In_1188,N_1251);
or U1772 (N_1772,N_1175,N_774);
nor U1773 (N_1773,N_950,N_1042);
nand U1774 (N_1774,N_1380,N_1229);
nand U1775 (N_1775,N_363,N_760);
xor U1776 (N_1776,N_1244,N_128);
nand U1777 (N_1777,N_1259,N_1294);
and U1778 (N_1778,In_185,In_2217);
nor U1779 (N_1779,N_653,In_1696);
xnor U1780 (N_1780,In_1059,In_2139);
nand U1781 (N_1781,N_1320,N_766);
or U1782 (N_1782,N_1240,In_1834);
nand U1783 (N_1783,In_714,In_249);
xnor U1784 (N_1784,In_196,N_1462);
nand U1785 (N_1785,N_897,N_970);
nor U1786 (N_1786,In_1417,In_1255);
or U1787 (N_1787,N_1295,N_564);
nor U1788 (N_1788,N_1352,In_1158);
and U1789 (N_1789,N_716,N_1486);
and U1790 (N_1790,N_690,In_1482);
xor U1791 (N_1791,N_1118,N_407);
nand U1792 (N_1792,N_1415,N_1336);
nor U1793 (N_1793,N_1025,N_665);
xor U1794 (N_1794,N_1388,N_1164);
nor U1795 (N_1795,In_2023,N_1273);
and U1796 (N_1796,In_280,N_1456);
xnor U1797 (N_1797,In_2376,In_0);
and U1798 (N_1798,N_1200,N_1017);
nand U1799 (N_1799,N_280,In_180);
nor U1800 (N_1800,In_644,N_795);
nor U1801 (N_1801,N_1215,N_1103);
and U1802 (N_1802,In_1100,In_2268);
and U1803 (N_1803,N_1262,In_330);
and U1804 (N_1804,N_1300,N_1129);
nor U1805 (N_1805,N_1227,N_1247);
nor U1806 (N_1806,N_1408,N_1054);
nand U1807 (N_1807,N_1100,N_798);
nor U1808 (N_1808,N_1250,In_1099);
xnor U1809 (N_1809,In_1084,N_13);
nand U1810 (N_1810,In_2244,N_762);
nand U1811 (N_1811,N_1069,N_1468);
nor U1812 (N_1812,In_807,N_1121);
nand U1813 (N_1813,N_1489,N_562);
nor U1814 (N_1814,N_991,N_782);
nand U1815 (N_1815,N_1333,N_493);
and U1816 (N_1816,In_1392,N_889);
or U1817 (N_1817,N_1279,In_1385);
nand U1818 (N_1818,N_568,In_2346);
xnor U1819 (N_1819,N_1038,In_1868);
xor U1820 (N_1820,N_1144,N_1230);
and U1821 (N_1821,N_1061,N_651);
xor U1822 (N_1822,In_1061,N_1083);
nand U1823 (N_1823,N_376,N_1008);
and U1824 (N_1824,In_1327,N_1192);
nor U1825 (N_1825,In_642,In_1988);
xnor U1826 (N_1826,N_370,In_67);
xor U1827 (N_1827,In_1067,N_507);
nor U1828 (N_1828,N_1039,In_510);
nand U1829 (N_1829,N_1166,N_784);
and U1830 (N_1830,N_1390,N_878);
or U1831 (N_1831,In_1983,N_1188);
xor U1832 (N_1832,N_511,N_1272);
nand U1833 (N_1833,N_318,N_1154);
xor U1834 (N_1834,N_1099,N_400);
xnor U1835 (N_1835,N_728,N_1231);
xnor U1836 (N_1836,N_1016,N_388);
and U1837 (N_1837,N_763,In_2309);
and U1838 (N_1838,In_908,In_988);
and U1839 (N_1839,N_1452,N_1233);
and U1840 (N_1840,In_68,N_1125);
nor U1841 (N_1841,In_183,N_1494);
nand U1842 (N_1842,In_652,N_753);
nand U1843 (N_1843,N_1068,N_1238);
nor U1844 (N_1844,N_689,N_948);
nor U1845 (N_1845,N_657,N_1116);
xnor U1846 (N_1846,N_1487,N_621);
nand U1847 (N_1847,N_1387,N_1145);
and U1848 (N_1848,N_1140,N_1426);
nand U1849 (N_1849,N_1318,N_1048);
nand U1850 (N_1850,N_1326,In_2160);
nor U1851 (N_1851,N_1391,N_1187);
and U1852 (N_1852,In_323,N_1019);
or U1853 (N_1853,N_718,N_504);
nor U1854 (N_1854,In_1974,N_1162);
or U1855 (N_1855,N_1353,N_1268);
nor U1856 (N_1856,N_365,N_44);
or U1857 (N_1857,In_1509,N_1335);
and U1858 (N_1858,In_1322,In_904);
and U1859 (N_1859,In_1274,N_1448);
nand U1860 (N_1860,N_917,N_1212);
xor U1861 (N_1861,N_617,N_968);
xnor U1862 (N_1862,N_1305,N_1288);
nor U1863 (N_1863,N_1457,N_1328);
xnor U1864 (N_1864,N_1495,In_1758);
or U1865 (N_1865,N_1132,In_1335);
or U1866 (N_1866,In_308,N_1469);
or U1867 (N_1867,N_697,N_1470);
nor U1868 (N_1868,In_599,N_512);
nand U1869 (N_1869,N_767,N_1237);
and U1870 (N_1870,N_725,In_1953);
xor U1871 (N_1871,N_821,In_1875);
nand U1872 (N_1872,N_1473,N_1397);
and U1873 (N_1873,N_1075,N_1170);
xor U1874 (N_1874,N_440,N_1296);
nand U1875 (N_1875,In_76,In_328);
or U1876 (N_1876,In_1414,In_1388);
or U1877 (N_1877,N_1475,N_720);
nand U1878 (N_1878,N_1453,N_1031);
xor U1879 (N_1879,N_1293,N_1139);
and U1880 (N_1880,N_982,N_1208);
nor U1881 (N_1881,N_1465,N_1464);
nand U1882 (N_1882,N_552,In_2088);
xor U1883 (N_1883,In_1781,N_1058);
xnor U1884 (N_1884,In_2247,In_834);
nor U1885 (N_1885,N_988,In_73);
nor U1886 (N_1886,N_1177,N_447);
xnor U1887 (N_1887,In_1007,N_1165);
xor U1888 (N_1888,N_1147,N_1467);
xor U1889 (N_1889,N_916,N_1399);
xnor U1890 (N_1890,N_1128,In_1688);
nor U1891 (N_1891,N_1482,In_81);
or U1892 (N_1892,N_667,N_1396);
nor U1893 (N_1893,N_814,In_2103);
and U1894 (N_1894,In_1476,N_1274);
xnor U1895 (N_1895,N_1160,N_1037);
nor U1896 (N_1896,N_1385,In_1091);
or U1897 (N_1897,N_1269,In_2028);
xnor U1898 (N_1898,In_1402,N_1219);
nand U1899 (N_1899,N_962,N_1297);
nand U1900 (N_1900,In_1879,N_783);
nand U1901 (N_1901,N_928,N_1422);
or U1902 (N_1902,In_436,In_2173);
or U1903 (N_1903,N_1427,N_1043);
nand U1904 (N_1904,N_1012,N_1001);
nor U1905 (N_1905,N_1299,N_1446);
xor U1906 (N_1906,N_1094,In_2399);
nand U1907 (N_1907,N_36,N_1102);
nor U1908 (N_1908,N_1040,N_838);
nand U1909 (N_1909,N_516,N_1278);
nor U1910 (N_1910,In_1973,N_1202);
nor U1911 (N_1911,N_1146,N_1478);
or U1912 (N_1912,N_1006,N_1496);
nand U1913 (N_1913,N_1291,N_208);
nor U1914 (N_1914,N_1096,N_1059);
nand U1915 (N_1915,In_780,In_1969);
and U1916 (N_1916,N_460,N_161);
and U1917 (N_1917,N_1301,In_314);
xor U1918 (N_1918,N_1271,N_868);
and U1919 (N_1919,N_652,In_2151);
nor U1920 (N_1920,In_276,N_1020);
or U1921 (N_1921,In_143,N_1471);
xnor U1922 (N_1922,In_1554,In_2137);
xnor U1923 (N_1923,N_1041,N_1081);
nor U1924 (N_1924,N_1073,N_1412);
nand U1925 (N_1925,N_859,N_1398);
and U1926 (N_1926,N_1204,N_1436);
xor U1927 (N_1927,N_1386,N_1356);
or U1928 (N_1928,N_788,In_2298);
or U1929 (N_1929,In_454,N_1142);
xor U1930 (N_1930,N_1149,In_166);
or U1931 (N_1931,N_1057,N_1378);
nor U1932 (N_1932,N_1255,N_1245);
nand U1933 (N_1933,N_683,In_969);
and U1934 (N_1934,In_1562,In_1544);
or U1935 (N_1935,In_1595,N_790);
nand U1936 (N_1936,In_1862,N_1363);
nor U1937 (N_1937,N_1093,N_1401);
xnor U1938 (N_1938,In_2388,In_1324);
nor U1939 (N_1939,N_994,N_976);
nand U1940 (N_1940,In_1093,N_1405);
and U1941 (N_1941,N_478,In_424);
nor U1942 (N_1942,N_845,N_1151);
nand U1943 (N_1943,N_804,N_1287);
or U1944 (N_1944,N_1441,N_1451);
xnor U1945 (N_1945,N_634,N_1298);
or U1946 (N_1946,In_1861,N_1376);
and U1947 (N_1947,N_1283,In_1805);
or U1948 (N_1948,N_1484,N_671);
nand U1949 (N_1949,In_2118,N_1365);
nand U1950 (N_1950,In_2471,In_58);
or U1951 (N_1951,N_1256,N_1191);
nor U1952 (N_1952,N_186,N_1091);
or U1953 (N_1953,N_827,N_639);
and U1954 (N_1954,N_1337,N_1023);
nand U1955 (N_1955,N_577,N_1466);
and U1956 (N_1956,In_842,N_723);
xor U1957 (N_1957,N_815,N_1076);
or U1958 (N_1958,N_231,N_637);
nand U1959 (N_1959,In_286,N_757);
nand U1960 (N_1960,N_305,N_38);
and U1961 (N_1961,In_2177,N_278);
or U1962 (N_1962,N_1119,In_656);
nand U1963 (N_1963,N_918,N_1416);
nand U1964 (N_1964,N_1372,N_893);
nor U1965 (N_1965,N_1046,N_1266);
or U1966 (N_1966,N_1400,N_658);
and U1967 (N_1967,N_1159,N_1123);
and U1968 (N_1968,In_1976,N_1035);
and U1969 (N_1969,N_1131,N_1080);
nand U1970 (N_1970,N_1362,N_1319);
and U1971 (N_1971,N_1292,N_1086);
or U1972 (N_1972,N_1155,N_1223);
and U1973 (N_1973,In_1114,N_259);
nand U1974 (N_1974,N_245,N_1033);
nor U1975 (N_1975,N_1364,N_922);
nor U1976 (N_1976,N_1089,N_886);
nor U1977 (N_1977,N_967,N_1220);
or U1978 (N_1978,N_1493,N_1195);
xor U1979 (N_1979,In_752,N_809);
xor U1980 (N_1980,In_1341,N_640);
or U1981 (N_1981,N_1411,N_1449);
or U1982 (N_1982,N_1003,N_1168);
nand U1983 (N_1983,N_140,In_246);
nor U1984 (N_1984,N_1010,In_1541);
nand U1985 (N_1985,N_554,N_214);
and U1986 (N_1986,N_109,N_1203);
xnor U1987 (N_1987,In_372,N_1242);
xor U1988 (N_1988,N_1375,N_1117);
nand U1989 (N_1989,N_1460,N_139);
and U1990 (N_1990,N_1134,N_1051);
xor U1991 (N_1991,N_1036,N_1270);
xnor U1992 (N_1992,N_1281,N_1206);
xor U1993 (N_1993,N_745,In_866);
or U1994 (N_1994,N_1324,N_1425);
or U1995 (N_1995,In_2371,N_1366);
xor U1996 (N_1996,N_1079,N_1052);
nor U1997 (N_1997,In_2364,N_1476);
nand U1998 (N_1998,N_1106,N_1115);
nand U1999 (N_1999,In_277,In_1205);
nand U2000 (N_2000,N_1656,N_1771);
xnor U2001 (N_2001,N_1929,N_1748);
nand U2002 (N_2002,N_1857,N_1514);
xor U2003 (N_2003,N_1724,N_1553);
and U2004 (N_2004,N_1997,N_1625);
and U2005 (N_2005,N_1945,N_1687);
nor U2006 (N_2006,N_1801,N_1933);
and U2007 (N_2007,N_1552,N_1793);
xnor U2008 (N_2008,N_1965,N_1557);
nor U2009 (N_2009,N_1858,N_1927);
nor U2010 (N_2010,N_1652,N_1838);
nor U2011 (N_2011,N_1706,N_1935);
or U2012 (N_2012,N_1718,N_1822);
or U2013 (N_2013,N_1735,N_1722);
nor U2014 (N_2014,N_1993,N_1797);
nor U2015 (N_2015,N_1977,N_1563);
nand U2016 (N_2016,N_1620,N_1518);
nor U2017 (N_2017,N_1526,N_1593);
or U2018 (N_2018,N_1504,N_1786);
and U2019 (N_2019,N_1930,N_1781);
xnor U2020 (N_2020,N_1598,N_1931);
and U2021 (N_2021,N_1626,N_1728);
or U2022 (N_2022,N_1795,N_1764);
nor U2023 (N_2023,N_1996,N_1916);
nor U2024 (N_2024,N_1988,N_1824);
nand U2025 (N_2025,N_1532,N_1684);
nor U2026 (N_2026,N_1805,N_1804);
xor U2027 (N_2027,N_1877,N_1716);
nand U2028 (N_2028,N_1729,N_1865);
nor U2029 (N_2029,N_1769,N_1899);
nand U2030 (N_2030,N_1530,N_1507);
or U2031 (N_2031,N_1703,N_1522);
and U2032 (N_2032,N_1803,N_1683);
and U2033 (N_2033,N_1566,N_1660);
xnor U2034 (N_2034,N_1647,N_1616);
xor U2035 (N_2035,N_1742,N_1898);
and U2036 (N_2036,N_1952,N_1770);
nor U2037 (N_2037,N_1905,N_1713);
nand U2038 (N_2038,N_1638,N_1776);
and U2039 (N_2039,N_1853,N_1813);
nor U2040 (N_2040,N_1697,N_1689);
nand U2041 (N_2041,N_1998,N_1873);
and U2042 (N_2042,N_1926,N_1704);
xnor U2043 (N_2043,N_1631,N_1774);
xnor U2044 (N_2044,N_1653,N_1709);
nor U2045 (N_2045,N_1794,N_1628);
or U2046 (N_2046,N_1634,N_1723);
nand U2047 (N_2047,N_1893,N_1740);
and U2048 (N_2048,N_1675,N_1880);
or U2049 (N_2049,N_1747,N_1731);
or U2050 (N_2050,N_1839,N_1758);
or U2051 (N_2051,N_1963,N_1934);
xnor U2052 (N_2052,N_1546,N_1627);
and U2053 (N_2053,N_1921,N_1955);
or U2054 (N_2054,N_1734,N_1649);
nor U2055 (N_2055,N_1529,N_1904);
or U2056 (N_2056,N_1698,N_1944);
or U2057 (N_2057,N_1919,N_1861);
and U2058 (N_2058,N_1701,N_1501);
or U2059 (N_2059,N_1784,N_1862);
and U2060 (N_2060,N_1702,N_1991);
or U2061 (N_2061,N_1937,N_1920);
nor U2062 (N_2062,N_1544,N_1572);
or U2063 (N_2063,N_1835,N_1915);
and U2064 (N_2064,N_1727,N_1881);
nand U2065 (N_2065,N_1644,N_1842);
or U2066 (N_2066,N_1502,N_1527);
xor U2067 (N_2067,N_1612,N_1579);
and U2068 (N_2068,N_1691,N_1978);
nand U2069 (N_2069,N_1782,N_1562);
or U2070 (N_2070,N_1609,N_1906);
and U2071 (N_2071,N_1954,N_1889);
nand U2072 (N_2072,N_1597,N_1744);
and U2073 (N_2073,N_1619,N_1985);
and U2074 (N_2074,N_1995,N_1536);
nor U2075 (N_2075,N_1632,N_1533);
nor U2076 (N_2076,N_1864,N_1743);
and U2077 (N_2077,N_1914,N_1615);
nor U2078 (N_2078,N_1556,N_1674);
xnor U2079 (N_2079,N_1953,N_1767);
xnor U2080 (N_2080,N_1922,N_1558);
nand U2081 (N_2081,N_1633,N_1655);
xnor U2082 (N_2082,N_1506,N_1848);
xor U2083 (N_2083,N_1975,N_1534);
and U2084 (N_2084,N_1986,N_1610);
nand U2085 (N_2085,N_1690,N_1732);
xnor U2086 (N_2086,N_1549,N_1902);
nand U2087 (N_2087,N_1867,N_1568);
nor U2088 (N_2088,N_1772,N_1539);
or U2089 (N_2089,N_1989,N_1999);
xor U2090 (N_2090,N_1923,N_1680);
xor U2091 (N_2091,N_1886,N_1583);
and U2092 (N_2092,N_1694,N_1810);
xnor U2093 (N_2093,N_1524,N_1773);
and U2094 (N_2094,N_1950,N_1979);
nand U2095 (N_2095,N_1688,N_1719);
and U2096 (N_2096,N_1948,N_1753);
xnor U2097 (N_2097,N_1721,N_1587);
nand U2098 (N_2098,N_1621,N_1511);
and U2099 (N_2099,N_1841,N_1882);
or U2100 (N_2100,N_1624,N_1708);
nand U2101 (N_2101,N_1783,N_1541);
nor U2102 (N_2102,N_1775,N_1692);
nor U2103 (N_2103,N_1778,N_1676);
nand U2104 (N_2104,N_1637,N_1543);
or U2105 (N_2105,N_1959,N_1830);
nand U2106 (N_2106,N_1798,N_1576);
or U2107 (N_2107,N_1984,N_1595);
nand U2108 (N_2108,N_1685,N_1754);
nand U2109 (N_2109,N_1700,N_1720);
xor U2110 (N_2110,N_1663,N_1763);
nor U2111 (N_2111,N_1715,N_1942);
xor U2112 (N_2112,N_1828,N_1911);
nand U2113 (N_2113,N_1642,N_1917);
xnor U2114 (N_2114,N_1976,N_1800);
or U2115 (N_2115,N_1849,N_1851);
nand U2116 (N_2116,N_1589,N_1714);
nand U2117 (N_2117,N_1973,N_1519);
and U2118 (N_2118,N_1641,N_1622);
nand U2119 (N_2119,N_1662,N_1693);
xnor U2120 (N_2120,N_1829,N_1515);
nor U2121 (N_2121,N_1580,N_1791);
and U2122 (N_2122,N_1608,N_1760);
or U2123 (N_2123,N_1779,N_1629);
nand U2124 (N_2124,N_1717,N_1573);
xor U2125 (N_2125,N_1913,N_1560);
nand U2126 (N_2126,N_1554,N_1705);
xnor U2127 (N_2127,N_1575,N_1594);
and U2128 (N_2128,N_1650,N_1503);
xnor U2129 (N_2129,N_1538,N_1605);
and U2130 (N_2130,N_1651,N_1799);
nor U2131 (N_2131,N_1752,N_1667);
nand U2132 (N_2132,N_1516,N_1564);
nand U2133 (N_2133,N_1618,N_1903);
nor U2134 (N_2134,N_1585,N_1817);
or U2135 (N_2135,N_1845,N_1757);
or U2136 (N_2136,N_1961,N_1547);
xor U2137 (N_2137,N_1592,N_1808);
nor U2138 (N_2138,N_1910,N_1699);
and U2139 (N_2139,N_1550,N_1982);
and U2140 (N_2140,N_1821,N_1970);
nor U2141 (N_2141,N_1751,N_1578);
nor U2142 (N_2142,N_1679,N_1648);
xnor U2143 (N_2143,N_1925,N_1548);
nand U2144 (N_2144,N_1811,N_1844);
xnor U2145 (N_2145,N_1577,N_1630);
nand U2146 (N_2146,N_1831,N_1909);
nor U2147 (N_2147,N_1636,N_1846);
or U2148 (N_2148,N_1951,N_1834);
or U2149 (N_2149,N_1654,N_1745);
or U2150 (N_2150,N_1792,N_1664);
or U2151 (N_2151,N_1866,N_1940);
nand U2152 (N_2152,N_1561,N_1766);
nor U2153 (N_2153,N_1957,N_1535);
or U2154 (N_2154,N_1990,N_1900);
or U2155 (N_2155,N_1939,N_1707);
xor U2156 (N_2156,N_1513,N_1540);
nand U2157 (N_2157,N_1780,N_1785);
xor U2158 (N_2158,N_1787,N_1924);
nor U2159 (N_2159,N_1969,N_1678);
xor U2160 (N_2160,N_1892,N_1545);
nand U2161 (N_2161,N_1823,N_1671);
and U2162 (N_2162,N_1872,N_1581);
or U2163 (N_2163,N_1512,N_1659);
nand U2164 (N_2164,N_1843,N_1711);
xor U2165 (N_2165,N_1509,N_1938);
xnor U2166 (N_2166,N_1869,N_1980);
and U2167 (N_2167,N_1555,N_1790);
xor U2168 (N_2168,N_1582,N_1755);
nand U2169 (N_2169,N_1603,N_1946);
xor U2170 (N_2170,N_1640,N_1569);
or U2171 (N_2171,N_1908,N_1531);
nor U2172 (N_2172,N_1852,N_1665);
nand U2173 (N_2173,N_1847,N_1570);
nor U2174 (N_2174,N_1896,N_1796);
or U2175 (N_2175,N_1762,N_1885);
xnor U2176 (N_2176,N_1874,N_1816);
xnor U2177 (N_2177,N_1571,N_1876);
nor U2178 (N_2178,N_1672,N_1981);
nor U2179 (N_2179,N_1907,N_1584);
nand U2180 (N_2180,N_1863,N_1737);
nor U2181 (N_2181,N_1606,N_1574);
or U2182 (N_2182,N_1756,N_1870);
or U2183 (N_2183,N_1854,N_1875);
nor U2184 (N_2184,N_1623,N_1635);
or U2185 (N_2185,N_1657,N_1528);
xnor U2186 (N_2186,N_1588,N_1825);
nor U2187 (N_2187,N_1517,N_1918);
or U2188 (N_2188,N_1895,N_1551);
or U2189 (N_2189,N_1681,N_1613);
or U2190 (N_2190,N_1668,N_1897);
and U2191 (N_2191,N_1523,N_1814);
nor U2192 (N_2192,N_1712,N_1645);
or U2193 (N_2193,N_1599,N_1971);
or U2194 (N_2194,N_1890,N_1710);
or U2195 (N_2195,N_1639,N_1967);
or U2196 (N_2196,N_1947,N_1928);
nor U2197 (N_2197,N_1520,N_1525);
nand U2198 (N_2198,N_1658,N_1868);
and U2199 (N_2199,N_1666,N_1661);
and U2200 (N_2200,N_1827,N_1510);
nor U2201 (N_2201,N_1695,N_1567);
nand U2202 (N_2202,N_1833,N_1819);
nand U2203 (N_2203,N_1932,N_1974);
nor U2204 (N_2204,N_1730,N_1891);
nor U2205 (N_2205,N_1994,N_1850);
nor U2206 (N_2206,N_1643,N_1941);
and U2207 (N_2207,N_1809,N_1815);
nand U2208 (N_2208,N_1812,N_1859);
xnor U2209 (N_2209,N_1670,N_1860);
nand U2210 (N_2210,N_1542,N_1887);
nor U2211 (N_2211,N_1559,N_1818);
nand U2212 (N_2212,N_1733,N_1768);
nor U2213 (N_2213,N_1601,N_1600);
or U2214 (N_2214,N_1820,N_1836);
or U2215 (N_2215,N_1958,N_1565);
xor U2216 (N_2216,N_1840,N_1960);
nor U2217 (N_2217,N_1741,N_1992);
nand U2218 (N_2218,N_1725,N_1962);
and U2219 (N_2219,N_1646,N_1682);
and U2220 (N_2220,N_1607,N_1901);
or U2221 (N_2221,N_1604,N_1591);
nand U2222 (N_2222,N_1883,N_1739);
nor U2223 (N_2223,N_1802,N_1807);
nand U2224 (N_2224,N_1806,N_1855);
xnor U2225 (N_2225,N_1888,N_1602);
xor U2226 (N_2226,N_1964,N_1738);
nor U2227 (N_2227,N_1749,N_1894);
xor U2228 (N_2228,N_1856,N_1611);
and U2229 (N_2229,N_1590,N_1746);
xor U2230 (N_2230,N_1826,N_1726);
or U2231 (N_2231,N_1521,N_1505);
and U2232 (N_2232,N_1968,N_1789);
and U2233 (N_2233,N_1677,N_1884);
or U2234 (N_2234,N_1879,N_1614);
and U2235 (N_2235,N_1669,N_1837);
or U2236 (N_2236,N_1788,N_1759);
nand U2237 (N_2237,N_1750,N_1943);
nand U2238 (N_2238,N_1966,N_1537);
or U2239 (N_2239,N_1761,N_1832);
and U2240 (N_2240,N_1736,N_1586);
xnor U2241 (N_2241,N_1500,N_1673);
xnor U2242 (N_2242,N_1972,N_1617);
xor U2243 (N_2243,N_1878,N_1508);
xor U2244 (N_2244,N_1596,N_1987);
nor U2245 (N_2245,N_1686,N_1949);
nor U2246 (N_2246,N_1871,N_1912);
xor U2247 (N_2247,N_1983,N_1777);
xor U2248 (N_2248,N_1765,N_1956);
xnor U2249 (N_2249,N_1936,N_1696);
or U2250 (N_2250,N_1939,N_1833);
or U2251 (N_2251,N_1821,N_1625);
nand U2252 (N_2252,N_1651,N_1791);
nor U2253 (N_2253,N_1889,N_1788);
and U2254 (N_2254,N_1700,N_1615);
nor U2255 (N_2255,N_1875,N_1825);
and U2256 (N_2256,N_1661,N_1729);
nor U2257 (N_2257,N_1842,N_1840);
and U2258 (N_2258,N_1921,N_1739);
nand U2259 (N_2259,N_1977,N_1521);
and U2260 (N_2260,N_1719,N_1843);
and U2261 (N_2261,N_1610,N_1673);
xnor U2262 (N_2262,N_1543,N_1995);
nand U2263 (N_2263,N_1862,N_1658);
nand U2264 (N_2264,N_1633,N_1995);
or U2265 (N_2265,N_1991,N_1651);
and U2266 (N_2266,N_1966,N_1526);
nor U2267 (N_2267,N_1566,N_1541);
nand U2268 (N_2268,N_1779,N_1812);
or U2269 (N_2269,N_1826,N_1581);
nand U2270 (N_2270,N_1555,N_1994);
or U2271 (N_2271,N_1514,N_1667);
or U2272 (N_2272,N_1574,N_1592);
and U2273 (N_2273,N_1611,N_1885);
xor U2274 (N_2274,N_1931,N_1605);
xnor U2275 (N_2275,N_1892,N_1893);
nor U2276 (N_2276,N_1995,N_1864);
or U2277 (N_2277,N_1679,N_1632);
nand U2278 (N_2278,N_1736,N_1810);
nand U2279 (N_2279,N_1523,N_1661);
and U2280 (N_2280,N_1629,N_1933);
xnor U2281 (N_2281,N_1583,N_1578);
or U2282 (N_2282,N_1637,N_1987);
and U2283 (N_2283,N_1541,N_1512);
nand U2284 (N_2284,N_1560,N_1525);
nand U2285 (N_2285,N_1842,N_1670);
nand U2286 (N_2286,N_1945,N_1959);
xnor U2287 (N_2287,N_1965,N_1891);
nand U2288 (N_2288,N_1793,N_1595);
xnor U2289 (N_2289,N_1572,N_1835);
nand U2290 (N_2290,N_1757,N_1726);
nor U2291 (N_2291,N_1640,N_1529);
and U2292 (N_2292,N_1592,N_1800);
xnor U2293 (N_2293,N_1679,N_1985);
xnor U2294 (N_2294,N_1972,N_1566);
xor U2295 (N_2295,N_1527,N_1826);
xor U2296 (N_2296,N_1815,N_1539);
nand U2297 (N_2297,N_1504,N_1741);
nand U2298 (N_2298,N_1864,N_1886);
or U2299 (N_2299,N_1633,N_1963);
or U2300 (N_2300,N_1689,N_1847);
or U2301 (N_2301,N_1838,N_1504);
nor U2302 (N_2302,N_1769,N_1889);
or U2303 (N_2303,N_1900,N_1605);
xnor U2304 (N_2304,N_1945,N_1685);
nand U2305 (N_2305,N_1800,N_1756);
and U2306 (N_2306,N_1543,N_1754);
xnor U2307 (N_2307,N_1707,N_1896);
xnor U2308 (N_2308,N_1502,N_1635);
nor U2309 (N_2309,N_1835,N_1736);
and U2310 (N_2310,N_1623,N_1737);
and U2311 (N_2311,N_1520,N_1714);
or U2312 (N_2312,N_1751,N_1949);
xor U2313 (N_2313,N_1500,N_1605);
nor U2314 (N_2314,N_1779,N_1815);
and U2315 (N_2315,N_1521,N_1975);
and U2316 (N_2316,N_1768,N_1589);
xor U2317 (N_2317,N_1737,N_1835);
or U2318 (N_2318,N_1865,N_1685);
nand U2319 (N_2319,N_1810,N_1879);
nand U2320 (N_2320,N_1557,N_1753);
nand U2321 (N_2321,N_1951,N_1945);
nand U2322 (N_2322,N_1692,N_1660);
or U2323 (N_2323,N_1781,N_1858);
nor U2324 (N_2324,N_1591,N_1981);
xor U2325 (N_2325,N_1739,N_1686);
nor U2326 (N_2326,N_1678,N_1931);
nand U2327 (N_2327,N_1643,N_1959);
nand U2328 (N_2328,N_1594,N_1532);
nand U2329 (N_2329,N_1534,N_1937);
and U2330 (N_2330,N_1544,N_1807);
and U2331 (N_2331,N_1533,N_1924);
and U2332 (N_2332,N_1869,N_1713);
xor U2333 (N_2333,N_1880,N_1924);
xor U2334 (N_2334,N_1818,N_1734);
and U2335 (N_2335,N_1722,N_1843);
and U2336 (N_2336,N_1686,N_1924);
and U2337 (N_2337,N_1966,N_1534);
nor U2338 (N_2338,N_1974,N_1645);
or U2339 (N_2339,N_1501,N_1806);
or U2340 (N_2340,N_1864,N_1881);
and U2341 (N_2341,N_1603,N_1657);
or U2342 (N_2342,N_1862,N_1943);
xnor U2343 (N_2343,N_1579,N_1816);
and U2344 (N_2344,N_1886,N_1690);
and U2345 (N_2345,N_1951,N_1673);
or U2346 (N_2346,N_1837,N_1845);
and U2347 (N_2347,N_1957,N_1543);
or U2348 (N_2348,N_1987,N_1911);
or U2349 (N_2349,N_1742,N_1665);
and U2350 (N_2350,N_1947,N_1536);
nor U2351 (N_2351,N_1501,N_1565);
or U2352 (N_2352,N_1707,N_1974);
nand U2353 (N_2353,N_1787,N_1928);
xor U2354 (N_2354,N_1509,N_1518);
xnor U2355 (N_2355,N_1993,N_1835);
or U2356 (N_2356,N_1566,N_1509);
or U2357 (N_2357,N_1573,N_1916);
nor U2358 (N_2358,N_1625,N_1596);
nand U2359 (N_2359,N_1915,N_1694);
or U2360 (N_2360,N_1974,N_1665);
or U2361 (N_2361,N_1750,N_1891);
and U2362 (N_2362,N_1678,N_1687);
xor U2363 (N_2363,N_1914,N_1545);
nand U2364 (N_2364,N_1605,N_1903);
nand U2365 (N_2365,N_1892,N_1508);
nor U2366 (N_2366,N_1757,N_1626);
nor U2367 (N_2367,N_1567,N_1918);
or U2368 (N_2368,N_1759,N_1914);
xor U2369 (N_2369,N_1744,N_1613);
nand U2370 (N_2370,N_1565,N_1905);
and U2371 (N_2371,N_1709,N_1612);
and U2372 (N_2372,N_1954,N_1622);
xnor U2373 (N_2373,N_1743,N_1985);
nand U2374 (N_2374,N_1687,N_1619);
nand U2375 (N_2375,N_1824,N_1625);
nor U2376 (N_2376,N_1801,N_1527);
and U2377 (N_2377,N_1663,N_1991);
nand U2378 (N_2378,N_1790,N_1590);
nand U2379 (N_2379,N_1992,N_1979);
xnor U2380 (N_2380,N_1603,N_1547);
nand U2381 (N_2381,N_1792,N_1825);
nor U2382 (N_2382,N_1537,N_1864);
and U2383 (N_2383,N_1518,N_1533);
or U2384 (N_2384,N_1938,N_1781);
nor U2385 (N_2385,N_1590,N_1546);
nor U2386 (N_2386,N_1931,N_1693);
nand U2387 (N_2387,N_1676,N_1953);
or U2388 (N_2388,N_1518,N_1908);
nor U2389 (N_2389,N_1999,N_1527);
or U2390 (N_2390,N_1641,N_1599);
and U2391 (N_2391,N_1659,N_1597);
and U2392 (N_2392,N_1586,N_1844);
and U2393 (N_2393,N_1814,N_1787);
and U2394 (N_2394,N_1795,N_1532);
or U2395 (N_2395,N_1509,N_1822);
and U2396 (N_2396,N_1595,N_1868);
and U2397 (N_2397,N_1511,N_1648);
nor U2398 (N_2398,N_1816,N_1903);
or U2399 (N_2399,N_1937,N_1844);
and U2400 (N_2400,N_1923,N_1724);
nand U2401 (N_2401,N_1948,N_1582);
and U2402 (N_2402,N_1952,N_1779);
nor U2403 (N_2403,N_1576,N_1954);
or U2404 (N_2404,N_1945,N_1997);
nand U2405 (N_2405,N_1835,N_1509);
and U2406 (N_2406,N_1997,N_1765);
nor U2407 (N_2407,N_1791,N_1828);
nand U2408 (N_2408,N_1956,N_1539);
nand U2409 (N_2409,N_1558,N_1802);
nor U2410 (N_2410,N_1957,N_1626);
or U2411 (N_2411,N_1997,N_1527);
nor U2412 (N_2412,N_1679,N_1943);
nand U2413 (N_2413,N_1527,N_1841);
xor U2414 (N_2414,N_1878,N_1518);
nor U2415 (N_2415,N_1621,N_1833);
and U2416 (N_2416,N_1791,N_1667);
xor U2417 (N_2417,N_1513,N_1740);
nor U2418 (N_2418,N_1642,N_1566);
xnor U2419 (N_2419,N_1934,N_1539);
nor U2420 (N_2420,N_1932,N_1582);
xnor U2421 (N_2421,N_1838,N_1591);
nor U2422 (N_2422,N_1897,N_1872);
nand U2423 (N_2423,N_1989,N_1837);
nor U2424 (N_2424,N_1630,N_1839);
nand U2425 (N_2425,N_1544,N_1945);
or U2426 (N_2426,N_1608,N_1522);
or U2427 (N_2427,N_1536,N_1881);
xor U2428 (N_2428,N_1770,N_1508);
xnor U2429 (N_2429,N_1862,N_1534);
nand U2430 (N_2430,N_1999,N_1586);
nor U2431 (N_2431,N_1585,N_1672);
and U2432 (N_2432,N_1521,N_1700);
or U2433 (N_2433,N_1705,N_1857);
nand U2434 (N_2434,N_1885,N_1780);
nor U2435 (N_2435,N_1669,N_1889);
or U2436 (N_2436,N_1828,N_1887);
nor U2437 (N_2437,N_1566,N_1731);
or U2438 (N_2438,N_1588,N_1579);
and U2439 (N_2439,N_1584,N_1545);
nor U2440 (N_2440,N_1620,N_1501);
xnor U2441 (N_2441,N_1702,N_1683);
and U2442 (N_2442,N_1628,N_1925);
nand U2443 (N_2443,N_1870,N_1967);
nor U2444 (N_2444,N_1643,N_1917);
nand U2445 (N_2445,N_1550,N_1721);
or U2446 (N_2446,N_1676,N_1771);
nand U2447 (N_2447,N_1961,N_1916);
and U2448 (N_2448,N_1616,N_1965);
or U2449 (N_2449,N_1843,N_1865);
nor U2450 (N_2450,N_1684,N_1836);
or U2451 (N_2451,N_1872,N_1552);
or U2452 (N_2452,N_1774,N_1793);
nor U2453 (N_2453,N_1650,N_1971);
nand U2454 (N_2454,N_1831,N_1980);
xor U2455 (N_2455,N_1517,N_1712);
xor U2456 (N_2456,N_1949,N_1947);
nand U2457 (N_2457,N_1549,N_1660);
nand U2458 (N_2458,N_1748,N_1958);
and U2459 (N_2459,N_1929,N_1785);
nand U2460 (N_2460,N_1806,N_1816);
xor U2461 (N_2461,N_1640,N_1600);
and U2462 (N_2462,N_1669,N_1860);
nand U2463 (N_2463,N_1678,N_1945);
nor U2464 (N_2464,N_1818,N_1707);
nor U2465 (N_2465,N_1747,N_1942);
nand U2466 (N_2466,N_1756,N_1942);
nor U2467 (N_2467,N_1718,N_1962);
and U2468 (N_2468,N_1605,N_1789);
or U2469 (N_2469,N_1880,N_1603);
nor U2470 (N_2470,N_1904,N_1986);
and U2471 (N_2471,N_1639,N_1889);
xnor U2472 (N_2472,N_1977,N_1720);
nand U2473 (N_2473,N_1526,N_1889);
and U2474 (N_2474,N_1856,N_1921);
nand U2475 (N_2475,N_1807,N_1539);
or U2476 (N_2476,N_1938,N_1859);
xor U2477 (N_2477,N_1756,N_1724);
nor U2478 (N_2478,N_1622,N_1704);
or U2479 (N_2479,N_1951,N_1734);
and U2480 (N_2480,N_1630,N_1715);
nor U2481 (N_2481,N_1580,N_1735);
or U2482 (N_2482,N_1644,N_1914);
and U2483 (N_2483,N_1834,N_1862);
nand U2484 (N_2484,N_1584,N_1646);
xor U2485 (N_2485,N_1785,N_1600);
xnor U2486 (N_2486,N_1917,N_1576);
nand U2487 (N_2487,N_1528,N_1958);
nand U2488 (N_2488,N_1948,N_1951);
or U2489 (N_2489,N_1589,N_1675);
nor U2490 (N_2490,N_1808,N_1942);
nand U2491 (N_2491,N_1907,N_1891);
or U2492 (N_2492,N_1519,N_1989);
xor U2493 (N_2493,N_1877,N_1571);
nor U2494 (N_2494,N_1644,N_1886);
nor U2495 (N_2495,N_1632,N_1806);
and U2496 (N_2496,N_1711,N_1828);
nor U2497 (N_2497,N_1865,N_1998);
and U2498 (N_2498,N_1514,N_1766);
or U2499 (N_2499,N_1628,N_1920);
or U2500 (N_2500,N_2021,N_2398);
and U2501 (N_2501,N_2238,N_2289);
or U2502 (N_2502,N_2296,N_2318);
nor U2503 (N_2503,N_2055,N_2427);
xor U2504 (N_2504,N_2388,N_2463);
xor U2505 (N_2505,N_2234,N_2267);
or U2506 (N_2506,N_2032,N_2274);
xnor U2507 (N_2507,N_2310,N_2473);
xor U2508 (N_2508,N_2103,N_2403);
xnor U2509 (N_2509,N_2303,N_2314);
and U2510 (N_2510,N_2038,N_2436);
xor U2511 (N_2511,N_2087,N_2125);
nand U2512 (N_2512,N_2494,N_2379);
or U2513 (N_2513,N_2043,N_2360);
xnor U2514 (N_2514,N_2011,N_2037);
nor U2515 (N_2515,N_2176,N_2340);
xnor U2516 (N_2516,N_2241,N_2257);
nor U2517 (N_2517,N_2299,N_2122);
or U2518 (N_2518,N_2407,N_2025);
xnor U2519 (N_2519,N_2005,N_2181);
nor U2520 (N_2520,N_2266,N_2107);
nor U2521 (N_2521,N_2474,N_2332);
xnor U2522 (N_2522,N_2121,N_2291);
nor U2523 (N_2523,N_2477,N_2232);
and U2524 (N_2524,N_2098,N_2189);
or U2525 (N_2525,N_2116,N_2111);
or U2526 (N_2526,N_2268,N_2183);
or U2527 (N_2527,N_2344,N_2158);
or U2528 (N_2528,N_2129,N_2497);
and U2529 (N_2529,N_2188,N_2182);
nand U2530 (N_2530,N_2109,N_2080);
xor U2531 (N_2531,N_2335,N_2321);
nand U2532 (N_2532,N_2365,N_2012);
and U2533 (N_2533,N_2311,N_2072);
nand U2534 (N_2534,N_2169,N_2399);
nand U2535 (N_2535,N_2465,N_2063);
and U2536 (N_2536,N_2393,N_2480);
nor U2537 (N_2537,N_2148,N_2307);
nand U2538 (N_2538,N_2325,N_2449);
or U2539 (N_2539,N_2155,N_2009);
and U2540 (N_2540,N_2359,N_2269);
nand U2541 (N_2541,N_2294,N_2115);
nor U2542 (N_2542,N_2371,N_2237);
or U2543 (N_2543,N_2434,N_2196);
and U2544 (N_2544,N_2397,N_2442);
or U2545 (N_2545,N_2472,N_2177);
xnor U2546 (N_2546,N_2285,N_2002);
xnor U2547 (N_2547,N_2099,N_2022);
nor U2548 (N_2548,N_2249,N_2230);
xnor U2549 (N_2549,N_2210,N_2225);
xor U2550 (N_2550,N_2271,N_2353);
xor U2551 (N_2551,N_2045,N_2491);
nand U2552 (N_2552,N_2137,N_2418);
and U2553 (N_2553,N_2413,N_2280);
or U2554 (N_2554,N_2165,N_2203);
nand U2555 (N_2555,N_2432,N_2346);
or U2556 (N_2556,N_2251,N_2255);
or U2557 (N_2557,N_2233,N_2488);
or U2558 (N_2558,N_2284,N_2205);
xor U2559 (N_2559,N_2222,N_2097);
nor U2560 (N_2560,N_2263,N_2049);
or U2561 (N_2561,N_2343,N_2164);
xor U2562 (N_2562,N_2133,N_2394);
and U2563 (N_2563,N_2014,N_2179);
nor U2564 (N_2564,N_2034,N_2193);
and U2565 (N_2565,N_2229,N_2059);
or U2566 (N_2566,N_2254,N_2073);
nand U2567 (N_2567,N_2185,N_2486);
or U2568 (N_2568,N_2243,N_2118);
nor U2569 (N_2569,N_2264,N_2157);
nor U2570 (N_2570,N_2101,N_2108);
nand U2571 (N_2571,N_2096,N_2128);
and U2572 (N_2572,N_2020,N_2430);
or U2573 (N_2573,N_2058,N_2240);
or U2574 (N_2574,N_2018,N_2368);
xor U2575 (N_2575,N_2373,N_2172);
nand U2576 (N_2576,N_2408,N_2074);
xor U2577 (N_2577,N_2091,N_2352);
nor U2578 (N_2578,N_2104,N_2161);
nor U2579 (N_2579,N_2057,N_2357);
nor U2580 (N_2580,N_2438,N_2355);
nand U2581 (N_2581,N_2075,N_2410);
nand U2582 (N_2582,N_2035,N_2324);
and U2583 (N_2583,N_2006,N_2351);
and U2584 (N_2584,N_2028,N_2019);
or U2585 (N_2585,N_2208,N_2146);
nor U2586 (N_2586,N_2452,N_2227);
or U2587 (N_2587,N_2275,N_2457);
nand U2588 (N_2588,N_2062,N_2286);
nand U2589 (N_2589,N_2127,N_2278);
or U2590 (N_2590,N_2067,N_2089);
and U2591 (N_2591,N_2455,N_2470);
nand U2592 (N_2592,N_2487,N_2444);
and U2593 (N_2593,N_2242,N_2260);
or U2594 (N_2594,N_2135,N_2202);
nor U2595 (N_2595,N_2467,N_2462);
or U2596 (N_2596,N_2124,N_2126);
xor U2597 (N_2597,N_2295,N_2156);
and U2598 (N_2598,N_2024,N_2342);
xnor U2599 (N_2599,N_2439,N_2380);
xnor U2600 (N_2600,N_2192,N_2117);
and U2601 (N_2601,N_2456,N_2492);
or U2602 (N_2602,N_2315,N_2329);
nand U2603 (N_2603,N_2304,N_2471);
nor U2604 (N_2604,N_2499,N_2419);
nor U2605 (N_2605,N_2458,N_2027);
nor U2606 (N_2606,N_2308,N_2010);
and U2607 (N_2607,N_2207,N_2231);
nand U2608 (N_2608,N_2029,N_2136);
nand U2609 (N_2609,N_2424,N_2114);
nand U2610 (N_2610,N_2498,N_2141);
nor U2611 (N_2611,N_2016,N_2008);
nand U2612 (N_2612,N_2461,N_2190);
nor U2613 (N_2613,N_2253,N_2377);
nand U2614 (N_2614,N_2065,N_2000);
and U2615 (N_2615,N_2212,N_2400);
nor U2616 (N_2616,N_2292,N_2282);
nor U2617 (N_2617,N_2316,N_2123);
or U2618 (N_2618,N_2447,N_2415);
xor U2619 (N_2619,N_2317,N_2036);
xor U2620 (N_2620,N_2453,N_2052);
and U2621 (N_2621,N_2119,N_2330);
nand U2622 (N_2622,N_2152,N_2198);
and U2623 (N_2623,N_2481,N_2175);
nand U2624 (N_2624,N_2451,N_2201);
or U2625 (N_2625,N_2159,N_2184);
xor U2626 (N_2626,N_2478,N_2076);
nand U2627 (N_2627,N_2044,N_2246);
xor U2628 (N_2628,N_2276,N_2160);
xnor U2629 (N_2629,N_2211,N_2250);
nand U2630 (N_2630,N_2079,N_2173);
and U2631 (N_2631,N_2421,N_2390);
or U2632 (N_2632,N_2042,N_2215);
nor U2633 (N_2633,N_2272,N_2445);
xnor U2634 (N_2634,N_2496,N_2077);
nand U2635 (N_2635,N_2088,N_2423);
nand U2636 (N_2636,N_2150,N_2450);
nor U2637 (N_2637,N_2085,N_2223);
xor U2638 (N_2638,N_2358,N_2056);
or U2639 (N_2639,N_2170,N_2139);
or U2640 (N_2640,N_2440,N_2347);
nand U2641 (N_2641,N_2218,N_2209);
nand U2642 (N_2642,N_2300,N_2084);
nor U2643 (N_2643,N_2051,N_2283);
xor U2644 (N_2644,N_2248,N_2206);
or U2645 (N_2645,N_2217,N_2245);
nor U2646 (N_2646,N_2348,N_2328);
xnor U2647 (N_2647,N_2140,N_2092);
or U2648 (N_2648,N_2420,N_2409);
xnor U2649 (N_2649,N_2401,N_2270);
xor U2650 (N_2650,N_2047,N_2171);
nor U2651 (N_2651,N_2252,N_2224);
and U2652 (N_2652,N_2485,N_2383);
or U2653 (N_2653,N_2186,N_2490);
nand U2654 (N_2654,N_2337,N_2138);
and U2655 (N_2655,N_2007,N_2244);
nor U2656 (N_2656,N_2031,N_2093);
nor U2657 (N_2657,N_2100,N_2105);
nor U2658 (N_2658,N_2259,N_2147);
and U2659 (N_2659,N_2066,N_2493);
and U2660 (N_2660,N_2213,N_2441);
and U2661 (N_2661,N_2279,N_2262);
or U2662 (N_2662,N_2195,N_2081);
nand U2663 (N_2663,N_2331,N_2163);
nor U2664 (N_2664,N_2375,N_2130);
nor U2665 (N_2665,N_2338,N_2023);
or U2666 (N_2666,N_2495,N_2306);
nor U2667 (N_2667,N_2443,N_2326);
nor U2668 (N_2668,N_2425,N_2131);
nor U2669 (N_2669,N_2416,N_2341);
nor U2670 (N_2670,N_2194,N_2385);
or U2671 (N_2671,N_2200,N_2017);
or U2672 (N_2672,N_2216,N_2174);
xnor U2673 (N_2673,N_2219,N_2313);
nand U2674 (N_2674,N_2345,N_2053);
and U2675 (N_2675,N_2214,N_2273);
or U2676 (N_2676,N_2149,N_2323);
and U2677 (N_2677,N_2030,N_2336);
and U2678 (N_2678,N_2431,N_2362);
xor U2679 (N_2679,N_2102,N_2144);
nor U2680 (N_2680,N_2113,N_2468);
xnor U2681 (N_2681,N_2327,N_2428);
nor U2682 (N_2682,N_2475,N_2405);
or U2683 (N_2683,N_2142,N_2082);
nand U2684 (N_2684,N_2162,N_2448);
and U2685 (N_2685,N_2277,N_2261);
and U2686 (N_2686,N_2039,N_2460);
or U2687 (N_2687,N_2064,N_2265);
xor U2688 (N_2688,N_2154,N_2466);
nand U2689 (N_2689,N_2435,N_2454);
xor U2690 (N_2690,N_2333,N_2083);
xor U2691 (N_2691,N_2414,N_2001);
nand U2692 (N_2692,N_2290,N_2422);
and U2693 (N_2693,N_2145,N_2363);
or U2694 (N_2694,N_2046,N_2178);
nand U2695 (N_2695,N_2143,N_2287);
xnor U2696 (N_2696,N_2220,N_2361);
or U2697 (N_2697,N_2404,N_2469);
and U2698 (N_2698,N_2464,N_2482);
nor U2699 (N_2699,N_2322,N_2112);
nor U2700 (N_2700,N_2429,N_2086);
nor U2701 (N_2701,N_2204,N_2180);
xor U2702 (N_2702,N_2476,N_2369);
nand U2703 (N_2703,N_2226,N_2256);
or U2704 (N_2704,N_2197,N_2048);
and U2705 (N_2705,N_2281,N_2258);
or U2706 (N_2706,N_2293,N_2372);
nor U2707 (N_2707,N_2134,N_2378);
xnor U2708 (N_2708,N_2026,N_2061);
xor U2709 (N_2709,N_2356,N_2221);
xnor U2710 (N_2710,N_2433,N_2187);
nand U2711 (N_2711,N_2376,N_2367);
and U2712 (N_2712,N_2334,N_2069);
nor U2713 (N_2713,N_2040,N_2349);
and U2714 (N_2714,N_2060,N_2297);
or U2715 (N_2715,N_2120,N_2068);
and U2716 (N_2716,N_2395,N_2396);
xnor U2717 (N_2717,N_2110,N_2391);
nor U2718 (N_2718,N_2191,N_2402);
and U2719 (N_2719,N_2071,N_2090);
nor U2720 (N_2720,N_2312,N_2132);
and U2721 (N_2721,N_2095,N_2054);
xnor U2722 (N_2722,N_2382,N_2320);
and U2723 (N_2723,N_2366,N_2389);
xnor U2724 (N_2724,N_2459,N_2381);
or U2725 (N_2725,N_2288,N_2479);
nor U2726 (N_2726,N_2070,N_2387);
xnor U2727 (N_2727,N_2483,N_2411);
nor U2728 (N_2728,N_2319,N_2151);
xor U2729 (N_2729,N_2106,N_2350);
and U2730 (N_2730,N_2003,N_2484);
nand U2731 (N_2731,N_2033,N_2302);
xor U2732 (N_2732,N_2446,N_2041);
nor U2733 (N_2733,N_2489,N_2412);
or U2734 (N_2734,N_2364,N_2339);
xor U2735 (N_2735,N_2301,N_2392);
nor U2736 (N_2736,N_2417,N_2199);
or U2737 (N_2737,N_2309,N_2384);
nor U2738 (N_2738,N_2050,N_2239);
nand U2739 (N_2739,N_2153,N_2247);
xnor U2740 (N_2740,N_2078,N_2236);
and U2741 (N_2741,N_2228,N_2354);
nor U2742 (N_2742,N_2437,N_2167);
or U2743 (N_2743,N_2235,N_2013);
or U2744 (N_2744,N_2168,N_2298);
or U2745 (N_2745,N_2015,N_2004);
xnor U2746 (N_2746,N_2406,N_2374);
or U2747 (N_2747,N_2426,N_2305);
xnor U2748 (N_2748,N_2370,N_2386);
xnor U2749 (N_2749,N_2094,N_2166);
xor U2750 (N_2750,N_2045,N_2475);
nand U2751 (N_2751,N_2453,N_2070);
nor U2752 (N_2752,N_2395,N_2381);
xor U2753 (N_2753,N_2227,N_2375);
and U2754 (N_2754,N_2123,N_2088);
nand U2755 (N_2755,N_2218,N_2175);
or U2756 (N_2756,N_2364,N_2370);
nor U2757 (N_2757,N_2015,N_2276);
xor U2758 (N_2758,N_2319,N_2081);
nor U2759 (N_2759,N_2437,N_2051);
or U2760 (N_2760,N_2404,N_2175);
or U2761 (N_2761,N_2067,N_2194);
xnor U2762 (N_2762,N_2268,N_2357);
and U2763 (N_2763,N_2290,N_2204);
and U2764 (N_2764,N_2121,N_2460);
or U2765 (N_2765,N_2218,N_2387);
nand U2766 (N_2766,N_2410,N_2246);
nor U2767 (N_2767,N_2029,N_2378);
xor U2768 (N_2768,N_2251,N_2091);
nand U2769 (N_2769,N_2238,N_2171);
nor U2770 (N_2770,N_2449,N_2342);
xnor U2771 (N_2771,N_2223,N_2233);
nand U2772 (N_2772,N_2021,N_2275);
nand U2773 (N_2773,N_2466,N_2036);
nand U2774 (N_2774,N_2064,N_2366);
and U2775 (N_2775,N_2065,N_2102);
nand U2776 (N_2776,N_2201,N_2452);
and U2777 (N_2777,N_2172,N_2226);
nand U2778 (N_2778,N_2120,N_2403);
xor U2779 (N_2779,N_2284,N_2483);
nand U2780 (N_2780,N_2255,N_2040);
and U2781 (N_2781,N_2354,N_2190);
and U2782 (N_2782,N_2253,N_2348);
and U2783 (N_2783,N_2293,N_2170);
or U2784 (N_2784,N_2281,N_2204);
nand U2785 (N_2785,N_2108,N_2475);
nand U2786 (N_2786,N_2239,N_2146);
nand U2787 (N_2787,N_2069,N_2404);
or U2788 (N_2788,N_2023,N_2129);
nand U2789 (N_2789,N_2111,N_2246);
and U2790 (N_2790,N_2286,N_2125);
xor U2791 (N_2791,N_2165,N_2234);
and U2792 (N_2792,N_2316,N_2150);
nor U2793 (N_2793,N_2026,N_2163);
xnor U2794 (N_2794,N_2043,N_2229);
nand U2795 (N_2795,N_2001,N_2016);
or U2796 (N_2796,N_2198,N_2328);
nand U2797 (N_2797,N_2056,N_2399);
xor U2798 (N_2798,N_2297,N_2329);
and U2799 (N_2799,N_2063,N_2110);
nand U2800 (N_2800,N_2117,N_2498);
and U2801 (N_2801,N_2426,N_2085);
or U2802 (N_2802,N_2205,N_2413);
and U2803 (N_2803,N_2074,N_2194);
nand U2804 (N_2804,N_2337,N_2286);
xor U2805 (N_2805,N_2190,N_2260);
or U2806 (N_2806,N_2359,N_2002);
nor U2807 (N_2807,N_2299,N_2111);
nor U2808 (N_2808,N_2118,N_2165);
nor U2809 (N_2809,N_2132,N_2425);
and U2810 (N_2810,N_2287,N_2437);
nor U2811 (N_2811,N_2461,N_2271);
and U2812 (N_2812,N_2033,N_2057);
and U2813 (N_2813,N_2367,N_2014);
and U2814 (N_2814,N_2341,N_2078);
nor U2815 (N_2815,N_2480,N_2384);
nor U2816 (N_2816,N_2413,N_2213);
nand U2817 (N_2817,N_2127,N_2090);
nand U2818 (N_2818,N_2119,N_2394);
and U2819 (N_2819,N_2040,N_2219);
nor U2820 (N_2820,N_2187,N_2499);
and U2821 (N_2821,N_2461,N_2017);
nand U2822 (N_2822,N_2019,N_2219);
xor U2823 (N_2823,N_2399,N_2449);
nand U2824 (N_2824,N_2008,N_2436);
nor U2825 (N_2825,N_2402,N_2238);
nand U2826 (N_2826,N_2050,N_2091);
or U2827 (N_2827,N_2333,N_2315);
nor U2828 (N_2828,N_2437,N_2050);
xor U2829 (N_2829,N_2132,N_2354);
nand U2830 (N_2830,N_2010,N_2136);
xor U2831 (N_2831,N_2108,N_2463);
nand U2832 (N_2832,N_2262,N_2253);
and U2833 (N_2833,N_2495,N_2284);
xnor U2834 (N_2834,N_2255,N_2277);
and U2835 (N_2835,N_2119,N_2495);
nor U2836 (N_2836,N_2471,N_2299);
or U2837 (N_2837,N_2060,N_2107);
or U2838 (N_2838,N_2320,N_2209);
nand U2839 (N_2839,N_2188,N_2326);
nand U2840 (N_2840,N_2499,N_2183);
xnor U2841 (N_2841,N_2440,N_2333);
nand U2842 (N_2842,N_2001,N_2254);
nor U2843 (N_2843,N_2427,N_2109);
or U2844 (N_2844,N_2045,N_2498);
and U2845 (N_2845,N_2073,N_2068);
nand U2846 (N_2846,N_2173,N_2346);
or U2847 (N_2847,N_2195,N_2263);
and U2848 (N_2848,N_2144,N_2183);
and U2849 (N_2849,N_2062,N_2449);
nand U2850 (N_2850,N_2077,N_2450);
and U2851 (N_2851,N_2216,N_2097);
and U2852 (N_2852,N_2192,N_2450);
or U2853 (N_2853,N_2482,N_2183);
xor U2854 (N_2854,N_2126,N_2097);
and U2855 (N_2855,N_2473,N_2362);
nand U2856 (N_2856,N_2209,N_2431);
nand U2857 (N_2857,N_2159,N_2391);
nor U2858 (N_2858,N_2036,N_2429);
nand U2859 (N_2859,N_2194,N_2467);
nor U2860 (N_2860,N_2126,N_2276);
nand U2861 (N_2861,N_2422,N_2406);
xor U2862 (N_2862,N_2084,N_2350);
nor U2863 (N_2863,N_2302,N_2242);
and U2864 (N_2864,N_2250,N_2055);
nor U2865 (N_2865,N_2498,N_2407);
and U2866 (N_2866,N_2230,N_2224);
and U2867 (N_2867,N_2409,N_2067);
or U2868 (N_2868,N_2138,N_2202);
nand U2869 (N_2869,N_2121,N_2227);
xnor U2870 (N_2870,N_2453,N_2102);
and U2871 (N_2871,N_2064,N_2458);
nand U2872 (N_2872,N_2095,N_2368);
nor U2873 (N_2873,N_2375,N_2422);
and U2874 (N_2874,N_2217,N_2182);
and U2875 (N_2875,N_2247,N_2385);
and U2876 (N_2876,N_2469,N_2113);
and U2877 (N_2877,N_2434,N_2375);
nor U2878 (N_2878,N_2061,N_2031);
nand U2879 (N_2879,N_2235,N_2193);
nor U2880 (N_2880,N_2103,N_2355);
or U2881 (N_2881,N_2415,N_2474);
nand U2882 (N_2882,N_2420,N_2126);
xnor U2883 (N_2883,N_2140,N_2249);
xnor U2884 (N_2884,N_2286,N_2081);
xor U2885 (N_2885,N_2246,N_2274);
xor U2886 (N_2886,N_2484,N_2057);
or U2887 (N_2887,N_2042,N_2475);
and U2888 (N_2888,N_2218,N_2324);
or U2889 (N_2889,N_2093,N_2042);
and U2890 (N_2890,N_2458,N_2018);
nor U2891 (N_2891,N_2302,N_2308);
nand U2892 (N_2892,N_2372,N_2381);
or U2893 (N_2893,N_2016,N_2291);
xor U2894 (N_2894,N_2133,N_2246);
and U2895 (N_2895,N_2122,N_2057);
xnor U2896 (N_2896,N_2457,N_2050);
nor U2897 (N_2897,N_2148,N_2029);
nand U2898 (N_2898,N_2031,N_2430);
and U2899 (N_2899,N_2275,N_2232);
nand U2900 (N_2900,N_2497,N_2464);
and U2901 (N_2901,N_2332,N_2427);
and U2902 (N_2902,N_2320,N_2123);
nand U2903 (N_2903,N_2439,N_2445);
or U2904 (N_2904,N_2478,N_2469);
nand U2905 (N_2905,N_2228,N_2319);
or U2906 (N_2906,N_2419,N_2335);
and U2907 (N_2907,N_2123,N_2214);
or U2908 (N_2908,N_2494,N_2093);
nor U2909 (N_2909,N_2284,N_2322);
and U2910 (N_2910,N_2328,N_2111);
nor U2911 (N_2911,N_2260,N_2476);
or U2912 (N_2912,N_2343,N_2211);
and U2913 (N_2913,N_2486,N_2310);
or U2914 (N_2914,N_2123,N_2197);
nor U2915 (N_2915,N_2217,N_2236);
or U2916 (N_2916,N_2080,N_2163);
or U2917 (N_2917,N_2448,N_2076);
xor U2918 (N_2918,N_2067,N_2190);
nand U2919 (N_2919,N_2061,N_2332);
nor U2920 (N_2920,N_2184,N_2458);
xnor U2921 (N_2921,N_2024,N_2335);
nand U2922 (N_2922,N_2210,N_2120);
or U2923 (N_2923,N_2051,N_2053);
xnor U2924 (N_2924,N_2092,N_2185);
or U2925 (N_2925,N_2284,N_2349);
xnor U2926 (N_2926,N_2036,N_2424);
or U2927 (N_2927,N_2111,N_2028);
xnor U2928 (N_2928,N_2151,N_2183);
and U2929 (N_2929,N_2432,N_2343);
xor U2930 (N_2930,N_2374,N_2163);
or U2931 (N_2931,N_2406,N_2046);
or U2932 (N_2932,N_2089,N_2164);
or U2933 (N_2933,N_2296,N_2474);
nor U2934 (N_2934,N_2007,N_2156);
xor U2935 (N_2935,N_2171,N_2174);
or U2936 (N_2936,N_2111,N_2379);
nand U2937 (N_2937,N_2309,N_2103);
nand U2938 (N_2938,N_2435,N_2380);
or U2939 (N_2939,N_2376,N_2296);
xor U2940 (N_2940,N_2460,N_2462);
nor U2941 (N_2941,N_2099,N_2357);
nand U2942 (N_2942,N_2245,N_2371);
xor U2943 (N_2943,N_2058,N_2052);
nor U2944 (N_2944,N_2088,N_2322);
xor U2945 (N_2945,N_2200,N_2423);
nor U2946 (N_2946,N_2030,N_2338);
nor U2947 (N_2947,N_2456,N_2022);
xnor U2948 (N_2948,N_2422,N_2040);
or U2949 (N_2949,N_2281,N_2431);
and U2950 (N_2950,N_2347,N_2290);
and U2951 (N_2951,N_2288,N_2145);
nand U2952 (N_2952,N_2181,N_2251);
nand U2953 (N_2953,N_2470,N_2304);
nand U2954 (N_2954,N_2251,N_2311);
nand U2955 (N_2955,N_2120,N_2479);
nand U2956 (N_2956,N_2197,N_2286);
nor U2957 (N_2957,N_2451,N_2115);
nor U2958 (N_2958,N_2393,N_2141);
nor U2959 (N_2959,N_2300,N_2006);
and U2960 (N_2960,N_2114,N_2385);
and U2961 (N_2961,N_2304,N_2090);
or U2962 (N_2962,N_2309,N_2119);
xor U2963 (N_2963,N_2261,N_2009);
nor U2964 (N_2964,N_2177,N_2036);
and U2965 (N_2965,N_2120,N_2198);
and U2966 (N_2966,N_2447,N_2025);
and U2967 (N_2967,N_2173,N_2024);
nand U2968 (N_2968,N_2488,N_2235);
nand U2969 (N_2969,N_2170,N_2028);
xor U2970 (N_2970,N_2395,N_2420);
nand U2971 (N_2971,N_2355,N_2443);
and U2972 (N_2972,N_2257,N_2091);
and U2973 (N_2973,N_2172,N_2179);
xnor U2974 (N_2974,N_2008,N_2004);
xor U2975 (N_2975,N_2340,N_2366);
nor U2976 (N_2976,N_2339,N_2075);
nand U2977 (N_2977,N_2210,N_2002);
nor U2978 (N_2978,N_2449,N_2217);
and U2979 (N_2979,N_2141,N_2478);
xor U2980 (N_2980,N_2494,N_2015);
nand U2981 (N_2981,N_2033,N_2006);
nor U2982 (N_2982,N_2144,N_2398);
xnor U2983 (N_2983,N_2485,N_2102);
xnor U2984 (N_2984,N_2200,N_2178);
nor U2985 (N_2985,N_2174,N_2404);
or U2986 (N_2986,N_2099,N_2389);
nand U2987 (N_2987,N_2487,N_2173);
and U2988 (N_2988,N_2097,N_2065);
xnor U2989 (N_2989,N_2252,N_2438);
or U2990 (N_2990,N_2089,N_2360);
nor U2991 (N_2991,N_2205,N_2190);
or U2992 (N_2992,N_2426,N_2176);
nor U2993 (N_2993,N_2277,N_2473);
nand U2994 (N_2994,N_2344,N_2212);
nor U2995 (N_2995,N_2260,N_2212);
nor U2996 (N_2996,N_2246,N_2148);
or U2997 (N_2997,N_2466,N_2376);
xor U2998 (N_2998,N_2065,N_2424);
nor U2999 (N_2999,N_2429,N_2488);
xor U3000 (N_3000,N_2519,N_2982);
nor U3001 (N_3001,N_2606,N_2694);
nor U3002 (N_3002,N_2575,N_2605);
and U3003 (N_3003,N_2507,N_2699);
or U3004 (N_3004,N_2763,N_2845);
nand U3005 (N_3005,N_2535,N_2934);
or U3006 (N_3006,N_2895,N_2750);
nand U3007 (N_3007,N_2928,N_2715);
xnor U3008 (N_3008,N_2508,N_2511);
xor U3009 (N_3009,N_2565,N_2783);
nand U3010 (N_3010,N_2992,N_2604);
or U3011 (N_3011,N_2995,N_2587);
or U3012 (N_3012,N_2899,N_2903);
or U3013 (N_3013,N_2680,N_2601);
nor U3014 (N_3014,N_2527,N_2850);
nand U3015 (N_3015,N_2720,N_2521);
and U3016 (N_3016,N_2738,N_2512);
and U3017 (N_3017,N_2517,N_2647);
or U3018 (N_3018,N_2841,N_2842);
nor U3019 (N_3019,N_2536,N_2724);
or U3020 (N_3020,N_2893,N_2655);
nor U3021 (N_3021,N_2642,N_2759);
and U3022 (N_3022,N_2676,N_2758);
nand U3023 (N_3023,N_2843,N_2986);
and U3024 (N_3024,N_2876,N_2697);
or U3025 (N_3025,N_2579,N_2892);
or U3026 (N_3026,N_2945,N_2785);
xor U3027 (N_3027,N_2765,N_2645);
nand U3028 (N_3028,N_2959,N_2880);
or U3029 (N_3029,N_2650,N_2796);
xnor U3030 (N_3030,N_2518,N_2701);
xor U3031 (N_3031,N_2526,N_2746);
nor U3032 (N_3032,N_2853,N_2687);
nor U3033 (N_3033,N_2585,N_2635);
nand U3034 (N_3034,N_2716,N_2848);
or U3035 (N_3035,N_2626,N_2686);
or U3036 (N_3036,N_2714,N_2542);
nor U3037 (N_3037,N_2778,N_2979);
nor U3038 (N_3038,N_2797,N_2833);
and U3039 (N_3039,N_2523,N_2669);
and U3040 (N_3040,N_2677,N_2886);
nand U3041 (N_3041,N_2855,N_2742);
or U3042 (N_3042,N_2832,N_2564);
nor U3043 (N_3043,N_2577,N_2653);
xnor U3044 (N_3044,N_2980,N_2555);
nor U3045 (N_3045,N_2904,N_2621);
and U3046 (N_3046,N_2811,N_2780);
xnor U3047 (N_3047,N_2978,N_2702);
nor U3048 (N_3048,N_2516,N_2703);
nor U3049 (N_3049,N_2556,N_2709);
xnor U3050 (N_3050,N_2840,N_2639);
or U3051 (N_3051,N_2659,N_2788);
or U3052 (N_3052,N_2533,N_2905);
or U3053 (N_3053,N_2509,N_2771);
xnor U3054 (N_3054,N_2551,N_2953);
nand U3055 (N_3055,N_2752,N_2657);
or U3056 (N_3056,N_2926,N_2863);
nor U3057 (N_3057,N_2884,N_2641);
nand U3058 (N_3058,N_2524,N_2736);
xor U3059 (N_3059,N_2543,N_2662);
or U3060 (N_3060,N_2914,N_2705);
and U3061 (N_3061,N_2902,N_2737);
nand U3062 (N_3062,N_2938,N_2611);
nor U3063 (N_3063,N_2515,N_2908);
and U3064 (N_3064,N_2830,N_2948);
nor U3065 (N_3065,N_2751,N_2671);
xor U3066 (N_3066,N_2609,N_2782);
and U3067 (N_3067,N_2727,N_2890);
nand U3068 (N_3068,N_2648,N_2970);
or U3069 (N_3069,N_2695,N_2915);
nand U3070 (N_3070,N_2576,N_2802);
and U3071 (N_3071,N_2907,N_2733);
nand U3072 (N_3072,N_2891,N_2969);
and U3073 (N_3073,N_2731,N_2897);
nand U3074 (N_3074,N_2949,N_2722);
nor U3075 (N_3075,N_2916,N_2684);
and U3076 (N_3076,N_2827,N_2568);
nor U3077 (N_3077,N_2852,N_2723);
or U3078 (N_3078,N_2660,N_2933);
or U3079 (N_3079,N_2944,N_2719);
nor U3080 (N_3080,N_2644,N_2779);
xor U3081 (N_3081,N_2814,N_2688);
nor U3082 (N_3082,N_2947,N_2707);
nand U3083 (N_3083,N_2623,N_2822);
nand U3084 (N_3084,N_2966,N_2839);
and U3085 (N_3085,N_2559,N_2756);
or U3086 (N_3086,N_2667,N_2652);
nor U3087 (N_3087,N_2844,N_2968);
nand U3088 (N_3088,N_2955,N_2815);
nand U3089 (N_3089,N_2627,N_2991);
nor U3090 (N_3090,N_2889,N_2962);
xnor U3091 (N_3091,N_2630,N_2794);
and U3092 (N_3092,N_2696,N_2808);
nand U3093 (N_3093,N_2874,N_2825);
xnor U3094 (N_3094,N_2504,N_2624);
or U3095 (N_3095,N_2574,N_2898);
nor U3096 (N_3096,N_2540,N_2869);
nand U3097 (N_3097,N_2865,N_2739);
or U3098 (N_3098,N_2649,N_2821);
and U3099 (N_3099,N_2681,N_2856);
or U3100 (N_3100,N_2679,N_2525);
xor U3101 (N_3101,N_2589,N_2793);
xnor U3102 (N_3102,N_2580,N_2646);
nor U3103 (N_3103,N_2661,N_2810);
xnor U3104 (N_3104,N_2761,N_2996);
nor U3105 (N_3105,N_2885,N_2954);
xor U3106 (N_3106,N_2873,N_2981);
and U3107 (N_3107,N_2625,N_2666);
xnor U3108 (N_3108,N_2561,N_2729);
xnor U3109 (N_3109,N_2633,N_2762);
or U3110 (N_3110,N_2673,N_2552);
nor U3111 (N_3111,N_2665,N_2870);
xnor U3112 (N_3112,N_2861,N_2741);
or U3113 (N_3113,N_2867,N_2730);
nand U3114 (N_3114,N_2828,N_2920);
or U3115 (N_3115,N_2501,N_2813);
and U3116 (N_3116,N_2610,N_2569);
or U3117 (N_3117,N_2941,N_2940);
nor U3118 (N_3118,N_2603,N_2913);
and U3119 (N_3119,N_2790,N_2997);
xor U3120 (N_3120,N_2859,N_2951);
nor U3121 (N_3121,N_2983,N_2616);
nor U3122 (N_3122,N_2798,N_2961);
and U3123 (N_3123,N_2860,N_2789);
nand U3124 (N_3124,N_2994,N_2573);
nor U3125 (N_3125,N_2682,N_2857);
and U3126 (N_3126,N_2943,N_2834);
or U3127 (N_3127,N_2503,N_2998);
and U3128 (N_3128,N_2692,N_2956);
nor U3129 (N_3129,N_2967,N_2987);
nor U3130 (N_3130,N_2831,N_2529);
nor U3131 (N_3131,N_2977,N_2505);
or U3132 (N_3132,N_2767,N_2749);
nor U3133 (N_3133,N_2562,N_2755);
and U3134 (N_3134,N_2617,N_2612);
xor U3135 (N_3135,N_2823,N_2868);
and U3136 (N_3136,N_2999,N_2598);
nor U3137 (N_3137,N_2544,N_2989);
and U3138 (N_3138,N_2651,N_2917);
nor U3139 (N_3139,N_2952,N_2957);
nor U3140 (N_3140,N_2541,N_2964);
nor U3141 (N_3141,N_2528,N_2613);
nor U3142 (N_3142,N_2781,N_2777);
nor U3143 (N_3143,N_2689,N_2620);
nand U3144 (N_3144,N_2801,N_2805);
nand U3145 (N_3145,N_2924,N_2818);
nand U3146 (N_3146,N_2710,N_2545);
or U3147 (N_3147,N_2608,N_2939);
or U3148 (N_3148,N_2872,N_2965);
and U3149 (N_3149,N_2974,N_2764);
nor U3150 (N_3150,N_2851,N_2592);
nor U3151 (N_3151,N_2600,N_2614);
and U3152 (N_3152,N_2734,N_2618);
nand U3153 (N_3153,N_2837,N_2588);
or U3154 (N_3154,N_2849,N_2572);
nand U3155 (N_3155,N_2550,N_2718);
and U3156 (N_3156,N_2975,N_2942);
nor U3157 (N_3157,N_2786,N_2678);
nor U3158 (N_3158,N_2776,N_2829);
and U3159 (N_3159,N_2583,N_2819);
and U3160 (N_3160,N_2950,N_2634);
and U3161 (N_3161,N_2591,N_2946);
or U3162 (N_3162,N_2602,N_2932);
or U3163 (N_3163,N_2988,N_2862);
nor U3164 (N_3164,N_2882,N_2704);
nor U3165 (N_3165,N_2663,N_2721);
nor U3166 (N_3166,N_2958,N_2735);
xor U3167 (N_3167,N_2976,N_2748);
xnor U3168 (N_3168,N_2581,N_2522);
nand U3169 (N_3169,N_2792,N_2510);
or U3170 (N_3170,N_2520,N_2769);
xor U3171 (N_3171,N_2875,N_2675);
or U3172 (N_3172,N_2570,N_2768);
and U3173 (N_3173,N_2566,N_2700);
nor U3174 (N_3174,N_2803,N_2685);
xnor U3175 (N_3175,N_2791,N_2910);
xor U3176 (N_3176,N_2674,N_2846);
nor U3177 (N_3177,N_2773,N_2547);
and U3178 (N_3178,N_2717,N_2930);
nand U3179 (N_3179,N_2909,N_2732);
and U3180 (N_3180,N_2972,N_2726);
xor U3181 (N_3181,N_2753,N_2963);
and U3182 (N_3182,N_2935,N_2537);
or U3183 (N_3183,N_2921,N_2539);
nor U3184 (N_3184,N_2668,N_2877);
xnor U3185 (N_3185,N_2772,N_2854);
nor U3186 (N_3186,N_2593,N_2806);
xor U3187 (N_3187,N_2900,N_2643);
or U3188 (N_3188,N_2774,N_2725);
xnor U3189 (N_3189,N_2858,N_2927);
nand U3190 (N_3190,N_2812,N_2881);
nor U3191 (N_3191,N_2629,N_2925);
or U3192 (N_3192,N_2538,N_2637);
nand U3193 (N_3193,N_2595,N_2800);
and U3194 (N_3194,N_2984,N_2607);
and U3195 (N_3195,N_2936,N_2864);
or U3196 (N_3196,N_2747,N_2632);
xnor U3197 (N_3197,N_2912,N_2919);
nand U3198 (N_3198,N_2622,N_2766);
or U3199 (N_3199,N_2658,N_2824);
or U3200 (N_3200,N_2582,N_2578);
and U3201 (N_3201,N_2656,N_2754);
xor U3202 (N_3202,N_2549,N_2514);
nand U3203 (N_3203,N_2553,N_2871);
or U3204 (N_3204,N_2971,N_2636);
and U3205 (N_3205,N_2728,N_2670);
nand U3206 (N_3206,N_2596,N_2590);
nand U3207 (N_3207,N_2619,N_2787);
or U3208 (N_3208,N_2554,N_2804);
nand U3209 (N_3209,N_2502,N_2799);
nand U3210 (N_3210,N_2664,N_2548);
or U3211 (N_3211,N_2615,N_2513);
and U3212 (N_3212,N_2532,N_2698);
xor U3213 (N_3213,N_2557,N_2929);
or U3214 (N_3214,N_2817,N_2847);
xor U3215 (N_3215,N_2993,N_2960);
nor U3216 (N_3216,N_2683,N_2745);
nor U3217 (N_3217,N_2631,N_2571);
nor U3218 (N_3218,N_2923,N_2584);
or U3219 (N_3219,N_2879,N_2628);
nand U3220 (N_3220,N_2937,N_2807);
or U3221 (N_3221,N_2836,N_2567);
nand U3222 (N_3222,N_2534,N_2896);
nor U3223 (N_3223,N_2784,N_2693);
and U3224 (N_3224,N_2638,N_2531);
nor U3225 (N_3225,N_2597,N_2560);
or U3226 (N_3226,N_2888,N_2558);
or U3227 (N_3227,N_2713,N_2712);
and U3228 (N_3228,N_2654,N_2599);
and U3229 (N_3229,N_2586,N_2922);
xor U3230 (N_3230,N_2795,N_2706);
nand U3231 (N_3231,N_2826,N_2866);
or U3232 (N_3232,N_2820,N_2743);
or U3233 (N_3233,N_2894,N_2887);
nand U3234 (N_3234,N_2760,N_2985);
xor U3235 (N_3235,N_2838,N_2640);
xor U3236 (N_3236,N_2816,N_2563);
nor U3237 (N_3237,N_2906,N_2672);
or U3238 (N_3238,N_2883,N_2973);
nand U3239 (N_3239,N_2775,N_2546);
nand U3240 (N_3240,N_2918,N_2500);
nand U3241 (N_3241,N_2744,N_2506);
nand U3242 (N_3242,N_2594,N_2708);
or U3243 (N_3243,N_2809,N_2878);
nor U3244 (N_3244,N_2690,N_2740);
or U3245 (N_3245,N_2911,N_2931);
xnor U3246 (N_3246,N_2530,N_2901);
nor U3247 (N_3247,N_2990,N_2711);
nor U3248 (N_3248,N_2835,N_2770);
xor U3249 (N_3249,N_2691,N_2757);
and U3250 (N_3250,N_2849,N_2895);
nand U3251 (N_3251,N_2873,N_2915);
xnor U3252 (N_3252,N_2609,N_2704);
nand U3253 (N_3253,N_2823,N_2610);
xor U3254 (N_3254,N_2658,N_2537);
nand U3255 (N_3255,N_2573,N_2705);
xor U3256 (N_3256,N_2778,N_2863);
and U3257 (N_3257,N_2919,N_2837);
nor U3258 (N_3258,N_2767,N_2727);
or U3259 (N_3259,N_2904,N_2539);
nand U3260 (N_3260,N_2563,N_2922);
or U3261 (N_3261,N_2834,N_2696);
nand U3262 (N_3262,N_2903,N_2598);
nor U3263 (N_3263,N_2739,N_2771);
nand U3264 (N_3264,N_2738,N_2630);
nand U3265 (N_3265,N_2611,N_2998);
xor U3266 (N_3266,N_2778,N_2836);
nor U3267 (N_3267,N_2520,N_2662);
xor U3268 (N_3268,N_2597,N_2868);
nand U3269 (N_3269,N_2741,N_2600);
nand U3270 (N_3270,N_2528,N_2591);
xnor U3271 (N_3271,N_2589,N_2911);
nor U3272 (N_3272,N_2625,N_2929);
nand U3273 (N_3273,N_2735,N_2881);
xor U3274 (N_3274,N_2570,N_2798);
nand U3275 (N_3275,N_2518,N_2993);
nand U3276 (N_3276,N_2857,N_2876);
or U3277 (N_3277,N_2683,N_2641);
nand U3278 (N_3278,N_2950,N_2821);
nor U3279 (N_3279,N_2587,N_2853);
nand U3280 (N_3280,N_2895,N_2721);
nand U3281 (N_3281,N_2813,N_2594);
nand U3282 (N_3282,N_2906,N_2552);
nor U3283 (N_3283,N_2648,N_2933);
and U3284 (N_3284,N_2906,N_2842);
nor U3285 (N_3285,N_2942,N_2555);
xor U3286 (N_3286,N_2719,N_2982);
and U3287 (N_3287,N_2825,N_2785);
or U3288 (N_3288,N_2989,N_2928);
or U3289 (N_3289,N_2847,N_2650);
and U3290 (N_3290,N_2951,N_2700);
or U3291 (N_3291,N_2736,N_2542);
nor U3292 (N_3292,N_2932,N_2936);
and U3293 (N_3293,N_2792,N_2833);
and U3294 (N_3294,N_2965,N_2754);
nor U3295 (N_3295,N_2749,N_2947);
and U3296 (N_3296,N_2671,N_2878);
nor U3297 (N_3297,N_2652,N_2811);
nand U3298 (N_3298,N_2623,N_2520);
xor U3299 (N_3299,N_2769,N_2567);
or U3300 (N_3300,N_2759,N_2646);
nor U3301 (N_3301,N_2584,N_2939);
nor U3302 (N_3302,N_2516,N_2951);
or U3303 (N_3303,N_2932,N_2789);
or U3304 (N_3304,N_2598,N_2883);
nor U3305 (N_3305,N_2554,N_2711);
xnor U3306 (N_3306,N_2739,N_2734);
nor U3307 (N_3307,N_2795,N_2703);
or U3308 (N_3308,N_2976,N_2614);
nor U3309 (N_3309,N_2584,N_2609);
nor U3310 (N_3310,N_2658,N_2784);
or U3311 (N_3311,N_2787,N_2941);
xnor U3312 (N_3312,N_2670,N_2873);
or U3313 (N_3313,N_2935,N_2870);
nor U3314 (N_3314,N_2860,N_2714);
xnor U3315 (N_3315,N_2847,N_2669);
nor U3316 (N_3316,N_2732,N_2538);
and U3317 (N_3317,N_2994,N_2585);
nor U3318 (N_3318,N_2995,N_2734);
xor U3319 (N_3319,N_2884,N_2865);
and U3320 (N_3320,N_2771,N_2663);
xnor U3321 (N_3321,N_2663,N_2735);
xnor U3322 (N_3322,N_2644,N_2674);
nor U3323 (N_3323,N_2841,N_2837);
and U3324 (N_3324,N_2713,N_2860);
and U3325 (N_3325,N_2955,N_2678);
nor U3326 (N_3326,N_2594,N_2508);
and U3327 (N_3327,N_2750,N_2681);
and U3328 (N_3328,N_2713,N_2700);
or U3329 (N_3329,N_2846,N_2875);
and U3330 (N_3330,N_2733,N_2832);
xor U3331 (N_3331,N_2807,N_2650);
nand U3332 (N_3332,N_2505,N_2543);
and U3333 (N_3333,N_2727,N_2936);
xor U3334 (N_3334,N_2797,N_2684);
nand U3335 (N_3335,N_2664,N_2740);
or U3336 (N_3336,N_2808,N_2686);
nor U3337 (N_3337,N_2794,N_2698);
xor U3338 (N_3338,N_2679,N_2964);
and U3339 (N_3339,N_2899,N_2790);
or U3340 (N_3340,N_2658,N_2742);
nand U3341 (N_3341,N_2732,N_2950);
or U3342 (N_3342,N_2614,N_2681);
xor U3343 (N_3343,N_2986,N_2688);
or U3344 (N_3344,N_2782,N_2537);
or U3345 (N_3345,N_2561,N_2607);
and U3346 (N_3346,N_2658,N_2571);
xnor U3347 (N_3347,N_2685,N_2520);
nor U3348 (N_3348,N_2903,N_2850);
or U3349 (N_3349,N_2986,N_2752);
nor U3350 (N_3350,N_2914,N_2926);
or U3351 (N_3351,N_2711,N_2687);
or U3352 (N_3352,N_2745,N_2580);
nand U3353 (N_3353,N_2885,N_2685);
and U3354 (N_3354,N_2646,N_2542);
nor U3355 (N_3355,N_2945,N_2593);
and U3356 (N_3356,N_2671,N_2777);
nor U3357 (N_3357,N_2870,N_2791);
and U3358 (N_3358,N_2515,N_2896);
xnor U3359 (N_3359,N_2638,N_2976);
nand U3360 (N_3360,N_2714,N_2929);
and U3361 (N_3361,N_2657,N_2723);
nand U3362 (N_3362,N_2506,N_2798);
nand U3363 (N_3363,N_2756,N_2527);
nor U3364 (N_3364,N_2889,N_2603);
and U3365 (N_3365,N_2764,N_2534);
nand U3366 (N_3366,N_2997,N_2641);
or U3367 (N_3367,N_2982,N_2962);
xnor U3368 (N_3368,N_2916,N_2986);
nand U3369 (N_3369,N_2789,N_2541);
and U3370 (N_3370,N_2665,N_2940);
nand U3371 (N_3371,N_2604,N_2978);
nand U3372 (N_3372,N_2709,N_2687);
and U3373 (N_3373,N_2665,N_2632);
nand U3374 (N_3374,N_2665,N_2920);
nand U3375 (N_3375,N_2947,N_2592);
xnor U3376 (N_3376,N_2798,N_2871);
nor U3377 (N_3377,N_2891,N_2702);
or U3378 (N_3378,N_2975,N_2851);
nor U3379 (N_3379,N_2837,N_2992);
xor U3380 (N_3380,N_2849,N_2816);
or U3381 (N_3381,N_2969,N_2953);
nand U3382 (N_3382,N_2750,N_2838);
xnor U3383 (N_3383,N_2635,N_2762);
and U3384 (N_3384,N_2969,N_2934);
nor U3385 (N_3385,N_2712,N_2631);
xnor U3386 (N_3386,N_2509,N_2911);
and U3387 (N_3387,N_2863,N_2829);
nand U3388 (N_3388,N_2511,N_2862);
nand U3389 (N_3389,N_2818,N_2798);
and U3390 (N_3390,N_2533,N_2525);
nand U3391 (N_3391,N_2677,N_2641);
xnor U3392 (N_3392,N_2916,N_2958);
and U3393 (N_3393,N_2746,N_2821);
xnor U3394 (N_3394,N_2739,N_2569);
nand U3395 (N_3395,N_2660,N_2890);
xnor U3396 (N_3396,N_2694,N_2896);
nand U3397 (N_3397,N_2932,N_2806);
xor U3398 (N_3398,N_2580,N_2784);
nor U3399 (N_3399,N_2624,N_2838);
and U3400 (N_3400,N_2903,N_2796);
nor U3401 (N_3401,N_2561,N_2638);
nand U3402 (N_3402,N_2660,N_2932);
and U3403 (N_3403,N_2916,N_2819);
xnor U3404 (N_3404,N_2545,N_2503);
nand U3405 (N_3405,N_2505,N_2684);
xnor U3406 (N_3406,N_2638,N_2862);
and U3407 (N_3407,N_2500,N_2871);
xnor U3408 (N_3408,N_2615,N_2999);
and U3409 (N_3409,N_2808,N_2781);
nor U3410 (N_3410,N_2962,N_2600);
and U3411 (N_3411,N_2517,N_2963);
or U3412 (N_3412,N_2558,N_2504);
and U3413 (N_3413,N_2842,N_2643);
nor U3414 (N_3414,N_2667,N_2801);
xnor U3415 (N_3415,N_2774,N_2787);
nor U3416 (N_3416,N_2671,N_2540);
nor U3417 (N_3417,N_2812,N_2870);
or U3418 (N_3418,N_2599,N_2673);
and U3419 (N_3419,N_2725,N_2957);
xor U3420 (N_3420,N_2560,N_2765);
nor U3421 (N_3421,N_2966,N_2799);
xor U3422 (N_3422,N_2961,N_2514);
and U3423 (N_3423,N_2587,N_2854);
nor U3424 (N_3424,N_2541,N_2834);
and U3425 (N_3425,N_2538,N_2761);
or U3426 (N_3426,N_2890,N_2655);
xnor U3427 (N_3427,N_2548,N_2904);
nand U3428 (N_3428,N_2903,N_2875);
nand U3429 (N_3429,N_2741,N_2763);
nand U3430 (N_3430,N_2671,N_2749);
or U3431 (N_3431,N_2808,N_2801);
nor U3432 (N_3432,N_2511,N_2514);
and U3433 (N_3433,N_2873,N_2991);
and U3434 (N_3434,N_2514,N_2706);
xnor U3435 (N_3435,N_2512,N_2863);
nand U3436 (N_3436,N_2923,N_2956);
or U3437 (N_3437,N_2623,N_2506);
or U3438 (N_3438,N_2855,N_2609);
xnor U3439 (N_3439,N_2981,N_2694);
nor U3440 (N_3440,N_2940,N_2711);
nand U3441 (N_3441,N_2618,N_2879);
or U3442 (N_3442,N_2650,N_2793);
xnor U3443 (N_3443,N_2804,N_2961);
and U3444 (N_3444,N_2657,N_2572);
xor U3445 (N_3445,N_2944,N_2887);
nor U3446 (N_3446,N_2867,N_2795);
and U3447 (N_3447,N_2729,N_2972);
nor U3448 (N_3448,N_2873,N_2767);
nand U3449 (N_3449,N_2949,N_2770);
and U3450 (N_3450,N_2506,N_2973);
nor U3451 (N_3451,N_2894,N_2891);
nor U3452 (N_3452,N_2912,N_2586);
nor U3453 (N_3453,N_2688,N_2941);
and U3454 (N_3454,N_2550,N_2603);
nor U3455 (N_3455,N_2509,N_2851);
or U3456 (N_3456,N_2976,N_2779);
nand U3457 (N_3457,N_2836,N_2942);
nand U3458 (N_3458,N_2760,N_2955);
or U3459 (N_3459,N_2874,N_2579);
nor U3460 (N_3460,N_2569,N_2789);
and U3461 (N_3461,N_2937,N_2633);
or U3462 (N_3462,N_2774,N_2944);
nand U3463 (N_3463,N_2642,N_2574);
nor U3464 (N_3464,N_2706,N_2658);
and U3465 (N_3465,N_2779,N_2771);
and U3466 (N_3466,N_2892,N_2832);
or U3467 (N_3467,N_2953,N_2758);
nand U3468 (N_3468,N_2686,N_2552);
nor U3469 (N_3469,N_2835,N_2848);
nor U3470 (N_3470,N_2573,N_2847);
nor U3471 (N_3471,N_2824,N_2921);
and U3472 (N_3472,N_2767,N_2929);
xnor U3473 (N_3473,N_2913,N_2993);
nor U3474 (N_3474,N_2688,N_2994);
and U3475 (N_3475,N_2893,N_2777);
nand U3476 (N_3476,N_2884,N_2577);
xor U3477 (N_3477,N_2513,N_2843);
nor U3478 (N_3478,N_2643,N_2905);
and U3479 (N_3479,N_2700,N_2542);
and U3480 (N_3480,N_2766,N_2571);
nor U3481 (N_3481,N_2798,N_2811);
nand U3482 (N_3482,N_2783,N_2806);
and U3483 (N_3483,N_2623,N_2982);
nor U3484 (N_3484,N_2941,N_2624);
nand U3485 (N_3485,N_2766,N_2947);
and U3486 (N_3486,N_2784,N_2884);
nand U3487 (N_3487,N_2818,N_2901);
nor U3488 (N_3488,N_2917,N_2965);
and U3489 (N_3489,N_2990,N_2843);
nand U3490 (N_3490,N_2877,N_2584);
or U3491 (N_3491,N_2592,N_2682);
xnor U3492 (N_3492,N_2841,N_2532);
nor U3493 (N_3493,N_2996,N_2618);
and U3494 (N_3494,N_2704,N_2954);
nand U3495 (N_3495,N_2998,N_2720);
and U3496 (N_3496,N_2815,N_2757);
and U3497 (N_3497,N_2999,N_2503);
xnor U3498 (N_3498,N_2816,N_2832);
nor U3499 (N_3499,N_2824,N_2624);
nor U3500 (N_3500,N_3115,N_3038);
or U3501 (N_3501,N_3257,N_3211);
or U3502 (N_3502,N_3084,N_3204);
nor U3503 (N_3503,N_3300,N_3382);
or U3504 (N_3504,N_3367,N_3111);
xor U3505 (N_3505,N_3030,N_3215);
or U3506 (N_3506,N_3416,N_3096);
and U3507 (N_3507,N_3010,N_3076);
and U3508 (N_3508,N_3092,N_3279);
and U3509 (N_3509,N_3481,N_3091);
or U3510 (N_3510,N_3389,N_3171);
or U3511 (N_3511,N_3289,N_3477);
or U3512 (N_3512,N_3060,N_3338);
nand U3513 (N_3513,N_3404,N_3241);
nor U3514 (N_3514,N_3445,N_3292);
or U3515 (N_3515,N_3497,N_3230);
and U3516 (N_3516,N_3028,N_3455);
nor U3517 (N_3517,N_3427,N_3400);
or U3518 (N_3518,N_3363,N_3244);
nor U3519 (N_3519,N_3172,N_3434);
or U3520 (N_3520,N_3381,N_3272);
nor U3521 (N_3521,N_3008,N_3044);
or U3522 (N_3522,N_3418,N_3261);
or U3523 (N_3523,N_3366,N_3225);
and U3524 (N_3524,N_3001,N_3190);
or U3525 (N_3525,N_3208,N_3488);
nand U3526 (N_3526,N_3471,N_3324);
xnor U3527 (N_3527,N_3331,N_3240);
or U3528 (N_3528,N_3407,N_3080);
and U3529 (N_3529,N_3421,N_3387);
and U3530 (N_3530,N_3436,N_3000);
nand U3531 (N_3531,N_3212,N_3026);
and U3532 (N_3532,N_3413,N_3169);
xnor U3533 (N_3533,N_3121,N_3016);
nand U3534 (N_3534,N_3068,N_3368);
xnor U3535 (N_3535,N_3403,N_3365);
and U3536 (N_3536,N_3429,N_3057);
and U3537 (N_3537,N_3414,N_3317);
xnor U3538 (N_3538,N_3428,N_3247);
and U3539 (N_3539,N_3491,N_3105);
nand U3540 (N_3540,N_3276,N_3246);
or U3541 (N_3541,N_3461,N_3263);
nand U3542 (N_3542,N_3320,N_3290);
xor U3543 (N_3543,N_3487,N_3219);
or U3544 (N_3544,N_3165,N_3166);
and U3545 (N_3545,N_3144,N_3405);
nand U3546 (N_3546,N_3378,N_3055);
and U3547 (N_3547,N_3221,N_3447);
nor U3548 (N_3548,N_3117,N_3262);
xnor U3549 (N_3549,N_3102,N_3081);
nand U3550 (N_3550,N_3056,N_3475);
nand U3551 (N_3551,N_3371,N_3451);
and U3552 (N_3552,N_3256,N_3196);
or U3553 (N_3553,N_3438,N_3316);
nor U3554 (N_3554,N_3299,N_3385);
xor U3555 (N_3555,N_3229,N_3499);
nand U3556 (N_3556,N_3234,N_3329);
xnor U3557 (N_3557,N_3003,N_3350);
xor U3558 (N_3558,N_3192,N_3349);
or U3559 (N_3559,N_3213,N_3138);
or U3560 (N_3560,N_3067,N_3151);
or U3561 (N_3561,N_3280,N_3089);
or U3562 (N_3562,N_3189,N_3046);
xor U3563 (N_3563,N_3128,N_3082);
nand U3564 (N_3564,N_3162,N_3402);
xor U3565 (N_3565,N_3069,N_3452);
or U3566 (N_3566,N_3109,N_3342);
or U3567 (N_3567,N_3195,N_3489);
xor U3568 (N_3568,N_3254,N_3410);
or U3569 (N_3569,N_3129,N_3466);
xor U3570 (N_3570,N_3090,N_3355);
nor U3571 (N_3571,N_3168,N_3012);
nor U3572 (N_3572,N_3137,N_3399);
nor U3573 (N_3573,N_3291,N_3142);
and U3574 (N_3574,N_3269,N_3116);
xor U3575 (N_3575,N_3470,N_3446);
xor U3576 (N_3576,N_3043,N_3153);
and U3577 (N_3577,N_3275,N_3130);
or U3578 (N_3578,N_3145,N_3025);
xor U3579 (N_3579,N_3235,N_3053);
xor U3580 (N_3580,N_3268,N_3370);
nor U3581 (N_3581,N_3435,N_3424);
nor U3582 (N_3582,N_3174,N_3449);
or U3583 (N_3583,N_3075,N_3364);
and U3584 (N_3584,N_3163,N_3126);
xor U3585 (N_3585,N_3267,N_3388);
or U3586 (N_3586,N_3356,N_3217);
or U3587 (N_3587,N_3431,N_3274);
or U3588 (N_3588,N_3415,N_3238);
or U3589 (N_3589,N_3253,N_3372);
nand U3590 (N_3590,N_3188,N_3191);
or U3591 (N_3591,N_3397,N_3018);
xnor U3592 (N_3592,N_3140,N_3223);
or U3593 (N_3593,N_3401,N_3309);
xor U3594 (N_3594,N_3118,N_3343);
or U3595 (N_3595,N_3311,N_3353);
nor U3596 (N_3596,N_3002,N_3373);
xor U3597 (N_3597,N_3377,N_3178);
or U3598 (N_3598,N_3450,N_3303);
nor U3599 (N_3599,N_3218,N_3333);
nand U3600 (N_3600,N_3308,N_3265);
nand U3601 (N_3601,N_3301,N_3182);
or U3602 (N_3602,N_3341,N_3017);
or U3603 (N_3603,N_3304,N_3061);
nand U3604 (N_3604,N_3490,N_3095);
xnor U3605 (N_3605,N_3348,N_3085);
nand U3606 (N_3606,N_3019,N_3480);
nor U3607 (N_3607,N_3205,N_3143);
and U3608 (N_3608,N_3242,N_3478);
nor U3609 (N_3609,N_3336,N_3245);
xnor U3610 (N_3610,N_3408,N_3023);
or U3611 (N_3611,N_3045,N_3332);
nor U3612 (N_3612,N_3237,N_3009);
and U3613 (N_3613,N_3422,N_3031);
xnor U3614 (N_3614,N_3058,N_3131);
or U3615 (N_3615,N_3093,N_3136);
nor U3616 (N_3616,N_3209,N_3305);
nand U3617 (N_3617,N_3285,N_3286);
and U3618 (N_3618,N_3006,N_3134);
xor U3619 (N_3619,N_3078,N_3119);
nand U3620 (N_3620,N_3203,N_3443);
xnor U3621 (N_3621,N_3393,N_3398);
or U3622 (N_3622,N_3411,N_3176);
or U3623 (N_3623,N_3351,N_3439);
and U3624 (N_3624,N_3049,N_3179);
nor U3625 (N_3625,N_3486,N_3050);
xor U3626 (N_3626,N_3098,N_3214);
and U3627 (N_3627,N_3493,N_3123);
or U3628 (N_3628,N_3295,N_3374);
or U3629 (N_3629,N_3483,N_3062);
nand U3630 (N_3630,N_3457,N_3021);
or U3631 (N_3631,N_3231,N_3150);
or U3632 (N_3632,N_3187,N_3484);
xnor U3633 (N_3633,N_3120,N_3482);
nand U3634 (N_3634,N_3141,N_3395);
and U3635 (N_3635,N_3432,N_3233);
xor U3636 (N_3636,N_3158,N_3293);
and U3637 (N_3637,N_3250,N_3236);
xnor U3638 (N_3638,N_3194,N_3032);
and U3639 (N_3639,N_3206,N_3015);
nor U3640 (N_3640,N_3321,N_3073);
or U3641 (N_3641,N_3177,N_3359);
or U3642 (N_3642,N_3281,N_3306);
or U3643 (N_3643,N_3464,N_3456);
and U3644 (N_3644,N_3079,N_3252);
nor U3645 (N_3645,N_3040,N_3148);
nand U3646 (N_3646,N_3270,N_3054);
nor U3647 (N_3647,N_3059,N_3051);
or U3648 (N_3648,N_3284,N_3347);
or U3649 (N_3649,N_3334,N_3201);
or U3650 (N_3650,N_3264,N_3282);
xor U3651 (N_3651,N_3227,N_3048);
nor U3652 (N_3652,N_3330,N_3473);
nor U3653 (N_3653,N_3394,N_3135);
nor U3654 (N_3654,N_3440,N_3161);
or U3655 (N_3655,N_3226,N_3022);
and U3656 (N_3656,N_3034,N_3094);
or U3657 (N_3657,N_3107,N_3114);
nand U3658 (N_3658,N_3020,N_3271);
xor U3659 (N_3659,N_3088,N_3033);
nand U3660 (N_3660,N_3083,N_3035);
nand U3661 (N_3661,N_3072,N_3185);
nand U3662 (N_3662,N_3492,N_3390);
nand U3663 (N_3663,N_3152,N_3360);
nor U3664 (N_3664,N_3474,N_3243);
nor U3665 (N_3665,N_3070,N_3318);
nor U3666 (N_3666,N_3175,N_3024);
nand U3667 (N_3667,N_3322,N_3124);
nor U3668 (N_3668,N_3065,N_3354);
xor U3669 (N_3669,N_3479,N_3409);
nor U3670 (N_3670,N_3296,N_3104);
and U3671 (N_3671,N_3005,N_3122);
nand U3672 (N_3672,N_3251,N_3287);
or U3673 (N_3673,N_3127,N_3004);
and U3674 (N_3674,N_3392,N_3071);
or U3675 (N_3675,N_3183,N_3278);
nor U3676 (N_3676,N_3323,N_3232);
nand U3677 (N_3677,N_3228,N_3302);
nand U3678 (N_3678,N_3462,N_3426);
xor U3679 (N_3679,N_3294,N_3042);
xnor U3680 (N_3680,N_3326,N_3222);
or U3681 (N_3681,N_3346,N_3260);
xor U3682 (N_3682,N_3448,N_3463);
xor U3683 (N_3683,N_3277,N_3248);
or U3684 (N_3684,N_3039,N_3200);
xor U3685 (N_3685,N_3273,N_3467);
nor U3686 (N_3686,N_3014,N_3027);
nor U3687 (N_3687,N_3412,N_3159);
or U3688 (N_3688,N_3101,N_3146);
nand U3689 (N_3689,N_3207,N_3425);
or U3690 (N_3690,N_3312,N_3454);
and U3691 (N_3691,N_3315,N_3186);
and U3692 (N_3692,N_3103,N_3419);
and U3693 (N_3693,N_3314,N_3327);
nand U3694 (N_3694,N_3406,N_3224);
xnor U3695 (N_3695,N_3197,N_3384);
xnor U3696 (N_3696,N_3340,N_3074);
or U3697 (N_3697,N_3011,N_3444);
nand U3698 (N_3698,N_3379,N_3202);
nor U3699 (N_3699,N_3173,N_3193);
or U3700 (N_3700,N_3157,N_3249);
nand U3701 (N_3701,N_3077,N_3459);
nor U3702 (N_3702,N_3441,N_3259);
xnor U3703 (N_3703,N_3112,N_3437);
nor U3704 (N_3704,N_3132,N_3352);
nand U3705 (N_3705,N_3258,N_3066);
xor U3706 (N_3706,N_3494,N_3375);
nor U3707 (N_3707,N_3430,N_3433);
xor U3708 (N_3708,N_3472,N_3380);
and U3709 (N_3709,N_3149,N_3335);
or U3710 (N_3710,N_3007,N_3154);
and U3711 (N_3711,N_3339,N_3041);
nor U3712 (N_3712,N_3337,N_3198);
xor U3713 (N_3713,N_3052,N_3458);
nor U3714 (N_3714,N_3139,N_3216);
or U3715 (N_3715,N_3199,N_3167);
xnor U3716 (N_3716,N_3013,N_3113);
or U3717 (N_3717,N_3106,N_3417);
nor U3718 (N_3718,N_3170,N_3180);
nor U3719 (N_3719,N_3255,N_3133);
xnor U3720 (N_3720,N_3362,N_3220);
nand U3721 (N_3721,N_3376,N_3160);
nand U3722 (N_3722,N_3476,N_3063);
nor U3723 (N_3723,N_3156,N_3086);
and U3724 (N_3724,N_3239,N_3453);
nor U3725 (N_3725,N_3099,N_3029);
or U3726 (N_3726,N_3361,N_3344);
and U3727 (N_3727,N_3036,N_3047);
xor U3728 (N_3728,N_3108,N_3420);
xnor U3729 (N_3729,N_3423,N_3442);
or U3730 (N_3730,N_3496,N_3210);
nand U3731 (N_3731,N_3110,N_3100);
nor U3732 (N_3732,N_3460,N_3184);
nor U3733 (N_3733,N_3147,N_3383);
nand U3734 (N_3734,N_3310,N_3325);
xnor U3735 (N_3735,N_3386,N_3495);
xor U3736 (N_3736,N_3485,N_3465);
nor U3737 (N_3737,N_3097,N_3266);
nor U3738 (N_3738,N_3064,N_3357);
xor U3739 (N_3739,N_3396,N_3468);
nor U3740 (N_3740,N_3313,N_3288);
nor U3741 (N_3741,N_3164,N_3037);
or U3742 (N_3742,N_3298,N_3369);
xnor U3743 (N_3743,N_3283,N_3391);
and U3744 (N_3744,N_3358,N_3087);
nor U3745 (N_3745,N_3297,N_3345);
nor U3746 (N_3746,N_3469,N_3125);
xnor U3747 (N_3747,N_3498,N_3328);
and U3748 (N_3748,N_3319,N_3155);
xnor U3749 (N_3749,N_3181,N_3307);
or U3750 (N_3750,N_3435,N_3472);
or U3751 (N_3751,N_3171,N_3413);
or U3752 (N_3752,N_3357,N_3473);
nand U3753 (N_3753,N_3223,N_3060);
and U3754 (N_3754,N_3003,N_3017);
nor U3755 (N_3755,N_3316,N_3362);
nand U3756 (N_3756,N_3242,N_3137);
or U3757 (N_3757,N_3391,N_3264);
nor U3758 (N_3758,N_3189,N_3302);
and U3759 (N_3759,N_3289,N_3264);
nand U3760 (N_3760,N_3426,N_3049);
or U3761 (N_3761,N_3462,N_3160);
nor U3762 (N_3762,N_3472,N_3406);
or U3763 (N_3763,N_3450,N_3193);
or U3764 (N_3764,N_3091,N_3021);
or U3765 (N_3765,N_3081,N_3293);
and U3766 (N_3766,N_3361,N_3210);
nand U3767 (N_3767,N_3305,N_3249);
and U3768 (N_3768,N_3239,N_3122);
nand U3769 (N_3769,N_3021,N_3167);
or U3770 (N_3770,N_3035,N_3335);
or U3771 (N_3771,N_3469,N_3311);
nand U3772 (N_3772,N_3352,N_3339);
and U3773 (N_3773,N_3361,N_3369);
nor U3774 (N_3774,N_3215,N_3304);
or U3775 (N_3775,N_3110,N_3048);
nand U3776 (N_3776,N_3092,N_3468);
xnor U3777 (N_3777,N_3392,N_3030);
or U3778 (N_3778,N_3333,N_3395);
nand U3779 (N_3779,N_3444,N_3418);
or U3780 (N_3780,N_3414,N_3402);
or U3781 (N_3781,N_3008,N_3178);
xnor U3782 (N_3782,N_3476,N_3146);
and U3783 (N_3783,N_3491,N_3313);
and U3784 (N_3784,N_3170,N_3387);
xnor U3785 (N_3785,N_3181,N_3059);
nor U3786 (N_3786,N_3437,N_3197);
and U3787 (N_3787,N_3131,N_3469);
nor U3788 (N_3788,N_3137,N_3116);
xnor U3789 (N_3789,N_3044,N_3359);
nand U3790 (N_3790,N_3480,N_3219);
nor U3791 (N_3791,N_3097,N_3046);
nand U3792 (N_3792,N_3199,N_3475);
nor U3793 (N_3793,N_3399,N_3030);
xor U3794 (N_3794,N_3014,N_3174);
nor U3795 (N_3795,N_3283,N_3436);
xor U3796 (N_3796,N_3421,N_3423);
and U3797 (N_3797,N_3293,N_3202);
nand U3798 (N_3798,N_3433,N_3408);
nor U3799 (N_3799,N_3204,N_3300);
or U3800 (N_3800,N_3135,N_3428);
or U3801 (N_3801,N_3105,N_3319);
or U3802 (N_3802,N_3407,N_3218);
or U3803 (N_3803,N_3402,N_3296);
and U3804 (N_3804,N_3063,N_3299);
nor U3805 (N_3805,N_3124,N_3429);
and U3806 (N_3806,N_3018,N_3413);
xor U3807 (N_3807,N_3370,N_3343);
nor U3808 (N_3808,N_3335,N_3129);
xnor U3809 (N_3809,N_3235,N_3021);
xor U3810 (N_3810,N_3321,N_3487);
nor U3811 (N_3811,N_3000,N_3246);
or U3812 (N_3812,N_3248,N_3355);
nor U3813 (N_3813,N_3437,N_3461);
nand U3814 (N_3814,N_3075,N_3435);
nor U3815 (N_3815,N_3110,N_3196);
and U3816 (N_3816,N_3391,N_3021);
or U3817 (N_3817,N_3412,N_3487);
and U3818 (N_3818,N_3052,N_3043);
nand U3819 (N_3819,N_3060,N_3402);
xor U3820 (N_3820,N_3025,N_3254);
and U3821 (N_3821,N_3443,N_3113);
nor U3822 (N_3822,N_3298,N_3004);
and U3823 (N_3823,N_3386,N_3313);
xnor U3824 (N_3824,N_3060,N_3099);
and U3825 (N_3825,N_3430,N_3241);
or U3826 (N_3826,N_3247,N_3345);
nor U3827 (N_3827,N_3346,N_3489);
xor U3828 (N_3828,N_3391,N_3073);
xnor U3829 (N_3829,N_3022,N_3385);
and U3830 (N_3830,N_3024,N_3394);
nand U3831 (N_3831,N_3497,N_3072);
and U3832 (N_3832,N_3012,N_3480);
nand U3833 (N_3833,N_3212,N_3395);
nand U3834 (N_3834,N_3247,N_3432);
and U3835 (N_3835,N_3485,N_3267);
and U3836 (N_3836,N_3450,N_3098);
xnor U3837 (N_3837,N_3449,N_3127);
nand U3838 (N_3838,N_3300,N_3165);
or U3839 (N_3839,N_3445,N_3158);
and U3840 (N_3840,N_3161,N_3054);
nand U3841 (N_3841,N_3379,N_3288);
nand U3842 (N_3842,N_3088,N_3468);
and U3843 (N_3843,N_3146,N_3329);
nand U3844 (N_3844,N_3063,N_3099);
nor U3845 (N_3845,N_3460,N_3242);
nand U3846 (N_3846,N_3138,N_3019);
xnor U3847 (N_3847,N_3177,N_3217);
nor U3848 (N_3848,N_3020,N_3094);
and U3849 (N_3849,N_3228,N_3077);
or U3850 (N_3850,N_3434,N_3402);
nor U3851 (N_3851,N_3132,N_3488);
nand U3852 (N_3852,N_3324,N_3237);
nor U3853 (N_3853,N_3182,N_3414);
or U3854 (N_3854,N_3382,N_3338);
and U3855 (N_3855,N_3039,N_3005);
nand U3856 (N_3856,N_3134,N_3105);
nand U3857 (N_3857,N_3105,N_3367);
or U3858 (N_3858,N_3192,N_3043);
xor U3859 (N_3859,N_3279,N_3126);
xnor U3860 (N_3860,N_3254,N_3296);
and U3861 (N_3861,N_3493,N_3093);
nor U3862 (N_3862,N_3460,N_3152);
xnor U3863 (N_3863,N_3354,N_3039);
or U3864 (N_3864,N_3446,N_3118);
nor U3865 (N_3865,N_3355,N_3233);
or U3866 (N_3866,N_3159,N_3240);
and U3867 (N_3867,N_3497,N_3360);
nand U3868 (N_3868,N_3397,N_3173);
nand U3869 (N_3869,N_3364,N_3045);
nand U3870 (N_3870,N_3336,N_3173);
nand U3871 (N_3871,N_3435,N_3338);
nor U3872 (N_3872,N_3028,N_3415);
xnor U3873 (N_3873,N_3092,N_3253);
or U3874 (N_3874,N_3198,N_3292);
and U3875 (N_3875,N_3249,N_3352);
or U3876 (N_3876,N_3112,N_3036);
and U3877 (N_3877,N_3302,N_3491);
and U3878 (N_3878,N_3318,N_3321);
xor U3879 (N_3879,N_3125,N_3189);
nor U3880 (N_3880,N_3055,N_3052);
and U3881 (N_3881,N_3098,N_3000);
nor U3882 (N_3882,N_3435,N_3073);
and U3883 (N_3883,N_3303,N_3318);
nor U3884 (N_3884,N_3022,N_3332);
nand U3885 (N_3885,N_3464,N_3127);
nor U3886 (N_3886,N_3319,N_3461);
nor U3887 (N_3887,N_3347,N_3409);
nor U3888 (N_3888,N_3141,N_3104);
nand U3889 (N_3889,N_3211,N_3078);
and U3890 (N_3890,N_3132,N_3415);
nor U3891 (N_3891,N_3184,N_3261);
nand U3892 (N_3892,N_3266,N_3304);
nor U3893 (N_3893,N_3247,N_3097);
nor U3894 (N_3894,N_3492,N_3073);
or U3895 (N_3895,N_3219,N_3400);
nand U3896 (N_3896,N_3185,N_3379);
nor U3897 (N_3897,N_3049,N_3029);
and U3898 (N_3898,N_3138,N_3336);
or U3899 (N_3899,N_3178,N_3254);
nand U3900 (N_3900,N_3047,N_3066);
or U3901 (N_3901,N_3468,N_3266);
or U3902 (N_3902,N_3065,N_3453);
and U3903 (N_3903,N_3366,N_3213);
or U3904 (N_3904,N_3487,N_3401);
xnor U3905 (N_3905,N_3256,N_3372);
nand U3906 (N_3906,N_3365,N_3234);
nand U3907 (N_3907,N_3104,N_3048);
and U3908 (N_3908,N_3431,N_3367);
or U3909 (N_3909,N_3170,N_3492);
xor U3910 (N_3910,N_3306,N_3031);
nor U3911 (N_3911,N_3006,N_3020);
nand U3912 (N_3912,N_3476,N_3243);
and U3913 (N_3913,N_3347,N_3489);
xor U3914 (N_3914,N_3313,N_3317);
and U3915 (N_3915,N_3258,N_3290);
nor U3916 (N_3916,N_3323,N_3134);
xor U3917 (N_3917,N_3209,N_3493);
xnor U3918 (N_3918,N_3098,N_3108);
nor U3919 (N_3919,N_3213,N_3379);
xnor U3920 (N_3920,N_3357,N_3337);
or U3921 (N_3921,N_3136,N_3137);
nand U3922 (N_3922,N_3171,N_3264);
and U3923 (N_3923,N_3084,N_3028);
nand U3924 (N_3924,N_3477,N_3022);
nor U3925 (N_3925,N_3145,N_3356);
nand U3926 (N_3926,N_3351,N_3011);
xor U3927 (N_3927,N_3122,N_3493);
nand U3928 (N_3928,N_3467,N_3498);
and U3929 (N_3929,N_3320,N_3356);
nand U3930 (N_3930,N_3187,N_3241);
xor U3931 (N_3931,N_3148,N_3030);
nand U3932 (N_3932,N_3272,N_3495);
xor U3933 (N_3933,N_3268,N_3050);
nor U3934 (N_3934,N_3143,N_3307);
nand U3935 (N_3935,N_3270,N_3138);
nor U3936 (N_3936,N_3220,N_3045);
or U3937 (N_3937,N_3455,N_3272);
or U3938 (N_3938,N_3472,N_3014);
or U3939 (N_3939,N_3476,N_3445);
and U3940 (N_3940,N_3267,N_3192);
xor U3941 (N_3941,N_3121,N_3064);
nand U3942 (N_3942,N_3032,N_3110);
and U3943 (N_3943,N_3468,N_3308);
xnor U3944 (N_3944,N_3309,N_3282);
nor U3945 (N_3945,N_3097,N_3434);
nor U3946 (N_3946,N_3274,N_3081);
xor U3947 (N_3947,N_3173,N_3105);
nand U3948 (N_3948,N_3019,N_3454);
xnor U3949 (N_3949,N_3424,N_3129);
or U3950 (N_3950,N_3297,N_3431);
xor U3951 (N_3951,N_3066,N_3380);
and U3952 (N_3952,N_3417,N_3353);
or U3953 (N_3953,N_3265,N_3446);
and U3954 (N_3954,N_3429,N_3477);
and U3955 (N_3955,N_3316,N_3386);
nor U3956 (N_3956,N_3465,N_3496);
nand U3957 (N_3957,N_3223,N_3181);
nand U3958 (N_3958,N_3298,N_3219);
nand U3959 (N_3959,N_3287,N_3090);
and U3960 (N_3960,N_3064,N_3247);
or U3961 (N_3961,N_3073,N_3199);
nand U3962 (N_3962,N_3356,N_3305);
or U3963 (N_3963,N_3139,N_3111);
nor U3964 (N_3964,N_3073,N_3420);
and U3965 (N_3965,N_3474,N_3004);
or U3966 (N_3966,N_3414,N_3430);
nor U3967 (N_3967,N_3388,N_3018);
nor U3968 (N_3968,N_3472,N_3193);
nand U3969 (N_3969,N_3487,N_3180);
or U3970 (N_3970,N_3313,N_3051);
xnor U3971 (N_3971,N_3237,N_3266);
nand U3972 (N_3972,N_3428,N_3200);
nand U3973 (N_3973,N_3132,N_3192);
and U3974 (N_3974,N_3082,N_3366);
nor U3975 (N_3975,N_3485,N_3147);
nor U3976 (N_3976,N_3472,N_3192);
and U3977 (N_3977,N_3165,N_3065);
and U3978 (N_3978,N_3022,N_3323);
xnor U3979 (N_3979,N_3207,N_3342);
and U3980 (N_3980,N_3087,N_3322);
and U3981 (N_3981,N_3165,N_3332);
xor U3982 (N_3982,N_3127,N_3403);
nand U3983 (N_3983,N_3397,N_3435);
nand U3984 (N_3984,N_3278,N_3160);
nand U3985 (N_3985,N_3112,N_3163);
or U3986 (N_3986,N_3004,N_3070);
nor U3987 (N_3987,N_3456,N_3229);
xor U3988 (N_3988,N_3095,N_3017);
and U3989 (N_3989,N_3165,N_3142);
or U3990 (N_3990,N_3491,N_3022);
xor U3991 (N_3991,N_3392,N_3231);
xnor U3992 (N_3992,N_3030,N_3277);
nor U3993 (N_3993,N_3205,N_3241);
xnor U3994 (N_3994,N_3380,N_3235);
nand U3995 (N_3995,N_3405,N_3412);
nand U3996 (N_3996,N_3394,N_3458);
and U3997 (N_3997,N_3200,N_3122);
or U3998 (N_3998,N_3031,N_3356);
and U3999 (N_3999,N_3239,N_3418);
and U4000 (N_4000,N_3902,N_3810);
nor U4001 (N_4001,N_3583,N_3764);
nand U4002 (N_4002,N_3646,N_3659);
and U4003 (N_4003,N_3808,N_3844);
nand U4004 (N_4004,N_3788,N_3536);
or U4005 (N_4005,N_3688,N_3930);
and U4006 (N_4006,N_3949,N_3801);
or U4007 (N_4007,N_3819,N_3911);
xnor U4008 (N_4008,N_3685,N_3709);
and U4009 (N_4009,N_3824,N_3775);
nand U4010 (N_4010,N_3779,N_3891);
xnor U4011 (N_4011,N_3777,N_3848);
xnor U4012 (N_4012,N_3741,N_3521);
xor U4013 (N_4013,N_3763,N_3768);
or U4014 (N_4014,N_3816,N_3931);
nand U4015 (N_4015,N_3580,N_3554);
and U4016 (N_4016,N_3660,N_3898);
and U4017 (N_4017,N_3956,N_3613);
or U4018 (N_4018,N_3591,N_3915);
and U4019 (N_4019,N_3622,N_3597);
nand U4020 (N_4020,N_3952,N_3705);
nor U4021 (N_4021,N_3567,N_3562);
and U4022 (N_4022,N_3720,N_3714);
nor U4023 (N_4023,N_3890,N_3595);
xor U4024 (N_4024,N_3652,N_3617);
nor U4025 (N_4025,N_3608,N_3811);
nand U4026 (N_4026,N_3533,N_3612);
xnor U4027 (N_4027,N_3843,N_3860);
or U4028 (N_4028,N_3570,N_3852);
and U4029 (N_4029,N_3537,N_3731);
and U4030 (N_4030,N_3706,N_3624);
nor U4031 (N_4031,N_3657,N_3512);
or U4032 (N_4032,N_3627,N_3557);
nor U4033 (N_4033,N_3614,N_3663);
nand U4034 (N_4034,N_3680,N_3851);
nand U4035 (N_4035,N_3645,N_3888);
or U4036 (N_4036,N_3935,N_3918);
and U4037 (N_4037,N_3710,N_3563);
and U4038 (N_4038,N_3750,N_3500);
xor U4039 (N_4039,N_3787,N_3826);
xnor U4040 (N_4040,N_3699,N_3618);
nand U4041 (N_4041,N_3790,N_3603);
and U4042 (N_4042,N_3789,N_3671);
nand U4043 (N_4043,N_3670,N_3786);
and U4044 (N_4044,N_3944,N_3961);
or U4045 (N_4045,N_3867,N_3765);
nand U4046 (N_4046,N_3859,N_3982);
xor U4047 (N_4047,N_3996,N_3964);
or U4048 (N_4048,N_3782,N_3637);
nand U4049 (N_4049,N_3836,N_3780);
nand U4050 (N_4050,N_3629,N_3650);
nor U4051 (N_4051,N_3544,N_3739);
or U4052 (N_4052,N_3639,N_3821);
nor U4053 (N_4053,N_3559,N_3529);
and U4054 (N_4054,N_3887,N_3980);
nand U4055 (N_4055,N_3674,N_3774);
and U4056 (N_4056,N_3968,N_3736);
and U4057 (N_4057,N_3681,N_3534);
or U4058 (N_4058,N_3885,N_3511);
or U4059 (N_4059,N_3679,N_3927);
xor U4060 (N_4060,N_3701,N_3879);
xnor U4061 (N_4061,N_3505,N_3740);
xor U4062 (N_4062,N_3545,N_3815);
nand U4063 (N_4063,N_3984,N_3926);
and U4064 (N_4064,N_3526,N_3566);
and U4065 (N_4065,N_3732,N_3593);
and U4066 (N_4066,N_3516,N_3835);
and U4067 (N_4067,N_3905,N_3582);
nor U4068 (N_4068,N_3793,N_3542);
nand U4069 (N_4069,N_3507,N_3753);
and U4070 (N_4070,N_3895,N_3623);
nor U4071 (N_4071,N_3937,N_3920);
nand U4072 (N_4072,N_3643,N_3922);
or U4073 (N_4073,N_3503,N_3619);
xnor U4074 (N_4074,N_3576,N_3609);
xnor U4075 (N_4075,N_3543,N_3717);
and U4076 (N_4076,N_3708,N_3584);
or U4077 (N_4077,N_3880,N_3822);
nor U4078 (N_4078,N_3812,N_3606);
nand U4079 (N_4079,N_3676,N_3939);
or U4080 (N_4080,N_3572,N_3738);
nand U4081 (N_4081,N_3658,N_3721);
and U4082 (N_4082,N_3995,N_3615);
and U4083 (N_4083,N_3901,N_3551);
or U4084 (N_4084,N_3975,N_3745);
nor U4085 (N_4085,N_3669,N_3501);
or U4086 (N_4086,N_3522,N_3625);
nor U4087 (N_4087,N_3938,N_3587);
nand U4088 (N_4088,N_3550,N_3517);
and U4089 (N_4089,N_3635,N_3698);
nand U4090 (N_4090,N_3896,N_3831);
nand U4091 (N_4091,N_3766,N_3571);
or U4092 (N_4092,N_3713,N_3735);
or U4093 (N_4093,N_3675,N_3596);
or U4094 (N_4094,N_3771,N_3796);
or U4095 (N_4095,N_3729,N_3588);
and U4096 (N_4096,N_3894,N_3523);
xnor U4097 (N_4097,N_3820,N_3702);
and U4098 (N_4098,N_3600,N_3838);
nor U4099 (N_4099,N_3797,N_3904);
or U4100 (N_4100,N_3513,N_3751);
nand U4101 (N_4101,N_3866,N_3954);
and U4102 (N_4102,N_3707,N_3863);
nand U4103 (N_4103,N_3997,N_3578);
or U4104 (N_4104,N_3704,N_3683);
or U4105 (N_4105,N_3743,N_3502);
nor U4106 (N_4106,N_3966,N_3817);
and U4107 (N_4107,N_3940,N_3869);
xor U4108 (N_4108,N_3794,N_3662);
nor U4109 (N_4109,N_3568,N_3579);
nand U4110 (N_4110,N_3804,N_3722);
and U4111 (N_4111,N_3634,N_3921);
or U4112 (N_4112,N_3733,N_3955);
nand U4113 (N_4113,N_3828,N_3827);
nand U4114 (N_4114,N_3876,N_3532);
nor U4115 (N_4115,N_3581,N_3971);
or U4116 (N_4116,N_3723,N_3983);
or U4117 (N_4117,N_3748,N_3549);
nand U4118 (N_4118,N_3728,N_3970);
or U4119 (N_4119,N_3610,N_3726);
or U4120 (N_4120,N_3590,N_3653);
or U4121 (N_4121,N_3691,N_3883);
nand U4122 (N_4122,N_3908,N_3712);
and U4123 (N_4123,N_3865,N_3607);
and U4124 (N_4124,N_3837,N_3686);
nor U4125 (N_4125,N_3945,N_3541);
nor U4126 (N_4126,N_3985,N_3781);
nand U4127 (N_4127,N_3626,N_3878);
and U4128 (N_4128,N_3700,N_3916);
xnor U4129 (N_4129,N_3834,N_3757);
and U4130 (N_4130,N_3520,N_3799);
nand U4131 (N_4131,N_3561,N_3974);
and U4132 (N_4132,N_3719,N_3933);
and U4133 (N_4133,N_3756,N_3785);
xor U4134 (N_4134,N_3839,N_3655);
and U4135 (N_4135,N_3642,N_3524);
nor U4136 (N_4136,N_3845,N_3759);
or U4137 (N_4137,N_3737,N_3752);
xnor U4138 (N_4138,N_3538,N_3525);
xnor U4139 (N_4139,N_3967,N_3684);
nor U4140 (N_4140,N_3932,N_3861);
and U4141 (N_4141,N_3641,N_3791);
or U4142 (N_4142,N_3560,N_3515);
or U4143 (N_4143,N_3925,N_3574);
nor U4144 (N_4144,N_3586,N_3656);
and U4145 (N_4145,N_3621,N_3565);
nand U4146 (N_4146,N_3856,N_3897);
nand U4147 (N_4147,N_3841,N_3903);
nor U4148 (N_4148,N_3783,N_3769);
and U4149 (N_4149,N_3923,N_3598);
nor U4150 (N_4150,N_3917,N_3747);
and U4151 (N_4151,N_3569,N_3847);
nor U4152 (N_4152,N_3957,N_3692);
or U4153 (N_4153,N_3514,N_3906);
or U4154 (N_4154,N_3889,N_3556);
and U4155 (N_4155,N_3849,N_3886);
and U4156 (N_4156,N_3953,N_3798);
or U4157 (N_4157,N_3928,N_3599);
or U4158 (N_4158,N_3840,N_3893);
xnor U4159 (N_4159,N_3802,N_3870);
nor U4160 (N_4160,N_3761,N_3539);
and U4161 (N_4161,N_3760,N_3825);
nor U4162 (N_4162,N_3724,N_3749);
nand U4163 (N_4163,N_3978,N_3850);
nor U4164 (N_4164,N_3672,N_3986);
nor U4165 (N_4165,N_3715,N_3881);
and U4166 (N_4166,N_3558,N_3972);
xor U4167 (N_4167,N_3547,N_3947);
xnor U4168 (N_4168,N_3899,N_3682);
nand U4169 (N_4169,N_3976,N_3994);
nor U4170 (N_4170,N_3689,N_3633);
and U4171 (N_4171,N_3546,N_3987);
xnor U4172 (N_4172,N_3969,N_3531);
and U4173 (N_4173,N_3585,N_3910);
nor U4174 (N_4174,N_3892,N_3548);
nand U4175 (N_4175,N_3973,N_3773);
nor U4176 (N_4176,N_3604,N_3992);
xnor U4177 (N_4177,N_3809,N_3711);
nor U4178 (N_4178,N_3725,N_3868);
nand U4179 (N_4179,N_3912,N_3784);
nor U4180 (N_4180,N_3508,N_3746);
nand U4181 (N_4181,N_3941,N_3666);
nand U4182 (N_4182,N_3929,N_3951);
xnor U4183 (N_4183,N_3846,N_3555);
xor U4184 (N_4184,N_3862,N_3716);
xor U4185 (N_4185,N_3742,N_3727);
xor U4186 (N_4186,N_3900,N_3668);
nand U4187 (N_4187,N_3778,N_3540);
nand U4188 (N_4188,N_3611,N_3872);
or U4189 (N_4189,N_3990,N_3772);
nand U4190 (N_4190,N_3943,N_3884);
xor U4191 (N_4191,N_3631,N_3665);
or U4192 (N_4192,N_3605,N_3807);
nor U4193 (N_4193,N_3770,N_3805);
nand U4194 (N_4194,N_3998,N_3506);
or U4195 (N_4195,N_3573,N_3767);
or U4196 (N_4196,N_3564,N_3988);
xor U4197 (N_4197,N_3762,N_3829);
nor U4198 (N_4198,N_3814,N_3664);
and U4199 (N_4199,N_3858,N_3909);
nand U4200 (N_4200,N_3882,N_3871);
nor U4201 (N_4201,N_3718,N_3877);
and U4202 (N_4202,N_3601,N_3553);
nor U4203 (N_4203,N_3661,N_3649);
or U4204 (N_4204,N_3832,N_3946);
nand U4205 (N_4205,N_3950,N_3528);
nand U4206 (N_4206,N_3758,N_3864);
nand U4207 (N_4207,N_3755,N_3963);
nand U4208 (N_4208,N_3813,N_3907);
and U4209 (N_4209,N_3962,N_3636);
and U4210 (N_4210,N_3942,N_3620);
nand U4211 (N_4211,N_3647,N_3504);
xor U4212 (N_4212,N_3575,N_3958);
or U4213 (N_4213,N_3913,N_3936);
nor U4214 (N_4214,N_3999,N_3640);
nor U4215 (N_4215,N_3509,N_3594);
and U4216 (N_4216,N_3800,N_3960);
and U4217 (N_4217,N_3519,N_3518);
or U4218 (N_4218,N_3687,N_3853);
nor U4219 (N_4219,N_3842,N_3694);
nor U4220 (N_4220,N_3616,N_3830);
nor U4221 (N_4221,N_3792,N_3754);
nand U4222 (N_4222,N_3527,N_3697);
xor U4223 (N_4223,N_3857,N_3833);
nand U4224 (N_4224,N_3638,N_3693);
or U4225 (N_4225,N_3577,N_3678);
xor U4226 (N_4226,N_3948,N_3979);
or U4227 (N_4227,N_3823,N_3696);
nor U4228 (N_4228,N_3703,N_3993);
nor U4229 (N_4229,N_3873,N_3977);
nor U4230 (N_4230,N_3806,N_3795);
or U4231 (N_4231,N_3648,N_3965);
and U4232 (N_4232,N_3934,N_3651);
and U4233 (N_4233,N_3630,N_3632);
nand U4234 (N_4234,N_3677,N_3959);
or U4235 (N_4235,N_3530,N_3991);
nor U4236 (N_4236,N_3854,N_3552);
xor U4237 (N_4237,N_3803,N_3919);
xnor U4238 (N_4238,N_3592,N_3695);
and U4239 (N_4239,N_3989,N_3690);
or U4240 (N_4240,N_3776,N_3730);
xor U4241 (N_4241,N_3644,N_3589);
nand U4242 (N_4242,N_3818,N_3535);
xor U4243 (N_4243,N_3875,N_3628);
nor U4244 (N_4244,N_3510,N_3654);
nand U4245 (N_4245,N_3744,N_3673);
nand U4246 (N_4246,N_3855,N_3667);
xor U4247 (N_4247,N_3734,N_3981);
or U4248 (N_4248,N_3874,N_3602);
xnor U4249 (N_4249,N_3924,N_3914);
nand U4250 (N_4250,N_3631,N_3938);
xnor U4251 (N_4251,N_3766,N_3532);
xor U4252 (N_4252,N_3757,N_3793);
xnor U4253 (N_4253,N_3617,N_3954);
and U4254 (N_4254,N_3694,N_3677);
and U4255 (N_4255,N_3992,N_3618);
and U4256 (N_4256,N_3864,N_3935);
or U4257 (N_4257,N_3685,N_3890);
nor U4258 (N_4258,N_3624,N_3909);
and U4259 (N_4259,N_3764,N_3970);
nand U4260 (N_4260,N_3657,N_3888);
xor U4261 (N_4261,N_3878,N_3823);
nand U4262 (N_4262,N_3768,N_3630);
nand U4263 (N_4263,N_3935,N_3659);
and U4264 (N_4264,N_3719,N_3763);
nor U4265 (N_4265,N_3587,N_3947);
or U4266 (N_4266,N_3768,N_3939);
or U4267 (N_4267,N_3741,N_3684);
xor U4268 (N_4268,N_3713,N_3794);
xor U4269 (N_4269,N_3726,N_3877);
or U4270 (N_4270,N_3727,N_3757);
or U4271 (N_4271,N_3730,N_3592);
or U4272 (N_4272,N_3818,N_3622);
and U4273 (N_4273,N_3874,N_3802);
nor U4274 (N_4274,N_3886,N_3836);
nor U4275 (N_4275,N_3964,N_3833);
xor U4276 (N_4276,N_3878,N_3761);
xnor U4277 (N_4277,N_3925,N_3899);
nand U4278 (N_4278,N_3813,N_3837);
or U4279 (N_4279,N_3883,N_3705);
xor U4280 (N_4280,N_3711,N_3593);
or U4281 (N_4281,N_3527,N_3942);
nor U4282 (N_4282,N_3515,N_3704);
nand U4283 (N_4283,N_3682,N_3530);
nor U4284 (N_4284,N_3585,N_3713);
xor U4285 (N_4285,N_3587,N_3718);
and U4286 (N_4286,N_3690,N_3764);
and U4287 (N_4287,N_3970,N_3601);
and U4288 (N_4288,N_3874,N_3512);
nand U4289 (N_4289,N_3588,N_3764);
nand U4290 (N_4290,N_3862,N_3712);
xnor U4291 (N_4291,N_3940,N_3511);
xnor U4292 (N_4292,N_3768,N_3716);
or U4293 (N_4293,N_3726,N_3901);
and U4294 (N_4294,N_3976,N_3947);
nand U4295 (N_4295,N_3510,N_3699);
nor U4296 (N_4296,N_3854,N_3757);
nand U4297 (N_4297,N_3850,N_3501);
nor U4298 (N_4298,N_3517,N_3753);
or U4299 (N_4299,N_3567,N_3775);
or U4300 (N_4300,N_3631,N_3728);
and U4301 (N_4301,N_3799,N_3677);
nand U4302 (N_4302,N_3510,N_3842);
nor U4303 (N_4303,N_3702,N_3665);
or U4304 (N_4304,N_3724,N_3828);
or U4305 (N_4305,N_3882,N_3543);
nor U4306 (N_4306,N_3560,N_3926);
xor U4307 (N_4307,N_3982,N_3757);
nor U4308 (N_4308,N_3607,N_3890);
nor U4309 (N_4309,N_3770,N_3860);
nor U4310 (N_4310,N_3557,N_3982);
nand U4311 (N_4311,N_3752,N_3782);
and U4312 (N_4312,N_3525,N_3664);
nand U4313 (N_4313,N_3692,N_3652);
and U4314 (N_4314,N_3709,N_3522);
nand U4315 (N_4315,N_3543,N_3790);
nor U4316 (N_4316,N_3706,N_3658);
nor U4317 (N_4317,N_3915,N_3948);
and U4318 (N_4318,N_3684,N_3998);
nand U4319 (N_4319,N_3692,N_3996);
or U4320 (N_4320,N_3890,N_3846);
nand U4321 (N_4321,N_3668,N_3627);
xnor U4322 (N_4322,N_3515,N_3867);
or U4323 (N_4323,N_3624,N_3972);
nand U4324 (N_4324,N_3903,N_3876);
xnor U4325 (N_4325,N_3800,N_3955);
nor U4326 (N_4326,N_3969,N_3919);
nand U4327 (N_4327,N_3950,N_3731);
or U4328 (N_4328,N_3743,N_3899);
nor U4329 (N_4329,N_3889,N_3649);
xnor U4330 (N_4330,N_3517,N_3577);
nand U4331 (N_4331,N_3732,N_3681);
or U4332 (N_4332,N_3919,N_3516);
xor U4333 (N_4333,N_3768,N_3901);
nand U4334 (N_4334,N_3573,N_3597);
or U4335 (N_4335,N_3819,N_3944);
and U4336 (N_4336,N_3880,N_3749);
xor U4337 (N_4337,N_3598,N_3786);
or U4338 (N_4338,N_3820,N_3855);
xnor U4339 (N_4339,N_3603,N_3878);
nor U4340 (N_4340,N_3892,N_3825);
nand U4341 (N_4341,N_3645,N_3590);
and U4342 (N_4342,N_3549,N_3615);
nor U4343 (N_4343,N_3806,N_3808);
and U4344 (N_4344,N_3671,N_3628);
xnor U4345 (N_4345,N_3694,N_3953);
nand U4346 (N_4346,N_3715,N_3861);
or U4347 (N_4347,N_3795,N_3615);
nor U4348 (N_4348,N_3682,N_3933);
nand U4349 (N_4349,N_3517,N_3899);
or U4350 (N_4350,N_3840,N_3515);
or U4351 (N_4351,N_3835,N_3756);
nand U4352 (N_4352,N_3809,N_3878);
xor U4353 (N_4353,N_3531,N_3751);
or U4354 (N_4354,N_3617,N_3594);
nand U4355 (N_4355,N_3640,N_3704);
xnor U4356 (N_4356,N_3704,N_3663);
nand U4357 (N_4357,N_3983,N_3532);
and U4358 (N_4358,N_3636,N_3567);
and U4359 (N_4359,N_3928,N_3566);
nor U4360 (N_4360,N_3669,N_3969);
nand U4361 (N_4361,N_3621,N_3535);
or U4362 (N_4362,N_3961,N_3922);
and U4363 (N_4363,N_3918,N_3812);
or U4364 (N_4364,N_3547,N_3508);
nor U4365 (N_4365,N_3500,N_3749);
xnor U4366 (N_4366,N_3685,N_3928);
or U4367 (N_4367,N_3919,N_3962);
nor U4368 (N_4368,N_3983,N_3653);
or U4369 (N_4369,N_3619,N_3860);
xnor U4370 (N_4370,N_3909,N_3835);
nand U4371 (N_4371,N_3819,N_3606);
nor U4372 (N_4372,N_3740,N_3795);
xnor U4373 (N_4373,N_3575,N_3610);
and U4374 (N_4374,N_3645,N_3672);
nand U4375 (N_4375,N_3671,N_3771);
and U4376 (N_4376,N_3567,N_3905);
xor U4377 (N_4377,N_3958,N_3525);
nor U4378 (N_4378,N_3599,N_3525);
xor U4379 (N_4379,N_3713,N_3631);
nor U4380 (N_4380,N_3847,N_3893);
or U4381 (N_4381,N_3614,N_3646);
nor U4382 (N_4382,N_3894,N_3912);
and U4383 (N_4383,N_3513,N_3883);
xor U4384 (N_4384,N_3666,N_3797);
nor U4385 (N_4385,N_3981,N_3928);
xnor U4386 (N_4386,N_3879,N_3747);
nor U4387 (N_4387,N_3607,N_3731);
nor U4388 (N_4388,N_3769,N_3964);
or U4389 (N_4389,N_3614,N_3652);
nand U4390 (N_4390,N_3552,N_3833);
and U4391 (N_4391,N_3607,N_3606);
and U4392 (N_4392,N_3986,N_3564);
or U4393 (N_4393,N_3834,N_3573);
nor U4394 (N_4394,N_3945,N_3907);
or U4395 (N_4395,N_3629,N_3944);
or U4396 (N_4396,N_3797,N_3814);
xor U4397 (N_4397,N_3948,N_3644);
nand U4398 (N_4398,N_3809,N_3949);
or U4399 (N_4399,N_3825,N_3955);
and U4400 (N_4400,N_3707,N_3943);
and U4401 (N_4401,N_3681,N_3787);
or U4402 (N_4402,N_3937,N_3957);
and U4403 (N_4403,N_3535,N_3852);
nor U4404 (N_4404,N_3634,N_3983);
and U4405 (N_4405,N_3790,N_3797);
nand U4406 (N_4406,N_3541,N_3801);
nor U4407 (N_4407,N_3944,N_3616);
nand U4408 (N_4408,N_3925,N_3623);
nand U4409 (N_4409,N_3853,N_3820);
nor U4410 (N_4410,N_3584,N_3878);
nor U4411 (N_4411,N_3592,N_3948);
xor U4412 (N_4412,N_3592,N_3781);
nand U4413 (N_4413,N_3692,N_3628);
or U4414 (N_4414,N_3646,N_3877);
and U4415 (N_4415,N_3659,N_3934);
nor U4416 (N_4416,N_3507,N_3745);
nand U4417 (N_4417,N_3669,N_3632);
or U4418 (N_4418,N_3972,N_3676);
nand U4419 (N_4419,N_3515,N_3832);
nor U4420 (N_4420,N_3703,N_3867);
and U4421 (N_4421,N_3635,N_3724);
and U4422 (N_4422,N_3967,N_3837);
nor U4423 (N_4423,N_3651,N_3770);
nor U4424 (N_4424,N_3678,N_3928);
nor U4425 (N_4425,N_3933,N_3884);
and U4426 (N_4426,N_3671,N_3641);
nor U4427 (N_4427,N_3875,N_3584);
and U4428 (N_4428,N_3770,N_3837);
nor U4429 (N_4429,N_3689,N_3814);
and U4430 (N_4430,N_3806,N_3648);
and U4431 (N_4431,N_3996,N_3691);
nand U4432 (N_4432,N_3993,N_3628);
and U4433 (N_4433,N_3703,N_3504);
nand U4434 (N_4434,N_3563,N_3632);
nand U4435 (N_4435,N_3995,N_3700);
nor U4436 (N_4436,N_3695,N_3713);
or U4437 (N_4437,N_3653,N_3585);
xnor U4438 (N_4438,N_3602,N_3806);
nor U4439 (N_4439,N_3669,N_3519);
xor U4440 (N_4440,N_3729,N_3920);
nor U4441 (N_4441,N_3642,N_3795);
or U4442 (N_4442,N_3942,N_3661);
nor U4443 (N_4443,N_3811,N_3765);
xnor U4444 (N_4444,N_3737,N_3869);
or U4445 (N_4445,N_3581,N_3587);
nand U4446 (N_4446,N_3825,N_3896);
and U4447 (N_4447,N_3933,N_3703);
nand U4448 (N_4448,N_3523,N_3625);
and U4449 (N_4449,N_3969,N_3536);
and U4450 (N_4450,N_3830,N_3608);
nand U4451 (N_4451,N_3998,N_3502);
or U4452 (N_4452,N_3577,N_3905);
or U4453 (N_4453,N_3842,N_3620);
nand U4454 (N_4454,N_3938,N_3825);
and U4455 (N_4455,N_3785,N_3697);
nor U4456 (N_4456,N_3950,N_3953);
nor U4457 (N_4457,N_3952,N_3811);
nor U4458 (N_4458,N_3612,N_3999);
nor U4459 (N_4459,N_3986,N_3782);
xnor U4460 (N_4460,N_3520,N_3871);
nor U4461 (N_4461,N_3961,N_3968);
and U4462 (N_4462,N_3880,N_3938);
nand U4463 (N_4463,N_3900,N_3762);
and U4464 (N_4464,N_3801,N_3917);
nand U4465 (N_4465,N_3919,N_3963);
or U4466 (N_4466,N_3786,N_3766);
nand U4467 (N_4467,N_3982,N_3603);
nand U4468 (N_4468,N_3680,N_3780);
nor U4469 (N_4469,N_3511,N_3923);
xnor U4470 (N_4470,N_3911,N_3764);
or U4471 (N_4471,N_3756,N_3670);
and U4472 (N_4472,N_3572,N_3892);
xnor U4473 (N_4473,N_3558,N_3928);
or U4474 (N_4474,N_3916,N_3719);
nor U4475 (N_4475,N_3792,N_3590);
or U4476 (N_4476,N_3693,N_3685);
nand U4477 (N_4477,N_3517,N_3530);
or U4478 (N_4478,N_3601,N_3786);
nor U4479 (N_4479,N_3683,N_3967);
or U4480 (N_4480,N_3578,N_3925);
xnor U4481 (N_4481,N_3511,N_3919);
and U4482 (N_4482,N_3995,N_3762);
xor U4483 (N_4483,N_3722,N_3651);
or U4484 (N_4484,N_3558,N_3645);
or U4485 (N_4485,N_3860,N_3928);
xnor U4486 (N_4486,N_3593,N_3911);
nor U4487 (N_4487,N_3559,N_3934);
nor U4488 (N_4488,N_3875,N_3501);
nand U4489 (N_4489,N_3885,N_3962);
or U4490 (N_4490,N_3599,N_3837);
and U4491 (N_4491,N_3683,N_3911);
and U4492 (N_4492,N_3639,N_3829);
nand U4493 (N_4493,N_3844,N_3933);
xor U4494 (N_4494,N_3914,N_3669);
nand U4495 (N_4495,N_3665,N_3874);
nor U4496 (N_4496,N_3753,N_3858);
or U4497 (N_4497,N_3681,N_3776);
xnor U4498 (N_4498,N_3618,N_3647);
nand U4499 (N_4499,N_3889,N_3957);
nor U4500 (N_4500,N_4312,N_4295);
xnor U4501 (N_4501,N_4409,N_4346);
nand U4502 (N_4502,N_4469,N_4484);
and U4503 (N_4503,N_4284,N_4476);
nand U4504 (N_4504,N_4459,N_4177);
nand U4505 (N_4505,N_4376,N_4398);
xnor U4506 (N_4506,N_4230,N_4478);
nand U4507 (N_4507,N_4142,N_4375);
nor U4508 (N_4508,N_4193,N_4122);
and U4509 (N_4509,N_4178,N_4045);
or U4510 (N_4510,N_4013,N_4436);
or U4511 (N_4511,N_4348,N_4446);
and U4512 (N_4512,N_4341,N_4447);
nor U4513 (N_4513,N_4118,N_4331);
nand U4514 (N_4514,N_4078,N_4004);
nor U4515 (N_4515,N_4379,N_4318);
nor U4516 (N_4516,N_4048,N_4019);
and U4517 (N_4517,N_4251,N_4268);
nand U4518 (N_4518,N_4070,N_4360);
xnor U4519 (N_4519,N_4305,N_4008);
nand U4520 (N_4520,N_4261,N_4067);
xnor U4521 (N_4521,N_4220,N_4498);
xor U4522 (N_4522,N_4417,N_4362);
nor U4523 (N_4523,N_4432,N_4011);
or U4524 (N_4524,N_4363,N_4244);
nor U4525 (N_4525,N_4014,N_4236);
and U4526 (N_4526,N_4077,N_4279);
or U4527 (N_4527,N_4396,N_4024);
or U4528 (N_4528,N_4160,N_4413);
or U4529 (N_4529,N_4247,N_4200);
nor U4530 (N_4530,N_4347,N_4442);
and U4531 (N_4531,N_4337,N_4336);
xnor U4532 (N_4532,N_4427,N_4387);
nand U4533 (N_4533,N_4315,N_4212);
nor U4534 (N_4534,N_4222,N_4445);
nor U4535 (N_4535,N_4324,N_4232);
and U4536 (N_4536,N_4405,N_4136);
xnor U4537 (N_4537,N_4113,N_4357);
xor U4538 (N_4538,N_4304,N_4040);
and U4539 (N_4539,N_4176,N_4235);
nand U4540 (N_4540,N_4429,N_4463);
nand U4541 (N_4541,N_4258,N_4089);
xnor U4542 (N_4542,N_4069,N_4397);
nand U4543 (N_4543,N_4455,N_4172);
nor U4544 (N_4544,N_4390,N_4195);
or U4545 (N_4545,N_4156,N_4086);
nand U4546 (N_4546,N_4219,N_4111);
xnor U4547 (N_4547,N_4050,N_4152);
and U4548 (N_4548,N_4350,N_4022);
nor U4549 (N_4549,N_4472,N_4248);
and U4550 (N_4550,N_4146,N_4483);
nor U4551 (N_4551,N_4344,N_4450);
or U4552 (N_4552,N_4494,N_4128);
and U4553 (N_4553,N_4148,N_4240);
or U4554 (N_4554,N_4028,N_4425);
nor U4555 (N_4555,N_4031,N_4290);
nor U4556 (N_4556,N_4353,N_4002);
and U4557 (N_4557,N_4161,N_4313);
nor U4558 (N_4558,N_4433,N_4402);
nor U4559 (N_4559,N_4093,N_4190);
xnor U4560 (N_4560,N_4253,N_4407);
and U4561 (N_4561,N_4391,N_4280);
xor U4562 (N_4562,N_4266,N_4215);
nand U4563 (N_4563,N_4189,N_4238);
nand U4564 (N_4564,N_4403,N_4415);
and U4565 (N_4565,N_4294,N_4202);
and U4566 (N_4566,N_4068,N_4198);
nand U4567 (N_4567,N_4199,N_4488);
and U4568 (N_4568,N_4486,N_4466);
and U4569 (N_4569,N_4435,N_4036);
nand U4570 (N_4570,N_4191,N_4372);
xor U4571 (N_4571,N_4026,N_4299);
xor U4572 (N_4572,N_4201,N_4231);
or U4573 (N_4573,N_4159,N_4053);
and U4574 (N_4574,N_4091,N_4493);
nor U4575 (N_4575,N_4110,N_4441);
and U4576 (N_4576,N_4083,N_4175);
nand U4577 (N_4577,N_4210,N_4216);
or U4578 (N_4578,N_4132,N_4151);
nand U4579 (N_4579,N_4420,N_4034);
or U4580 (N_4580,N_4119,N_4325);
xor U4581 (N_4581,N_4271,N_4241);
nand U4582 (N_4582,N_4303,N_4073);
nor U4583 (N_4583,N_4009,N_4096);
xnor U4584 (N_4584,N_4367,N_4006);
or U4585 (N_4585,N_4120,N_4129);
or U4586 (N_4586,N_4381,N_4452);
nor U4587 (N_4587,N_4492,N_4204);
xnor U4588 (N_4588,N_4007,N_4197);
xnor U4589 (N_4589,N_4016,N_4426);
and U4590 (N_4590,N_4187,N_4449);
and U4591 (N_4591,N_4474,N_4252);
xor U4592 (N_4592,N_4227,N_4479);
nand U4593 (N_4593,N_4264,N_4029);
nor U4594 (N_4594,N_4371,N_4419);
or U4595 (N_4595,N_4229,N_4207);
and U4596 (N_4596,N_4010,N_4317);
or U4597 (N_4597,N_4226,N_4267);
nor U4598 (N_4598,N_4327,N_4233);
nand U4599 (N_4599,N_4246,N_4000);
nand U4600 (N_4600,N_4168,N_4465);
nand U4601 (N_4601,N_4460,N_4395);
nand U4602 (N_4602,N_4326,N_4174);
nand U4603 (N_4603,N_4170,N_4150);
or U4604 (N_4604,N_4351,N_4464);
or U4605 (N_4605,N_4046,N_4328);
and U4606 (N_4606,N_4075,N_4308);
and U4607 (N_4607,N_4361,N_4355);
or U4608 (N_4608,N_4203,N_4301);
or U4609 (N_4609,N_4329,N_4408);
and U4610 (N_4610,N_4289,N_4237);
xnor U4611 (N_4611,N_4477,N_4393);
or U4612 (N_4612,N_4074,N_4404);
nand U4613 (N_4613,N_4349,N_4414);
or U4614 (N_4614,N_4462,N_4056);
xor U4615 (N_4615,N_4491,N_4342);
or U4616 (N_4616,N_4225,N_4154);
and U4617 (N_4617,N_4054,N_4380);
nor U4618 (N_4618,N_4256,N_4275);
nor U4619 (N_4619,N_4082,N_4033);
and U4620 (N_4620,N_4439,N_4133);
and U4621 (N_4621,N_4223,N_4311);
xnor U4622 (N_4622,N_4260,N_4287);
and U4623 (N_4623,N_4292,N_4386);
xor U4624 (N_4624,N_4468,N_4181);
or U4625 (N_4625,N_4106,N_4412);
and U4626 (N_4626,N_4416,N_4027);
and U4627 (N_4627,N_4400,N_4140);
xor U4628 (N_4628,N_4265,N_4081);
or U4629 (N_4629,N_4080,N_4126);
nand U4630 (N_4630,N_4316,N_4323);
and U4631 (N_4631,N_4319,N_4164);
nor U4632 (N_4632,N_4457,N_4208);
and U4633 (N_4633,N_4281,N_4064);
nand U4634 (N_4634,N_4188,N_4012);
and U4635 (N_4635,N_4072,N_4257);
and U4636 (N_4636,N_4343,N_4103);
or U4637 (N_4637,N_4333,N_4017);
and U4638 (N_4638,N_4021,N_4043);
or U4639 (N_4639,N_4388,N_4141);
nand U4640 (N_4640,N_4489,N_4114);
and U4641 (N_4641,N_4144,N_4421);
or U4642 (N_4642,N_4431,N_4286);
nand U4643 (N_4643,N_4157,N_4377);
nand U4644 (N_4644,N_4123,N_4352);
and U4645 (N_4645,N_4035,N_4480);
xor U4646 (N_4646,N_4125,N_4307);
or U4647 (N_4647,N_4003,N_4038);
nor U4648 (N_4648,N_4098,N_4254);
nand U4649 (N_4649,N_4471,N_4167);
or U4650 (N_4650,N_4205,N_4411);
or U4651 (N_4651,N_4255,N_4100);
nor U4652 (N_4652,N_4166,N_4213);
nand U4653 (N_4653,N_4183,N_4061);
or U4654 (N_4654,N_4139,N_4039);
nor U4655 (N_4655,N_4276,N_4099);
nor U4656 (N_4656,N_4134,N_4209);
and U4657 (N_4657,N_4242,N_4196);
or U4658 (N_4658,N_4456,N_4298);
nand U4659 (N_4659,N_4116,N_4076);
or U4660 (N_4660,N_4025,N_4030);
xor U4661 (N_4661,N_4153,N_4273);
or U4662 (N_4662,N_4454,N_4218);
nand U4663 (N_4663,N_4293,N_4461);
nand U4664 (N_4664,N_4041,N_4145);
xnor U4665 (N_4665,N_4079,N_4368);
and U4666 (N_4666,N_4481,N_4018);
and U4667 (N_4667,N_4165,N_4105);
and U4668 (N_4668,N_4163,N_4487);
nand U4669 (N_4669,N_4023,N_4135);
xor U4670 (N_4670,N_4071,N_4345);
and U4671 (N_4671,N_4044,N_4097);
nor U4672 (N_4672,N_4259,N_4364);
and U4673 (N_4673,N_4149,N_4370);
xor U4674 (N_4674,N_4084,N_4066);
nand U4675 (N_4675,N_4042,N_4310);
nor U4676 (N_4676,N_4121,N_4117);
or U4677 (N_4677,N_4032,N_4055);
or U4678 (N_4678,N_4047,N_4297);
nor U4679 (N_4679,N_4049,N_4262);
or U4680 (N_4680,N_4389,N_4302);
or U4681 (N_4681,N_4060,N_4101);
or U4682 (N_4682,N_4224,N_4422);
xor U4683 (N_4683,N_4185,N_4162);
xor U4684 (N_4684,N_4094,N_4438);
or U4685 (N_4685,N_4158,N_4057);
xnor U4686 (N_4686,N_4130,N_4321);
xnor U4687 (N_4687,N_4037,N_4496);
nor U4688 (N_4688,N_4102,N_4340);
nor U4689 (N_4689,N_4320,N_4155);
or U4690 (N_4690,N_4374,N_4495);
and U4691 (N_4691,N_4108,N_4051);
xnor U4692 (N_4692,N_4288,N_4090);
xor U4693 (N_4693,N_4499,N_4282);
and U4694 (N_4694,N_4369,N_4383);
xnor U4695 (N_4695,N_4410,N_4087);
or U4696 (N_4696,N_4485,N_4270);
nand U4697 (N_4697,N_4206,N_4497);
nor U4698 (N_4698,N_4444,N_4467);
and U4699 (N_4699,N_4385,N_4274);
nand U4700 (N_4700,N_4243,N_4092);
nor U4701 (N_4701,N_4291,N_4314);
and U4702 (N_4702,N_4179,N_4285);
nor U4703 (N_4703,N_4239,N_4428);
nand U4704 (N_4704,N_4180,N_4338);
and U4705 (N_4705,N_4424,N_4131);
nand U4706 (N_4706,N_4115,N_4058);
xnor U4707 (N_4707,N_4490,N_4354);
nor U4708 (N_4708,N_4334,N_4448);
xor U4709 (N_4709,N_4194,N_4399);
xor U4710 (N_4710,N_4112,N_4147);
nor U4711 (N_4711,N_4137,N_4211);
nand U4712 (N_4712,N_4382,N_4062);
or U4713 (N_4713,N_4365,N_4430);
xnor U4714 (N_4714,N_4423,N_4283);
and U4715 (N_4715,N_4182,N_4339);
nor U4716 (N_4716,N_4228,N_4214);
nand U4717 (N_4717,N_4221,N_4020);
nand U4718 (N_4718,N_4245,N_4309);
nand U4719 (N_4719,N_4406,N_4109);
xor U4720 (N_4720,N_4127,N_4453);
and U4721 (N_4721,N_4278,N_4104);
or U4722 (N_4722,N_4088,N_4359);
or U4723 (N_4723,N_4107,N_4475);
nand U4724 (N_4724,N_4143,N_4473);
nand U4725 (N_4725,N_4272,N_4217);
nor U4726 (N_4726,N_4063,N_4234);
nor U4727 (N_4727,N_4138,N_4330);
or U4728 (N_4728,N_4184,N_4059);
nor U4729 (N_4729,N_4296,N_4171);
xor U4730 (N_4730,N_4249,N_4384);
and U4731 (N_4731,N_4001,N_4394);
and U4732 (N_4732,N_4269,N_4332);
or U4733 (N_4733,N_4458,N_4401);
xor U4734 (N_4734,N_4482,N_4443);
or U4735 (N_4735,N_4356,N_4015);
nand U4736 (N_4736,N_4366,N_4005);
nand U4737 (N_4737,N_4306,N_4470);
or U4738 (N_4738,N_4263,N_4437);
nand U4739 (N_4739,N_4322,N_4250);
nor U4740 (N_4740,N_4124,N_4358);
xnor U4741 (N_4741,N_4173,N_4300);
nor U4742 (N_4742,N_4095,N_4451);
xor U4743 (N_4743,N_4378,N_4434);
nor U4744 (N_4744,N_4373,N_4065);
nand U4745 (N_4745,N_4169,N_4186);
nor U4746 (N_4746,N_4440,N_4052);
and U4747 (N_4747,N_4085,N_4335);
xor U4748 (N_4748,N_4277,N_4418);
or U4749 (N_4749,N_4192,N_4392);
and U4750 (N_4750,N_4158,N_4477);
and U4751 (N_4751,N_4247,N_4046);
xor U4752 (N_4752,N_4105,N_4460);
or U4753 (N_4753,N_4382,N_4360);
or U4754 (N_4754,N_4159,N_4221);
nor U4755 (N_4755,N_4191,N_4308);
xor U4756 (N_4756,N_4296,N_4334);
nand U4757 (N_4757,N_4348,N_4037);
nor U4758 (N_4758,N_4037,N_4207);
or U4759 (N_4759,N_4476,N_4486);
nand U4760 (N_4760,N_4347,N_4084);
nand U4761 (N_4761,N_4324,N_4071);
nand U4762 (N_4762,N_4185,N_4447);
or U4763 (N_4763,N_4060,N_4362);
nor U4764 (N_4764,N_4149,N_4309);
or U4765 (N_4765,N_4352,N_4300);
nand U4766 (N_4766,N_4424,N_4177);
nor U4767 (N_4767,N_4117,N_4142);
nand U4768 (N_4768,N_4335,N_4469);
nand U4769 (N_4769,N_4305,N_4223);
and U4770 (N_4770,N_4384,N_4324);
xnor U4771 (N_4771,N_4052,N_4011);
nand U4772 (N_4772,N_4082,N_4488);
nand U4773 (N_4773,N_4497,N_4231);
nand U4774 (N_4774,N_4241,N_4048);
and U4775 (N_4775,N_4209,N_4446);
and U4776 (N_4776,N_4117,N_4429);
xor U4777 (N_4777,N_4093,N_4272);
nor U4778 (N_4778,N_4484,N_4150);
nor U4779 (N_4779,N_4074,N_4345);
or U4780 (N_4780,N_4235,N_4310);
and U4781 (N_4781,N_4117,N_4188);
or U4782 (N_4782,N_4364,N_4200);
xnor U4783 (N_4783,N_4280,N_4138);
nor U4784 (N_4784,N_4253,N_4060);
xor U4785 (N_4785,N_4048,N_4101);
nand U4786 (N_4786,N_4376,N_4067);
and U4787 (N_4787,N_4054,N_4216);
and U4788 (N_4788,N_4480,N_4438);
nand U4789 (N_4789,N_4224,N_4119);
nand U4790 (N_4790,N_4298,N_4459);
nand U4791 (N_4791,N_4446,N_4444);
nor U4792 (N_4792,N_4217,N_4278);
xnor U4793 (N_4793,N_4458,N_4141);
nand U4794 (N_4794,N_4435,N_4423);
nor U4795 (N_4795,N_4360,N_4421);
nor U4796 (N_4796,N_4269,N_4154);
and U4797 (N_4797,N_4104,N_4488);
and U4798 (N_4798,N_4295,N_4317);
or U4799 (N_4799,N_4497,N_4089);
nor U4800 (N_4800,N_4383,N_4128);
and U4801 (N_4801,N_4045,N_4305);
xor U4802 (N_4802,N_4419,N_4230);
or U4803 (N_4803,N_4357,N_4056);
and U4804 (N_4804,N_4199,N_4406);
nor U4805 (N_4805,N_4205,N_4181);
nor U4806 (N_4806,N_4001,N_4434);
or U4807 (N_4807,N_4059,N_4020);
or U4808 (N_4808,N_4344,N_4015);
nor U4809 (N_4809,N_4135,N_4100);
and U4810 (N_4810,N_4349,N_4377);
nand U4811 (N_4811,N_4150,N_4324);
nor U4812 (N_4812,N_4235,N_4260);
xor U4813 (N_4813,N_4277,N_4424);
xor U4814 (N_4814,N_4267,N_4102);
and U4815 (N_4815,N_4057,N_4202);
nor U4816 (N_4816,N_4293,N_4363);
nor U4817 (N_4817,N_4351,N_4247);
nor U4818 (N_4818,N_4292,N_4064);
nand U4819 (N_4819,N_4299,N_4497);
xor U4820 (N_4820,N_4345,N_4073);
nand U4821 (N_4821,N_4355,N_4412);
nand U4822 (N_4822,N_4255,N_4478);
or U4823 (N_4823,N_4432,N_4466);
xor U4824 (N_4824,N_4081,N_4171);
nor U4825 (N_4825,N_4070,N_4352);
nor U4826 (N_4826,N_4122,N_4052);
or U4827 (N_4827,N_4292,N_4141);
nor U4828 (N_4828,N_4114,N_4349);
and U4829 (N_4829,N_4406,N_4498);
or U4830 (N_4830,N_4224,N_4059);
and U4831 (N_4831,N_4370,N_4306);
xor U4832 (N_4832,N_4042,N_4374);
nand U4833 (N_4833,N_4277,N_4062);
or U4834 (N_4834,N_4068,N_4373);
xor U4835 (N_4835,N_4036,N_4241);
and U4836 (N_4836,N_4297,N_4197);
nor U4837 (N_4837,N_4085,N_4091);
nand U4838 (N_4838,N_4078,N_4060);
nor U4839 (N_4839,N_4483,N_4312);
and U4840 (N_4840,N_4292,N_4454);
and U4841 (N_4841,N_4249,N_4030);
nor U4842 (N_4842,N_4415,N_4481);
and U4843 (N_4843,N_4262,N_4401);
or U4844 (N_4844,N_4272,N_4241);
xor U4845 (N_4845,N_4144,N_4328);
and U4846 (N_4846,N_4085,N_4423);
nor U4847 (N_4847,N_4458,N_4327);
nand U4848 (N_4848,N_4436,N_4249);
nor U4849 (N_4849,N_4413,N_4415);
nand U4850 (N_4850,N_4101,N_4035);
or U4851 (N_4851,N_4013,N_4328);
or U4852 (N_4852,N_4405,N_4436);
or U4853 (N_4853,N_4197,N_4393);
or U4854 (N_4854,N_4048,N_4189);
or U4855 (N_4855,N_4302,N_4056);
or U4856 (N_4856,N_4217,N_4178);
nor U4857 (N_4857,N_4459,N_4251);
nand U4858 (N_4858,N_4483,N_4141);
nand U4859 (N_4859,N_4072,N_4058);
and U4860 (N_4860,N_4154,N_4460);
and U4861 (N_4861,N_4050,N_4071);
nor U4862 (N_4862,N_4123,N_4274);
and U4863 (N_4863,N_4108,N_4317);
nor U4864 (N_4864,N_4163,N_4028);
and U4865 (N_4865,N_4323,N_4132);
nor U4866 (N_4866,N_4153,N_4138);
nor U4867 (N_4867,N_4092,N_4239);
xor U4868 (N_4868,N_4201,N_4273);
xnor U4869 (N_4869,N_4378,N_4487);
nor U4870 (N_4870,N_4396,N_4201);
nor U4871 (N_4871,N_4281,N_4060);
nor U4872 (N_4872,N_4093,N_4253);
nor U4873 (N_4873,N_4197,N_4401);
and U4874 (N_4874,N_4402,N_4396);
xor U4875 (N_4875,N_4423,N_4060);
and U4876 (N_4876,N_4384,N_4464);
or U4877 (N_4877,N_4169,N_4389);
or U4878 (N_4878,N_4004,N_4235);
and U4879 (N_4879,N_4194,N_4011);
or U4880 (N_4880,N_4467,N_4165);
nand U4881 (N_4881,N_4045,N_4030);
and U4882 (N_4882,N_4371,N_4241);
xor U4883 (N_4883,N_4392,N_4329);
xnor U4884 (N_4884,N_4009,N_4375);
or U4885 (N_4885,N_4467,N_4447);
or U4886 (N_4886,N_4023,N_4017);
and U4887 (N_4887,N_4329,N_4117);
and U4888 (N_4888,N_4448,N_4114);
nor U4889 (N_4889,N_4238,N_4212);
or U4890 (N_4890,N_4132,N_4025);
nor U4891 (N_4891,N_4334,N_4493);
nor U4892 (N_4892,N_4120,N_4255);
nor U4893 (N_4893,N_4410,N_4221);
nand U4894 (N_4894,N_4011,N_4373);
nor U4895 (N_4895,N_4210,N_4234);
and U4896 (N_4896,N_4492,N_4168);
or U4897 (N_4897,N_4277,N_4251);
nor U4898 (N_4898,N_4140,N_4090);
xnor U4899 (N_4899,N_4021,N_4167);
nor U4900 (N_4900,N_4016,N_4131);
or U4901 (N_4901,N_4360,N_4425);
xnor U4902 (N_4902,N_4497,N_4283);
nor U4903 (N_4903,N_4365,N_4404);
xnor U4904 (N_4904,N_4441,N_4498);
nand U4905 (N_4905,N_4313,N_4483);
nor U4906 (N_4906,N_4476,N_4115);
nand U4907 (N_4907,N_4204,N_4300);
nor U4908 (N_4908,N_4428,N_4422);
nand U4909 (N_4909,N_4116,N_4113);
xnor U4910 (N_4910,N_4047,N_4214);
xor U4911 (N_4911,N_4423,N_4103);
or U4912 (N_4912,N_4071,N_4119);
and U4913 (N_4913,N_4391,N_4385);
xor U4914 (N_4914,N_4466,N_4401);
and U4915 (N_4915,N_4022,N_4258);
nand U4916 (N_4916,N_4205,N_4344);
and U4917 (N_4917,N_4172,N_4475);
nand U4918 (N_4918,N_4252,N_4256);
and U4919 (N_4919,N_4237,N_4172);
nand U4920 (N_4920,N_4448,N_4139);
xor U4921 (N_4921,N_4285,N_4379);
or U4922 (N_4922,N_4441,N_4160);
nor U4923 (N_4923,N_4298,N_4096);
nor U4924 (N_4924,N_4283,N_4417);
and U4925 (N_4925,N_4197,N_4363);
or U4926 (N_4926,N_4233,N_4250);
or U4927 (N_4927,N_4221,N_4179);
nor U4928 (N_4928,N_4199,N_4070);
or U4929 (N_4929,N_4446,N_4219);
xor U4930 (N_4930,N_4411,N_4405);
nand U4931 (N_4931,N_4023,N_4058);
nand U4932 (N_4932,N_4233,N_4293);
xnor U4933 (N_4933,N_4130,N_4350);
and U4934 (N_4934,N_4167,N_4362);
nand U4935 (N_4935,N_4334,N_4211);
nand U4936 (N_4936,N_4393,N_4487);
or U4937 (N_4937,N_4006,N_4275);
nand U4938 (N_4938,N_4075,N_4063);
or U4939 (N_4939,N_4310,N_4328);
nor U4940 (N_4940,N_4273,N_4200);
or U4941 (N_4941,N_4061,N_4329);
or U4942 (N_4942,N_4156,N_4376);
xnor U4943 (N_4943,N_4237,N_4296);
and U4944 (N_4944,N_4269,N_4085);
or U4945 (N_4945,N_4207,N_4070);
or U4946 (N_4946,N_4083,N_4350);
or U4947 (N_4947,N_4482,N_4263);
nor U4948 (N_4948,N_4329,N_4231);
xor U4949 (N_4949,N_4418,N_4347);
nand U4950 (N_4950,N_4223,N_4301);
xnor U4951 (N_4951,N_4182,N_4043);
nor U4952 (N_4952,N_4361,N_4449);
nand U4953 (N_4953,N_4183,N_4477);
nand U4954 (N_4954,N_4198,N_4410);
nand U4955 (N_4955,N_4455,N_4234);
nand U4956 (N_4956,N_4157,N_4432);
nor U4957 (N_4957,N_4205,N_4019);
nand U4958 (N_4958,N_4092,N_4101);
or U4959 (N_4959,N_4324,N_4459);
or U4960 (N_4960,N_4219,N_4306);
or U4961 (N_4961,N_4352,N_4433);
nor U4962 (N_4962,N_4133,N_4386);
nor U4963 (N_4963,N_4025,N_4448);
or U4964 (N_4964,N_4155,N_4199);
nor U4965 (N_4965,N_4287,N_4090);
nand U4966 (N_4966,N_4283,N_4274);
nor U4967 (N_4967,N_4248,N_4164);
xor U4968 (N_4968,N_4357,N_4475);
and U4969 (N_4969,N_4035,N_4087);
or U4970 (N_4970,N_4283,N_4335);
nor U4971 (N_4971,N_4418,N_4393);
or U4972 (N_4972,N_4089,N_4092);
nand U4973 (N_4973,N_4304,N_4136);
nand U4974 (N_4974,N_4407,N_4233);
xnor U4975 (N_4975,N_4460,N_4042);
and U4976 (N_4976,N_4365,N_4103);
nand U4977 (N_4977,N_4034,N_4213);
nand U4978 (N_4978,N_4162,N_4329);
and U4979 (N_4979,N_4199,N_4172);
or U4980 (N_4980,N_4364,N_4400);
or U4981 (N_4981,N_4486,N_4415);
nor U4982 (N_4982,N_4491,N_4071);
and U4983 (N_4983,N_4066,N_4202);
nand U4984 (N_4984,N_4331,N_4292);
nor U4985 (N_4985,N_4417,N_4452);
or U4986 (N_4986,N_4293,N_4499);
and U4987 (N_4987,N_4198,N_4039);
nor U4988 (N_4988,N_4039,N_4275);
xor U4989 (N_4989,N_4157,N_4398);
nand U4990 (N_4990,N_4092,N_4083);
or U4991 (N_4991,N_4134,N_4467);
and U4992 (N_4992,N_4309,N_4344);
and U4993 (N_4993,N_4358,N_4300);
nor U4994 (N_4994,N_4440,N_4162);
nand U4995 (N_4995,N_4226,N_4423);
or U4996 (N_4996,N_4311,N_4069);
xor U4997 (N_4997,N_4036,N_4097);
nor U4998 (N_4998,N_4237,N_4333);
or U4999 (N_4999,N_4061,N_4473);
xnor U5000 (N_5000,N_4714,N_4807);
or U5001 (N_5001,N_4747,N_4880);
xor U5002 (N_5002,N_4854,N_4943);
xor U5003 (N_5003,N_4611,N_4975);
and U5004 (N_5004,N_4543,N_4628);
xor U5005 (N_5005,N_4990,N_4554);
nor U5006 (N_5006,N_4555,N_4727);
nor U5007 (N_5007,N_4849,N_4671);
and U5008 (N_5008,N_4558,N_4841);
and U5009 (N_5009,N_4837,N_4514);
nor U5010 (N_5010,N_4636,N_4673);
and U5011 (N_5011,N_4893,N_4592);
nor U5012 (N_5012,N_4683,N_4662);
xnor U5013 (N_5013,N_4742,N_4879);
nor U5014 (N_5014,N_4559,N_4594);
xor U5015 (N_5015,N_4979,N_4719);
and U5016 (N_5016,N_4538,N_4780);
or U5017 (N_5017,N_4964,N_4732);
and U5018 (N_5018,N_4899,N_4755);
nand U5019 (N_5019,N_4947,N_4878);
and U5020 (N_5020,N_4697,N_4877);
xnor U5021 (N_5021,N_4756,N_4677);
or U5022 (N_5022,N_4960,N_4888);
xor U5023 (N_5023,N_4778,N_4912);
xor U5024 (N_5024,N_4895,N_4630);
or U5025 (N_5025,N_4796,N_4501);
nor U5026 (N_5026,N_4651,N_4550);
or U5027 (N_5027,N_4822,N_4918);
xor U5028 (N_5028,N_4632,N_4506);
and U5029 (N_5029,N_4761,N_4509);
and U5030 (N_5030,N_4871,N_4722);
xnor U5031 (N_5031,N_4534,N_4634);
xor U5032 (N_5032,N_4900,N_4825);
and U5033 (N_5033,N_4643,N_4766);
xnor U5034 (N_5034,N_4513,N_4887);
or U5035 (N_5035,N_4640,N_4711);
and U5036 (N_5036,N_4522,N_4998);
or U5037 (N_5037,N_4954,N_4674);
or U5038 (N_5038,N_4901,N_4903);
nor U5039 (N_5039,N_4838,N_4539);
and U5040 (N_5040,N_4799,N_4801);
nor U5041 (N_5041,N_4731,N_4598);
nor U5042 (N_5042,N_4569,N_4813);
xor U5043 (N_5043,N_4852,N_4627);
nand U5044 (N_5044,N_4929,N_4916);
and U5045 (N_5045,N_4988,N_4763);
nand U5046 (N_5046,N_4886,N_4610);
xor U5047 (N_5047,N_4641,N_4845);
xnor U5048 (N_5048,N_4659,N_4890);
or U5049 (N_5049,N_4795,N_4804);
nand U5050 (N_5050,N_4941,N_4521);
and U5051 (N_5051,N_4810,N_4779);
nand U5052 (N_5052,N_4721,N_4696);
xor U5053 (N_5053,N_4782,N_4664);
and U5054 (N_5054,N_4737,N_4987);
or U5055 (N_5055,N_4760,N_4533);
and U5056 (N_5056,N_4773,N_4787);
and U5057 (N_5057,N_4821,N_4607);
and U5058 (N_5058,N_4638,N_4648);
nand U5059 (N_5059,N_4580,N_4812);
and U5060 (N_5060,N_4847,N_4604);
or U5061 (N_5061,N_4973,N_4743);
xnor U5062 (N_5062,N_4986,N_4827);
nor U5063 (N_5063,N_4736,N_4974);
nor U5064 (N_5064,N_4842,N_4919);
and U5065 (N_5065,N_4968,N_4589);
nor U5066 (N_5066,N_4991,N_4599);
nand U5067 (N_5067,N_4794,N_4826);
and U5068 (N_5068,N_4819,N_4527);
xnor U5069 (N_5069,N_4791,N_4989);
and U5070 (N_5070,N_4959,N_4944);
and U5071 (N_5071,N_4889,N_4585);
and U5072 (N_5072,N_4586,N_4823);
or U5073 (N_5073,N_4980,N_4524);
nor U5074 (N_5074,N_4818,N_4925);
nor U5075 (N_5075,N_4875,N_4902);
nand U5076 (N_5076,N_4920,N_4820);
xor U5077 (N_5077,N_4931,N_4713);
nor U5078 (N_5078,N_4617,N_4578);
nand U5079 (N_5079,N_4689,N_4897);
nand U5080 (N_5080,N_4690,N_4999);
xor U5081 (N_5081,N_4562,N_4684);
xor U5082 (N_5082,N_4802,N_4809);
or U5083 (N_5083,N_4525,N_4882);
or U5084 (N_5084,N_4772,N_4734);
nand U5085 (N_5085,N_4551,N_4588);
xnor U5086 (N_5086,N_4762,N_4557);
nor U5087 (N_5087,N_4831,N_4996);
or U5088 (N_5088,N_4603,N_4751);
and U5089 (N_5089,N_4981,N_4595);
or U5090 (N_5090,N_4940,N_4858);
nand U5091 (N_5091,N_4518,N_4952);
nand U5092 (N_5092,N_4574,N_4962);
nand U5093 (N_5093,N_4503,N_4631);
and U5094 (N_5094,N_4656,N_4834);
and U5095 (N_5095,N_4507,N_4950);
nor U5096 (N_5096,N_4548,N_4767);
or U5097 (N_5097,N_4769,N_4654);
nand U5098 (N_5098,N_4618,N_4606);
xor U5099 (N_5099,N_4695,N_4730);
xor U5100 (N_5100,N_4701,N_4612);
xnor U5101 (N_5101,N_4765,N_4520);
or U5102 (N_5102,N_4857,N_4913);
nor U5103 (N_5103,N_4698,N_4536);
or U5104 (N_5104,N_4932,N_4789);
or U5105 (N_5105,N_4705,N_4945);
nand U5106 (N_5106,N_4572,N_4775);
nand U5107 (N_5107,N_4982,N_4560);
and U5108 (N_5108,N_4786,N_4680);
nand U5109 (N_5109,N_4934,N_4844);
nor U5110 (N_5110,N_4939,N_4771);
and U5111 (N_5111,N_4862,N_4670);
xor U5112 (N_5112,N_4904,N_4971);
nand U5113 (N_5113,N_4839,N_4754);
and U5114 (N_5114,N_4564,N_4587);
nand U5115 (N_5115,N_4508,N_4957);
xnor U5116 (N_5116,N_4785,N_4647);
xnor U5117 (N_5117,N_4573,N_4679);
xnor U5118 (N_5118,N_4921,N_4556);
nor U5119 (N_5119,N_4675,N_4545);
or U5120 (N_5120,N_4639,N_4579);
and U5121 (N_5121,N_4876,N_4790);
xor U5122 (N_5122,N_4884,N_4652);
or U5123 (N_5123,N_4745,N_4828);
or U5124 (N_5124,N_4622,N_4972);
and U5125 (N_5125,N_4800,N_4541);
nand U5126 (N_5126,N_4702,N_4924);
or U5127 (N_5127,N_4891,N_4729);
nor U5128 (N_5128,N_4927,N_4892);
nand U5129 (N_5129,N_4911,N_4657);
or U5130 (N_5130,N_4576,N_4535);
and U5131 (N_5131,N_4709,N_4992);
nor U5132 (N_5132,N_4649,N_4609);
nand U5133 (N_5133,N_4582,N_4777);
xnor U5134 (N_5134,N_4600,N_4568);
or U5135 (N_5135,N_4859,N_4874);
xnor U5136 (N_5136,N_4566,N_4868);
nor U5137 (N_5137,N_4946,N_4629);
or U5138 (N_5138,N_4704,N_4829);
nor U5139 (N_5139,N_4860,N_4505);
nand U5140 (N_5140,N_4735,N_4577);
or U5141 (N_5141,N_4863,N_4542);
and U5142 (N_5142,N_4978,N_4753);
nand U5143 (N_5143,N_4726,N_4633);
xor U5144 (N_5144,N_4898,N_4855);
nand U5145 (N_5145,N_4956,N_4805);
and U5146 (N_5146,N_4936,N_4720);
or U5147 (N_5147,N_4915,N_4846);
and U5148 (N_5148,N_4835,N_4798);
nor U5149 (N_5149,N_4710,N_4870);
and U5150 (N_5150,N_4510,N_4626);
nand U5151 (N_5151,N_4864,N_4803);
or U5152 (N_5152,N_4758,N_4750);
nand U5153 (N_5153,N_4565,N_4700);
and U5154 (N_5154,N_4861,N_4824);
and U5155 (N_5155,N_4832,N_4853);
xnor U5156 (N_5156,N_4850,N_4644);
nor U5157 (N_5157,N_4792,N_4757);
xor U5158 (N_5158,N_4993,N_4694);
nor U5159 (N_5159,N_4984,N_4517);
nor U5160 (N_5160,N_4867,N_4770);
or U5161 (N_5161,N_4584,N_4693);
or U5162 (N_5162,N_4816,N_4646);
xor U5163 (N_5163,N_4635,N_4699);
xor U5164 (N_5164,N_4793,N_4917);
nand U5165 (N_5165,N_4797,N_4723);
or U5166 (N_5166,N_4601,N_4531);
or U5167 (N_5167,N_4865,N_4930);
and U5168 (N_5168,N_4567,N_4937);
xnor U5169 (N_5169,N_4781,N_4687);
xnor U5170 (N_5170,N_4910,N_4716);
or U5171 (N_5171,N_4688,N_4752);
xor U5172 (N_5172,N_4969,N_4881);
xnor U5173 (N_5173,N_4977,N_4661);
xnor U5174 (N_5174,N_4749,N_4856);
xnor U5175 (N_5175,N_4815,N_4669);
nor U5176 (N_5176,N_4866,N_4963);
xnor U5177 (N_5177,N_4894,N_4616);
or U5178 (N_5178,N_4540,N_4570);
and U5179 (N_5179,N_4676,N_4808);
xor U5180 (N_5180,N_4914,N_4608);
and U5181 (N_5181,N_4715,N_4970);
xnor U5182 (N_5182,N_4537,N_4613);
nor U5183 (N_5183,N_4666,N_4907);
or U5184 (N_5184,N_4788,N_4806);
or U5185 (N_5185,N_4967,N_4830);
or U5186 (N_5186,N_4833,N_4624);
nor U5187 (N_5187,N_4544,N_4949);
nand U5188 (N_5188,N_4685,N_4995);
and U5189 (N_5189,N_4733,N_4681);
nor U5190 (N_5190,N_4528,N_4707);
and U5191 (N_5191,N_4909,N_4836);
or U5192 (N_5192,N_4935,N_4906);
nor U5193 (N_5193,N_4843,N_4668);
or U5194 (N_5194,N_4840,N_4615);
and U5195 (N_5195,N_4547,N_4642);
or U5196 (N_5196,N_4516,N_4728);
nor U5197 (N_5197,N_4994,N_4660);
and U5198 (N_5198,N_4908,N_4817);
xnor U5199 (N_5199,N_4645,N_4885);
nand U5200 (N_5200,N_4500,N_4602);
nand U5201 (N_5201,N_4511,N_4741);
and U5202 (N_5202,N_4953,N_4552);
or U5203 (N_5203,N_4515,N_4614);
or U5204 (N_5204,N_4658,N_4759);
or U5205 (N_5205,N_4965,N_4623);
and U5206 (N_5206,N_4637,N_4896);
or U5207 (N_5207,N_4961,N_4512);
and U5208 (N_5208,N_4703,N_4619);
xor U5209 (N_5209,N_4571,N_4814);
and U5210 (N_5210,N_4682,N_4625);
or U5211 (N_5211,N_4575,N_4655);
nor U5212 (N_5212,N_4948,N_4958);
or U5213 (N_5213,N_4581,N_4708);
nand U5214 (N_5214,N_4739,N_4593);
xor U5215 (N_5215,N_4997,N_4869);
and U5216 (N_5216,N_4764,N_4663);
xor U5217 (N_5217,N_4678,N_4596);
nand U5218 (N_5218,N_4553,N_4621);
nor U5219 (N_5219,N_4740,N_4590);
and U5220 (N_5220,N_4922,N_4717);
and U5221 (N_5221,N_4620,N_4768);
and U5222 (N_5222,N_4583,N_4597);
nand U5223 (N_5223,N_4691,N_4976);
xor U5224 (N_5224,N_4783,N_4724);
nand U5225 (N_5225,N_4738,N_4951);
nor U5226 (N_5226,N_4672,N_4872);
xor U5227 (N_5227,N_4985,N_4563);
nand U5228 (N_5228,N_4938,N_4546);
xnor U5229 (N_5229,N_4665,N_4653);
nor U5230 (N_5230,N_4650,N_4873);
nor U5231 (N_5231,N_4923,N_4725);
nor U5232 (N_5232,N_4955,N_4811);
or U5233 (N_5233,N_4776,N_4942);
nor U5234 (N_5234,N_4706,N_4692);
and U5235 (N_5235,N_4526,N_4746);
and U5236 (N_5236,N_4532,N_4529);
xor U5237 (N_5237,N_4519,N_4851);
or U5238 (N_5238,N_4523,N_4549);
or U5239 (N_5239,N_4667,N_4748);
xor U5240 (N_5240,N_4605,N_4712);
or U5241 (N_5241,N_4530,N_4933);
and U5242 (N_5242,N_4905,N_4502);
nand U5243 (N_5243,N_4784,N_4928);
or U5244 (N_5244,N_4774,N_4926);
or U5245 (N_5245,N_4504,N_4718);
xnor U5246 (N_5246,N_4686,N_4883);
xnor U5247 (N_5247,N_4591,N_4744);
xnor U5248 (N_5248,N_4848,N_4561);
and U5249 (N_5249,N_4966,N_4983);
and U5250 (N_5250,N_4840,N_4617);
and U5251 (N_5251,N_4773,N_4664);
xnor U5252 (N_5252,N_4958,N_4915);
or U5253 (N_5253,N_4538,N_4814);
and U5254 (N_5254,N_4612,N_4986);
nand U5255 (N_5255,N_4670,N_4744);
or U5256 (N_5256,N_4957,N_4657);
or U5257 (N_5257,N_4891,N_4722);
nand U5258 (N_5258,N_4662,N_4630);
nor U5259 (N_5259,N_4550,N_4681);
nor U5260 (N_5260,N_4633,N_4502);
and U5261 (N_5261,N_4848,N_4971);
and U5262 (N_5262,N_4654,N_4776);
or U5263 (N_5263,N_4639,N_4945);
nor U5264 (N_5264,N_4908,N_4840);
and U5265 (N_5265,N_4856,N_4532);
or U5266 (N_5266,N_4556,N_4508);
nand U5267 (N_5267,N_4987,N_4759);
and U5268 (N_5268,N_4960,N_4805);
nor U5269 (N_5269,N_4703,N_4978);
nand U5270 (N_5270,N_4863,N_4794);
or U5271 (N_5271,N_4837,N_4925);
and U5272 (N_5272,N_4925,N_4701);
and U5273 (N_5273,N_4982,N_4709);
nand U5274 (N_5274,N_4628,N_4820);
nand U5275 (N_5275,N_4954,N_4732);
nand U5276 (N_5276,N_4566,N_4819);
or U5277 (N_5277,N_4606,N_4815);
xor U5278 (N_5278,N_4654,N_4961);
nor U5279 (N_5279,N_4670,N_4906);
nor U5280 (N_5280,N_4698,N_4734);
nand U5281 (N_5281,N_4512,N_4576);
xor U5282 (N_5282,N_4555,N_4960);
xor U5283 (N_5283,N_4778,N_4510);
or U5284 (N_5284,N_4956,N_4848);
nand U5285 (N_5285,N_4953,N_4901);
or U5286 (N_5286,N_4748,N_4991);
and U5287 (N_5287,N_4823,N_4605);
nor U5288 (N_5288,N_4797,N_4595);
or U5289 (N_5289,N_4782,N_4742);
xnor U5290 (N_5290,N_4971,N_4942);
nand U5291 (N_5291,N_4505,N_4508);
nor U5292 (N_5292,N_4688,N_4720);
nand U5293 (N_5293,N_4609,N_4772);
or U5294 (N_5294,N_4648,N_4708);
and U5295 (N_5295,N_4848,N_4853);
nand U5296 (N_5296,N_4795,N_4582);
xnor U5297 (N_5297,N_4511,N_4531);
nand U5298 (N_5298,N_4862,N_4985);
or U5299 (N_5299,N_4536,N_4510);
and U5300 (N_5300,N_4938,N_4639);
nand U5301 (N_5301,N_4591,N_4545);
and U5302 (N_5302,N_4657,N_4503);
and U5303 (N_5303,N_4793,N_4559);
or U5304 (N_5304,N_4555,N_4926);
and U5305 (N_5305,N_4804,N_4537);
nand U5306 (N_5306,N_4997,N_4561);
nor U5307 (N_5307,N_4929,N_4626);
nand U5308 (N_5308,N_4800,N_4894);
and U5309 (N_5309,N_4658,N_4511);
nand U5310 (N_5310,N_4782,N_4709);
nor U5311 (N_5311,N_4883,N_4724);
xor U5312 (N_5312,N_4634,N_4615);
or U5313 (N_5313,N_4943,N_4830);
nor U5314 (N_5314,N_4794,N_4619);
nand U5315 (N_5315,N_4684,N_4966);
xor U5316 (N_5316,N_4623,N_4926);
nand U5317 (N_5317,N_4856,N_4727);
and U5318 (N_5318,N_4742,N_4715);
nand U5319 (N_5319,N_4598,N_4556);
xor U5320 (N_5320,N_4524,N_4706);
and U5321 (N_5321,N_4825,N_4891);
nand U5322 (N_5322,N_4826,N_4542);
nor U5323 (N_5323,N_4787,N_4794);
and U5324 (N_5324,N_4601,N_4786);
nor U5325 (N_5325,N_4790,N_4993);
or U5326 (N_5326,N_4830,N_4608);
or U5327 (N_5327,N_4539,N_4839);
and U5328 (N_5328,N_4870,N_4746);
nand U5329 (N_5329,N_4941,N_4846);
nor U5330 (N_5330,N_4825,N_4567);
nor U5331 (N_5331,N_4875,N_4719);
xnor U5332 (N_5332,N_4845,N_4740);
and U5333 (N_5333,N_4644,N_4812);
xor U5334 (N_5334,N_4578,N_4703);
and U5335 (N_5335,N_4964,N_4840);
or U5336 (N_5336,N_4616,N_4669);
nor U5337 (N_5337,N_4960,N_4832);
nand U5338 (N_5338,N_4755,N_4595);
nand U5339 (N_5339,N_4804,N_4799);
xnor U5340 (N_5340,N_4530,N_4816);
xor U5341 (N_5341,N_4710,N_4522);
nor U5342 (N_5342,N_4677,N_4981);
xor U5343 (N_5343,N_4872,N_4952);
nand U5344 (N_5344,N_4744,N_4995);
nand U5345 (N_5345,N_4816,N_4511);
nand U5346 (N_5346,N_4605,N_4909);
xnor U5347 (N_5347,N_4941,N_4981);
nor U5348 (N_5348,N_4870,N_4503);
nand U5349 (N_5349,N_4622,N_4942);
or U5350 (N_5350,N_4908,N_4693);
and U5351 (N_5351,N_4720,N_4976);
nor U5352 (N_5352,N_4543,N_4948);
xor U5353 (N_5353,N_4684,N_4644);
nor U5354 (N_5354,N_4886,N_4936);
nor U5355 (N_5355,N_4810,N_4688);
xnor U5356 (N_5356,N_4561,N_4635);
or U5357 (N_5357,N_4518,N_4864);
or U5358 (N_5358,N_4675,N_4609);
or U5359 (N_5359,N_4616,N_4841);
nor U5360 (N_5360,N_4505,N_4642);
nor U5361 (N_5361,N_4979,N_4887);
nand U5362 (N_5362,N_4645,N_4817);
xor U5363 (N_5363,N_4675,N_4582);
and U5364 (N_5364,N_4704,N_4888);
xor U5365 (N_5365,N_4789,N_4727);
or U5366 (N_5366,N_4946,N_4623);
xor U5367 (N_5367,N_4604,N_4606);
xor U5368 (N_5368,N_4751,N_4520);
nand U5369 (N_5369,N_4867,N_4638);
nor U5370 (N_5370,N_4654,N_4798);
xnor U5371 (N_5371,N_4647,N_4714);
and U5372 (N_5372,N_4764,N_4522);
and U5373 (N_5373,N_4590,N_4794);
or U5374 (N_5374,N_4864,N_4779);
nand U5375 (N_5375,N_4704,N_4993);
xnor U5376 (N_5376,N_4771,N_4547);
nand U5377 (N_5377,N_4566,N_4646);
nand U5378 (N_5378,N_4848,N_4984);
xor U5379 (N_5379,N_4974,N_4566);
nor U5380 (N_5380,N_4985,N_4800);
nand U5381 (N_5381,N_4604,N_4551);
nor U5382 (N_5382,N_4895,N_4912);
xor U5383 (N_5383,N_4823,N_4761);
or U5384 (N_5384,N_4863,N_4844);
or U5385 (N_5385,N_4915,N_4624);
nor U5386 (N_5386,N_4658,N_4630);
nor U5387 (N_5387,N_4760,N_4777);
nor U5388 (N_5388,N_4688,N_4871);
xnor U5389 (N_5389,N_4849,N_4581);
xnor U5390 (N_5390,N_4870,N_4518);
and U5391 (N_5391,N_4727,N_4923);
nor U5392 (N_5392,N_4545,N_4719);
or U5393 (N_5393,N_4647,N_4537);
and U5394 (N_5394,N_4934,N_4574);
or U5395 (N_5395,N_4510,N_4679);
nor U5396 (N_5396,N_4758,N_4614);
or U5397 (N_5397,N_4909,N_4704);
nand U5398 (N_5398,N_4881,N_4991);
and U5399 (N_5399,N_4664,N_4505);
xor U5400 (N_5400,N_4999,N_4958);
or U5401 (N_5401,N_4787,N_4655);
or U5402 (N_5402,N_4567,N_4617);
or U5403 (N_5403,N_4599,N_4698);
xor U5404 (N_5404,N_4635,N_4693);
nor U5405 (N_5405,N_4668,N_4868);
nor U5406 (N_5406,N_4577,N_4977);
nor U5407 (N_5407,N_4607,N_4710);
xnor U5408 (N_5408,N_4865,N_4983);
or U5409 (N_5409,N_4502,N_4642);
xor U5410 (N_5410,N_4801,N_4625);
nand U5411 (N_5411,N_4528,N_4699);
nand U5412 (N_5412,N_4601,N_4515);
nand U5413 (N_5413,N_4894,N_4633);
nor U5414 (N_5414,N_4843,N_4636);
nor U5415 (N_5415,N_4647,N_4528);
xnor U5416 (N_5416,N_4515,N_4708);
nor U5417 (N_5417,N_4592,N_4658);
xnor U5418 (N_5418,N_4836,N_4958);
xnor U5419 (N_5419,N_4741,N_4814);
nor U5420 (N_5420,N_4935,N_4713);
or U5421 (N_5421,N_4633,N_4774);
and U5422 (N_5422,N_4962,N_4532);
and U5423 (N_5423,N_4658,N_4833);
xor U5424 (N_5424,N_4904,N_4842);
nand U5425 (N_5425,N_4599,N_4576);
nor U5426 (N_5426,N_4807,N_4540);
or U5427 (N_5427,N_4864,N_4736);
xnor U5428 (N_5428,N_4901,N_4628);
and U5429 (N_5429,N_4893,N_4783);
nand U5430 (N_5430,N_4845,N_4982);
and U5431 (N_5431,N_4681,N_4797);
xor U5432 (N_5432,N_4506,N_4817);
and U5433 (N_5433,N_4811,N_4640);
or U5434 (N_5434,N_4598,N_4849);
or U5435 (N_5435,N_4902,N_4824);
and U5436 (N_5436,N_4738,N_4748);
or U5437 (N_5437,N_4862,N_4894);
nor U5438 (N_5438,N_4548,N_4870);
xnor U5439 (N_5439,N_4723,N_4839);
nor U5440 (N_5440,N_4909,N_4812);
and U5441 (N_5441,N_4845,N_4589);
nor U5442 (N_5442,N_4665,N_4690);
nand U5443 (N_5443,N_4839,N_4583);
and U5444 (N_5444,N_4685,N_4895);
and U5445 (N_5445,N_4763,N_4502);
nor U5446 (N_5446,N_4500,N_4753);
nand U5447 (N_5447,N_4530,N_4788);
and U5448 (N_5448,N_4910,N_4946);
xor U5449 (N_5449,N_4511,N_4738);
nand U5450 (N_5450,N_4521,N_4904);
and U5451 (N_5451,N_4648,N_4869);
and U5452 (N_5452,N_4843,N_4915);
xor U5453 (N_5453,N_4978,N_4924);
and U5454 (N_5454,N_4762,N_4516);
or U5455 (N_5455,N_4693,N_4833);
nand U5456 (N_5456,N_4748,N_4834);
nor U5457 (N_5457,N_4903,N_4966);
nand U5458 (N_5458,N_4872,N_4900);
nor U5459 (N_5459,N_4661,N_4940);
or U5460 (N_5460,N_4692,N_4889);
xor U5461 (N_5461,N_4821,N_4601);
xor U5462 (N_5462,N_4900,N_4507);
xnor U5463 (N_5463,N_4756,N_4747);
nand U5464 (N_5464,N_4618,N_4919);
or U5465 (N_5465,N_4996,N_4761);
or U5466 (N_5466,N_4534,N_4527);
and U5467 (N_5467,N_4959,N_4853);
xor U5468 (N_5468,N_4959,N_4770);
and U5469 (N_5469,N_4857,N_4904);
and U5470 (N_5470,N_4897,N_4619);
and U5471 (N_5471,N_4917,N_4739);
nor U5472 (N_5472,N_4892,N_4756);
nor U5473 (N_5473,N_4791,N_4936);
nand U5474 (N_5474,N_4840,N_4846);
nand U5475 (N_5475,N_4802,N_4811);
xnor U5476 (N_5476,N_4995,N_4643);
nor U5477 (N_5477,N_4997,N_4995);
and U5478 (N_5478,N_4946,N_4899);
or U5479 (N_5479,N_4626,N_4556);
xnor U5480 (N_5480,N_4752,N_4952);
xnor U5481 (N_5481,N_4512,N_4614);
xor U5482 (N_5482,N_4625,N_4884);
and U5483 (N_5483,N_4669,N_4749);
nor U5484 (N_5484,N_4971,N_4835);
and U5485 (N_5485,N_4889,N_4716);
nand U5486 (N_5486,N_4543,N_4530);
nand U5487 (N_5487,N_4670,N_4915);
xnor U5488 (N_5488,N_4809,N_4963);
nand U5489 (N_5489,N_4687,N_4999);
and U5490 (N_5490,N_4935,N_4832);
and U5491 (N_5491,N_4972,N_4865);
and U5492 (N_5492,N_4541,N_4830);
or U5493 (N_5493,N_4600,N_4734);
and U5494 (N_5494,N_4883,N_4513);
or U5495 (N_5495,N_4528,N_4654);
nor U5496 (N_5496,N_4536,N_4892);
or U5497 (N_5497,N_4540,N_4805);
or U5498 (N_5498,N_4897,N_4969);
or U5499 (N_5499,N_4883,N_4745);
nand U5500 (N_5500,N_5134,N_5079);
or U5501 (N_5501,N_5164,N_5109);
and U5502 (N_5502,N_5437,N_5274);
nor U5503 (N_5503,N_5220,N_5102);
nand U5504 (N_5504,N_5105,N_5275);
nor U5505 (N_5505,N_5222,N_5315);
nor U5506 (N_5506,N_5231,N_5090);
nand U5507 (N_5507,N_5070,N_5168);
or U5508 (N_5508,N_5343,N_5451);
nand U5509 (N_5509,N_5279,N_5373);
nor U5510 (N_5510,N_5013,N_5365);
and U5511 (N_5511,N_5285,N_5172);
xnor U5512 (N_5512,N_5160,N_5304);
and U5513 (N_5513,N_5156,N_5421);
and U5514 (N_5514,N_5397,N_5417);
nand U5515 (N_5515,N_5449,N_5040);
nand U5516 (N_5516,N_5225,N_5265);
and U5517 (N_5517,N_5133,N_5051);
nor U5518 (N_5518,N_5122,N_5277);
or U5519 (N_5519,N_5428,N_5376);
nand U5520 (N_5520,N_5310,N_5065);
nor U5521 (N_5521,N_5224,N_5186);
nand U5522 (N_5522,N_5347,N_5472);
nand U5523 (N_5523,N_5015,N_5498);
nand U5524 (N_5524,N_5250,N_5114);
xnor U5525 (N_5525,N_5151,N_5107);
xor U5526 (N_5526,N_5414,N_5434);
xor U5527 (N_5527,N_5366,N_5111);
nand U5528 (N_5528,N_5263,N_5100);
or U5529 (N_5529,N_5426,N_5104);
and U5530 (N_5530,N_5423,N_5321);
xnor U5531 (N_5531,N_5063,N_5311);
nor U5532 (N_5532,N_5495,N_5470);
nand U5533 (N_5533,N_5142,N_5061);
nand U5534 (N_5534,N_5386,N_5001);
nor U5535 (N_5535,N_5429,N_5077);
nor U5536 (N_5536,N_5064,N_5149);
or U5537 (N_5537,N_5328,N_5112);
nor U5538 (N_5538,N_5488,N_5244);
nand U5539 (N_5539,N_5214,N_5062);
nor U5540 (N_5540,N_5413,N_5184);
nor U5541 (N_5541,N_5076,N_5067);
nand U5542 (N_5542,N_5033,N_5054);
and U5543 (N_5543,N_5045,N_5095);
and U5544 (N_5544,N_5368,N_5273);
and U5545 (N_5545,N_5035,N_5302);
xnor U5546 (N_5546,N_5471,N_5409);
and U5547 (N_5547,N_5097,N_5034);
nand U5548 (N_5548,N_5210,N_5454);
nor U5549 (N_5549,N_5336,N_5329);
nand U5550 (N_5550,N_5401,N_5180);
nor U5551 (N_5551,N_5226,N_5233);
and U5552 (N_5552,N_5075,N_5126);
xor U5553 (N_5553,N_5374,N_5125);
nor U5554 (N_5554,N_5453,N_5084);
nor U5555 (N_5555,N_5016,N_5405);
nor U5556 (N_5556,N_5476,N_5467);
nor U5557 (N_5557,N_5206,N_5031);
nand U5558 (N_5558,N_5003,N_5269);
nor U5559 (N_5559,N_5309,N_5412);
and U5560 (N_5560,N_5249,N_5389);
nand U5561 (N_5561,N_5357,N_5139);
nand U5562 (N_5562,N_5348,N_5262);
nand U5563 (N_5563,N_5294,N_5096);
or U5564 (N_5564,N_5036,N_5438);
xor U5565 (N_5565,N_5485,N_5021);
nor U5566 (N_5566,N_5286,N_5110);
xnor U5567 (N_5567,N_5327,N_5137);
nand U5568 (N_5568,N_5318,N_5018);
and U5569 (N_5569,N_5439,N_5176);
nand U5570 (N_5570,N_5173,N_5213);
nor U5571 (N_5571,N_5243,N_5322);
and U5572 (N_5572,N_5420,N_5085);
xnor U5573 (N_5573,N_5404,N_5130);
or U5574 (N_5574,N_5246,N_5431);
nor U5575 (N_5575,N_5161,N_5227);
nor U5576 (N_5576,N_5446,N_5195);
or U5577 (N_5577,N_5291,N_5332);
and U5578 (N_5578,N_5254,N_5422);
nand U5579 (N_5579,N_5144,N_5146);
nand U5580 (N_5580,N_5006,N_5375);
or U5581 (N_5581,N_5387,N_5167);
xnor U5582 (N_5582,N_5435,N_5427);
or U5583 (N_5583,N_5266,N_5433);
and U5584 (N_5584,N_5325,N_5153);
or U5585 (N_5585,N_5020,N_5333);
nand U5586 (N_5586,N_5120,N_5185);
and U5587 (N_5587,N_5166,N_5356);
xor U5588 (N_5588,N_5152,N_5209);
xor U5589 (N_5589,N_5457,N_5359);
nand U5590 (N_5590,N_5379,N_5352);
xor U5591 (N_5591,N_5190,N_5255);
and U5592 (N_5592,N_5253,N_5484);
and U5593 (N_5593,N_5290,N_5086);
and U5594 (N_5594,N_5008,N_5300);
and U5595 (N_5595,N_5074,N_5101);
xnor U5596 (N_5596,N_5355,N_5478);
xor U5597 (N_5597,N_5205,N_5236);
nand U5598 (N_5598,N_5459,N_5115);
and U5599 (N_5599,N_5030,N_5344);
xnor U5600 (N_5600,N_5448,N_5402);
nor U5601 (N_5601,N_5022,N_5340);
nor U5602 (N_5602,N_5023,N_5464);
xnor U5603 (N_5603,N_5394,N_5460);
or U5604 (N_5604,N_5043,N_5271);
nor U5605 (N_5605,N_5462,N_5466);
or U5606 (N_5606,N_5301,N_5408);
or U5607 (N_5607,N_5248,N_5455);
nor U5608 (N_5608,N_5261,N_5014);
xor U5609 (N_5609,N_5432,N_5251);
nand U5610 (N_5610,N_5444,N_5278);
nand U5611 (N_5611,N_5191,N_5298);
and U5612 (N_5612,N_5007,N_5053);
or U5613 (N_5613,N_5135,N_5393);
xor U5614 (N_5614,N_5025,N_5383);
or U5615 (N_5615,N_5313,N_5046);
xor U5616 (N_5616,N_5192,N_5369);
nand U5617 (N_5617,N_5479,N_5145);
xnor U5618 (N_5618,N_5042,N_5335);
nand U5619 (N_5619,N_5430,N_5299);
and U5620 (N_5620,N_5496,N_5252);
and U5621 (N_5621,N_5371,N_5163);
or U5622 (N_5622,N_5232,N_5204);
and U5623 (N_5623,N_5113,N_5403);
nand U5624 (N_5624,N_5489,N_5307);
xor U5625 (N_5625,N_5406,N_5492);
or U5626 (N_5626,N_5159,N_5364);
nand U5627 (N_5627,N_5187,N_5268);
and U5628 (N_5628,N_5181,N_5038);
or U5629 (N_5629,N_5239,N_5055);
or U5630 (N_5630,N_5229,N_5039);
nor U5631 (N_5631,N_5400,N_5098);
xnor U5632 (N_5632,N_5380,N_5486);
xnor U5633 (N_5633,N_5258,N_5092);
nor U5634 (N_5634,N_5456,N_5238);
nor U5635 (N_5635,N_5491,N_5330);
and U5636 (N_5636,N_5490,N_5169);
xor U5637 (N_5637,N_5060,N_5463);
xnor U5638 (N_5638,N_5494,N_5284);
xnor U5639 (N_5639,N_5044,N_5080);
and U5640 (N_5640,N_5103,N_5497);
and U5641 (N_5641,N_5068,N_5287);
nor U5642 (N_5642,N_5201,N_5468);
nand U5643 (N_5643,N_5019,N_5481);
nand U5644 (N_5644,N_5245,N_5048);
xnor U5645 (N_5645,N_5424,N_5257);
nand U5646 (N_5646,N_5320,N_5323);
and U5647 (N_5647,N_5155,N_5223);
nand U5648 (N_5648,N_5211,N_5199);
nand U5649 (N_5649,N_5367,N_5419);
nand U5650 (N_5650,N_5240,N_5469);
and U5651 (N_5651,N_5087,N_5477);
nand U5652 (N_5652,N_5041,N_5132);
and U5653 (N_5653,N_5017,N_5136);
or U5654 (N_5654,N_5078,N_5351);
nor U5655 (N_5655,N_5150,N_5140);
and U5656 (N_5656,N_5372,N_5212);
or U5657 (N_5657,N_5147,N_5121);
nand U5658 (N_5658,N_5306,N_5395);
nand U5659 (N_5659,N_5131,N_5475);
and U5660 (N_5660,N_5083,N_5215);
nor U5661 (N_5661,N_5465,N_5081);
nand U5662 (N_5662,N_5200,N_5119);
nand U5663 (N_5663,N_5411,N_5000);
xnor U5664 (N_5664,N_5093,N_5058);
and U5665 (N_5665,N_5337,N_5117);
nor U5666 (N_5666,N_5218,N_5237);
and U5667 (N_5667,N_5363,N_5171);
xor U5668 (N_5668,N_5452,N_5174);
nand U5669 (N_5669,N_5073,N_5342);
xor U5670 (N_5670,N_5407,N_5312);
xnor U5671 (N_5671,N_5148,N_5235);
nand U5672 (N_5672,N_5388,N_5267);
or U5673 (N_5673,N_5303,N_5179);
nand U5674 (N_5674,N_5256,N_5183);
or U5675 (N_5675,N_5099,N_5341);
nor U5676 (N_5676,N_5382,N_5319);
nor U5677 (N_5677,N_5260,N_5370);
xnor U5678 (N_5678,N_5004,N_5123);
nor U5679 (N_5679,N_5138,N_5334);
nand U5680 (N_5680,N_5499,N_5272);
or U5681 (N_5681,N_5094,N_5443);
and U5682 (N_5682,N_5118,N_5165);
nand U5683 (N_5683,N_5188,N_5230);
nor U5684 (N_5684,N_5202,N_5349);
nand U5685 (N_5685,N_5441,N_5416);
nor U5686 (N_5686,N_5182,N_5141);
or U5687 (N_5687,N_5331,N_5339);
or U5688 (N_5688,N_5047,N_5089);
or U5689 (N_5689,N_5392,N_5354);
and U5690 (N_5690,N_5436,N_5203);
nor U5691 (N_5691,N_5196,N_5360);
nand U5692 (N_5692,N_5338,N_5276);
xor U5693 (N_5693,N_5281,N_5066);
xor U5694 (N_5694,N_5295,N_5296);
nand U5695 (N_5695,N_5057,N_5129);
or U5696 (N_5696,N_5072,N_5217);
xor U5697 (N_5697,N_5378,N_5162);
or U5698 (N_5698,N_5059,N_5005);
nor U5699 (N_5699,N_5415,N_5106);
and U5700 (N_5700,N_5308,N_5208);
or U5701 (N_5701,N_5399,N_5127);
nor U5702 (N_5702,N_5450,N_5293);
and U5703 (N_5703,N_5088,N_5474);
and U5704 (N_5704,N_5193,N_5410);
or U5705 (N_5705,N_5082,N_5280);
xor U5706 (N_5706,N_5346,N_5247);
or U5707 (N_5707,N_5241,N_5011);
or U5708 (N_5708,N_5050,N_5297);
or U5709 (N_5709,N_5197,N_5390);
nor U5710 (N_5710,N_5483,N_5361);
xnor U5711 (N_5711,N_5157,N_5385);
nor U5712 (N_5712,N_5010,N_5398);
or U5713 (N_5713,N_5024,N_5108);
nor U5714 (N_5714,N_5228,N_5305);
xor U5715 (N_5715,N_5447,N_5049);
xor U5716 (N_5716,N_5353,N_5377);
nand U5717 (N_5717,N_5158,N_5052);
nor U5718 (N_5718,N_5292,N_5154);
xnor U5719 (N_5719,N_5259,N_5009);
and U5720 (N_5720,N_5314,N_5289);
nor U5721 (N_5721,N_5116,N_5445);
nand U5722 (N_5722,N_5317,N_5170);
or U5723 (N_5723,N_5216,N_5069);
nand U5724 (N_5724,N_5124,N_5487);
nor U5725 (N_5725,N_5324,N_5071);
and U5726 (N_5726,N_5425,N_5270);
and U5727 (N_5727,N_5027,N_5461);
nor U5728 (N_5728,N_5283,N_5242);
and U5729 (N_5729,N_5194,N_5282);
nand U5730 (N_5730,N_5381,N_5391);
nor U5731 (N_5731,N_5143,N_5418);
xor U5732 (N_5732,N_5091,N_5037);
or U5733 (N_5733,N_5128,N_5482);
and U5734 (N_5734,N_5345,N_5326);
xor U5735 (N_5735,N_5442,N_5012);
and U5736 (N_5736,N_5316,N_5002);
or U5737 (N_5737,N_5358,N_5219);
nor U5738 (N_5738,N_5175,N_5026);
nand U5739 (N_5739,N_5384,N_5264);
nor U5740 (N_5740,N_5198,N_5458);
nand U5741 (N_5741,N_5362,N_5473);
or U5742 (N_5742,N_5189,N_5234);
nor U5743 (N_5743,N_5178,N_5396);
nand U5744 (N_5744,N_5493,N_5350);
and U5745 (N_5745,N_5221,N_5028);
nor U5746 (N_5746,N_5480,N_5288);
or U5747 (N_5747,N_5056,N_5440);
nand U5748 (N_5748,N_5029,N_5177);
nor U5749 (N_5749,N_5032,N_5207);
or U5750 (N_5750,N_5494,N_5139);
nor U5751 (N_5751,N_5018,N_5233);
and U5752 (N_5752,N_5101,N_5290);
or U5753 (N_5753,N_5058,N_5211);
nor U5754 (N_5754,N_5334,N_5164);
nor U5755 (N_5755,N_5138,N_5234);
nand U5756 (N_5756,N_5287,N_5189);
and U5757 (N_5757,N_5374,N_5069);
nor U5758 (N_5758,N_5142,N_5237);
xnor U5759 (N_5759,N_5201,N_5251);
xnor U5760 (N_5760,N_5247,N_5010);
nor U5761 (N_5761,N_5143,N_5226);
nor U5762 (N_5762,N_5240,N_5147);
and U5763 (N_5763,N_5471,N_5042);
nand U5764 (N_5764,N_5354,N_5286);
or U5765 (N_5765,N_5406,N_5497);
or U5766 (N_5766,N_5441,N_5232);
nand U5767 (N_5767,N_5490,N_5297);
nor U5768 (N_5768,N_5277,N_5316);
and U5769 (N_5769,N_5359,N_5149);
xnor U5770 (N_5770,N_5041,N_5301);
nand U5771 (N_5771,N_5240,N_5472);
nand U5772 (N_5772,N_5128,N_5493);
nor U5773 (N_5773,N_5022,N_5399);
nor U5774 (N_5774,N_5491,N_5250);
or U5775 (N_5775,N_5365,N_5343);
and U5776 (N_5776,N_5296,N_5368);
nor U5777 (N_5777,N_5039,N_5323);
xnor U5778 (N_5778,N_5295,N_5162);
and U5779 (N_5779,N_5067,N_5218);
or U5780 (N_5780,N_5187,N_5215);
or U5781 (N_5781,N_5481,N_5015);
nand U5782 (N_5782,N_5044,N_5450);
nor U5783 (N_5783,N_5401,N_5358);
xnor U5784 (N_5784,N_5025,N_5034);
or U5785 (N_5785,N_5282,N_5428);
nor U5786 (N_5786,N_5332,N_5328);
and U5787 (N_5787,N_5018,N_5091);
nand U5788 (N_5788,N_5354,N_5200);
and U5789 (N_5789,N_5414,N_5413);
and U5790 (N_5790,N_5101,N_5333);
or U5791 (N_5791,N_5199,N_5053);
or U5792 (N_5792,N_5340,N_5242);
xnor U5793 (N_5793,N_5181,N_5205);
and U5794 (N_5794,N_5100,N_5033);
xnor U5795 (N_5795,N_5271,N_5479);
and U5796 (N_5796,N_5058,N_5172);
nor U5797 (N_5797,N_5264,N_5060);
nand U5798 (N_5798,N_5473,N_5347);
or U5799 (N_5799,N_5190,N_5361);
xor U5800 (N_5800,N_5112,N_5193);
nand U5801 (N_5801,N_5372,N_5249);
nand U5802 (N_5802,N_5460,N_5276);
nor U5803 (N_5803,N_5020,N_5264);
xor U5804 (N_5804,N_5012,N_5014);
nor U5805 (N_5805,N_5341,N_5438);
xor U5806 (N_5806,N_5060,N_5340);
nand U5807 (N_5807,N_5127,N_5471);
nand U5808 (N_5808,N_5212,N_5122);
xnor U5809 (N_5809,N_5325,N_5266);
xnor U5810 (N_5810,N_5109,N_5070);
or U5811 (N_5811,N_5357,N_5153);
or U5812 (N_5812,N_5244,N_5174);
or U5813 (N_5813,N_5042,N_5413);
xor U5814 (N_5814,N_5055,N_5262);
or U5815 (N_5815,N_5398,N_5045);
xnor U5816 (N_5816,N_5154,N_5326);
nor U5817 (N_5817,N_5017,N_5004);
and U5818 (N_5818,N_5149,N_5477);
nand U5819 (N_5819,N_5281,N_5371);
nand U5820 (N_5820,N_5421,N_5285);
or U5821 (N_5821,N_5099,N_5120);
or U5822 (N_5822,N_5423,N_5044);
xnor U5823 (N_5823,N_5090,N_5425);
xnor U5824 (N_5824,N_5335,N_5471);
xor U5825 (N_5825,N_5134,N_5250);
xnor U5826 (N_5826,N_5149,N_5320);
nor U5827 (N_5827,N_5359,N_5104);
and U5828 (N_5828,N_5420,N_5194);
nand U5829 (N_5829,N_5047,N_5297);
or U5830 (N_5830,N_5436,N_5163);
or U5831 (N_5831,N_5366,N_5326);
and U5832 (N_5832,N_5246,N_5091);
nor U5833 (N_5833,N_5122,N_5405);
xor U5834 (N_5834,N_5375,N_5474);
and U5835 (N_5835,N_5089,N_5421);
or U5836 (N_5836,N_5134,N_5076);
nand U5837 (N_5837,N_5150,N_5254);
nor U5838 (N_5838,N_5480,N_5316);
nor U5839 (N_5839,N_5193,N_5088);
and U5840 (N_5840,N_5312,N_5241);
nand U5841 (N_5841,N_5249,N_5335);
nand U5842 (N_5842,N_5260,N_5095);
nand U5843 (N_5843,N_5082,N_5484);
xnor U5844 (N_5844,N_5101,N_5093);
and U5845 (N_5845,N_5405,N_5032);
nand U5846 (N_5846,N_5436,N_5272);
xor U5847 (N_5847,N_5427,N_5323);
nor U5848 (N_5848,N_5406,N_5265);
and U5849 (N_5849,N_5172,N_5198);
xor U5850 (N_5850,N_5063,N_5261);
or U5851 (N_5851,N_5206,N_5377);
nand U5852 (N_5852,N_5258,N_5347);
and U5853 (N_5853,N_5034,N_5334);
xor U5854 (N_5854,N_5059,N_5077);
and U5855 (N_5855,N_5002,N_5355);
or U5856 (N_5856,N_5383,N_5348);
nor U5857 (N_5857,N_5314,N_5189);
nor U5858 (N_5858,N_5201,N_5331);
nand U5859 (N_5859,N_5074,N_5051);
nor U5860 (N_5860,N_5227,N_5152);
xnor U5861 (N_5861,N_5431,N_5335);
or U5862 (N_5862,N_5149,N_5160);
or U5863 (N_5863,N_5437,N_5076);
and U5864 (N_5864,N_5327,N_5073);
or U5865 (N_5865,N_5194,N_5160);
nor U5866 (N_5866,N_5233,N_5191);
nor U5867 (N_5867,N_5066,N_5087);
and U5868 (N_5868,N_5488,N_5283);
nand U5869 (N_5869,N_5074,N_5038);
or U5870 (N_5870,N_5217,N_5414);
and U5871 (N_5871,N_5191,N_5008);
or U5872 (N_5872,N_5298,N_5329);
or U5873 (N_5873,N_5267,N_5038);
xnor U5874 (N_5874,N_5194,N_5199);
and U5875 (N_5875,N_5083,N_5326);
nand U5876 (N_5876,N_5175,N_5121);
or U5877 (N_5877,N_5107,N_5270);
nand U5878 (N_5878,N_5297,N_5128);
or U5879 (N_5879,N_5001,N_5492);
or U5880 (N_5880,N_5312,N_5094);
or U5881 (N_5881,N_5156,N_5302);
nor U5882 (N_5882,N_5400,N_5421);
nand U5883 (N_5883,N_5150,N_5123);
or U5884 (N_5884,N_5425,N_5122);
nand U5885 (N_5885,N_5433,N_5078);
nand U5886 (N_5886,N_5133,N_5388);
nand U5887 (N_5887,N_5089,N_5091);
nand U5888 (N_5888,N_5086,N_5351);
and U5889 (N_5889,N_5113,N_5114);
nand U5890 (N_5890,N_5008,N_5236);
nor U5891 (N_5891,N_5024,N_5435);
nand U5892 (N_5892,N_5121,N_5484);
nor U5893 (N_5893,N_5170,N_5479);
xor U5894 (N_5894,N_5261,N_5370);
nor U5895 (N_5895,N_5297,N_5028);
xor U5896 (N_5896,N_5104,N_5235);
or U5897 (N_5897,N_5236,N_5054);
nand U5898 (N_5898,N_5218,N_5271);
nor U5899 (N_5899,N_5171,N_5002);
nand U5900 (N_5900,N_5215,N_5301);
and U5901 (N_5901,N_5117,N_5265);
or U5902 (N_5902,N_5038,N_5405);
or U5903 (N_5903,N_5435,N_5294);
nor U5904 (N_5904,N_5466,N_5037);
and U5905 (N_5905,N_5062,N_5162);
and U5906 (N_5906,N_5028,N_5112);
xnor U5907 (N_5907,N_5288,N_5192);
or U5908 (N_5908,N_5338,N_5241);
xnor U5909 (N_5909,N_5408,N_5484);
nand U5910 (N_5910,N_5070,N_5098);
and U5911 (N_5911,N_5110,N_5049);
xnor U5912 (N_5912,N_5335,N_5011);
and U5913 (N_5913,N_5174,N_5302);
or U5914 (N_5914,N_5207,N_5462);
nand U5915 (N_5915,N_5197,N_5032);
and U5916 (N_5916,N_5304,N_5348);
xnor U5917 (N_5917,N_5088,N_5318);
nand U5918 (N_5918,N_5417,N_5425);
xnor U5919 (N_5919,N_5459,N_5113);
nand U5920 (N_5920,N_5467,N_5252);
or U5921 (N_5921,N_5182,N_5434);
nand U5922 (N_5922,N_5064,N_5398);
and U5923 (N_5923,N_5464,N_5200);
and U5924 (N_5924,N_5011,N_5208);
xnor U5925 (N_5925,N_5481,N_5233);
and U5926 (N_5926,N_5049,N_5053);
nand U5927 (N_5927,N_5066,N_5201);
xnor U5928 (N_5928,N_5267,N_5065);
or U5929 (N_5929,N_5125,N_5080);
or U5930 (N_5930,N_5125,N_5150);
xor U5931 (N_5931,N_5404,N_5236);
xnor U5932 (N_5932,N_5129,N_5058);
or U5933 (N_5933,N_5235,N_5444);
or U5934 (N_5934,N_5217,N_5237);
xnor U5935 (N_5935,N_5358,N_5290);
nor U5936 (N_5936,N_5243,N_5354);
and U5937 (N_5937,N_5220,N_5209);
nor U5938 (N_5938,N_5048,N_5015);
nor U5939 (N_5939,N_5009,N_5190);
nor U5940 (N_5940,N_5171,N_5285);
nand U5941 (N_5941,N_5169,N_5387);
and U5942 (N_5942,N_5367,N_5334);
nand U5943 (N_5943,N_5037,N_5117);
xnor U5944 (N_5944,N_5048,N_5249);
and U5945 (N_5945,N_5285,N_5374);
nor U5946 (N_5946,N_5386,N_5421);
nor U5947 (N_5947,N_5303,N_5464);
and U5948 (N_5948,N_5327,N_5357);
or U5949 (N_5949,N_5024,N_5182);
nor U5950 (N_5950,N_5218,N_5486);
nand U5951 (N_5951,N_5358,N_5259);
xnor U5952 (N_5952,N_5449,N_5015);
xor U5953 (N_5953,N_5172,N_5363);
nor U5954 (N_5954,N_5459,N_5132);
xor U5955 (N_5955,N_5061,N_5223);
nor U5956 (N_5956,N_5470,N_5390);
or U5957 (N_5957,N_5483,N_5113);
xnor U5958 (N_5958,N_5443,N_5229);
or U5959 (N_5959,N_5195,N_5309);
xor U5960 (N_5960,N_5131,N_5351);
xnor U5961 (N_5961,N_5307,N_5469);
nor U5962 (N_5962,N_5160,N_5349);
xnor U5963 (N_5963,N_5259,N_5453);
or U5964 (N_5964,N_5289,N_5243);
xor U5965 (N_5965,N_5394,N_5190);
nor U5966 (N_5966,N_5076,N_5061);
nand U5967 (N_5967,N_5329,N_5437);
nor U5968 (N_5968,N_5494,N_5470);
xor U5969 (N_5969,N_5420,N_5355);
nor U5970 (N_5970,N_5199,N_5413);
nand U5971 (N_5971,N_5305,N_5166);
nor U5972 (N_5972,N_5372,N_5009);
nor U5973 (N_5973,N_5208,N_5275);
and U5974 (N_5974,N_5281,N_5099);
xnor U5975 (N_5975,N_5388,N_5336);
and U5976 (N_5976,N_5261,N_5255);
xnor U5977 (N_5977,N_5417,N_5028);
xnor U5978 (N_5978,N_5341,N_5232);
nor U5979 (N_5979,N_5284,N_5185);
xor U5980 (N_5980,N_5303,N_5496);
xor U5981 (N_5981,N_5068,N_5157);
and U5982 (N_5982,N_5196,N_5379);
xnor U5983 (N_5983,N_5300,N_5319);
or U5984 (N_5984,N_5392,N_5189);
nor U5985 (N_5985,N_5000,N_5423);
nor U5986 (N_5986,N_5323,N_5447);
or U5987 (N_5987,N_5324,N_5088);
and U5988 (N_5988,N_5151,N_5178);
nor U5989 (N_5989,N_5417,N_5328);
nand U5990 (N_5990,N_5007,N_5359);
xor U5991 (N_5991,N_5381,N_5482);
or U5992 (N_5992,N_5065,N_5206);
nand U5993 (N_5993,N_5437,N_5162);
xor U5994 (N_5994,N_5167,N_5181);
and U5995 (N_5995,N_5117,N_5001);
nand U5996 (N_5996,N_5416,N_5177);
xor U5997 (N_5997,N_5040,N_5264);
or U5998 (N_5998,N_5478,N_5472);
nand U5999 (N_5999,N_5428,N_5133);
nor U6000 (N_6000,N_5539,N_5594);
and U6001 (N_6001,N_5642,N_5981);
nand U6002 (N_6002,N_5752,N_5927);
nand U6003 (N_6003,N_5734,N_5649);
nor U6004 (N_6004,N_5794,N_5588);
or U6005 (N_6005,N_5589,N_5839);
nand U6006 (N_6006,N_5658,N_5540);
xor U6007 (N_6007,N_5703,N_5699);
nand U6008 (N_6008,N_5747,N_5807);
and U6009 (N_6009,N_5942,N_5898);
or U6010 (N_6010,N_5505,N_5951);
nand U6011 (N_6011,N_5680,N_5726);
nand U6012 (N_6012,N_5862,N_5626);
and U6013 (N_6013,N_5965,N_5834);
nor U6014 (N_6014,N_5549,N_5547);
nor U6015 (N_6015,N_5619,N_5556);
nor U6016 (N_6016,N_5976,N_5673);
and U6017 (N_6017,N_5706,N_5688);
nor U6018 (N_6018,N_5584,N_5801);
or U6019 (N_6019,N_5859,N_5596);
and U6020 (N_6020,N_5779,N_5676);
xor U6021 (N_6021,N_5691,N_5892);
xnor U6022 (N_6022,N_5756,N_5795);
or U6023 (N_6023,N_5724,N_5929);
nor U6024 (N_6024,N_5915,N_5617);
xnor U6025 (N_6025,N_5534,N_5879);
nand U6026 (N_6026,N_5887,N_5907);
nand U6027 (N_6027,N_5912,N_5525);
nand U6028 (N_6028,N_5854,N_5620);
nor U6029 (N_6029,N_5817,N_5911);
nor U6030 (N_6030,N_5868,N_5704);
nor U6031 (N_6031,N_5624,N_5934);
nand U6032 (N_6032,N_5733,N_5906);
or U6033 (N_6033,N_5785,N_5622);
nor U6034 (N_6034,N_5996,N_5857);
xor U6035 (N_6035,N_5994,N_5742);
and U6036 (N_6036,N_5806,N_5618);
or U6037 (N_6037,N_5820,N_5761);
or U6038 (N_6038,N_5708,N_5792);
and U6039 (N_6039,N_5998,N_5616);
xor U6040 (N_6040,N_5864,N_5844);
and U6041 (N_6041,N_5652,N_5836);
xor U6042 (N_6042,N_5579,N_5563);
nor U6043 (N_6043,N_5664,N_5861);
nand U6044 (N_6044,N_5827,N_5928);
nand U6045 (N_6045,N_5885,N_5790);
nor U6046 (N_6046,N_5926,N_5709);
xnor U6047 (N_6047,N_5608,N_5557);
xnor U6048 (N_6048,N_5808,N_5644);
and U6049 (N_6049,N_5908,N_5646);
or U6050 (N_6050,N_5787,N_5560);
nand U6051 (N_6051,N_5753,N_5871);
nor U6052 (N_6052,N_5848,N_5899);
and U6053 (N_6053,N_5901,N_5502);
nor U6054 (N_6054,N_5692,N_5975);
nand U6055 (N_6055,N_5886,N_5980);
nor U6056 (N_6056,N_5812,N_5741);
nor U6057 (N_6057,N_5973,N_5705);
nor U6058 (N_6058,N_5754,N_5865);
xor U6059 (N_6059,N_5972,N_5826);
xor U6060 (N_6060,N_5512,N_5968);
nor U6061 (N_6061,N_5755,N_5781);
or U6062 (N_6062,N_5774,N_5920);
nor U6063 (N_6063,N_5757,N_5598);
nand U6064 (N_6064,N_5894,N_5772);
nor U6065 (N_6065,N_5938,N_5610);
nor U6066 (N_6066,N_5648,N_5881);
or U6067 (N_6067,N_5650,N_5576);
or U6068 (N_6068,N_5611,N_5759);
xor U6069 (N_6069,N_5518,N_5668);
xnor U6070 (N_6070,N_5728,N_5986);
xnor U6071 (N_6071,N_5535,N_5717);
nor U6072 (N_6072,N_5590,N_5948);
or U6073 (N_6073,N_5985,N_5916);
and U6074 (N_6074,N_5918,N_5974);
nand U6075 (N_6075,N_5701,N_5566);
xor U6076 (N_6076,N_5883,N_5950);
and U6077 (N_6077,N_5647,N_5758);
or U6078 (N_6078,N_5609,N_5946);
nor U6079 (N_6079,N_5884,N_5874);
nor U6080 (N_6080,N_5803,N_5681);
nand U6081 (N_6081,N_5696,N_5570);
nand U6082 (N_6082,N_5878,N_5924);
and U6083 (N_6083,N_5635,N_5727);
nor U6084 (N_6084,N_5775,N_5822);
or U6085 (N_6085,N_5813,N_5506);
nor U6086 (N_6086,N_5777,N_5569);
xnor U6087 (N_6087,N_5613,N_5583);
nand U6088 (N_6088,N_5850,N_5532);
and U6089 (N_6089,N_5625,N_5670);
nand U6090 (N_6090,N_5723,N_5627);
nor U6091 (N_6091,N_5931,N_5846);
nor U6092 (N_6092,N_5716,N_5645);
and U6093 (N_6093,N_5640,N_5592);
nand U6094 (N_6094,N_5623,N_5661);
and U6095 (N_6095,N_5783,N_5678);
nand U6096 (N_6096,N_5815,N_5538);
nand U6097 (N_6097,N_5914,N_5863);
and U6098 (N_6098,N_5621,N_5930);
nand U6099 (N_6099,N_5529,N_5963);
xnor U6100 (N_6100,N_5541,N_5572);
and U6101 (N_6101,N_5653,N_5749);
or U6102 (N_6102,N_5612,N_5721);
nand U6103 (N_6103,N_5903,N_5764);
nand U6104 (N_6104,N_5891,N_5511);
xor U6105 (N_6105,N_5939,N_5900);
nand U6106 (N_6106,N_5677,N_5660);
xor U6107 (N_6107,N_5551,N_5768);
and U6108 (N_6108,N_5888,N_5545);
nor U6109 (N_6109,N_5604,N_5933);
xnor U6110 (N_6110,N_5543,N_5542);
or U6111 (N_6111,N_5987,N_5970);
and U6112 (N_6112,N_5770,N_5521);
nand U6113 (N_6113,N_5687,N_5568);
nor U6114 (N_6114,N_5639,N_5513);
nand U6115 (N_6115,N_5776,N_5530);
or U6116 (N_6116,N_5956,N_5867);
or U6117 (N_6117,N_5936,N_5905);
xor U6118 (N_6118,N_5830,N_5841);
and U6119 (N_6119,N_5837,N_5522);
xor U6120 (N_6120,N_5913,N_5607);
xor U6121 (N_6121,N_5595,N_5602);
xnor U6122 (N_6122,N_5791,N_5880);
nor U6123 (N_6123,N_5788,N_5944);
xnor U6124 (N_6124,N_5597,N_5665);
nor U6125 (N_6125,N_5722,N_5711);
and U6126 (N_6126,N_5707,N_5809);
nor U6127 (N_6127,N_5860,N_5760);
nand U6128 (N_6128,N_5831,N_5666);
and U6129 (N_6129,N_5869,N_5955);
nor U6130 (N_6130,N_5667,N_5750);
or U6131 (N_6131,N_5958,N_5698);
nand U6132 (N_6132,N_5737,N_5577);
and U6133 (N_6133,N_5751,N_5524);
nor U6134 (N_6134,N_5743,N_5531);
xnor U6135 (N_6135,N_5634,N_5585);
nor U6136 (N_6136,N_5997,N_5546);
or U6137 (N_6137,N_5840,N_5810);
xor U6138 (N_6138,N_5636,N_5957);
or U6139 (N_6139,N_5565,N_5533);
and U6140 (N_6140,N_5700,N_5941);
xnor U6141 (N_6141,N_5519,N_5605);
xor U6142 (N_6142,N_5904,N_5744);
xor U6143 (N_6143,N_5993,N_5954);
xor U6144 (N_6144,N_5895,N_5897);
or U6145 (N_6145,N_5952,N_5537);
or U6146 (N_6146,N_5849,N_5919);
xor U6147 (N_6147,N_5989,N_5995);
xnor U6148 (N_6148,N_5659,N_5990);
or U6149 (N_6149,N_5953,N_5714);
and U6150 (N_6150,N_5674,N_5890);
xnor U6151 (N_6151,N_5715,N_5977);
and U6152 (N_6152,N_5567,N_5882);
nand U6153 (N_6153,N_5838,N_5988);
xnor U6154 (N_6154,N_5949,N_5835);
or U6155 (N_6155,N_5935,N_5638);
xor U6156 (N_6156,N_5654,N_5571);
nor U6157 (N_6157,N_5922,N_5765);
xor U6158 (N_6158,N_5829,N_5599);
and U6159 (N_6159,N_5961,N_5690);
xnor U6160 (N_6160,N_5999,N_5964);
xor U6161 (N_6161,N_5694,N_5784);
xnor U6162 (N_6162,N_5960,N_5866);
and U6163 (N_6163,N_5693,N_5702);
nand U6164 (N_6164,N_5771,N_5876);
nand U6165 (N_6165,N_5889,N_5739);
xnor U6166 (N_6166,N_5695,N_5766);
nand U6167 (N_6167,N_5982,N_5736);
nand U6168 (N_6168,N_5713,N_5656);
nand U6169 (N_6169,N_5762,N_5798);
xor U6170 (N_6170,N_5655,N_5679);
and U6171 (N_6171,N_5503,N_5730);
nand U6172 (N_6172,N_5923,N_5821);
and U6173 (N_6173,N_5548,N_5828);
nor U6174 (N_6174,N_5526,N_5552);
xnor U6175 (N_6175,N_5553,N_5501);
xnor U6176 (N_6176,N_5991,N_5825);
and U6177 (N_6177,N_5824,N_5735);
and U6178 (N_6178,N_5561,N_5978);
and U6179 (N_6179,N_5629,N_5797);
and U6180 (N_6180,N_5818,N_5558);
nor U6181 (N_6181,N_5651,N_5685);
or U6182 (N_6182,N_5575,N_5528);
nand U6183 (N_6183,N_5962,N_5778);
and U6184 (N_6184,N_5729,N_5940);
nor U6185 (N_6185,N_5921,N_5718);
nor U6186 (N_6186,N_5580,N_5740);
nor U6187 (N_6187,N_5591,N_5870);
and U6188 (N_6188,N_5581,N_5966);
or U6189 (N_6189,N_5632,N_5682);
and U6190 (N_6190,N_5833,N_5637);
and U6191 (N_6191,N_5536,N_5748);
and U6192 (N_6192,N_5793,N_5816);
and U6193 (N_6193,N_5507,N_5802);
xnor U6194 (N_6194,N_5631,N_5773);
and U6195 (N_6195,N_5814,N_5767);
and U6196 (N_6196,N_5663,N_5855);
and U6197 (N_6197,N_5845,N_5712);
and U6198 (N_6198,N_5550,N_5804);
xnor U6199 (N_6199,N_5858,N_5710);
xor U6200 (N_6200,N_5601,N_5943);
nand U6201 (N_6201,N_5852,N_5947);
or U6202 (N_6202,N_5725,N_5983);
or U6203 (N_6203,N_5662,N_5800);
xor U6204 (N_6204,N_5600,N_5508);
xnor U6205 (N_6205,N_5945,N_5811);
and U6206 (N_6206,N_5877,N_5769);
and U6207 (N_6207,N_5843,N_5853);
xor U6208 (N_6208,N_5520,N_5516);
nand U6209 (N_6209,N_5875,N_5902);
nand U6210 (N_6210,N_5910,N_5669);
or U6211 (N_6211,N_5925,N_5562);
nand U6212 (N_6212,N_5805,N_5932);
and U6213 (N_6213,N_5657,N_5582);
nor U6214 (N_6214,N_5633,N_5745);
xnor U6215 (N_6215,N_5504,N_5893);
or U6216 (N_6216,N_5510,N_5683);
or U6217 (N_6217,N_5523,N_5896);
nor U6218 (N_6218,N_5917,N_5782);
nor U6219 (N_6219,N_5780,N_5672);
or U6220 (N_6220,N_5832,N_5971);
or U6221 (N_6221,N_5689,N_5732);
or U6222 (N_6222,N_5675,N_5628);
or U6223 (N_6223,N_5796,N_5979);
nand U6224 (N_6224,N_5641,N_5719);
nor U6225 (N_6225,N_5555,N_5574);
nor U6226 (N_6226,N_5564,N_5614);
nand U6227 (N_6227,N_5873,N_5799);
nand U6228 (N_6228,N_5514,N_5544);
or U6229 (N_6229,N_5587,N_5603);
nand U6230 (N_6230,N_5559,N_5738);
and U6231 (N_6231,N_5527,N_5643);
and U6232 (N_6232,N_5856,N_5517);
or U6233 (N_6233,N_5686,N_5746);
nor U6234 (N_6234,N_5573,N_5554);
or U6235 (N_6235,N_5763,N_5909);
or U6236 (N_6236,N_5842,N_5509);
or U6237 (N_6237,N_5789,N_5586);
xor U6238 (N_6238,N_5937,N_5823);
or U6239 (N_6239,N_5615,N_5515);
xnor U6240 (N_6240,N_5671,N_5851);
nor U6241 (N_6241,N_5819,N_5967);
nor U6242 (N_6242,N_5992,N_5731);
xor U6243 (N_6243,N_5500,N_5720);
xnor U6244 (N_6244,N_5697,N_5606);
nor U6245 (N_6245,N_5593,N_5786);
nor U6246 (N_6246,N_5578,N_5684);
and U6247 (N_6247,N_5984,N_5969);
and U6248 (N_6248,N_5630,N_5872);
nand U6249 (N_6249,N_5847,N_5959);
xnor U6250 (N_6250,N_5591,N_5571);
and U6251 (N_6251,N_5997,N_5860);
nor U6252 (N_6252,N_5976,N_5721);
and U6253 (N_6253,N_5592,N_5630);
nand U6254 (N_6254,N_5998,N_5584);
and U6255 (N_6255,N_5937,N_5503);
or U6256 (N_6256,N_5994,N_5753);
xnor U6257 (N_6257,N_5624,N_5693);
nor U6258 (N_6258,N_5592,N_5609);
or U6259 (N_6259,N_5934,N_5897);
xor U6260 (N_6260,N_5530,N_5945);
and U6261 (N_6261,N_5938,N_5698);
nand U6262 (N_6262,N_5540,N_5556);
or U6263 (N_6263,N_5505,N_5887);
nand U6264 (N_6264,N_5812,N_5822);
or U6265 (N_6265,N_5983,N_5839);
and U6266 (N_6266,N_5856,N_5871);
nor U6267 (N_6267,N_5513,N_5940);
and U6268 (N_6268,N_5895,N_5755);
xor U6269 (N_6269,N_5698,N_5795);
xor U6270 (N_6270,N_5964,N_5671);
and U6271 (N_6271,N_5510,N_5886);
nor U6272 (N_6272,N_5546,N_5661);
xor U6273 (N_6273,N_5584,N_5503);
nand U6274 (N_6274,N_5703,N_5795);
nor U6275 (N_6275,N_5633,N_5605);
nor U6276 (N_6276,N_5853,N_5718);
nor U6277 (N_6277,N_5568,N_5999);
or U6278 (N_6278,N_5634,N_5842);
nand U6279 (N_6279,N_5587,N_5845);
nand U6280 (N_6280,N_5823,N_5810);
or U6281 (N_6281,N_5817,N_5520);
xor U6282 (N_6282,N_5994,N_5637);
nand U6283 (N_6283,N_5555,N_5626);
nor U6284 (N_6284,N_5912,N_5910);
nand U6285 (N_6285,N_5830,N_5506);
and U6286 (N_6286,N_5898,N_5582);
or U6287 (N_6287,N_5941,N_5863);
or U6288 (N_6288,N_5659,N_5930);
and U6289 (N_6289,N_5679,N_5736);
nand U6290 (N_6290,N_5736,N_5770);
xnor U6291 (N_6291,N_5739,N_5878);
or U6292 (N_6292,N_5580,N_5590);
nor U6293 (N_6293,N_5984,N_5791);
and U6294 (N_6294,N_5703,N_5875);
xor U6295 (N_6295,N_5976,N_5975);
nor U6296 (N_6296,N_5633,N_5971);
and U6297 (N_6297,N_5840,N_5877);
xnor U6298 (N_6298,N_5771,N_5849);
xor U6299 (N_6299,N_5824,N_5566);
xor U6300 (N_6300,N_5636,N_5728);
xor U6301 (N_6301,N_5940,N_5928);
and U6302 (N_6302,N_5538,N_5891);
nor U6303 (N_6303,N_5676,N_5876);
and U6304 (N_6304,N_5872,N_5851);
and U6305 (N_6305,N_5766,N_5526);
and U6306 (N_6306,N_5910,N_5594);
nand U6307 (N_6307,N_5980,N_5650);
xnor U6308 (N_6308,N_5594,N_5804);
xnor U6309 (N_6309,N_5560,N_5786);
nand U6310 (N_6310,N_5576,N_5951);
nor U6311 (N_6311,N_5539,N_5798);
xor U6312 (N_6312,N_5581,N_5727);
nor U6313 (N_6313,N_5511,N_5786);
nor U6314 (N_6314,N_5811,N_5594);
or U6315 (N_6315,N_5737,N_5932);
and U6316 (N_6316,N_5673,N_5935);
or U6317 (N_6317,N_5975,N_5703);
and U6318 (N_6318,N_5658,N_5857);
and U6319 (N_6319,N_5601,N_5969);
nor U6320 (N_6320,N_5753,N_5890);
or U6321 (N_6321,N_5917,N_5830);
or U6322 (N_6322,N_5718,N_5588);
and U6323 (N_6323,N_5674,N_5682);
nand U6324 (N_6324,N_5667,N_5907);
nand U6325 (N_6325,N_5631,N_5912);
and U6326 (N_6326,N_5985,N_5809);
nor U6327 (N_6327,N_5779,N_5617);
xor U6328 (N_6328,N_5784,N_5940);
xor U6329 (N_6329,N_5971,N_5864);
nand U6330 (N_6330,N_5812,N_5915);
nand U6331 (N_6331,N_5619,N_5600);
xnor U6332 (N_6332,N_5979,N_5964);
nor U6333 (N_6333,N_5906,N_5625);
or U6334 (N_6334,N_5847,N_5611);
nor U6335 (N_6335,N_5803,N_5696);
xor U6336 (N_6336,N_5948,N_5695);
or U6337 (N_6337,N_5864,N_5827);
and U6338 (N_6338,N_5989,N_5609);
xnor U6339 (N_6339,N_5634,N_5521);
xnor U6340 (N_6340,N_5687,N_5811);
nor U6341 (N_6341,N_5752,N_5551);
nand U6342 (N_6342,N_5975,N_5606);
xnor U6343 (N_6343,N_5659,N_5785);
xnor U6344 (N_6344,N_5658,N_5849);
nand U6345 (N_6345,N_5719,N_5825);
xnor U6346 (N_6346,N_5572,N_5640);
and U6347 (N_6347,N_5654,N_5721);
xor U6348 (N_6348,N_5572,N_5729);
xnor U6349 (N_6349,N_5687,N_5755);
and U6350 (N_6350,N_5873,N_5576);
or U6351 (N_6351,N_5798,N_5977);
xor U6352 (N_6352,N_5511,N_5904);
xnor U6353 (N_6353,N_5902,N_5572);
or U6354 (N_6354,N_5649,N_5678);
and U6355 (N_6355,N_5768,N_5576);
or U6356 (N_6356,N_5644,N_5567);
xor U6357 (N_6357,N_5896,N_5996);
or U6358 (N_6358,N_5518,N_5810);
nand U6359 (N_6359,N_5794,N_5803);
nand U6360 (N_6360,N_5889,N_5718);
nand U6361 (N_6361,N_5944,N_5751);
and U6362 (N_6362,N_5993,N_5530);
nand U6363 (N_6363,N_5613,N_5930);
nand U6364 (N_6364,N_5567,N_5611);
nor U6365 (N_6365,N_5753,N_5855);
nand U6366 (N_6366,N_5804,N_5693);
nor U6367 (N_6367,N_5809,N_5950);
xnor U6368 (N_6368,N_5947,N_5911);
xor U6369 (N_6369,N_5597,N_5593);
and U6370 (N_6370,N_5655,N_5941);
or U6371 (N_6371,N_5656,N_5980);
or U6372 (N_6372,N_5617,N_5935);
and U6373 (N_6373,N_5830,N_5984);
nand U6374 (N_6374,N_5932,N_5626);
xor U6375 (N_6375,N_5554,N_5848);
xor U6376 (N_6376,N_5517,N_5996);
xor U6377 (N_6377,N_5628,N_5882);
or U6378 (N_6378,N_5922,N_5612);
nand U6379 (N_6379,N_5968,N_5815);
nand U6380 (N_6380,N_5536,N_5932);
nor U6381 (N_6381,N_5808,N_5714);
nand U6382 (N_6382,N_5806,N_5551);
and U6383 (N_6383,N_5597,N_5799);
xor U6384 (N_6384,N_5803,N_5624);
nand U6385 (N_6385,N_5592,N_5551);
nor U6386 (N_6386,N_5517,N_5510);
xnor U6387 (N_6387,N_5552,N_5754);
nor U6388 (N_6388,N_5534,N_5565);
and U6389 (N_6389,N_5798,N_5783);
xor U6390 (N_6390,N_5671,N_5630);
nand U6391 (N_6391,N_5713,N_5710);
and U6392 (N_6392,N_5739,N_5602);
nor U6393 (N_6393,N_5686,N_5843);
nor U6394 (N_6394,N_5741,N_5515);
nand U6395 (N_6395,N_5795,N_5808);
and U6396 (N_6396,N_5587,N_5984);
or U6397 (N_6397,N_5501,N_5932);
nor U6398 (N_6398,N_5740,N_5915);
or U6399 (N_6399,N_5768,N_5950);
nor U6400 (N_6400,N_5615,N_5760);
nand U6401 (N_6401,N_5656,N_5852);
or U6402 (N_6402,N_5976,N_5926);
and U6403 (N_6403,N_5575,N_5555);
or U6404 (N_6404,N_5796,N_5716);
nor U6405 (N_6405,N_5528,N_5678);
and U6406 (N_6406,N_5642,N_5878);
or U6407 (N_6407,N_5592,N_5683);
nand U6408 (N_6408,N_5572,N_5955);
or U6409 (N_6409,N_5697,N_5940);
xor U6410 (N_6410,N_5727,N_5905);
nand U6411 (N_6411,N_5915,N_5693);
or U6412 (N_6412,N_5705,N_5877);
nor U6413 (N_6413,N_5708,N_5848);
nor U6414 (N_6414,N_5993,N_5686);
or U6415 (N_6415,N_5509,N_5803);
nor U6416 (N_6416,N_5524,N_5874);
nand U6417 (N_6417,N_5586,N_5660);
xor U6418 (N_6418,N_5505,N_5868);
and U6419 (N_6419,N_5944,N_5614);
or U6420 (N_6420,N_5589,N_5614);
nor U6421 (N_6421,N_5657,N_5649);
or U6422 (N_6422,N_5525,N_5682);
nand U6423 (N_6423,N_5549,N_5683);
nand U6424 (N_6424,N_5629,N_5596);
nor U6425 (N_6425,N_5748,N_5729);
nand U6426 (N_6426,N_5508,N_5648);
or U6427 (N_6427,N_5733,N_5624);
or U6428 (N_6428,N_5539,N_5986);
or U6429 (N_6429,N_5996,N_5974);
and U6430 (N_6430,N_5680,N_5798);
nor U6431 (N_6431,N_5684,N_5825);
or U6432 (N_6432,N_5732,N_5766);
xor U6433 (N_6433,N_5984,N_5893);
nor U6434 (N_6434,N_5508,N_5727);
nand U6435 (N_6435,N_5522,N_5601);
nor U6436 (N_6436,N_5842,N_5998);
nand U6437 (N_6437,N_5583,N_5770);
and U6438 (N_6438,N_5847,N_5967);
nor U6439 (N_6439,N_5619,N_5854);
nor U6440 (N_6440,N_5919,N_5787);
nor U6441 (N_6441,N_5965,N_5516);
nor U6442 (N_6442,N_5567,N_5847);
nand U6443 (N_6443,N_5957,N_5972);
and U6444 (N_6444,N_5690,N_5782);
and U6445 (N_6445,N_5649,N_5993);
nor U6446 (N_6446,N_5769,N_5536);
nor U6447 (N_6447,N_5606,N_5736);
or U6448 (N_6448,N_5850,N_5692);
nor U6449 (N_6449,N_5709,N_5802);
or U6450 (N_6450,N_5854,N_5922);
and U6451 (N_6451,N_5970,N_5673);
nor U6452 (N_6452,N_5728,N_5547);
nand U6453 (N_6453,N_5875,N_5590);
nand U6454 (N_6454,N_5553,N_5911);
or U6455 (N_6455,N_5820,N_5799);
nor U6456 (N_6456,N_5540,N_5747);
nand U6457 (N_6457,N_5527,N_5759);
xor U6458 (N_6458,N_5956,N_5621);
nor U6459 (N_6459,N_5947,N_5973);
and U6460 (N_6460,N_5570,N_5547);
nand U6461 (N_6461,N_5533,N_5982);
nand U6462 (N_6462,N_5605,N_5557);
and U6463 (N_6463,N_5974,N_5624);
or U6464 (N_6464,N_5656,N_5720);
xnor U6465 (N_6465,N_5517,N_5559);
and U6466 (N_6466,N_5707,N_5841);
xor U6467 (N_6467,N_5828,N_5556);
xnor U6468 (N_6468,N_5602,N_5624);
or U6469 (N_6469,N_5734,N_5622);
nand U6470 (N_6470,N_5699,N_5841);
or U6471 (N_6471,N_5764,N_5929);
xnor U6472 (N_6472,N_5645,N_5636);
or U6473 (N_6473,N_5948,N_5605);
xnor U6474 (N_6474,N_5852,N_5606);
and U6475 (N_6475,N_5765,N_5842);
and U6476 (N_6476,N_5558,N_5715);
nor U6477 (N_6477,N_5750,N_5650);
and U6478 (N_6478,N_5900,N_5805);
nor U6479 (N_6479,N_5739,N_5644);
or U6480 (N_6480,N_5952,N_5654);
nand U6481 (N_6481,N_5565,N_5919);
and U6482 (N_6482,N_5906,N_5945);
xnor U6483 (N_6483,N_5537,N_5832);
nor U6484 (N_6484,N_5549,N_5765);
or U6485 (N_6485,N_5632,N_5716);
or U6486 (N_6486,N_5673,N_5572);
xnor U6487 (N_6487,N_5966,N_5905);
and U6488 (N_6488,N_5535,N_5679);
or U6489 (N_6489,N_5706,N_5940);
and U6490 (N_6490,N_5711,N_5798);
nand U6491 (N_6491,N_5540,N_5867);
or U6492 (N_6492,N_5694,N_5723);
xor U6493 (N_6493,N_5937,N_5854);
or U6494 (N_6494,N_5571,N_5831);
or U6495 (N_6495,N_5937,N_5668);
and U6496 (N_6496,N_5648,N_5603);
nor U6497 (N_6497,N_5504,N_5656);
xnor U6498 (N_6498,N_5602,N_5648);
or U6499 (N_6499,N_5615,N_5981);
nand U6500 (N_6500,N_6330,N_6159);
and U6501 (N_6501,N_6471,N_6056);
or U6502 (N_6502,N_6388,N_6078);
and U6503 (N_6503,N_6194,N_6331);
xnor U6504 (N_6504,N_6235,N_6303);
and U6505 (N_6505,N_6483,N_6404);
nand U6506 (N_6506,N_6354,N_6366);
or U6507 (N_6507,N_6424,N_6148);
nor U6508 (N_6508,N_6131,N_6048);
nor U6509 (N_6509,N_6248,N_6410);
or U6510 (N_6510,N_6461,N_6152);
nand U6511 (N_6511,N_6329,N_6000);
or U6512 (N_6512,N_6326,N_6193);
xnor U6513 (N_6513,N_6263,N_6072);
xor U6514 (N_6514,N_6157,N_6151);
nor U6515 (N_6515,N_6055,N_6239);
xnor U6516 (N_6516,N_6062,N_6409);
nor U6517 (N_6517,N_6422,N_6381);
xor U6518 (N_6518,N_6003,N_6024);
nor U6519 (N_6519,N_6082,N_6467);
and U6520 (N_6520,N_6480,N_6423);
xnor U6521 (N_6521,N_6445,N_6380);
or U6522 (N_6522,N_6304,N_6237);
nor U6523 (N_6523,N_6134,N_6198);
nand U6524 (N_6524,N_6034,N_6027);
nand U6525 (N_6525,N_6324,N_6188);
nand U6526 (N_6526,N_6236,N_6207);
nor U6527 (N_6527,N_6013,N_6323);
nand U6528 (N_6528,N_6438,N_6083);
and U6529 (N_6529,N_6120,N_6377);
or U6530 (N_6530,N_6183,N_6214);
nor U6531 (N_6531,N_6349,N_6232);
nand U6532 (N_6532,N_6124,N_6096);
nand U6533 (N_6533,N_6099,N_6125);
or U6534 (N_6534,N_6435,N_6311);
xor U6535 (N_6535,N_6308,N_6261);
nand U6536 (N_6536,N_6250,N_6032);
nor U6537 (N_6537,N_6167,N_6118);
nand U6538 (N_6538,N_6455,N_6184);
nor U6539 (N_6539,N_6243,N_6314);
and U6540 (N_6540,N_6446,N_6029);
and U6541 (N_6541,N_6249,N_6337);
and U6542 (N_6542,N_6466,N_6498);
and U6543 (N_6543,N_6154,N_6225);
nor U6544 (N_6544,N_6357,N_6020);
xor U6545 (N_6545,N_6475,N_6028);
nor U6546 (N_6546,N_6174,N_6278);
and U6547 (N_6547,N_6292,N_6295);
and U6548 (N_6548,N_6320,N_6169);
nand U6549 (N_6549,N_6402,N_6224);
and U6550 (N_6550,N_6210,N_6037);
nor U6551 (N_6551,N_6453,N_6310);
or U6552 (N_6552,N_6177,N_6080);
and U6553 (N_6553,N_6254,N_6156);
xor U6554 (N_6554,N_6244,N_6265);
nor U6555 (N_6555,N_6077,N_6274);
or U6556 (N_6556,N_6367,N_6260);
nand U6557 (N_6557,N_6021,N_6211);
nand U6558 (N_6558,N_6073,N_6421);
or U6559 (N_6559,N_6428,N_6222);
xnor U6560 (N_6560,N_6081,N_6494);
or U6561 (N_6561,N_6065,N_6439);
nand U6562 (N_6562,N_6229,N_6089);
xnor U6563 (N_6563,N_6299,N_6040);
nand U6564 (N_6564,N_6164,N_6012);
and U6565 (N_6565,N_6087,N_6086);
xor U6566 (N_6566,N_6001,N_6362);
xor U6567 (N_6567,N_6495,N_6440);
nor U6568 (N_6568,N_6059,N_6142);
nor U6569 (N_6569,N_6473,N_6117);
nand U6570 (N_6570,N_6202,N_6327);
nand U6571 (N_6571,N_6460,N_6312);
nor U6572 (N_6572,N_6420,N_6288);
or U6573 (N_6573,N_6178,N_6487);
nor U6574 (N_6574,N_6146,N_6352);
and U6575 (N_6575,N_6479,N_6060);
nor U6576 (N_6576,N_6196,N_6114);
xor U6577 (N_6577,N_6465,N_6341);
or U6578 (N_6578,N_6205,N_6140);
nor U6579 (N_6579,N_6245,N_6429);
nor U6580 (N_6580,N_6128,N_6338);
or U6581 (N_6581,N_6328,N_6301);
or U6582 (N_6582,N_6256,N_6348);
xnor U6583 (N_6583,N_6126,N_6259);
xnor U6584 (N_6584,N_6302,N_6097);
or U6585 (N_6585,N_6276,N_6147);
nor U6586 (N_6586,N_6300,N_6436);
xnor U6587 (N_6587,N_6216,N_6233);
and U6588 (N_6588,N_6345,N_6332);
nor U6589 (N_6589,N_6297,N_6171);
xor U6590 (N_6590,N_6155,N_6355);
or U6591 (N_6591,N_6234,N_6018);
and U6592 (N_6592,N_6092,N_6127);
and U6593 (N_6593,N_6286,N_6283);
xnor U6594 (N_6594,N_6005,N_6291);
nor U6595 (N_6595,N_6135,N_6163);
or U6596 (N_6596,N_6449,N_6411);
nor U6597 (N_6597,N_6110,N_6069);
xnor U6598 (N_6598,N_6206,N_6113);
nor U6599 (N_6599,N_6353,N_6294);
xor U6600 (N_6600,N_6342,N_6387);
or U6601 (N_6601,N_6363,N_6122);
and U6602 (N_6602,N_6384,N_6419);
and U6603 (N_6603,N_6149,N_6334);
nand U6604 (N_6604,N_6144,N_6053);
or U6605 (N_6605,N_6186,N_6153);
and U6606 (N_6606,N_6112,N_6485);
or U6607 (N_6607,N_6322,N_6185);
or U6608 (N_6608,N_6133,N_6270);
xor U6609 (N_6609,N_6488,N_6165);
nand U6610 (N_6610,N_6390,N_6346);
or U6611 (N_6611,N_6022,N_6405);
nor U6612 (N_6612,N_6090,N_6042);
or U6613 (N_6613,N_6437,N_6463);
nor U6614 (N_6614,N_6431,N_6006);
or U6615 (N_6615,N_6425,N_6396);
nor U6616 (N_6616,N_6102,N_6212);
xor U6617 (N_6617,N_6187,N_6158);
nor U6618 (N_6618,N_6373,N_6279);
and U6619 (N_6619,N_6298,N_6452);
nand U6620 (N_6620,N_6103,N_6190);
xnor U6621 (N_6621,N_6030,N_6019);
nand U6622 (N_6622,N_6317,N_6319);
and U6623 (N_6623,N_6038,N_6119);
and U6624 (N_6624,N_6010,N_6365);
and U6625 (N_6625,N_6192,N_6079);
nand U6626 (N_6626,N_6025,N_6258);
xnor U6627 (N_6627,N_6486,N_6277);
xnor U6628 (N_6628,N_6189,N_6071);
xor U6629 (N_6629,N_6011,N_6255);
or U6630 (N_6630,N_6014,N_6307);
and U6631 (N_6631,N_6238,N_6015);
xor U6632 (N_6632,N_6393,N_6172);
nand U6633 (N_6633,N_6161,N_6399);
or U6634 (N_6634,N_6371,N_6374);
xor U6635 (N_6635,N_6061,N_6418);
nor U6636 (N_6636,N_6477,N_6182);
and U6637 (N_6637,N_6413,N_6378);
nand U6638 (N_6638,N_6379,N_6284);
nor U6639 (N_6639,N_6444,N_6457);
or U6640 (N_6640,N_6344,N_6442);
xor U6641 (N_6641,N_6497,N_6271);
xor U6642 (N_6642,N_6252,N_6215);
nor U6643 (N_6643,N_6228,N_6336);
xor U6644 (N_6644,N_6383,N_6335);
nor U6645 (N_6645,N_6241,N_6407);
or U6646 (N_6646,N_6166,N_6121);
or U6647 (N_6647,N_6068,N_6031);
and U6648 (N_6648,N_6458,N_6051);
and U6649 (N_6649,N_6004,N_6339);
xor U6650 (N_6650,N_6039,N_6430);
and U6651 (N_6651,N_6052,N_6076);
or U6652 (N_6652,N_6070,N_6191);
and U6653 (N_6653,N_6492,N_6347);
nor U6654 (N_6654,N_6100,N_6231);
nand U6655 (N_6655,N_6451,N_6476);
xnor U6656 (N_6656,N_6478,N_6035);
or U6657 (N_6657,N_6129,N_6481);
and U6658 (N_6658,N_6287,N_6054);
xnor U6659 (N_6659,N_6414,N_6257);
nand U6660 (N_6660,N_6408,N_6130);
xor U6661 (N_6661,N_6240,N_6468);
or U6662 (N_6662,N_6143,N_6281);
nor U6663 (N_6663,N_6176,N_6496);
nor U6664 (N_6664,N_6098,N_6204);
nand U6665 (N_6665,N_6085,N_6470);
nand U6666 (N_6666,N_6401,N_6115);
and U6667 (N_6667,N_6104,N_6391);
and U6668 (N_6668,N_6201,N_6358);
nand U6669 (N_6669,N_6067,N_6064);
nor U6670 (N_6670,N_6008,N_6325);
nand U6671 (N_6671,N_6385,N_6179);
nor U6672 (N_6672,N_6262,N_6200);
nor U6673 (N_6673,N_6269,N_6441);
nand U6674 (N_6674,N_6023,N_6175);
xor U6675 (N_6675,N_6017,N_6199);
nand U6676 (N_6676,N_6219,N_6246);
and U6677 (N_6677,N_6482,N_6181);
xnor U6678 (N_6678,N_6132,N_6046);
nand U6679 (N_6679,N_6321,N_6221);
or U6680 (N_6680,N_6168,N_6406);
nand U6681 (N_6681,N_6375,N_6180);
or U6682 (N_6682,N_6462,N_6432);
and U6683 (N_6683,N_6472,N_6305);
xnor U6684 (N_6684,N_6107,N_6111);
or U6685 (N_6685,N_6002,N_6369);
or U6686 (N_6686,N_6106,N_6386);
nand U6687 (N_6687,N_6108,N_6091);
or U6688 (N_6688,N_6370,N_6218);
xor U6689 (N_6689,N_6109,N_6397);
or U6690 (N_6690,N_6266,N_6036);
xor U6691 (N_6691,N_6251,N_6289);
and U6692 (N_6692,N_6203,N_6490);
xnor U6693 (N_6693,N_6075,N_6350);
nor U6694 (N_6694,N_6415,N_6427);
nor U6695 (N_6695,N_6491,N_6093);
and U6696 (N_6696,N_6450,N_6309);
nand U6697 (N_6697,N_6223,N_6434);
and U6698 (N_6698,N_6376,N_6045);
nand U6699 (N_6699,N_6489,N_6137);
nand U6700 (N_6700,N_6273,N_6058);
nor U6701 (N_6701,N_6416,N_6084);
nor U6702 (N_6702,N_6459,N_6041);
and U6703 (N_6703,N_6316,N_6499);
or U6704 (N_6704,N_6394,N_6464);
xnor U6705 (N_6705,N_6293,N_6290);
nand U6706 (N_6706,N_6275,N_6368);
xnor U6707 (N_6707,N_6116,N_6443);
nand U6708 (N_6708,N_6026,N_6095);
nand U6709 (N_6709,N_6433,N_6389);
and U6710 (N_6710,N_6050,N_6264);
and U6711 (N_6711,N_6209,N_6139);
nand U6712 (N_6712,N_6138,N_6094);
nand U6713 (N_6713,N_6484,N_6049);
nand U6714 (N_6714,N_6474,N_6063);
nor U6715 (N_6715,N_6066,N_6173);
and U6716 (N_6716,N_6356,N_6306);
nand U6717 (N_6717,N_6282,N_6469);
xor U6718 (N_6718,N_6412,N_6247);
nor U6719 (N_6719,N_6101,N_6007);
or U6720 (N_6720,N_6047,N_6242);
nand U6721 (N_6721,N_6296,N_6145);
and U6722 (N_6722,N_6313,N_6398);
xnor U6723 (N_6723,N_6272,N_6088);
nor U6724 (N_6724,N_6403,N_6267);
nor U6725 (N_6725,N_6340,N_6136);
nor U6726 (N_6726,N_6454,N_6493);
nand U6727 (N_6727,N_6016,N_6057);
nor U6728 (N_6728,N_6456,N_6220);
xor U6729 (N_6729,N_6105,N_6364);
and U6730 (N_6730,N_6123,N_6285);
nand U6731 (N_6731,N_6360,N_6033);
nand U6732 (N_6732,N_6343,N_6141);
nand U6733 (N_6733,N_6253,N_6400);
xnor U6734 (N_6734,N_6226,N_6043);
nor U6735 (N_6735,N_6208,N_6009);
or U6736 (N_6736,N_6197,N_6227);
or U6737 (N_6737,N_6230,N_6213);
nor U6738 (N_6738,N_6195,N_6426);
nand U6739 (N_6739,N_6268,N_6044);
nor U6740 (N_6740,N_6333,N_6150);
xnor U6741 (N_6741,N_6395,N_6217);
xor U6742 (N_6742,N_6417,N_6162);
nand U6743 (N_6743,N_6361,N_6318);
xnor U6744 (N_6744,N_6372,N_6359);
or U6745 (N_6745,N_6382,N_6448);
nor U6746 (N_6746,N_6160,N_6315);
nor U6747 (N_6747,N_6074,N_6280);
xnor U6748 (N_6748,N_6351,N_6447);
xor U6749 (N_6749,N_6392,N_6170);
nor U6750 (N_6750,N_6070,N_6100);
or U6751 (N_6751,N_6235,N_6079);
xor U6752 (N_6752,N_6227,N_6361);
nand U6753 (N_6753,N_6162,N_6282);
nor U6754 (N_6754,N_6323,N_6314);
and U6755 (N_6755,N_6118,N_6002);
nand U6756 (N_6756,N_6017,N_6194);
or U6757 (N_6757,N_6442,N_6151);
or U6758 (N_6758,N_6278,N_6368);
or U6759 (N_6759,N_6484,N_6456);
and U6760 (N_6760,N_6193,N_6302);
and U6761 (N_6761,N_6462,N_6279);
nor U6762 (N_6762,N_6294,N_6477);
nor U6763 (N_6763,N_6237,N_6102);
nor U6764 (N_6764,N_6103,N_6251);
nand U6765 (N_6765,N_6005,N_6248);
or U6766 (N_6766,N_6438,N_6437);
xnor U6767 (N_6767,N_6223,N_6188);
nor U6768 (N_6768,N_6004,N_6436);
nand U6769 (N_6769,N_6050,N_6161);
or U6770 (N_6770,N_6288,N_6222);
nor U6771 (N_6771,N_6381,N_6031);
xnor U6772 (N_6772,N_6168,N_6007);
nor U6773 (N_6773,N_6005,N_6410);
nand U6774 (N_6774,N_6308,N_6051);
and U6775 (N_6775,N_6361,N_6255);
nor U6776 (N_6776,N_6303,N_6043);
or U6777 (N_6777,N_6253,N_6097);
nand U6778 (N_6778,N_6108,N_6454);
nor U6779 (N_6779,N_6278,N_6170);
or U6780 (N_6780,N_6075,N_6110);
nor U6781 (N_6781,N_6159,N_6048);
xor U6782 (N_6782,N_6191,N_6016);
and U6783 (N_6783,N_6089,N_6026);
nand U6784 (N_6784,N_6033,N_6131);
and U6785 (N_6785,N_6182,N_6311);
nand U6786 (N_6786,N_6102,N_6211);
xor U6787 (N_6787,N_6176,N_6100);
or U6788 (N_6788,N_6237,N_6480);
nand U6789 (N_6789,N_6325,N_6302);
nand U6790 (N_6790,N_6433,N_6141);
or U6791 (N_6791,N_6270,N_6278);
and U6792 (N_6792,N_6417,N_6020);
nand U6793 (N_6793,N_6153,N_6092);
nor U6794 (N_6794,N_6300,N_6378);
nand U6795 (N_6795,N_6460,N_6174);
xnor U6796 (N_6796,N_6436,N_6094);
or U6797 (N_6797,N_6394,N_6110);
nor U6798 (N_6798,N_6194,N_6243);
and U6799 (N_6799,N_6273,N_6002);
nor U6800 (N_6800,N_6439,N_6477);
xnor U6801 (N_6801,N_6134,N_6386);
and U6802 (N_6802,N_6471,N_6183);
nor U6803 (N_6803,N_6452,N_6411);
or U6804 (N_6804,N_6106,N_6227);
or U6805 (N_6805,N_6462,N_6292);
and U6806 (N_6806,N_6262,N_6171);
nor U6807 (N_6807,N_6353,N_6183);
nand U6808 (N_6808,N_6415,N_6044);
xnor U6809 (N_6809,N_6019,N_6423);
nand U6810 (N_6810,N_6380,N_6424);
or U6811 (N_6811,N_6196,N_6418);
and U6812 (N_6812,N_6307,N_6071);
or U6813 (N_6813,N_6238,N_6352);
nor U6814 (N_6814,N_6487,N_6308);
nor U6815 (N_6815,N_6023,N_6180);
xnor U6816 (N_6816,N_6111,N_6018);
nor U6817 (N_6817,N_6226,N_6197);
xnor U6818 (N_6818,N_6492,N_6482);
or U6819 (N_6819,N_6418,N_6170);
or U6820 (N_6820,N_6091,N_6463);
nor U6821 (N_6821,N_6100,N_6455);
or U6822 (N_6822,N_6405,N_6365);
nor U6823 (N_6823,N_6300,N_6457);
xnor U6824 (N_6824,N_6139,N_6159);
or U6825 (N_6825,N_6410,N_6192);
xor U6826 (N_6826,N_6058,N_6365);
and U6827 (N_6827,N_6142,N_6097);
and U6828 (N_6828,N_6359,N_6311);
and U6829 (N_6829,N_6243,N_6281);
or U6830 (N_6830,N_6358,N_6010);
or U6831 (N_6831,N_6492,N_6263);
nand U6832 (N_6832,N_6467,N_6167);
and U6833 (N_6833,N_6086,N_6083);
xnor U6834 (N_6834,N_6252,N_6017);
or U6835 (N_6835,N_6446,N_6249);
and U6836 (N_6836,N_6067,N_6301);
or U6837 (N_6837,N_6441,N_6312);
nand U6838 (N_6838,N_6240,N_6143);
and U6839 (N_6839,N_6157,N_6197);
xnor U6840 (N_6840,N_6222,N_6424);
nand U6841 (N_6841,N_6461,N_6438);
nand U6842 (N_6842,N_6052,N_6478);
or U6843 (N_6843,N_6462,N_6416);
nor U6844 (N_6844,N_6110,N_6440);
nand U6845 (N_6845,N_6335,N_6412);
nor U6846 (N_6846,N_6101,N_6237);
xnor U6847 (N_6847,N_6013,N_6122);
nor U6848 (N_6848,N_6088,N_6251);
and U6849 (N_6849,N_6380,N_6225);
nor U6850 (N_6850,N_6375,N_6024);
or U6851 (N_6851,N_6295,N_6408);
nor U6852 (N_6852,N_6282,N_6007);
nand U6853 (N_6853,N_6447,N_6378);
and U6854 (N_6854,N_6489,N_6076);
and U6855 (N_6855,N_6061,N_6330);
and U6856 (N_6856,N_6373,N_6292);
nand U6857 (N_6857,N_6035,N_6227);
nand U6858 (N_6858,N_6159,N_6333);
nand U6859 (N_6859,N_6441,N_6301);
and U6860 (N_6860,N_6267,N_6464);
xor U6861 (N_6861,N_6116,N_6391);
nand U6862 (N_6862,N_6256,N_6075);
or U6863 (N_6863,N_6158,N_6475);
nor U6864 (N_6864,N_6239,N_6223);
nor U6865 (N_6865,N_6372,N_6036);
nand U6866 (N_6866,N_6478,N_6077);
or U6867 (N_6867,N_6448,N_6097);
nor U6868 (N_6868,N_6249,N_6454);
or U6869 (N_6869,N_6144,N_6278);
xnor U6870 (N_6870,N_6128,N_6041);
or U6871 (N_6871,N_6110,N_6290);
xor U6872 (N_6872,N_6134,N_6064);
nand U6873 (N_6873,N_6191,N_6006);
nand U6874 (N_6874,N_6402,N_6307);
and U6875 (N_6875,N_6194,N_6001);
and U6876 (N_6876,N_6478,N_6078);
xor U6877 (N_6877,N_6311,N_6484);
nand U6878 (N_6878,N_6441,N_6227);
nor U6879 (N_6879,N_6499,N_6043);
or U6880 (N_6880,N_6248,N_6398);
nor U6881 (N_6881,N_6147,N_6264);
and U6882 (N_6882,N_6205,N_6432);
nor U6883 (N_6883,N_6285,N_6095);
nand U6884 (N_6884,N_6152,N_6475);
xor U6885 (N_6885,N_6438,N_6301);
and U6886 (N_6886,N_6194,N_6046);
or U6887 (N_6887,N_6472,N_6444);
nand U6888 (N_6888,N_6341,N_6337);
and U6889 (N_6889,N_6360,N_6120);
nand U6890 (N_6890,N_6140,N_6244);
nand U6891 (N_6891,N_6233,N_6072);
nand U6892 (N_6892,N_6410,N_6160);
or U6893 (N_6893,N_6009,N_6362);
and U6894 (N_6894,N_6013,N_6084);
and U6895 (N_6895,N_6190,N_6471);
and U6896 (N_6896,N_6171,N_6306);
and U6897 (N_6897,N_6028,N_6117);
or U6898 (N_6898,N_6110,N_6390);
or U6899 (N_6899,N_6419,N_6080);
nor U6900 (N_6900,N_6330,N_6121);
nand U6901 (N_6901,N_6059,N_6238);
or U6902 (N_6902,N_6432,N_6331);
nor U6903 (N_6903,N_6432,N_6126);
or U6904 (N_6904,N_6047,N_6025);
nor U6905 (N_6905,N_6391,N_6485);
or U6906 (N_6906,N_6314,N_6445);
and U6907 (N_6907,N_6222,N_6197);
xor U6908 (N_6908,N_6490,N_6014);
or U6909 (N_6909,N_6460,N_6106);
nand U6910 (N_6910,N_6030,N_6389);
xor U6911 (N_6911,N_6250,N_6068);
and U6912 (N_6912,N_6245,N_6322);
and U6913 (N_6913,N_6469,N_6443);
or U6914 (N_6914,N_6136,N_6495);
or U6915 (N_6915,N_6217,N_6382);
and U6916 (N_6916,N_6318,N_6384);
xor U6917 (N_6917,N_6025,N_6276);
or U6918 (N_6918,N_6491,N_6440);
nor U6919 (N_6919,N_6188,N_6016);
nand U6920 (N_6920,N_6255,N_6426);
nor U6921 (N_6921,N_6203,N_6195);
nor U6922 (N_6922,N_6263,N_6170);
and U6923 (N_6923,N_6400,N_6094);
and U6924 (N_6924,N_6295,N_6296);
nor U6925 (N_6925,N_6221,N_6488);
or U6926 (N_6926,N_6059,N_6017);
xor U6927 (N_6927,N_6148,N_6192);
nand U6928 (N_6928,N_6211,N_6265);
nand U6929 (N_6929,N_6415,N_6489);
nand U6930 (N_6930,N_6324,N_6230);
nor U6931 (N_6931,N_6084,N_6174);
nor U6932 (N_6932,N_6144,N_6450);
xnor U6933 (N_6933,N_6408,N_6494);
xor U6934 (N_6934,N_6259,N_6139);
xor U6935 (N_6935,N_6072,N_6419);
and U6936 (N_6936,N_6004,N_6441);
or U6937 (N_6937,N_6243,N_6196);
or U6938 (N_6938,N_6335,N_6455);
or U6939 (N_6939,N_6498,N_6412);
nand U6940 (N_6940,N_6137,N_6088);
and U6941 (N_6941,N_6085,N_6097);
nand U6942 (N_6942,N_6413,N_6081);
or U6943 (N_6943,N_6450,N_6315);
and U6944 (N_6944,N_6286,N_6094);
and U6945 (N_6945,N_6299,N_6124);
nor U6946 (N_6946,N_6085,N_6291);
or U6947 (N_6947,N_6165,N_6040);
and U6948 (N_6948,N_6152,N_6340);
xnor U6949 (N_6949,N_6402,N_6159);
nand U6950 (N_6950,N_6085,N_6407);
nand U6951 (N_6951,N_6480,N_6036);
nor U6952 (N_6952,N_6396,N_6019);
and U6953 (N_6953,N_6071,N_6486);
nand U6954 (N_6954,N_6466,N_6369);
and U6955 (N_6955,N_6170,N_6183);
and U6956 (N_6956,N_6248,N_6366);
nor U6957 (N_6957,N_6257,N_6244);
xor U6958 (N_6958,N_6425,N_6257);
nand U6959 (N_6959,N_6076,N_6041);
nand U6960 (N_6960,N_6060,N_6470);
or U6961 (N_6961,N_6049,N_6237);
and U6962 (N_6962,N_6051,N_6423);
nor U6963 (N_6963,N_6100,N_6280);
and U6964 (N_6964,N_6029,N_6250);
nor U6965 (N_6965,N_6207,N_6301);
and U6966 (N_6966,N_6260,N_6070);
xor U6967 (N_6967,N_6330,N_6197);
or U6968 (N_6968,N_6443,N_6170);
and U6969 (N_6969,N_6233,N_6276);
nor U6970 (N_6970,N_6252,N_6336);
or U6971 (N_6971,N_6272,N_6288);
nand U6972 (N_6972,N_6051,N_6495);
nor U6973 (N_6973,N_6407,N_6330);
nor U6974 (N_6974,N_6218,N_6047);
xnor U6975 (N_6975,N_6395,N_6446);
or U6976 (N_6976,N_6135,N_6348);
xor U6977 (N_6977,N_6262,N_6202);
xor U6978 (N_6978,N_6341,N_6064);
nand U6979 (N_6979,N_6115,N_6458);
nor U6980 (N_6980,N_6229,N_6472);
nor U6981 (N_6981,N_6173,N_6153);
or U6982 (N_6982,N_6347,N_6210);
and U6983 (N_6983,N_6215,N_6228);
or U6984 (N_6984,N_6409,N_6010);
and U6985 (N_6985,N_6188,N_6387);
and U6986 (N_6986,N_6116,N_6461);
nor U6987 (N_6987,N_6298,N_6371);
nor U6988 (N_6988,N_6453,N_6268);
and U6989 (N_6989,N_6036,N_6415);
nor U6990 (N_6990,N_6397,N_6006);
or U6991 (N_6991,N_6153,N_6149);
xor U6992 (N_6992,N_6033,N_6281);
nand U6993 (N_6993,N_6377,N_6498);
nand U6994 (N_6994,N_6253,N_6356);
nand U6995 (N_6995,N_6249,N_6005);
nor U6996 (N_6996,N_6213,N_6493);
and U6997 (N_6997,N_6338,N_6154);
xor U6998 (N_6998,N_6405,N_6317);
xor U6999 (N_6999,N_6099,N_6036);
nor U7000 (N_7000,N_6863,N_6767);
or U7001 (N_7001,N_6773,N_6821);
nor U7002 (N_7002,N_6528,N_6763);
nor U7003 (N_7003,N_6749,N_6544);
or U7004 (N_7004,N_6655,N_6661);
nand U7005 (N_7005,N_6728,N_6822);
or U7006 (N_7006,N_6825,N_6599);
xnor U7007 (N_7007,N_6628,N_6594);
xor U7008 (N_7008,N_6940,N_6941);
or U7009 (N_7009,N_6560,N_6748);
nand U7010 (N_7010,N_6747,N_6914);
or U7011 (N_7011,N_6675,N_6917);
nor U7012 (N_7012,N_6589,N_6903);
nand U7013 (N_7013,N_6627,N_6870);
nand U7014 (N_7014,N_6558,N_6952);
xnor U7015 (N_7015,N_6673,N_6760);
nor U7016 (N_7016,N_6835,N_6935);
nor U7017 (N_7017,N_6624,N_6851);
or U7018 (N_7018,N_6567,N_6788);
or U7019 (N_7019,N_6686,N_6768);
nor U7020 (N_7020,N_6826,N_6808);
nand U7021 (N_7021,N_6846,N_6575);
nand U7022 (N_7022,N_6755,N_6720);
nor U7023 (N_7023,N_6994,N_6910);
xnor U7024 (N_7024,N_6695,N_6936);
nor U7025 (N_7025,N_6705,N_6644);
nor U7026 (N_7026,N_6895,N_6996);
or U7027 (N_7027,N_6754,N_6885);
xor U7028 (N_7028,N_6837,N_6850);
or U7029 (N_7029,N_6897,N_6904);
and U7030 (N_7030,N_6569,N_6777);
and U7031 (N_7031,N_6953,N_6758);
nor U7032 (N_7032,N_6789,N_6770);
nor U7033 (N_7033,N_6666,N_6981);
nand U7034 (N_7034,N_6992,N_6798);
nand U7035 (N_7035,N_6933,N_6593);
nor U7036 (N_7036,N_6919,N_6576);
nor U7037 (N_7037,N_6510,N_6949);
xnor U7038 (N_7038,N_6684,N_6968);
and U7039 (N_7039,N_6871,N_6657);
or U7040 (N_7040,N_6838,N_6750);
and U7041 (N_7041,N_6667,N_6659);
xnor U7042 (N_7042,N_6916,N_6557);
nor U7043 (N_7043,N_6784,N_6762);
nand U7044 (N_7044,N_6988,N_6840);
and U7045 (N_7045,N_6813,N_6950);
nor U7046 (N_7046,N_6900,N_6712);
and U7047 (N_7047,N_6793,N_6766);
nor U7048 (N_7048,N_6847,N_6960);
or U7049 (N_7049,N_6797,N_6591);
nor U7050 (N_7050,N_6946,N_6753);
or U7051 (N_7051,N_6639,N_6527);
or U7052 (N_7052,N_6504,N_6991);
or U7053 (N_7053,N_6564,N_6783);
and U7054 (N_7054,N_6679,N_6725);
nor U7055 (N_7055,N_6577,N_6807);
or U7056 (N_7056,N_6868,N_6891);
nand U7057 (N_7057,N_6764,N_6631);
or U7058 (N_7058,N_6948,N_6608);
nor U7059 (N_7059,N_6774,N_6892);
xnor U7060 (N_7060,N_6611,N_6610);
and U7061 (N_7061,N_6615,N_6939);
and U7062 (N_7062,N_6723,N_6967);
or U7063 (N_7063,N_6596,N_6697);
xnor U7064 (N_7064,N_6606,N_6781);
nor U7065 (N_7065,N_6721,N_6523);
xnor U7066 (N_7066,N_6964,N_6573);
nor U7067 (N_7067,N_6713,N_6894);
nand U7068 (N_7068,N_6621,N_6524);
nand U7069 (N_7069,N_6539,N_6632);
nor U7070 (N_7070,N_6787,N_6913);
nor U7071 (N_7071,N_6526,N_6711);
nor U7072 (N_7072,N_6683,N_6799);
xnor U7073 (N_7073,N_6654,N_6827);
and U7074 (N_7074,N_6906,N_6926);
nand U7075 (N_7075,N_6884,N_6566);
nand U7076 (N_7076,N_6902,N_6603);
nor U7077 (N_7077,N_6972,N_6693);
nand U7078 (N_7078,N_6898,N_6701);
and U7079 (N_7079,N_6974,N_6842);
or U7080 (N_7080,N_6987,N_6522);
nor U7081 (N_7081,N_6928,N_6961);
nand U7082 (N_7082,N_6700,N_6841);
and U7083 (N_7083,N_6865,N_6636);
nand U7084 (N_7084,N_6989,N_6809);
xor U7085 (N_7085,N_6899,N_6735);
nor U7086 (N_7086,N_6857,N_6844);
nor U7087 (N_7087,N_6699,N_6739);
or U7088 (N_7088,N_6872,N_6722);
and U7089 (N_7089,N_6796,N_6732);
or U7090 (N_7090,N_6530,N_6970);
nand U7091 (N_7091,N_6612,N_6958);
nor U7092 (N_7092,N_6779,N_6811);
or U7093 (N_7093,N_6703,N_6652);
or U7094 (N_7094,N_6640,N_6518);
xor U7095 (N_7095,N_6782,N_6506);
and U7096 (N_7096,N_6890,N_6918);
nor U7097 (N_7097,N_6927,N_6617);
or U7098 (N_7098,N_6819,N_6944);
or U7099 (N_7099,N_6543,N_6555);
xor U7100 (N_7100,N_6859,N_6889);
nor U7101 (N_7101,N_6924,N_6795);
nand U7102 (N_7102,N_6529,N_6715);
nor U7103 (N_7103,N_6647,N_6586);
or U7104 (N_7104,N_6814,N_6832);
xor U7105 (N_7105,N_6601,N_6828);
or U7106 (N_7106,N_6546,N_6729);
xor U7107 (N_7107,N_6947,N_6909);
xor U7108 (N_7108,N_6930,N_6867);
and U7109 (N_7109,N_6716,N_6737);
nand U7110 (N_7110,N_6545,N_6873);
or U7111 (N_7111,N_6780,N_6669);
or U7112 (N_7112,N_6696,N_6502);
or U7113 (N_7113,N_6790,N_6671);
or U7114 (N_7114,N_6641,N_6771);
and U7115 (N_7115,N_6775,N_6761);
or U7116 (N_7116,N_6574,N_6551);
and U7117 (N_7117,N_6525,N_6810);
nand U7118 (N_7118,N_6800,N_6507);
or U7119 (N_7119,N_6681,N_6658);
xnor U7120 (N_7120,N_6533,N_6578);
and U7121 (N_7121,N_6689,N_6938);
nor U7122 (N_7122,N_6687,N_6839);
or U7123 (N_7123,N_6806,N_6532);
xor U7124 (N_7124,N_6776,N_6547);
xnor U7125 (N_7125,N_6500,N_6643);
nand U7126 (N_7126,N_6619,N_6559);
or U7127 (N_7127,N_6975,N_6665);
nand U7128 (N_7128,N_6887,N_6668);
or U7129 (N_7129,N_6794,N_6911);
nor U7130 (N_7130,N_6549,N_6959);
and U7131 (N_7131,N_6688,N_6538);
nor U7132 (N_7132,N_6923,N_6605);
xor U7133 (N_7133,N_6934,N_6583);
and U7134 (N_7134,N_6702,N_6585);
nor U7135 (N_7135,N_6678,N_6620);
xnor U7136 (N_7136,N_6664,N_6509);
nand U7137 (N_7137,N_6874,N_6756);
and U7138 (N_7138,N_6600,N_6912);
nor U7139 (N_7139,N_6663,N_6519);
or U7140 (N_7140,N_6932,N_6957);
and U7141 (N_7141,N_6694,N_6517);
xor U7142 (N_7142,N_6646,N_6623);
or U7143 (N_7143,N_6733,N_6531);
nor U7144 (N_7144,N_6690,N_6896);
nand U7145 (N_7145,N_6581,N_6893);
and U7146 (N_7146,N_6503,N_6740);
nand U7147 (N_7147,N_6830,N_6922);
nor U7148 (N_7148,N_6986,N_6805);
nand U7149 (N_7149,N_6542,N_6786);
nor U7150 (N_7150,N_6829,N_6804);
nand U7151 (N_7151,N_6820,N_6717);
nand U7152 (N_7152,N_6855,N_6993);
xnor U7153 (N_7153,N_6937,N_6979);
and U7154 (N_7154,N_6719,N_6757);
nor U7155 (N_7155,N_6843,N_6536);
or U7156 (N_7156,N_6877,N_6505);
xnor U7157 (N_7157,N_6718,N_6625);
and U7158 (N_7158,N_6812,N_6598);
or U7159 (N_7159,N_6751,N_6556);
nand U7160 (N_7160,N_6571,N_6582);
or U7161 (N_7161,N_6866,N_6744);
nand U7162 (N_7162,N_6609,N_6584);
xnor U7163 (N_7163,N_6965,N_6633);
and U7164 (N_7164,N_6626,N_6836);
or U7165 (N_7165,N_6604,N_6710);
nor U7166 (N_7166,N_6672,N_6561);
nand U7167 (N_7167,N_6513,N_6685);
nor U7168 (N_7168,N_6514,N_6511);
and U7169 (N_7169,N_6929,N_6920);
or U7170 (N_7170,N_6709,N_6976);
and U7171 (N_7171,N_6515,N_6691);
or U7172 (N_7172,N_6879,N_6580);
xnor U7173 (N_7173,N_6572,N_6864);
nand U7174 (N_7174,N_6548,N_6618);
nor U7175 (N_7175,N_6951,N_6971);
and U7176 (N_7176,N_6590,N_6802);
xor U7177 (N_7177,N_6676,N_6995);
nand U7178 (N_7178,N_6845,N_6521);
or U7179 (N_7179,N_6653,N_6831);
nor U7180 (N_7180,N_6680,N_6818);
and U7181 (N_7181,N_6925,N_6942);
xor U7182 (N_7182,N_6724,N_6833);
xor U7183 (N_7183,N_6982,N_6734);
xnor U7184 (N_7184,N_6662,N_6956);
and U7185 (N_7185,N_6848,N_6607);
and U7186 (N_7186,N_6597,N_6858);
nand U7187 (N_7187,N_6704,N_6645);
nand U7188 (N_7188,N_6563,N_6656);
or U7189 (N_7189,N_6772,N_6651);
or U7190 (N_7190,N_6962,N_6803);
xor U7191 (N_7191,N_6708,N_6512);
and U7192 (N_7192,N_6706,N_6540);
nand U7193 (N_7193,N_6856,N_6905);
nor U7194 (N_7194,N_6769,N_6943);
xnor U7195 (N_7195,N_6554,N_6650);
xnor U7196 (N_7196,N_6614,N_6587);
nand U7197 (N_7197,N_6537,N_6985);
nor U7198 (N_7198,N_6516,N_6876);
xor U7199 (N_7199,N_6908,N_6778);
and U7200 (N_7200,N_6736,N_6973);
nor U7201 (N_7201,N_6634,N_6550);
nand U7202 (N_7202,N_6860,N_6570);
or U7203 (N_7203,N_6853,N_6714);
nand U7204 (N_7204,N_6823,N_6854);
nor U7205 (N_7205,N_6997,N_6815);
nand U7206 (N_7206,N_6743,N_6955);
nor U7207 (N_7207,N_6595,N_6726);
nand U7208 (N_7208,N_6727,N_6535);
nand U7209 (N_7209,N_6978,N_6963);
nor U7210 (N_7210,N_6852,N_6579);
nor U7211 (N_7211,N_6745,N_6875);
nand U7212 (N_7212,N_6785,N_6801);
or U7213 (N_7213,N_6742,N_6738);
and U7214 (N_7214,N_6670,N_6501);
and U7215 (N_7215,N_6999,N_6980);
or U7216 (N_7216,N_6707,N_6969);
or U7217 (N_7217,N_6752,N_6954);
and U7218 (N_7218,N_6966,N_6637);
nor U7219 (N_7219,N_6886,N_6834);
and U7220 (N_7220,N_6592,N_6881);
nor U7221 (N_7221,N_6677,N_6588);
or U7222 (N_7222,N_6552,N_6622);
or U7223 (N_7223,N_6945,N_6862);
nand U7224 (N_7224,N_6629,N_6824);
and U7225 (N_7225,N_6731,N_6534);
or U7226 (N_7226,N_6730,N_6816);
nor U7227 (N_7227,N_6541,N_6791);
nand U7228 (N_7228,N_6817,N_6983);
and U7229 (N_7229,N_6792,N_6682);
and U7230 (N_7230,N_6921,N_6616);
xor U7231 (N_7231,N_6613,N_6901);
or U7232 (N_7232,N_6869,N_6698);
and U7233 (N_7233,N_6998,N_6888);
nand U7234 (N_7234,N_6553,N_6849);
nand U7235 (N_7235,N_6915,N_6520);
nand U7236 (N_7236,N_6880,N_6630);
nor U7237 (N_7237,N_6649,N_6882);
nor U7238 (N_7238,N_6674,N_6602);
nand U7239 (N_7239,N_6692,N_6878);
nor U7240 (N_7240,N_6990,N_6638);
nor U7241 (N_7241,N_6508,N_6642);
and U7242 (N_7242,N_6759,N_6883);
xor U7243 (N_7243,N_6741,N_6648);
nor U7244 (N_7244,N_6907,N_6660);
and U7245 (N_7245,N_6635,N_6568);
xor U7246 (N_7246,N_6931,N_6746);
nand U7247 (N_7247,N_6562,N_6861);
or U7248 (N_7248,N_6977,N_6984);
or U7249 (N_7249,N_6765,N_6565);
nor U7250 (N_7250,N_6676,N_6959);
nor U7251 (N_7251,N_6510,N_6834);
xor U7252 (N_7252,N_6597,N_6974);
and U7253 (N_7253,N_6540,N_6672);
xor U7254 (N_7254,N_6569,N_6597);
xor U7255 (N_7255,N_6548,N_6630);
xnor U7256 (N_7256,N_6799,N_6585);
and U7257 (N_7257,N_6513,N_6569);
nand U7258 (N_7258,N_6558,N_6810);
xor U7259 (N_7259,N_6681,N_6938);
and U7260 (N_7260,N_6894,N_6828);
nor U7261 (N_7261,N_6648,N_6538);
nor U7262 (N_7262,N_6748,N_6788);
or U7263 (N_7263,N_6702,N_6797);
nor U7264 (N_7264,N_6873,N_6619);
nand U7265 (N_7265,N_6603,N_6826);
and U7266 (N_7266,N_6804,N_6557);
and U7267 (N_7267,N_6551,N_6793);
or U7268 (N_7268,N_6584,N_6985);
nand U7269 (N_7269,N_6500,N_6762);
xnor U7270 (N_7270,N_6770,N_6952);
xor U7271 (N_7271,N_6896,N_6715);
xor U7272 (N_7272,N_6974,N_6581);
nand U7273 (N_7273,N_6535,N_6834);
xor U7274 (N_7274,N_6802,N_6846);
nor U7275 (N_7275,N_6920,N_6818);
nand U7276 (N_7276,N_6776,N_6900);
and U7277 (N_7277,N_6507,N_6729);
or U7278 (N_7278,N_6962,N_6661);
nand U7279 (N_7279,N_6851,N_6804);
or U7280 (N_7280,N_6746,N_6679);
nand U7281 (N_7281,N_6558,N_6617);
or U7282 (N_7282,N_6747,N_6839);
and U7283 (N_7283,N_6570,N_6618);
or U7284 (N_7284,N_6719,N_6899);
or U7285 (N_7285,N_6790,N_6850);
or U7286 (N_7286,N_6539,N_6651);
xor U7287 (N_7287,N_6673,N_6647);
or U7288 (N_7288,N_6613,N_6961);
nor U7289 (N_7289,N_6769,N_6721);
xnor U7290 (N_7290,N_6734,N_6550);
xor U7291 (N_7291,N_6827,N_6612);
xor U7292 (N_7292,N_6775,N_6603);
or U7293 (N_7293,N_6600,N_6886);
or U7294 (N_7294,N_6723,N_6791);
xnor U7295 (N_7295,N_6979,N_6906);
and U7296 (N_7296,N_6505,N_6677);
nor U7297 (N_7297,N_6743,N_6545);
and U7298 (N_7298,N_6941,N_6620);
nand U7299 (N_7299,N_6621,N_6795);
nor U7300 (N_7300,N_6938,N_6996);
and U7301 (N_7301,N_6661,N_6859);
or U7302 (N_7302,N_6586,N_6572);
nor U7303 (N_7303,N_6782,N_6671);
and U7304 (N_7304,N_6888,N_6896);
or U7305 (N_7305,N_6907,N_6936);
nor U7306 (N_7306,N_6844,N_6725);
nand U7307 (N_7307,N_6514,N_6989);
xnor U7308 (N_7308,N_6900,N_6644);
or U7309 (N_7309,N_6512,N_6534);
nand U7310 (N_7310,N_6723,N_6525);
nand U7311 (N_7311,N_6656,N_6890);
nor U7312 (N_7312,N_6602,N_6503);
or U7313 (N_7313,N_6664,N_6690);
nand U7314 (N_7314,N_6834,N_6725);
or U7315 (N_7315,N_6701,N_6508);
nand U7316 (N_7316,N_6715,N_6586);
and U7317 (N_7317,N_6983,N_6763);
nand U7318 (N_7318,N_6887,N_6570);
xnor U7319 (N_7319,N_6970,N_6931);
nand U7320 (N_7320,N_6561,N_6764);
nand U7321 (N_7321,N_6663,N_6955);
nand U7322 (N_7322,N_6576,N_6974);
or U7323 (N_7323,N_6743,N_6807);
or U7324 (N_7324,N_6752,N_6609);
nor U7325 (N_7325,N_6765,N_6931);
nor U7326 (N_7326,N_6869,N_6678);
xnor U7327 (N_7327,N_6606,N_6747);
and U7328 (N_7328,N_6888,N_6717);
or U7329 (N_7329,N_6862,N_6686);
nor U7330 (N_7330,N_6564,N_6877);
xor U7331 (N_7331,N_6537,N_6813);
nor U7332 (N_7332,N_6529,N_6561);
or U7333 (N_7333,N_6865,N_6776);
or U7334 (N_7334,N_6738,N_6575);
nor U7335 (N_7335,N_6579,N_6790);
or U7336 (N_7336,N_6667,N_6700);
xor U7337 (N_7337,N_6779,N_6692);
nand U7338 (N_7338,N_6869,N_6689);
and U7339 (N_7339,N_6701,N_6583);
or U7340 (N_7340,N_6918,N_6839);
or U7341 (N_7341,N_6685,N_6951);
or U7342 (N_7342,N_6926,N_6750);
and U7343 (N_7343,N_6509,N_6523);
or U7344 (N_7344,N_6893,N_6908);
and U7345 (N_7345,N_6654,N_6761);
nor U7346 (N_7346,N_6881,N_6564);
and U7347 (N_7347,N_6569,N_6623);
and U7348 (N_7348,N_6837,N_6913);
and U7349 (N_7349,N_6943,N_6941);
and U7350 (N_7350,N_6829,N_6963);
xor U7351 (N_7351,N_6891,N_6918);
nand U7352 (N_7352,N_6965,N_6781);
nand U7353 (N_7353,N_6808,N_6952);
or U7354 (N_7354,N_6896,N_6862);
and U7355 (N_7355,N_6664,N_6822);
nand U7356 (N_7356,N_6699,N_6870);
nor U7357 (N_7357,N_6881,N_6679);
nor U7358 (N_7358,N_6866,N_6805);
and U7359 (N_7359,N_6707,N_6672);
nor U7360 (N_7360,N_6754,N_6663);
or U7361 (N_7361,N_6917,N_6729);
or U7362 (N_7362,N_6625,N_6927);
xnor U7363 (N_7363,N_6851,N_6993);
or U7364 (N_7364,N_6989,N_6505);
nand U7365 (N_7365,N_6838,N_6775);
xnor U7366 (N_7366,N_6800,N_6577);
xnor U7367 (N_7367,N_6874,N_6741);
and U7368 (N_7368,N_6632,N_6542);
nand U7369 (N_7369,N_6873,N_6656);
and U7370 (N_7370,N_6776,N_6825);
nand U7371 (N_7371,N_6860,N_6700);
nor U7372 (N_7372,N_6716,N_6797);
xnor U7373 (N_7373,N_6943,N_6926);
nor U7374 (N_7374,N_6589,N_6803);
or U7375 (N_7375,N_6644,N_6778);
or U7376 (N_7376,N_6574,N_6837);
and U7377 (N_7377,N_6995,N_6992);
nor U7378 (N_7378,N_6742,N_6866);
and U7379 (N_7379,N_6691,N_6660);
nand U7380 (N_7380,N_6711,N_6787);
xnor U7381 (N_7381,N_6795,N_6640);
or U7382 (N_7382,N_6603,N_6853);
nor U7383 (N_7383,N_6795,N_6643);
xor U7384 (N_7384,N_6760,N_6823);
nor U7385 (N_7385,N_6524,N_6831);
xnor U7386 (N_7386,N_6928,N_6855);
nor U7387 (N_7387,N_6793,N_6700);
xnor U7388 (N_7388,N_6954,N_6670);
nor U7389 (N_7389,N_6956,N_6673);
nor U7390 (N_7390,N_6591,N_6942);
and U7391 (N_7391,N_6836,N_6770);
nand U7392 (N_7392,N_6646,N_6641);
nand U7393 (N_7393,N_6574,N_6972);
and U7394 (N_7394,N_6660,N_6721);
and U7395 (N_7395,N_6640,N_6636);
or U7396 (N_7396,N_6952,N_6749);
or U7397 (N_7397,N_6894,N_6517);
and U7398 (N_7398,N_6579,N_6869);
xor U7399 (N_7399,N_6658,N_6685);
nor U7400 (N_7400,N_6838,N_6589);
and U7401 (N_7401,N_6946,N_6929);
or U7402 (N_7402,N_6687,N_6762);
nand U7403 (N_7403,N_6540,N_6927);
nand U7404 (N_7404,N_6549,N_6741);
nand U7405 (N_7405,N_6534,N_6732);
xnor U7406 (N_7406,N_6679,N_6633);
nand U7407 (N_7407,N_6797,N_6690);
nand U7408 (N_7408,N_6563,N_6588);
nand U7409 (N_7409,N_6683,N_6632);
nor U7410 (N_7410,N_6615,N_6707);
and U7411 (N_7411,N_6586,N_6728);
nor U7412 (N_7412,N_6761,N_6668);
and U7413 (N_7413,N_6543,N_6722);
and U7414 (N_7414,N_6738,N_6774);
nor U7415 (N_7415,N_6608,N_6911);
nand U7416 (N_7416,N_6634,N_6901);
nand U7417 (N_7417,N_6677,N_6570);
xnor U7418 (N_7418,N_6517,N_6792);
xnor U7419 (N_7419,N_6811,N_6595);
xnor U7420 (N_7420,N_6575,N_6656);
xor U7421 (N_7421,N_6607,N_6816);
nor U7422 (N_7422,N_6740,N_6536);
xor U7423 (N_7423,N_6933,N_6823);
and U7424 (N_7424,N_6629,N_6963);
xor U7425 (N_7425,N_6847,N_6940);
xor U7426 (N_7426,N_6806,N_6840);
nand U7427 (N_7427,N_6653,N_6566);
or U7428 (N_7428,N_6730,N_6964);
or U7429 (N_7429,N_6630,N_6899);
or U7430 (N_7430,N_6761,N_6757);
nor U7431 (N_7431,N_6513,N_6789);
and U7432 (N_7432,N_6908,N_6995);
nand U7433 (N_7433,N_6783,N_6820);
or U7434 (N_7434,N_6530,N_6515);
and U7435 (N_7435,N_6553,N_6662);
nor U7436 (N_7436,N_6649,N_6519);
nor U7437 (N_7437,N_6977,N_6542);
or U7438 (N_7438,N_6508,N_6972);
nor U7439 (N_7439,N_6726,N_6976);
and U7440 (N_7440,N_6507,N_6741);
and U7441 (N_7441,N_6599,N_6882);
xnor U7442 (N_7442,N_6665,N_6937);
and U7443 (N_7443,N_6726,N_6845);
nor U7444 (N_7444,N_6609,N_6728);
and U7445 (N_7445,N_6927,N_6958);
or U7446 (N_7446,N_6952,N_6852);
or U7447 (N_7447,N_6818,N_6901);
nand U7448 (N_7448,N_6827,N_6697);
or U7449 (N_7449,N_6806,N_6602);
nand U7450 (N_7450,N_6853,N_6979);
nand U7451 (N_7451,N_6831,N_6886);
nor U7452 (N_7452,N_6816,N_6639);
and U7453 (N_7453,N_6583,N_6900);
or U7454 (N_7454,N_6954,N_6691);
or U7455 (N_7455,N_6809,N_6782);
and U7456 (N_7456,N_6505,N_6515);
nand U7457 (N_7457,N_6682,N_6966);
nor U7458 (N_7458,N_6795,N_6521);
xor U7459 (N_7459,N_6510,N_6844);
nor U7460 (N_7460,N_6514,N_6699);
nand U7461 (N_7461,N_6917,N_6680);
or U7462 (N_7462,N_6849,N_6688);
or U7463 (N_7463,N_6730,N_6607);
xnor U7464 (N_7464,N_6693,N_6748);
nor U7465 (N_7465,N_6810,N_6923);
or U7466 (N_7466,N_6882,N_6698);
nand U7467 (N_7467,N_6560,N_6758);
nor U7468 (N_7468,N_6552,N_6531);
xnor U7469 (N_7469,N_6823,N_6532);
xnor U7470 (N_7470,N_6924,N_6596);
or U7471 (N_7471,N_6634,N_6647);
xnor U7472 (N_7472,N_6899,N_6593);
nor U7473 (N_7473,N_6635,N_6927);
or U7474 (N_7474,N_6638,N_6652);
or U7475 (N_7475,N_6942,N_6527);
xor U7476 (N_7476,N_6588,N_6596);
nand U7477 (N_7477,N_6863,N_6830);
or U7478 (N_7478,N_6669,N_6929);
nand U7479 (N_7479,N_6870,N_6871);
and U7480 (N_7480,N_6812,N_6681);
nand U7481 (N_7481,N_6553,N_6511);
xor U7482 (N_7482,N_6903,N_6708);
and U7483 (N_7483,N_6797,N_6508);
xor U7484 (N_7484,N_6608,N_6958);
xnor U7485 (N_7485,N_6980,N_6580);
or U7486 (N_7486,N_6540,N_6802);
or U7487 (N_7487,N_6510,N_6716);
or U7488 (N_7488,N_6650,N_6802);
xor U7489 (N_7489,N_6994,N_6658);
nand U7490 (N_7490,N_6535,N_6784);
or U7491 (N_7491,N_6692,N_6944);
and U7492 (N_7492,N_6935,N_6898);
nor U7493 (N_7493,N_6862,N_6729);
or U7494 (N_7494,N_6703,N_6742);
and U7495 (N_7495,N_6705,N_6756);
or U7496 (N_7496,N_6612,N_6806);
or U7497 (N_7497,N_6984,N_6949);
xnor U7498 (N_7498,N_6956,N_6543);
or U7499 (N_7499,N_6579,N_6926);
or U7500 (N_7500,N_7382,N_7280);
and U7501 (N_7501,N_7306,N_7246);
and U7502 (N_7502,N_7424,N_7353);
nand U7503 (N_7503,N_7465,N_7021);
and U7504 (N_7504,N_7232,N_7368);
and U7505 (N_7505,N_7176,N_7401);
or U7506 (N_7506,N_7073,N_7298);
nor U7507 (N_7507,N_7239,N_7242);
nor U7508 (N_7508,N_7264,N_7127);
xnor U7509 (N_7509,N_7484,N_7463);
or U7510 (N_7510,N_7468,N_7215);
nor U7511 (N_7511,N_7235,N_7479);
xor U7512 (N_7512,N_7376,N_7388);
or U7513 (N_7513,N_7128,N_7076);
and U7514 (N_7514,N_7352,N_7301);
or U7515 (N_7515,N_7348,N_7065);
xor U7516 (N_7516,N_7360,N_7358);
nor U7517 (N_7517,N_7174,N_7123);
or U7518 (N_7518,N_7198,N_7109);
xor U7519 (N_7519,N_7008,N_7071);
xnor U7520 (N_7520,N_7053,N_7346);
nand U7521 (N_7521,N_7207,N_7419);
and U7522 (N_7522,N_7381,N_7228);
nand U7523 (N_7523,N_7034,N_7044);
xnor U7524 (N_7524,N_7085,N_7278);
nand U7525 (N_7525,N_7254,N_7316);
or U7526 (N_7526,N_7212,N_7236);
xnor U7527 (N_7527,N_7377,N_7384);
xor U7528 (N_7528,N_7051,N_7456);
nand U7529 (N_7529,N_7092,N_7320);
nor U7530 (N_7530,N_7192,N_7119);
or U7531 (N_7531,N_7074,N_7366);
xor U7532 (N_7532,N_7116,N_7031);
nor U7533 (N_7533,N_7057,N_7422);
and U7534 (N_7534,N_7488,N_7300);
nor U7535 (N_7535,N_7035,N_7441);
nor U7536 (N_7536,N_7025,N_7299);
nand U7537 (N_7537,N_7446,N_7194);
and U7538 (N_7538,N_7030,N_7131);
nor U7539 (N_7539,N_7169,N_7343);
nor U7540 (N_7540,N_7062,N_7233);
xnor U7541 (N_7541,N_7361,N_7165);
and U7542 (N_7542,N_7371,N_7181);
nor U7543 (N_7543,N_7262,N_7311);
or U7544 (N_7544,N_7155,N_7022);
nand U7545 (N_7545,N_7494,N_7158);
xor U7546 (N_7546,N_7244,N_7309);
nor U7547 (N_7547,N_7394,N_7187);
nand U7548 (N_7548,N_7277,N_7037);
xor U7549 (N_7549,N_7237,N_7032);
nand U7550 (N_7550,N_7010,N_7349);
and U7551 (N_7551,N_7136,N_7436);
xor U7552 (N_7552,N_7435,N_7493);
xor U7553 (N_7553,N_7243,N_7407);
nand U7554 (N_7554,N_7213,N_7279);
xor U7555 (N_7555,N_7081,N_7075);
xor U7556 (N_7556,N_7362,N_7240);
and U7557 (N_7557,N_7470,N_7006);
or U7558 (N_7558,N_7414,N_7383);
xnor U7559 (N_7559,N_7400,N_7129);
or U7560 (N_7560,N_7270,N_7045);
xor U7561 (N_7561,N_7378,N_7390);
and U7562 (N_7562,N_7266,N_7147);
or U7563 (N_7563,N_7221,N_7372);
nor U7564 (N_7564,N_7173,N_7137);
nand U7565 (N_7565,N_7043,N_7427);
and U7566 (N_7566,N_7012,N_7157);
xnor U7567 (N_7567,N_7229,N_7061);
and U7568 (N_7568,N_7079,N_7024);
xor U7569 (N_7569,N_7354,N_7249);
nor U7570 (N_7570,N_7196,N_7370);
or U7571 (N_7571,N_7340,N_7448);
or U7572 (N_7572,N_7029,N_7195);
and U7573 (N_7573,N_7175,N_7047);
nor U7574 (N_7574,N_7313,N_7052);
xor U7575 (N_7575,N_7337,N_7009);
or U7576 (N_7576,N_7283,N_7184);
or U7577 (N_7577,N_7201,N_7310);
nor U7578 (N_7578,N_7087,N_7408);
or U7579 (N_7579,N_7102,N_7151);
and U7580 (N_7580,N_7159,N_7342);
nand U7581 (N_7581,N_7106,N_7039);
and U7582 (N_7582,N_7190,N_7486);
xnor U7583 (N_7583,N_7185,N_7013);
xor U7584 (N_7584,N_7296,N_7002);
nor U7585 (N_7585,N_7007,N_7124);
nor U7586 (N_7586,N_7373,N_7095);
nand U7587 (N_7587,N_7336,N_7125);
and U7588 (N_7588,N_7023,N_7485);
nand U7589 (N_7589,N_7223,N_7001);
nand U7590 (N_7590,N_7405,N_7292);
or U7591 (N_7591,N_7150,N_7058);
or U7592 (N_7592,N_7259,N_7210);
and U7593 (N_7593,N_7209,N_7252);
xnor U7594 (N_7594,N_7255,N_7154);
nor U7595 (N_7595,N_7345,N_7459);
or U7596 (N_7596,N_7303,N_7206);
xor U7597 (N_7597,N_7224,N_7417);
xnor U7598 (N_7598,N_7049,N_7261);
xor U7599 (N_7599,N_7433,N_7046);
or U7600 (N_7600,N_7458,N_7449);
nand U7601 (N_7601,N_7028,N_7420);
nor U7602 (N_7602,N_7171,N_7250);
nor U7603 (N_7603,N_7481,N_7096);
nand U7604 (N_7604,N_7117,N_7308);
nand U7605 (N_7605,N_7330,N_7005);
nand U7606 (N_7606,N_7347,N_7273);
nand U7607 (N_7607,N_7122,N_7097);
or U7608 (N_7608,N_7080,N_7466);
or U7609 (N_7609,N_7317,N_7335);
nand U7610 (N_7610,N_7395,N_7197);
nor U7611 (N_7611,N_7359,N_7398);
and U7612 (N_7612,N_7186,N_7231);
or U7613 (N_7613,N_7163,N_7480);
nand U7614 (N_7614,N_7130,N_7048);
or U7615 (N_7615,N_7018,N_7225);
xnor U7616 (N_7616,N_7226,N_7385);
or U7617 (N_7617,N_7072,N_7139);
or U7618 (N_7618,N_7134,N_7403);
nor U7619 (N_7619,N_7247,N_7302);
nor U7620 (N_7620,N_7329,N_7219);
or U7621 (N_7621,N_7418,N_7295);
nor U7622 (N_7622,N_7341,N_7364);
nand U7623 (N_7623,N_7434,N_7275);
xnor U7624 (N_7624,N_7357,N_7100);
xor U7625 (N_7625,N_7016,N_7258);
xnor U7626 (N_7626,N_7033,N_7082);
nor U7627 (N_7627,N_7211,N_7166);
or U7628 (N_7628,N_7497,N_7487);
nor U7629 (N_7629,N_7220,N_7443);
nor U7630 (N_7630,N_7289,N_7339);
nand U7631 (N_7631,N_7406,N_7386);
xnor U7632 (N_7632,N_7202,N_7482);
or U7633 (N_7633,N_7396,N_7321);
xor U7634 (N_7634,N_7293,N_7003);
xnor U7635 (N_7635,N_7307,N_7068);
or U7636 (N_7636,N_7274,N_7036);
or U7637 (N_7637,N_7115,N_7241);
xnor U7638 (N_7638,N_7291,N_7344);
xor U7639 (N_7639,N_7338,N_7204);
and U7640 (N_7640,N_7491,N_7294);
or U7641 (N_7641,N_7440,N_7140);
and U7642 (N_7642,N_7409,N_7326);
nor U7643 (N_7643,N_7217,N_7462);
nand U7644 (N_7644,N_7457,N_7064);
and U7645 (N_7645,N_7251,N_7234);
nand U7646 (N_7646,N_7020,N_7084);
and U7647 (N_7647,N_7438,N_7170);
or U7648 (N_7648,N_7467,N_7411);
and U7649 (N_7649,N_7365,N_7474);
and U7650 (N_7650,N_7268,N_7415);
xnor U7651 (N_7651,N_7112,N_7322);
nor U7652 (N_7652,N_7067,N_7426);
xnor U7653 (N_7653,N_7297,N_7138);
and U7654 (N_7654,N_7105,N_7141);
or U7655 (N_7655,N_7077,N_7056);
and U7656 (N_7656,N_7253,N_7256);
or U7657 (N_7657,N_7152,N_7069);
and U7658 (N_7658,N_7121,N_7319);
or U7659 (N_7659,N_7282,N_7019);
nand U7660 (N_7660,N_7327,N_7189);
or U7661 (N_7661,N_7014,N_7355);
nand U7662 (N_7662,N_7450,N_7496);
nand U7663 (N_7663,N_7055,N_7286);
nand U7664 (N_7664,N_7333,N_7478);
nor U7665 (N_7665,N_7476,N_7113);
xnor U7666 (N_7666,N_7290,N_7090);
nand U7667 (N_7667,N_7284,N_7432);
nor U7668 (N_7668,N_7379,N_7040);
and U7669 (N_7669,N_7059,N_7318);
nor U7670 (N_7670,N_7285,N_7111);
xnor U7671 (N_7671,N_7227,N_7063);
nand U7672 (N_7672,N_7107,N_7177);
and U7673 (N_7673,N_7315,N_7332);
and U7674 (N_7674,N_7042,N_7135);
xnor U7675 (N_7675,N_7182,N_7089);
and U7676 (N_7676,N_7464,N_7091);
xnor U7677 (N_7677,N_7161,N_7054);
or U7678 (N_7678,N_7499,N_7216);
nor U7679 (N_7679,N_7205,N_7203);
nor U7680 (N_7680,N_7167,N_7222);
nand U7681 (N_7681,N_7011,N_7445);
and U7682 (N_7682,N_7451,N_7188);
nand U7683 (N_7683,N_7200,N_7144);
nand U7684 (N_7684,N_7421,N_7389);
and U7685 (N_7685,N_7269,N_7410);
nor U7686 (N_7686,N_7126,N_7413);
or U7687 (N_7687,N_7015,N_7444);
nor U7688 (N_7688,N_7331,N_7245);
nor U7689 (N_7689,N_7118,N_7145);
and U7690 (N_7690,N_7455,N_7108);
nor U7691 (N_7691,N_7325,N_7066);
and U7692 (N_7692,N_7399,N_7180);
nor U7693 (N_7693,N_7490,N_7142);
nand U7694 (N_7694,N_7238,N_7199);
xor U7695 (N_7695,N_7439,N_7168);
nor U7696 (N_7696,N_7367,N_7000);
or U7697 (N_7697,N_7070,N_7489);
xnor U7698 (N_7698,N_7369,N_7156);
nor U7699 (N_7699,N_7387,N_7402);
nor U7700 (N_7700,N_7038,N_7263);
or U7701 (N_7701,N_7397,N_7143);
and U7702 (N_7702,N_7428,N_7447);
or U7703 (N_7703,N_7351,N_7356);
xor U7704 (N_7704,N_7230,N_7492);
nor U7705 (N_7705,N_7453,N_7208);
xor U7706 (N_7706,N_7477,N_7017);
nand U7707 (N_7707,N_7271,N_7257);
nor U7708 (N_7708,N_7179,N_7324);
and U7709 (N_7709,N_7281,N_7193);
nand U7710 (N_7710,N_7146,N_7248);
and U7711 (N_7711,N_7312,N_7276);
and U7712 (N_7712,N_7148,N_7114);
nand U7713 (N_7713,N_7483,N_7287);
nor U7714 (N_7714,N_7393,N_7363);
xnor U7715 (N_7715,N_7495,N_7218);
xnor U7716 (N_7716,N_7164,N_7172);
nor U7717 (N_7717,N_7120,N_7094);
nor U7718 (N_7718,N_7460,N_7412);
nor U7719 (N_7719,N_7391,N_7429);
nand U7720 (N_7720,N_7267,N_7026);
xnor U7721 (N_7721,N_7475,N_7191);
or U7722 (N_7722,N_7103,N_7093);
nand U7723 (N_7723,N_7304,N_7041);
and U7724 (N_7724,N_7454,N_7323);
and U7725 (N_7725,N_7423,N_7431);
or U7726 (N_7726,N_7098,N_7374);
xor U7727 (N_7727,N_7004,N_7160);
and U7728 (N_7728,N_7442,N_7088);
xnor U7729 (N_7729,N_7265,N_7050);
nand U7730 (N_7730,N_7452,N_7153);
xnor U7731 (N_7731,N_7214,N_7162);
xnor U7732 (N_7732,N_7375,N_7425);
nand U7733 (N_7733,N_7101,N_7083);
and U7734 (N_7734,N_7334,N_7473);
nor U7735 (N_7735,N_7416,N_7110);
nand U7736 (N_7736,N_7272,N_7471);
or U7737 (N_7737,N_7461,N_7132);
and U7738 (N_7738,N_7099,N_7350);
xor U7739 (N_7739,N_7328,N_7380);
and U7740 (N_7740,N_7149,N_7305);
nand U7741 (N_7741,N_7498,N_7104);
xnor U7742 (N_7742,N_7392,N_7060);
and U7743 (N_7743,N_7469,N_7430);
xnor U7744 (N_7744,N_7027,N_7133);
and U7745 (N_7745,N_7288,N_7437);
nand U7746 (N_7746,N_7086,N_7183);
xor U7747 (N_7747,N_7260,N_7178);
or U7748 (N_7748,N_7404,N_7078);
and U7749 (N_7749,N_7314,N_7472);
nand U7750 (N_7750,N_7402,N_7297);
nor U7751 (N_7751,N_7187,N_7227);
and U7752 (N_7752,N_7286,N_7236);
xor U7753 (N_7753,N_7051,N_7052);
nor U7754 (N_7754,N_7275,N_7472);
nor U7755 (N_7755,N_7016,N_7332);
xnor U7756 (N_7756,N_7153,N_7143);
nand U7757 (N_7757,N_7386,N_7402);
and U7758 (N_7758,N_7098,N_7334);
nor U7759 (N_7759,N_7141,N_7393);
and U7760 (N_7760,N_7384,N_7353);
or U7761 (N_7761,N_7007,N_7211);
and U7762 (N_7762,N_7489,N_7181);
or U7763 (N_7763,N_7440,N_7343);
xor U7764 (N_7764,N_7175,N_7222);
and U7765 (N_7765,N_7099,N_7468);
nand U7766 (N_7766,N_7321,N_7133);
nand U7767 (N_7767,N_7269,N_7120);
and U7768 (N_7768,N_7123,N_7403);
xnor U7769 (N_7769,N_7413,N_7202);
and U7770 (N_7770,N_7165,N_7239);
nand U7771 (N_7771,N_7071,N_7086);
xor U7772 (N_7772,N_7162,N_7187);
nor U7773 (N_7773,N_7050,N_7042);
xor U7774 (N_7774,N_7267,N_7064);
nand U7775 (N_7775,N_7471,N_7060);
xnor U7776 (N_7776,N_7370,N_7444);
or U7777 (N_7777,N_7040,N_7167);
nand U7778 (N_7778,N_7193,N_7300);
nand U7779 (N_7779,N_7345,N_7352);
nor U7780 (N_7780,N_7306,N_7262);
or U7781 (N_7781,N_7248,N_7043);
xnor U7782 (N_7782,N_7347,N_7396);
nor U7783 (N_7783,N_7458,N_7141);
nor U7784 (N_7784,N_7479,N_7325);
nor U7785 (N_7785,N_7269,N_7360);
nand U7786 (N_7786,N_7061,N_7449);
nor U7787 (N_7787,N_7370,N_7194);
or U7788 (N_7788,N_7058,N_7498);
xnor U7789 (N_7789,N_7169,N_7398);
and U7790 (N_7790,N_7423,N_7106);
xnor U7791 (N_7791,N_7245,N_7370);
xor U7792 (N_7792,N_7447,N_7029);
and U7793 (N_7793,N_7102,N_7362);
or U7794 (N_7794,N_7440,N_7170);
nand U7795 (N_7795,N_7302,N_7235);
nand U7796 (N_7796,N_7445,N_7331);
or U7797 (N_7797,N_7195,N_7132);
xor U7798 (N_7798,N_7208,N_7248);
nor U7799 (N_7799,N_7016,N_7072);
xnor U7800 (N_7800,N_7076,N_7402);
nand U7801 (N_7801,N_7167,N_7215);
and U7802 (N_7802,N_7024,N_7348);
or U7803 (N_7803,N_7445,N_7033);
xor U7804 (N_7804,N_7274,N_7238);
nor U7805 (N_7805,N_7418,N_7254);
and U7806 (N_7806,N_7469,N_7096);
nor U7807 (N_7807,N_7293,N_7065);
nand U7808 (N_7808,N_7094,N_7028);
xor U7809 (N_7809,N_7127,N_7386);
nand U7810 (N_7810,N_7064,N_7320);
xor U7811 (N_7811,N_7272,N_7473);
or U7812 (N_7812,N_7016,N_7436);
nand U7813 (N_7813,N_7199,N_7483);
xor U7814 (N_7814,N_7166,N_7406);
and U7815 (N_7815,N_7273,N_7133);
xor U7816 (N_7816,N_7197,N_7005);
and U7817 (N_7817,N_7205,N_7353);
nor U7818 (N_7818,N_7356,N_7342);
xnor U7819 (N_7819,N_7015,N_7495);
xnor U7820 (N_7820,N_7249,N_7417);
or U7821 (N_7821,N_7415,N_7250);
nand U7822 (N_7822,N_7021,N_7490);
nand U7823 (N_7823,N_7010,N_7115);
nand U7824 (N_7824,N_7263,N_7215);
or U7825 (N_7825,N_7010,N_7144);
nand U7826 (N_7826,N_7448,N_7413);
xnor U7827 (N_7827,N_7470,N_7394);
xnor U7828 (N_7828,N_7382,N_7316);
and U7829 (N_7829,N_7104,N_7283);
or U7830 (N_7830,N_7270,N_7237);
nand U7831 (N_7831,N_7130,N_7059);
nand U7832 (N_7832,N_7059,N_7221);
nand U7833 (N_7833,N_7118,N_7296);
or U7834 (N_7834,N_7062,N_7217);
or U7835 (N_7835,N_7089,N_7233);
and U7836 (N_7836,N_7353,N_7306);
or U7837 (N_7837,N_7097,N_7192);
xor U7838 (N_7838,N_7410,N_7207);
xnor U7839 (N_7839,N_7176,N_7360);
xnor U7840 (N_7840,N_7362,N_7379);
or U7841 (N_7841,N_7461,N_7049);
nor U7842 (N_7842,N_7233,N_7361);
xnor U7843 (N_7843,N_7378,N_7067);
and U7844 (N_7844,N_7031,N_7099);
nand U7845 (N_7845,N_7225,N_7485);
xnor U7846 (N_7846,N_7450,N_7145);
xor U7847 (N_7847,N_7089,N_7018);
xor U7848 (N_7848,N_7249,N_7363);
or U7849 (N_7849,N_7038,N_7279);
or U7850 (N_7850,N_7344,N_7390);
xnor U7851 (N_7851,N_7133,N_7226);
or U7852 (N_7852,N_7310,N_7293);
or U7853 (N_7853,N_7306,N_7197);
xnor U7854 (N_7854,N_7012,N_7426);
nand U7855 (N_7855,N_7217,N_7142);
or U7856 (N_7856,N_7175,N_7299);
or U7857 (N_7857,N_7320,N_7032);
or U7858 (N_7858,N_7188,N_7355);
xnor U7859 (N_7859,N_7243,N_7263);
xnor U7860 (N_7860,N_7238,N_7469);
xnor U7861 (N_7861,N_7377,N_7017);
or U7862 (N_7862,N_7092,N_7382);
or U7863 (N_7863,N_7393,N_7051);
nand U7864 (N_7864,N_7099,N_7363);
or U7865 (N_7865,N_7131,N_7027);
nor U7866 (N_7866,N_7014,N_7152);
and U7867 (N_7867,N_7212,N_7288);
xor U7868 (N_7868,N_7296,N_7481);
nor U7869 (N_7869,N_7464,N_7076);
nor U7870 (N_7870,N_7119,N_7098);
nor U7871 (N_7871,N_7120,N_7356);
xnor U7872 (N_7872,N_7241,N_7363);
nand U7873 (N_7873,N_7307,N_7078);
nand U7874 (N_7874,N_7010,N_7099);
or U7875 (N_7875,N_7178,N_7244);
nor U7876 (N_7876,N_7408,N_7379);
xor U7877 (N_7877,N_7164,N_7123);
xnor U7878 (N_7878,N_7478,N_7190);
nor U7879 (N_7879,N_7278,N_7125);
or U7880 (N_7880,N_7214,N_7403);
nor U7881 (N_7881,N_7056,N_7111);
and U7882 (N_7882,N_7427,N_7082);
nor U7883 (N_7883,N_7036,N_7472);
and U7884 (N_7884,N_7447,N_7199);
xor U7885 (N_7885,N_7322,N_7348);
xor U7886 (N_7886,N_7074,N_7222);
nor U7887 (N_7887,N_7287,N_7435);
and U7888 (N_7888,N_7362,N_7384);
and U7889 (N_7889,N_7103,N_7158);
or U7890 (N_7890,N_7490,N_7012);
and U7891 (N_7891,N_7020,N_7354);
and U7892 (N_7892,N_7411,N_7279);
and U7893 (N_7893,N_7449,N_7232);
xor U7894 (N_7894,N_7436,N_7276);
xor U7895 (N_7895,N_7273,N_7378);
nor U7896 (N_7896,N_7179,N_7036);
and U7897 (N_7897,N_7141,N_7052);
and U7898 (N_7898,N_7494,N_7475);
nand U7899 (N_7899,N_7115,N_7056);
and U7900 (N_7900,N_7470,N_7227);
nand U7901 (N_7901,N_7236,N_7453);
or U7902 (N_7902,N_7142,N_7364);
or U7903 (N_7903,N_7104,N_7213);
and U7904 (N_7904,N_7499,N_7152);
nand U7905 (N_7905,N_7116,N_7394);
nor U7906 (N_7906,N_7155,N_7054);
or U7907 (N_7907,N_7435,N_7219);
nor U7908 (N_7908,N_7180,N_7380);
and U7909 (N_7909,N_7309,N_7029);
nand U7910 (N_7910,N_7162,N_7303);
nor U7911 (N_7911,N_7148,N_7497);
xnor U7912 (N_7912,N_7125,N_7116);
nand U7913 (N_7913,N_7226,N_7240);
xnor U7914 (N_7914,N_7200,N_7371);
or U7915 (N_7915,N_7333,N_7317);
nor U7916 (N_7916,N_7052,N_7042);
and U7917 (N_7917,N_7340,N_7382);
or U7918 (N_7918,N_7106,N_7461);
and U7919 (N_7919,N_7122,N_7405);
and U7920 (N_7920,N_7279,N_7392);
or U7921 (N_7921,N_7233,N_7437);
nor U7922 (N_7922,N_7497,N_7119);
xnor U7923 (N_7923,N_7137,N_7290);
nand U7924 (N_7924,N_7221,N_7439);
nor U7925 (N_7925,N_7436,N_7008);
nand U7926 (N_7926,N_7342,N_7499);
nand U7927 (N_7927,N_7464,N_7161);
nor U7928 (N_7928,N_7400,N_7096);
or U7929 (N_7929,N_7202,N_7214);
or U7930 (N_7930,N_7082,N_7087);
xnor U7931 (N_7931,N_7453,N_7041);
nand U7932 (N_7932,N_7451,N_7415);
nor U7933 (N_7933,N_7134,N_7078);
nand U7934 (N_7934,N_7364,N_7420);
or U7935 (N_7935,N_7148,N_7141);
or U7936 (N_7936,N_7246,N_7149);
and U7937 (N_7937,N_7224,N_7491);
or U7938 (N_7938,N_7300,N_7308);
nand U7939 (N_7939,N_7276,N_7045);
xnor U7940 (N_7940,N_7297,N_7223);
and U7941 (N_7941,N_7196,N_7222);
xnor U7942 (N_7942,N_7117,N_7011);
nand U7943 (N_7943,N_7285,N_7294);
xor U7944 (N_7944,N_7091,N_7331);
or U7945 (N_7945,N_7199,N_7331);
or U7946 (N_7946,N_7457,N_7334);
nand U7947 (N_7947,N_7348,N_7004);
xnor U7948 (N_7948,N_7179,N_7050);
and U7949 (N_7949,N_7125,N_7477);
nor U7950 (N_7950,N_7202,N_7112);
xnor U7951 (N_7951,N_7064,N_7494);
nor U7952 (N_7952,N_7425,N_7227);
nor U7953 (N_7953,N_7145,N_7409);
or U7954 (N_7954,N_7027,N_7496);
nand U7955 (N_7955,N_7195,N_7226);
xor U7956 (N_7956,N_7402,N_7026);
nor U7957 (N_7957,N_7232,N_7172);
nor U7958 (N_7958,N_7025,N_7189);
nor U7959 (N_7959,N_7363,N_7471);
nand U7960 (N_7960,N_7474,N_7260);
nor U7961 (N_7961,N_7450,N_7338);
or U7962 (N_7962,N_7165,N_7411);
nand U7963 (N_7963,N_7478,N_7270);
nor U7964 (N_7964,N_7116,N_7175);
or U7965 (N_7965,N_7415,N_7343);
nor U7966 (N_7966,N_7152,N_7251);
nor U7967 (N_7967,N_7437,N_7294);
and U7968 (N_7968,N_7322,N_7064);
nand U7969 (N_7969,N_7335,N_7130);
and U7970 (N_7970,N_7170,N_7453);
nor U7971 (N_7971,N_7201,N_7115);
or U7972 (N_7972,N_7387,N_7467);
or U7973 (N_7973,N_7045,N_7252);
nand U7974 (N_7974,N_7438,N_7069);
nor U7975 (N_7975,N_7321,N_7079);
xor U7976 (N_7976,N_7384,N_7387);
xnor U7977 (N_7977,N_7363,N_7389);
nor U7978 (N_7978,N_7164,N_7246);
nand U7979 (N_7979,N_7314,N_7031);
or U7980 (N_7980,N_7354,N_7494);
or U7981 (N_7981,N_7112,N_7118);
or U7982 (N_7982,N_7083,N_7211);
nor U7983 (N_7983,N_7143,N_7434);
xor U7984 (N_7984,N_7135,N_7400);
xor U7985 (N_7985,N_7295,N_7375);
and U7986 (N_7986,N_7045,N_7072);
nand U7987 (N_7987,N_7375,N_7434);
and U7988 (N_7988,N_7043,N_7346);
or U7989 (N_7989,N_7375,N_7341);
xor U7990 (N_7990,N_7278,N_7309);
xor U7991 (N_7991,N_7456,N_7148);
or U7992 (N_7992,N_7279,N_7174);
and U7993 (N_7993,N_7418,N_7456);
or U7994 (N_7994,N_7210,N_7481);
nand U7995 (N_7995,N_7006,N_7123);
xnor U7996 (N_7996,N_7238,N_7209);
and U7997 (N_7997,N_7138,N_7396);
xor U7998 (N_7998,N_7143,N_7141);
and U7999 (N_7999,N_7356,N_7136);
or U8000 (N_8000,N_7559,N_7584);
and U8001 (N_8001,N_7526,N_7688);
xor U8002 (N_8002,N_7988,N_7921);
or U8003 (N_8003,N_7519,N_7621);
nand U8004 (N_8004,N_7969,N_7743);
and U8005 (N_8005,N_7539,N_7785);
or U8006 (N_8006,N_7847,N_7624);
xnor U8007 (N_8007,N_7843,N_7596);
and U8008 (N_8008,N_7855,N_7907);
and U8009 (N_8009,N_7853,N_7659);
xnor U8010 (N_8010,N_7990,N_7642);
nand U8011 (N_8011,N_7595,N_7657);
and U8012 (N_8012,N_7963,N_7766);
nand U8013 (N_8013,N_7927,N_7706);
or U8014 (N_8014,N_7972,N_7626);
xor U8015 (N_8015,N_7586,N_7506);
nor U8016 (N_8016,N_7793,N_7955);
xor U8017 (N_8017,N_7512,N_7958);
xor U8018 (N_8018,N_7560,N_7860);
xor U8019 (N_8019,N_7655,N_7938);
nand U8020 (N_8020,N_7720,N_7679);
or U8021 (N_8021,N_7827,N_7692);
nor U8022 (N_8022,N_7518,N_7825);
nor U8023 (N_8023,N_7664,N_7632);
or U8024 (N_8024,N_7856,N_7760);
xor U8025 (N_8025,N_7643,N_7630);
nand U8026 (N_8026,N_7635,N_7757);
nor U8027 (N_8027,N_7752,N_7895);
or U8028 (N_8028,N_7826,N_7590);
and U8029 (N_8029,N_7831,N_7984);
xnor U8030 (N_8030,N_7686,N_7604);
or U8031 (N_8031,N_7929,N_7603);
and U8032 (N_8032,N_7803,N_7607);
nand U8033 (N_8033,N_7501,N_7613);
and U8034 (N_8034,N_7934,N_7931);
or U8035 (N_8035,N_7978,N_7837);
nand U8036 (N_8036,N_7742,N_7776);
xnor U8037 (N_8037,N_7583,N_7858);
or U8038 (N_8038,N_7845,N_7571);
nor U8039 (N_8039,N_7730,N_7591);
xor U8040 (N_8040,N_7924,N_7939);
xor U8041 (N_8041,N_7817,N_7919);
nand U8042 (N_8042,N_7592,N_7581);
and U8043 (N_8043,N_7683,N_7649);
xnor U8044 (N_8044,N_7662,N_7541);
nand U8045 (N_8045,N_7995,N_7503);
nor U8046 (N_8046,N_7795,N_7648);
nand U8047 (N_8047,N_7734,N_7561);
xnor U8048 (N_8048,N_7891,N_7737);
xor U8049 (N_8049,N_7680,N_7703);
and U8050 (N_8050,N_7544,N_7770);
nor U8051 (N_8051,N_7666,N_7741);
xnor U8052 (N_8052,N_7677,N_7530);
and U8053 (N_8053,N_7773,N_7693);
nand U8054 (N_8054,N_7868,N_7510);
nor U8055 (N_8055,N_7925,N_7896);
nand U8056 (N_8056,N_7889,N_7521);
nor U8057 (N_8057,N_7728,N_7660);
nor U8058 (N_8058,N_7790,N_7698);
nand U8059 (N_8059,N_7517,N_7550);
and U8060 (N_8060,N_7876,N_7739);
nand U8061 (N_8061,N_7753,N_7951);
and U8062 (N_8062,N_7977,N_7610);
nor U8063 (N_8063,N_7534,N_7904);
xnor U8064 (N_8064,N_7552,N_7669);
and U8065 (N_8065,N_7736,N_7765);
nor U8066 (N_8066,N_7543,N_7614);
xnor U8067 (N_8067,N_7983,N_7522);
or U8068 (N_8068,N_7789,N_7898);
or U8069 (N_8069,N_7999,N_7818);
xnor U8070 (N_8070,N_7909,N_7771);
xor U8071 (N_8071,N_7875,N_7796);
nor U8072 (N_8072,N_7536,N_7641);
and U8073 (N_8073,N_7943,N_7717);
xor U8074 (N_8074,N_7574,N_7502);
nor U8075 (N_8075,N_7754,N_7707);
nor U8076 (N_8076,N_7869,N_7948);
xnor U8077 (N_8077,N_7525,N_7779);
nor U8078 (N_8078,N_7986,N_7528);
or U8079 (N_8079,N_7859,N_7578);
or U8080 (N_8080,N_7829,N_7886);
or U8081 (N_8081,N_7953,N_7663);
nand U8082 (N_8082,N_7968,N_7711);
nor U8083 (N_8083,N_7846,N_7874);
nor U8084 (N_8084,N_7775,N_7797);
and U8085 (N_8085,N_7533,N_7619);
nand U8086 (N_8086,N_7594,N_7638);
nand U8087 (N_8087,N_7637,N_7640);
nor U8088 (N_8088,N_7602,N_7567);
nor U8089 (N_8089,N_7598,N_7622);
or U8090 (N_8090,N_7933,N_7675);
nand U8091 (N_8091,N_7674,N_7993);
nand U8092 (N_8092,N_7917,N_7894);
and U8093 (N_8093,N_7836,N_7877);
or U8094 (N_8094,N_7850,N_7885);
xor U8095 (N_8095,N_7838,N_7722);
xor U8096 (N_8096,N_7940,N_7802);
nand U8097 (N_8097,N_7962,N_7961);
nand U8098 (N_8098,N_7918,N_7715);
nor U8099 (N_8099,N_7892,N_7806);
nand U8100 (N_8100,N_7794,N_7723);
nor U8101 (N_8101,N_7589,N_7758);
or U8102 (N_8102,N_7593,N_7769);
or U8103 (N_8103,N_7611,N_7937);
or U8104 (N_8104,N_7980,N_7672);
nand U8105 (N_8105,N_7947,N_7699);
and U8106 (N_8106,N_7970,N_7705);
xnor U8107 (N_8107,N_7587,N_7944);
and U8108 (N_8108,N_7982,N_7685);
nor U8109 (N_8109,N_7694,N_7799);
and U8110 (N_8110,N_7966,N_7879);
xnor U8111 (N_8111,N_7507,N_7744);
or U8112 (N_8112,N_7644,N_7971);
nand U8113 (N_8113,N_7609,N_7727);
xor U8114 (N_8114,N_7565,N_7628);
xnor U8115 (N_8115,N_7905,N_7992);
or U8116 (N_8116,N_7996,N_7652);
nor U8117 (N_8117,N_7661,N_7634);
nor U8118 (N_8118,N_7857,N_7945);
and U8119 (N_8119,N_7524,N_7973);
and U8120 (N_8120,N_7646,N_7665);
nor U8121 (N_8121,N_7941,N_7656);
or U8122 (N_8122,N_7805,N_7923);
nand U8123 (N_8123,N_7700,N_7513);
xor U8124 (N_8124,N_7515,N_7862);
or U8125 (N_8125,N_7920,N_7960);
or U8126 (N_8126,N_7801,N_7828);
xor U8127 (N_8127,N_7901,N_7788);
and U8128 (N_8128,N_7668,N_7936);
and U8129 (N_8129,N_7618,N_7822);
and U8130 (N_8130,N_7888,N_7952);
or U8131 (N_8131,N_7710,N_7819);
or U8132 (N_8132,N_7684,N_7562);
xor U8133 (N_8133,N_7508,N_7784);
or U8134 (N_8134,N_7865,N_7772);
or U8135 (N_8135,N_7697,N_7903);
or U8136 (N_8136,N_7570,N_7636);
xor U8137 (N_8137,N_7890,N_7712);
nand U8138 (N_8138,N_7946,N_7902);
xnor U8139 (N_8139,N_7912,N_7690);
nand U8140 (N_8140,N_7620,N_7568);
and U8141 (N_8141,N_7556,N_7516);
xor U8142 (N_8142,N_7523,N_7840);
or U8143 (N_8143,N_7732,N_7812);
or U8144 (N_8144,N_7884,N_7695);
xor U8145 (N_8145,N_7740,N_7658);
nand U8146 (N_8146,N_7748,N_7866);
and U8147 (N_8147,N_7849,N_7798);
xor U8148 (N_8148,N_7551,N_7792);
xor U8149 (N_8149,N_7554,N_7930);
nand U8150 (N_8150,N_7910,N_7815);
xor U8151 (N_8151,N_7500,N_7616);
or U8152 (N_8152,N_7639,N_7738);
and U8153 (N_8153,N_7670,N_7633);
or U8154 (N_8154,N_7735,N_7564);
nor U8155 (N_8155,N_7600,N_7957);
and U8156 (N_8156,N_7935,N_7509);
xor U8157 (N_8157,N_7881,N_7916);
nor U8158 (N_8158,N_7768,N_7749);
and U8159 (N_8159,N_7708,N_7914);
nor U8160 (N_8160,N_7667,N_7676);
and U8161 (N_8161,N_7804,N_7976);
nor U8162 (N_8162,N_7612,N_7725);
nand U8163 (N_8163,N_7867,N_7761);
nor U8164 (N_8164,N_7959,N_7553);
or U8165 (N_8165,N_7733,N_7535);
nand U8166 (N_8166,N_7580,N_7950);
nand U8167 (N_8167,N_7576,N_7780);
nand U8168 (N_8168,N_7650,N_7864);
xnor U8169 (N_8169,N_7702,N_7563);
or U8170 (N_8170,N_7608,N_7689);
or U8171 (N_8171,N_7900,N_7504);
or U8172 (N_8172,N_7540,N_7873);
or U8173 (N_8173,N_7954,N_7701);
or U8174 (N_8174,N_7747,N_7716);
xor U8175 (N_8175,N_7645,N_7691);
xor U8176 (N_8176,N_7994,N_7729);
nor U8177 (N_8177,N_7746,N_7520);
nor U8178 (N_8178,N_7572,N_7615);
nor U8179 (N_8179,N_7985,N_7719);
or U8180 (N_8180,N_7915,N_7908);
nand U8181 (N_8181,N_7721,N_7756);
xor U8182 (N_8182,N_7546,N_7820);
nand U8183 (N_8183,N_7991,N_7627);
xnor U8184 (N_8184,N_7835,N_7778);
nand U8185 (N_8185,N_7505,N_7841);
xnor U8186 (N_8186,N_7763,N_7678);
xor U8187 (N_8187,N_7605,N_7555);
nor U8188 (N_8188,N_7532,N_7870);
and U8189 (N_8189,N_7872,N_7582);
nand U8190 (N_8190,N_7871,N_7671);
and U8191 (N_8191,N_7852,N_7549);
nand U8192 (N_8192,N_7704,N_7511);
nor U8193 (N_8193,N_7979,N_7767);
nand U8194 (N_8194,N_7893,N_7844);
nor U8195 (N_8195,N_7623,N_7786);
nor U8196 (N_8196,N_7682,N_7588);
nor U8197 (N_8197,N_7751,N_7573);
and U8198 (N_8198,N_7724,N_7783);
nor U8199 (N_8199,N_7547,N_7809);
nand U8200 (N_8200,N_7687,N_7830);
xor U8201 (N_8201,N_7606,N_7601);
or U8202 (N_8202,N_7514,N_7949);
nand U8203 (N_8203,N_7529,N_7956);
or U8204 (N_8204,N_7597,N_7709);
xnor U8205 (N_8205,N_7777,N_7654);
and U8206 (N_8206,N_7527,N_7537);
nor U8207 (N_8207,N_7625,N_7851);
nor U8208 (N_8208,N_7926,N_7808);
nor U8209 (N_8209,N_7599,N_7782);
and U8210 (N_8210,N_7617,N_7651);
xnor U8211 (N_8211,N_7989,N_7755);
and U8212 (N_8212,N_7807,N_7913);
or U8213 (N_8213,N_7883,N_7897);
or U8214 (N_8214,N_7631,N_7545);
or U8215 (N_8215,N_7629,N_7987);
nand U8216 (N_8216,N_7557,N_7653);
xnor U8217 (N_8217,N_7811,N_7942);
and U8218 (N_8218,N_7928,N_7713);
nand U8219 (N_8219,N_7774,N_7899);
or U8220 (N_8220,N_7575,N_7731);
and U8221 (N_8221,N_7854,N_7696);
nand U8222 (N_8222,N_7566,N_7832);
or U8223 (N_8223,N_7548,N_7558);
and U8224 (N_8224,N_7882,N_7781);
xnor U8225 (N_8225,N_7823,N_7647);
and U8226 (N_8226,N_7878,N_7810);
or U8227 (N_8227,N_7759,N_7764);
nand U8228 (N_8228,N_7911,N_7967);
xor U8229 (N_8229,N_7814,N_7718);
or U8230 (N_8230,N_7861,N_7998);
or U8231 (N_8231,N_7800,N_7842);
and U8232 (N_8232,N_7863,N_7714);
xor U8233 (N_8233,N_7922,N_7932);
xor U8234 (N_8234,N_7821,N_7813);
xor U8235 (N_8235,N_7585,N_7762);
and U8236 (N_8236,N_7964,N_7569);
nand U8237 (N_8237,N_7975,N_7974);
or U8238 (N_8238,N_7997,N_7745);
nand U8239 (N_8239,N_7906,N_7681);
nand U8240 (N_8240,N_7839,N_7816);
xnor U8241 (N_8241,N_7538,N_7579);
nor U8242 (N_8242,N_7880,N_7531);
xnor U8243 (N_8243,N_7787,N_7834);
nand U8244 (N_8244,N_7887,N_7824);
nor U8245 (N_8245,N_7542,N_7833);
and U8246 (N_8246,N_7791,N_7848);
nand U8247 (N_8247,N_7673,N_7577);
and U8248 (N_8248,N_7981,N_7750);
nor U8249 (N_8249,N_7965,N_7726);
nor U8250 (N_8250,N_7706,N_7909);
nor U8251 (N_8251,N_7794,N_7529);
nand U8252 (N_8252,N_7871,N_7864);
nand U8253 (N_8253,N_7724,N_7558);
or U8254 (N_8254,N_7639,N_7592);
and U8255 (N_8255,N_7771,N_7887);
and U8256 (N_8256,N_7549,N_7693);
xor U8257 (N_8257,N_7901,N_7584);
nand U8258 (N_8258,N_7656,N_7814);
xnor U8259 (N_8259,N_7893,N_7688);
nor U8260 (N_8260,N_7677,N_7557);
and U8261 (N_8261,N_7592,N_7813);
and U8262 (N_8262,N_7568,N_7582);
nor U8263 (N_8263,N_7587,N_7809);
nor U8264 (N_8264,N_7995,N_7622);
nor U8265 (N_8265,N_7545,N_7828);
nand U8266 (N_8266,N_7667,N_7863);
nor U8267 (N_8267,N_7584,N_7678);
nor U8268 (N_8268,N_7980,N_7790);
and U8269 (N_8269,N_7716,N_7759);
nand U8270 (N_8270,N_7986,N_7864);
nand U8271 (N_8271,N_7776,N_7615);
or U8272 (N_8272,N_7616,N_7928);
nor U8273 (N_8273,N_7655,N_7669);
nand U8274 (N_8274,N_7649,N_7700);
xnor U8275 (N_8275,N_7633,N_7616);
xor U8276 (N_8276,N_7794,N_7670);
nand U8277 (N_8277,N_7929,N_7932);
xnor U8278 (N_8278,N_7895,N_7595);
or U8279 (N_8279,N_7976,N_7519);
nor U8280 (N_8280,N_7636,N_7832);
xnor U8281 (N_8281,N_7506,N_7571);
or U8282 (N_8282,N_7854,N_7820);
nand U8283 (N_8283,N_7929,N_7806);
xnor U8284 (N_8284,N_7925,N_7542);
nand U8285 (N_8285,N_7808,N_7873);
and U8286 (N_8286,N_7539,N_7900);
and U8287 (N_8287,N_7582,N_7668);
and U8288 (N_8288,N_7637,N_7975);
nand U8289 (N_8289,N_7539,N_7724);
nand U8290 (N_8290,N_7528,N_7826);
xnor U8291 (N_8291,N_7589,N_7937);
nor U8292 (N_8292,N_7900,N_7808);
nand U8293 (N_8293,N_7916,N_7828);
xnor U8294 (N_8294,N_7827,N_7862);
and U8295 (N_8295,N_7952,N_7594);
nor U8296 (N_8296,N_7517,N_7623);
and U8297 (N_8297,N_7664,N_7734);
xor U8298 (N_8298,N_7903,N_7642);
and U8299 (N_8299,N_7554,N_7820);
nand U8300 (N_8300,N_7770,N_7599);
nand U8301 (N_8301,N_7769,N_7784);
and U8302 (N_8302,N_7719,N_7727);
and U8303 (N_8303,N_7985,N_7708);
nand U8304 (N_8304,N_7704,N_7715);
or U8305 (N_8305,N_7725,N_7520);
xor U8306 (N_8306,N_7525,N_7798);
and U8307 (N_8307,N_7717,N_7687);
nand U8308 (N_8308,N_7947,N_7726);
nand U8309 (N_8309,N_7982,N_7535);
or U8310 (N_8310,N_7542,N_7706);
nand U8311 (N_8311,N_7860,N_7792);
xnor U8312 (N_8312,N_7924,N_7991);
and U8313 (N_8313,N_7899,N_7834);
nand U8314 (N_8314,N_7732,N_7783);
or U8315 (N_8315,N_7815,N_7895);
xnor U8316 (N_8316,N_7981,N_7893);
and U8317 (N_8317,N_7642,N_7779);
nor U8318 (N_8318,N_7594,N_7899);
and U8319 (N_8319,N_7839,N_7587);
xor U8320 (N_8320,N_7712,N_7583);
xor U8321 (N_8321,N_7617,N_7600);
nand U8322 (N_8322,N_7548,N_7504);
or U8323 (N_8323,N_7629,N_7686);
nor U8324 (N_8324,N_7842,N_7965);
nor U8325 (N_8325,N_7597,N_7969);
or U8326 (N_8326,N_7723,N_7790);
or U8327 (N_8327,N_7676,N_7733);
xnor U8328 (N_8328,N_7530,N_7587);
nand U8329 (N_8329,N_7898,N_7727);
or U8330 (N_8330,N_7760,N_7511);
nand U8331 (N_8331,N_7983,N_7887);
nor U8332 (N_8332,N_7605,N_7779);
xor U8333 (N_8333,N_7810,N_7589);
xnor U8334 (N_8334,N_7837,N_7952);
and U8335 (N_8335,N_7935,N_7627);
or U8336 (N_8336,N_7892,N_7580);
xnor U8337 (N_8337,N_7854,N_7643);
nor U8338 (N_8338,N_7573,N_7858);
nand U8339 (N_8339,N_7722,N_7931);
nand U8340 (N_8340,N_7661,N_7859);
and U8341 (N_8341,N_7518,N_7756);
and U8342 (N_8342,N_7772,N_7877);
nor U8343 (N_8343,N_7602,N_7865);
xnor U8344 (N_8344,N_7831,N_7998);
or U8345 (N_8345,N_7624,N_7511);
nand U8346 (N_8346,N_7774,N_7945);
and U8347 (N_8347,N_7866,N_7843);
xor U8348 (N_8348,N_7617,N_7813);
or U8349 (N_8349,N_7919,N_7946);
nand U8350 (N_8350,N_7671,N_7938);
or U8351 (N_8351,N_7891,N_7924);
and U8352 (N_8352,N_7822,N_7827);
and U8353 (N_8353,N_7684,N_7849);
nor U8354 (N_8354,N_7544,N_7577);
nand U8355 (N_8355,N_7691,N_7883);
or U8356 (N_8356,N_7790,N_7511);
nand U8357 (N_8357,N_7606,N_7872);
or U8358 (N_8358,N_7644,N_7841);
nor U8359 (N_8359,N_7886,N_7839);
or U8360 (N_8360,N_7999,N_7813);
nor U8361 (N_8361,N_7667,N_7959);
or U8362 (N_8362,N_7661,N_7919);
and U8363 (N_8363,N_7755,N_7714);
nand U8364 (N_8364,N_7950,N_7836);
and U8365 (N_8365,N_7850,N_7743);
and U8366 (N_8366,N_7866,N_7523);
xnor U8367 (N_8367,N_7765,N_7669);
or U8368 (N_8368,N_7660,N_7851);
xor U8369 (N_8369,N_7537,N_7778);
or U8370 (N_8370,N_7630,N_7580);
and U8371 (N_8371,N_7939,N_7860);
or U8372 (N_8372,N_7935,N_7732);
or U8373 (N_8373,N_7695,N_7886);
nor U8374 (N_8374,N_7660,N_7692);
xnor U8375 (N_8375,N_7716,N_7500);
or U8376 (N_8376,N_7562,N_7641);
nand U8377 (N_8377,N_7802,N_7862);
nand U8378 (N_8378,N_7657,N_7758);
nand U8379 (N_8379,N_7536,N_7911);
xor U8380 (N_8380,N_7734,N_7922);
and U8381 (N_8381,N_7752,N_7933);
nand U8382 (N_8382,N_7533,N_7890);
and U8383 (N_8383,N_7739,N_7632);
nand U8384 (N_8384,N_7776,N_7700);
nor U8385 (N_8385,N_7570,N_7523);
xnor U8386 (N_8386,N_7902,N_7665);
or U8387 (N_8387,N_7545,N_7718);
nand U8388 (N_8388,N_7590,N_7810);
xnor U8389 (N_8389,N_7881,N_7858);
nand U8390 (N_8390,N_7648,N_7529);
nand U8391 (N_8391,N_7863,N_7825);
xnor U8392 (N_8392,N_7819,N_7812);
nor U8393 (N_8393,N_7977,N_7891);
nand U8394 (N_8394,N_7790,N_7719);
and U8395 (N_8395,N_7502,N_7819);
or U8396 (N_8396,N_7544,N_7775);
and U8397 (N_8397,N_7930,N_7949);
and U8398 (N_8398,N_7849,N_7569);
nand U8399 (N_8399,N_7620,N_7764);
xnor U8400 (N_8400,N_7521,N_7695);
or U8401 (N_8401,N_7774,N_7534);
xnor U8402 (N_8402,N_7827,N_7646);
and U8403 (N_8403,N_7529,N_7672);
nand U8404 (N_8404,N_7820,N_7561);
nor U8405 (N_8405,N_7974,N_7902);
or U8406 (N_8406,N_7515,N_7870);
xor U8407 (N_8407,N_7631,N_7763);
xor U8408 (N_8408,N_7695,N_7830);
xnor U8409 (N_8409,N_7856,N_7947);
or U8410 (N_8410,N_7650,N_7774);
and U8411 (N_8411,N_7606,N_7721);
xnor U8412 (N_8412,N_7671,N_7772);
and U8413 (N_8413,N_7554,N_7534);
xor U8414 (N_8414,N_7999,N_7854);
or U8415 (N_8415,N_7612,N_7539);
xor U8416 (N_8416,N_7658,N_7617);
xnor U8417 (N_8417,N_7622,N_7645);
and U8418 (N_8418,N_7554,N_7528);
and U8419 (N_8419,N_7943,N_7910);
xnor U8420 (N_8420,N_7803,N_7911);
or U8421 (N_8421,N_7777,N_7753);
nor U8422 (N_8422,N_7773,N_7893);
or U8423 (N_8423,N_7684,N_7688);
and U8424 (N_8424,N_7506,N_7595);
xor U8425 (N_8425,N_7541,N_7572);
and U8426 (N_8426,N_7837,N_7856);
xor U8427 (N_8427,N_7867,N_7643);
or U8428 (N_8428,N_7726,N_7715);
and U8429 (N_8429,N_7899,N_7698);
nand U8430 (N_8430,N_7633,N_7927);
xor U8431 (N_8431,N_7672,N_7716);
and U8432 (N_8432,N_7815,N_7921);
or U8433 (N_8433,N_7539,N_7672);
or U8434 (N_8434,N_7735,N_7512);
and U8435 (N_8435,N_7819,N_7632);
nand U8436 (N_8436,N_7947,N_7734);
nand U8437 (N_8437,N_7593,N_7558);
xnor U8438 (N_8438,N_7744,N_7655);
or U8439 (N_8439,N_7778,N_7641);
and U8440 (N_8440,N_7686,N_7783);
nor U8441 (N_8441,N_7626,N_7870);
nor U8442 (N_8442,N_7576,N_7817);
nor U8443 (N_8443,N_7797,N_7714);
nor U8444 (N_8444,N_7986,N_7784);
and U8445 (N_8445,N_7828,N_7565);
nor U8446 (N_8446,N_7731,N_7789);
or U8447 (N_8447,N_7578,N_7939);
or U8448 (N_8448,N_7537,N_7597);
nor U8449 (N_8449,N_7611,N_7930);
nand U8450 (N_8450,N_7804,N_7523);
nand U8451 (N_8451,N_7629,N_7537);
and U8452 (N_8452,N_7904,N_7943);
and U8453 (N_8453,N_7750,N_7895);
and U8454 (N_8454,N_7656,N_7803);
nor U8455 (N_8455,N_7949,N_7543);
and U8456 (N_8456,N_7829,N_7838);
nand U8457 (N_8457,N_7934,N_7671);
or U8458 (N_8458,N_7875,N_7569);
and U8459 (N_8459,N_7903,N_7739);
xor U8460 (N_8460,N_7902,N_7699);
nor U8461 (N_8461,N_7512,N_7951);
nor U8462 (N_8462,N_7855,N_7771);
and U8463 (N_8463,N_7645,N_7604);
and U8464 (N_8464,N_7679,N_7670);
nor U8465 (N_8465,N_7780,N_7897);
xor U8466 (N_8466,N_7797,N_7839);
nor U8467 (N_8467,N_7592,N_7655);
nor U8468 (N_8468,N_7901,N_7607);
nand U8469 (N_8469,N_7766,N_7943);
or U8470 (N_8470,N_7736,N_7674);
nor U8471 (N_8471,N_7891,N_7535);
nand U8472 (N_8472,N_7554,N_7737);
nor U8473 (N_8473,N_7732,N_7501);
xnor U8474 (N_8474,N_7636,N_7544);
and U8475 (N_8475,N_7603,N_7538);
or U8476 (N_8476,N_7626,N_7577);
nor U8477 (N_8477,N_7778,N_7644);
xnor U8478 (N_8478,N_7535,N_7996);
xnor U8479 (N_8479,N_7762,N_7941);
nor U8480 (N_8480,N_7758,N_7679);
nand U8481 (N_8481,N_7546,N_7630);
and U8482 (N_8482,N_7572,N_7549);
nor U8483 (N_8483,N_7924,N_7797);
and U8484 (N_8484,N_7687,N_7915);
nand U8485 (N_8485,N_7685,N_7785);
and U8486 (N_8486,N_7746,N_7531);
nand U8487 (N_8487,N_7843,N_7884);
nor U8488 (N_8488,N_7857,N_7962);
nand U8489 (N_8489,N_7639,N_7999);
or U8490 (N_8490,N_7835,N_7745);
xor U8491 (N_8491,N_7769,N_7915);
xor U8492 (N_8492,N_7988,N_7687);
and U8493 (N_8493,N_7611,N_7763);
and U8494 (N_8494,N_7569,N_7793);
nand U8495 (N_8495,N_7525,N_7894);
and U8496 (N_8496,N_7795,N_7556);
or U8497 (N_8497,N_7916,N_7550);
and U8498 (N_8498,N_7861,N_7558);
nor U8499 (N_8499,N_7570,N_7771);
and U8500 (N_8500,N_8284,N_8311);
or U8501 (N_8501,N_8169,N_8058);
and U8502 (N_8502,N_8033,N_8130);
xor U8503 (N_8503,N_8466,N_8011);
nor U8504 (N_8504,N_8110,N_8316);
nor U8505 (N_8505,N_8382,N_8159);
nor U8506 (N_8506,N_8376,N_8264);
nand U8507 (N_8507,N_8137,N_8030);
and U8508 (N_8508,N_8401,N_8411);
xnor U8509 (N_8509,N_8226,N_8420);
xor U8510 (N_8510,N_8083,N_8002);
xor U8511 (N_8511,N_8131,N_8270);
nor U8512 (N_8512,N_8409,N_8414);
or U8513 (N_8513,N_8079,N_8357);
nor U8514 (N_8514,N_8475,N_8190);
nor U8515 (N_8515,N_8218,N_8071);
nand U8516 (N_8516,N_8108,N_8305);
and U8517 (N_8517,N_8047,N_8326);
or U8518 (N_8518,N_8034,N_8297);
or U8519 (N_8519,N_8049,N_8486);
nand U8520 (N_8520,N_8201,N_8118);
or U8521 (N_8521,N_8280,N_8374);
and U8522 (N_8522,N_8439,N_8485);
nand U8523 (N_8523,N_8246,N_8199);
xnor U8524 (N_8524,N_8082,N_8333);
nor U8525 (N_8525,N_8105,N_8360);
xnor U8526 (N_8526,N_8327,N_8153);
and U8527 (N_8527,N_8278,N_8061);
xnor U8528 (N_8528,N_8286,N_8216);
and U8529 (N_8529,N_8234,N_8000);
nand U8530 (N_8530,N_8174,N_8152);
xor U8531 (N_8531,N_8455,N_8309);
or U8532 (N_8532,N_8390,N_8472);
or U8533 (N_8533,N_8410,N_8233);
and U8534 (N_8534,N_8255,N_8138);
or U8535 (N_8535,N_8340,N_8194);
nand U8536 (N_8536,N_8303,N_8171);
and U8537 (N_8537,N_8059,N_8368);
and U8538 (N_8538,N_8039,N_8249);
or U8539 (N_8539,N_8408,N_8349);
xnor U8540 (N_8540,N_8282,N_8175);
and U8541 (N_8541,N_8307,N_8447);
and U8542 (N_8542,N_8165,N_8170);
and U8543 (N_8543,N_8470,N_8177);
or U8544 (N_8544,N_8172,N_8224);
xor U8545 (N_8545,N_8151,N_8457);
or U8546 (N_8546,N_8413,N_8210);
nand U8547 (N_8547,N_8028,N_8239);
and U8548 (N_8548,N_8375,N_8240);
nand U8549 (N_8549,N_8492,N_8302);
nand U8550 (N_8550,N_8022,N_8109);
or U8551 (N_8551,N_8162,N_8188);
and U8552 (N_8552,N_8250,N_8460);
xor U8553 (N_8553,N_8356,N_8057);
nor U8554 (N_8554,N_8098,N_8388);
nand U8555 (N_8555,N_8236,N_8317);
xor U8556 (N_8556,N_8383,N_8001);
or U8557 (N_8557,N_8352,N_8467);
nor U8558 (N_8558,N_8436,N_8180);
or U8559 (N_8559,N_8417,N_8362);
xnor U8560 (N_8560,N_8018,N_8148);
xor U8561 (N_8561,N_8269,N_8381);
and U8562 (N_8562,N_8456,N_8046);
nor U8563 (N_8563,N_8244,N_8115);
nand U8564 (N_8564,N_8281,N_8013);
and U8565 (N_8565,N_8335,N_8154);
nand U8566 (N_8566,N_8418,N_8076);
nand U8567 (N_8567,N_8161,N_8331);
or U8568 (N_8568,N_8396,N_8009);
or U8569 (N_8569,N_8443,N_8119);
or U8570 (N_8570,N_8142,N_8363);
and U8571 (N_8571,N_8067,N_8050);
nor U8572 (N_8572,N_8095,N_8123);
nand U8573 (N_8573,N_8181,N_8310);
and U8574 (N_8574,N_8484,N_8193);
or U8575 (N_8575,N_8025,N_8279);
and U8576 (N_8576,N_8112,N_8160);
nand U8577 (N_8577,N_8451,N_8043);
nor U8578 (N_8578,N_8425,N_8196);
nand U8579 (N_8579,N_8394,N_8256);
nor U8580 (N_8580,N_8008,N_8386);
nor U8581 (N_8581,N_8052,N_8415);
nor U8582 (N_8582,N_8324,N_8321);
nand U8583 (N_8583,N_8041,N_8191);
nand U8584 (N_8584,N_8145,N_8441);
nor U8585 (N_8585,N_8406,N_8107);
nand U8586 (N_8586,N_8100,N_8099);
xnor U8587 (N_8587,N_8312,N_8035);
nand U8588 (N_8588,N_8068,N_8176);
xor U8589 (N_8589,N_8274,N_8481);
nand U8590 (N_8590,N_8392,N_8208);
nand U8591 (N_8591,N_8084,N_8446);
nor U8592 (N_8592,N_8200,N_8010);
nor U8593 (N_8593,N_8081,N_8277);
xnor U8594 (N_8594,N_8351,N_8487);
and U8595 (N_8595,N_8393,N_8053);
nor U8596 (N_8596,N_8319,N_8021);
nor U8597 (N_8597,N_8135,N_8299);
nand U8598 (N_8598,N_8207,N_8213);
nor U8599 (N_8599,N_8495,N_8065);
xor U8600 (N_8600,N_8354,N_8449);
xor U8601 (N_8601,N_8294,N_8254);
xnor U8602 (N_8602,N_8498,N_8285);
and U8603 (N_8603,N_8214,N_8132);
or U8604 (N_8604,N_8347,N_8399);
xor U8605 (N_8605,N_8404,N_8163);
xor U8606 (N_8606,N_8229,N_8044);
nand U8607 (N_8607,N_8377,N_8471);
and U8608 (N_8608,N_8045,N_8124);
nor U8609 (N_8609,N_8345,N_8338);
xor U8610 (N_8610,N_8243,N_8267);
and U8611 (N_8611,N_8221,N_8339);
nor U8612 (N_8612,N_8343,N_8150);
nor U8613 (N_8613,N_8007,N_8004);
and U8614 (N_8614,N_8231,N_8320);
nor U8615 (N_8615,N_8093,N_8038);
xnor U8616 (N_8616,N_8295,N_8440);
nand U8617 (N_8617,N_8097,N_8230);
nand U8618 (N_8618,N_8369,N_8155);
or U8619 (N_8619,N_8266,N_8265);
or U8620 (N_8620,N_8127,N_8276);
xnor U8621 (N_8621,N_8334,N_8458);
nor U8622 (N_8622,N_8330,N_8087);
xor U8623 (N_8623,N_8168,N_8085);
or U8624 (N_8624,N_8419,N_8431);
and U8625 (N_8625,N_8006,N_8158);
nor U8626 (N_8626,N_8227,N_8074);
and U8627 (N_8627,N_8062,N_8157);
or U8628 (N_8628,N_8016,N_8423);
and U8629 (N_8629,N_8070,N_8206);
nand U8630 (N_8630,N_8156,N_8003);
or U8631 (N_8631,N_8042,N_8040);
nor U8632 (N_8632,N_8017,N_8198);
xnor U8633 (N_8633,N_8433,N_8477);
or U8634 (N_8634,N_8427,N_8189);
nor U8635 (N_8635,N_8064,N_8453);
nor U8636 (N_8636,N_8090,N_8140);
nor U8637 (N_8637,N_8048,N_8219);
and U8638 (N_8638,N_8054,N_8459);
nor U8639 (N_8639,N_8407,N_8027);
nand U8640 (N_8640,N_8091,N_8461);
xor U8641 (N_8641,N_8397,N_8126);
nand U8642 (N_8642,N_8032,N_8251);
xnor U8643 (N_8643,N_8232,N_8121);
nand U8644 (N_8644,N_8204,N_8488);
xor U8645 (N_8645,N_8426,N_8092);
nand U8646 (N_8646,N_8350,N_8403);
nand U8647 (N_8647,N_8480,N_8066);
or U8648 (N_8648,N_8257,N_8183);
nand U8649 (N_8649,N_8104,N_8454);
and U8650 (N_8650,N_8179,N_8385);
nand U8651 (N_8651,N_8308,N_8117);
nor U8652 (N_8652,N_8103,N_8056);
nand U8653 (N_8653,N_8372,N_8258);
nand U8654 (N_8654,N_8078,N_8400);
nand U8655 (N_8655,N_8075,N_8490);
nor U8656 (N_8656,N_8149,N_8398);
nand U8657 (N_8657,N_8370,N_8434);
nand U8658 (N_8658,N_8102,N_8187);
or U8659 (N_8659,N_8186,N_8055);
and U8660 (N_8660,N_8364,N_8291);
xnor U8661 (N_8661,N_8217,N_8469);
nand U8662 (N_8662,N_8012,N_8205);
xor U8663 (N_8663,N_8342,N_8337);
xor U8664 (N_8664,N_8445,N_8318);
or U8665 (N_8665,N_8479,N_8476);
xor U8666 (N_8666,N_8432,N_8086);
xor U8667 (N_8667,N_8468,N_8391);
nor U8668 (N_8668,N_8366,N_8422);
nand U8669 (N_8669,N_8300,N_8080);
nand U8670 (N_8670,N_8273,N_8379);
or U8671 (N_8671,N_8405,N_8228);
nand U8672 (N_8672,N_8139,N_8128);
or U8673 (N_8673,N_8106,N_8212);
nor U8674 (N_8674,N_8353,N_8395);
nand U8675 (N_8675,N_8144,N_8164);
xnor U8676 (N_8676,N_8125,N_8314);
or U8677 (N_8677,N_8328,N_8336);
and U8678 (N_8678,N_8329,N_8129);
nand U8679 (N_8679,N_8024,N_8088);
nor U8680 (N_8680,N_8195,N_8094);
xor U8681 (N_8681,N_8489,N_8442);
xor U8682 (N_8682,N_8421,N_8373);
nand U8683 (N_8683,N_8346,N_8323);
xnor U8684 (N_8684,N_8167,N_8192);
nand U8685 (N_8685,N_8037,N_8301);
or U8686 (N_8686,N_8253,N_8245);
xor U8687 (N_8687,N_8252,N_8332);
or U8688 (N_8688,N_8452,N_8378);
nor U8689 (N_8689,N_8412,N_8499);
nand U8690 (N_8690,N_8133,N_8304);
xor U8691 (N_8691,N_8387,N_8268);
or U8692 (N_8692,N_8435,N_8497);
xor U8693 (N_8693,N_8341,N_8325);
nor U8694 (N_8694,N_8113,N_8122);
or U8695 (N_8695,N_8361,N_8178);
nor U8696 (N_8696,N_8429,N_8315);
xor U8697 (N_8697,N_8272,N_8073);
nor U8698 (N_8698,N_8464,N_8197);
nor U8699 (N_8699,N_8344,N_8023);
nand U8700 (N_8700,N_8348,N_8225);
nor U8701 (N_8701,N_8051,N_8215);
or U8702 (N_8702,N_8029,N_8494);
or U8703 (N_8703,N_8120,N_8491);
nor U8704 (N_8704,N_8202,N_8203);
nor U8705 (N_8705,N_8298,N_8211);
nand U8706 (N_8706,N_8237,N_8288);
and U8707 (N_8707,N_8096,N_8367);
nor U8708 (N_8708,N_8444,N_8262);
or U8709 (N_8709,N_8241,N_8146);
xor U8710 (N_8710,N_8292,N_8063);
xor U8711 (N_8711,N_8166,N_8290);
or U8712 (N_8712,N_8060,N_8283);
and U8713 (N_8713,N_8293,N_8474);
nor U8714 (N_8714,N_8136,N_8259);
or U8715 (N_8715,N_8371,N_8384);
and U8716 (N_8716,N_8141,N_8380);
nand U8717 (N_8717,N_8275,N_8020);
nand U8718 (N_8718,N_8365,N_8069);
and U8719 (N_8719,N_8465,N_8263);
or U8720 (N_8720,N_8359,N_8306);
and U8721 (N_8721,N_8182,N_8242);
nand U8722 (N_8722,N_8185,N_8089);
nand U8723 (N_8723,N_8478,N_8116);
nor U8724 (N_8724,N_8111,N_8031);
or U8725 (N_8725,N_8438,N_8313);
and U8726 (N_8726,N_8261,N_8271);
nor U8727 (N_8727,N_8462,N_8222);
xor U8728 (N_8728,N_8019,N_8238);
nor U8729 (N_8729,N_8450,N_8026);
nor U8730 (N_8730,N_8184,N_8463);
nor U8731 (N_8731,N_8289,N_8260);
or U8732 (N_8732,N_8114,N_8014);
xnor U8733 (N_8733,N_8358,N_8296);
xor U8734 (N_8734,N_8437,N_8424);
or U8735 (N_8735,N_8287,N_8430);
nand U8736 (N_8736,N_8483,N_8248);
xor U8737 (N_8737,N_8209,N_8005);
nor U8738 (N_8738,N_8247,N_8173);
or U8739 (N_8739,N_8322,N_8235);
and U8740 (N_8740,N_8220,N_8072);
nand U8741 (N_8741,N_8473,N_8077);
nand U8742 (N_8742,N_8101,N_8496);
nor U8743 (N_8743,N_8355,N_8428);
or U8744 (N_8744,N_8416,N_8134);
nor U8745 (N_8745,N_8147,N_8493);
xnor U8746 (N_8746,N_8143,N_8036);
nand U8747 (N_8747,N_8389,N_8448);
nand U8748 (N_8748,N_8223,N_8482);
nand U8749 (N_8749,N_8402,N_8015);
nand U8750 (N_8750,N_8060,N_8437);
nor U8751 (N_8751,N_8471,N_8249);
nand U8752 (N_8752,N_8294,N_8061);
nand U8753 (N_8753,N_8360,N_8086);
and U8754 (N_8754,N_8406,N_8475);
nand U8755 (N_8755,N_8125,N_8425);
nand U8756 (N_8756,N_8054,N_8436);
nand U8757 (N_8757,N_8009,N_8354);
nor U8758 (N_8758,N_8444,N_8240);
nor U8759 (N_8759,N_8108,N_8475);
xnor U8760 (N_8760,N_8335,N_8486);
nor U8761 (N_8761,N_8259,N_8409);
nor U8762 (N_8762,N_8041,N_8198);
nor U8763 (N_8763,N_8332,N_8487);
or U8764 (N_8764,N_8135,N_8104);
and U8765 (N_8765,N_8398,N_8092);
nand U8766 (N_8766,N_8316,N_8409);
or U8767 (N_8767,N_8157,N_8195);
nand U8768 (N_8768,N_8030,N_8247);
or U8769 (N_8769,N_8107,N_8353);
xnor U8770 (N_8770,N_8147,N_8486);
or U8771 (N_8771,N_8482,N_8392);
xnor U8772 (N_8772,N_8325,N_8247);
nand U8773 (N_8773,N_8173,N_8096);
and U8774 (N_8774,N_8305,N_8340);
and U8775 (N_8775,N_8393,N_8182);
xnor U8776 (N_8776,N_8497,N_8228);
or U8777 (N_8777,N_8031,N_8210);
nor U8778 (N_8778,N_8076,N_8222);
or U8779 (N_8779,N_8283,N_8155);
and U8780 (N_8780,N_8400,N_8004);
or U8781 (N_8781,N_8249,N_8486);
and U8782 (N_8782,N_8480,N_8095);
xor U8783 (N_8783,N_8334,N_8379);
nor U8784 (N_8784,N_8054,N_8453);
nand U8785 (N_8785,N_8260,N_8464);
or U8786 (N_8786,N_8088,N_8406);
xnor U8787 (N_8787,N_8019,N_8316);
nand U8788 (N_8788,N_8267,N_8273);
or U8789 (N_8789,N_8481,N_8069);
xor U8790 (N_8790,N_8319,N_8354);
or U8791 (N_8791,N_8016,N_8115);
nor U8792 (N_8792,N_8057,N_8288);
or U8793 (N_8793,N_8283,N_8062);
nand U8794 (N_8794,N_8337,N_8478);
xnor U8795 (N_8795,N_8205,N_8226);
xnor U8796 (N_8796,N_8382,N_8303);
xnor U8797 (N_8797,N_8092,N_8046);
xnor U8798 (N_8798,N_8397,N_8065);
or U8799 (N_8799,N_8282,N_8465);
or U8800 (N_8800,N_8301,N_8463);
xor U8801 (N_8801,N_8323,N_8197);
nand U8802 (N_8802,N_8069,N_8160);
xor U8803 (N_8803,N_8156,N_8162);
xor U8804 (N_8804,N_8411,N_8494);
or U8805 (N_8805,N_8446,N_8431);
or U8806 (N_8806,N_8429,N_8469);
xnor U8807 (N_8807,N_8133,N_8277);
nand U8808 (N_8808,N_8432,N_8349);
nor U8809 (N_8809,N_8170,N_8038);
xor U8810 (N_8810,N_8353,N_8135);
and U8811 (N_8811,N_8237,N_8052);
nor U8812 (N_8812,N_8239,N_8338);
and U8813 (N_8813,N_8434,N_8060);
nand U8814 (N_8814,N_8339,N_8426);
nand U8815 (N_8815,N_8396,N_8326);
nor U8816 (N_8816,N_8316,N_8125);
or U8817 (N_8817,N_8145,N_8380);
or U8818 (N_8818,N_8136,N_8396);
or U8819 (N_8819,N_8199,N_8457);
nor U8820 (N_8820,N_8441,N_8015);
xor U8821 (N_8821,N_8282,N_8131);
xor U8822 (N_8822,N_8004,N_8062);
xnor U8823 (N_8823,N_8256,N_8090);
and U8824 (N_8824,N_8315,N_8246);
or U8825 (N_8825,N_8006,N_8464);
nand U8826 (N_8826,N_8365,N_8003);
xnor U8827 (N_8827,N_8036,N_8482);
xnor U8828 (N_8828,N_8210,N_8411);
nor U8829 (N_8829,N_8485,N_8035);
or U8830 (N_8830,N_8172,N_8236);
xor U8831 (N_8831,N_8359,N_8131);
nor U8832 (N_8832,N_8397,N_8336);
xor U8833 (N_8833,N_8195,N_8065);
or U8834 (N_8834,N_8069,N_8197);
nor U8835 (N_8835,N_8208,N_8323);
or U8836 (N_8836,N_8415,N_8186);
or U8837 (N_8837,N_8348,N_8441);
nor U8838 (N_8838,N_8134,N_8201);
xor U8839 (N_8839,N_8152,N_8347);
and U8840 (N_8840,N_8200,N_8227);
xnor U8841 (N_8841,N_8416,N_8271);
xnor U8842 (N_8842,N_8347,N_8472);
nand U8843 (N_8843,N_8415,N_8244);
and U8844 (N_8844,N_8103,N_8102);
and U8845 (N_8845,N_8446,N_8126);
xnor U8846 (N_8846,N_8471,N_8334);
nor U8847 (N_8847,N_8113,N_8207);
and U8848 (N_8848,N_8233,N_8091);
xor U8849 (N_8849,N_8300,N_8352);
or U8850 (N_8850,N_8129,N_8131);
nand U8851 (N_8851,N_8202,N_8186);
nor U8852 (N_8852,N_8103,N_8066);
and U8853 (N_8853,N_8155,N_8214);
or U8854 (N_8854,N_8039,N_8272);
or U8855 (N_8855,N_8463,N_8133);
nand U8856 (N_8856,N_8386,N_8385);
xor U8857 (N_8857,N_8216,N_8471);
nand U8858 (N_8858,N_8270,N_8115);
xnor U8859 (N_8859,N_8333,N_8394);
and U8860 (N_8860,N_8446,N_8066);
nor U8861 (N_8861,N_8104,N_8285);
nand U8862 (N_8862,N_8411,N_8324);
and U8863 (N_8863,N_8219,N_8266);
or U8864 (N_8864,N_8388,N_8143);
or U8865 (N_8865,N_8003,N_8285);
nand U8866 (N_8866,N_8172,N_8019);
nand U8867 (N_8867,N_8254,N_8044);
nand U8868 (N_8868,N_8013,N_8047);
nor U8869 (N_8869,N_8153,N_8413);
nand U8870 (N_8870,N_8487,N_8030);
nor U8871 (N_8871,N_8198,N_8386);
nand U8872 (N_8872,N_8166,N_8432);
xor U8873 (N_8873,N_8100,N_8440);
or U8874 (N_8874,N_8108,N_8231);
xnor U8875 (N_8875,N_8236,N_8352);
nor U8876 (N_8876,N_8314,N_8218);
or U8877 (N_8877,N_8150,N_8392);
nand U8878 (N_8878,N_8434,N_8354);
and U8879 (N_8879,N_8346,N_8223);
nor U8880 (N_8880,N_8005,N_8271);
xor U8881 (N_8881,N_8023,N_8180);
or U8882 (N_8882,N_8425,N_8422);
nor U8883 (N_8883,N_8109,N_8301);
nor U8884 (N_8884,N_8238,N_8317);
nor U8885 (N_8885,N_8432,N_8266);
and U8886 (N_8886,N_8424,N_8348);
and U8887 (N_8887,N_8492,N_8357);
nand U8888 (N_8888,N_8321,N_8152);
or U8889 (N_8889,N_8096,N_8380);
and U8890 (N_8890,N_8483,N_8175);
and U8891 (N_8891,N_8087,N_8260);
nor U8892 (N_8892,N_8246,N_8255);
xor U8893 (N_8893,N_8266,N_8418);
nor U8894 (N_8894,N_8315,N_8019);
or U8895 (N_8895,N_8411,N_8402);
and U8896 (N_8896,N_8213,N_8255);
nor U8897 (N_8897,N_8408,N_8233);
nand U8898 (N_8898,N_8273,N_8155);
xor U8899 (N_8899,N_8046,N_8114);
nand U8900 (N_8900,N_8481,N_8358);
nand U8901 (N_8901,N_8247,N_8404);
or U8902 (N_8902,N_8180,N_8064);
and U8903 (N_8903,N_8032,N_8134);
nand U8904 (N_8904,N_8140,N_8187);
and U8905 (N_8905,N_8278,N_8483);
and U8906 (N_8906,N_8019,N_8323);
xor U8907 (N_8907,N_8445,N_8307);
nand U8908 (N_8908,N_8004,N_8219);
and U8909 (N_8909,N_8286,N_8360);
xor U8910 (N_8910,N_8045,N_8031);
nor U8911 (N_8911,N_8468,N_8292);
or U8912 (N_8912,N_8219,N_8484);
nand U8913 (N_8913,N_8356,N_8472);
xnor U8914 (N_8914,N_8015,N_8381);
and U8915 (N_8915,N_8114,N_8258);
or U8916 (N_8916,N_8429,N_8354);
nor U8917 (N_8917,N_8079,N_8269);
nand U8918 (N_8918,N_8059,N_8015);
xor U8919 (N_8919,N_8495,N_8202);
xnor U8920 (N_8920,N_8032,N_8021);
nand U8921 (N_8921,N_8293,N_8461);
nand U8922 (N_8922,N_8278,N_8181);
nand U8923 (N_8923,N_8382,N_8021);
and U8924 (N_8924,N_8277,N_8303);
and U8925 (N_8925,N_8102,N_8291);
xor U8926 (N_8926,N_8071,N_8338);
nand U8927 (N_8927,N_8315,N_8304);
and U8928 (N_8928,N_8046,N_8431);
and U8929 (N_8929,N_8240,N_8192);
nand U8930 (N_8930,N_8232,N_8472);
or U8931 (N_8931,N_8355,N_8455);
xor U8932 (N_8932,N_8049,N_8221);
xnor U8933 (N_8933,N_8203,N_8465);
xnor U8934 (N_8934,N_8112,N_8036);
or U8935 (N_8935,N_8394,N_8483);
xor U8936 (N_8936,N_8338,N_8186);
nand U8937 (N_8937,N_8062,N_8063);
and U8938 (N_8938,N_8268,N_8372);
and U8939 (N_8939,N_8311,N_8478);
nor U8940 (N_8940,N_8467,N_8244);
or U8941 (N_8941,N_8269,N_8419);
and U8942 (N_8942,N_8221,N_8215);
and U8943 (N_8943,N_8263,N_8446);
nand U8944 (N_8944,N_8195,N_8410);
and U8945 (N_8945,N_8260,N_8309);
xor U8946 (N_8946,N_8314,N_8222);
xor U8947 (N_8947,N_8070,N_8074);
or U8948 (N_8948,N_8486,N_8045);
xnor U8949 (N_8949,N_8380,N_8408);
and U8950 (N_8950,N_8458,N_8042);
nor U8951 (N_8951,N_8376,N_8481);
nor U8952 (N_8952,N_8498,N_8331);
nand U8953 (N_8953,N_8414,N_8249);
and U8954 (N_8954,N_8439,N_8494);
nand U8955 (N_8955,N_8274,N_8209);
xor U8956 (N_8956,N_8443,N_8125);
xnor U8957 (N_8957,N_8046,N_8272);
or U8958 (N_8958,N_8174,N_8251);
xnor U8959 (N_8959,N_8497,N_8476);
xor U8960 (N_8960,N_8185,N_8252);
and U8961 (N_8961,N_8001,N_8030);
and U8962 (N_8962,N_8487,N_8190);
xnor U8963 (N_8963,N_8049,N_8092);
nor U8964 (N_8964,N_8078,N_8202);
and U8965 (N_8965,N_8320,N_8016);
nand U8966 (N_8966,N_8310,N_8092);
or U8967 (N_8967,N_8079,N_8300);
nor U8968 (N_8968,N_8145,N_8355);
or U8969 (N_8969,N_8409,N_8309);
nand U8970 (N_8970,N_8415,N_8234);
and U8971 (N_8971,N_8330,N_8442);
nor U8972 (N_8972,N_8074,N_8210);
and U8973 (N_8973,N_8026,N_8137);
nor U8974 (N_8974,N_8249,N_8165);
and U8975 (N_8975,N_8127,N_8296);
nor U8976 (N_8976,N_8368,N_8484);
and U8977 (N_8977,N_8228,N_8273);
nor U8978 (N_8978,N_8025,N_8134);
nor U8979 (N_8979,N_8261,N_8058);
and U8980 (N_8980,N_8479,N_8333);
and U8981 (N_8981,N_8060,N_8288);
nand U8982 (N_8982,N_8013,N_8091);
nand U8983 (N_8983,N_8135,N_8379);
nor U8984 (N_8984,N_8217,N_8415);
and U8985 (N_8985,N_8231,N_8219);
nor U8986 (N_8986,N_8433,N_8067);
or U8987 (N_8987,N_8214,N_8422);
nor U8988 (N_8988,N_8086,N_8071);
nor U8989 (N_8989,N_8394,N_8254);
xnor U8990 (N_8990,N_8481,N_8434);
and U8991 (N_8991,N_8036,N_8497);
or U8992 (N_8992,N_8121,N_8363);
and U8993 (N_8993,N_8474,N_8186);
xnor U8994 (N_8994,N_8231,N_8002);
nand U8995 (N_8995,N_8094,N_8073);
nand U8996 (N_8996,N_8355,N_8001);
and U8997 (N_8997,N_8245,N_8131);
and U8998 (N_8998,N_8081,N_8213);
or U8999 (N_8999,N_8005,N_8198);
xnor U9000 (N_9000,N_8760,N_8829);
and U9001 (N_9001,N_8837,N_8508);
nor U9002 (N_9002,N_8613,N_8570);
and U9003 (N_9003,N_8581,N_8878);
xor U9004 (N_9004,N_8935,N_8907);
nor U9005 (N_9005,N_8506,N_8709);
xor U9006 (N_9006,N_8763,N_8729);
and U9007 (N_9007,N_8942,N_8710);
nand U9008 (N_9008,N_8993,N_8732);
and U9009 (N_9009,N_8784,N_8800);
or U9010 (N_9010,N_8597,N_8568);
nand U9011 (N_9011,N_8847,N_8670);
nor U9012 (N_9012,N_8913,N_8814);
xnor U9013 (N_9013,N_8534,N_8662);
and U9014 (N_9014,N_8676,N_8767);
or U9015 (N_9015,N_8781,N_8545);
and U9016 (N_9016,N_8538,N_8957);
nand U9017 (N_9017,N_8695,N_8787);
or U9018 (N_9018,N_8778,N_8811);
and U9019 (N_9019,N_8572,N_8702);
and U9020 (N_9020,N_8832,N_8815);
and U9021 (N_9021,N_8647,N_8902);
or U9022 (N_9022,N_8697,N_8773);
xnor U9023 (N_9023,N_8877,N_8794);
nand U9024 (N_9024,N_8565,N_8549);
or U9025 (N_9025,N_8827,N_8685);
xor U9026 (N_9026,N_8922,N_8866);
or U9027 (N_9027,N_8514,N_8511);
nand U9028 (N_9028,N_8901,N_8680);
nand U9029 (N_9029,N_8688,N_8980);
or U9030 (N_9030,N_8985,N_8655);
and U9031 (N_9031,N_8937,N_8677);
nand U9032 (N_9032,N_8616,N_8965);
xnor U9033 (N_9033,N_8700,N_8660);
nor U9034 (N_9034,N_8588,N_8560);
nand U9035 (N_9035,N_8524,N_8654);
and U9036 (N_9036,N_8924,N_8584);
nor U9037 (N_9037,N_8961,N_8605);
and U9038 (N_9038,N_8822,N_8667);
and U9039 (N_9039,N_8651,N_8635);
or U9040 (N_9040,N_8772,N_8983);
or U9041 (N_9041,N_8683,N_8792);
or U9042 (N_9042,N_8589,N_8898);
and U9043 (N_9043,N_8868,N_8759);
or U9044 (N_9044,N_8958,N_8741);
nor U9045 (N_9045,N_8909,N_8520);
xor U9046 (N_9046,N_8779,N_8641);
nor U9047 (N_9047,N_8795,N_8876);
nor U9048 (N_9048,N_8887,N_8665);
and U9049 (N_9049,N_8675,N_8559);
or U9050 (N_9050,N_8531,N_8970);
or U9051 (N_9051,N_8879,N_8602);
nand U9052 (N_9052,N_8528,N_8736);
nand U9053 (N_9053,N_8894,N_8558);
nand U9054 (N_9054,N_8798,N_8543);
and U9055 (N_9055,N_8755,N_8610);
or U9056 (N_9056,N_8889,N_8706);
and U9057 (N_9057,N_8502,N_8599);
and U9058 (N_9058,N_8673,N_8933);
and U9059 (N_9059,N_8649,N_8843);
and U9060 (N_9060,N_8928,N_8750);
nor U9061 (N_9061,N_8940,N_8854);
and U9062 (N_9062,N_8834,N_8758);
or U9063 (N_9063,N_8927,N_8842);
xor U9064 (N_9064,N_8845,N_8972);
nand U9065 (N_9065,N_8557,N_8517);
nor U9066 (N_9066,N_8780,N_8804);
and U9067 (N_9067,N_8672,N_8592);
nor U9068 (N_9068,N_8640,N_8810);
xor U9069 (N_9069,N_8960,N_8872);
or U9070 (N_9070,N_8747,N_8663);
nand U9071 (N_9071,N_8619,N_8802);
or U9072 (N_9072,N_8918,N_8659);
or U9073 (N_9073,N_8608,N_8949);
or U9074 (N_9074,N_8809,N_8537);
xnor U9075 (N_9075,N_8578,N_8875);
xnor U9076 (N_9076,N_8874,N_8626);
xor U9077 (N_9077,N_8733,N_8699);
or U9078 (N_9078,N_8527,N_8686);
or U9079 (N_9079,N_8938,N_8586);
nand U9080 (N_9080,N_8519,N_8783);
nor U9081 (N_9081,N_8751,N_8745);
nand U9082 (N_9082,N_8535,N_8712);
nor U9083 (N_9083,N_8791,N_8807);
and U9084 (N_9084,N_8547,N_8861);
nor U9085 (N_9085,N_8645,N_8738);
xnor U9086 (N_9086,N_8777,N_8835);
xnor U9087 (N_9087,N_8906,N_8696);
and U9088 (N_9088,N_8513,N_8575);
xnor U9089 (N_9089,N_8959,N_8540);
or U9090 (N_9090,N_8943,N_8657);
xor U9091 (N_9091,N_8652,N_8982);
nor U9092 (N_9092,N_8515,N_8737);
nand U9093 (N_9093,N_8512,N_8704);
or U9094 (N_9094,N_8687,N_8742);
and U9095 (N_9095,N_8743,N_8618);
or U9096 (N_9096,N_8669,N_8542);
xnor U9097 (N_9097,N_8816,N_8674);
and U9098 (N_9098,N_8689,N_8721);
and U9099 (N_9099,N_8853,N_8881);
and U9100 (N_9100,N_8808,N_8871);
xnor U9101 (N_9101,N_8668,N_8595);
or U9102 (N_9102,N_8653,N_8757);
nand U9103 (N_9103,N_8701,N_8756);
nor U9104 (N_9104,N_8503,N_8555);
and U9105 (N_9105,N_8833,N_8846);
nand U9106 (N_9106,N_8782,N_8786);
and U9107 (N_9107,N_8978,N_8968);
and U9108 (N_9108,N_8698,N_8614);
and U9109 (N_9109,N_8691,N_8604);
nand U9110 (N_9110,N_8880,N_8591);
nand U9111 (N_9111,N_8716,N_8646);
nor U9112 (N_9112,N_8761,N_8830);
nor U9113 (N_9113,N_8857,N_8639);
nor U9114 (N_9114,N_8941,N_8799);
nand U9115 (N_9115,N_8931,N_8921);
xor U9116 (N_9116,N_8582,N_8577);
xor U9117 (N_9117,N_8867,N_8529);
nand U9118 (N_9118,N_8951,N_8740);
xor U9119 (N_9119,N_8671,N_8911);
or U9120 (N_9120,N_8892,N_8950);
xnor U9121 (N_9121,N_8554,N_8914);
and U9122 (N_9122,N_8539,N_8828);
xor U9123 (N_9123,N_8936,N_8724);
nor U9124 (N_9124,N_8826,N_8932);
nand U9125 (N_9125,N_8548,N_8988);
or U9126 (N_9126,N_8583,N_8630);
xor U9127 (N_9127,N_8963,N_8908);
nand U9128 (N_9128,N_8730,N_8703);
nand U9129 (N_9129,N_8728,N_8637);
nand U9130 (N_9130,N_8998,N_8770);
or U9131 (N_9131,N_8598,N_8899);
and U9132 (N_9132,N_8530,N_8930);
and U9133 (N_9133,N_8812,N_8771);
nor U9134 (N_9134,N_8962,N_8522);
nor U9135 (N_9135,N_8536,N_8650);
or U9136 (N_9136,N_8720,N_8805);
nor U9137 (N_9137,N_8882,N_8885);
nor U9138 (N_9138,N_8790,N_8574);
and U9139 (N_9139,N_8974,N_8831);
nand U9140 (N_9140,N_8863,N_8523);
nand U9141 (N_9141,N_8516,N_8994);
xnor U9142 (N_9142,N_8768,N_8748);
and U9143 (N_9143,N_8955,N_8886);
and U9144 (N_9144,N_8573,N_8693);
and U9145 (N_9145,N_8579,N_8617);
nand U9146 (N_9146,N_8855,N_8681);
nor U9147 (N_9147,N_8897,N_8825);
xor U9148 (N_9148,N_8905,N_8566);
nor U9149 (N_9149,N_8838,N_8569);
or U9150 (N_9150,N_8904,N_8788);
nor U9151 (N_9151,N_8563,N_8916);
nor U9152 (N_9152,N_8900,N_8851);
nor U9153 (N_9153,N_8501,N_8923);
or U9154 (N_9154,N_8509,N_8769);
nor U9155 (N_9155,N_8552,N_8731);
or U9156 (N_9156,N_8926,N_8708);
nand U9157 (N_9157,N_8919,N_8858);
nor U9158 (N_9158,N_8797,N_8521);
nor U9159 (N_9159,N_8801,N_8644);
nand U9160 (N_9160,N_8947,N_8884);
nor U9161 (N_9161,N_8550,N_8986);
xor U9162 (N_9162,N_8609,N_8992);
or U9163 (N_9163,N_8896,N_8623);
nor U9164 (N_9164,N_8722,N_8607);
xor U9165 (N_9165,N_8796,N_8526);
nand U9166 (N_9166,N_8723,N_8628);
nand U9167 (N_9167,N_8561,N_8991);
or U9168 (N_9168,N_8859,N_8713);
and U9169 (N_9169,N_8964,N_8603);
and U9170 (N_9170,N_8622,N_8803);
or U9171 (N_9171,N_8611,N_8925);
nand U9172 (N_9172,N_8594,N_8507);
xnor U9173 (N_9173,N_8564,N_8966);
nor U9174 (N_9174,N_8785,N_8819);
or U9175 (N_9175,N_8711,N_8870);
nand U9176 (N_9176,N_8590,N_8500);
nand U9177 (N_9177,N_8553,N_8956);
nand U9178 (N_9178,N_8969,N_8541);
or U9179 (N_9179,N_8839,N_8585);
or U9180 (N_9180,N_8580,N_8690);
and U9181 (N_9181,N_8775,N_8694);
and U9182 (N_9182,N_8726,N_8633);
nor U9183 (N_9183,N_8817,N_8656);
or U9184 (N_9184,N_8606,N_8944);
nor U9185 (N_9185,N_8890,N_8648);
nand U9186 (N_9186,N_8620,N_8824);
or U9187 (N_9187,N_8504,N_8789);
nand U9188 (N_9188,N_8975,N_8642);
nor U9189 (N_9189,N_8735,N_8596);
nor U9190 (N_9190,N_8734,N_8762);
nor U9191 (N_9191,N_8952,N_8634);
nor U9192 (N_9192,N_8510,N_8915);
nand U9193 (N_9193,N_8849,N_8954);
or U9194 (N_9194,N_8967,N_8840);
nor U9195 (N_9195,N_8891,N_8869);
and U9196 (N_9196,N_8749,N_8636);
nand U9197 (N_9197,N_8912,N_8627);
or U9198 (N_9198,N_8895,N_8518);
nand U9199 (N_9199,N_8679,N_8571);
nor U9200 (N_9200,N_8984,N_8989);
nor U9201 (N_9201,N_8546,N_8638);
nor U9202 (N_9202,N_8692,N_8666);
or U9203 (N_9203,N_8764,N_8551);
xor U9204 (N_9204,N_8893,N_8727);
xor U9205 (N_9205,N_8836,N_8865);
nor U9206 (N_9206,N_8841,N_8682);
xnor U9207 (N_9207,N_8714,N_8664);
nand U9208 (N_9208,N_8766,N_8739);
xor U9209 (N_9209,N_8920,N_8615);
xor U9210 (N_9210,N_8621,N_8976);
nor U9211 (N_9211,N_8939,N_8883);
nand U9212 (N_9212,N_8848,N_8973);
or U9213 (N_9213,N_8562,N_8567);
xnor U9214 (N_9214,N_8860,N_8945);
or U9215 (N_9215,N_8888,N_8707);
xor U9216 (N_9216,N_8658,N_8776);
or U9217 (N_9217,N_8533,N_8844);
or U9218 (N_9218,N_8544,N_8820);
and U9219 (N_9219,N_8601,N_8505);
nor U9220 (N_9220,N_8532,N_8996);
xnor U9221 (N_9221,N_8981,N_8813);
xnor U9222 (N_9222,N_8873,N_8821);
and U9223 (N_9223,N_8823,N_8971);
xnor U9224 (N_9224,N_8725,N_8862);
and U9225 (N_9225,N_8903,N_8718);
xnor U9226 (N_9226,N_8910,N_8995);
xor U9227 (N_9227,N_8856,N_8864);
or U9228 (N_9228,N_8746,N_8754);
nor U9229 (N_9229,N_8997,N_8765);
nor U9230 (N_9230,N_8987,N_8631);
nor U9231 (N_9231,N_8600,N_8999);
or U9232 (N_9232,N_8525,N_8806);
and U9233 (N_9233,N_8684,N_8705);
and U9234 (N_9234,N_8953,N_8715);
xor U9235 (N_9235,N_8990,N_8752);
nand U9236 (N_9236,N_8629,N_8587);
nand U9237 (N_9237,N_8576,N_8946);
nand U9238 (N_9238,N_8593,N_8948);
xor U9239 (N_9239,N_8850,N_8929);
nor U9240 (N_9240,N_8719,N_8852);
nor U9241 (N_9241,N_8744,N_8917);
or U9242 (N_9242,N_8556,N_8624);
xor U9243 (N_9243,N_8612,N_8678);
and U9244 (N_9244,N_8934,N_8643);
nand U9245 (N_9245,N_8753,N_8774);
xnor U9246 (N_9246,N_8977,N_8793);
nand U9247 (N_9247,N_8717,N_8625);
xor U9248 (N_9248,N_8979,N_8661);
nand U9249 (N_9249,N_8632,N_8818);
nand U9250 (N_9250,N_8763,N_8567);
nand U9251 (N_9251,N_8748,N_8505);
xnor U9252 (N_9252,N_8825,N_8777);
and U9253 (N_9253,N_8702,N_8794);
xnor U9254 (N_9254,N_8688,N_8665);
nand U9255 (N_9255,N_8582,N_8876);
nand U9256 (N_9256,N_8533,N_8720);
and U9257 (N_9257,N_8678,N_8722);
nor U9258 (N_9258,N_8960,N_8888);
and U9259 (N_9259,N_8853,N_8730);
or U9260 (N_9260,N_8991,N_8583);
nor U9261 (N_9261,N_8730,N_8908);
and U9262 (N_9262,N_8780,N_8741);
or U9263 (N_9263,N_8817,N_8583);
or U9264 (N_9264,N_8939,N_8850);
nand U9265 (N_9265,N_8541,N_8651);
and U9266 (N_9266,N_8512,N_8964);
xnor U9267 (N_9267,N_8590,N_8899);
nor U9268 (N_9268,N_8822,N_8929);
nor U9269 (N_9269,N_8771,N_8784);
or U9270 (N_9270,N_8554,N_8829);
xor U9271 (N_9271,N_8873,N_8624);
or U9272 (N_9272,N_8567,N_8849);
nor U9273 (N_9273,N_8510,N_8818);
or U9274 (N_9274,N_8759,N_8615);
xor U9275 (N_9275,N_8536,N_8586);
nor U9276 (N_9276,N_8545,N_8927);
nor U9277 (N_9277,N_8874,N_8943);
xnor U9278 (N_9278,N_8658,N_8859);
xnor U9279 (N_9279,N_8827,N_8757);
nand U9280 (N_9280,N_8987,N_8709);
and U9281 (N_9281,N_8630,N_8950);
nor U9282 (N_9282,N_8830,N_8717);
xor U9283 (N_9283,N_8646,N_8814);
or U9284 (N_9284,N_8731,N_8967);
and U9285 (N_9285,N_8751,N_8656);
and U9286 (N_9286,N_8658,N_8796);
or U9287 (N_9287,N_8877,N_8590);
nand U9288 (N_9288,N_8895,N_8528);
and U9289 (N_9289,N_8765,N_8936);
and U9290 (N_9290,N_8535,N_8549);
or U9291 (N_9291,N_8592,N_8600);
and U9292 (N_9292,N_8834,N_8968);
xor U9293 (N_9293,N_8731,N_8634);
nand U9294 (N_9294,N_8717,N_8794);
nor U9295 (N_9295,N_8764,N_8654);
nand U9296 (N_9296,N_8840,N_8806);
and U9297 (N_9297,N_8628,N_8539);
and U9298 (N_9298,N_8655,N_8553);
and U9299 (N_9299,N_8608,N_8944);
nor U9300 (N_9300,N_8853,N_8743);
and U9301 (N_9301,N_8941,N_8637);
nor U9302 (N_9302,N_8937,N_8830);
nand U9303 (N_9303,N_8736,N_8571);
nand U9304 (N_9304,N_8511,N_8776);
xor U9305 (N_9305,N_8855,N_8972);
and U9306 (N_9306,N_8747,N_8706);
xor U9307 (N_9307,N_8790,N_8632);
xor U9308 (N_9308,N_8891,N_8647);
nor U9309 (N_9309,N_8999,N_8949);
and U9310 (N_9310,N_8531,N_8620);
or U9311 (N_9311,N_8575,N_8982);
nor U9312 (N_9312,N_8779,N_8678);
xnor U9313 (N_9313,N_8995,N_8894);
or U9314 (N_9314,N_8954,N_8761);
xnor U9315 (N_9315,N_8900,N_8608);
nor U9316 (N_9316,N_8699,N_8640);
or U9317 (N_9317,N_8813,N_8965);
nor U9318 (N_9318,N_8850,N_8798);
and U9319 (N_9319,N_8694,N_8684);
or U9320 (N_9320,N_8714,N_8519);
xor U9321 (N_9321,N_8870,N_8702);
nand U9322 (N_9322,N_8533,N_8889);
xor U9323 (N_9323,N_8746,N_8593);
or U9324 (N_9324,N_8527,N_8979);
and U9325 (N_9325,N_8683,N_8760);
nor U9326 (N_9326,N_8758,N_8541);
nor U9327 (N_9327,N_8861,N_8634);
or U9328 (N_9328,N_8683,N_8904);
nor U9329 (N_9329,N_8678,N_8693);
xor U9330 (N_9330,N_8624,N_8535);
nand U9331 (N_9331,N_8636,N_8560);
nand U9332 (N_9332,N_8905,N_8707);
xor U9333 (N_9333,N_8991,N_8994);
and U9334 (N_9334,N_8942,N_8886);
nand U9335 (N_9335,N_8655,N_8545);
or U9336 (N_9336,N_8734,N_8531);
or U9337 (N_9337,N_8588,N_8774);
nand U9338 (N_9338,N_8898,N_8811);
or U9339 (N_9339,N_8869,N_8707);
and U9340 (N_9340,N_8607,N_8709);
nor U9341 (N_9341,N_8992,N_8569);
nand U9342 (N_9342,N_8726,N_8508);
nor U9343 (N_9343,N_8940,N_8826);
or U9344 (N_9344,N_8999,N_8920);
or U9345 (N_9345,N_8513,N_8673);
and U9346 (N_9346,N_8840,N_8821);
and U9347 (N_9347,N_8800,N_8535);
or U9348 (N_9348,N_8605,N_8629);
xnor U9349 (N_9349,N_8775,N_8656);
or U9350 (N_9350,N_8762,N_8774);
xor U9351 (N_9351,N_8859,N_8847);
xnor U9352 (N_9352,N_8911,N_8750);
nor U9353 (N_9353,N_8977,N_8934);
nor U9354 (N_9354,N_8739,N_8635);
or U9355 (N_9355,N_8705,N_8501);
or U9356 (N_9356,N_8852,N_8877);
or U9357 (N_9357,N_8517,N_8877);
nand U9358 (N_9358,N_8801,N_8967);
xnor U9359 (N_9359,N_8643,N_8945);
or U9360 (N_9360,N_8748,N_8855);
or U9361 (N_9361,N_8748,N_8648);
and U9362 (N_9362,N_8590,N_8570);
xnor U9363 (N_9363,N_8881,N_8731);
xor U9364 (N_9364,N_8997,N_8510);
nand U9365 (N_9365,N_8950,N_8710);
and U9366 (N_9366,N_8904,N_8937);
and U9367 (N_9367,N_8682,N_8891);
or U9368 (N_9368,N_8624,N_8635);
nor U9369 (N_9369,N_8630,N_8701);
or U9370 (N_9370,N_8546,N_8910);
xor U9371 (N_9371,N_8814,N_8984);
nor U9372 (N_9372,N_8677,N_8986);
or U9373 (N_9373,N_8669,N_8612);
nand U9374 (N_9374,N_8551,N_8532);
or U9375 (N_9375,N_8639,N_8602);
xnor U9376 (N_9376,N_8515,N_8649);
or U9377 (N_9377,N_8998,N_8672);
nand U9378 (N_9378,N_8786,N_8894);
xor U9379 (N_9379,N_8950,N_8577);
nand U9380 (N_9380,N_8699,N_8654);
nand U9381 (N_9381,N_8528,N_8844);
xor U9382 (N_9382,N_8661,N_8578);
or U9383 (N_9383,N_8565,N_8795);
nand U9384 (N_9384,N_8877,N_8614);
xnor U9385 (N_9385,N_8582,N_8619);
xnor U9386 (N_9386,N_8650,N_8826);
or U9387 (N_9387,N_8980,N_8568);
nand U9388 (N_9388,N_8814,N_8584);
and U9389 (N_9389,N_8576,N_8956);
and U9390 (N_9390,N_8991,N_8802);
and U9391 (N_9391,N_8908,N_8922);
or U9392 (N_9392,N_8722,N_8688);
and U9393 (N_9393,N_8909,N_8533);
or U9394 (N_9394,N_8656,N_8806);
xnor U9395 (N_9395,N_8972,N_8567);
nand U9396 (N_9396,N_8898,N_8750);
and U9397 (N_9397,N_8947,N_8609);
nor U9398 (N_9398,N_8561,N_8671);
and U9399 (N_9399,N_8971,N_8824);
nand U9400 (N_9400,N_8619,N_8907);
nor U9401 (N_9401,N_8911,N_8847);
or U9402 (N_9402,N_8852,N_8806);
and U9403 (N_9403,N_8873,N_8526);
xor U9404 (N_9404,N_8526,N_8584);
nor U9405 (N_9405,N_8960,N_8946);
xor U9406 (N_9406,N_8864,N_8817);
xor U9407 (N_9407,N_8780,N_8976);
nor U9408 (N_9408,N_8577,N_8652);
xor U9409 (N_9409,N_8997,N_8976);
nand U9410 (N_9410,N_8696,N_8630);
and U9411 (N_9411,N_8970,N_8727);
nand U9412 (N_9412,N_8854,N_8745);
xnor U9413 (N_9413,N_8989,N_8958);
xnor U9414 (N_9414,N_8504,N_8844);
and U9415 (N_9415,N_8551,N_8708);
nand U9416 (N_9416,N_8617,N_8541);
nand U9417 (N_9417,N_8685,N_8922);
and U9418 (N_9418,N_8911,N_8913);
and U9419 (N_9419,N_8714,N_8652);
nand U9420 (N_9420,N_8570,N_8855);
nand U9421 (N_9421,N_8961,N_8626);
nand U9422 (N_9422,N_8631,N_8580);
or U9423 (N_9423,N_8926,N_8510);
nor U9424 (N_9424,N_8597,N_8594);
nor U9425 (N_9425,N_8792,N_8610);
nand U9426 (N_9426,N_8938,N_8706);
or U9427 (N_9427,N_8952,N_8589);
and U9428 (N_9428,N_8658,N_8890);
or U9429 (N_9429,N_8868,N_8708);
nor U9430 (N_9430,N_8882,N_8714);
nor U9431 (N_9431,N_8654,N_8523);
xnor U9432 (N_9432,N_8651,N_8747);
xnor U9433 (N_9433,N_8645,N_8603);
nand U9434 (N_9434,N_8881,N_8545);
xor U9435 (N_9435,N_8550,N_8534);
xor U9436 (N_9436,N_8743,N_8975);
nor U9437 (N_9437,N_8538,N_8859);
or U9438 (N_9438,N_8895,N_8894);
nor U9439 (N_9439,N_8550,N_8958);
xnor U9440 (N_9440,N_8669,N_8665);
or U9441 (N_9441,N_8817,N_8814);
nand U9442 (N_9442,N_8656,N_8528);
nor U9443 (N_9443,N_8983,N_8746);
xnor U9444 (N_9444,N_8940,N_8735);
nand U9445 (N_9445,N_8906,N_8550);
nand U9446 (N_9446,N_8628,N_8715);
nor U9447 (N_9447,N_8628,N_8765);
nand U9448 (N_9448,N_8969,N_8670);
nand U9449 (N_9449,N_8597,N_8914);
xor U9450 (N_9450,N_8596,N_8579);
and U9451 (N_9451,N_8925,N_8992);
xnor U9452 (N_9452,N_8594,N_8503);
or U9453 (N_9453,N_8683,N_8836);
nand U9454 (N_9454,N_8923,N_8833);
xnor U9455 (N_9455,N_8670,N_8895);
or U9456 (N_9456,N_8754,N_8837);
xor U9457 (N_9457,N_8921,N_8777);
or U9458 (N_9458,N_8813,N_8793);
nand U9459 (N_9459,N_8689,N_8606);
nand U9460 (N_9460,N_8934,N_8558);
xor U9461 (N_9461,N_8910,N_8641);
and U9462 (N_9462,N_8600,N_8912);
nor U9463 (N_9463,N_8756,N_8688);
nand U9464 (N_9464,N_8902,N_8788);
and U9465 (N_9465,N_8712,N_8636);
nand U9466 (N_9466,N_8920,N_8657);
nand U9467 (N_9467,N_8774,N_8840);
nor U9468 (N_9468,N_8556,N_8598);
or U9469 (N_9469,N_8910,N_8908);
or U9470 (N_9470,N_8665,N_8700);
and U9471 (N_9471,N_8844,N_8675);
nor U9472 (N_9472,N_8603,N_8817);
and U9473 (N_9473,N_8625,N_8849);
xor U9474 (N_9474,N_8607,N_8984);
xor U9475 (N_9475,N_8926,N_8537);
xor U9476 (N_9476,N_8583,N_8834);
and U9477 (N_9477,N_8735,N_8937);
xnor U9478 (N_9478,N_8594,N_8936);
or U9479 (N_9479,N_8544,N_8931);
or U9480 (N_9480,N_8959,N_8565);
or U9481 (N_9481,N_8636,N_8902);
nor U9482 (N_9482,N_8731,N_8812);
nor U9483 (N_9483,N_8739,N_8979);
and U9484 (N_9484,N_8504,N_8529);
nand U9485 (N_9485,N_8981,N_8736);
nor U9486 (N_9486,N_8945,N_8603);
or U9487 (N_9487,N_8570,N_8544);
and U9488 (N_9488,N_8991,N_8591);
or U9489 (N_9489,N_8846,N_8546);
xnor U9490 (N_9490,N_8898,N_8565);
or U9491 (N_9491,N_8519,N_8527);
nand U9492 (N_9492,N_8596,N_8973);
nand U9493 (N_9493,N_8963,N_8671);
nor U9494 (N_9494,N_8969,N_8907);
xor U9495 (N_9495,N_8885,N_8675);
nand U9496 (N_9496,N_8580,N_8892);
nand U9497 (N_9497,N_8502,N_8762);
xor U9498 (N_9498,N_8571,N_8530);
nand U9499 (N_9499,N_8807,N_8532);
and U9500 (N_9500,N_9157,N_9049);
or U9501 (N_9501,N_9364,N_9032);
or U9502 (N_9502,N_9040,N_9428);
and U9503 (N_9503,N_9248,N_9077);
xnor U9504 (N_9504,N_9115,N_9084);
and U9505 (N_9505,N_9346,N_9222);
nor U9506 (N_9506,N_9477,N_9490);
xor U9507 (N_9507,N_9168,N_9373);
xor U9508 (N_9508,N_9113,N_9182);
nor U9509 (N_9509,N_9270,N_9274);
nor U9510 (N_9510,N_9436,N_9127);
or U9511 (N_9511,N_9010,N_9489);
or U9512 (N_9512,N_9067,N_9474);
xnor U9513 (N_9513,N_9357,N_9259);
and U9514 (N_9514,N_9305,N_9273);
xnor U9515 (N_9515,N_9348,N_9355);
xnor U9516 (N_9516,N_9386,N_9241);
and U9517 (N_9517,N_9136,N_9382);
nand U9518 (N_9518,N_9470,N_9186);
xor U9519 (N_9519,N_9197,N_9023);
xnor U9520 (N_9520,N_9288,N_9371);
nand U9521 (N_9521,N_9362,N_9233);
and U9522 (N_9522,N_9140,N_9108);
or U9523 (N_9523,N_9327,N_9178);
nand U9524 (N_9524,N_9253,N_9063);
xor U9525 (N_9525,N_9004,N_9167);
or U9526 (N_9526,N_9413,N_9225);
nand U9527 (N_9527,N_9478,N_9419);
nand U9528 (N_9528,N_9358,N_9158);
xnor U9529 (N_9529,N_9333,N_9393);
and U9530 (N_9530,N_9202,N_9149);
or U9531 (N_9531,N_9070,N_9237);
and U9532 (N_9532,N_9006,N_9073);
nor U9533 (N_9533,N_9204,N_9352);
nor U9534 (N_9534,N_9121,N_9163);
xor U9535 (N_9535,N_9142,N_9174);
xnor U9536 (N_9536,N_9418,N_9492);
and U9537 (N_9537,N_9071,N_9043);
nor U9538 (N_9538,N_9155,N_9164);
xnor U9539 (N_9539,N_9190,N_9018);
or U9540 (N_9540,N_9302,N_9338);
nor U9541 (N_9541,N_9435,N_9031);
and U9542 (N_9542,N_9440,N_9332);
and U9543 (N_9543,N_9195,N_9154);
xor U9544 (N_9544,N_9465,N_9090);
or U9545 (N_9545,N_9014,N_9452);
or U9546 (N_9546,N_9317,N_9320);
and U9547 (N_9547,N_9254,N_9251);
and U9548 (N_9548,N_9238,N_9231);
nor U9549 (N_9549,N_9279,N_9214);
or U9550 (N_9550,N_9122,N_9161);
nand U9551 (N_9551,N_9235,N_9125);
nand U9552 (N_9552,N_9187,N_9116);
nor U9553 (N_9553,N_9030,N_9118);
nor U9554 (N_9554,N_9480,N_9497);
nor U9555 (N_9555,N_9488,N_9379);
nor U9556 (N_9556,N_9001,N_9138);
xor U9557 (N_9557,N_9337,N_9455);
or U9558 (N_9558,N_9261,N_9111);
or U9559 (N_9559,N_9196,N_9258);
or U9560 (N_9560,N_9313,N_9271);
nor U9561 (N_9561,N_9209,N_9124);
xnor U9562 (N_9562,N_9325,N_9473);
nand U9563 (N_9563,N_9495,N_9385);
or U9564 (N_9564,N_9434,N_9091);
xnor U9565 (N_9565,N_9285,N_9165);
and U9566 (N_9566,N_9276,N_9297);
or U9567 (N_9567,N_9060,N_9398);
and U9568 (N_9568,N_9079,N_9089);
nand U9569 (N_9569,N_9130,N_9395);
nor U9570 (N_9570,N_9099,N_9104);
xnor U9571 (N_9571,N_9052,N_9016);
or U9572 (N_9572,N_9374,N_9074);
nand U9573 (N_9573,N_9055,N_9384);
or U9574 (N_9574,N_9042,N_9180);
or U9575 (N_9575,N_9494,N_9101);
or U9576 (N_9576,N_9432,N_9107);
nand U9577 (N_9577,N_9098,N_9039);
and U9578 (N_9578,N_9024,N_9240);
nand U9579 (N_9579,N_9345,N_9114);
or U9580 (N_9580,N_9021,N_9422);
or U9581 (N_9581,N_9137,N_9106);
or U9582 (N_9582,N_9017,N_9466);
nand U9583 (N_9583,N_9076,N_9402);
and U9584 (N_9584,N_9380,N_9416);
and U9585 (N_9585,N_9227,N_9472);
or U9586 (N_9586,N_9173,N_9252);
nor U9587 (N_9587,N_9400,N_9341);
or U9588 (N_9588,N_9212,N_9189);
xnor U9589 (N_9589,N_9292,N_9405);
nand U9590 (N_9590,N_9131,N_9047);
nand U9591 (N_9591,N_9429,N_9095);
or U9592 (N_9592,N_9062,N_9061);
xor U9593 (N_9593,N_9399,N_9449);
and U9594 (N_9594,N_9065,N_9007);
xor U9595 (N_9595,N_9299,N_9456);
xnor U9596 (N_9596,N_9105,N_9457);
or U9597 (N_9597,N_9414,N_9217);
nor U9598 (N_9598,N_9289,N_9126);
nand U9599 (N_9599,N_9284,N_9257);
nand U9600 (N_9600,N_9044,N_9179);
nor U9601 (N_9601,N_9499,N_9396);
and U9602 (N_9602,N_9476,N_9319);
or U9603 (N_9603,N_9236,N_9367);
nor U9604 (N_9604,N_9128,N_9051);
and U9605 (N_9605,N_9314,N_9239);
nand U9606 (N_9606,N_9461,N_9135);
nand U9607 (N_9607,N_9378,N_9147);
xnor U9608 (N_9608,N_9117,N_9308);
xor U9609 (N_9609,N_9339,N_9304);
xnor U9610 (N_9610,N_9109,N_9340);
or U9611 (N_9611,N_9467,N_9205);
nand U9612 (N_9612,N_9309,N_9048);
nand U9613 (N_9613,N_9272,N_9224);
xor U9614 (N_9614,N_9387,N_9265);
and U9615 (N_9615,N_9143,N_9451);
and U9616 (N_9616,N_9268,N_9218);
and U9617 (N_9617,N_9496,N_9059);
and U9618 (N_9618,N_9471,N_9420);
or U9619 (N_9619,N_9283,N_9331);
xnor U9620 (N_9620,N_9294,N_9360);
and U9621 (N_9621,N_9232,N_9376);
nor U9622 (N_9622,N_9356,N_9056);
nand U9623 (N_9623,N_9086,N_9183);
xor U9624 (N_9624,N_9094,N_9354);
nor U9625 (N_9625,N_9353,N_9406);
or U9626 (N_9626,N_9003,N_9483);
and U9627 (N_9627,N_9038,N_9119);
or U9628 (N_9628,N_9170,N_9306);
nand U9629 (N_9629,N_9026,N_9041);
nand U9630 (N_9630,N_9475,N_9366);
or U9631 (N_9631,N_9200,N_9193);
nand U9632 (N_9632,N_9000,N_9390);
nor U9633 (N_9633,N_9444,N_9343);
xor U9634 (N_9634,N_9072,N_9141);
xnor U9635 (N_9635,N_9370,N_9267);
and U9636 (N_9636,N_9249,N_9152);
nand U9637 (N_9637,N_9321,N_9287);
or U9638 (N_9638,N_9050,N_9391);
nor U9639 (N_9639,N_9162,N_9151);
nor U9640 (N_9640,N_9087,N_9329);
xnor U9641 (N_9641,N_9171,N_9498);
or U9642 (N_9642,N_9198,N_9463);
or U9643 (N_9643,N_9092,N_9447);
xnor U9644 (N_9644,N_9129,N_9081);
and U9645 (N_9645,N_9250,N_9361);
or U9646 (N_9646,N_9057,N_9377);
and U9647 (N_9647,N_9369,N_9372);
and U9648 (N_9648,N_9433,N_9424);
nand U9649 (N_9649,N_9002,N_9011);
or U9650 (N_9650,N_9278,N_9083);
xnor U9651 (N_9651,N_9491,N_9303);
xor U9652 (N_9652,N_9192,N_9020);
nand U9653 (N_9653,N_9409,N_9365);
nand U9654 (N_9654,N_9479,N_9394);
or U9655 (N_9655,N_9295,N_9410);
nand U9656 (N_9656,N_9028,N_9110);
or U9657 (N_9657,N_9335,N_9166);
nor U9658 (N_9658,N_9013,N_9347);
xor U9659 (N_9659,N_9426,N_9260);
and U9660 (N_9660,N_9228,N_9234);
nand U9661 (N_9661,N_9160,N_9493);
nand U9662 (N_9662,N_9363,N_9342);
xor U9663 (N_9663,N_9069,N_9458);
nor U9664 (N_9664,N_9008,N_9188);
xor U9665 (N_9665,N_9243,N_9185);
xor U9666 (N_9666,N_9009,N_9134);
nand U9667 (N_9667,N_9423,N_9263);
nor U9668 (N_9668,N_9034,N_9427);
nand U9669 (N_9669,N_9176,N_9025);
xnor U9670 (N_9670,N_9407,N_9159);
xnor U9671 (N_9671,N_9229,N_9266);
xor U9672 (N_9672,N_9037,N_9033);
or U9673 (N_9673,N_9112,N_9281);
nand U9674 (N_9674,N_9027,N_9213);
nand U9675 (N_9675,N_9169,N_9242);
and U9676 (N_9676,N_9156,N_9307);
nand U9677 (N_9677,N_9397,N_9103);
and U9678 (N_9678,N_9264,N_9350);
nand U9679 (N_9679,N_9298,N_9330);
or U9680 (N_9680,N_9191,N_9445);
or U9681 (N_9681,N_9417,N_9153);
and U9682 (N_9682,N_9256,N_9215);
nand U9683 (N_9683,N_9146,N_9058);
and U9684 (N_9684,N_9068,N_9208);
nor U9685 (N_9685,N_9139,N_9301);
and U9686 (N_9686,N_9085,N_9311);
xor U9687 (N_9687,N_9053,N_9066);
nand U9688 (N_9688,N_9184,N_9255);
or U9689 (N_9689,N_9210,N_9282);
and U9690 (N_9690,N_9132,N_9207);
nor U9691 (N_9691,N_9230,N_9097);
or U9692 (N_9692,N_9381,N_9262);
nor U9693 (N_9693,N_9296,N_9148);
nor U9694 (N_9694,N_9312,N_9269);
or U9695 (N_9695,N_9448,N_9482);
or U9696 (N_9696,N_9464,N_9012);
and U9697 (N_9697,N_9468,N_9383);
or U9698 (N_9698,N_9438,N_9421);
xor U9699 (N_9699,N_9247,N_9401);
and U9700 (N_9700,N_9453,N_9064);
or U9701 (N_9701,N_9203,N_9080);
or U9702 (N_9702,N_9144,N_9430);
nor U9703 (N_9703,N_9462,N_9145);
xor U9704 (N_9704,N_9469,N_9280);
xnor U9705 (N_9705,N_9323,N_9005);
xor U9706 (N_9706,N_9442,N_9439);
nand U9707 (N_9707,N_9315,N_9293);
xnor U9708 (N_9708,N_9310,N_9088);
or U9709 (N_9709,N_9133,N_9223);
xor U9710 (N_9710,N_9441,N_9316);
and U9711 (N_9711,N_9326,N_9368);
nor U9712 (N_9712,N_9450,N_9351);
and U9713 (N_9713,N_9318,N_9029);
nand U9714 (N_9714,N_9392,N_9035);
or U9715 (N_9715,N_9359,N_9246);
xnor U9716 (N_9716,N_9388,N_9460);
xor U9717 (N_9717,N_9054,N_9150);
or U9718 (N_9718,N_9181,N_9075);
xnor U9719 (N_9719,N_9201,N_9425);
nand U9720 (N_9720,N_9022,N_9291);
nor U9721 (N_9721,N_9199,N_9486);
or U9722 (N_9722,N_9172,N_9045);
xor U9723 (N_9723,N_9485,N_9211);
or U9724 (N_9724,N_9226,N_9437);
nand U9725 (N_9725,N_9120,N_9015);
nor U9726 (N_9726,N_9082,N_9322);
or U9727 (N_9727,N_9344,N_9349);
and U9728 (N_9728,N_9487,N_9046);
nor U9729 (N_9729,N_9336,N_9093);
nand U9730 (N_9730,N_9286,N_9328);
nor U9731 (N_9731,N_9411,N_9443);
xnor U9732 (N_9732,N_9375,N_9036);
xnor U9733 (N_9733,N_9408,N_9220);
xnor U9734 (N_9734,N_9177,N_9459);
nand U9735 (N_9735,N_9389,N_9403);
nor U9736 (N_9736,N_9123,N_9019);
and U9737 (N_9737,N_9481,N_9431);
nand U9738 (N_9738,N_9277,N_9404);
and U9739 (N_9739,N_9102,N_9415);
nand U9740 (N_9740,N_9412,N_9334);
and U9741 (N_9741,N_9245,N_9078);
xnor U9742 (N_9742,N_9221,N_9175);
or U9743 (N_9743,N_9216,N_9454);
and U9744 (N_9744,N_9206,N_9194);
and U9745 (N_9745,N_9100,N_9484);
xor U9746 (N_9746,N_9096,N_9300);
nand U9747 (N_9747,N_9446,N_9290);
xnor U9748 (N_9748,N_9275,N_9244);
nand U9749 (N_9749,N_9219,N_9324);
nand U9750 (N_9750,N_9032,N_9242);
nand U9751 (N_9751,N_9183,N_9013);
and U9752 (N_9752,N_9297,N_9178);
xor U9753 (N_9753,N_9007,N_9286);
and U9754 (N_9754,N_9498,N_9477);
nand U9755 (N_9755,N_9350,N_9149);
or U9756 (N_9756,N_9452,N_9488);
and U9757 (N_9757,N_9449,N_9334);
nand U9758 (N_9758,N_9158,N_9040);
nor U9759 (N_9759,N_9289,N_9177);
and U9760 (N_9760,N_9100,N_9243);
or U9761 (N_9761,N_9258,N_9045);
xnor U9762 (N_9762,N_9069,N_9415);
or U9763 (N_9763,N_9064,N_9441);
xnor U9764 (N_9764,N_9197,N_9141);
nor U9765 (N_9765,N_9333,N_9050);
xor U9766 (N_9766,N_9219,N_9143);
xnor U9767 (N_9767,N_9151,N_9026);
and U9768 (N_9768,N_9303,N_9197);
or U9769 (N_9769,N_9251,N_9239);
nor U9770 (N_9770,N_9469,N_9402);
and U9771 (N_9771,N_9094,N_9015);
nand U9772 (N_9772,N_9498,N_9323);
nor U9773 (N_9773,N_9434,N_9355);
nand U9774 (N_9774,N_9448,N_9417);
nor U9775 (N_9775,N_9221,N_9050);
and U9776 (N_9776,N_9056,N_9175);
nor U9777 (N_9777,N_9065,N_9434);
and U9778 (N_9778,N_9437,N_9154);
and U9779 (N_9779,N_9442,N_9183);
nor U9780 (N_9780,N_9442,N_9376);
and U9781 (N_9781,N_9427,N_9064);
nand U9782 (N_9782,N_9171,N_9336);
or U9783 (N_9783,N_9064,N_9236);
and U9784 (N_9784,N_9265,N_9229);
xnor U9785 (N_9785,N_9384,N_9136);
xor U9786 (N_9786,N_9431,N_9138);
nand U9787 (N_9787,N_9113,N_9367);
nand U9788 (N_9788,N_9169,N_9385);
or U9789 (N_9789,N_9231,N_9201);
xor U9790 (N_9790,N_9157,N_9000);
nor U9791 (N_9791,N_9282,N_9493);
nand U9792 (N_9792,N_9301,N_9017);
or U9793 (N_9793,N_9181,N_9380);
or U9794 (N_9794,N_9012,N_9449);
nor U9795 (N_9795,N_9071,N_9356);
nand U9796 (N_9796,N_9180,N_9417);
and U9797 (N_9797,N_9247,N_9437);
xor U9798 (N_9798,N_9228,N_9185);
xor U9799 (N_9799,N_9467,N_9127);
nand U9800 (N_9800,N_9165,N_9018);
nand U9801 (N_9801,N_9005,N_9472);
nand U9802 (N_9802,N_9119,N_9033);
or U9803 (N_9803,N_9489,N_9316);
and U9804 (N_9804,N_9271,N_9424);
xnor U9805 (N_9805,N_9462,N_9084);
or U9806 (N_9806,N_9439,N_9338);
xnor U9807 (N_9807,N_9061,N_9117);
nor U9808 (N_9808,N_9058,N_9210);
or U9809 (N_9809,N_9269,N_9308);
nor U9810 (N_9810,N_9306,N_9065);
or U9811 (N_9811,N_9031,N_9321);
nor U9812 (N_9812,N_9068,N_9436);
nand U9813 (N_9813,N_9073,N_9256);
or U9814 (N_9814,N_9448,N_9456);
xor U9815 (N_9815,N_9498,N_9160);
xor U9816 (N_9816,N_9137,N_9112);
nor U9817 (N_9817,N_9027,N_9383);
and U9818 (N_9818,N_9193,N_9021);
nor U9819 (N_9819,N_9255,N_9085);
or U9820 (N_9820,N_9325,N_9446);
and U9821 (N_9821,N_9182,N_9259);
nor U9822 (N_9822,N_9244,N_9047);
or U9823 (N_9823,N_9382,N_9302);
xor U9824 (N_9824,N_9331,N_9209);
or U9825 (N_9825,N_9421,N_9315);
xnor U9826 (N_9826,N_9287,N_9389);
or U9827 (N_9827,N_9443,N_9355);
nand U9828 (N_9828,N_9272,N_9101);
xor U9829 (N_9829,N_9116,N_9454);
or U9830 (N_9830,N_9013,N_9235);
and U9831 (N_9831,N_9295,N_9150);
nor U9832 (N_9832,N_9008,N_9476);
nor U9833 (N_9833,N_9130,N_9010);
or U9834 (N_9834,N_9483,N_9297);
or U9835 (N_9835,N_9361,N_9268);
nor U9836 (N_9836,N_9242,N_9168);
nor U9837 (N_9837,N_9193,N_9038);
xnor U9838 (N_9838,N_9106,N_9101);
nand U9839 (N_9839,N_9323,N_9106);
and U9840 (N_9840,N_9445,N_9243);
nor U9841 (N_9841,N_9384,N_9103);
and U9842 (N_9842,N_9403,N_9353);
nand U9843 (N_9843,N_9147,N_9257);
and U9844 (N_9844,N_9302,N_9459);
nor U9845 (N_9845,N_9332,N_9462);
xnor U9846 (N_9846,N_9118,N_9235);
or U9847 (N_9847,N_9225,N_9406);
nor U9848 (N_9848,N_9157,N_9136);
or U9849 (N_9849,N_9128,N_9080);
xor U9850 (N_9850,N_9230,N_9232);
nor U9851 (N_9851,N_9187,N_9180);
and U9852 (N_9852,N_9125,N_9422);
nand U9853 (N_9853,N_9144,N_9223);
and U9854 (N_9854,N_9469,N_9331);
and U9855 (N_9855,N_9357,N_9309);
nor U9856 (N_9856,N_9293,N_9279);
xnor U9857 (N_9857,N_9155,N_9347);
xor U9858 (N_9858,N_9254,N_9206);
or U9859 (N_9859,N_9207,N_9160);
nor U9860 (N_9860,N_9334,N_9138);
nor U9861 (N_9861,N_9034,N_9418);
or U9862 (N_9862,N_9491,N_9025);
and U9863 (N_9863,N_9163,N_9479);
xnor U9864 (N_9864,N_9290,N_9480);
nand U9865 (N_9865,N_9097,N_9274);
or U9866 (N_9866,N_9047,N_9117);
or U9867 (N_9867,N_9478,N_9127);
or U9868 (N_9868,N_9210,N_9258);
and U9869 (N_9869,N_9187,N_9249);
nor U9870 (N_9870,N_9235,N_9334);
and U9871 (N_9871,N_9094,N_9077);
nor U9872 (N_9872,N_9158,N_9008);
or U9873 (N_9873,N_9249,N_9467);
nand U9874 (N_9874,N_9294,N_9476);
and U9875 (N_9875,N_9256,N_9349);
nand U9876 (N_9876,N_9175,N_9248);
xnor U9877 (N_9877,N_9428,N_9331);
nor U9878 (N_9878,N_9453,N_9080);
or U9879 (N_9879,N_9284,N_9076);
nor U9880 (N_9880,N_9002,N_9225);
xor U9881 (N_9881,N_9106,N_9496);
or U9882 (N_9882,N_9233,N_9089);
xor U9883 (N_9883,N_9113,N_9412);
and U9884 (N_9884,N_9370,N_9395);
xnor U9885 (N_9885,N_9481,N_9244);
and U9886 (N_9886,N_9050,N_9321);
or U9887 (N_9887,N_9364,N_9018);
nand U9888 (N_9888,N_9340,N_9360);
nand U9889 (N_9889,N_9212,N_9034);
nand U9890 (N_9890,N_9464,N_9069);
nor U9891 (N_9891,N_9329,N_9051);
nand U9892 (N_9892,N_9000,N_9146);
nor U9893 (N_9893,N_9091,N_9104);
xnor U9894 (N_9894,N_9249,N_9496);
and U9895 (N_9895,N_9017,N_9494);
nor U9896 (N_9896,N_9166,N_9277);
and U9897 (N_9897,N_9227,N_9164);
or U9898 (N_9898,N_9048,N_9004);
or U9899 (N_9899,N_9089,N_9077);
or U9900 (N_9900,N_9257,N_9153);
or U9901 (N_9901,N_9332,N_9335);
and U9902 (N_9902,N_9468,N_9085);
and U9903 (N_9903,N_9340,N_9121);
and U9904 (N_9904,N_9155,N_9203);
xor U9905 (N_9905,N_9116,N_9030);
or U9906 (N_9906,N_9083,N_9121);
xnor U9907 (N_9907,N_9076,N_9495);
xnor U9908 (N_9908,N_9436,N_9378);
xnor U9909 (N_9909,N_9438,N_9106);
xor U9910 (N_9910,N_9457,N_9185);
or U9911 (N_9911,N_9474,N_9240);
xnor U9912 (N_9912,N_9174,N_9240);
nor U9913 (N_9913,N_9027,N_9268);
and U9914 (N_9914,N_9119,N_9302);
nand U9915 (N_9915,N_9392,N_9335);
nand U9916 (N_9916,N_9264,N_9415);
nor U9917 (N_9917,N_9243,N_9108);
nand U9918 (N_9918,N_9395,N_9013);
and U9919 (N_9919,N_9465,N_9386);
nand U9920 (N_9920,N_9088,N_9009);
or U9921 (N_9921,N_9254,N_9334);
xor U9922 (N_9922,N_9114,N_9353);
or U9923 (N_9923,N_9406,N_9017);
and U9924 (N_9924,N_9061,N_9392);
nor U9925 (N_9925,N_9160,N_9126);
and U9926 (N_9926,N_9471,N_9053);
or U9927 (N_9927,N_9169,N_9473);
and U9928 (N_9928,N_9104,N_9013);
nand U9929 (N_9929,N_9244,N_9283);
nand U9930 (N_9930,N_9289,N_9176);
nor U9931 (N_9931,N_9006,N_9483);
nand U9932 (N_9932,N_9043,N_9389);
nand U9933 (N_9933,N_9046,N_9039);
or U9934 (N_9934,N_9457,N_9188);
nand U9935 (N_9935,N_9265,N_9003);
xnor U9936 (N_9936,N_9327,N_9437);
nand U9937 (N_9937,N_9470,N_9083);
and U9938 (N_9938,N_9029,N_9256);
or U9939 (N_9939,N_9314,N_9090);
nor U9940 (N_9940,N_9480,N_9018);
and U9941 (N_9941,N_9362,N_9075);
and U9942 (N_9942,N_9483,N_9312);
and U9943 (N_9943,N_9000,N_9362);
xnor U9944 (N_9944,N_9385,N_9410);
nand U9945 (N_9945,N_9271,N_9028);
or U9946 (N_9946,N_9226,N_9284);
and U9947 (N_9947,N_9213,N_9166);
nor U9948 (N_9948,N_9428,N_9054);
and U9949 (N_9949,N_9271,N_9225);
or U9950 (N_9950,N_9117,N_9026);
xor U9951 (N_9951,N_9409,N_9429);
and U9952 (N_9952,N_9378,N_9235);
nand U9953 (N_9953,N_9428,N_9213);
nor U9954 (N_9954,N_9138,N_9413);
xor U9955 (N_9955,N_9254,N_9352);
nand U9956 (N_9956,N_9149,N_9289);
xnor U9957 (N_9957,N_9088,N_9444);
nand U9958 (N_9958,N_9468,N_9182);
nor U9959 (N_9959,N_9185,N_9035);
and U9960 (N_9960,N_9472,N_9467);
xnor U9961 (N_9961,N_9043,N_9477);
and U9962 (N_9962,N_9398,N_9203);
nand U9963 (N_9963,N_9028,N_9314);
or U9964 (N_9964,N_9260,N_9320);
nand U9965 (N_9965,N_9140,N_9350);
and U9966 (N_9966,N_9359,N_9332);
xor U9967 (N_9967,N_9393,N_9037);
or U9968 (N_9968,N_9182,N_9368);
and U9969 (N_9969,N_9037,N_9407);
or U9970 (N_9970,N_9083,N_9478);
nor U9971 (N_9971,N_9060,N_9317);
nor U9972 (N_9972,N_9089,N_9043);
nor U9973 (N_9973,N_9108,N_9414);
nor U9974 (N_9974,N_9094,N_9119);
nor U9975 (N_9975,N_9270,N_9212);
or U9976 (N_9976,N_9085,N_9304);
or U9977 (N_9977,N_9383,N_9168);
and U9978 (N_9978,N_9349,N_9486);
or U9979 (N_9979,N_9014,N_9147);
and U9980 (N_9980,N_9035,N_9468);
and U9981 (N_9981,N_9279,N_9424);
and U9982 (N_9982,N_9492,N_9144);
xor U9983 (N_9983,N_9461,N_9070);
xnor U9984 (N_9984,N_9250,N_9085);
or U9985 (N_9985,N_9402,N_9226);
or U9986 (N_9986,N_9233,N_9071);
xnor U9987 (N_9987,N_9144,N_9149);
nand U9988 (N_9988,N_9179,N_9077);
xnor U9989 (N_9989,N_9367,N_9259);
xnor U9990 (N_9990,N_9224,N_9340);
or U9991 (N_9991,N_9433,N_9164);
or U9992 (N_9992,N_9040,N_9366);
or U9993 (N_9993,N_9425,N_9401);
nand U9994 (N_9994,N_9349,N_9104);
nor U9995 (N_9995,N_9263,N_9180);
and U9996 (N_9996,N_9388,N_9247);
xnor U9997 (N_9997,N_9103,N_9482);
nor U9998 (N_9998,N_9204,N_9405);
or U9999 (N_9999,N_9319,N_9087);
xor U10000 (N_10000,N_9715,N_9691);
and U10001 (N_10001,N_9783,N_9719);
xnor U10002 (N_10002,N_9577,N_9571);
nand U10003 (N_10003,N_9982,N_9600);
and U10004 (N_10004,N_9500,N_9739);
nand U10005 (N_10005,N_9697,N_9879);
nor U10006 (N_10006,N_9544,N_9661);
and U10007 (N_10007,N_9798,N_9606);
and U10008 (N_10008,N_9504,N_9550);
xnor U10009 (N_10009,N_9682,N_9732);
or U10010 (N_10010,N_9973,N_9863);
nor U10011 (N_10011,N_9918,N_9935);
or U10012 (N_10012,N_9887,N_9727);
nor U10013 (N_10013,N_9745,N_9842);
or U10014 (N_10014,N_9692,N_9969);
and U10015 (N_10015,N_9924,N_9898);
nor U10016 (N_10016,N_9743,N_9911);
and U10017 (N_10017,N_9940,N_9519);
or U10018 (N_10018,N_9567,N_9736);
nor U10019 (N_10019,N_9582,N_9938);
nand U10020 (N_10020,N_9520,N_9585);
xor U10021 (N_10021,N_9716,N_9978);
xnor U10022 (N_10022,N_9722,N_9613);
nor U10023 (N_10023,N_9654,N_9584);
nor U10024 (N_10024,N_9547,N_9649);
nand U10025 (N_10025,N_9781,N_9916);
and U10026 (N_10026,N_9862,N_9787);
nand U10027 (N_10027,N_9737,N_9501);
xor U10028 (N_10028,N_9778,N_9912);
xnor U10029 (N_10029,N_9677,N_9789);
nand U10030 (N_10030,N_9891,N_9833);
xor U10031 (N_10031,N_9994,N_9826);
nand U10032 (N_10032,N_9535,N_9557);
nor U10033 (N_10033,N_9770,N_9983);
or U10034 (N_10034,N_9925,N_9937);
nor U10035 (N_10035,N_9603,N_9839);
xor U10036 (N_10036,N_9946,N_9533);
and U10037 (N_10037,N_9922,N_9755);
nand U10038 (N_10038,N_9871,N_9694);
nand U10039 (N_10039,N_9805,N_9549);
nand U10040 (N_10040,N_9790,N_9655);
nor U10041 (N_10041,N_9966,N_9810);
and U10042 (N_10042,N_9629,N_9553);
and U10043 (N_10043,N_9536,N_9792);
nand U10044 (N_10044,N_9950,N_9534);
or U10045 (N_10045,N_9506,N_9985);
xor U10046 (N_10046,N_9611,N_9769);
and U10047 (N_10047,N_9546,N_9929);
and U10048 (N_10048,N_9517,N_9949);
nand U10049 (N_10049,N_9788,N_9742);
or U10050 (N_10050,N_9927,N_9815);
and U10051 (N_10051,N_9644,N_9817);
or U10052 (N_10052,N_9882,N_9643);
or U10053 (N_10053,N_9884,N_9888);
or U10054 (N_10054,N_9897,N_9873);
or U10055 (N_10055,N_9867,N_9824);
or U10056 (N_10056,N_9576,N_9690);
or U10057 (N_10057,N_9541,N_9712);
and U10058 (N_10058,N_9754,N_9591);
or U10059 (N_10059,N_9797,N_9895);
nand U10060 (N_10060,N_9751,N_9799);
and U10061 (N_10061,N_9726,N_9931);
and U10062 (N_10062,N_9944,N_9532);
xor U10063 (N_10063,N_9740,N_9572);
or U10064 (N_10064,N_9568,N_9669);
and U10065 (N_10065,N_9951,N_9926);
nor U10066 (N_10066,N_9673,N_9723);
nor U10067 (N_10067,N_9832,N_9821);
and U10068 (N_10068,N_9554,N_9779);
nand U10069 (N_10069,N_9999,N_9609);
or U10070 (N_10070,N_9594,N_9791);
nor U10071 (N_10071,N_9820,N_9988);
nand U10072 (N_10072,N_9957,N_9593);
nor U10073 (N_10073,N_9637,N_9590);
and U10074 (N_10074,N_9843,N_9774);
nor U10075 (N_10075,N_9616,N_9914);
or U10076 (N_10076,N_9980,N_9991);
xor U10077 (N_10077,N_9858,N_9809);
and U10078 (N_10078,N_9869,N_9777);
nor U10079 (N_10079,N_9563,N_9639);
or U10080 (N_10080,N_9962,N_9538);
and U10081 (N_10081,N_9556,N_9967);
or U10082 (N_10082,N_9640,N_9756);
and U10083 (N_10083,N_9623,N_9685);
nor U10084 (N_10084,N_9921,N_9525);
or U10085 (N_10085,N_9984,N_9959);
nor U10086 (N_10086,N_9527,N_9717);
xor U10087 (N_10087,N_9964,N_9886);
nor U10088 (N_10088,N_9972,N_9860);
xnor U10089 (N_10089,N_9711,N_9877);
nand U10090 (N_10090,N_9808,N_9857);
nor U10091 (N_10091,N_9859,N_9955);
and U10092 (N_10092,N_9581,N_9829);
or U10093 (N_10093,N_9656,N_9958);
xor U10094 (N_10094,N_9870,N_9846);
and U10095 (N_10095,N_9678,N_9511);
xor U10096 (N_10096,N_9695,N_9622);
or U10097 (N_10097,N_9725,N_9653);
nand U10098 (N_10098,N_9811,N_9773);
nor U10099 (N_10099,N_9936,N_9713);
and U10100 (N_10100,N_9705,N_9990);
and U10101 (N_10101,N_9981,N_9865);
nor U10102 (N_10102,N_9845,N_9698);
xnor U10103 (N_10103,N_9907,N_9971);
xor U10104 (N_10104,N_9813,N_9841);
xnor U10105 (N_10105,N_9632,N_9524);
xor U10106 (N_10106,N_9825,N_9834);
or U10107 (N_10107,N_9552,N_9665);
xnor U10108 (N_10108,N_9741,N_9529);
nor U10109 (N_10109,N_9744,N_9646);
and U10110 (N_10110,N_9560,N_9776);
xor U10111 (N_10111,N_9531,N_9802);
xor U10112 (N_10112,N_9615,N_9509);
nor U10113 (N_10113,N_9618,N_9848);
xnor U10114 (N_10114,N_9861,N_9566);
nand U10115 (N_10115,N_9793,N_9747);
or U10116 (N_10116,N_9522,N_9555);
and U10117 (N_10117,N_9619,N_9565);
xnor U10118 (N_10118,N_9704,N_9672);
or U10119 (N_10119,N_9823,N_9666);
xnor U10120 (N_10120,N_9952,N_9617);
and U10121 (N_10121,N_9947,N_9683);
or U10122 (N_10122,N_9707,N_9763);
and U10123 (N_10123,N_9610,N_9923);
or U10124 (N_10124,N_9956,N_9700);
or U10125 (N_10125,N_9749,N_9510);
nand U10126 (N_10126,N_9892,N_9784);
or U10127 (N_10127,N_9574,N_9729);
or U10128 (N_10128,N_9919,N_9597);
xnor U10129 (N_10129,N_9573,N_9569);
nand U10130 (N_10130,N_9598,N_9807);
or U10131 (N_10131,N_9900,N_9987);
xor U10132 (N_10132,N_9814,N_9976);
xor U10133 (N_10133,N_9889,N_9890);
or U10134 (N_10134,N_9831,N_9875);
nand U10135 (N_10135,N_9589,N_9735);
xor U10136 (N_10136,N_9954,N_9696);
xor U10137 (N_10137,N_9915,N_9641);
nor U10138 (N_10138,N_9904,N_9782);
and U10139 (N_10139,N_9688,N_9633);
nand U10140 (N_10140,N_9515,N_9930);
xnor U10141 (N_10141,N_9605,N_9934);
and U10142 (N_10142,N_9852,N_9753);
and U10143 (N_10143,N_9965,N_9562);
nand U10144 (N_10144,N_9849,N_9801);
xor U10145 (N_10145,N_9503,N_9680);
nor U10146 (N_10146,N_9868,N_9724);
and U10147 (N_10147,N_9939,N_9986);
nand U10148 (N_10148,N_9681,N_9595);
nor U10149 (N_10149,N_9561,N_9775);
xnor U10150 (N_10150,N_9539,N_9658);
xor U10151 (N_10151,N_9850,N_9670);
nor U10152 (N_10152,N_9507,N_9602);
or U10153 (N_10153,N_9804,N_9762);
and U10154 (N_10154,N_9620,N_9627);
and U10155 (N_10155,N_9731,N_9837);
or U10156 (N_10156,N_9878,N_9866);
xor U10157 (N_10157,N_9812,N_9634);
nor U10158 (N_10158,N_9883,N_9730);
nand U10159 (N_10159,N_9827,N_9570);
xnor U10160 (N_10160,N_9578,N_9512);
and U10161 (N_10161,N_9785,N_9702);
nand U10162 (N_10162,N_9943,N_9575);
nand U10163 (N_10163,N_9652,N_9899);
or U10164 (N_10164,N_9953,N_9945);
nor U10165 (N_10165,N_9701,N_9601);
nor U10166 (N_10166,N_9638,N_9662);
and U10167 (N_10167,N_9709,N_9625);
nand U10168 (N_10168,N_9989,N_9963);
and U10169 (N_10169,N_9767,N_9995);
xnor U10170 (N_10170,N_9671,N_9579);
or U10171 (N_10171,N_9803,N_9559);
nand U10172 (N_10172,N_9961,N_9720);
or U10173 (N_10173,N_9548,N_9614);
nand U10174 (N_10174,N_9816,N_9772);
xor U10175 (N_10175,N_9795,N_9822);
nand U10176 (N_10176,N_9663,N_9800);
or U10177 (N_10177,N_9583,N_9628);
nand U10178 (N_10178,N_9970,N_9657);
or U10179 (N_10179,N_9942,N_9847);
nand U10180 (N_10180,N_9830,N_9513);
nor U10181 (N_10181,N_9604,N_9645);
xnor U10182 (N_10182,N_9505,N_9881);
nor U10183 (N_10183,N_9855,N_9896);
xor U10184 (N_10184,N_9844,N_9708);
xnor U10185 (N_10185,N_9818,N_9684);
nor U10186 (N_10186,N_9530,N_9718);
xor U10187 (N_10187,N_9901,N_9710);
nor U10188 (N_10188,N_9968,N_9838);
xor U10189 (N_10189,N_9612,N_9693);
nand U10190 (N_10190,N_9521,N_9920);
or U10191 (N_10191,N_9746,N_9748);
nor U10192 (N_10192,N_9586,N_9840);
nor U10193 (N_10193,N_9659,N_9523);
xor U10194 (N_10194,N_9948,N_9906);
and U10195 (N_10195,N_9721,N_9771);
and U10196 (N_10196,N_9836,N_9630);
nand U10197 (N_10197,N_9979,N_9508);
xor U10198 (N_10198,N_9786,N_9624);
and U10199 (N_10199,N_9806,N_9941);
xnor U10200 (N_10200,N_9766,N_9765);
or U10201 (N_10201,N_9706,N_9768);
nand U10202 (N_10202,N_9545,N_9993);
nor U10203 (N_10203,N_9679,N_9856);
and U10204 (N_10204,N_9752,N_9526);
and U10205 (N_10205,N_9880,N_9917);
or U10206 (N_10206,N_9757,N_9885);
nand U10207 (N_10207,N_9794,N_9893);
and U10208 (N_10208,N_9908,N_9699);
nor U10209 (N_10209,N_9905,N_9997);
and U10210 (N_10210,N_9872,N_9703);
and U10211 (N_10211,N_9760,N_9642);
nand U10212 (N_10212,N_9902,N_9714);
nor U10213 (N_10213,N_9728,N_9607);
nand U10214 (N_10214,N_9733,N_9631);
xor U10215 (N_10215,N_9758,N_9502);
xor U10216 (N_10216,N_9608,N_9580);
nand U10217 (N_10217,N_9996,N_9668);
nand U10218 (N_10218,N_9780,N_9516);
xnor U10219 (N_10219,N_9528,N_9974);
and U10220 (N_10220,N_9635,N_9854);
nor U10221 (N_10221,N_9626,N_9759);
nand U10222 (N_10222,N_9761,N_9542);
nand U10223 (N_10223,N_9588,N_9551);
nand U10224 (N_10224,N_9636,N_9960);
or U10225 (N_10225,N_9664,N_9998);
or U10226 (N_10226,N_9853,N_9819);
nand U10227 (N_10227,N_9592,N_9764);
xor U10228 (N_10228,N_9599,N_9992);
xnor U10229 (N_10229,N_9894,N_9828);
and U10230 (N_10230,N_9933,N_9909);
or U10231 (N_10231,N_9734,N_9667);
nand U10232 (N_10232,N_9648,N_9587);
nor U10233 (N_10233,N_9537,N_9876);
nor U10234 (N_10234,N_9910,N_9913);
nand U10235 (N_10235,N_9675,N_9518);
nor U10236 (N_10236,N_9835,N_9650);
nor U10237 (N_10237,N_9874,N_9738);
xnor U10238 (N_10238,N_9660,N_9851);
and U10239 (N_10239,N_9621,N_9932);
nor U10240 (N_10240,N_9977,N_9564);
nor U10241 (N_10241,N_9674,N_9687);
nor U10242 (N_10242,N_9689,N_9676);
xor U10243 (N_10243,N_9864,N_9540);
and U10244 (N_10244,N_9686,N_9903);
nand U10245 (N_10245,N_9647,N_9596);
nor U10246 (N_10246,N_9543,N_9750);
and U10247 (N_10247,N_9975,N_9514);
and U10248 (N_10248,N_9558,N_9928);
nand U10249 (N_10249,N_9796,N_9651);
or U10250 (N_10250,N_9514,N_9799);
and U10251 (N_10251,N_9702,N_9971);
and U10252 (N_10252,N_9899,N_9915);
and U10253 (N_10253,N_9785,N_9504);
xor U10254 (N_10254,N_9927,N_9866);
nand U10255 (N_10255,N_9530,N_9589);
nand U10256 (N_10256,N_9588,N_9544);
or U10257 (N_10257,N_9806,N_9504);
xnor U10258 (N_10258,N_9736,N_9657);
nand U10259 (N_10259,N_9701,N_9505);
nand U10260 (N_10260,N_9956,N_9958);
and U10261 (N_10261,N_9510,N_9642);
or U10262 (N_10262,N_9590,N_9670);
nor U10263 (N_10263,N_9857,N_9933);
or U10264 (N_10264,N_9549,N_9630);
and U10265 (N_10265,N_9979,N_9899);
nor U10266 (N_10266,N_9832,N_9989);
and U10267 (N_10267,N_9886,N_9845);
or U10268 (N_10268,N_9926,N_9838);
nor U10269 (N_10269,N_9990,N_9748);
nor U10270 (N_10270,N_9737,N_9923);
nand U10271 (N_10271,N_9617,N_9711);
xnor U10272 (N_10272,N_9634,N_9626);
or U10273 (N_10273,N_9885,N_9561);
or U10274 (N_10274,N_9697,N_9883);
or U10275 (N_10275,N_9738,N_9989);
xor U10276 (N_10276,N_9680,N_9822);
xor U10277 (N_10277,N_9954,N_9951);
or U10278 (N_10278,N_9980,N_9663);
or U10279 (N_10279,N_9897,N_9631);
xor U10280 (N_10280,N_9564,N_9684);
xor U10281 (N_10281,N_9614,N_9619);
and U10282 (N_10282,N_9815,N_9768);
and U10283 (N_10283,N_9552,N_9810);
xor U10284 (N_10284,N_9671,N_9700);
nor U10285 (N_10285,N_9681,N_9947);
xnor U10286 (N_10286,N_9801,N_9566);
xnor U10287 (N_10287,N_9612,N_9666);
nand U10288 (N_10288,N_9720,N_9920);
and U10289 (N_10289,N_9937,N_9868);
or U10290 (N_10290,N_9734,N_9995);
and U10291 (N_10291,N_9763,N_9857);
nor U10292 (N_10292,N_9867,N_9666);
nor U10293 (N_10293,N_9716,N_9662);
nand U10294 (N_10294,N_9849,N_9640);
or U10295 (N_10295,N_9588,N_9886);
and U10296 (N_10296,N_9957,N_9930);
or U10297 (N_10297,N_9672,N_9620);
nor U10298 (N_10298,N_9631,N_9984);
nand U10299 (N_10299,N_9666,N_9813);
nand U10300 (N_10300,N_9881,N_9947);
xnor U10301 (N_10301,N_9868,N_9606);
nand U10302 (N_10302,N_9558,N_9904);
or U10303 (N_10303,N_9733,N_9564);
nand U10304 (N_10304,N_9866,N_9510);
nor U10305 (N_10305,N_9899,N_9780);
nor U10306 (N_10306,N_9701,N_9775);
nor U10307 (N_10307,N_9501,N_9531);
xnor U10308 (N_10308,N_9717,N_9685);
or U10309 (N_10309,N_9686,N_9748);
and U10310 (N_10310,N_9644,N_9794);
xor U10311 (N_10311,N_9898,N_9754);
or U10312 (N_10312,N_9766,N_9545);
xor U10313 (N_10313,N_9901,N_9980);
xnor U10314 (N_10314,N_9970,N_9681);
and U10315 (N_10315,N_9731,N_9624);
or U10316 (N_10316,N_9522,N_9747);
and U10317 (N_10317,N_9735,N_9772);
xnor U10318 (N_10318,N_9939,N_9529);
or U10319 (N_10319,N_9869,N_9741);
or U10320 (N_10320,N_9664,N_9520);
or U10321 (N_10321,N_9607,N_9755);
nand U10322 (N_10322,N_9898,N_9842);
and U10323 (N_10323,N_9698,N_9899);
or U10324 (N_10324,N_9622,N_9888);
or U10325 (N_10325,N_9767,N_9642);
nor U10326 (N_10326,N_9739,N_9964);
or U10327 (N_10327,N_9636,N_9897);
and U10328 (N_10328,N_9599,N_9601);
and U10329 (N_10329,N_9993,N_9705);
xor U10330 (N_10330,N_9696,N_9657);
nor U10331 (N_10331,N_9701,N_9602);
nor U10332 (N_10332,N_9645,N_9715);
nand U10333 (N_10333,N_9612,N_9740);
nand U10334 (N_10334,N_9875,N_9776);
or U10335 (N_10335,N_9692,N_9735);
and U10336 (N_10336,N_9641,N_9677);
and U10337 (N_10337,N_9620,N_9656);
or U10338 (N_10338,N_9579,N_9607);
xnor U10339 (N_10339,N_9824,N_9796);
nand U10340 (N_10340,N_9582,N_9511);
nor U10341 (N_10341,N_9711,N_9574);
nor U10342 (N_10342,N_9950,N_9768);
and U10343 (N_10343,N_9772,N_9908);
xor U10344 (N_10344,N_9753,N_9641);
nand U10345 (N_10345,N_9800,N_9674);
nor U10346 (N_10346,N_9755,N_9756);
nor U10347 (N_10347,N_9910,N_9800);
nand U10348 (N_10348,N_9836,N_9694);
or U10349 (N_10349,N_9865,N_9715);
nor U10350 (N_10350,N_9684,N_9968);
nor U10351 (N_10351,N_9740,N_9939);
or U10352 (N_10352,N_9608,N_9985);
xor U10353 (N_10353,N_9872,N_9755);
nor U10354 (N_10354,N_9902,N_9797);
nand U10355 (N_10355,N_9657,N_9877);
nor U10356 (N_10356,N_9867,N_9664);
nand U10357 (N_10357,N_9616,N_9955);
and U10358 (N_10358,N_9805,N_9764);
xnor U10359 (N_10359,N_9691,N_9729);
xor U10360 (N_10360,N_9532,N_9670);
or U10361 (N_10361,N_9510,N_9806);
and U10362 (N_10362,N_9961,N_9898);
and U10363 (N_10363,N_9808,N_9806);
or U10364 (N_10364,N_9679,N_9620);
and U10365 (N_10365,N_9753,N_9515);
nor U10366 (N_10366,N_9620,N_9531);
or U10367 (N_10367,N_9525,N_9633);
or U10368 (N_10368,N_9897,N_9989);
and U10369 (N_10369,N_9591,N_9558);
and U10370 (N_10370,N_9707,N_9948);
and U10371 (N_10371,N_9999,N_9684);
nor U10372 (N_10372,N_9779,N_9527);
nor U10373 (N_10373,N_9980,N_9844);
xnor U10374 (N_10374,N_9841,N_9723);
nor U10375 (N_10375,N_9826,N_9698);
and U10376 (N_10376,N_9898,N_9565);
nor U10377 (N_10377,N_9577,N_9983);
nand U10378 (N_10378,N_9782,N_9999);
and U10379 (N_10379,N_9656,N_9773);
and U10380 (N_10380,N_9821,N_9691);
or U10381 (N_10381,N_9706,N_9908);
nor U10382 (N_10382,N_9783,N_9799);
nand U10383 (N_10383,N_9581,N_9722);
xnor U10384 (N_10384,N_9556,N_9853);
xnor U10385 (N_10385,N_9728,N_9553);
and U10386 (N_10386,N_9789,N_9757);
nand U10387 (N_10387,N_9518,N_9843);
or U10388 (N_10388,N_9508,N_9923);
nand U10389 (N_10389,N_9966,N_9814);
xnor U10390 (N_10390,N_9745,N_9549);
or U10391 (N_10391,N_9694,N_9968);
or U10392 (N_10392,N_9937,N_9766);
xnor U10393 (N_10393,N_9631,N_9746);
nand U10394 (N_10394,N_9628,N_9925);
or U10395 (N_10395,N_9633,N_9711);
xor U10396 (N_10396,N_9982,N_9613);
and U10397 (N_10397,N_9898,N_9513);
nor U10398 (N_10398,N_9916,N_9597);
nand U10399 (N_10399,N_9868,N_9732);
nor U10400 (N_10400,N_9788,N_9624);
and U10401 (N_10401,N_9659,N_9833);
or U10402 (N_10402,N_9657,N_9928);
nand U10403 (N_10403,N_9734,N_9928);
and U10404 (N_10404,N_9831,N_9705);
and U10405 (N_10405,N_9560,N_9747);
nor U10406 (N_10406,N_9885,N_9662);
xnor U10407 (N_10407,N_9971,N_9511);
xnor U10408 (N_10408,N_9761,N_9654);
xnor U10409 (N_10409,N_9552,N_9678);
and U10410 (N_10410,N_9656,N_9542);
and U10411 (N_10411,N_9751,N_9806);
nor U10412 (N_10412,N_9699,N_9907);
or U10413 (N_10413,N_9571,N_9696);
and U10414 (N_10414,N_9520,N_9875);
nand U10415 (N_10415,N_9827,N_9893);
xor U10416 (N_10416,N_9817,N_9762);
and U10417 (N_10417,N_9695,N_9694);
xnor U10418 (N_10418,N_9517,N_9888);
nor U10419 (N_10419,N_9608,N_9640);
or U10420 (N_10420,N_9839,N_9764);
nand U10421 (N_10421,N_9715,N_9760);
nand U10422 (N_10422,N_9695,N_9617);
or U10423 (N_10423,N_9896,N_9839);
nand U10424 (N_10424,N_9808,N_9739);
xor U10425 (N_10425,N_9764,N_9978);
or U10426 (N_10426,N_9656,N_9705);
and U10427 (N_10427,N_9739,N_9546);
or U10428 (N_10428,N_9905,N_9507);
xor U10429 (N_10429,N_9514,N_9597);
nor U10430 (N_10430,N_9586,N_9859);
and U10431 (N_10431,N_9517,N_9720);
nand U10432 (N_10432,N_9845,N_9561);
xor U10433 (N_10433,N_9777,N_9954);
xnor U10434 (N_10434,N_9853,N_9900);
nand U10435 (N_10435,N_9959,N_9569);
nor U10436 (N_10436,N_9646,N_9844);
nand U10437 (N_10437,N_9969,N_9655);
xor U10438 (N_10438,N_9955,N_9829);
xor U10439 (N_10439,N_9643,N_9507);
or U10440 (N_10440,N_9950,N_9588);
nor U10441 (N_10441,N_9565,N_9939);
and U10442 (N_10442,N_9647,N_9513);
nand U10443 (N_10443,N_9924,N_9949);
nor U10444 (N_10444,N_9640,N_9809);
xnor U10445 (N_10445,N_9776,N_9648);
and U10446 (N_10446,N_9552,N_9948);
or U10447 (N_10447,N_9591,N_9803);
nor U10448 (N_10448,N_9641,N_9929);
and U10449 (N_10449,N_9500,N_9932);
xnor U10450 (N_10450,N_9944,N_9877);
xnor U10451 (N_10451,N_9819,N_9647);
nor U10452 (N_10452,N_9746,N_9943);
nor U10453 (N_10453,N_9792,N_9563);
nor U10454 (N_10454,N_9674,N_9963);
nand U10455 (N_10455,N_9676,N_9500);
or U10456 (N_10456,N_9773,N_9698);
or U10457 (N_10457,N_9599,N_9716);
or U10458 (N_10458,N_9996,N_9786);
and U10459 (N_10459,N_9826,N_9516);
xor U10460 (N_10460,N_9721,N_9515);
and U10461 (N_10461,N_9723,N_9550);
nand U10462 (N_10462,N_9547,N_9965);
and U10463 (N_10463,N_9563,N_9904);
nand U10464 (N_10464,N_9708,N_9763);
or U10465 (N_10465,N_9867,N_9658);
or U10466 (N_10466,N_9634,N_9719);
and U10467 (N_10467,N_9894,N_9668);
nor U10468 (N_10468,N_9559,N_9906);
nor U10469 (N_10469,N_9827,N_9819);
and U10470 (N_10470,N_9665,N_9940);
xor U10471 (N_10471,N_9864,N_9692);
and U10472 (N_10472,N_9615,N_9836);
xor U10473 (N_10473,N_9783,N_9584);
nor U10474 (N_10474,N_9806,N_9988);
nor U10475 (N_10475,N_9904,N_9624);
nand U10476 (N_10476,N_9895,N_9762);
nand U10477 (N_10477,N_9712,N_9777);
or U10478 (N_10478,N_9575,N_9971);
and U10479 (N_10479,N_9615,N_9570);
nand U10480 (N_10480,N_9776,N_9527);
nand U10481 (N_10481,N_9994,N_9610);
and U10482 (N_10482,N_9616,N_9742);
or U10483 (N_10483,N_9805,N_9968);
nor U10484 (N_10484,N_9848,N_9673);
nor U10485 (N_10485,N_9960,N_9706);
or U10486 (N_10486,N_9747,N_9760);
nor U10487 (N_10487,N_9856,N_9924);
xor U10488 (N_10488,N_9845,N_9880);
or U10489 (N_10489,N_9797,N_9635);
and U10490 (N_10490,N_9945,N_9540);
nand U10491 (N_10491,N_9859,N_9862);
nand U10492 (N_10492,N_9833,N_9613);
xor U10493 (N_10493,N_9664,N_9877);
and U10494 (N_10494,N_9841,N_9552);
xnor U10495 (N_10495,N_9936,N_9891);
and U10496 (N_10496,N_9975,N_9610);
and U10497 (N_10497,N_9857,N_9696);
or U10498 (N_10498,N_9703,N_9609);
and U10499 (N_10499,N_9802,N_9576);
nand U10500 (N_10500,N_10205,N_10283);
nand U10501 (N_10501,N_10336,N_10015);
and U10502 (N_10502,N_10134,N_10268);
xnor U10503 (N_10503,N_10092,N_10369);
or U10504 (N_10504,N_10257,N_10400);
nor U10505 (N_10505,N_10351,N_10344);
nor U10506 (N_10506,N_10495,N_10364);
nor U10507 (N_10507,N_10222,N_10168);
or U10508 (N_10508,N_10408,N_10014);
nand U10509 (N_10509,N_10062,N_10010);
nor U10510 (N_10510,N_10278,N_10108);
or U10511 (N_10511,N_10035,N_10341);
xnor U10512 (N_10512,N_10183,N_10357);
or U10513 (N_10513,N_10102,N_10387);
and U10514 (N_10514,N_10325,N_10041);
xnor U10515 (N_10515,N_10398,N_10361);
nand U10516 (N_10516,N_10352,N_10424);
or U10517 (N_10517,N_10358,N_10499);
and U10518 (N_10518,N_10300,N_10438);
or U10519 (N_10519,N_10468,N_10294);
nand U10520 (N_10520,N_10101,N_10224);
or U10521 (N_10521,N_10025,N_10310);
nor U10522 (N_10522,N_10354,N_10078);
nand U10523 (N_10523,N_10086,N_10421);
and U10524 (N_10524,N_10251,N_10220);
nor U10525 (N_10525,N_10345,N_10428);
nand U10526 (N_10526,N_10083,N_10047);
xnor U10527 (N_10527,N_10489,N_10055);
or U10528 (N_10528,N_10353,N_10274);
nand U10529 (N_10529,N_10399,N_10296);
nand U10530 (N_10530,N_10256,N_10311);
nor U10531 (N_10531,N_10233,N_10116);
nor U10532 (N_10532,N_10470,N_10021);
and U10533 (N_10533,N_10415,N_10390);
or U10534 (N_10534,N_10243,N_10201);
or U10535 (N_10535,N_10330,N_10079);
nor U10536 (N_10536,N_10309,N_10263);
and U10537 (N_10537,N_10248,N_10136);
nor U10538 (N_10538,N_10488,N_10044);
and U10539 (N_10539,N_10405,N_10419);
xor U10540 (N_10540,N_10322,N_10163);
nand U10541 (N_10541,N_10223,N_10464);
nor U10542 (N_10542,N_10288,N_10362);
or U10543 (N_10543,N_10197,N_10125);
nand U10544 (N_10544,N_10249,N_10135);
and U10545 (N_10545,N_10377,N_10221);
nor U10546 (N_10546,N_10157,N_10308);
xnor U10547 (N_10547,N_10113,N_10122);
or U10548 (N_10548,N_10207,N_10187);
nor U10549 (N_10549,N_10131,N_10038);
nand U10550 (N_10550,N_10121,N_10462);
or U10551 (N_10551,N_10320,N_10191);
or U10552 (N_10552,N_10427,N_10127);
nor U10553 (N_10553,N_10384,N_10180);
nor U10554 (N_10554,N_10067,N_10472);
and U10555 (N_10555,N_10327,N_10313);
xor U10556 (N_10556,N_10279,N_10328);
and U10557 (N_10557,N_10453,N_10449);
or U10558 (N_10558,N_10392,N_10213);
nand U10559 (N_10559,N_10291,N_10396);
nor U10560 (N_10560,N_10228,N_10185);
xnor U10561 (N_10561,N_10171,N_10450);
nor U10562 (N_10562,N_10232,N_10217);
nor U10563 (N_10563,N_10199,N_10318);
and U10564 (N_10564,N_10496,N_10203);
nand U10565 (N_10565,N_10479,N_10343);
or U10566 (N_10566,N_10019,N_10052);
nor U10567 (N_10567,N_10467,N_10254);
nand U10568 (N_10568,N_10179,N_10093);
nand U10569 (N_10569,N_10323,N_10460);
nand U10570 (N_10570,N_10247,N_10103);
or U10571 (N_10571,N_10020,N_10258);
and U10572 (N_10572,N_10097,N_10487);
nand U10573 (N_10573,N_10246,N_10012);
nand U10574 (N_10574,N_10039,N_10461);
nand U10575 (N_10575,N_10099,N_10429);
xnor U10576 (N_10576,N_10435,N_10478);
and U10577 (N_10577,N_10034,N_10480);
nand U10578 (N_10578,N_10490,N_10030);
nand U10579 (N_10579,N_10446,N_10161);
nor U10580 (N_10580,N_10253,N_10264);
nor U10581 (N_10581,N_10080,N_10447);
and U10582 (N_10582,N_10418,N_10314);
xnor U10583 (N_10583,N_10089,N_10476);
nand U10584 (N_10584,N_10389,N_10365);
and U10585 (N_10585,N_10347,N_10188);
nor U10586 (N_10586,N_10219,N_10403);
or U10587 (N_10587,N_10494,N_10049);
nor U10588 (N_10588,N_10042,N_10349);
nand U10589 (N_10589,N_10401,N_10106);
nand U10590 (N_10590,N_10346,N_10053);
nor U10591 (N_10591,N_10360,N_10153);
and U10592 (N_10592,N_10481,N_10455);
xor U10593 (N_10593,N_10192,N_10027);
xor U10594 (N_10594,N_10209,N_10287);
nand U10595 (N_10595,N_10165,N_10022);
xor U10596 (N_10596,N_10404,N_10002);
nor U10597 (N_10597,N_10332,N_10011);
nand U10598 (N_10598,N_10214,N_10160);
xor U10599 (N_10599,N_10457,N_10059);
nor U10600 (N_10600,N_10230,N_10056);
or U10601 (N_10601,N_10120,N_10198);
xnor U10602 (N_10602,N_10226,N_10141);
xor U10603 (N_10603,N_10094,N_10193);
xor U10604 (N_10604,N_10211,N_10355);
xnor U10605 (N_10605,N_10497,N_10350);
xnor U10606 (N_10606,N_10043,N_10096);
nand U10607 (N_10607,N_10087,N_10437);
or U10608 (N_10608,N_10144,N_10172);
nor U10609 (N_10609,N_10442,N_10269);
or U10610 (N_10610,N_10498,N_10371);
or U10611 (N_10611,N_10471,N_10315);
and U10612 (N_10612,N_10182,N_10088);
nand U10613 (N_10613,N_10382,N_10169);
or U10614 (N_10614,N_10436,N_10110);
and U10615 (N_10615,N_10206,N_10340);
and U10616 (N_10616,N_10218,N_10434);
nor U10617 (N_10617,N_10175,N_10189);
and U10618 (N_10618,N_10037,N_10393);
xor U10619 (N_10619,N_10381,N_10054);
nand U10620 (N_10620,N_10149,N_10109);
nand U10621 (N_10621,N_10299,N_10372);
nand U10622 (N_10622,N_10319,N_10138);
or U10623 (N_10623,N_10081,N_10007);
or U10624 (N_10624,N_10284,N_10252);
or U10625 (N_10625,N_10276,N_10312);
nor U10626 (N_10626,N_10301,N_10298);
or U10627 (N_10627,N_10454,N_10317);
nor U10628 (N_10628,N_10376,N_10003);
nand U10629 (N_10629,N_10184,N_10281);
nand U10630 (N_10630,N_10431,N_10412);
nor U10631 (N_10631,N_10413,N_10245);
nor U10632 (N_10632,N_10237,N_10072);
xnor U10633 (N_10633,N_10273,N_10005);
nor U10634 (N_10634,N_10162,N_10225);
nor U10635 (N_10635,N_10366,N_10178);
nand U10636 (N_10636,N_10064,N_10045);
nor U10637 (N_10637,N_10235,N_10028);
nor U10638 (N_10638,N_10140,N_10114);
nor U10639 (N_10639,N_10255,N_10069);
and U10640 (N_10640,N_10440,N_10176);
or U10641 (N_10641,N_10417,N_10058);
nand U10642 (N_10642,N_10367,N_10290);
nand U10643 (N_10643,N_10491,N_10304);
xnor U10644 (N_10644,N_10166,N_10227);
or U10645 (N_10645,N_10482,N_10050);
or U10646 (N_10646,N_10448,N_10280);
or U10647 (N_10647,N_10137,N_10375);
nor U10648 (N_10648,N_10293,N_10402);
and U10649 (N_10649,N_10128,N_10167);
or U10650 (N_10650,N_10240,N_10456);
and U10651 (N_10651,N_10333,N_10445);
xnor U10652 (N_10652,N_10407,N_10238);
or U10653 (N_10653,N_10383,N_10076);
or U10654 (N_10654,N_10379,N_10229);
nor U10655 (N_10655,N_10380,N_10119);
xor U10656 (N_10656,N_10430,N_10395);
nor U10657 (N_10657,N_10316,N_10152);
xnor U10658 (N_10658,N_10117,N_10324);
or U10659 (N_10659,N_10443,N_10065);
or U10660 (N_10660,N_10164,N_10391);
nand U10661 (N_10661,N_10277,N_10406);
nor U10662 (N_10662,N_10029,N_10452);
nand U10663 (N_10663,N_10426,N_10334);
xnor U10664 (N_10664,N_10173,N_10373);
nand U10665 (N_10665,N_10126,N_10433);
xor U10666 (N_10666,N_10463,N_10051);
and U10667 (N_10667,N_10239,N_10331);
nand U10668 (N_10668,N_10008,N_10026);
or U10669 (N_10669,N_10104,N_10212);
or U10670 (N_10670,N_10196,N_10394);
nor U10671 (N_10671,N_10145,N_10174);
and U10672 (N_10672,N_10204,N_10105);
or U10673 (N_10673,N_10321,N_10326);
xnor U10674 (N_10674,N_10414,N_10484);
nand U10675 (N_10675,N_10474,N_10063);
or U10676 (N_10676,N_10465,N_10210);
and U10677 (N_10677,N_10285,N_10292);
and U10678 (N_10678,N_10057,N_10095);
nor U10679 (N_10679,N_10100,N_10425);
and U10680 (N_10680,N_10170,N_10143);
and U10681 (N_10681,N_10441,N_10148);
nor U10682 (N_10682,N_10388,N_10208);
xor U10683 (N_10683,N_10397,N_10270);
xor U10684 (N_10684,N_10335,N_10339);
xor U10685 (N_10685,N_10473,N_10216);
xor U10686 (N_10686,N_10459,N_10146);
nor U10687 (N_10687,N_10195,N_10082);
nand U10688 (N_10688,N_10156,N_10374);
or U10689 (N_10689,N_10337,N_10307);
xor U10690 (N_10690,N_10004,N_10023);
and U10691 (N_10691,N_10286,N_10018);
nor U10692 (N_10692,N_10244,N_10423);
and U10693 (N_10693,N_10439,N_10272);
xnor U10694 (N_10694,N_10370,N_10071);
nand U10695 (N_10695,N_10469,N_10031);
and U10696 (N_10696,N_10385,N_10139);
or U10697 (N_10697,N_10090,N_10066);
or U10698 (N_10698,N_10009,N_10420);
xor U10699 (N_10699,N_10061,N_10215);
nor U10700 (N_10700,N_10302,N_10202);
or U10701 (N_10701,N_10342,N_10150);
nor U10702 (N_10702,N_10260,N_10070);
xor U10703 (N_10703,N_10130,N_10036);
xnor U10704 (N_10704,N_10084,N_10085);
or U10705 (N_10705,N_10262,N_10118);
or U10706 (N_10706,N_10410,N_10475);
nand U10707 (N_10707,N_10068,N_10231);
nor U10708 (N_10708,N_10142,N_10123);
nor U10709 (N_10709,N_10261,N_10266);
nand U10710 (N_10710,N_10305,N_10024);
or U10711 (N_10711,N_10048,N_10451);
nand U10712 (N_10712,N_10483,N_10091);
nor U10713 (N_10713,N_10074,N_10073);
and U10714 (N_10714,N_10485,N_10098);
or U10715 (N_10715,N_10329,N_10409);
nand U10716 (N_10716,N_10242,N_10234);
nor U10717 (N_10717,N_10016,N_10107);
xnor U10718 (N_10718,N_10297,N_10416);
and U10719 (N_10719,N_10493,N_10458);
and U10720 (N_10720,N_10378,N_10303);
and U10721 (N_10721,N_10006,N_10432);
and U10722 (N_10722,N_10115,N_10075);
nand U10723 (N_10723,N_10111,N_10147);
nor U10724 (N_10724,N_10492,N_10154);
or U10725 (N_10725,N_10000,N_10060);
xnor U10726 (N_10726,N_10181,N_10158);
nor U10727 (N_10727,N_10275,N_10013);
nor U10728 (N_10728,N_10444,N_10259);
nor U10729 (N_10729,N_10368,N_10411);
or U10730 (N_10730,N_10236,N_10250);
and U10731 (N_10731,N_10356,N_10265);
xor U10732 (N_10732,N_10241,N_10177);
and U10733 (N_10733,N_10386,N_10338);
or U10734 (N_10734,N_10077,N_10133);
nand U10735 (N_10735,N_10040,N_10486);
nand U10736 (N_10736,N_10124,N_10190);
xor U10737 (N_10737,N_10200,N_10348);
nor U10738 (N_10738,N_10289,N_10194);
xnor U10739 (N_10739,N_10033,N_10363);
nand U10740 (N_10740,N_10132,N_10186);
or U10741 (N_10741,N_10001,N_10282);
or U10742 (N_10742,N_10129,N_10422);
nor U10743 (N_10743,N_10159,N_10267);
xor U10744 (N_10744,N_10017,N_10112);
and U10745 (N_10745,N_10151,N_10155);
nor U10746 (N_10746,N_10295,N_10359);
and U10747 (N_10747,N_10271,N_10046);
xor U10748 (N_10748,N_10306,N_10477);
nand U10749 (N_10749,N_10466,N_10032);
or U10750 (N_10750,N_10368,N_10062);
nand U10751 (N_10751,N_10127,N_10450);
nor U10752 (N_10752,N_10144,N_10493);
xor U10753 (N_10753,N_10310,N_10407);
and U10754 (N_10754,N_10176,N_10022);
or U10755 (N_10755,N_10443,N_10095);
nand U10756 (N_10756,N_10390,N_10498);
and U10757 (N_10757,N_10057,N_10243);
nand U10758 (N_10758,N_10479,N_10475);
or U10759 (N_10759,N_10272,N_10341);
and U10760 (N_10760,N_10304,N_10056);
xnor U10761 (N_10761,N_10307,N_10071);
nand U10762 (N_10762,N_10449,N_10344);
or U10763 (N_10763,N_10293,N_10046);
and U10764 (N_10764,N_10343,N_10333);
or U10765 (N_10765,N_10202,N_10323);
and U10766 (N_10766,N_10046,N_10487);
nand U10767 (N_10767,N_10085,N_10173);
nor U10768 (N_10768,N_10106,N_10192);
or U10769 (N_10769,N_10018,N_10498);
nand U10770 (N_10770,N_10191,N_10198);
nand U10771 (N_10771,N_10400,N_10444);
or U10772 (N_10772,N_10487,N_10442);
xor U10773 (N_10773,N_10198,N_10322);
xnor U10774 (N_10774,N_10401,N_10018);
nand U10775 (N_10775,N_10207,N_10142);
nand U10776 (N_10776,N_10171,N_10072);
nand U10777 (N_10777,N_10488,N_10439);
and U10778 (N_10778,N_10070,N_10363);
nor U10779 (N_10779,N_10362,N_10114);
and U10780 (N_10780,N_10301,N_10194);
nand U10781 (N_10781,N_10353,N_10182);
or U10782 (N_10782,N_10290,N_10481);
nand U10783 (N_10783,N_10244,N_10439);
nor U10784 (N_10784,N_10242,N_10161);
nor U10785 (N_10785,N_10338,N_10247);
xor U10786 (N_10786,N_10373,N_10117);
nand U10787 (N_10787,N_10089,N_10291);
nand U10788 (N_10788,N_10454,N_10462);
xor U10789 (N_10789,N_10001,N_10188);
nand U10790 (N_10790,N_10327,N_10067);
xor U10791 (N_10791,N_10344,N_10265);
and U10792 (N_10792,N_10394,N_10089);
nand U10793 (N_10793,N_10408,N_10092);
or U10794 (N_10794,N_10171,N_10332);
xor U10795 (N_10795,N_10388,N_10029);
or U10796 (N_10796,N_10214,N_10094);
nor U10797 (N_10797,N_10401,N_10413);
xnor U10798 (N_10798,N_10339,N_10492);
nor U10799 (N_10799,N_10402,N_10350);
nand U10800 (N_10800,N_10349,N_10295);
or U10801 (N_10801,N_10383,N_10415);
and U10802 (N_10802,N_10390,N_10109);
nor U10803 (N_10803,N_10240,N_10176);
and U10804 (N_10804,N_10342,N_10353);
and U10805 (N_10805,N_10010,N_10108);
nor U10806 (N_10806,N_10326,N_10413);
nand U10807 (N_10807,N_10355,N_10170);
or U10808 (N_10808,N_10415,N_10177);
and U10809 (N_10809,N_10017,N_10276);
or U10810 (N_10810,N_10433,N_10008);
nor U10811 (N_10811,N_10044,N_10081);
nand U10812 (N_10812,N_10187,N_10318);
or U10813 (N_10813,N_10384,N_10159);
and U10814 (N_10814,N_10209,N_10016);
or U10815 (N_10815,N_10450,N_10431);
nor U10816 (N_10816,N_10149,N_10320);
nand U10817 (N_10817,N_10273,N_10031);
nor U10818 (N_10818,N_10447,N_10395);
nand U10819 (N_10819,N_10185,N_10444);
and U10820 (N_10820,N_10183,N_10269);
xor U10821 (N_10821,N_10214,N_10222);
and U10822 (N_10822,N_10050,N_10314);
nor U10823 (N_10823,N_10084,N_10286);
xnor U10824 (N_10824,N_10175,N_10270);
or U10825 (N_10825,N_10183,N_10094);
and U10826 (N_10826,N_10406,N_10353);
or U10827 (N_10827,N_10022,N_10211);
and U10828 (N_10828,N_10055,N_10222);
and U10829 (N_10829,N_10124,N_10389);
nand U10830 (N_10830,N_10391,N_10340);
or U10831 (N_10831,N_10264,N_10392);
nand U10832 (N_10832,N_10139,N_10389);
xor U10833 (N_10833,N_10179,N_10007);
and U10834 (N_10834,N_10037,N_10467);
or U10835 (N_10835,N_10024,N_10437);
nor U10836 (N_10836,N_10421,N_10071);
nand U10837 (N_10837,N_10459,N_10150);
nand U10838 (N_10838,N_10319,N_10325);
nor U10839 (N_10839,N_10230,N_10124);
nand U10840 (N_10840,N_10413,N_10235);
nand U10841 (N_10841,N_10343,N_10300);
or U10842 (N_10842,N_10383,N_10294);
nor U10843 (N_10843,N_10306,N_10327);
and U10844 (N_10844,N_10020,N_10088);
nand U10845 (N_10845,N_10101,N_10057);
nor U10846 (N_10846,N_10187,N_10106);
or U10847 (N_10847,N_10019,N_10173);
or U10848 (N_10848,N_10045,N_10237);
nor U10849 (N_10849,N_10444,N_10049);
nand U10850 (N_10850,N_10428,N_10161);
and U10851 (N_10851,N_10278,N_10133);
nand U10852 (N_10852,N_10325,N_10205);
nor U10853 (N_10853,N_10381,N_10398);
and U10854 (N_10854,N_10275,N_10114);
nand U10855 (N_10855,N_10487,N_10119);
nand U10856 (N_10856,N_10001,N_10273);
nand U10857 (N_10857,N_10100,N_10002);
nand U10858 (N_10858,N_10133,N_10245);
or U10859 (N_10859,N_10276,N_10188);
or U10860 (N_10860,N_10496,N_10407);
and U10861 (N_10861,N_10279,N_10274);
nor U10862 (N_10862,N_10351,N_10348);
nor U10863 (N_10863,N_10474,N_10123);
nor U10864 (N_10864,N_10269,N_10203);
xor U10865 (N_10865,N_10029,N_10426);
nor U10866 (N_10866,N_10164,N_10314);
and U10867 (N_10867,N_10267,N_10191);
nand U10868 (N_10868,N_10161,N_10358);
or U10869 (N_10869,N_10401,N_10312);
nor U10870 (N_10870,N_10022,N_10200);
and U10871 (N_10871,N_10348,N_10126);
and U10872 (N_10872,N_10205,N_10370);
and U10873 (N_10873,N_10353,N_10039);
xor U10874 (N_10874,N_10126,N_10386);
xnor U10875 (N_10875,N_10342,N_10060);
and U10876 (N_10876,N_10081,N_10446);
nor U10877 (N_10877,N_10330,N_10477);
nor U10878 (N_10878,N_10174,N_10120);
nor U10879 (N_10879,N_10117,N_10395);
nor U10880 (N_10880,N_10241,N_10285);
nand U10881 (N_10881,N_10274,N_10499);
and U10882 (N_10882,N_10192,N_10448);
nor U10883 (N_10883,N_10446,N_10285);
nand U10884 (N_10884,N_10039,N_10212);
nand U10885 (N_10885,N_10127,N_10265);
nor U10886 (N_10886,N_10059,N_10165);
and U10887 (N_10887,N_10179,N_10202);
and U10888 (N_10888,N_10032,N_10345);
xnor U10889 (N_10889,N_10108,N_10460);
nand U10890 (N_10890,N_10322,N_10223);
and U10891 (N_10891,N_10360,N_10359);
and U10892 (N_10892,N_10289,N_10135);
nor U10893 (N_10893,N_10253,N_10455);
nand U10894 (N_10894,N_10417,N_10259);
nand U10895 (N_10895,N_10384,N_10190);
and U10896 (N_10896,N_10116,N_10076);
or U10897 (N_10897,N_10314,N_10398);
xor U10898 (N_10898,N_10189,N_10469);
or U10899 (N_10899,N_10293,N_10284);
xor U10900 (N_10900,N_10180,N_10231);
nand U10901 (N_10901,N_10090,N_10142);
nor U10902 (N_10902,N_10281,N_10439);
xnor U10903 (N_10903,N_10174,N_10166);
nor U10904 (N_10904,N_10319,N_10035);
nand U10905 (N_10905,N_10110,N_10419);
nor U10906 (N_10906,N_10347,N_10106);
xor U10907 (N_10907,N_10016,N_10123);
nor U10908 (N_10908,N_10251,N_10461);
nor U10909 (N_10909,N_10121,N_10226);
nand U10910 (N_10910,N_10263,N_10100);
and U10911 (N_10911,N_10272,N_10014);
or U10912 (N_10912,N_10329,N_10079);
and U10913 (N_10913,N_10434,N_10103);
and U10914 (N_10914,N_10208,N_10490);
xnor U10915 (N_10915,N_10133,N_10430);
and U10916 (N_10916,N_10024,N_10155);
xnor U10917 (N_10917,N_10270,N_10376);
nor U10918 (N_10918,N_10426,N_10499);
or U10919 (N_10919,N_10248,N_10335);
or U10920 (N_10920,N_10258,N_10419);
or U10921 (N_10921,N_10165,N_10457);
or U10922 (N_10922,N_10063,N_10155);
nand U10923 (N_10923,N_10201,N_10157);
and U10924 (N_10924,N_10206,N_10359);
xor U10925 (N_10925,N_10258,N_10310);
or U10926 (N_10926,N_10332,N_10308);
nand U10927 (N_10927,N_10028,N_10057);
and U10928 (N_10928,N_10234,N_10461);
and U10929 (N_10929,N_10478,N_10268);
and U10930 (N_10930,N_10466,N_10236);
and U10931 (N_10931,N_10124,N_10313);
and U10932 (N_10932,N_10263,N_10453);
or U10933 (N_10933,N_10117,N_10193);
nor U10934 (N_10934,N_10167,N_10219);
or U10935 (N_10935,N_10024,N_10398);
and U10936 (N_10936,N_10346,N_10110);
nand U10937 (N_10937,N_10186,N_10188);
nand U10938 (N_10938,N_10084,N_10074);
and U10939 (N_10939,N_10111,N_10249);
xnor U10940 (N_10940,N_10372,N_10485);
nor U10941 (N_10941,N_10284,N_10238);
and U10942 (N_10942,N_10001,N_10253);
xor U10943 (N_10943,N_10458,N_10260);
nand U10944 (N_10944,N_10277,N_10142);
nor U10945 (N_10945,N_10016,N_10096);
and U10946 (N_10946,N_10159,N_10280);
nor U10947 (N_10947,N_10474,N_10492);
nor U10948 (N_10948,N_10445,N_10085);
xnor U10949 (N_10949,N_10084,N_10464);
xor U10950 (N_10950,N_10152,N_10250);
nor U10951 (N_10951,N_10154,N_10413);
nand U10952 (N_10952,N_10357,N_10064);
nand U10953 (N_10953,N_10097,N_10129);
xor U10954 (N_10954,N_10383,N_10454);
or U10955 (N_10955,N_10009,N_10289);
nand U10956 (N_10956,N_10124,N_10180);
xor U10957 (N_10957,N_10361,N_10192);
nand U10958 (N_10958,N_10132,N_10112);
xor U10959 (N_10959,N_10234,N_10417);
nand U10960 (N_10960,N_10243,N_10230);
nand U10961 (N_10961,N_10177,N_10329);
and U10962 (N_10962,N_10492,N_10340);
nand U10963 (N_10963,N_10009,N_10147);
xor U10964 (N_10964,N_10361,N_10240);
nor U10965 (N_10965,N_10114,N_10442);
nand U10966 (N_10966,N_10446,N_10014);
nor U10967 (N_10967,N_10157,N_10240);
xor U10968 (N_10968,N_10182,N_10226);
nor U10969 (N_10969,N_10497,N_10025);
xnor U10970 (N_10970,N_10445,N_10064);
and U10971 (N_10971,N_10319,N_10073);
nand U10972 (N_10972,N_10041,N_10175);
and U10973 (N_10973,N_10151,N_10025);
and U10974 (N_10974,N_10038,N_10083);
and U10975 (N_10975,N_10437,N_10307);
and U10976 (N_10976,N_10140,N_10202);
and U10977 (N_10977,N_10415,N_10090);
or U10978 (N_10978,N_10143,N_10427);
nor U10979 (N_10979,N_10342,N_10010);
nand U10980 (N_10980,N_10480,N_10470);
and U10981 (N_10981,N_10371,N_10302);
or U10982 (N_10982,N_10405,N_10036);
xnor U10983 (N_10983,N_10094,N_10435);
nand U10984 (N_10984,N_10234,N_10146);
nand U10985 (N_10985,N_10339,N_10386);
nor U10986 (N_10986,N_10129,N_10316);
or U10987 (N_10987,N_10310,N_10245);
or U10988 (N_10988,N_10486,N_10407);
and U10989 (N_10989,N_10353,N_10397);
nor U10990 (N_10990,N_10025,N_10471);
and U10991 (N_10991,N_10016,N_10119);
nand U10992 (N_10992,N_10462,N_10252);
and U10993 (N_10993,N_10492,N_10158);
nand U10994 (N_10994,N_10490,N_10084);
nand U10995 (N_10995,N_10427,N_10240);
xnor U10996 (N_10996,N_10126,N_10118);
and U10997 (N_10997,N_10223,N_10018);
xor U10998 (N_10998,N_10145,N_10149);
nand U10999 (N_10999,N_10303,N_10391);
or U11000 (N_11000,N_10880,N_10999);
or U11001 (N_11001,N_10734,N_10700);
nand U11002 (N_11002,N_10678,N_10799);
and U11003 (N_11003,N_10570,N_10770);
nor U11004 (N_11004,N_10783,N_10583);
nor U11005 (N_11005,N_10832,N_10865);
or U11006 (N_11006,N_10981,N_10983);
nor U11007 (N_11007,N_10871,N_10636);
nor U11008 (N_11008,N_10898,N_10905);
nand U11009 (N_11009,N_10691,N_10584);
or U11010 (N_11010,N_10607,N_10712);
xnor U11011 (N_11011,N_10746,N_10568);
and U11012 (N_11012,N_10856,N_10842);
xnor U11013 (N_11013,N_10903,N_10904);
or U11014 (N_11014,N_10502,N_10657);
xnor U11015 (N_11015,N_10915,N_10768);
and U11016 (N_11016,N_10971,N_10989);
xor U11017 (N_11017,N_10776,N_10914);
xor U11018 (N_11018,N_10763,N_10752);
nor U11019 (N_11019,N_10585,N_10806);
xnor U11020 (N_11020,N_10870,N_10567);
nand U11021 (N_11021,N_10522,N_10658);
nand U11022 (N_11022,N_10702,N_10716);
and U11023 (N_11023,N_10955,N_10759);
nand U11024 (N_11024,N_10860,N_10850);
nor U11025 (N_11025,N_10608,N_10721);
xor U11026 (N_11026,N_10647,N_10614);
nor U11027 (N_11027,N_10782,N_10911);
or U11028 (N_11028,N_10674,N_10679);
and U11029 (N_11029,N_10505,N_10848);
nand U11030 (N_11030,N_10566,N_10830);
and U11031 (N_11031,N_10857,N_10698);
nand U11032 (N_11032,N_10808,N_10589);
xor U11033 (N_11033,N_10573,N_10652);
xnor U11034 (N_11034,N_10977,N_10535);
nor U11035 (N_11035,N_10798,N_10660);
or U11036 (N_11036,N_10533,N_10801);
xnor U11037 (N_11037,N_10662,N_10601);
or U11038 (N_11038,N_10552,N_10580);
or U11039 (N_11039,N_10667,N_10627);
xnor U11040 (N_11040,N_10844,N_10953);
and U11041 (N_11041,N_10938,N_10664);
or U11042 (N_11042,N_10772,N_10612);
and U11043 (N_11043,N_10827,N_10883);
nor U11044 (N_11044,N_10939,N_10531);
nand U11045 (N_11045,N_10536,N_10990);
or U11046 (N_11046,N_10895,N_10790);
nor U11047 (N_11047,N_10908,N_10996);
and U11048 (N_11048,N_10766,N_10569);
nor U11049 (N_11049,N_10820,N_10896);
nor U11050 (N_11050,N_10900,N_10738);
nor U11051 (N_11051,N_10773,N_10602);
or U11052 (N_11052,N_10845,N_10872);
or U11053 (N_11053,N_10594,N_10866);
nand U11054 (N_11054,N_10688,N_10651);
nand U11055 (N_11055,N_10694,N_10854);
nand U11056 (N_11056,N_10600,N_10864);
nor U11057 (N_11057,N_10980,N_10737);
or U11058 (N_11058,N_10878,N_10730);
nand U11059 (N_11059,N_10736,N_10598);
or U11060 (N_11060,N_10982,N_10809);
or U11061 (N_11061,N_10745,N_10912);
nand U11062 (N_11062,N_10910,N_10917);
nand U11063 (N_11063,N_10648,N_10606);
nor U11064 (N_11064,N_10693,N_10978);
nand U11065 (N_11065,N_10574,N_10692);
and U11066 (N_11066,N_10720,N_10788);
or U11067 (N_11067,N_10909,N_10689);
xnor U11068 (N_11068,N_10932,N_10529);
or U11069 (N_11069,N_10735,N_10774);
or U11070 (N_11070,N_10951,N_10840);
xnor U11071 (N_11071,N_10604,N_10890);
nor U11072 (N_11072,N_10637,N_10513);
or U11073 (N_11073,N_10644,N_10524);
or U11074 (N_11074,N_10538,N_10653);
and U11075 (N_11075,N_10560,N_10673);
or U11076 (N_11076,N_10676,N_10668);
and U11077 (N_11077,N_10632,N_10944);
and U11078 (N_11078,N_10791,N_10672);
and U11079 (N_11079,N_10509,N_10595);
or U11080 (N_11080,N_10754,N_10544);
xor U11081 (N_11081,N_10706,N_10597);
and U11082 (N_11082,N_10765,N_10994);
or U11083 (N_11083,N_10695,N_10764);
nor U11084 (N_11084,N_10555,N_10512);
and U11085 (N_11085,N_10748,N_10590);
nor U11086 (N_11086,N_10891,N_10897);
and U11087 (N_11087,N_10811,N_10749);
nor U11088 (N_11088,N_10943,N_10501);
nand U11089 (N_11089,N_10525,N_10936);
xnor U11090 (N_11090,N_10515,N_10686);
nor U11091 (N_11091,N_10579,N_10665);
and U11092 (N_11092,N_10642,N_10817);
or U11093 (N_11093,N_10941,N_10521);
nor U11094 (N_11094,N_10704,N_10993);
nand U11095 (N_11095,N_10863,N_10714);
nand U11096 (N_11096,N_10725,N_10804);
or U11097 (N_11097,N_10611,N_10847);
and U11098 (N_11098,N_10805,N_10922);
and U11099 (N_11099,N_10519,N_10859);
xor U11100 (N_11100,N_10596,N_10862);
nor U11101 (N_11101,N_10718,N_10901);
nor U11102 (N_11102,N_10687,N_10528);
and U11103 (N_11103,N_10879,N_10532);
xnor U11104 (N_11104,N_10875,N_10794);
and U11105 (N_11105,N_10979,N_10719);
or U11106 (N_11106,N_10797,N_10884);
nand U11107 (N_11107,N_10551,N_10699);
and U11108 (N_11108,N_10629,N_10630);
nand U11109 (N_11109,N_10813,N_10886);
and U11110 (N_11110,N_10684,N_10670);
and U11111 (N_11111,N_10591,N_10581);
nand U11112 (N_11112,N_10708,N_10825);
nor U11113 (N_11113,N_10504,N_10920);
xor U11114 (N_11114,N_10923,N_10998);
nor U11115 (N_11115,N_10666,N_10887);
nand U11116 (N_11116,N_10743,N_10619);
or U11117 (N_11117,N_10609,N_10624);
xnor U11118 (N_11118,N_10617,N_10625);
or U11119 (N_11119,N_10534,N_10545);
and U11120 (N_11120,N_10973,N_10728);
or U11121 (N_11121,N_10899,N_10960);
or U11122 (N_11122,N_10937,N_10655);
xor U11123 (N_11123,N_10778,N_10711);
nand U11124 (N_11124,N_10829,N_10739);
xor U11125 (N_11125,N_10959,N_10967);
nand U11126 (N_11126,N_10918,N_10924);
and U11127 (N_11127,N_10577,N_10751);
or U11128 (N_11128,N_10514,N_10946);
and U11129 (N_11129,N_10709,N_10603);
xor U11130 (N_11130,N_10965,N_10760);
xor U11131 (N_11131,N_10777,N_10775);
or U11132 (N_11132,N_10869,N_10784);
and U11133 (N_11133,N_10926,N_10838);
or U11134 (N_11134,N_10893,N_10613);
or U11135 (N_11135,N_10565,N_10543);
xnor U11136 (N_11136,N_10582,N_10523);
or U11137 (N_11137,N_10940,N_10962);
and U11138 (N_11138,N_10843,N_10701);
nor U11139 (N_11139,N_10762,N_10690);
xor U11140 (N_11140,N_10852,N_10826);
or U11141 (N_11141,N_10818,N_10952);
or U11142 (N_11142,N_10628,N_10623);
or U11143 (N_11143,N_10508,N_10753);
nand U11144 (N_11144,N_10800,N_10575);
xor U11145 (N_11145,N_10507,N_10785);
xor U11146 (N_11146,N_10705,N_10835);
xnor U11147 (N_11147,N_10605,N_10795);
nor U11148 (N_11148,N_10968,N_10781);
and U11149 (N_11149,N_10554,N_10511);
xnor U11150 (N_11150,N_10592,N_10550);
or U11151 (N_11151,N_10894,N_10779);
and U11152 (N_11152,N_10916,N_10927);
nor U11153 (N_11153,N_10517,N_10995);
xor U11154 (N_11154,N_10954,N_10834);
nand U11155 (N_11155,N_10931,N_10950);
or U11156 (N_11156,N_10787,N_10729);
nand U11157 (N_11157,N_10621,N_10685);
nor U11158 (N_11158,N_10558,N_10855);
or U11159 (N_11159,N_10867,N_10518);
or U11160 (N_11160,N_10726,N_10564);
and U11161 (N_11161,N_10537,N_10933);
and U11162 (N_11162,N_10727,N_10970);
nor U11163 (N_11163,N_10618,N_10682);
xor U11164 (N_11164,N_10925,N_10683);
and U11165 (N_11165,N_10733,N_10821);
or U11166 (N_11166,N_10542,N_10526);
xnor U11167 (N_11167,N_10930,N_10945);
and U11168 (N_11168,N_10530,N_10576);
or U11169 (N_11169,N_10731,N_10771);
and U11170 (N_11170,N_10547,N_10541);
or U11171 (N_11171,N_10957,N_10812);
and U11172 (N_11172,N_10755,N_10640);
xor U11173 (N_11173,N_10643,N_10814);
xor U11174 (N_11174,N_10974,N_10680);
xor U11175 (N_11175,N_10969,N_10626);
or U11176 (N_11176,N_10562,N_10822);
nand U11177 (N_11177,N_10988,N_10928);
or U11178 (N_11178,N_10885,N_10756);
nor U11179 (N_11179,N_10747,N_10540);
nor U11180 (N_11180,N_10559,N_10861);
nor U11181 (N_11181,N_10921,N_10561);
nand U11182 (N_11182,N_10527,N_10549);
or U11183 (N_11183,N_10586,N_10713);
xor U11184 (N_11184,N_10539,N_10656);
nand U11185 (N_11185,N_10992,N_10669);
nand U11186 (N_11186,N_10557,N_10744);
nand U11187 (N_11187,N_10837,N_10520);
and U11188 (N_11188,N_10947,N_10659);
and U11189 (N_11189,N_10750,N_10675);
xor U11190 (N_11190,N_10997,N_10757);
xnor U11191 (N_11191,N_10638,N_10697);
and U11192 (N_11192,N_10723,N_10984);
nor U11193 (N_11193,N_10503,N_10906);
or U11194 (N_11194,N_10563,N_10789);
nor U11195 (N_11195,N_10696,N_10615);
xnor U11196 (N_11196,N_10722,N_10635);
nand U11197 (N_11197,N_10741,N_10645);
nand U11198 (N_11198,N_10786,N_10961);
and U11199 (N_11199,N_10792,N_10831);
nand U11200 (N_11200,N_10677,N_10929);
and U11201 (N_11201,N_10853,N_10976);
nand U11202 (N_11202,N_10966,N_10681);
nand U11203 (N_11203,N_10841,N_10949);
nand U11204 (N_11204,N_10717,N_10654);
and U11205 (N_11205,N_10810,N_10987);
or U11206 (N_11206,N_10815,N_10913);
or U11207 (N_11207,N_10849,N_10631);
and U11208 (N_11208,N_10803,N_10616);
or U11209 (N_11209,N_10761,N_10858);
xnor U11210 (N_11210,N_10587,N_10593);
nand U11211 (N_11211,N_10874,N_10942);
nor U11212 (N_11212,N_10548,N_10572);
nor U11213 (N_11213,N_10546,N_10715);
nor U11214 (N_11214,N_10902,N_10724);
nand U11215 (N_11215,N_10599,N_10740);
or U11216 (N_11216,N_10622,N_10868);
nor U11217 (N_11217,N_10500,N_10892);
xor U11218 (N_11218,N_10510,N_10671);
or U11219 (N_11219,N_10963,N_10649);
nor U11220 (N_11220,N_10758,N_10663);
and U11221 (N_11221,N_10889,N_10641);
nor U11222 (N_11222,N_10578,N_10661);
and U11223 (N_11223,N_10846,N_10991);
nand U11224 (N_11224,N_10707,N_10972);
or U11225 (N_11225,N_10948,N_10639);
xnor U11226 (N_11226,N_10793,N_10710);
nand U11227 (N_11227,N_10934,N_10556);
nor U11228 (N_11228,N_10802,N_10824);
or U11229 (N_11229,N_10881,N_10633);
or U11230 (N_11230,N_10732,N_10882);
nand U11231 (N_11231,N_10819,N_10767);
and U11232 (N_11232,N_10634,N_10769);
nand U11233 (N_11233,N_10836,N_10610);
nor U11234 (N_11234,N_10985,N_10620);
xnor U11235 (N_11235,N_10851,N_10919);
nand U11236 (N_11236,N_10877,N_10935);
or U11237 (N_11237,N_10964,N_10956);
nor U11238 (N_11238,N_10888,N_10828);
nand U11239 (N_11239,N_10516,N_10839);
or U11240 (N_11240,N_10907,N_10571);
nand U11241 (N_11241,N_10876,N_10650);
nand U11242 (N_11242,N_10975,N_10742);
nand U11243 (N_11243,N_10796,N_10816);
xnor U11244 (N_11244,N_10986,N_10506);
and U11245 (N_11245,N_10833,N_10780);
xor U11246 (N_11246,N_10958,N_10823);
and U11247 (N_11247,N_10646,N_10873);
xnor U11248 (N_11248,N_10703,N_10588);
xnor U11249 (N_11249,N_10553,N_10807);
nor U11250 (N_11250,N_10730,N_10629);
xnor U11251 (N_11251,N_10811,N_10807);
xor U11252 (N_11252,N_10925,N_10644);
and U11253 (N_11253,N_10891,N_10577);
and U11254 (N_11254,N_10734,N_10586);
nand U11255 (N_11255,N_10625,N_10811);
or U11256 (N_11256,N_10599,N_10679);
nor U11257 (N_11257,N_10798,N_10709);
or U11258 (N_11258,N_10900,N_10699);
xor U11259 (N_11259,N_10979,N_10565);
nor U11260 (N_11260,N_10647,N_10795);
and U11261 (N_11261,N_10918,N_10585);
or U11262 (N_11262,N_10538,N_10682);
or U11263 (N_11263,N_10662,N_10658);
and U11264 (N_11264,N_10509,N_10519);
nand U11265 (N_11265,N_10533,N_10655);
or U11266 (N_11266,N_10778,N_10751);
nor U11267 (N_11267,N_10927,N_10779);
and U11268 (N_11268,N_10724,N_10590);
xor U11269 (N_11269,N_10576,N_10910);
and U11270 (N_11270,N_10733,N_10514);
xnor U11271 (N_11271,N_10985,N_10561);
nor U11272 (N_11272,N_10686,N_10681);
or U11273 (N_11273,N_10816,N_10763);
and U11274 (N_11274,N_10948,N_10935);
or U11275 (N_11275,N_10716,N_10582);
nor U11276 (N_11276,N_10905,N_10902);
nor U11277 (N_11277,N_10797,N_10964);
or U11278 (N_11278,N_10678,N_10945);
nor U11279 (N_11279,N_10821,N_10909);
nand U11280 (N_11280,N_10795,N_10666);
xnor U11281 (N_11281,N_10937,N_10611);
or U11282 (N_11282,N_10996,N_10951);
or U11283 (N_11283,N_10955,N_10666);
nor U11284 (N_11284,N_10657,N_10824);
nor U11285 (N_11285,N_10969,N_10756);
or U11286 (N_11286,N_10757,N_10790);
or U11287 (N_11287,N_10964,N_10795);
nand U11288 (N_11288,N_10553,N_10950);
nand U11289 (N_11289,N_10839,N_10845);
xnor U11290 (N_11290,N_10915,N_10921);
xnor U11291 (N_11291,N_10843,N_10691);
nor U11292 (N_11292,N_10669,N_10689);
and U11293 (N_11293,N_10789,N_10769);
or U11294 (N_11294,N_10587,N_10542);
xor U11295 (N_11295,N_10829,N_10636);
or U11296 (N_11296,N_10968,N_10586);
or U11297 (N_11297,N_10644,N_10906);
nand U11298 (N_11298,N_10592,N_10969);
xnor U11299 (N_11299,N_10623,N_10662);
or U11300 (N_11300,N_10806,N_10660);
nor U11301 (N_11301,N_10900,N_10988);
or U11302 (N_11302,N_10574,N_10547);
nor U11303 (N_11303,N_10814,N_10521);
or U11304 (N_11304,N_10850,N_10641);
nor U11305 (N_11305,N_10818,N_10740);
nand U11306 (N_11306,N_10587,N_10533);
nand U11307 (N_11307,N_10692,N_10771);
nor U11308 (N_11308,N_10503,N_10600);
and U11309 (N_11309,N_10798,N_10922);
or U11310 (N_11310,N_10670,N_10708);
xnor U11311 (N_11311,N_10703,N_10724);
nor U11312 (N_11312,N_10840,N_10809);
or U11313 (N_11313,N_10638,N_10701);
nor U11314 (N_11314,N_10564,N_10762);
or U11315 (N_11315,N_10729,N_10604);
nor U11316 (N_11316,N_10712,N_10770);
or U11317 (N_11317,N_10909,N_10975);
nand U11318 (N_11318,N_10972,N_10750);
nand U11319 (N_11319,N_10816,N_10636);
nor U11320 (N_11320,N_10602,N_10870);
nand U11321 (N_11321,N_10594,N_10582);
and U11322 (N_11322,N_10726,N_10779);
nor U11323 (N_11323,N_10624,N_10634);
nand U11324 (N_11324,N_10533,N_10609);
nor U11325 (N_11325,N_10974,N_10552);
xnor U11326 (N_11326,N_10917,N_10744);
xor U11327 (N_11327,N_10681,N_10573);
and U11328 (N_11328,N_10580,N_10557);
or U11329 (N_11329,N_10502,N_10970);
or U11330 (N_11330,N_10747,N_10526);
and U11331 (N_11331,N_10673,N_10882);
nor U11332 (N_11332,N_10817,N_10605);
or U11333 (N_11333,N_10594,N_10558);
nor U11334 (N_11334,N_10503,N_10642);
nand U11335 (N_11335,N_10691,N_10786);
and U11336 (N_11336,N_10752,N_10813);
nor U11337 (N_11337,N_10707,N_10955);
and U11338 (N_11338,N_10970,N_10572);
nand U11339 (N_11339,N_10502,N_10685);
nand U11340 (N_11340,N_10657,N_10625);
nor U11341 (N_11341,N_10734,N_10659);
nor U11342 (N_11342,N_10944,N_10747);
or U11343 (N_11343,N_10896,N_10985);
or U11344 (N_11344,N_10994,N_10559);
xor U11345 (N_11345,N_10933,N_10528);
and U11346 (N_11346,N_10791,N_10683);
nor U11347 (N_11347,N_10820,N_10659);
or U11348 (N_11348,N_10876,N_10610);
nor U11349 (N_11349,N_10962,N_10774);
or U11350 (N_11350,N_10925,N_10785);
nor U11351 (N_11351,N_10645,N_10808);
nand U11352 (N_11352,N_10672,N_10663);
nand U11353 (N_11353,N_10722,N_10757);
nand U11354 (N_11354,N_10889,N_10668);
nand U11355 (N_11355,N_10766,N_10956);
and U11356 (N_11356,N_10582,N_10767);
nor U11357 (N_11357,N_10681,N_10524);
nand U11358 (N_11358,N_10542,N_10878);
nand U11359 (N_11359,N_10695,N_10974);
or U11360 (N_11360,N_10950,N_10581);
and U11361 (N_11361,N_10886,N_10849);
xor U11362 (N_11362,N_10689,N_10922);
nor U11363 (N_11363,N_10505,N_10908);
nor U11364 (N_11364,N_10675,N_10500);
or U11365 (N_11365,N_10834,N_10889);
and U11366 (N_11366,N_10981,N_10562);
xor U11367 (N_11367,N_10789,N_10718);
and U11368 (N_11368,N_10714,N_10532);
nand U11369 (N_11369,N_10984,N_10761);
nand U11370 (N_11370,N_10740,N_10951);
or U11371 (N_11371,N_10627,N_10591);
nand U11372 (N_11372,N_10660,N_10630);
nor U11373 (N_11373,N_10618,N_10593);
and U11374 (N_11374,N_10967,N_10809);
or U11375 (N_11375,N_10908,N_10714);
nand U11376 (N_11376,N_10900,N_10844);
or U11377 (N_11377,N_10649,N_10555);
nor U11378 (N_11378,N_10613,N_10756);
nand U11379 (N_11379,N_10696,N_10778);
nand U11380 (N_11380,N_10621,N_10512);
nand U11381 (N_11381,N_10825,N_10999);
nor U11382 (N_11382,N_10677,N_10913);
nor U11383 (N_11383,N_10839,N_10530);
nand U11384 (N_11384,N_10746,N_10645);
nor U11385 (N_11385,N_10548,N_10957);
or U11386 (N_11386,N_10971,N_10939);
or U11387 (N_11387,N_10627,N_10559);
or U11388 (N_11388,N_10682,N_10849);
or U11389 (N_11389,N_10900,N_10962);
nand U11390 (N_11390,N_10710,N_10808);
xnor U11391 (N_11391,N_10963,N_10721);
nor U11392 (N_11392,N_10727,N_10521);
and U11393 (N_11393,N_10986,N_10900);
nor U11394 (N_11394,N_10688,N_10757);
xnor U11395 (N_11395,N_10603,N_10526);
or U11396 (N_11396,N_10912,N_10815);
nand U11397 (N_11397,N_10660,N_10780);
or U11398 (N_11398,N_10942,N_10783);
xnor U11399 (N_11399,N_10666,N_10629);
xor U11400 (N_11400,N_10639,N_10708);
and U11401 (N_11401,N_10690,N_10984);
or U11402 (N_11402,N_10981,N_10504);
xnor U11403 (N_11403,N_10948,N_10730);
and U11404 (N_11404,N_10786,N_10799);
nor U11405 (N_11405,N_10728,N_10938);
nor U11406 (N_11406,N_10560,N_10817);
xor U11407 (N_11407,N_10842,N_10927);
nand U11408 (N_11408,N_10753,N_10965);
or U11409 (N_11409,N_10654,N_10634);
xor U11410 (N_11410,N_10510,N_10685);
xor U11411 (N_11411,N_10764,N_10893);
nand U11412 (N_11412,N_10555,N_10549);
xor U11413 (N_11413,N_10795,N_10517);
nor U11414 (N_11414,N_10974,N_10532);
or U11415 (N_11415,N_10605,N_10661);
nor U11416 (N_11416,N_10608,N_10904);
nand U11417 (N_11417,N_10525,N_10806);
and U11418 (N_11418,N_10795,N_10669);
xnor U11419 (N_11419,N_10843,N_10942);
and U11420 (N_11420,N_10902,N_10975);
xnor U11421 (N_11421,N_10953,N_10642);
or U11422 (N_11422,N_10793,N_10997);
or U11423 (N_11423,N_10935,N_10743);
nand U11424 (N_11424,N_10915,N_10700);
nor U11425 (N_11425,N_10804,N_10510);
xor U11426 (N_11426,N_10892,N_10617);
nor U11427 (N_11427,N_10716,N_10913);
and U11428 (N_11428,N_10683,N_10916);
and U11429 (N_11429,N_10880,N_10849);
nand U11430 (N_11430,N_10601,N_10667);
nand U11431 (N_11431,N_10918,N_10954);
xor U11432 (N_11432,N_10960,N_10511);
nand U11433 (N_11433,N_10770,N_10505);
and U11434 (N_11434,N_10605,N_10984);
xor U11435 (N_11435,N_10852,N_10748);
or U11436 (N_11436,N_10840,N_10705);
and U11437 (N_11437,N_10920,N_10676);
or U11438 (N_11438,N_10542,N_10862);
and U11439 (N_11439,N_10658,N_10653);
and U11440 (N_11440,N_10607,N_10514);
xor U11441 (N_11441,N_10990,N_10525);
nand U11442 (N_11442,N_10517,N_10954);
and U11443 (N_11443,N_10500,N_10737);
xnor U11444 (N_11444,N_10885,N_10763);
nor U11445 (N_11445,N_10898,N_10996);
nor U11446 (N_11446,N_10555,N_10899);
or U11447 (N_11447,N_10841,N_10631);
or U11448 (N_11448,N_10682,N_10704);
xnor U11449 (N_11449,N_10501,N_10892);
nand U11450 (N_11450,N_10883,N_10938);
and U11451 (N_11451,N_10594,N_10949);
and U11452 (N_11452,N_10534,N_10550);
and U11453 (N_11453,N_10758,N_10806);
and U11454 (N_11454,N_10699,N_10710);
or U11455 (N_11455,N_10539,N_10970);
or U11456 (N_11456,N_10579,N_10843);
xor U11457 (N_11457,N_10888,N_10623);
nor U11458 (N_11458,N_10578,N_10931);
or U11459 (N_11459,N_10694,N_10514);
or U11460 (N_11460,N_10705,N_10587);
nand U11461 (N_11461,N_10715,N_10891);
nor U11462 (N_11462,N_10643,N_10927);
nor U11463 (N_11463,N_10820,N_10537);
and U11464 (N_11464,N_10839,N_10736);
and U11465 (N_11465,N_10957,N_10847);
xor U11466 (N_11466,N_10888,N_10599);
or U11467 (N_11467,N_10517,N_10550);
and U11468 (N_11468,N_10857,N_10599);
xnor U11469 (N_11469,N_10963,N_10748);
nand U11470 (N_11470,N_10992,N_10944);
or U11471 (N_11471,N_10564,N_10739);
nor U11472 (N_11472,N_10827,N_10661);
xnor U11473 (N_11473,N_10663,N_10838);
xnor U11474 (N_11474,N_10580,N_10756);
nor U11475 (N_11475,N_10554,N_10707);
nor U11476 (N_11476,N_10517,N_10684);
and U11477 (N_11477,N_10973,N_10925);
xnor U11478 (N_11478,N_10793,N_10597);
nand U11479 (N_11479,N_10735,N_10530);
and U11480 (N_11480,N_10705,N_10871);
nor U11481 (N_11481,N_10743,N_10844);
nor U11482 (N_11482,N_10948,N_10890);
xor U11483 (N_11483,N_10947,N_10653);
or U11484 (N_11484,N_10663,N_10993);
nand U11485 (N_11485,N_10560,N_10718);
or U11486 (N_11486,N_10638,N_10581);
and U11487 (N_11487,N_10809,N_10643);
or U11488 (N_11488,N_10968,N_10770);
nand U11489 (N_11489,N_10977,N_10544);
nand U11490 (N_11490,N_10837,N_10890);
nand U11491 (N_11491,N_10706,N_10975);
or U11492 (N_11492,N_10982,N_10907);
nor U11493 (N_11493,N_10899,N_10888);
xor U11494 (N_11494,N_10681,N_10551);
nand U11495 (N_11495,N_10637,N_10526);
nor U11496 (N_11496,N_10556,N_10940);
nand U11497 (N_11497,N_10559,N_10560);
and U11498 (N_11498,N_10536,N_10714);
xor U11499 (N_11499,N_10969,N_10958);
or U11500 (N_11500,N_11057,N_11099);
and U11501 (N_11501,N_11480,N_11268);
xor U11502 (N_11502,N_11018,N_11237);
xnor U11503 (N_11503,N_11136,N_11132);
or U11504 (N_11504,N_11294,N_11088);
or U11505 (N_11505,N_11329,N_11409);
xnor U11506 (N_11506,N_11179,N_11241);
nor U11507 (N_11507,N_11193,N_11277);
nor U11508 (N_11508,N_11116,N_11246);
and U11509 (N_11509,N_11448,N_11081);
nor U11510 (N_11510,N_11162,N_11374);
xor U11511 (N_11511,N_11417,N_11146);
or U11512 (N_11512,N_11168,N_11157);
xnor U11513 (N_11513,N_11189,N_11263);
xnor U11514 (N_11514,N_11231,N_11342);
and U11515 (N_11515,N_11164,N_11210);
nand U11516 (N_11516,N_11289,N_11302);
nor U11517 (N_11517,N_11100,N_11346);
and U11518 (N_11518,N_11258,N_11188);
or U11519 (N_11519,N_11438,N_11256);
nor U11520 (N_11520,N_11488,N_11058);
and U11521 (N_11521,N_11083,N_11320);
or U11522 (N_11522,N_11222,N_11357);
xnor U11523 (N_11523,N_11013,N_11330);
nor U11524 (N_11524,N_11327,N_11355);
and U11525 (N_11525,N_11412,N_11197);
and U11526 (N_11526,N_11159,N_11254);
and U11527 (N_11527,N_11235,N_11475);
nand U11528 (N_11528,N_11025,N_11219);
nor U11529 (N_11529,N_11447,N_11174);
nor U11530 (N_11530,N_11322,N_11353);
xnor U11531 (N_11531,N_11075,N_11005);
nor U11532 (N_11532,N_11082,N_11175);
nor U11533 (N_11533,N_11416,N_11308);
xor U11534 (N_11534,N_11388,N_11170);
or U11535 (N_11535,N_11269,N_11207);
or U11536 (N_11536,N_11242,N_11031);
xnor U11537 (N_11537,N_11128,N_11483);
nor U11538 (N_11538,N_11473,N_11095);
xor U11539 (N_11539,N_11017,N_11395);
nand U11540 (N_11540,N_11087,N_11065);
or U11541 (N_11541,N_11153,N_11354);
nand U11542 (N_11542,N_11348,N_11117);
nand U11543 (N_11543,N_11295,N_11339);
nor U11544 (N_11544,N_11150,N_11171);
xor U11545 (N_11545,N_11421,N_11201);
nand U11546 (N_11546,N_11465,N_11366);
nand U11547 (N_11547,N_11215,N_11037);
or U11548 (N_11548,N_11212,N_11143);
xnor U11549 (N_11549,N_11273,N_11103);
nor U11550 (N_11550,N_11209,N_11107);
and U11551 (N_11551,N_11042,N_11108);
or U11552 (N_11552,N_11078,N_11109);
and U11553 (N_11553,N_11454,N_11457);
nand U11554 (N_11554,N_11259,N_11461);
nand U11555 (N_11555,N_11009,N_11120);
or U11556 (N_11556,N_11424,N_11093);
and U11557 (N_11557,N_11455,N_11048);
and U11558 (N_11558,N_11185,N_11314);
and U11559 (N_11559,N_11040,N_11034);
nand U11560 (N_11560,N_11003,N_11267);
and U11561 (N_11561,N_11344,N_11002);
nor U11562 (N_11562,N_11247,N_11436);
xor U11563 (N_11563,N_11152,N_11063);
xnor U11564 (N_11564,N_11446,N_11300);
or U11565 (N_11565,N_11274,N_11482);
and U11566 (N_11566,N_11049,N_11485);
nor U11567 (N_11567,N_11379,N_11323);
or U11568 (N_11568,N_11262,N_11264);
or U11569 (N_11569,N_11377,N_11499);
xor U11570 (N_11570,N_11122,N_11383);
or U11571 (N_11571,N_11324,N_11196);
or U11572 (N_11572,N_11008,N_11206);
xnor U11573 (N_11573,N_11123,N_11358);
xnor U11574 (N_11574,N_11054,N_11004);
nand U11575 (N_11575,N_11481,N_11279);
nor U11576 (N_11576,N_11035,N_11144);
and U11577 (N_11577,N_11290,N_11378);
and U11578 (N_11578,N_11403,N_11453);
and U11579 (N_11579,N_11331,N_11486);
nand U11580 (N_11580,N_11376,N_11177);
and U11581 (N_11581,N_11211,N_11158);
nor U11582 (N_11582,N_11167,N_11362);
nand U11583 (N_11583,N_11444,N_11394);
nand U11584 (N_11584,N_11350,N_11372);
or U11585 (N_11585,N_11073,N_11024);
and U11586 (N_11586,N_11156,N_11045);
nand U11587 (N_11587,N_11317,N_11006);
and U11588 (N_11588,N_11126,N_11079);
xor U11589 (N_11589,N_11076,N_11370);
and U11590 (N_11590,N_11187,N_11284);
and U11591 (N_11591,N_11134,N_11133);
or U11592 (N_11592,N_11112,N_11288);
or U11593 (N_11593,N_11142,N_11272);
or U11594 (N_11594,N_11026,N_11229);
nand U11595 (N_11595,N_11479,N_11463);
nand U11596 (N_11596,N_11343,N_11494);
nand U11597 (N_11597,N_11135,N_11102);
nor U11598 (N_11598,N_11028,N_11077);
nor U11599 (N_11599,N_11449,N_11255);
or U11600 (N_11600,N_11292,N_11176);
and U11601 (N_11601,N_11000,N_11181);
xnor U11602 (N_11602,N_11094,N_11293);
nor U11603 (N_11603,N_11437,N_11022);
nand U11604 (N_11604,N_11154,N_11385);
nand U11605 (N_11605,N_11228,N_11326);
xnor U11606 (N_11606,N_11356,N_11335);
or U11607 (N_11607,N_11307,N_11425);
nand U11608 (N_11608,N_11271,N_11418);
and U11609 (N_11609,N_11487,N_11275);
or U11610 (N_11610,N_11129,N_11405);
nand U11611 (N_11611,N_11234,N_11309);
xor U11612 (N_11612,N_11172,N_11408);
nand U11613 (N_11613,N_11404,N_11224);
and U11614 (N_11614,N_11382,N_11423);
xnor U11615 (N_11615,N_11462,N_11451);
nand U11616 (N_11616,N_11019,N_11352);
nor U11617 (N_11617,N_11299,N_11336);
nor U11618 (N_11618,N_11380,N_11249);
xor U11619 (N_11619,N_11396,N_11141);
xor U11620 (N_11620,N_11315,N_11384);
or U11621 (N_11621,N_11127,N_11029);
nor U11622 (N_11622,N_11422,N_11431);
nand U11623 (N_11623,N_11051,N_11226);
and U11624 (N_11624,N_11092,N_11021);
or U11625 (N_11625,N_11166,N_11464);
xnor U11626 (N_11626,N_11411,N_11347);
nand U11627 (N_11627,N_11470,N_11068);
xnor U11628 (N_11628,N_11435,N_11469);
nand U11629 (N_11629,N_11182,N_11399);
nor U11630 (N_11630,N_11496,N_11137);
nor U11631 (N_11631,N_11270,N_11276);
nand U11632 (N_11632,N_11280,N_11038);
nor U11633 (N_11633,N_11478,N_11476);
or U11634 (N_11634,N_11253,N_11227);
nand U11635 (N_11635,N_11204,N_11086);
and U11636 (N_11636,N_11043,N_11311);
xor U11637 (N_11637,N_11221,N_11105);
nor U11638 (N_11638,N_11340,N_11066);
nor U11639 (N_11639,N_11287,N_11367);
nand U11640 (N_11640,N_11124,N_11349);
nor U11641 (N_11641,N_11248,N_11080);
nor U11642 (N_11642,N_11419,N_11061);
xor U11643 (N_11643,N_11191,N_11318);
nor U11644 (N_11644,N_11303,N_11363);
xnor U11645 (N_11645,N_11130,N_11452);
nor U11646 (N_11646,N_11381,N_11345);
and U11647 (N_11647,N_11319,N_11433);
or U11648 (N_11648,N_11398,N_11218);
and U11649 (N_11649,N_11055,N_11460);
nand U11650 (N_11650,N_11466,N_11337);
or U11651 (N_11651,N_11285,N_11244);
and U11652 (N_11652,N_11429,N_11402);
and U11653 (N_11653,N_11427,N_11430);
xor U11654 (N_11654,N_11239,N_11202);
nor U11655 (N_11655,N_11012,N_11371);
nor U11656 (N_11656,N_11217,N_11261);
xnor U11657 (N_11657,N_11401,N_11139);
nor U11658 (N_11658,N_11467,N_11203);
nor U11659 (N_11659,N_11145,N_11312);
xor U11660 (N_11660,N_11151,N_11072);
or U11661 (N_11661,N_11016,N_11140);
xor U11662 (N_11662,N_11369,N_11493);
or U11663 (N_11663,N_11328,N_11097);
or U11664 (N_11664,N_11434,N_11291);
or U11665 (N_11665,N_11148,N_11165);
nor U11666 (N_11666,N_11147,N_11495);
nand U11667 (N_11667,N_11050,N_11230);
xnor U11668 (N_11668,N_11007,N_11039);
and U11669 (N_11669,N_11085,N_11014);
nor U11670 (N_11670,N_11064,N_11118);
or U11671 (N_11671,N_11477,N_11413);
nand U11672 (N_11672,N_11059,N_11089);
and U11673 (N_11673,N_11397,N_11426);
nor U11674 (N_11674,N_11233,N_11407);
or U11675 (N_11675,N_11360,N_11046);
xor U11676 (N_11676,N_11432,N_11298);
nand U11677 (N_11677,N_11101,N_11027);
nor U11678 (N_11678,N_11232,N_11121);
nor U11679 (N_11679,N_11020,N_11296);
or U11680 (N_11680,N_11266,N_11060);
nor U11681 (N_11681,N_11361,N_11334);
or U11682 (N_11682,N_11163,N_11186);
or U11683 (N_11683,N_11115,N_11313);
nand U11684 (N_11684,N_11220,N_11110);
and U11685 (N_11685,N_11074,N_11238);
and U11686 (N_11686,N_11199,N_11439);
and U11687 (N_11687,N_11410,N_11200);
nand U11688 (N_11688,N_11067,N_11443);
or U11689 (N_11689,N_11216,N_11490);
nor U11690 (N_11690,N_11033,N_11090);
nor U11691 (N_11691,N_11011,N_11056);
xor U11692 (N_11692,N_11282,N_11316);
and U11693 (N_11693,N_11471,N_11149);
xor U11694 (N_11694,N_11458,N_11459);
nor U11695 (N_11695,N_11386,N_11304);
xor U11696 (N_11696,N_11332,N_11070);
nand U11697 (N_11697,N_11010,N_11098);
xor U11698 (N_11698,N_11032,N_11190);
xor U11699 (N_11699,N_11492,N_11265);
nor U11700 (N_11700,N_11180,N_11389);
and U11701 (N_11701,N_11113,N_11178);
nor U11702 (N_11702,N_11243,N_11183);
nor U11703 (N_11703,N_11062,N_11257);
nand U11704 (N_11704,N_11041,N_11138);
or U11705 (N_11705,N_11415,N_11400);
nor U11706 (N_11706,N_11030,N_11364);
or U11707 (N_11707,N_11091,N_11375);
nor U11708 (N_11708,N_11359,N_11023);
nand U11709 (N_11709,N_11161,N_11297);
xnor U11710 (N_11710,N_11205,N_11406);
or U11711 (N_11711,N_11440,N_11044);
xnor U11712 (N_11712,N_11192,N_11223);
and U11713 (N_11713,N_11392,N_11368);
xnor U11714 (N_11714,N_11001,N_11160);
nor U11715 (N_11715,N_11260,N_11213);
nor U11716 (N_11716,N_11155,N_11321);
nor U11717 (N_11717,N_11420,N_11084);
nor U11718 (N_11718,N_11169,N_11391);
or U11719 (N_11719,N_11310,N_11365);
and U11720 (N_11720,N_11096,N_11125);
xnor U11721 (N_11721,N_11281,N_11053);
nor U11722 (N_11722,N_11472,N_11131);
nand U11723 (N_11723,N_11214,N_11036);
xnor U11724 (N_11724,N_11445,N_11278);
or U11725 (N_11725,N_11236,N_11441);
nand U11726 (N_11726,N_11497,N_11245);
xnor U11727 (N_11727,N_11184,N_11208);
nand U11728 (N_11728,N_11173,N_11283);
or U11729 (N_11729,N_11069,N_11195);
nand U11730 (N_11730,N_11194,N_11286);
or U11731 (N_11731,N_11414,N_11442);
nor U11732 (N_11732,N_11047,N_11428);
nand U11733 (N_11733,N_11252,N_11119);
or U11734 (N_11734,N_11052,N_11071);
nand U11735 (N_11735,N_11306,N_11225);
or U11736 (N_11736,N_11393,N_11351);
nand U11737 (N_11737,N_11333,N_11474);
or U11738 (N_11738,N_11104,N_11468);
nand U11739 (N_11739,N_11491,N_11240);
nand U11740 (N_11740,N_11114,N_11325);
nor U11741 (N_11741,N_11387,N_11373);
nor U11742 (N_11742,N_11301,N_11305);
nor U11743 (N_11743,N_11338,N_11489);
or U11744 (N_11744,N_11106,N_11198);
nor U11745 (N_11745,N_11341,N_11450);
and U11746 (N_11746,N_11390,N_11111);
nor U11747 (N_11747,N_11015,N_11498);
nor U11748 (N_11748,N_11484,N_11456);
and U11749 (N_11749,N_11251,N_11250);
xnor U11750 (N_11750,N_11429,N_11469);
nor U11751 (N_11751,N_11012,N_11065);
nand U11752 (N_11752,N_11202,N_11255);
nand U11753 (N_11753,N_11229,N_11020);
nor U11754 (N_11754,N_11396,N_11044);
nand U11755 (N_11755,N_11018,N_11067);
or U11756 (N_11756,N_11063,N_11053);
and U11757 (N_11757,N_11336,N_11175);
nand U11758 (N_11758,N_11054,N_11297);
and U11759 (N_11759,N_11372,N_11284);
nor U11760 (N_11760,N_11297,N_11063);
nor U11761 (N_11761,N_11122,N_11270);
and U11762 (N_11762,N_11464,N_11434);
nand U11763 (N_11763,N_11236,N_11075);
nor U11764 (N_11764,N_11390,N_11339);
nor U11765 (N_11765,N_11075,N_11139);
or U11766 (N_11766,N_11400,N_11379);
xnor U11767 (N_11767,N_11465,N_11230);
xor U11768 (N_11768,N_11072,N_11132);
or U11769 (N_11769,N_11156,N_11383);
nand U11770 (N_11770,N_11487,N_11165);
xor U11771 (N_11771,N_11175,N_11414);
xnor U11772 (N_11772,N_11018,N_11315);
nand U11773 (N_11773,N_11205,N_11327);
nor U11774 (N_11774,N_11006,N_11492);
nand U11775 (N_11775,N_11251,N_11069);
nand U11776 (N_11776,N_11230,N_11245);
or U11777 (N_11777,N_11256,N_11334);
or U11778 (N_11778,N_11190,N_11008);
or U11779 (N_11779,N_11415,N_11101);
and U11780 (N_11780,N_11392,N_11002);
nand U11781 (N_11781,N_11422,N_11419);
nand U11782 (N_11782,N_11018,N_11434);
nand U11783 (N_11783,N_11315,N_11034);
xor U11784 (N_11784,N_11292,N_11320);
nor U11785 (N_11785,N_11128,N_11291);
and U11786 (N_11786,N_11183,N_11288);
and U11787 (N_11787,N_11009,N_11220);
xnor U11788 (N_11788,N_11349,N_11206);
xor U11789 (N_11789,N_11120,N_11087);
nor U11790 (N_11790,N_11087,N_11179);
or U11791 (N_11791,N_11037,N_11498);
nor U11792 (N_11792,N_11083,N_11247);
and U11793 (N_11793,N_11371,N_11119);
nor U11794 (N_11794,N_11385,N_11026);
and U11795 (N_11795,N_11125,N_11153);
nor U11796 (N_11796,N_11003,N_11483);
xor U11797 (N_11797,N_11400,N_11450);
xnor U11798 (N_11798,N_11448,N_11275);
xor U11799 (N_11799,N_11262,N_11089);
nor U11800 (N_11800,N_11063,N_11136);
nor U11801 (N_11801,N_11004,N_11443);
and U11802 (N_11802,N_11304,N_11193);
or U11803 (N_11803,N_11103,N_11061);
or U11804 (N_11804,N_11108,N_11282);
or U11805 (N_11805,N_11481,N_11177);
nand U11806 (N_11806,N_11087,N_11108);
xor U11807 (N_11807,N_11174,N_11390);
and U11808 (N_11808,N_11258,N_11153);
or U11809 (N_11809,N_11183,N_11349);
nand U11810 (N_11810,N_11040,N_11155);
xnor U11811 (N_11811,N_11263,N_11254);
and U11812 (N_11812,N_11327,N_11426);
nor U11813 (N_11813,N_11079,N_11272);
and U11814 (N_11814,N_11304,N_11317);
and U11815 (N_11815,N_11288,N_11222);
and U11816 (N_11816,N_11457,N_11030);
xnor U11817 (N_11817,N_11005,N_11497);
nand U11818 (N_11818,N_11318,N_11047);
nand U11819 (N_11819,N_11302,N_11455);
xnor U11820 (N_11820,N_11472,N_11369);
nand U11821 (N_11821,N_11363,N_11314);
nor U11822 (N_11822,N_11313,N_11053);
and U11823 (N_11823,N_11160,N_11003);
or U11824 (N_11824,N_11320,N_11219);
nor U11825 (N_11825,N_11066,N_11198);
nor U11826 (N_11826,N_11167,N_11419);
nor U11827 (N_11827,N_11304,N_11218);
and U11828 (N_11828,N_11120,N_11145);
nor U11829 (N_11829,N_11044,N_11309);
xnor U11830 (N_11830,N_11202,N_11367);
nor U11831 (N_11831,N_11042,N_11276);
nor U11832 (N_11832,N_11478,N_11373);
xor U11833 (N_11833,N_11275,N_11094);
nand U11834 (N_11834,N_11217,N_11220);
nand U11835 (N_11835,N_11346,N_11208);
nor U11836 (N_11836,N_11018,N_11280);
nand U11837 (N_11837,N_11325,N_11123);
nor U11838 (N_11838,N_11046,N_11459);
nor U11839 (N_11839,N_11174,N_11184);
nor U11840 (N_11840,N_11391,N_11090);
nand U11841 (N_11841,N_11294,N_11447);
nand U11842 (N_11842,N_11447,N_11155);
nand U11843 (N_11843,N_11342,N_11346);
and U11844 (N_11844,N_11421,N_11473);
or U11845 (N_11845,N_11087,N_11059);
nand U11846 (N_11846,N_11366,N_11278);
nand U11847 (N_11847,N_11351,N_11211);
nand U11848 (N_11848,N_11113,N_11185);
or U11849 (N_11849,N_11233,N_11249);
xnor U11850 (N_11850,N_11334,N_11180);
or U11851 (N_11851,N_11236,N_11470);
nand U11852 (N_11852,N_11082,N_11455);
xor U11853 (N_11853,N_11477,N_11486);
or U11854 (N_11854,N_11078,N_11499);
nand U11855 (N_11855,N_11003,N_11481);
or U11856 (N_11856,N_11083,N_11133);
nor U11857 (N_11857,N_11012,N_11195);
and U11858 (N_11858,N_11150,N_11292);
nor U11859 (N_11859,N_11291,N_11341);
xnor U11860 (N_11860,N_11331,N_11345);
and U11861 (N_11861,N_11220,N_11499);
and U11862 (N_11862,N_11238,N_11231);
or U11863 (N_11863,N_11347,N_11119);
nor U11864 (N_11864,N_11086,N_11035);
nand U11865 (N_11865,N_11273,N_11139);
nand U11866 (N_11866,N_11232,N_11252);
or U11867 (N_11867,N_11210,N_11354);
nor U11868 (N_11868,N_11361,N_11024);
nor U11869 (N_11869,N_11415,N_11344);
or U11870 (N_11870,N_11097,N_11082);
nor U11871 (N_11871,N_11234,N_11469);
or U11872 (N_11872,N_11042,N_11325);
or U11873 (N_11873,N_11204,N_11080);
nor U11874 (N_11874,N_11396,N_11268);
xor U11875 (N_11875,N_11182,N_11327);
nor U11876 (N_11876,N_11100,N_11458);
nand U11877 (N_11877,N_11420,N_11461);
or U11878 (N_11878,N_11282,N_11046);
nor U11879 (N_11879,N_11445,N_11315);
nand U11880 (N_11880,N_11475,N_11423);
xor U11881 (N_11881,N_11423,N_11042);
or U11882 (N_11882,N_11044,N_11466);
xnor U11883 (N_11883,N_11420,N_11466);
xor U11884 (N_11884,N_11214,N_11405);
or U11885 (N_11885,N_11417,N_11095);
nor U11886 (N_11886,N_11465,N_11471);
and U11887 (N_11887,N_11304,N_11358);
xor U11888 (N_11888,N_11304,N_11310);
nand U11889 (N_11889,N_11382,N_11260);
nand U11890 (N_11890,N_11444,N_11096);
nand U11891 (N_11891,N_11452,N_11144);
nand U11892 (N_11892,N_11224,N_11351);
and U11893 (N_11893,N_11346,N_11305);
nor U11894 (N_11894,N_11076,N_11030);
or U11895 (N_11895,N_11186,N_11414);
nand U11896 (N_11896,N_11265,N_11174);
nor U11897 (N_11897,N_11288,N_11402);
and U11898 (N_11898,N_11333,N_11337);
xor U11899 (N_11899,N_11355,N_11371);
and U11900 (N_11900,N_11340,N_11107);
nand U11901 (N_11901,N_11153,N_11075);
or U11902 (N_11902,N_11332,N_11347);
nor U11903 (N_11903,N_11262,N_11305);
or U11904 (N_11904,N_11475,N_11310);
and U11905 (N_11905,N_11324,N_11233);
or U11906 (N_11906,N_11343,N_11239);
and U11907 (N_11907,N_11415,N_11133);
and U11908 (N_11908,N_11488,N_11321);
or U11909 (N_11909,N_11431,N_11090);
xor U11910 (N_11910,N_11129,N_11116);
or U11911 (N_11911,N_11283,N_11177);
xor U11912 (N_11912,N_11281,N_11171);
xnor U11913 (N_11913,N_11078,N_11379);
xnor U11914 (N_11914,N_11146,N_11075);
and U11915 (N_11915,N_11292,N_11331);
or U11916 (N_11916,N_11268,N_11105);
xor U11917 (N_11917,N_11383,N_11307);
and U11918 (N_11918,N_11037,N_11149);
and U11919 (N_11919,N_11372,N_11027);
nand U11920 (N_11920,N_11363,N_11412);
or U11921 (N_11921,N_11375,N_11440);
xor U11922 (N_11922,N_11485,N_11151);
or U11923 (N_11923,N_11270,N_11444);
nor U11924 (N_11924,N_11209,N_11431);
nor U11925 (N_11925,N_11101,N_11411);
nor U11926 (N_11926,N_11328,N_11245);
nor U11927 (N_11927,N_11214,N_11459);
nand U11928 (N_11928,N_11244,N_11269);
or U11929 (N_11929,N_11234,N_11145);
xor U11930 (N_11930,N_11108,N_11137);
nor U11931 (N_11931,N_11124,N_11202);
nor U11932 (N_11932,N_11070,N_11006);
nand U11933 (N_11933,N_11098,N_11400);
xor U11934 (N_11934,N_11108,N_11318);
and U11935 (N_11935,N_11314,N_11285);
nor U11936 (N_11936,N_11343,N_11299);
nor U11937 (N_11937,N_11296,N_11493);
or U11938 (N_11938,N_11339,N_11143);
xnor U11939 (N_11939,N_11493,N_11462);
and U11940 (N_11940,N_11272,N_11248);
or U11941 (N_11941,N_11106,N_11073);
nand U11942 (N_11942,N_11046,N_11014);
or U11943 (N_11943,N_11194,N_11378);
nand U11944 (N_11944,N_11182,N_11067);
or U11945 (N_11945,N_11327,N_11399);
nand U11946 (N_11946,N_11247,N_11250);
and U11947 (N_11947,N_11267,N_11369);
or U11948 (N_11948,N_11087,N_11403);
and U11949 (N_11949,N_11288,N_11382);
nor U11950 (N_11950,N_11415,N_11424);
or U11951 (N_11951,N_11025,N_11084);
and U11952 (N_11952,N_11055,N_11316);
nand U11953 (N_11953,N_11032,N_11138);
xor U11954 (N_11954,N_11087,N_11201);
nor U11955 (N_11955,N_11095,N_11212);
and U11956 (N_11956,N_11112,N_11401);
xnor U11957 (N_11957,N_11220,N_11370);
xor U11958 (N_11958,N_11100,N_11014);
xor U11959 (N_11959,N_11209,N_11183);
xor U11960 (N_11960,N_11060,N_11327);
nor U11961 (N_11961,N_11085,N_11405);
and U11962 (N_11962,N_11389,N_11173);
or U11963 (N_11963,N_11136,N_11331);
xnor U11964 (N_11964,N_11196,N_11405);
and U11965 (N_11965,N_11497,N_11265);
nand U11966 (N_11966,N_11371,N_11097);
nand U11967 (N_11967,N_11017,N_11255);
or U11968 (N_11968,N_11139,N_11320);
and U11969 (N_11969,N_11152,N_11373);
and U11970 (N_11970,N_11319,N_11109);
xnor U11971 (N_11971,N_11136,N_11455);
xnor U11972 (N_11972,N_11049,N_11298);
nand U11973 (N_11973,N_11443,N_11054);
and U11974 (N_11974,N_11104,N_11252);
nor U11975 (N_11975,N_11072,N_11494);
nand U11976 (N_11976,N_11137,N_11046);
xor U11977 (N_11977,N_11188,N_11017);
xnor U11978 (N_11978,N_11121,N_11005);
xor U11979 (N_11979,N_11262,N_11064);
nand U11980 (N_11980,N_11480,N_11289);
or U11981 (N_11981,N_11446,N_11481);
and U11982 (N_11982,N_11451,N_11343);
nand U11983 (N_11983,N_11406,N_11253);
nor U11984 (N_11984,N_11407,N_11230);
nor U11985 (N_11985,N_11368,N_11083);
nand U11986 (N_11986,N_11303,N_11473);
nor U11987 (N_11987,N_11273,N_11105);
xor U11988 (N_11988,N_11443,N_11387);
nor U11989 (N_11989,N_11200,N_11112);
or U11990 (N_11990,N_11400,N_11251);
xor U11991 (N_11991,N_11355,N_11220);
nor U11992 (N_11992,N_11269,N_11079);
nor U11993 (N_11993,N_11014,N_11344);
nor U11994 (N_11994,N_11223,N_11329);
and U11995 (N_11995,N_11167,N_11211);
xor U11996 (N_11996,N_11404,N_11147);
nand U11997 (N_11997,N_11027,N_11140);
or U11998 (N_11998,N_11150,N_11239);
nand U11999 (N_11999,N_11231,N_11016);
or U12000 (N_12000,N_11610,N_11919);
and U12001 (N_12001,N_11548,N_11698);
or U12002 (N_12002,N_11724,N_11668);
nand U12003 (N_12003,N_11705,N_11750);
nand U12004 (N_12004,N_11793,N_11974);
or U12005 (N_12005,N_11747,N_11581);
xnor U12006 (N_12006,N_11611,N_11700);
xnor U12007 (N_12007,N_11887,N_11563);
nand U12008 (N_12008,N_11876,N_11915);
or U12009 (N_12009,N_11766,N_11802);
xor U12010 (N_12010,N_11886,N_11808);
nor U12011 (N_12011,N_11920,N_11716);
nor U12012 (N_12012,N_11647,N_11769);
or U12013 (N_12013,N_11636,N_11584);
nand U12014 (N_12014,N_11737,N_11839);
xor U12015 (N_12015,N_11586,N_11777);
or U12016 (N_12016,N_11711,N_11686);
nor U12017 (N_12017,N_11691,N_11707);
or U12018 (N_12018,N_11824,N_11863);
and U12019 (N_12019,N_11812,N_11794);
xnor U12020 (N_12020,N_11799,N_11814);
and U12021 (N_12021,N_11651,N_11529);
nand U12022 (N_12022,N_11846,N_11740);
and U12023 (N_12023,N_11569,N_11931);
or U12024 (N_12024,N_11615,N_11639);
nand U12025 (N_12025,N_11888,N_11632);
or U12026 (N_12026,N_11922,N_11709);
nor U12027 (N_12027,N_11852,N_11589);
or U12028 (N_12028,N_11753,N_11717);
nand U12029 (N_12029,N_11556,N_11981);
nand U12030 (N_12030,N_11907,N_11619);
and U12031 (N_12031,N_11689,N_11593);
xor U12032 (N_12032,N_11996,N_11576);
xor U12033 (N_12033,N_11829,N_11507);
or U12034 (N_12034,N_11741,N_11801);
nand U12035 (N_12035,N_11976,N_11746);
nand U12036 (N_12036,N_11889,N_11940);
nand U12037 (N_12037,N_11729,N_11764);
or U12038 (N_12038,N_11966,N_11675);
nor U12039 (N_12039,N_11778,N_11834);
nor U12040 (N_12040,N_11932,N_11558);
or U12041 (N_12041,N_11728,N_11736);
xor U12042 (N_12042,N_11528,N_11683);
xnor U12043 (N_12043,N_11849,N_11553);
nor U12044 (N_12044,N_11540,N_11743);
nand U12045 (N_12045,N_11787,N_11962);
xnor U12046 (N_12046,N_11873,N_11826);
and U12047 (N_12047,N_11550,N_11993);
or U12048 (N_12048,N_11665,N_11527);
nor U12049 (N_12049,N_11908,N_11513);
or U12050 (N_12050,N_11843,N_11935);
nand U12051 (N_12051,N_11518,N_11930);
nor U12052 (N_12052,N_11688,N_11784);
nor U12053 (N_12053,N_11702,N_11517);
and U12054 (N_12054,N_11795,N_11768);
nand U12055 (N_12055,N_11516,N_11678);
xor U12056 (N_12056,N_11770,N_11850);
and U12057 (N_12057,N_11629,N_11631);
xor U12058 (N_12058,N_11898,N_11775);
or U12059 (N_12059,N_11872,N_11859);
or U12060 (N_12060,N_11882,N_11945);
nand U12061 (N_12061,N_11579,N_11505);
or U12062 (N_12062,N_11519,N_11551);
or U12063 (N_12063,N_11625,N_11995);
nand U12064 (N_12064,N_11616,N_11714);
nand U12065 (N_12065,N_11896,N_11537);
or U12066 (N_12066,N_11645,N_11967);
nand U12067 (N_12067,N_11726,N_11654);
and U12068 (N_12068,N_11817,N_11554);
xnor U12069 (N_12069,N_11597,N_11971);
nor U12070 (N_12070,N_11699,N_11687);
or U12071 (N_12071,N_11851,N_11612);
and U12072 (N_12072,N_11963,N_11938);
nand U12073 (N_12073,N_11533,N_11899);
or U12074 (N_12074,N_11900,N_11599);
or U12075 (N_12075,N_11695,N_11941);
or U12076 (N_12076,N_11649,N_11622);
xnor U12077 (N_12077,N_11708,N_11942);
nand U12078 (N_12078,N_11818,N_11975);
nand U12079 (N_12079,N_11578,N_11911);
or U12080 (N_12080,N_11662,N_11564);
nand U12081 (N_12081,N_11666,N_11992);
and U12082 (N_12082,N_11706,N_11844);
nand U12083 (N_12083,N_11943,N_11523);
xor U12084 (N_12084,N_11653,N_11701);
xnor U12085 (N_12085,N_11570,N_11500);
or U12086 (N_12086,N_11830,N_11792);
xor U12087 (N_12087,N_11956,N_11557);
nor U12088 (N_12088,N_11738,N_11949);
and U12089 (N_12089,N_11833,N_11811);
nand U12090 (N_12090,N_11803,N_11957);
and U12091 (N_12091,N_11660,N_11825);
nor U12092 (N_12092,N_11572,N_11562);
nor U12093 (N_12093,N_11838,N_11565);
xnor U12094 (N_12094,N_11539,N_11953);
or U12095 (N_12095,N_11685,N_11914);
nor U12096 (N_12096,N_11970,N_11635);
nor U12097 (N_12097,N_11917,N_11693);
nand U12098 (N_12098,N_11715,N_11878);
or U12099 (N_12099,N_11828,N_11771);
xor U12100 (N_12100,N_11982,N_11968);
and U12101 (N_12101,N_11655,N_11774);
nor U12102 (N_12102,N_11623,N_11514);
nand U12103 (N_12103,N_11865,N_11567);
or U12104 (N_12104,N_11588,N_11577);
xor U12105 (N_12105,N_11861,N_11955);
nor U12106 (N_12106,N_11763,N_11674);
nor U12107 (N_12107,N_11515,N_11696);
nand U12108 (N_12108,N_11906,N_11789);
nand U12109 (N_12109,N_11845,N_11959);
nor U12110 (N_12110,N_11697,N_11961);
nand U12111 (N_12111,N_11532,N_11827);
nor U12112 (N_12112,N_11909,N_11512);
or U12113 (N_12113,N_11721,N_11690);
or U12114 (N_12114,N_11742,N_11980);
nor U12115 (N_12115,N_11837,N_11779);
or U12116 (N_12116,N_11857,N_11757);
xor U12117 (N_12117,N_11734,N_11791);
nand U12118 (N_12118,N_11832,N_11821);
xnor U12119 (N_12119,N_11761,N_11637);
xor U12120 (N_12120,N_11985,N_11841);
or U12121 (N_12121,N_11783,N_11646);
nor U12122 (N_12122,N_11751,N_11999);
nand U12123 (N_12123,N_11923,N_11890);
nor U12124 (N_12124,N_11679,N_11680);
and U12125 (N_12125,N_11641,N_11864);
xnor U12126 (N_12126,N_11607,N_11542);
nor U12127 (N_12127,N_11511,N_11652);
nor U12128 (N_12128,N_11969,N_11541);
nand U12129 (N_12129,N_11835,N_11998);
or U12130 (N_12130,N_11853,N_11813);
and U12131 (N_12131,N_11620,N_11823);
or U12132 (N_12132,N_11718,N_11643);
nor U12133 (N_12133,N_11848,N_11991);
nor U12134 (N_12134,N_11965,N_11809);
xor U12135 (N_12135,N_11663,N_11952);
xnor U12136 (N_12136,N_11804,N_11633);
and U12137 (N_12137,N_11805,N_11608);
or U12138 (N_12138,N_11526,N_11884);
and U12139 (N_12139,N_11797,N_11860);
or U12140 (N_12140,N_11862,N_11676);
or U12141 (N_12141,N_11658,N_11925);
nor U12142 (N_12142,N_11543,N_11807);
or U12143 (N_12143,N_11671,N_11561);
nand U12144 (N_12144,N_11885,N_11524);
and U12145 (N_12145,N_11937,N_11710);
and U12146 (N_12146,N_11587,N_11781);
or U12147 (N_12147,N_11547,N_11847);
nor U12148 (N_12148,N_11936,N_11739);
and U12149 (N_12149,N_11720,N_11544);
and U12150 (N_12150,N_11765,N_11510);
or U12151 (N_12151,N_11592,N_11947);
xor U12152 (N_12152,N_11571,N_11582);
or U12153 (N_12153,N_11522,N_11595);
nand U12154 (N_12154,N_11559,N_11600);
nor U12155 (N_12155,N_11933,N_11549);
and U12156 (N_12156,N_11806,N_11950);
or U12157 (N_12157,N_11546,N_11722);
nor U12158 (N_12158,N_11928,N_11881);
or U12159 (N_12159,N_11921,N_11723);
and U12160 (N_12160,N_11583,N_11883);
nor U12161 (N_12161,N_11732,N_11972);
and U12162 (N_12162,N_11703,N_11756);
or U12163 (N_12163,N_11630,N_11901);
nand U12164 (N_12164,N_11867,N_11912);
or U12165 (N_12165,N_11712,N_11964);
nand U12166 (N_12166,N_11854,N_11893);
xor U12167 (N_12167,N_11997,N_11606);
or U12168 (N_12168,N_11749,N_11910);
nand U12169 (N_12169,N_11585,N_11684);
nor U12170 (N_12170,N_11856,N_11874);
nor U12171 (N_12171,N_11868,N_11816);
nand U12172 (N_12172,N_11754,N_11875);
nand U12173 (N_12173,N_11895,N_11744);
nand U12174 (N_12174,N_11642,N_11618);
xor U12175 (N_12175,N_11673,N_11939);
xnor U12176 (N_12176,N_11661,N_11785);
xor U12177 (N_12177,N_11798,N_11903);
xnor U12178 (N_12178,N_11638,N_11934);
nor U12179 (N_12179,N_11694,N_11815);
nand U12180 (N_12180,N_11796,N_11790);
nand U12181 (N_12181,N_11820,N_11656);
and U12182 (N_12182,N_11767,N_11759);
nor U12183 (N_12183,N_11560,N_11946);
nor U12184 (N_12184,N_11755,N_11502);
xnor U12185 (N_12185,N_11552,N_11840);
nor U12186 (N_12186,N_11760,N_11948);
xor U12187 (N_12187,N_11776,N_11509);
nand U12188 (N_12188,N_11979,N_11520);
xor U12189 (N_12189,N_11780,N_11904);
and U12190 (N_12190,N_11855,N_11704);
nor U12191 (N_12191,N_11628,N_11892);
nor U12192 (N_12192,N_11842,N_11566);
nand U12193 (N_12193,N_11989,N_11929);
nand U12194 (N_12194,N_11782,N_11535);
or U12195 (N_12195,N_11918,N_11988);
xnor U12196 (N_12196,N_11733,N_11748);
and U12197 (N_12197,N_11869,N_11731);
nand U12198 (N_12198,N_11555,N_11978);
and U12199 (N_12199,N_11905,N_11727);
xor U12200 (N_12200,N_11670,N_11621);
xor U12201 (N_12201,N_11667,N_11627);
xor U12202 (N_12202,N_11508,N_11536);
xnor U12203 (N_12203,N_11605,N_11598);
or U12204 (N_12204,N_11987,N_11538);
nand U12205 (N_12205,N_11603,N_11819);
xor U12206 (N_12206,N_11719,N_11692);
xor U12207 (N_12207,N_11530,N_11596);
nor U12208 (N_12208,N_11973,N_11640);
and U12209 (N_12209,N_11870,N_11822);
or U12210 (N_12210,N_11773,N_11677);
nand U12211 (N_12211,N_11531,N_11927);
nor U12212 (N_12212,N_11871,N_11879);
and U12213 (N_12213,N_11877,N_11573);
and U12214 (N_12214,N_11503,N_11568);
or U12215 (N_12215,N_11624,N_11594);
nand U12216 (N_12216,N_11983,N_11664);
xor U12217 (N_12217,N_11534,N_11506);
nand U12218 (N_12218,N_11713,N_11902);
or U12219 (N_12219,N_11916,N_11810);
nor U12220 (N_12220,N_11958,N_11772);
nand U12221 (N_12221,N_11659,N_11575);
xor U12222 (N_12222,N_11650,N_11545);
nor U12223 (N_12223,N_11891,N_11681);
nor U12224 (N_12224,N_11648,N_11800);
nor U12225 (N_12225,N_11574,N_11758);
nor U12226 (N_12226,N_11897,N_11672);
nand U12227 (N_12227,N_11836,N_11954);
xnor U12228 (N_12228,N_11924,N_11960);
nor U12229 (N_12229,N_11590,N_11626);
nor U12230 (N_12230,N_11669,N_11591);
nor U12231 (N_12231,N_11866,N_11501);
nor U12232 (N_12232,N_11644,N_11858);
or U12233 (N_12233,N_11634,N_11880);
or U12234 (N_12234,N_11977,N_11986);
and U12235 (N_12235,N_11788,N_11831);
and U12236 (N_12236,N_11762,N_11752);
and U12237 (N_12237,N_11913,N_11745);
or U12238 (N_12238,N_11609,N_11951);
or U12239 (N_12239,N_11682,N_11894);
nor U12240 (N_12240,N_11601,N_11602);
nor U12241 (N_12241,N_11525,N_11735);
nand U12242 (N_12242,N_11944,N_11521);
nand U12243 (N_12243,N_11984,N_11994);
nor U12244 (N_12244,N_11504,N_11786);
or U12245 (N_12245,N_11613,N_11580);
nor U12246 (N_12246,N_11926,N_11725);
and U12247 (N_12247,N_11990,N_11617);
nand U12248 (N_12248,N_11604,N_11614);
and U12249 (N_12249,N_11730,N_11657);
and U12250 (N_12250,N_11770,N_11991);
xnor U12251 (N_12251,N_11671,N_11868);
nor U12252 (N_12252,N_11790,N_11780);
nand U12253 (N_12253,N_11929,N_11655);
nor U12254 (N_12254,N_11784,N_11637);
nor U12255 (N_12255,N_11755,N_11799);
and U12256 (N_12256,N_11882,N_11859);
and U12257 (N_12257,N_11808,N_11989);
nor U12258 (N_12258,N_11921,N_11681);
and U12259 (N_12259,N_11738,N_11925);
xnor U12260 (N_12260,N_11770,N_11940);
and U12261 (N_12261,N_11973,N_11551);
xnor U12262 (N_12262,N_11516,N_11970);
or U12263 (N_12263,N_11999,N_11904);
nor U12264 (N_12264,N_11726,N_11634);
nand U12265 (N_12265,N_11932,N_11918);
xnor U12266 (N_12266,N_11946,N_11731);
nand U12267 (N_12267,N_11821,N_11554);
nor U12268 (N_12268,N_11850,N_11883);
and U12269 (N_12269,N_11588,N_11897);
and U12270 (N_12270,N_11740,N_11930);
nor U12271 (N_12271,N_11995,N_11710);
nand U12272 (N_12272,N_11840,N_11795);
nand U12273 (N_12273,N_11585,N_11607);
and U12274 (N_12274,N_11943,N_11986);
xnor U12275 (N_12275,N_11898,N_11615);
nand U12276 (N_12276,N_11835,N_11973);
or U12277 (N_12277,N_11816,N_11716);
xor U12278 (N_12278,N_11627,N_11524);
nand U12279 (N_12279,N_11834,N_11830);
or U12280 (N_12280,N_11914,N_11884);
nor U12281 (N_12281,N_11649,N_11845);
or U12282 (N_12282,N_11907,N_11877);
or U12283 (N_12283,N_11850,N_11648);
nand U12284 (N_12284,N_11998,N_11503);
nor U12285 (N_12285,N_11989,N_11863);
or U12286 (N_12286,N_11550,N_11767);
and U12287 (N_12287,N_11766,N_11933);
xor U12288 (N_12288,N_11670,N_11806);
nor U12289 (N_12289,N_11825,N_11731);
or U12290 (N_12290,N_11681,N_11611);
nor U12291 (N_12291,N_11785,N_11738);
or U12292 (N_12292,N_11891,N_11702);
or U12293 (N_12293,N_11541,N_11669);
nor U12294 (N_12294,N_11988,N_11942);
nand U12295 (N_12295,N_11769,N_11914);
nand U12296 (N_12296,N_11580,N_11895);
or U12297 (N_12297,N_11903,N_11555);
nand U12298 (N_12298,N_11726,N_11820);
or U12299 (N_12299,N_11885,N_11714);
nand U12300 (N_12300,N_11874,N_11513);
and U12301 (N_12301,N_11981,N_11885);
xnor U12302 (N_12302,N_11882,N_11595);
nand U12303 (N_12303,N_11551,N_11964);
and U12304 (N_12304,N_11675,N_11822);
nor U12305 (N_12305,N_11959,N_11994);
xor U12306 (N_12306,N_11811,N_11563);
xnor U12307 (N_12307,N_11522,N_11795);
or U12308 (N_12308,N_11919,N_11910);
nand U12309 (N_12309,N_11721,N_11546);
and U12310 (N_12310,N_11658,N_11762);
xor U12311 (N_12311,N_11578,N_11541);
and U12312 (N_12312,N_11631,N_11889);
xor U12313 (N_12313,N_11866,N_11619);
nor U12314 (N_12314,N_11745,N_11866);
or U12315 (N_12315,N_11799,N_11722);
nor U12316 (N_12316,N_11723,N_11729);
xnor U12317 (N_12317,N_11571,N_11511);
and U12318 (N_12318,N_11823,N_11934);
xnor U12319 (N_12319,N_11617,N_11785);
xor U12320 (N_12320,N_11952,N_11789);
xnor U12321 (N_12321,N_11931,N_11712);
or U12322 (N_12322,N_11976,N_11622);
or U12323 (N_12323,N_11915,N_11669);
nand U12324 (N_12324,N_11989,N_11916);
and U12325 (N_12325,N_11562,N_11506);
and U12326 (N_12326,N_11819,N_11623);
nor U12327 (N_12327,N_11866,N_11574);
nand U12328 (N_12328,N_11759,N_11922);
and U12329 (N_12329,N_11990,N_11748);
or U12330 (N_12330,N_11710,N_11872);
xor U12331 (N_12331,N_11653,N_11889);
nand U12332 (N_12332,N_11930,N_11889);
nor U12333 (N_12333,N_11600,N_11695);
or U12334 (N_12334,N_11666,N_11676);
nor U12335 (N_12335,N_11813,N_11712);
xnor U12336 (N_12336,N_11879,N_11571);
and U12337 (N_12337,N_11549,N_11924);
xnor U12338 (N_12338,N_11889,N_11587);
nor U12339 (N_12339,N_11711,N_11668);
or U12340 (N_12340,N_11585,N_11584);
xor U12341 (N_12341,N_11524,N_11997);
nor U12342 (N_12342,N_11694,N_11566);
nor U12343 (N_12343,N_11533,N_11757);
nor U12344 (N_12344,N_11721,N_11930);
or U12345 (N_12345,N_11587,N_11909);
or U12346 (N_12346,N_11560,N_11633);
and U12347 (N_12347,N_11754,N_11876);
or U12348 (N_12348,N_11981,N_11571);
or U12349 (N_12349,N_11962,N_11966);
or U12350 (N_12350,N_11569,N_11769);
nor U12351 (N_12351,N_11652,N_11995);
or U12352 (N_12352,N_11849,N_11818);
xnor U12353 (N_12353,N_11676,N_11518);
or U12354 (N_12354,N_11794,N_11979);
xnor U12355 (N_12355,N_11541,N_11933);
nand U12356 (N_12356,N_11696,N_11795);
nor U12357 (N_12357,N_11905,N_11536);
or U12358 (N_12358,N_11959,N_11740);
xor U12359 (N_12359,N_11719,N_11776);
nor U12360 (N_12360,N_11576,N_11633);
nand U12361 (N_12361,N_11536,N_11848);
or U12362 (N_12362,N_11640,N_11997);
nand U12363 (N_12363,N_11857,N_11548);
nor U12364 (N_12364,N_11635,N_11558);
or U12365 (N_12365,N_11967,N_11703);
or U12366 (N_12366,N_11553,N_11894);
or U12367 (N_12367,N_11723,N_11986);
or U12368 (N_12368,N_11781,N_11916);
or U12369 (N_12369,N_11978,N_11609);
xor U12370 (N_12370,N_11878,N_11986);
or U12371 (N_12371,N_11638,N_11849);
and U12372 (N_12372,N_11933,N_11619);
nor U12373 (N_12373,N_11721,N_11583);
or U12374 (N_12374,N_11861,N_11651);
and U12375 (N_12375,N_11641,N_11702);
and U12376 (N_12376,N_11896,N_11870);
xor U12377 (N_12377,N_11681,N_11719);
nand U12378 (N_12378,N_11550,N_11551);
nor U12379 (N_12379,N_11918,N_11758);
nand U12380 (N_12380,N_11551,N_11871);
or U12381 (N_12381,N_11810,N_11727);
xor U12382 (N_12382,N_11794,N_11784);
xnor U12383 (N_12383,N_11856,N_11712);
and U12384 (N_12384,N_11840,N_11713);
and U12385 (N_12385,N_11951,N_11790);
nor U12386 (N_12386,N_11881,N_11520);
nor U12387 (N_12387,N_11859,N_11681);
and U12388 (N_12388,N_11953,N_11698);
and U12389 (N_12389,N_11820,N_11861);
or U12390 (N_12390,N_11641,N_11516);
or U12391 (N_12391,N_11895,N_11871);
nand U12392 (N_12392,N_11501,N_11696);
or U12393 (N_12393,N_11579,N_11833);
or U12394 (N_12394,N_11898,N_11918);
xnor U12395 (N_12395,N_11664,N_11942);
or U12396 (N_12396,N_11811,N_11574);
and U12397 (N_12397,N_11849,N_11511);
and U12398 (N_12398,N_11948,N_11912);
and U12399 (N_12399,N_11663,N_11753);
nand U12400 (N_12400,N_11541,N_11687);
nor U12401 (N_12401,N_11919,N_11543);
or U12402 (N_12402,N_11741,N_11609);
and U12403 (N_12403,N_11821,N_11646);
or U12404 (N_12404,N_11506,N_11789);
xor U12405 (N_12405,N_11658,N_11568);
nor U12406 (N_12406,N_11882,N_11624);
xor U12407 (N_12407,N_11734,N_11859);
nand U12408 (N_12408,N_11589,N_11580);
nor U12409 (N_12409,N_11705,N_11587);
xnor U12410 (N_12410,N_11649,N_11979);
or U12411 (N_12411,N_11714,N_11909);
nand U12412 (N_12412,N_11561,N_11915);
xor U12413 (N_12413,N_11921,N_11606);
and U12414 (N_12414,N_11533,N_11629);
nor U12415 (N_12415,N_11825,N_11552);
xnor U12416 (N_12416,N_11621,N_11886);
or U12417 (N_12417,N_11873,N_11788);
nor U12418 (N_12418,N_11662,N_11850);
or U12419 (N_12419,N_11804,N_11634);
and U12420 (N_12420,N_11944,N_11592);
nor U12421 (N_12421,N_11769,N_11594);
nand U12422 (N_12422,N_11823,N_11725);
xnor U12423 (N_12423,N_11581,N_11624);
and U12424 (N_12424,N_11518,N_11771);
or U12425 (N_12425,N_11783,N_11770);
xnor U12426 (N_12426,N_11636,N_11558);
or U12427 (N_12427,N_11690,N_11594);
xor U12428 (N_12428,N_11652,N_11961);
xnor U12429 (N_12429,N_11761,N_11558);
nand U12430 (N_12430,N_11925,N_11886);
xor U12431 (N_12431,N_11822,N_11547);
nand U12432 (N_12432,N_11702,N_11700);
nor U12433 (N_12433,N_11650,N_11786);
or U12434 (N_12434,N_11636,N_11758);
nor U12435 (N_12435,N_11918,N_11897);
or U12436 (N_12436,N_11773,N_11518);
or U12437 (N_12437,N_11564,N_11998);
or U12438 (N_12438,N_11695,N_11936);
nor U12439 (N_12439,N_11617,N_11923);
or U12440 (N_12440,N_11641,N_11994);
and U12441 (N_12441,N_11671,N_11640);
nand U12442 (N_12442,N_11645,N_11601);
nand U12443 (N_12443,N_11829,N_11887);
nor U12444 (N_12444,N_11661,N_11573);
or U12445 (N_12445,N_11965,N_11796);
or U12446 (N_12446,N_11707,N_11639);
or U12447 (N_12447,N_11543,N_11604);
and U12448 (N_12448,N_11628,N_11832);
or U12449 (N_12449,N_11679,N_11857);
or U12450 (N_12450,N_11608,N_11867);
xnor U12451 (N_12451,N_11634,N_11706);
nor U12452 (N_12452,N_11986,N_11684);
nand U12453 (N_12453,N_11738,N_11966);
nand U12454 (N_12454,N_11769,N_11759);
or U12455 (N_12455,N_11543,N_11866);
or U12456 (N_12456,N_11749,N_11855);
or U12457 (N_12457,N_11925,N_11967);
nand U12458 (N_12458,N_11968,N_11587);
or U12459 (N_12459,N_11926,N_11960);
nor U12460 (N_12460,N_11939,N_11646);
nand U12461 (N_12461,N_11548,N_11593);
nand U12462 (N_12462,N_11889,N_11765);
nor U12463 (N_12463,N_11613,N_11683);
and U12464 (N_12464,N_11975,N_11973);
and U12465 (N_12465,N_11987,N_11631);
or U12466 (N_12466,N_11820,N_11516);
or U12467 (N_12467,N_11740,N_11505);
xnor U12468 (N_12468,N_11591,N_11965);
xor U12469 (N_12469,N_11531,N_11590);
xor U12470 (N_12470,N_11708,N_11912);
nand U12471 (N_12471,N_11939,N_11511);
nand U12472 (N_12472,N_11647,N_11987);
and U12473 (N_12473,N_11549,N_11709);
xor U12474 (N_12474,N_11739,N_11982);
or U12475 (N_12475,N_11688,N_11909);
nor U12476 (N_12476,N_11765,N_11811);
xor U12477 (N_12477,N_11940,N_11735);
xnor U12478 (N_12478,N_11663,N_11630);
xnor U12479 (N_12479,N_11976,N_11587);
nand U12480 (N_12480,N_11978,N_11810);
nor U12481 (N_12481,N_11841,N_11530);
nand U12482 (N_12482,N_11671,N_11696);
nor U12483 (N_12483,N_11860,N_11956);
nor U12484 (N_12484,N_11952,N_11708);
nor U12485 (N_12485,N_11516,N_11623);
xnor U12486 (N_12486,N_11827,N_11587);
xor U12487 (N_12487,N_11522,N_11613);
nand U12488 (N_12488,N_11609,N_11748);
xnor U12489 (N_12489,N_11695,N_11891);
or U12490 (N_12490,N_11613,N_11943);
nand U12491 (N_12491,N_11685,N_11913);
nor U12492 (N_12492,N_11994,N_11972);
and U12493 (N_12493,N_11906,N_11715);
xnor U12494 (N_12494,N_11903,N_11728);
and U12495 (N_12495,N_11619,N_11795);
xor U12496 (N_12496,N_11586,N_11990);
or U12497 (N_12497,N_11983,N_11796);
nand U12498 (N_12498,N_11621,N_11627);
or U12499 (N_12499,N_11988,N_11648);
nor U12500 (N_12500,N_12020,N_12191);
or U12501 (N_12501,N_12490,N_12031);
xnor U12502 (N_12502,N_12331,N_12400);
nor U12503 (N_12503,N_12295,N_12156);
or U12504 (N_12504,N_12014,N_12403);
xnor U12505 (N_12505,N_12284,N_12259);
xnor U12506 (N_12506,N_12055,N_12015);
or U12507 (N_12507,N_12057,N_12000);
xor U12508 (N_12508,N_12499,N_12145);
nand U12509 (N_12509,N_12243,N_12354);
xnor U12510 (N_12510,N_12387,N_12073);
and U12511 (N_12511,N_12365,N_12464);
and U12512 (N_12512,N_12416,N_12377);
and U12513 (N_12513,N_12363,N_12061);
nand U12514 (N_12514,N_12407,N_12336);
and U12515 (N_12515,N_12192,N_12009);
or U12516 (N_12516,N_12189,N_12263);
or U12517 (N_12517,N_12376,N_12090);
and U12518 (N_12518,N_12019,N_12271);
and U12519 (N_12519,N_12094,N_12116);
or U12520 (N_12520,N_12476,N_12091);
nor U12521 (N_12521,N_12383,N_12240);
nor U12522 (N_12522,N_12484,N_12109);
and U12523 (N_12523,N_12186,N_12333);
and U12524 (N_12524,N_12062,N_12451);
or U12525 (N_12525,N_12158,N_12279);
or U12526 (N_12526,N_12213,N_12220);
nand U12527 (N_12527,N_12232,N_12030);
and U12528 (N_12528,N_12023,N_12493);
or U12529 (N_12529,N_12436,N_12349);
xor U12530 (N_12530,N_12150,N_12248);
nor U12531 (N_12531,N_12390,N_12486);
or U12532 (N_12532,N_12256,N_12360);
nand U12533 (N_12533,N_12133,N_12102);
nor U12534 (N_12534,N_12089,N_12082);
xor U12535 (N_12535,N_12087,N_12016);
xnor U12536 (N_12536,N_12335,N_12478);
nand U12537 (N_12537,N_12364,N_12179);
nor U12538 (N_12538,N_12027,N_12495);
nor U12539 (N_12539,N_12404,N_12337);
or U12540 (N_12540,N_12434,N_12151);
or U12541 (N_12541,N_12190,N_12462);
nand U12542 (N_12542,N_12497,N_12393);
xor U12543 (N_12543,N_12329,N_12247);
and U12544 (N_12544,N_12018,N_12473);
nand U12545 (N_12545,N_12110,N_12032);
and U12546 (N_12546,N_12276,N_12260);
nor U12547 (N_12547,N_12305,N_12483);
nor U12548 (N_12548,N_12198,N_12037);
and U12549 (N_12549,N_12058,N_12002);
or U12550 (N_12550,N_12041,N_12107);
nand U12551 (N_12551,N_12154,N_12021);
nor U12552 (N_12552,N_12246,N_12153);
or U12553 (N_12553,N_12471,N_12217);
nand U12554 (N_12554,N_12085,N_12439);
nand U12555 (N_12555,N_12472,N_12098);
nor U12556 (N_12556,N_12287,N_12128);
and U12557 (N_12557,N_12137,N_12035);
nand U12558 (N_12558,N_12309,N_12435);
xnor U12559 (N_12559,N_12011,N_12103);
nor U12560 (N_12560,N_12455,N_12264);
nor U12561 (N_12561,N_12034,N_12199);
nand U12562 (N_12562,N_12443,N_12406);
xor U12563 (N_12563,N_12125,N_12429);
nor U12564 (N_12564,N_12398,N_12299);
or U12565 (N_12565,N_12193,N_12143);
nor U12566 (N_12566,N_12005,N_12080);
xor U12567 (N_12567,N_12384,N_12095);
and U12568 (N_12568,N_12173,N_12036);
or U12569 (N_12569,N_12210,N_12008);
nor U12570 (N_12570,N_12350,N_12083);
and U12571 (N_12571,N_12071,N_12209);
xor U12572 (N_12572,N_12458,N_12282);
xnor U12573 (N_12573,N_12289,N_12466);
and U12574 (N_12574,N_12274,N_12187);
or U12575 (N_12575,N_12425,N_12319);
and U12576 (N_12576,N_12341,N_12268);
xor U12577 (N_12577,N_12127,N_12045);
or U12578 (N_12578,N_12060,N_12132);
xnor U12579 (N_12579,N_12120,N_12303);
nor U12580 (N_12580,N_12409,N_12068);
xor U12581 (N_12581,N_12223,N_12170);
or U12582 (N_12582,N_12211,N_12053);
nand U12583 (N_12583,N_12301,N_12092);
nand U12584 (N_12584,N_12351,N_12226);
nand U12585 (N_12585,N_12347,N_12488);
or U12586 (N_12586,N_12395,N_12134);
or U12587 (N_12587,N_12261,N_12361);
nand U12588 (N_12588,N_12188,N_12148);
xnor U12589 (N_12589,N_12196,N_12251);
nand U12590 (N_12590,N_12169,N_12147);
xor U12591 (N_12591,N_12175,N_12221);
and U12592 (N_12592,N_12206,N_12070);
xor U12593 (N_12593,N_12121,N_12355);
and U12594 (N_12594,N_12026,N_12205);
or U12595 (N_12595,N_12059,N_12266);
or U12596 (N_12596,N_12230,N_12423);
nand U12597 (N_12597,N_12040,N_12123);
nand U12598 (N_12598,N_12104,N_12456);
nor U12599 (N_12599,N_12212,N_12039);
and U12600 (N_12600,N_12272,N_12482);
nor U12601 (N_12601,N_12049,N_12064);
or U12602 (N_12602,N_12214,N_12370);
or U12603 (N_12603,N_12431,N_12433);
nand U12604 (N_12604,N_12181,N_12146);
xor U12605 (N_12605,N_12385,N_12022);
and U12606 (N_12606,N_12200,N_12491);
xor U12607 (N_12607,N_12255,N_12017);
and U12608 (N_12608,N_12167,N_12496);
nand U12609 (N_12609,N_12316,N_12204);
or U12610 (N_12610,N_12281,N_12369);
xor U12611 (N_12611,N_12010,N_12114);
or U12612 (N_12612,N_12302,N_12166);
nand U12613 (N_12613,N_12029,N_12463);
and U12614 (N_12614,N_12296,N_12371);
nand U12615 (N_12615,N_12313,N_12420);
nor U12616 (N_12616,N_12131,N_12163);
nor U12617 (N_12617,N_12469,N_12076);
nand U12618 (N_12618,N_12426,N_12448);
xnor U12619 (N_12619,N_12298,N_12234);
or U12620 (N_12620,N_12449,N_12438);
and U12621 (N_12621,N_12267,N_12291);
or U12622 (N_12622,N_12208,N_12228);
xnor U12623 (N_12623,N_12388,N_12402);
nand U12624 (N_12624,N_12440,N_12124);
nand U12625 (N_12625,N_12072,N_12216);
nor U12626 (N_12626,N_12328,N_12465);
nor U12627 (N_12627,N_12115,N_12066);
xnor U12628 (N_12628,N_12392,N_12344);
xnor U12629 (N_12629,N_12273,N_12269);
xnor U12630 (N_12630,N_12479,N_12280);
and U12631 (N_12631,N_12489,N_12047);
nor U12632 (N_12632,N_12157,N_12419);
and U12633 (N_12633,N_12461,N_12160);
or U12634 (N_12634,N_12318,N_12088);
xnor U12635 (N_12635,N_12277,N_12437);
nor U12636 (N_12636,N_12044,N_12381);
nand U12637 (N_12637,N_12346,N_12470);
xnor U12638 (N_12638,N_12475,N_12174);
xnor U12639 (N_12639,N_12498,N_12038);
nor U12640 (N_12640,N_12013,N_12164);
nand U12641 (N_12641,N_12324,N_12441);
xnor U12642 (N_12642,N_12112,N_12445);
nand U12643 (N_12643,N_12321,N_12326);
xnor U12644 (N_12644,N_12306,N_12339);
and U12645 (N_12645,N_12450,N_12063);
xor U12646 (N_12646,N_12081,N_12315);
nor U12647 (N_12647,N_12399,N_12258);
nor U12648 (N_12648,N_12046,N_12359);
nor U12649 (N_12649,N_12097,N_12467);
or U12650 (N_12650,N_12065,N_12074);
nand U12651 (N_12651,N_12378,N_12161);
nor U12652 (N_12652,N_12159,N_12386);
xor U12653 (N_12653,N_12474,N_12093);
xnor U12654 (N_12654,N_12307,N_12136);
and U12655 (N_12655,N_12004,N_12101);
and U12656 (N_12656,N_12428,N_12139);
xor U12657 (N_12657,N_12086,N_12001);
xnor U12658 (N_12658,N_12487,N_12135);
xor U12659 (N_12659,N_12096,N_12140);
nor U12660 (N_12660,N_12494,N_12007);
nand U12661 (N_12661,N_12270,N_12119);
nor U12662 (N_12662,N_12457,N_12492);
nand U12663 (N_12663,N_12084,N_12310);
or U12664 (N_12664,N_12345,N_12460);
xor U12665 (N_12665,N_12452,N_12410);
and U12666 (N_12666,N_12138,N_12481);
nor U12667 (N_12667,N_12442,N_12311);
nand U12668 (N_12668,N_12118,N_12257);
nor U12669 (N_12669,N_12236,N_12184);
nand U12670 (N_12670,N_12389,N_12180);
or U12671 (N_12671,N_12283,N_12185);
nand U12672 (N_12672,N_12033,N_12394);
and U12673 (N_12673,N_12012,N_12485);
or U12674 (N_12674,N_12067,N_12300);
or U12675 (N_12675,N_12444,N_12254);
or U12676 (N_12676,N_12312,N_12340);
and U12677 (N_12677,N_12366,N_12362);
nand U12678 (N_12678,N_12353,N_12265);
and U12679 (N_12679,N_12242,N_12382);
xor U12680 (N_12680,N_12231,N_12342);
nor U12681 (N_12681,N_12227,N_12100);
nand U12682 (N_12682,N_12320,N_12024);
or U12683 (N_12683,N_12142,N_12197);
or U12684 (N_12684,N_12446,N_12178);
or U12685 (N_12685,N_12144,N_12126);
or U12686 (N_12686,N_12308,N_12468);
nor U12687 (N_12687,N_12380,N_12050);
and U12688 (N_12688,N_12357,N_12413);
nand U12689 (N_12689,N_12079,N_12338);
nor U12690 (N_12690,N_12453,N_12348);
nor U12691 (N_12691,N_12391,N_12052);
nand U12692 (N_12692,N_12373,N_12297);
and U12693 (N_12693,N_12224,N_12372);
nand U12694 (N_12694,N_12412,N_12415);
or U12695 (N_12695,N_12042,N_12414);
xnor U12696 (N_12696,N_12327,N_12253);
or U12697 (N_12697,N_12105,N_12334);
and U12698 (N_12698,N_12317,N_12106);
nor U12699 (N_12699,N_12152,N_12245);
and U12700 (N_12700,N_12219,N_12237);
nor U12701 (N_12701,N_12293,N_12422);
or U12702 (N_12702,N_12275,N_12238);
nand U12703 (N_12703,N_12235,N_12447);
nand U12704 (N_12704,N_12367,N_12172);
nand U12705 (N_12705,N_12454,N_12292);
nor U12706 (N_12706,N_12430,N_12477);
or U12707 (N_12707,N_12207,N_12028);
and U12708 (N_12708,N_12048,N_12075);
nand U12709 (N_12709,N_12294,N_12330);
and U12710 (N_12710,N_12262,N_12168);
xnor U12711 (N_12711,N_12252,N_12314);
and U12712 (N_12712,N_12288,N_12025);
nand U12713 (N_12713,N_12323,N_12356);
or U12714 (N_12714,N_12069,N_12077);
and U12715 (N_12715,N_12285,N_12286);
nor U12716 (N_12716,N_12149,N_12215);
or U12717 (N_12717,N_12352,N_12162);
and U12718 (N_12718,N_12202,N_12405);
nand U12719 (N_12719,N_12078,N_12225);
xnor U12720 (N_12720,N_12233,N_12222);
or U12721 (N_12721,N_12343,N_12141);
nor U12722 (N_12722,N_12396,N_12290);
or U12723 (N_12723,N_12241,N_12111);
or U12724 (N_12724,N_12003,N_12043);
nor U12725 (N_12725,N_12099,N_12122);
or U12726 (N_12726,N_12278,N_12201);
and U12727 (N_12727,N_12056,N_12418);
and U12728 (N_12728,N_12421,N_12417);
nor U12729 (N_12729,N_12375,N_12249);
nor U12730 (N_12730,N_12130,N_12424);
or U12731 (N_12731,N_12054,N_12325);
nand U12732 (N_12732,N_12250,N_12155);
nand U12733 (N_12733,N_12176,N_12480);
or U12734 (N_12734,N_12401,N_12332);
xnor U12735 (N_12735,N_12427,N_12194);
xnor U12736 (N_12736,N_12229,N_12368);
nand U12737 (N_12737,N_12218,N_12408);
xor U12738 (N_12738,N_12129,N_12432);
nor U12739 (N_12739,N_12177,N_12195);
and U12740 (N_12740,N_12397,N_12374);
and U12741 (N_12741,N_12051,N_12459);
nor U12742 (N_12742,N_12322,N_12006);
nor U12743 (N_12743,N_12117,N_12203);
nor U12744 (N_12744,N_12182,N_12108);
xnor U12745 (N_12745,N_12411,N_12113);
xor U12746 (N_12746,N_12379,N_12304);
xor U12747 (N_12747,N_12171,N_12358);
xnor U12748 (N_12748,N_12165,N_12239);
or U12749 (N_12749,N_12183,N_12244);
nand U12750 (N_12750,N_12190,N_12178);
nor U12751 (N_12751,N_12316,N_12091);
or U12752 (N_12752,N_12364,N_12369);
or U12753 (N_12753,N_12198,N_12428);
and U12754 (N_12754,N_12225,N_12381);
nand U12755 (N_12755,N_12249,N_12069);
or U12756 (N_12756,N_12486,N_12482);
xor U12757 (N_12757,N_12033,N_12197);
and U12758 (N_12758,N_12054,N_12365);
nor U12759 (N_12759,N_12157,N_12142);
xnor U12760 (N_12760,N_12283,N_12425);
nor U12761 (N_12761,N_12441,N_12406);
nor U12762 (N_12762,N_12169,N_12042);
or U12763 (N_12763,N_12154,N_12215);
and U12764 (N_12764,N_12395,N_12465);
or U12765 (N_12765,N_12119,N_12333);
and U12766 (N_12766,N_12276,N_12298);
xnor U12767 (N_12767,N_12016,N_12060);
and U12768 (N_12768,N_12223,N_12242);
xor U12769 (N_12769,N_12435,N_12038);
xnor U12770 (N_12770,N_12112,N_12199);
nand U12771 (N_12771,N_12242,N_12352);
nand U12772 (N_12772,N_12019,N_12059);
or U12773 (N_12773,N_12059,N_12111);
or U12774 (N_12774,N_12428,N_12427);
or U12775 (N_12775,N_12445,N_12407);
nor U12776 (N_12776,N_12414,N_12176);
nand U12777 (N_12777,N_12048,N_12130);
nand U12778 (N_12778,N_12201,N_12339);
or U12779 (N_12779,N_12008,N_12484);
nor U12780 (N_12780,N_12056,N_12042);
and U12781 (N_12781,N_12317,N_12078);
or U12782 (N_12782,N_12390,N_12369);
or U12783 (N_12783,N_12025,N_12090);
or U12784 (N_12784,N_12383,N_12095);
or U12785 (N_12785,N_12499,N_12237);
nor U12786 (N_12786,N_12109,N_12300);
nand U12787 (N_12787,N_12065,N_12232);
nand U12788 (N_12788,N_12086,N_12306);
nand U12789 (N_12789,N_12192,N_12345);
or U12790 (N_12790,N_12026,N_12169);
nand U12791 (N_12791,N_12058,N_12472);
and U12792 (N_12792,N_12115,N_12129);
xnor U12793 (N_12793,N_12436,N_12228);
nand U12794 (N_12794,N_12074,N_12367);
nor U12795 (N_12795,N_12258,N_12101);
nand U12796 (N_12796,N_12094,N_12377);
and U12797 (N_12797,N_12460,N_12335);
nand U12798 (N_12798,N_12280,N_12438);
or U12799 (N_12799,N_12191,N_12281);
and U12800 (N_12800,N_12377,N_12156);
nand U12801 (N_12801,N_12135,N_12213);
nand U12802 (N_12802,N_12137,N_12133);
and U12803 (N_12803,N_12409,N_12117);
xnor U12804 (N_12804,N_12466,N_12198);
nand U12805 (N_12805,N_12362,N_12018);
xnor U12806 (N_12806,N_12413,N_12118);
and U12807 (N_12807,N_12170,N_12236);
and U12808 (N_12808,N_12389,N_12463);
or U12809 (N_12809,N_12442,N_12056);
and U12810 (N_12810,N_12364,N_12123);
xor U12811 (N_12811,N_12034,N_12214);
nand U12812 (N_12812,N_12336,N_12301);
and U12813 (N_12813,N_12410,N_12085);
xor U12814 (N_12814,N_12424,N_12233);
nand U12815 (N_12815,N_12459,N_12173);
or U12816 (N_12816,N_12258,N_12134);
or U12817 (N_12817,N_12271,N_12110);
and U12818 (N_12818,N_12113,N_12207);
or U12819 (N_12819,N_12061,N_12021);
xor U12820 (N_12820,N_12318,N_12029);
xnor U12821 (N_12821,N_12447,N_12102);
nand U12822 (N_12822,N_12487,N_12232);
nor U12823 (N_12823,N_12426,N_12461);
and U12824 (N_12824,N_12147,N_12470);
nor U12825 (N_12825,N_12209,N_12378);
and U12826 (N_12826,N_12045,N_12121);
xnor U12827 (N_12827,N_12252,N_12036);
and U12828 (N_12828,N_12284,N_12079);
and U12829 (N_12829,N_12172,N_12029);
and U12830 (N_12830,N_12417,N_12235);
xor U12831 (N_12831,N_12456,N_12303);
or U12832 (N_12832,N_12377,N_12347);
nand U12833 (N_12833,N_12006,N_12120);
nand U12834 (N_12834,N_12142,N_12292);
and U12835 (N_12835,N_12010,N_12058);
nand U12836 (N_12836,N_12314,N_12167);
and U12837 (N_12837,N_12422,N_12301);
nand U12838 (N_12838,N_12026,N_12320);
nor U12839 (N_12839,N_12300,N_12043);
or U12840 (N_12840,N_12051,N_12219);
and U12841 (N_12841,N_12479,N_12400);
or U12842 (N_12842,N_12190,N_12304);
nor U12843 (N_12843,N_12148,N_12440);
nand U12844 (N_12844,N_12463,N_12145);
and U12845 (N_12845,N_12014,N_12130);
or U12846 (N_12846,N_12088,N_12496);
nor U12847 (N_12847,N_12498,N_12050);
or U12848 (N_12848,N_12051,N_12101);
and U12849 (N_12849,N_12366,N_12051);
nor U12850 (N_12850,N_12475,N_12224);
xor U12851 (N_12851,N_12366,N_12137);
nor U12852 (N_12852,N_12133,N_12398);
xnor U12853 (N_12853,N_12314,N_12123);
or U12854 (N_12854,N_12468,N_12193);
and U12855 (N_12855,N_12036,N_12055);
nand U12856 (N_12856,N_12334,N_12263);
nand U12857 (N_12857,N_12403,N_12333);
and U12858 (N_12858,N_12287,N_12334);
nand U12859 (N_12859,N_12222,N_12496);
xor U12860 (N_12860,N_12474,N_12133);
or U12861 (N_12861,N_12383,N_12025);
or U12862 (N_12862,N_12113,N_12370);
or U12863 (N_12863,N_12139,N_12403);
and U12864 (N_12864,N_12151,N_12485);
nor U12865 (N_12865,N_12494,N_12175);
xor U12866 (N_12866,N_12149,N_12128);
xor U12867 (N_12867,N_12282,N_12467);
nand U12868 (N_12868,N_12300,N_12474);
xor U12869 (N_12869,N_12327,N_12456);
nand U12870 (N_12870,N_12380,N_12329);
nor U12871 (N_12871,N_12145,N_12302);
nand U12872 (N_12872,N_12124,N_12024);
or U12873 (N_12873,N_12448,N_12386);
nor U12874 (N_12874,N_12222,N_12490);
xnor U12875 (N_12875,N_12130,N_12341);
nand U12876 (N_12876,N_12356,N_12139);
nand U12877 (N_12877,N_12263,N_12273);
xor U12878 (N_12878,N_12356,N_12401);
and U12879 (N_12879,N_12332,N_12131);
xor U12880 (N_12880,N_12065,N_12372);
nand U12881 (N_12881,N_12266,N_12229);
xor U12882 (N_12882,N_12044,N_12378);
nand U12883 (N_12883,N_12024,N_12209);
nand U12884 (N_12884,N_12052,N_12198);
xor U12885 (N_12885,N_12119,N_12092);
nand U12886 (N_12886,N_12211,N_12109);
and U12887 (N_12887,N_12289,N_12444);
xnor U12888 (N_12888,N_12402,N_12410);
or U12889 (N_12889,N_12118,N_12343);
or U12890 (N_12890,N_12459,N_12415);
and U12891 (N_12891,N_12020,N_12195);
and U12892 (N_12892,N_12222,N_12074);
nand U12893 (N_12893,N_12143,N_12479);
nand U12894 (N_12894,N_12188,N_12475);
xnor U12895 (N_12895,N_12422,N_12446);
nand U12896 (N_12896,N_12086,N_12205);
xor U12897 (N_12897,N_12051,N_12152);
and U12898 (N_12898,N_12138,N_12111);
and U12899 (N_12899,N_12125,N_12340);
nand U12900 (N_12900,N_12365,N_12386);
and U12901 (N_12901,N_12387,N_12376);
and U12902 (N_12902,N_12434,N_12098);
or U12903 (N_12903,N_12366,N_12402);
nor U12904 (N_12904,N_12189,N_12082);
or U12905 (N_12905,N_12222,N_12225);
or U12906 (N_12906,N_12031,N_12308);
xor U12907 (N_12907,N_12445,N_12472);
nand U12908 (N_12908,N_12129,N_12229);
nand U12909 (N_12909,N_12411,N_12176);
or U12910 (N_12910,N_12398,N_12406);
and U12911 (N_12911,N_12462,N_12047);
or U12912 (N_12912,N_12353,N_12345);
xnor U12913 (N_12913,N_12298,N_12046);
xor U12914 (N_12914,N_12173,N_12352);
and U12915 (N_12915,N_12390,N_12066);
nor U12916 (N_12916,N_12044,N_12247);
or U12917 (N_12917,N_12373,N_12323);
nand U12918 (N_12918,N_12397,N_12345);
xor U12919 (N_12919,N_12220,N_12480);
nand U12920 (N_12920,N_12188,N_12015);
or U12921 (N_12921,N_12246,N_12307);
or U12922 (N_12922,N_12390,N_12490);
and U12923 (N_12923,N_12130,N_12088);
or U12924 (N_12924,N_12428,N_12142);
nand U12925 (N_12925,N_12269,N_12390);
nor U12926 (N_12926,N_12304,N_12347);
or U12927 (N_12927,N_12031,N_12351);
or U12928 (N_12928,N_12368,N_12381);
and U12929 (N_12929,N_12476,N_12318);
xnor U12930 (N_12930,N_12381,N_12197);
nand U12931 (N_12931,N_12295,N_12481);
xor U12932 (N_12932,N_12226,N_12342);
and U12933 (N_12933,N_12009,N_12197);
xnor U12934 (N_12934,N_12465,N_12426);
xor U12935 (N_12935,N_12467,N_12216);
xor U12936 (N_12936,N_12153,N_12012);
or U12937 (N_12937,N_12233,N_12088);
or U12938 (N_12938,N_12240,N_12342);
nor U12939 (N_12939,N_12154,N_12066);
xor U12940 (N_12940,N_12275,N_12114);
and U12941 (N_12941,N_12190,N_12478);
and U12942 (N_12942,N_12276,N_12005);
xnor U12943 (N_12943,N_12321,N_12236);
and U12944 (N_12944,N_12336,N_12432);
and U12945 (N_12945,N_12278,N_12188);
xor U12946 (N_12946,N_12213,N_12238);
nor U12947 (N_12947,N_12484,N_12257);
nor U12948 (N_12948,N_12218,N_12121);
and U12949 (N_12949,N_12395,N_12101);
nand U12950 (N_12950,N_12165,N_12285);
or U12951 (N_12951,N_12314,N_12390);
and U12952 (N_12952,N_12157,N_12216);
or U12953 (N_12953,N_12089,N_12154);
nand U12954 (N_12954,N_12400,N_12495);
and U12955 (N_12955,N_12353,N_12403);
nand U12956 (N_12956,N_12213,N_12419);
or U12957 (N_12957,N_12240,N_12097);
nand U12958 (N_12958,N_12396,N_12184);
xnor U12959 (N_12959,N_12212,N_12080);
xnor U12960 (N_12960,N_12159,N_12242);
nand U12961 (N_12961,N_12451,N_12453);
xor U12962 (N_12962,N_12374,N_12188);
nor U12963 (N_12963,N_12044,N_12229);
nor U12964 (N_12964,N_12328,N_12247);
nor U12965 (N_12965,N_12459,N_12306);
and U12966 (N_12966,N_12167,N_12465);
nand U12967 (N_12967,N_12262,N_12228);
nor U12968 (N_12968,N_12375,N_12234);
xnor U12969 (N_12969,N_12385,N_12084);
nand U12970 (N_12970,N_12007,N_12218);
nor U12971 (N_12971,N_12211,N_12382);
nor U12972 (N_12972,N_12278,N_12143);
nand U12973 (N_12973,N_12353,N_12065);
nand U12974 (N_12974,N_12002,N_12311);
or U12975 (N_12975,N_12257,N_12151);
nor U12976 (N_12976,N_12293,N_12012);
nor U12977 (N_12977,N_12097,N_12378);
nor U12978 (N_12978,N_12009,N_12485);
and U12979 (N_12979,N_12275,N_12268);
nor U12980 (N_12980,N_12218,N_12220);
or U12981 (N_12981,N_12334,N_12270);
and U12982 (N_12982,N_12472,N_12147);
nor U12983 (N_12983,N_12438,N_12412);
nor U12984 (N_12984,N_12230,N_12486);
and U12985 (N_12985,N_12257,N_12368);
xnor U12986 (N_12986,N_12286,N_12169);
xor U12987 (N_12987,N_12155,N_12019);
nand U12988 (N_12988,N_12452,N_12172);
xnor U12989 (N_12989,N_12279,N_12061);
nand U12990 (N_12990,N_12471,N_12429);
xor U12991 (N_12991,N_12376,N_12267);
and U12992 (N_12992,N_12326,N_12051);
xor U12993 (N_12993,N_12137,N_12297);
or U12994 (N_12994,N_12422,N_12027);
or U12995 (N_12995,N_12326,N_12231);
or U12996 (N_12996,N_12026,N_12036);
xor U12997 (N_12997,N_12405,N_12471);
nor U12998 (N_12998,N_12477,N_12360);
xor U12999 (N_12999,N_12374,N_12447);
xor U13000 (N_13000,N_12706,N_12858);
or U13001 (N_13001,N_12804,N_12595);
nand U13002 (N_13002,N_12880,N_12619);
nand U13003 (N_13003,N_12782,N_12932);
xor U13004 (N_13004,N_12814,N_12790);
nor U13005 (N_13005,N_12751,N_12660);
nand U13006 (N_13006,N_12950,N_12999);
or U13007 (N_13007,N_12991,N_12519);
nor U13008 (N_13008,N_12979,N_12635);
nand U13009 (N_13009,N_12652,N_12793);
nor U13010 (N_13010,N_12864,N_12733);
nand U13011 (N_13011,N_12511,N_12621);
nor U13012 (N_13012,N_12678,N_12644);
nor U13013 (N_13013,N_12745,N_12926);
or U13014 (N_13014,N_12759,N_12765);
nand U13015 (N_13015,N_12590,N_12761);
or U13016 (N_13016,N_12506,N_12549);
nor U13017 (N_13017,N_12885,N_12539);
and U13018 (N_13018,N_12515,N_12617);
nand U13019 (N_13019,N_12851,N_12871);
nor U13020 (N_13020,N_12682,N_12625);
xor U13021 (N_13021,N_12683,N_12696);
or U13022 (N_13022,N_12965,N_12879);
or U13023 (N_13023,N_12513,N_12943);
or U13024 (N_13024,N_12768,N_12591);
xor U13025 (N_13025,N_12921,N_12523);
nand U13026 (N_13026,N_12666,N_12764);
or U13027 (N_13027,N_12658,N_12822);
and U13028 (N_13028,N_12839,N_12630);
xnor U13029 (N_13029,N_12976,N_12620);
nor U13030 (N_13030,N_12556,N_12972);
xnor U13031 (N_13031,N_12785,N_12881);
and U13032 (N_13032,N_12604,N_12889);
nor U13033 (N_13033,N_12998,N_12656);
or U13034 (N_13034,N_12651,N_12674);
nor U13035 (N_13035,N_12989,N_12925);
and U13036 (N_13036,N_12747,N_12542);
xnor U13037 (N_13037,N_12525,N_12909);
nor U13038 (N_13038,N_12895,N_12888);
and U13039 (N_13039,N_12918,N_12924);
nor U13040 (N_13040,N_12748,N_12521);
and U13041 (N_13041,N_12994,N_12891);
or U13042 (N_13042,N_12802,N_12899);
xnor U13043 (N_13043,N_12754,N_12900);
or U13044 (N_13044,N_12529,N_12964);
or U13045 (N_13045,N_12775,N_12801);
nor U13046 (N_13046,N_12912,N_12984);
or U13047 (N_13047,N_12783,N_12601);
nor U13048 (N_13048,N_12948,N_12520);
nand U13049 (N_13049,N_12739,N_12993);
nand U13050 (N_13050,N_12530,N_12954);
and U13051 (N_13051,N_12574,N_12770);
and U13052 (N_13052,N_12815,N_12548);
nand U13053 (N_13053,N_12892,N_12813);
and U13054 (N_13054,N_12585,N_12531);
nor U13055 (N_13055,N_12659,N_12504);
or U13056 (N_13056,N_12740,N_12843);
or U13057 (N_13057,N_12809,N_12634);
nor U13058 (N_13058,N_12526,N_12812);
or U13059 (N_13059,N_12896,N_12821);
or U13060 (N_13060,N_12949,N_12704);
and U13061 (N_13061,N_12712,N_12631);
xnor U13062 (N_13062,N_12772,N_12586);
xor U13063 (N_13063,N_12942,N_12614);
and U13064 (N_13064,N_12654,N_12805);
and U13065 (N_13065,N_12616,N_12850);
and U13066 (N_13066,N_12705,N_12940);
or U13067 (N_13067,N_12811,N_12675);
or U13068 (N_13068,N_12834,N_12847);
or U13069 (N_13069,N_12581,N_12597);
and U13070 (N_13070,N_12509,N_12600);
nand U13071 (N_13071,N_12780,N_12941);
or U13072 (N_13072,N_12981,N_12958);
nand U13073 (N_13073,N_12810,N_12860);
or U13074 (N_13074,N_12919,N_12632);
xor U13075 (N_13075,N_12898,N_12605);
xor U13076 (N_13076,N_12800,N_12671);
or U13077 (N_13077,N_12835,N_12612);
or U13078 (N_13078,N_12622,N_12707);
nor U13079 (N_13079,N_12870,N_12787);
nor U13080 (N_13080,N_12867,N_12829);
xnor U13081 (N_13081,N_12746,N_12732);
nand U13082 (N_13082,N_12749,N_12956);
nor U13083 (N_13083,N_12645,N_12594);
nand U13084 (N_13084,N_12767,N_12663);
nor U13085 (N_13085,N_12697,N_12778);
and U13086 (N_13086,N_12611,N_12971);
or U13087 (N_13087,N_12615,N_12987);
and U13088 (N_13088,N_12866,N_12758);
nand U13089 (N_13089,N_12514,N_12568);
xnor U13090 (N_13090,N_12587,N_12657);
nand U13091 (N_13091,N_12540,N_12545);
xnor U13092 (N_13092,N_12827,N_12575);
xor U13093 (N_13093,N_12708,N_12555);
nor U13094 (N_13094,N_12788,N_12757);
xnor U13095 (N_13095,N_12524,N_12840);
xor U13096 (N_13096,N_12823,N_12856);
nor U13097 (N_13097,N_12922,N_12570);
and U13098 (N_13098,N_12838,N_12854);
and U13099 (N_13099,N_12502,N_12522);
and U13100 (N_13100,N_12853,N_12642);
or U13101 (N_13101,N_12893,N_12546);
or U13102 (N_13102,N_12518,N_12565);
and U13103 (N_13103,N_12558,N_12983);
nor U13104 (N_13104,N_12716,N_12974);
and U13105 (N_13105,N_12828,N_12884);
or U13106 (N_13106,N_12537,N_12677);
and U13107 (N_13107,N_12820,N_12527);
nor U13108 (N_13108,N_12737,N_12640);
xor U13109 (N_13109,N_12848,N_12613);
or U13110 (N_13110,N_12966,N_12734);
nand U13111 (N_13111,N_12883,N_12653);
nor U13112 (N_13112,N_12859,N_12992);
nor U13113 (N_13113,N_12583,N_12725);
or U13114 (N_13114,N_12936,N_12503);
or U13115 (N_13115,N_12953,N_12929);
or U13116 (N_13116,N_12855,N_12934);
xor U13117 (N_13117,N_12512,N_12544);
and U13118 (N_13118,N_12661,N_12698);
or U13119 (N_13119,N_12554,N_12774);
nor U13120 (N_13120,N_12844,N_12862);
or U13121 (N_13121,N_12903,N_12536);
and U13122 (N_13122,N_12599,N_12711);
nor U13123 (N_13123,N_12627,N_12636);
and U13124 (N_13124,N_12562,N_12593);
nor U13125 (N_13125,N_12869,N_12608);
nor U13126 (N_13126,N_12559,N_12927);
nand U13127 (N_13127,N_12904,N_12873);
nand U13128 (N_13128,N_12908,N_12715);
or U13129 (N_13129,N_12944,N_12959);
nand U13130 (N_13130,N_12569,N_12670);
nor U13131 (N_13131,N_12730,N_12628);
nand U13132 (N_13132,N_12500,N_12731);
nor U13133 (N_13133,N_12985,N_12863);
nor U13134 (N_13134,N_12945,N_12508);
and U13135 (N_13135,N_12803,N_12607);
nor U13136 (N_13136,N_12849,N_12962);
xnor U13137 (N_13137,N_12639,N_12997);
nand U13138 (N_13138,N_12799,N_12664);
and U13139 (N_13139,N_12824,N_12741);
and U13140 (N_13140,N_12794,N_12996);
xnor U13141 (N_13141,N_12550,N_12669);
xnor U13142 (N_13142,N_12763,N_12626);
and U13143 (N_13143,N_12955,N_12872);
nor U13144 (N_13144,N_12938,N_12875);
or U13145 (N_13145,N_12750,N_12641);
xnor U13146 (N_13146,N_12781,N_12786);
nor U13147 (N_13147,N_12609,N_12906);
nor U13148 (N_13148,N_12973,N_12700);
or U13149 (N_13149,N_12744,N_12655);
or U13150 (N_13150,N_12833,N_12886);
nor U13151 (N_13151,N_12582,N_12543);
nor U13152 (N_13152,N_12967,N_12982);
or U13153 (N_13153,N_12578,N_12687);
nand U13154 (N_13154,N_12907,N_12894);
or U13155 (N_13155,N_12784,N_12986);
xor U13156 (N_13156,N_12714,N_12818);
nand U13157 (N_13157,N_12951,N_12905);
nor U13158 (N_13158,N_12576,N_12501);
xor U13159 (N_13159,N_12939,N_12773);
or U13160 (N_13160,N_12566,N_12728);
and U13161 (N_13161,N_12792,N_12742);
and U13162 (N_13162,N_12723,N_12977);
nor U13163 (N_13163,N_12975,N_12830);
or U13164 (N_13164,N_12807,N_12933);
nand U13165 (N_13165,N_12685,N_12673);
or U13166 (N_13166,N_12533,N_12692);
and U13167 (N_13167,N_12686,N_12680);
nand U13168 (N_13168,N_12573,N_12861);
nor U13169 (N_13169,N_12688,N_12571);
xnor U13170 (N_13170,N_12534,N_12897);
and U13171 (N_13171,N_12695,N_12797);
nor U13172 (N_13172,N_12720,N_12755);
and U13173 (N_13173,N_12703,N_12946);
or U13174 (N_13174,N_12567,N_12738);
xnor U13175 (N_13175,N_12505,N_12541);
or U13176 (N_13176,N_12960,N_12817);
and U13177 (N_13177,N_12588,N_12980);
xnor U13178 (N_13178,N_12920,N_12769);
and U13179 (N_13179,N_12845,N_12721);
nand U13180 (N_13180,N_12563,N_12719);
nor U13181 (N_13181,N_12910,N_12650);
nand U13182 (N_13182,N_12766,N_12667);
nand U13183 (N_13183,N_12798,N_12836);
nand U13184 (N_13184,N_12557,N_12507);
nand U13185 (N_13185,N_12572,N_12694);
nor U13186 (N_13186,N_12681,N_12832);
nand U13187 (N_13187,N_12825,N_12961);
and U13188 (N_13188,N_12887,N_12726);
or U13189 (N_13189,N_12729,N_12679);
nand U13190 (N_13190,N_12935,N_12646);
nor U13191 (N_13191,N_12624,N_12710);
nor U13192 (N_13192,N_12865,N_12779);
nor U13193 (N_13193,N_12735,N_12874);
nand U13194 (N_13194,N_12672,N_12831);
nor U13195 (N_13195,N_12930,N_12618);
nand U13196 (N_13196,N_12796,N_12701);
or U13197 (N_13197,N_12647,N_12722);
and U13198 (N_13198,N_12789,N_12819);
nand U13199 (N_13199,N_12995,N_12806);
and U13200 (N_13200,N_12913,N_12517);
nand U13201 (N_13201,N_12771,N_12547);
xor U13202 (N_13202,N_12516,N_12528);
xor U13203 (N_13203,N_12643,N_12978);
nor U13204 (N_13204,N_12676,N_12753);
nand U13205 (N_13205,N_12691,N_12963);
nor U13206 (N_13206,N_12990,N_12957);
xor U13207 (N_13207,N_12752,N_12876);
nor U13208 (N_13208,N_12602,N_12648);
nand U13209 (N_13209,N_12551,N_12841);
nor U13210 (N_13210,N_12917,N_12510);
nor U13211 (N_13211,N_12842,N_12902);
or U13212 (N_13212,N_12606,N_12577);
and U13213 (N_13213,N_12736,N_12743);
nand U13214 (N_13214,N_12727,N_12580);
and U13215 (N_13215,N_12564,N_12532);
and U13216 (N_13216,N_12603,N_12552);
nand U13217 (N_13217,N_12756,N_12762);
xnor U13218 (N_13218,N_12901,N_12791);
nand U13219 (N_13219,N_12535,N_12584);
nor U13220 (N_13220,N_12713,N_12988);
nor U13221 (N_13221,N_12633,N_12560);
and U13222 (N_13222,N_12665,N_12969);
xnor U13223 (N_13223,N_12553,N_12699);
nor U13224 (N_13224,N_12637,N_12776);
nand U13225 (N_13225,N_12968,N_12684);
and U13226 (N_13226,N_12914,N_12852);
and U13227 (N_13227,N_12837,N_12931);
nor U13228 (N_13228,N_12649,N_12808);
nand U13229 (N_13229,N_12846,N_12598);
nor U13230 (N_13230,N_12868,N_12693);
nor U13231 (N_13231,N_12857,N_12878);
or U13232 (N_13232,N_12724,N_12561);
or U13233 (N_13233,N_12916,N_12911);
and U13234 (N_13234,N_12826,N_12610);
xnor U13235 (N_13235,N_12717,N_12947);
and U13236 (N_13236,N_12718,N_12596);
or U13237 (N_13237,N_12702,N_12662);
and U13238 (N_13238,N_12579,N_12690);
or U13239 (N_13239,N_12709,N_12777);
and U13240 (N_13240,N_12760,N_12538);
or U13241 (N_13241,N_12668,N_12623);
or U13242 (N_13242,N_12915,N_12638);
or U13243 (N_13243,N_12928,N_12816);
or U13244 (N_13244,N_12923,N_12589);
and U13245 (N_13245,N_12592,N_12689);
nor U13246 (N_13246,N_12795,N_12629);
nand U13247 (N_13247,N_12882,N_12890);
nor U13248 (N_13248,N_12970,N_12952);
nor U13249 (N_13249,N_12877,N_12937);
and U13250 (N_13250,N_12796,N_12901);
nand U13251 (N_13251,N_12535,N_12883);
nand U13252 (N_13252,N_12983,N_12596);
and U13253 (N_13253,N_12726,N_12945);
nor U13254 (N_13254,N_12567,N_12627);
nor U13255 (N_13255,N_12864,N_12555);
nor U13256 (N_13256,N_12987,N_12699);
xor U13257 (N_13257,N_12914,N_12982);
or U13258 (N_13258,N_12569,N_12845);
or U13259 (N_13259,N_12806,N_12720);
nand U13260 (N_13260,N_12970,N_12732);
nor U13261 (N_13261,N_12822,N_12595);
nand U13262 (N_13262,N_12614,N_12912);
or U13263 (N_13263,N_12643,N_12897);
nand U13264 (N_13264,N_12740,N_12710);
nor U13265 (N_13265,N_12880,N_12669);
xor U13266 (N_13266,N_12509,N_12938);
nor U13267 (N_13267,N_12765,N_12578);
xor U13268 (N_13268,N_12741,N_12991);
xor U13269 (N_13269,N_12794,N_12617);
xor U13270 (N_13270,N_12548,N_12971);
and U13271 (N_13271,N_12843,N_12618);
and U13272 (N_13272,N_12540,N_12841);
nor U13273 (N_13273,N_12716,N_12515);
and U13274 (N_13274,N_12809,N_12622);
xor U13275 (N_13275,N_12846,N_12627);
and U13276 (N_13276,N_12794,N_12684);
and U13277 (N_13277,N_12850,N_12697);
xor U13278 (N_13278,N_12857,N_12788);
xnor U13279 (N_13279,N_12695,N_12863);
and U13280 (N_13280,N_12523,N_12606);
nor U13281 (N_13281,N_12585,N_12546);
nand U13282 (N_13282,N_12652,N_12957);
and U13283 (N_13283,N_12632,N_12801);
nand U13284 (N_13284,N_12962,N_12715);
and U13285 (N_13285,N_12671,N_12596);
and U13286 (N_13286,N_12630,N_12776);
xnor U13287 (N_13287,N_12868,N_12660);
and U13288 (N_13288,N_12542,N_12778);
and U13289 (N_13289,N_12927,N_12518);
nor U13290 (N_13290,N_12543,N_12987);
or U13291 (N_13291,N_12960,N_12517);
nand U13292 (N_13292,N_12627,N_12925);
nor U13293 (N_13293,N_12926,N_12620);
xnor U13294 (N_13294,N_12535,N_12930);
or U13295 (N_13295,N_12638,N_12770);
xor U13296 (N_13296,N_12869,N_12694);
nor U13297 (N_13297,N_12941,N_12516);
nor U13298 (N_13298,N_12942,N_12966);
xor U13299 (N_13299,N_12571,N_12696);
or U13300 (N_13300,N_12882,N_12556);
nand U13301 (N_13301,N_12816,N_12814);
or U13302 (N_13302,N_12604,N_12677);
nand U13303 (N_13303,N_12619,N_12793);
nand U13304 (N_13304,N_12749,N_12733);
or U13305 (N_13305,N_12637,N_12564);
xor U13306 (N_13306,N_12779,N_12965);
xnor U13307 (N_13307,N_12617,N_12573);
nand U13308 (N_13308,N_12718,N_12981);
nand U13309 (N_13309,N_12666,N_12846);
xor U13310 (N_13310,N_12698,N_12793);
nor U13311 (N_13311,N_12935,N_12600);
nor U13312 (N_13312,N_12823,N_12661);
nand U13313 (N_13313,N_12551,N_12567);
xnor U13314 (N_13314,N_12871,N_12743);
or U13315 (N_13315,N_12692,N_12964);
nand U13316 (N_13316,N_12769,N_12676);
and U13317 (N_13317,N_12685,N_12897);
and U13318 (N_13318,N_12707,N_12826);
and U13319 (N_13319,N_12700,N_12995);
or U13320 (N_13320,N_12831,N_12760);
nor U13321 (N_13321,N_12616,N_12908);
and U13322 (N_13322,N_12595,N_12722);
nand U13323 (N_13323,N_12892,N_12596);
xor U13324 (N_13324,N_12806,N_12627);
and U13325 (N_13325,N_12602,N_12608);
or U13326 (N_13326,N_12781,N_12910);
xnor U13327 (N_13327,N_12678,N_12705);
nor U13328 (N_13328,N_12959,N_12779);
or U13329 (N_13329,N_12611,N_12636);
xnor U13330 (N_13330,N_12584,N_12709);
nand U13331 (N_13331,N_12513,N_12975);
xor U13332 (N_13332,N_12518,N_12682);
or U13333 (N_13333,N_12716,N_12637);
and U13334 (N_13334,N_12846,N_12739);
or U13335 (N_13335,N_12627,N_12755);
and U13336 (N_13336,N_12842,N_12834);
xnor U13337 (N_13337,N_12854,N_12529);
nand U13338 (N_13338,N_12953,N_12944);
and U13339 (N_13339,N_12857,N_12511);
nand U13340 (N_13340,N_12657,N_12894);
xnor U13341 (N_13341,N_12876,N_12557);
nor U13342 (N_13342,N_12995,N_12721);
or U13343 (N_13343,N_12948,N_12518);
nand U13344 (N_13344,N_12516,N_12633);
nand U13345 (N_13345,N_12534,N_12877);
and U13346 (N_13346,N_12888,N_12795);
or U13347 (N_13347,N_12621,N_12559);
or U13348 (N_13348,N_12534,N_12927);
or U13349 (N_13349,N_12920,N_12594);
nand U13350 (N_13350,N_12862,N_12722);
or U13351 (N_13351,N_12527,N_12714);
nand U13352 (N_13352,N_12502,N_12770);
xnor U13353 (N_13353,N_12760,N_12733);
nor U13354 (N_13354,N_12831,N_12752);
and U13355 (N_13355,N_12950,N_12681);
xnor U13356 (N_13356,N_12573,N_12910);
xor U13357 (N_13357,N_12799,N_12541);
or U13358 (N_13358,N_12731,N_12637);
xor U13359 (N_13359,N_12626,N_12802);
and U13360 (N_13360,N_12950,N_12796);
or U13361 (N_13361,N_12570,N_12594);
xnor U13362 (N_13362,N_12661,N_12601);
nand U13363 (N_13363,N_12744,N_12820);
xor U13364 (N_13364,N_12515,N_12674);
nor U13365 (N_13365,N_12677,N_12725);
or U13366 (N_13366,N_12602,N_12843);
and U13367 (N_13367,N_12858,N_12829);
nand U13368 (N_13368,N_12620,N_12638);
nand U13369 (N_13369,N_12650,N_12937);
or U13370 (N_13370,N_12626,N_12945);
xor U13371 (N_13371,N_12567,N_12630);
nor U13372 (N_13372,N_12716,N_12525);
nor U13373 (N_13373,N_12981,N_12974);
and U13374 (N_13374,N_12590,N_12560);
nand U13375 (N_13375,N_12936,N_12975);
nand U13376 (N_13376,N_12910,N_12808);
xnor U13377 (N_13377,N_12501,N_12565);
and U13378 (N_13378,N_12744,N_12919);
and U13379 (N_13379,N_12557,N_12671);
xnor U13380 (N_13380,N_12843,N_12951);
nor U13381 (N_13381,N_12513,N_12573);
or U13382 (N_13382,N_12689,N_12783);
and U13383 (N_13383,N_12608,N_12777);
or U13384 (N_13384,N_12775,N_12964);
nand U13385 (N_13385,N_12662,N_12632);
xnor U13386 (N_13386,N_12968,N_12537);
xnor U13387 (N_13387,N_12794,N_12804);
and U13388 (N_13388,N_12987,N_12759);
xor U13389 (N_13389,N_12954,N_12748);
and U13390 (N_13390,N_12810,N_12633);
nand U13391 (N_13391,N_12519,N_12693);
and U13392 (N_13392,N_12557,N_12826);
nand U13393 (N_13393,N_12846,N_12872);
nand U13394 (N_13394,N_12545,N_12862);
and U13395 (N_13395,N_12502,N_12585);
nand U13396 (N_13396,N_12744,N_12894);
nand U13397 (N_13397,N_12516,N_12960);
and U13398 (N_13398,N_12672,N_12684);
and U13399 (N_13399,N_12993,N_12604);
and U13400 (N_13400,N_12892,N_12798);
and U13401 (N_13401,N_12821,N_12850);
or U13402 (N_13402,N_12783,N_12754);
or U13403 (N_13403,N_12872,N_12733);
xnor U13404 (N_13404,N_12583,N_12560);
nor U13405 (N_13405,N_12627,N_12993);
and U13406 (N_13406,N_12525,N_12930);
nand U13407 (N_13407,N_12635,N_12841);
xnor U13408 (N_13408,N_12576,N_12903);
or U13409 (N_13409,N_12638,N_12934);
nand U13410 (N_13410,N_12695,N_12712);
or U13411 (N_13411,N_12923,N_12603);
or U13412 (N_13412,N_12852,N_12687);
nor U13413 (N_13413,N_12546,N_12759);
xor U13414 (N_13414,N_12955,N_12960);
nor U13415 (N_13415,N_12824,N_12927);
xor U13416 (N_13416,N_12567,N_12792);
and U13417 (N_13417,N_12538,N_12630);
nor U13418 (N_13418,N_12596,N_12955);
nand U13419 (N_13419,N_12579,N_12637);
nor U13420 (N_13420,N_12773,N_12566);
nand U13421 (N_13421,N_12677,N_12669);
nor U13422 (N_13422,N_12815,N_12943);
or U13423 (N_13423,N_12764,N_12965);
xor U13424 (N_13424,N_12622,N_12501);
or U13425 (N_13425,N_12982,N_12887);
xor U13426 (N_13426,N_12914,N_12653);
nor U13427 (N_13427,N_12855,N_12573);
and U13428 (N_13428,N_12620,N_12806);
nor U13429 (N_13429,N_12597,N_12518);
xnor U13430 (N_13430,N_12612,N_12939);
nand U13431 (N_13431,N_12937,N_12914);
nor U13432 (N_13432,N_12814,N_12588);
xnor U13433 (N_13433,N_12713,N_12725);
or U13434 (N_13434,N_12689,N_12673);
nand U13435 (N_13435,N_12894,N_12748);
and U13436 (N_13436,N_12740,N_12557);
nor U13437 (N_13437,N_12592,N_12868);
or U13438 (N_13438,N_12722,N_12926);
nor U13439 (N_13439,N_12503,N_12676);
nand U13440 (N_13440,N_12815,N_12762);
xor U13441 (N_13441,N_12729,N_12802);
nand U13442 (N_13442,N_12962,N_12772);
xnor U13443 (N_13443,N_12717,N_12769);
xnor U13444 (N_13444,N_12595,N_12836);
nand U13445 (N_13445,N_12648,N_12973);
and U13446 (N_13446,N_12650,N_12526);
or U13447 (N_13447,N_12794,N_12867);
or U13448 (N_13448,N_12796,N_12837);
nor U13449 (N_13449,N_12912,N_12764);
or U13450 (N_13450,N_12898,N_12808);
and U13451 (N_13451,N_12908,N_12941);
nand U13452 (N_13452,N_12626,N_12930);
nor U13453 (N_13453,N_12789,N_12920);
and U13454 (N_13454,N_12927,N_12706);
and U13455 (N_13455,N_12598,N_12735);
xor U13456 (N_13456,N_12852,N_12531);
nor U13457 (N_13457,N_12720,N_12916);
or U13458 (N_13458,N_12513,N_12899);
nor U13459 (N_13459,N_12790,N_12513);
nand U13460 (N_13460,N_12514,N_12684);
nand U13461 (N_13461,N_12744,N_12978);
nor U13462 (N_13462,N_12713,N_12853);
or U13463 (N_13463,N_12813,N_12964);
nand U13464 (N_13464,N_12786,N_12830);
or U13465 (N_13465,N_12631,N_12844);
and U13466 (N_13466,N_12946,N_12878);
xnor U13467 (N_13467,N_12574,N_12591);
xnor U13468 (N_13468,N_12808,N_12856);
or U13469 (N_13469,N_12572,N_12680);
xnor U13470 (N_13470,N_12547,N_12696);
nor U13471 (N_13471,N_12977,N_12792);
nor U13472 (N_13472,N_12904,N_12828);
and U13473 (N_13473,N_12534,N_12543);
or U13474 (N_13474,N_12676,N_12811);
xnor U13475 (N_13475,N_12679,N_12796);
nand U13476 (N_13476,N_12739,N_12875);
or U13477 (N_13477,N_12697,N_12837);
nand U13478 (N_13478,N_12981,N_12950);
or U13479 (N_13479,N_12525,N_12666);
and U13480 (N_13480,N_12617,N_12971);
nor U13481 (N_13481,N_12558,N_12551);
and U13482 (N_13482,N_12910,N_12715);
xnor U13483 (N_13483,N_12750,N_12582);
nand U13484 (N_13484,N_12760,N_12854);
and U13485 (N_13485,N_12764,N_12851);
or U13486 (N_13486,N_12868,N_12793);
and U13487 (N_13487,N_12909,N_12565);
nand U13488 (N_13488,N_12840,N_12953);
and U13489 (N_13489,N_12931,N_12582);
or U13490 (N_13490,N_12822,N_12596);
and U13491 (N_13491,N_12836,N_12523);
and U13492 (N_13492,N_12790,N_12763);
or U13493 (N_13493,N_12504,N_12738);
and U13494 (N_13494,N_12544,N_12923);
xnor U13495 (N_13495,N_12957,N_12913);
xor U13496 (N_13496,N_12848,N_12688);
or U13497 (N_13497,N_12589,N_12846);
nor U13498 (N_13498,N_12635,N_12973);
nor U13499 (N_13499,N_12705,N_12583);
nor U13500 (N_13500,N_13388,N_13219);
or U13501 (N_13501,N_13181,N_13302);
nor U13502 (N_13502,N_13487,N_13089);
or U13503 (N_13503,N_13150,N_13298);
or U13504 (N_13504,N_13254,N_13083);
or U13505 (N_13505,N_13060,N_13224);
nor U13506 (N_13506,N_13095,N_13435);
and U13507 (N_13507,N_13253,N_13395);
or U13508 (N_13508,N_13015,N_13047);
xnor U13509 (N_13509,N_13304,N_13188);
or U13510 (N_13510,N_13292,N_13202);
nand U13511 (N_13511,N_13094,N_13494);
nor U13512 (N_13512,N_13495,N_13081);
or U13513 (N_13513,N_13330,N_13403);
xnor U13514 (N_13514,N_13082,N_13427);
nor U13515 (N_13515,N_13469,N_13258);
and U13516 (N_13516,N_13165,N_13305);
xnor U13517 (N_13517,N_13438,N_13448);
and U13518 (N_13518,N_13325,N_13420);
xor U13519 (N_13519,N_13274,N_13499);
nand U13520 (N_13520,N_13361,N_13363);
nor U13521 (N_13521,N_13024,N_13451);
and U13522 (N_13522,N_13116,N_13446);
nand U13523 (N_13523,N_13185,N_13239);
and U13524 (N_13524,N_13107,N_13008);
nand U13525 (N_13525,N_13322,N_13108);
and U13526 (N_13526,N_13231,N_13402);
xnor U13527 (N_13527,N_13085,N_13168);
xnor U13528 (N_13528,N_13382,N_13467);
and U13529 (N_13529,N_13009,N_13485);
and U13530 (N_13530,N_13232,N_13179);
xnor U13531 (N_13531,N_13244,N_13104);
and U13532 (N_13532,N_13412,N_13425);
nor U13533 (N_13533,N_13045,N_13040);
xor U13534 (N_13534,N_13048,N_13352);
nand U13535 (N_13535,N_13262,N_13068);
and U13536 (N_13536,N_13197,N_13221);
nor U13537 (N_13537,N_13404,N_13041);
and U13538 (N_13538,N_13250,N_13144);
xnor U13539 (N_13539,N_13006,N_13398);
nand U13540 (N_13540,N_13037,N_13337);
and U13541 (N_13541,N_13242,N_13209);
nand U13542 (N_13542,N_13272,N_13328);
nor U13543 (N_13543,N_13090,N_13285);
xor U13544 (N_13544,N_13025,N_13183);
or U13545 (N_13545,N_13133,N_13236);
nand U13546 (N_13546,N_13259,N_13155);
or U13547 (N_13547,N_13129,N_13443);
or U13548 (N_13548,N_13028,N_13369);
xor U13549 (N_13549,N_13473,N_13338);
nor U13550 (N_13550,N_13163,N_13249);
xor U13551 (N_13551,N_13289,N_13329);
or U13552 (N_13552,N_13201,N_13158);
and U13553 (N_13553,N_13211,N_13429);
xor U13554 (N_13554,N_13383,N_13479);
nor U13555 (N_13555,N_13314,N_13145);
xor U13556 (N_13556,N_13489,N_13303);
xor U13557 (N_13557,N_13324,N_13235);
nand U13558 (N_13558,N_13036,N_13121);
and U13559 (N_13559,N_13125,N_13152);
nor U13560 (N_13560,N_13416,N_13445);
and U13561 (N_13561,N_13111,N_13349);
nand U13562 (N_13562,N_13205,N_13021);
nand U13563 (N_13563,N_13423,N_13441);
or U13564 (N_13564,N_13186,N_13140);
nand U13565 (N_13565,N_13280,N_13268);
nor U13566 (N_13566,N_13342,N_13424);
xor U13567 (N_13567,N_13460,N_13273);
and U13568 (N_13568,N_13167,N_13478);
and U13569 (N_13569,N_13379,N_13012);
nand U13570 (N_13570,N_13044,N_13000);
xnor U13571 (N_13571,N_13295,N_13252);
or U13572 (N_13572,N_13360,N_13245);
or U13573 (N_13573,N_13112,N_13365);
and U13574 (N_13574,N_13137,N_13464);
xnor U13575 (N_13575,N_13411,N_13146);
nand U13576 (N_13576,N_13456,N_13477);
and U13577 (N_13577,N_13226,N_13332);
nand U13578 (N_13578,N_13043,N_13059);
nor U13579 (N_13579,N_13476,N_13393);
or U13580 (N_13580,N_13340,N_13434);
xor U13581 (N_13581,N_13051,N_13153);
nand U13582 (N_13582,N_13005,N_13046);
xnor U13583 (N_13583,N_13141,N_13031);
or U13584 (N_13584,N_13066,N_13331);
nor U13585 (N_13585,N_13091,N_13011);
nor U13586 (N_13586,N_13099,N_13058);
xor U13587 (N_13587,N_13269,N_13010);
and U13588 (N_13588,N_13171,N_13243);
xnor U13589 (N_13589,N_13463,N_13333);
nand U13590 (N_13590,N_13439,N_13161);
nor U13591 (N_13591,N_13247,N_13394);
xnor U13592 (N_13592,N_13049,N_13222);
or U13593 (N_13593,N_13013,N_13070);
or U13594 (N_13594,N_13400,N_13054);
and U13595 (N_13595,N_13454,N_13364);
nand U13596 (N_13596,N_13182,N_13026);
nor U13597 (N_13597,N_13149,N_13173);
or U13598 (N_13598,N_13255,N_13038);
xor U13599 (N_13599,N_13312,N_13447);
nor U13600 (N_13600,N_13359,N_13297);
and U13601 (N_13601,N_13271,N_13452);
nor U13602 (N_13602,N_13080,N_13263);
xor U13603 (N_13603,N_13466,N_13376);
nand U13604 (N_13604,N_13296,N_13117);
or U13605 (N_13605,N_13288,N_13234);
or U13606 (N_13606,N_13122,N_13350);
nand U13607 (N_13607,N_13213,N_13284);
or U13608 (N_13608,N_13367,N_13334);
nand U13609 (N_13609,N_13097,N_13490);
and U13610 (N_13610,N_13033,N_13374);
nor U13611 (N_13611,N_13283,N_13237);
or U13612 (N_13612,N_13159,N_13194);
and U13613 (N_13613,N_13053,N_13124);
xor U13614 (N_13614,N_13310,N_13355);
or U13615 (N_13615,N_13214,N_13264);
nand U13616 (N_13616,N_13078,N_13462);
or U13617 (N_13617,N_13136,N_13093);
nor U13618 (N_13618,N_13131,N_13381);
nand U13619 (N_13619,N_13087,N_13135);
nor U13620 (N_13620,N_13301,N_13413);
and U13621 (N_13621,N_13279,N_13132);
xor U13622 (N_13622,N_13321,N_13278);
or U13623 (N_13623,N_13386,N_13139);
xnor U13624 (N_13624,N_13248,N_13019);
nor U13625 (N_13625,N_13414,N_13436);
xnor U13626 (N_13626,N_13323,N_13127);
and U13627 (N_13627,N_13126,N_13007);
nor U13628 (N_13628,N_13343,N_13071);
xor U13629 (N_13629,N_13105,N_13061);
and U13630 (N_13630,N_13375,N_13428);
xnor U13631 (N_13631,N_13461,N_13014);
and U13632 (N_13632,N_13029,N_13092);
nor U13633 (N_13633,N_13180,N_13335);
nand U13634 (N_13634,N_13432,N_13178);
nand U13635 (N_13635,N_13472,N_13246);
or U13636 (N_13636,N_13317,N_13098);
nor U13637 (N_13637,N_13372,N_13327);
and U13638 (N_13638,N_13184,N_13415);
xor U13639 (N_13639,N_13294,N_13120);
nor U13640 (N_13640,N_13308,N_13187);
xor U13641 (N_13641,N_13370,N_13318);
and U13642 (N_13642,N_13486,N_13172);
nor U13643 (N_13643,N_13399,N_13326);
nand U13644 (N_13644,N_13204,N_13260);
xnor U13645 (N_13645,N_13138,N_13151);
or U13646 (N_13646,N_13063,N_13039);
nand U13647 (N_13647,N_13371,N_13032);
and U13648 (N_13648,N_13164,N_13227);
nor U13649 (N_13649,N_13421,N_13437);
nand U13650 (N_13650,N_13101,N_13482);
nor U13651 (N_13651,N_13341,N_13459);
nor U13652 (N_13652,N_13366,N_13348);
and U13653 (N_13653,N_13387,N_13241);
nand U13654 (N_13654,N_13450,N_13346);
or U13655 (N_13655,N_13162,N_13453);
and U13656 (N_13656,N_13190,N_13076);
or U13657 (N_13657,N_13405,N_13240);
nor U13658 (N_13658,N_13391,N_13203);
and U13659 (N_13659,N_13483,N_13390);
or U13660 (N_13660,N_13238,N_13073);
nand U13661 (N_13661,N_13215,N_13216);
or U13662 (N_13662,N_13431,N_13481);
nand U13663 (N_13663,N_13113,N_13493);
nor U13664 (N_13664,N_13142,N_13079);
nand U13665 (N_13665,N_13444,N_13052);
and U13666 (N_13666,N_13470,N_13336);
xor U13667 (N_13667,N_13380,N_13075);
nor U13668 (N_13668,N_13373,N_13267);
nor U13669 (N_13669,N_13115,N_13480);
and U13670 (N_13670,N_13384,N_13358);
or U13671 (N_13671,N_13488,N_13293);
nor U13672 (N_13672,N_13418,N_13458);
and U13673 (N_13673,N_13315,N_13103);
or U13674 (N_13674,N_13407,N_13287);
or U13675 (N_13675,N_13134,N_13004);
and U13676 (N_13676,N_13277,N_13106);
nand U13677 (N_13677,N_13016,N_13195);
or U13678 (N_13678,N_13177,N_13147);
nor U13679 (N_13679,N_13062,N_13286);
nand U13680 (N_13680,N_13497,N_13491);
nand U13681 (N_13681,N_13422,N_13110);
or U13682 (N_13682,N_13055,N_13148);
and U13683 (N_13683,N_13406,N_13256);
nor U13684 (N_13684,N_13154,N_13389);
and U13685 (N_13685,N_13449,N_13492);
and U13686 (N_13686,N_13199,N_13198);
and U13687 (N_13687,N_13397,N_13409);
and U13688 (N_13688,N_13291,N_13313);
or U13689 (N_13689,N_13096,N_13193);
nor U13690 (N_13690,N_13316,N_13030);
nor U13691 (N_13691,N_13210,N_13022);
nand U13692 (N_13692,N_13498,N_13086);
xnor U13693 (N_13693,N_13212,N_13067);
xor U13694 (N_13694,N_13118,N_13396);
nor U13695 (N_13695,N_13484,N_13109);
xor U13696 (N_13696,N_13306,N_13378);
or U13697 (N_13697,N_13282,N_13192);
and U13698 (N_13698,N_13206,N_13351);
or U13699 (N_13699,N_13169,N_13339);
and U13700 (N_13700,N_13344,N_13225);
xor U13701 (N_13701,N_13002,N_13440);
and U13702 (N_13702,N_13320,N_13156);
and U13703 (N_13703,N_13077,N_13228);
nand U13704 (N_13704,N_13057,N_13207);
xor U13705 (N_13705,N_13417,N_13354);
xor U13706 (N_13706,N_13196,N_13307);
xnor U13707 (N_13707,N_13275,N_13299);
xnor U13708 (N_13708,N_13347,N_13257);
nand U13709 (N_13709,N_13074,N_13276);
nand U13710 (N_13710,N_13065,N_13233);
xor U13711 (N_13711,N_13281,N_13377);
xor U13712 (N_13712,N_13023,N_13468);
xor U13713 (N_13713,N_13408,N_13119);
nand U13714 (N_13714,N_13084,N_13189);
nor U13715 (N_13715,N_13392,N_13200);
and U13716 (N_13716,N_13017,N_13166);
or U13717 (N_13717,N_13319,N_13170);
nand U13718 (N_13718,N_13300,N_13102);
nor U13719 (N_13719,N_13191,N_13069);
and U13720 (N_13720,N_13160,N_13474);
and U13721 (N_13721,N_13130,N_13442);
nand U13722 (N_13722,N_13027,N_13353);
or U13723 (N_13723,N_13128,N_13035);
or U13724 (N_13724,N_13100,N_13266);
nand U13725 (N_13725,N_13229,N_13496);
or U13726 (N_13726,N_13174,N_13143);
xor U13727 (N_13727,N_13356,N_13311);
nor U13728 (N_13728,N_13457,N_13003);
nand U13729 (N_13729,N_13218,N_13220);
and U13730 (N_13730,N_13455,N_13042);
or U13731 (N_13731,N_13018,N_13433);
or U13732 (N_13732,N_13001,N_13072);
xor U13733 (N_13733,N_13419,N_13251);
or U13734 (N_13734,N_13471,N_13357);
nand U13735 (N_13735,N_13064,N_13401);
or U13736 (N_13736,N_13020,N_13345);
and U13737 (N_13737,N_13426,N_13223);
or U13738 (N_13738,N_13034,N_13362);
nor U13739 (N_13739,N_13088,N_13230);
or U13740 (N_13740,N_13114,N_13157);
xnor U13741 (N_13741,N_13410,N_13056);
nand U13742 (N_13742,N_13430,N_13123);
nor U13743 (N_13743,N_13465,N_13385);
nor U13744 (N_13744,N_13050,N_13270);
and U13745 (N_13745,N_13265,N_13475);
nand U13746 (N_13746,N_13261,N_13217);
and U13747 (N_13747,N_13368,N_13176);
and U13748 (N_13748,N_13309,N_13175);
nor U13749 (N_13749,N_13208,N_13290);
and U13750 (N_13750,N_13038,N_13370);
or U13751 (N_13751,N_13426,N_13210);
and U13752 (N_13752,N_13015,N_13430);
nand U13753 (N_13753,N_13275,N_13323);
or U13754 (N_13754,N_13296,N_13010);
xor U13755 (N_13755,N_13466,N_13430);
and U13756 (N_13756,N_13398,N_13137);
and U13757 (N_13757,N_13269,N_13012);
and U13758 (N_13758,N_13054,N_13121);
nor U13759 (N_13759,N_13463,N_13155);
xnor U13760 (N_13760,N_13335,N_13192);
nand U13761 (N_13761,N_13473,N_13064);
or U13762 (N_13762,N_13418,N_13159);
or U13763 (N_13763,N_13493,N_13253);
nor U13764 (N_13764,N_13184,N_13114);
nor U13765 (N_13765,N_13202,N_13413);
nand U13766 (N_13766,N_13035,N_13029);
or U13767 (N_13767,N_13396,N_13027);
xnor U13768 (N_13768,N_13378,N_13162);
and U13769 (N_13769,N_13111,N_13239);
nor U13770 (N_13770,N_13250,N_13098);
nor U13771 (N_13771,N_13497,N_13311);
nand U13772 (N_13772,N_13426,N_13017);
nand U13773 (N_13773,N_13124,N_13350);
nor U13774 (N_13774,N_13045,N_13152);
xnor U13775 (N_13775,N_13281,N_13405);
and U13776 (N_13776,N_13195,N_13159);
xor U13777 (N_13777,N_13028,N_13399);
and U13778 (N_13778,N_13014,N_13197);
and U13779 (N_13779,N_13114,N_13468);
and U13780 (N_13780,N_13442,N_13063);
and U13781 (N_13781,N_13350,N_13245);
nor U13782 (N_13782,N_13499,N_13481);
and U13783 (N_13783,N_13050,N_13480);
and U13784 (N_13784,N_13043,N_13039);
nor U13785 (N_13785,N_13401,N_13316);
nand U13786 (N_13786,N_13033,N_13158);
nor U13787 (N_13787,N_13429,N_13158);
xnor U13788 (N_13788,N_13372,N_13369);
or U13789 (N_13789,N_13387,N_13161);
and U13790 (N_13790,N_13489,N_13146);
and U13791 (N_13791,N_13384,N_13359);
xor U13792 (N_13792,N_13097,N_13335);
and U13793 (N_13793,N_13143,N_13478);
xor U13794 (N_13794,N_13050,N_13379);
nand U13795 (N_13795,N_13395,N_13293);
nor U13796 (N_13796,N_13164,N_13093);
nor U13797 (N_13797,N_13371,N_13028);
and U13798 (N_13798,N_13052,N_13474);
nand U13799 (N_13799,N_13243,N_13300);
xnor U13800 (N_13800,N_13217,N_13271);
xor U13801 (N_13801,N_13456,N_13062);
or U13802 (N_13802,N_13306,N_13232);
nor U13803 (N_13803,N_13201,N_13439);
xor U13804 (N_13804,N_13031,N_13115);
nand U13805 (N_13805,N_13402,N_13029);
nand U13806 (N_13806,N_13202,N_13124);
or U13807 (N_13807,N_13024,N_13023);
or U13808 (N_13808,N_13498,N_13352);
nor U13809 (N_13809,N_13070,N_13241);
nor U13810 (N_13810,N_13393,N_13499);
or U13811 (N_13811,N_13197,N_13422);
nor U13812 (N_13812,N_13087,N_13371);
nand U13813 (N_13813,N_13165,N_13186);
or U13814 (N_13814,N_13161,N_13269);
xor U13815 (N_13815,N_13360,N_13257);
and U13816 (N_13816,N_13040,N_13454);
and U13817 (N_13817,N_13477,N_13308);
nand U13818 (N_13818,N_13098,N_13299);
nand U13819 (N_13819,N_13341,N_13497);
nor U13820 (N_13820,N_13055,N_13255);
nor U13821 (N_13821,N_13277,N_13464);
or U13822 (N_13822,N_13294,N_13110);
and U13823 (N_13823,N_13175,N_13440);
nand U13824 (N_13824,N_13103,N_13353);
nand U13825 (N_13825,N_13230,N_13118);
xor U13826 (N_13826,N_13003,N_13428);
or U13827 (N_13827,N_13347,N_13165);
or U13828 (N_13828,N_13479,N_13010);
and U13829 (N_13829,N_13094,N_13211);
nor U13830 (N_13830,N_13349,N_13324);
nand U13831 (N_13831,N_13260,N_13061);
xnor U13832 (N_13832,N_13383,N_13139);
nor U13833 (N_13833,N_13410,N_13161);
nand U13834 (N_13834,N_13439,N_13303);
or U13835 (N_13835,N_13306,N_13271);
xor U13836 (N_13836,N_13078,N_13032);
nand U13837 (N_13837,N_13005,N_13421);
nand U13838 (N_13838,N_13122,N_13335);
or U13839 (N_13839,N_13498,N_13188);
nand U13840 (N_13840,N_13364,N_13300);
nor U13841 (N_13841,N_13139,N_13289);
xnor U13842 (N_13842,N_13439,N_13053);
xnor U13843 (N_13843,N_13331,N_13278);
nand U13844 (N_13844,N_13362,N_13088);
nand U13845 (N_13845,N_13159,N_13229);
and U13846 (N_13846,N_13163,N_13196);
nand U13847 (N_13847,N_13383,N_13475);
nand U13848 (N_13848,N_13424,N_13406);
nor U13849 (N_13849,N_13083,N_13221);
and U13850 (N_13850,N_13204,N_13219);
or U13851 (N_13851,N_13302,N_13439);
or U13852 (N_13852,N_13163,N_13262);
nand U13853 (N_13853,N_13461,N_13011);
nor U13854 (N_13854,N_13164,N_13221);
and U13855 (N_13855,N_13093,N_13412);
or U13856 (N_13856,N_13472,N_13456);
xor U13857 (N_13857,N_13206,N_13232);
xnor U13858 (N_13858,N_13224,N_13208);
xor U13859 (N_13859,N_13263,N_13171);
and U13860 (N_13860,N_13116,N_13102);
or U13861 (N_13861,N_13009,N_13358);
nand U13862 (N_13862,N_13380,N_13390);
xnor U13863 (N_13863,N_13349,N_13278);
xor U13864 (N_13864,N_13099,N_13019);
nand U13865 (N_13865,N_13499,N_13208);
and U13866 (N_13866,N_13029,N_13245);
or U13867 (N_13867,N_13225,N_13450);
and U13868 (N_13868,N_13016,N_13349);
nand U13869 (N_13869,N_13487,N_13485);
or U13870 (N_13870,N_13235,N_13281);
nand U13871 (N_13871,N_13003,N_13291);
xor U13872 (N_13872,N_13375,N_13455);
nor U13873 (N_13873,N_13186,N_13092);
or U13874 (N_13874,N_13388,N_13197);
or U13875 (N_13875,N_13302,N_13005);
nand U13876 (N_13876,N_13249,N_13067);
xnor U13877 (N_13877,N_13118,N_13241);
or U13878 (N_13878,N_13070,N_13285);
nand U13879 (N_13879,N_13048,N_13231);
nand U13880 (N_13880,N_13285,N_13407);
nor U13881 (N_13881,N_13112,N_13382);
nand U13882 (N_13882,N_13426,N_13152);
nand U13883 (N_13883,N_13478,N_13292);
xnor U13884 (N_13884,N_13054,N_13411);
or U13885 (N_13885,N_13049,N_13052);
or U13886 (N_13886,N_13253,N_13372);
nor U13887 (N_13887,N_13100,N_13310);
nor U13888 (N_13888,N_13492,N_13092);
nor U13889 (N_13889,N_13246,N_13358);
xor U13890 (N_13890,N_13134,N_13025);
and U13891 (N_13891,N_13373,N_13032);
xnor U13892 (N_13892,N_13450,N_13386);
and U13893 (N_13893,N_13024,N_13040);
or U13894 (N_13894,N_13312,N_13010);
xnor U13895 (N_13895,N_13191,N_13143);
and U13896 (N_13896,N_13413,N_13135);
nand U13897 (N_13897,N_13370,N_13067);
and U13898 (N_13898,N_13176,N_13094);
or U13899 (N_13899,N_13099,N_13330);
nand U13900 (N_13900,N_13398,N_13112);
nor U13901 (N_13901,N_13229,N_13413);
and U13902 (N_13902,N_13420,N_13423);
and U13903 (N_13903,N_13110,N_13343);
nor U13904 (N_13904,N_13029,N_13319);
nand U13905 (N_13905,N_13462,N_13197);
or U13906 (N_13906,N_13036,N_13103);
and U13907 (N_13907,N_13280,N_13459);
and U13908 (N_13908,N_13440,N_13266);
and U13909 (N_13909,N_13110,N_13290);
or U13910 (N_13910,N_13259,N_13046);
and U13911 (N_13911,N_13153,N_13249);
xnor U13912 (N_13912,N_13194,N_13489);
nor U13913 (N_13913,N_13385,N_13464);
nor U13914 (N_13914,N_13373,N_13183);
or U13915 (N_13915,N_13256,N_13009);
xor U13916 (N_13916,N_13356,N_13070);
or U13917 (N_13917,N_13210,N_13447);
or U13918 (N_13918,N_13280,N_13151);
nand U13919 (N_13919,N_13004,N_13294);
xnor U13920 (N_13920,N_13273,N_13432);
nor U13921 (N_13921,N_13158,N_13422);
xor U13922 (N_13922,N_13427,N_13462);
nand U13923 (N_13923,N_13151,N_13335);
xor U13924 (N_13924,N_13459,N_13026);
nor U13925 (N_13925,N_13197,N_13468);
or U13926 (N_13926,N_13411,N_13393);
nand U13927 (N_13927,N_13316,N_13414);
and U13928 (N_13928,N_13034,N_13051);
xor U13929 (N_13929,N_13259,N_13060);
or U13930 (N_13930,N_13154,N_13302);
nor U13931 (N_13931,N_13188,N_13419);
nor U13932 (N_13932,N_13297,N_13248);
xnor U13933 (N_13933,N_13121,N_13269);
xor U13934 (N_13934,N_13438,N_13012);
nand U13935 (N_13935,N_13462,N_13072);
nand U13936 (N_13936,N_13103,N_13435);
or U13937 (N_13937,N_13436,N_13359);
and U13938 (N_13938,N_13068,N_13272);
or U13939 (N_13939,N_13496,N_13242);
nor U13940 (N_13940,N_13299,N_13023);
or U13941 (N_13941,N_13107,N_13295);
and U13942 (N_13942,N_13399,N_13226);
nor U13943 (N_13943,N_13236,N_13060);
or U13944 (N_13944,N_13167,N_13418);
nand U13945 (N_13945,N_13028,N_13088);
nor U13946 (N_13946,N_13368,N_13156);
xor U13947 (N_13947,N_13441,N_13199);
and U13948 (N_13948,N_13123,N_13091);
or U13949 (N_13949,N_13236,N_13258);
xor U13950 (N_13950,N_13477,N_13128);
nand U13951 (N_13951,N_13423,N_13101);
and U13952 (N_13952,N_13205,N_13499);
nor U13953 (N_13953,N_13165,N_13467);
or U13954 (N_13954,N_13117,N_13494);
xnor U13955 (N_13955,N_13230,N_13418);
nor U13956 (N_13956,N_13452,N_13281);
nor U13957 (N_13957,N_13342,N_13234);
xnor U13958 (N_13958,N_13191,N_13247);
and U13959 (N_13959,N_13129,N_13338);
xor U13960 (N_13960,N_13077,N_13355);
nand U13961 (N_13961,N_13282,N_13190);
or U13962 (N_13962,N_13135,N_13168);
xor U13963 (N_13963,N_13131,N_13198);
and U13964 (N_13964,N_13307,N_13397);
or U13965 (N_13965,N_13203,N_13345);
or U13966 (N_13966,N_13020,N_13267);
nor U13967 (N_13967,N_13053,N_13028);
and U13968 (N_13968,N_13056,N_13017);
or U13969 (N_13969,N_13206,N_13166);
and U13970 (N_13970,N_13063,N_13201);
nor U13971 (N_13971,N_13112,N_13303);
nand U13972 (N_13972,N_13357,N_13216);
nand U13973 (N_13973,N_13265,N_13395);
or U13974 (N_13974,N_13414,N_13409);
and U13975 (N_13975,N_13392,N_13485);
xor U13976 (N_13976,N_13476,N_13030);
nand U13977 (N_13977,N_13082,N_13360);
nand U13978 (N_13978,N_13385,N_13135);
nand U13979 (N_13979,N_13289,N_13413);
and U13980 (N_13980,N_13413,N_13196);
xor U13981 (N_13981,N_13180,N_13266);
nor U13982 (N_13982,N_13131,N_13269);
and U13983 (N_13983,N_13293,N_13177);
or U13984 (N_13984,N_13066,N_13393);
and U13985 (N_13985,N_13025,N_13447);
and U13986 (N_13986,N_13006,N_13216);
nand U13987 (N_13987,N_13039,N_13317);
nand U13988 (N_13988,N_13420,N_13161);
nor U13989 (N_13989,N_13265,N_13132);
and U13990 (N_13990,N_13196,N_13229);
nor U13991 (N_13991,N_13339,N_13232);
nand U13992 (N_13992,N_13389,N_13324);
nand U13993 (N_13993,N_13390,N_13371);
nor U13994 (N_13994,N_13280,N_13242);
and U13995 (N_13995,N_13352,N_13115);
nor U13996 (N_13996,N_13084,N_13396);
or U13997 (N_13997,N_13391,N_13446);
xnor U13998 (N_13998,N_13122,N_13478);
and U13999 (N_13999,N_13245,N_13183);
nand U14000 (N_14000,N_13505,N_13515);
or U14001 (N_14001,N_13606,N_13504);
nor U14002 (N_14002,N_13632,N_13751);
nor U14003 (N_14003,N_13781,N_13686);
nand U14004 (N_14004,N_13996,N_13784);
and U14005 (N_14005,N_13720,N_13862);
or U14006 (N_14006,N_13994,N_13818);
xor U14007 (N_14007,N_13611,N_13876);
and U14008 (N_14008,N_13870,N_13652);
xnor U14009 (N_14009,N_13900,N_13806);
and U14010 (N_14010,N_13835,N_13893);
and U14011 (N_14011,N_13620,N_13953);
nor U14012 (N_14012,N_13816,N_13526);
and U14013 (N_14013,N_13985,N_13624);
xor U14014 (N_14014,N_13634,N_13861);
or U14015 (N_14015,N_13901,N_13952);
nor U14016 (N_14016,N_13626,N_13650);
nor U14017 (N_14017,N_13666,N_13590);
or U14018 (N_14018,N_13548,N_13978);
or U14019 (N_14019,N_13792,N_13727);
nand U14020 (N_14020,N_13556,N_13763);
and U14021 (N_14021,N_13938,N_13575);
nand U14022 (N_14022,N_13932,N_13649);
nand U14023 (N_14023,N_13612,N_13857);
nand U14024 (N_14024,N_13529,N_13712);
and U14025 (N_14025,N_13676,N_13716);
nand U14026 (N_14026,N_13780,N_13608);
nand U14027 (N_14027,N_13790,N_13815);
nand U14028 (N_14028,N_13977,N_13694);
nor U14029 (N_14029,N_13885,N_13655);
and U14030 (N_14030,N_13629,N_13776);
or U14031 (N_14031,N_13638,N_13964);
nand U14032 (N_14032,N_13565,N_13843);
xor U14033 (N_14033,N_13558,N_13623);
xor U14034 (N_14034,N_13759,N_13966);
nor U14035 (N_14035,N_13967,N_13576);
nor U14036 (N_14036,N_13510,N_13588);
nand U14037 (N_14037,N_13808,N_13661);
xnor U14038 (N_14038,N_13890,N_13867);
xnor U14039 (N_14039,N_13521,N_13768);
or U14040 (N_14040,N_13602,N_13975);
or U14041 (N_14041,N_13577,N_13791);
xnor U14042 (N_14042,N_13704,N_13825);
nand U14043 (N_14043,N_13618,N_13936);
nor U14044 (N_14044,N_13884,N_13562);
nor U14045 (N_14045,N_13929,N_13918);
and U14046 (N_14046,N_13925,N_13758);
or U14047 (N_14047,N_13810,N_13860);
and U14048 (N_14048,N_13761,N_13729);
nand U14049 (N_14049,N_13696,N_13863);
nor U14050 (N_14050,N_13997,N_13789);
xnor U14051 (N_14051,N_13713,N_13923);
or U14052 (N_14052,N_13514,N_13689);
nor U14053 (N_14053,N_13728,N_13598);
nor U14054 (N_14054,N_13766,N_13697);
and U14055 (N_14055,N_13786,N_13663);
or U14056 (N_14056,N_13886,N_13995);
and U14057 (N_14057,N_13783,N_13841);
nand U14058 (N_14058,N_13855,N_13507);
and U14059 (N_14059,N_13594,N_13684);
nor U14060 (N_14060,N_13714,N_13685);
and U14061 (N_14061,N_13927,N_13669);
xnor U14062 (N_14062,N_13836,N_13633);
and U14063 (N_14063,N_13584,N_13693);
nor U14064 (N_14064,N_13683,N_13859);
and U14065 (N_14065,N_13957,N_13813);
xor U14066 (N_14066,N_13844,N_13769);
nand U14067 (N_14067,N_13544,N_13617);
or U14068 (N_14068,N_13847,N_13858);
or U14069 (N_14069,N_13738,N_13563);
xor U14070 (N_14070,N_13775,N_13948);
xor U14071 (N_14071,N_13681,N_13963);
xor U14072 (N_14072,N_13750,N_13910);
nor U14073 (N_14073,N_13917,N_13960);
and U14074 (N_14074,N_13915,N_13873);
nand U14075 (N_14075,N_13880,N_13959);
and U14076 (N_14076,N_13962,N_13842);
nor U14077 (N_14077,N_13907,N_13670);
nand U14078 (N_14078,N_13903,N_13587);
nor U14079 (N_14079,N_13930,N_13990);
and U14080 (N_14080,N_13767,N_13567);
or U14081 (N_14081,N_13703,N_13673);
nor U14082 (N_14082,N_13688,N_13945);
xnor U14083 (N_14083,N_13969,N_13840);
nor U14084 (N_14084,N_13586,N_13531);
and U14085 (N_14085,N_13949,N_13872);
xor U14086 (N_14086,N_13664,N_13811);
and U14087 (N_14087,N_13545,N_13849);
or U14088 (N_14088,N_13668,N_13739);
nand U14089 (N_14089,N_13896,N_13679);
nand U14090 (N_14090,N_13943,N_13797);
nor U14091 (N_14091,N_13935,N_13740);
nor U14092 (N_14092,N_13541,N_13782);
and U14093 (N_14093,N_13830,N_13603);
xor U14094 (N_14094,N_13534,N_13610);
nand U14095 (N_14095,N_13804,N_13939);
or U14096 (N_14096,N_13581,N_13640);
and U14097 (N_14097,N_13875,N_13878);
or U14098 (N_14098,N_13674,N_13513);
xor U14099 (N_14099,N_13799,N_13956);
nand U14100 (N_14100,N_13905,N_13546);
and U14101 (N_14101,N_13656,N_13627);
nand U14102 (N_14102,N_13998,N_13805);
nand U14103 (N_14103,N_13730,N_13735);
nor U14104 (N_14104,N_13942,N_13591);
nor U14105 (N_14105,N_13502,N_13981);
nand U14106 (N_14106,N_13695,N_13538);
nor U14107 (N_14107,N_13527,N_13865);
or U14108 (N_14108,N_13993,N_13573);
nor U14109 (N_14109,N_13746,N_13986);
and U14110 (N_14110,N_13654,N_13671);
xnor U14111 (N_14111,N_13785,N_13765);
nand U14112 (N_14112,N_13937,N_13748);
nand U14113 (N_14113,N_13651,N_13928);
nor U14114 (N_14114,N_13579,N_13913);
and U14115 (N_14115,N_13778,N_13642);
and U14116 (N_14116,N_13940,N_13823);
nor U14117 (N_14117,N_13822,N_13987);
xnor U14118 (N_14118,N_13757,N_13687);
nor U14119 (N_14119,N_13850,N_13523);
nand U14120 (N_14120,N_13906,N_13922);
nand U14121 (N_14121,N_13795,N_13657);
and U14122 (N_14122,N_13647,N_13547);
xor U14123 (N_14123,N_13803,N_13574);
xor U14124 (N_14124,N_13570,N_13801);
and U14125 (N_14125,N_13535,N_13691);
or U14126 (N_14126,N_13838,N_13934);
and U14127 (N_14127,N_13616,N_13516);
or U14128 (N_14128,N_13734,N_13800);
nor U14129 (N_14129,N_13724,N_13719);
nand U14130 (N_14130,N_13871,N_13503);
nand U14131 (N_14131,N_13889,N_13821);
or U14132 (N_14132,N_13709,N_13585);
xor U14133 (N_14133,N_13931,N_13530);
xor U14134 (N_14134,N_13607,N_13677);
xor U14135 (N_14135,N_13914,N_13852);
nand U14136 (N_14136,N_13895,N_13756);
and U14137 (N_14137,N_13974,N_13817);
xor U14138 (N_14138,N_13794,N_13777);
or U14139 (N_14139,N_13592,N_13736);
xor U14140 (N_14140,N_13643,N_13965);
nor U14141 (N_14141,N_13500,N_13899);
nand U14142 (N_14142,N_13645,N_13764);
xor U14143 (N_14143,N_13571,N_13846);
and U14144 (N_14144,N_13636,N_13774);
xnor U14145 (N_14145,N_13812,N_13733);
and U14146 (N_14146,N_13658,N_13798);
nand U14147 (N_14147,N_13628,N_13506);
xnor U14148 (N_14148,N_13509,N_13793);
or U14149 (N_14149,N_13557,N_13722);
xor U14150 (N_14150,N_13705,N_13542);
nand U14151 (N_14151,N_13824,N_13725);
nand U14152 (N_14152,N_13596,N_13770);
nor U14153 (N_14153,N_13980,N_13971);
xnor U14154 (N_14154,N_13522,N_13864);
nand U14155 (N_14155,N_13702,N_13622);
nand U14156 (N_14156,N_13991,N_13891);
and U14157 (N_14157,N_13779,N_13583);
xor U14158 (N_14158,N_13614,N_13726);
or U14159 (N_14159,N_13692,N_13667);
nor U14160 (N_14160,N_13662,N_13552);
or U14161 (N_14161,N_13946,N_13630);
or U14162 (N_14162,N_13600,N_13992);
nor U14163 (N_14163,N_13827,N_13517);
nor U14164 (N_14164,N_13831,N_13731);
nand U14165 (N_14165,N_13680,N_13635);
or U14166 (N_14166,N_13648,N_13659);
and U14167 (N_14167,N_13951,N_13569);
and U14168 (N_14168,N_13868,N_13839);
xor U14169 (N_14169,N_13837,N_13999);
nand U14170 (N_14170,N_13958,N_13723);
or U14171 (N_14171,N_13989,N_13787);
nor U14172 (N_14172,N_13621,N_13845);
xor U14173 (N_14173,N_13721,N_13988);
nor U14174 (N_14174,N_13856,N_13568);
or U14175 (N_14175,N_13718,N_13737);
or U14176 (N_14176,N_13888,N_13754);
and U14177 (N_14177,N_13540,N_13698);
xnor U14178 (N_14178,N_13897,N_13747);
nor U14179 (N_14179,N_13894,N_13706);
xnor U14180 (N_14180,N_13566,N_13834);
or U14181 (N_14181,N_13543,N_13707);
nand U14182 (N_14182,N_13933,N_13973);
or U14183 (N_14183,N_13771,N_13788);
or U14184 (N_14184,N_13954,N_13532);
nor U14185 (N_14185,N_13605,N_13537);
or U14186 (N_14186,N_13699,N_13807);
and U14187 (N_14187,N_13520,N_13604);
xor U14188 (N_14188,N_13809,N_13550);
xor U14189 (N_14189,N_13715,N_13961);
and U14190 (N_14190,N_13637,N_13753);
and U14191 (N_14191,N_13911,N_13814);
nor U14192 (N_14192,N_13665,N_13660);
xnor U14193 (N_14193,N_13882,N_13613);
or U14194 (N_14194,N_13902,N_13559);
nor U14195 (N_14195,N_13518,N_13755);
nand U14196 (N_14196,N_13732,N_13682);
or U14197 (N_14197,N_13549,N_13773);
or U14198 (N_14198,N_13625,N_13982);
nand U14199 (N_14199,N_13820,N_13599);
nor U14200 (N_14200,N_13920,N_13832);
nand U14201 (N_14201,N_13833,N_13701);
or U14202 (N_14202,N_13597,N_13877);
nand U14203 (N_14203,N_13672,N_13589);
and U14204 (N_14204,N_13887,N_13869);
xnor U14205 (N_14205,N_13560,N_13879);
nor U14206 (N_14206,N_13826,N_13554);
or U14207 (N_14207,N_13580,N_13950);
nor U14208 (N_14208,N_13519,N_13508);
or U14209 (N_14209,N_13743,N_13898);
nor U14210 (N_14210,N_13926,N_13572);
and U14211 (N_14211,N_13646,N_13916);
nand U14212 (N_14212,N_13912,N_13919);
xor U14213 (N_14213,N_13710,N_13536);
and U14214 (N_14214,N_13690,N_13595);
nor U14215 (N_14215,N_13524,N_13609);
nor U14216 (N_14216,N_13909,N_13553);
and U14217 (N_14217,N_13851,N_13979);
nor U14218 (N_14218,N_13874,N_13760);
and U14219 (N_14219,N_13802,N_13883);
xnor U14220 (N_14220,N_13854,N_13970);
nor U14221 (N_14221,N_13892,N_13976);
and U14222 (N_14222,N_13955,N_13908);
or U14223 (N_14223,N_13578,N_13752);
nor U14224 (N_14224,N_13866,N_13631);
and U14225 (N_14225,N_13564,N_13749);
nand U14226 (N_14226,N_13742,N_13528);
nand U14227 (N_14227,N_13848,N_13708);
xor U14228 (N_14228,N_13641,N_13921);
and U14229 (N_14229,N_13947,N_13711);
xor U14230 (N_14230,N_13762,N_13582);
or U14231 (N_14231,N_13853,N_13593);
nor U14232 (N_14232,N_13533,N_13512);
or U14233 (N_14233,N_13700,N_13675);
or U14234 (N_14234,N_13819,N_13619);
nor U14235 (N_14235,N_13601,N_13741);
nand U14236 (N_14236,N_13511,N_13717);
or U14237 (N_14237,N_13539,N_13904);
and U14238 (N_14238,N_13944,N_13678);
nand U14239 (N_14239,N_13551,N_13615);
nand U14240 (N_14240,N_13941,N_13555);
and U14241 (N_14241,N_13561,N_13653);
or U14242 (N_14242,N_13501,N_13829);
or U14243 (N_14243,N_13796,N_13984);
or U14244 (N_14244,N_13968,N_13744);
xnor U14245 (N_14245,N_13828,N_13881);
or U14246 (N_14246,N_13924,N_13745);
and U14247 (N_14247,N_13772,N_13972);
and U14248 (N_14248,N_13644,N_13639);
or U14249 (N_14249,N_13983,N_13525);
or U14250 (N_14250,N_13963,N_13727);
xor U14251 (N_14251,N_13528,N_13994);
or U14252 (N_14252,N_13522,N_13828);
nor U14253 (N_14253,N_13793,N_13526);
xnor U14254 (N_14254,N_13999,N_13867);
nor U14255 (N_14255,N_13545,N_13619);
xor U14256 (N_14256,N_13894,N_13508);
xnor U14257 (N_14257,N_13500,N_13943);
or U14258 (N_14258,N_13525,N_13559);
or U14259 (N_14259,N_13927,N_13511);
or U14260 (N_14260,N_13859,N_13802);
xor U14261 (N_14261,N_13505,N_13645);
and U14262 (N_14262,N_13759,N_13556);
and U14263 (N_14263,N_13606,N_13701);
and U14264 (N_14264,N_13810,N_13671);
xor U14265 (N_14265,N_13771,N_13630);
and U14266 (N_14266,N_13936,N_13731);
xor U14267 (N_14267,N_13851,N_13526);
or U14268 (N_14268,N_13564,N_13942);
and U14269 (N_14269,N_13842,N_13774);
nor U14270 (N_14270,N_13927,N_13607);
and U14271 (N_14271,N_13728,N_13507);
or U14272 (N_14272,N_13909,N_13933);
nand U14273 (N_14273,N_13819,N_13896);
nand U14274 (N_14274,N_13848,N_13554);
nand U14275 (N_14275,N_13901,N_13992);
and U14276 (N_14276,N_13692,N_13803);
or U14277 (N_14277,N_13649,N_13846);
nand U14278 (N_14278,N_13978,N_13864);
nor U14279 (N_14279,N_13661,N_13614);
or U14280 (N_14280,N_13569,N_13842);
or U14281 (N_14281,N_13966,N_13914);
or U14282 (N_14282,N_13741,N_13827);
nor U14283 (N_14283,N_13785,N_13871);
nand U14284 (N_14284,N_13713,N_13802);
and U14285 (N_14285,N_13686,N_13992);
or U14286 (N_14286,N_13692,N_13621);
nor U14287 (N_14287,N_13510,N_13638);
xor U14288 (N_14288,N_13944,N_13938);
or U14289 (N_14289,N_13810,N_13565);
and U14290 (N_14290,N_13731,N_13735);
nand U14291 (N_14291,N_13524,N_13565);
and U14292 (N_14292,N_13752,N_13549);
xor U14293 (N_14293,N_13928,N_13648);
or U14294 (N_14294,N_13880,N_13758);
or U14295 (N_14295,N_13759,N_13895);
or U14296 (N_14296,N_13750,N_13737);
xnor U14297 (N_14297,N_13639,N_13768);
nand U14298 (N_14298,N_13532,N_13819);
xor U14299 (N_14299,N_13912,N_13807);
nand U14300 (N_14300,N_13768,N_13917);
and U14301 (N_14301,N_13924,N_13568);
or U14302 (N_14302,N_13501,N_13588);
xnor U14303 (N_14303,N_13972,N_13645);
and U14304 (N_14304,N_13709,N_13513);
or U14305 (N_14305,N_13581,N_13694);
nor U14306 (N_14306,N_13822,N_13684);
nor U14307 (N_14307,N_13567,N_13638);
or U14308 (N_14308,N_13805,N_13627);
and U14309 (N_14309,N_13732,N_13685);
xor U14310 (N_14310,N_13532,N_13797);
nand U14311 (N_14311,N_13744,N_13567);
xnor U14312 (N_14312,N_13669,N_13756);
xor U14313 (N_14313,N_13518,N_13678);
and U14314 (N_14314,N_13583,N_13952);
nand U14315 (N_14315,N_13594,N_13908);
or U14316 (N_14316,N_13647,N_13953);
or U14317 (N_14317,N_13869,N_13813);
xnor U14318 (N_14318,N_13746,N_13677);
xor U14319 (N_14319,N_13850,N_13620);
xor U14320 (N_14320,N_13558,N_13586);
and U14321 (N_14321,N_13516,N_13697);
nor U14322 (N_14322,N_13981,N_13532);
nor U14323 (N_14323,N_13757,N_13571);
xnor U14324 (N_14324,N_13744,N_13729);
and U14325 (N_14325,N_13506,N_13527);
and U14326 (N_14326,N_13632,N_13597);
xnor U14327 (N_14327,N_13618,N_13731);
and U14328 (N_14328,N_13761,N_13721);
nor U14329 (N_14329,N_13699,N_13873);
nand U14330 (N_14330,N_13538,N_13636);
xor U14331 (N_14331,N_13602,N_13726);
xor U14332 (N_14332,N_13518,N_13551);
nand U14333 (N_14333,N_13503,N_13601);
nor U14334 (N_14334,N_13918,N_13986);
xor U14335 (N_14335,N_13632,N_13578);
nand U14336 (N_14336,N_13589,N_13827);
nand U14337 (N_14337,N_13501,N_13641);
or U14338 (N_14338,N_13538,N_13744);
and U14339 (N_14339,N_13559,N_13576);
xnor U14340 (N_14340,N_13603,N_13614);
or U14341 (N_14341,N_13921,N_13792);
nor U14342 (N_14342,N_13504,N_13884);
nand U14343 (N_14343,N_13965,N_13856);
and U14344 (N_14344,N_13677,N_13649);
nand U14345 (N_14345,N_13884,N_13791);
and U14346 (N_14346,N_13689,N_13703);
nand U14347 (N_14347,N_13556,N_13994);
and U14348 (N_14348,N_13857,N_13683);
and U14349 (N_14349,N_13884,N_13758);
nand U14350 (N_14350,N_13783,N_13815);
xnor U14351 (N_14351,N_13725,N_13683);
xnor U14352 (N_14352,N_13561,N_13656);
or U14353 (N_14353,N_13533,N_13930);
and U14354 (N_14354,N_13623,N_13698);
xor U14355 (N_14355,N_13609,N_13817);
and U14356 (N_14356,N_13974,N_13829);
nor U14357 (N_14357,N_13902,N_13934);
nand U14358 (N_14358,N_13904,N_13573);
and U14359 (N_14359,N_13838,N_13540);
or U14360 (N_14360,N_13826,N_13561);
and U14361 (N_14361,N_13791,N_13533);
nor U14362 (N_14362,N_13747,N_13885);
nor U14363 (N_14363,N_13984,N_13972);
and U14364 (N_14364,N_13925,N_13739);
xnor U14365 (N_14365,N_13984,N_13944);
xor U14366 (N_14366,N_13816,N_13709);
and U14367 (N_14367,N_13893,N_13591);
xnor U14368 (N_14368,N_13955,N_13830);
and U14369 (N_14369,N_13986,N_13862);
xnor U14370 (N_14370,N_13507,N_13863);
nor U14371 (N_14371,N_13571,N_13761);
or U14372 (N_14372,N_13721,N_13620);
nand U14373 (N_14373,N_13633,N_13904);
nor U14374 (N_14374,N_13676,N_13789);
nor U14375 (N_14375,N_13820,N_13859);
xnor U14376 (N_14376,N_13718,N_13728);
nor U14377 (N_14377,N_13749,N_13944);
xnor U14378 (N_14378,N_13839,N_13593);
nor U14379 (N_14379,N_13652,N_13704);
xnor U14380 (N_14380,N_13818,N_13981);
and U14381 (N_14381,N_13870,N_13802);
or U14382 (N_14382,N_13867,N_13513);
nor U14383 (N_14383,N_13956,N_13988);
and U14384 (N_14384,N_13507,N_13922);
xor U14385 (N_14385,N_13858,N_13893);
or U14386 (N_14386,N_13959,N_13833);
nor U14387 (N_14387,N_13728,N_13826);
nand U14388 (N_14388,N_13965,N_13850);
nand U14389 (N_14389,N_13783,N_13684);
nor U14390 (N_14390,N_13702,N_13665);
xnor U14391 (N_14391,N_13600,N_13717);
nor U14392 (N_14392,N_13764,N_13755);
nand U14393 (N_14393,N_13950,N_13705);
and U14394 (N_14394,N_13856,N_13735);
nor U14395 (N_14395,N_13799,N_13524);
xor U14396 (N_14396,N_13934,N_13548);
or U14397 (N_14397,N_13681,N_13747);
nand U14398 (N_14398,N_13697,N_13590);
and U14399 (N_14399,N_13733,N_13585);
and U14400 (N_14400,N_13668,N_13828);
or U14401 (N_14401,N_13729,N_13623);
and U14402 (N_14402,N_13723,N_13947);
and U14403 (N_14403,N_13788,N_13839);
or U14404 (N_14404,N_13672,N_13513);
nor U14405 (N_14405,N_13548,N_13606);
xnor U14406 (N_14406,N_13610,N_13785);
and U14407 (N_14407,N_13925,N_13549);
nand U14408 (N_14408,N_13515,N_13513);
xor U14409 (N_14409,N_13822,N_13630);
nor U14410 (N_14410,N_13514,N_13730);
nand U14411 (N_14411,N_13695,N_13558);
nor U14412 (N_14412,N_13614,N_13946);
and U14413 (N_14413,N_13844,N_13835);
nand U14414 (N_14414,N_13669,N_13619);
nor U14415 (N_14415,N_13955,N_13739);
nand U14416 (N_14416,N_13647,N_13599);
nor U14417 (N_14417,N_13850,N_13908);
xnor U14418 (N_14418,N_13920,N_13684);
or U14419 (N_14419,N_13613,N_13588);
nor U14420 (N_14420,N_13540,N_13961);
xnor U14421 (N_14421,N_13652,N_13505);
xor U14422 (N_14422,N_13857,N_13756);
and U14423 (N_14423,N_13817,N_13683);
xnor U14424 (N_14424,N_13607,N_13909);
or U14425 (N_14425,N_13507,N_13943);
and U14426 (N_14426,N_13905,N_13932);
or U14427 (N_14427,N_13678,N_13541);
xnor U14428 (N_14428,N_13985,N_13875);
nand U14429 (N_14429,N_13525,N_13536);
or U14430 (N_14430,N_13501,N_13562);
or U14431 (N_14431,N_13977,N_13759);
nor U14432 (N_14432,N_13599,N_13866);
and U14433 (N_14433,N_13530,N_13863);
xnor U14434 (N_14434,N_13671,N_13981);
nor U14435 (N_14435,N_13680,N_13958);
nor U14436 (N_14436,N_13958,N_13567);
or U14437 (N_14437,N_13696,N_13909);
and U14438 (N_14438,N_13777,N_13743);
and U14439 (N_14439,N_13888,N_13925);
or U14440 (N_14440,N_13788,N_13524);
and U14441 (N_14441,N_13839,N_13825);
and U14442 (N_14442,N_13801,N_13551);
nor U14443 (N_14443,N_13920,N_13956);
nor U14444 (N_14444,N_13948,N_13539);
and U14445 (N_14445,N_13683,N_13671);
and U14446 (N_14446,N_13978,N_13633);
nand U14447 (N_14447,N_13687,N_13620);
or U14448 (N_14448,N_13978,N_13824);
and U14449 (N_14449,N_13661,N_13883);
nand U14450 (N_14450,N_13882,N_13699);
nor U14451 (N_14451,N_13798,N_13620);
and U14452 (N_14452,N_13826,N_13903);
and U14453 (N_14453,N_13694,N_13670);
xnor U14454 (N_14454,N_13718,N_13502);
xnor U14455 (N_14455,N_13509,N_13530);
nor U14456 (N_14456,N_13617,N_13805);
or U14457 (N_14457,N_13792,N_13942);
nor U14458 (N_14458,N_13893,N_13682);
nor U14459 (N_14459,N_13620,N_13919);
or U14460 (N_14460,N_13882,N_13959);
nand U14461 (N_14461,N_13861,N_13530);
nor U14462 (N_14462,N_13812,N_13748);
or U14463 (N_14463,N_13693,N_13536);
xor U14464 (N_14464,N_13730,N_13674);
nor U14465 (N_14465,N_13637,N_13943);
nand U14466 (N_14466,N_13855,N_13715);
xor U14467 (N_14467,N_13916,N_13961);
or U14468 (N_14468,N_13825,N_13960);
nand U14469 (N_14469,N_13786,N_13674);
and U14470 (N_14470,N_13565,N_13737);
nand U14471 (N_14471,N_13609,N_13675);
nor U14472 (N_14472,N_13592,N_13694);
nor U14473 (N_14473,N_13828,N_13659);
xor U14474 (N_14474,N_13579,N_13834);
or U14475 (N_14475,N_13673,N_13988);
nand U14476 (N_14476,N_13861,N_13928);
xnor U14477 (N_14477,N_13892,N_13681);
and U14478 (N_14478,N_13573,N_13689);
nand U14479 (N_14479,N_13963,N_13739);
xor U14480 (N_14480,N_13558,N_13637);
and U14481 (N_14481,N_13743,N_13926);
nand U14482 (N_14482,N_13705,N_13766);
nand U14483 (N_14483,N_13721,N_13803);
and U14484 (N_14484,N_13854,N_13837);
or U14485 (N_14485,N_13518,N_13945);
or U14486 (N_14486,N_13865,N_13762);
or U14487 (N_14487,N_13773,N_13874);
nand U14488 (N_14488,N_13550,N_13519);
xnor U14489 (N_14489,N_13746,N_13682);
and U14490 (N_14490,N_13728,N_13758);
and U14491 (N_14491,N_13855,N_13700);
and U14492 (N_14492,N_13515,N_13575);
nand U14493 (N_14493,N_13942,N_13965);
or U14494 (N_14494,N_13547,N_13865);
and U14495 (N_14495,N_13771,N_13747);
nand U14496 (N_14496,N_13701,N_13597);
nor U14497 (N_14497,N_13515,N_13715);
xnor U14498 (N_14498,N_13887,N_13979);
and U14499 (N_14499,N_13960,N_13554);
and U14500 (N_14500,N_14103,N_14010);
or U14501 (N_14501,N_14362,N_14310);
and U14502 (N_14502,N_14458,N_14283);
xnor U14503 (N_14503,N_14339,N_14089);
or U14504 (N_14504,N_14135,N_14265);
or U14505 (N_14505,N_14222,N_14376);
nand U14506 (N_14506,N_14360,N_14083);
and U14507 (N_14507,N_14436,N_14217);
or U14508 (N_14508,N_14345,N_14357);
xnor U14509 (N_14509,N_14142,N_14261);
nor U14510 (N_14510,N_14391,N_14335);
xnor U14511 (N_14511,N_14324,N_14406);
nand U14512 (N_14512,N_14320,N_14277);
xor U14513 (N_14513,N_14100,N_14491);
nand U14514 (N_14514,N_14461,N_14132);
or U14515 (N_14515,N_14386,N_14157);
or U14516 (N_14516,N_14166,N_14290);
nor U14517 (N_14517,N_14190,N_14229);
or U14518 (N_14518,N_14221,N_14005);
nand U14519 (N_14519,N_14359,N_14060);
nand U14520 (N_14520,N_14304,N_14289);
nand U14521 (N_14521,N_14457,N_14479);
nand U14522 (N_14522,N_14446,N_14216);
xnor U14523 (N_14523,N_14331,N_14119);
or U14524 (N_14524,N_14378,N_14169);
or U14525 (N_14525,N_14058,N_14305);
nand U14526 (N_14526,N_14243,N_14269);
nand U14527 (N_14527,N_14450,N_14381);
xor U14528 (N_14528,N_14490,N_14355);
nor U14529 (N_14529,N_14470,N_14205);
or U14530 (N_14530,N_14498,N_14061);
or U14531 (N_14531,N_14039,N_14480);
and U14532 (N_14532,N_14088,N_14388);
nor U14533 (N_14533,N_14076,N_14227);
and U14534 (N_14534,N_14240,N_14233);
xor U14535 (N_14535,N_14348,N_14108);
and U14536 (N_14536,N_14160,N_14434);
nor U14537 (N_14537,N_14390,N_14318);
nor U14538 (N_14538,N_14091,N_14031);
and U14539 (N_14539,N_14315,N_14412);
xor U14540 (N_14540,N_14057,N_14319);
xnor U14541 (N_14541,N_14257,N_14371);
and U14542 (N_14542,N_14188,N_14116);
nand U14543 (N_14543,N_14198,N_14447);
xnor U14544 (N_14544,N_14373,N_14299);
nor U14545 (N_14545,N_14260,N_14045);
nand U14546 (N_14546,N_14332,N_14475);
nor U14547 (N_14547,N_14080,N_14051);
nor U14548 (N_14548,N_14115,N_14467);
or U14549 (N_14549,N_14140,N_14201);
nand U14550 (N_14550,N_14311,N_14273);
or U14551 (N_14551,N_14050,N_14044);
and U14552 (N_14552,N_14220,N_14055);
nor U14553 (N_14553,N_14382,N_14481);
and U14554 (N_14554,N_14469,N_14397);
or U14555 (N_14555,N_14230,N_14191);
xor U14556 (N_14556,N_14016,N_14268);
or U14557 (N_14557,N_14471,N_14018);
nand U14558 (N_14558,N_14292,N_14123);
xor U14559 (N_14559,N_14054,N_14099);
xor U14560 (N_14560,N_14263,N_14394);
xnor U14561 (N_14561,N_14437,N_14293);
or U14562 (N_14562,N_14183,N_14241);
and U14563 (N_14563,N_14254,N_14445);
nor U14564 (N_14564,N_14365,N_14189);
or U14565 (N_14565,N_14392,N_14175);
and U14566 (N_14566,N_14170,N_14047);
and U14567 (N_14567,N_14377,N_14225);
nand U14568 (N_14568,N_14462,N_14401);
or U14569 (N_14569,N_14246,N_14025);
and U14570 (N_14570,N_14167,N_14426);
nand U14571 (N_14571,N_14094,N_14027);
and U14572 (N_14572,N_14215,N_14164);
xor U14573 (N_14573,N_14042,N_14452);
nand U14574 (N_14574,N_14330,N_14297);
or U14575 (N_14575,N_14049,N_14264);
nor U14576 (N_14576,N_14499,N_14294);
nor U14577 (N_14577,N_14405,N_14137);
and U14578 (N_14578,N_14300,N_14125);
or U14579 (N_14579,N_14008,N_14148);
nor U14580 (N_14580,N_14145,N_14237);
xor U14581 (N_14581,N_14180,N_14464);
or U14582 (N_14582,N_14033,N_14255);
or U14583 (N_14583,N_14107,N_14333);
nor U14584 (N_14584,N_14231,N_14338);
nand U14585 (N_14585,N_14326,N_14483);
nor U14586 (N_14586,N_14364,N_14417);
nor U14587 (N_14587,N_14029,N_14440);
nor U14588 (N_14588,N_14021,N_14347);
and U14589 (N_14589,N_14195,N_14149);
nand U14590 (N_14590,N_14428,N_14172);
nor U14591 (N_14591,N_14262,N_14317);
xor U14592 (N_14592,N_14036,N_14374);
and U14593 (N_14593,N_14072,N_14423);
xor U14594 (N_14594,N_14109,N_14134);
nor U14595 (N_14595,N_14030,N_14282);
and U14596 (N_14596,N_14112,N_14207);
and U14597 (N_14597,N_14303,N_14126);
or U14598 (N_14598,N_14070,N_14380);
xnor U14599 (N_14599,N_14385,N_14007);
and U14600 (N_14600,N_14040,N_14298);
xor U14601 (N_14601,N_14443,N_14253);
nor U14602 (N_14602,N_14403,N_14000);
nand U14603 (N_14603,N_14308,N_14474);
and U14604 (N_14604,N_14037,N_14302);
and U14605 (N_14605,N_14313,N_14287);
xnor U14606 (N_14606,N_14346,N_14141);
or U14607 (N_14607,N_14307,N_14418);
xor U14608 (N_14608,N_14017,N_14489);
nor U14609 (N_14609,N_14204,N_14131);
or U14610 (N_14610,N_14492,N_14150);
and U14611 (N_14611,N_14156,N_14448);
nand U14612 (N_14612,N_14473,N_14267);
nand U14613 (N_14613,N_14223,N_14138);
xnor U14614 (N_14614,N_14214,N_14465);
nand U14615 (N_14615,N_14079,N_14349);
or U14616 (N_14616,N_14487,N_14419);
or U14617 (N_14617,N_14139,N_14059);
nand U14618 (N_14618,N_14463,N_14117);
nand U14619 (N_14619,N_14168,N_14001);
and U14620 (N_14620,N_14466,N_14478);
nand U14621 (N_14621,N_14363,N_14092);
xor U14622 (N_14622,N_14093,N_14232);
nor U14623 (N_14623,N_14351,N_14398);
nand U14624 (N_14624,N_14206,N_14194);
nor U14625 (N_14625,N_14043,N_14155);
nand U14626 (N_14626,N_14105,N_14200);
xor U14627 (N_14627,N_14323,N_14258);
nor U14628 (N_14628,N_14098,N_14210);
nor U14629 (N_14629,N_14130,N_14366);
and U14630 (N_14630,N_14078,N_14372);
or U14631 (N_14631,N_14369,N_14329);
or U14632 (N_14632,N_14411,N_14336);
or U14633 (N_14633,N_14022,N_14414);
xor U14634 (N_14634,N_14396,N_14352);
nor U14635 (N_14635,N_14178,N_14291);
nor U14636 (N_14636,N_14484,N_14438);
nand U14637 (N_14637,N_14306,N_14006);
nor U14638 (N_14638,N_14028,N_14409);
nor U14639 (N_14639,N_14035,N_14375);
or U14640 (N_14640,N_14090,N_14358);
and U14641 (N_14641,N_14041,N_14482);
and U14642 (N_14642,N_14361,N_14176);
xnor U14643 (N_14643,N_14325,N_14128);
and U14644 (N_14644,N_14337,N_14309);
xnor U14645 (N_14645,N_14424,N_14328);
and U14646 (N_14646,N_14496,N_14165);
and U14647 (N_14647,N_14278,N_14387);
nand U14648 (N_14648,N_14250,N_14288);
or U14649 (N_14649,N_14075,N_14235);
nor U14650 (N_14650,N_14065,N_14082);
nor U14651 (N_14651,N_14236,N_14173);
and U14652 (N_14652,N_14185,N_14399);
or U14653 (N_14653,N_14367,N_14276);
xor U14654 (N_14654,N_14129,N_14281);
or U14655 (N_14655,N_14182,N_14468);
nand U14656 (N_14656,N_14284,N_14177);
nor U14657 (N_14657,N_14350,N_14003);
nor U14658 (N_14658,N_14096,N_14181);
or U14659 (N_14659,N_14454,N_14136);
or U14660 (N_14660,N_14422,N_14486);
and U14661 (N_14661,N_14013,N_14111);
nor U14662 (N_14662,N_14151,N_14420);
and U14663 (N_14663,N_14296,N_14400);
and U14664 (N_14664,N_14113,N_14071);
and U14665 (N_14665,N_14285,N_14015);
or U14666 (N_14666,N_14012,N_14280);
xnor U14667 (N_14667,N_14034,N_14073);
nand U14668 (N_14668,N_14106,N_14407);
xor U14669 (N_14669,N_14192,N_14066);
xnor U14670 (N_14670,N_14162,N_14147);
xnor U14671 (N_14671,N_14408,N_14161);
or U14672 (N_14672,N_14179,N_14327);
nand U14673 (N_14673,N_14046,N_14154);
nand U14674 (N_14674,N_14270,N_14014);
nand U14675 (N_14675,N_14024,N_14272);
nand U14676 (N_14676,N_14444,N_14416);
or U14677 (N_14677,N_14095,N_14354);
or U14678 (N_14678,N_14238,N_14455);
xnor U14679 (N_14679,N_14218,N_14228);
xor U14680 (N_14680,N_14067,N_14477);
xor U14681 (N_14681,N_14384,N_14431);
and U14682 (N_14682,N_14493,N_14342);
xnor U14683 (N_14683,N_14146,N_14274);
or U14684 (N_14684,N_14286,N_14251);
nor U14685 (N_14685,N_14197,N_14144);
and U14686 (N_14686,N_14085,N_14341);
nor U14687 (N_14687,N_14442,N_14171);
nor U14688 (N_14688,N_14494,N_14026);
nor U14689 (N_14689,N_14402,N_14202);
nor U14690 (N_14690,N_14224,N_14433);
nand U14691 (N_14691,N_14213,N_14032);
and U14692 (N_14692,N_14495,N_14019);
xor U14693 (N_14693,N_14389,N_14211);
or U14694 (N_14694,N_14226,N_14084);
nor U14695 (N_14695,N_14456,N_14193);
or U14696 (N_14696,N_14020,N_14248);
nor U14697 (N_14697,N_14485,N_14356);
nor U14698 (N_14698,N_14184,N_14203);
nor U14699 (N_14699,N_14104,N_14322);
xor U14700 (N_14700,N_14209,N_14343);
and U14701 (N_14701,N_14383,N_14245);
nand U14702 (N_14702,N_14038,N_14159);
or U14703 (N_14703,N_14081,N_14114);
nand U14704 (N_14704,N_14124,N_14208);
or U14705 (N_14705,N_14314,N_14295);
and U14706 (N_14706,N_14143,N_14275);
nand U14707 (N_14707,N_14404,N_14425);
and U14708 (N_14708,N_14158,N_14064);
and U14709 (N_14709,N_14212,N_14252);
and U14710 (N_14710,N_14097,N_14023);
nand U14711 (N_14711,N_14497,N_14110);
and U14712 (N_14712,N_14009,N_14174);
and U14713 (N_14713,N_14234,N_14087);
or U14714 (N_14714,N_14476,N_14102);
or U14715 (N_14715,N_14393,N_14249);
nor U14716 (N_14716,N_14063,N_14199);
nand U14717 (N_14717,N_14186,N_14413);
and U14718 (N_14718,N_14122,N_14163);
xor U14719 (N_14719,N_14279,N_14052);
nor U14720 (N_14720,N_14353,N_14316);
and U14721 (N_14721,N_14415,N_14133);
or U14722 (N_14722,N_14062,N_14077);
nor U14723 (N_14723,N_14451,N_14048);
xor U14724 (N_14724,N_14053,N_14395);
xnor U14725 (N_14725,N_14056,N_14256);
nor U14726 (N_14726,N_14459,N_14271);
or U14727 (N_14727,N_14344,N_14247);
nor U14728 (N_14728,N_14069,N_14086);
nand U14729 (N_14729,N_14488,N_14187);
nor U14730 (N_14730,N_14439,N_14370);
xnor U14731 (N_14731,N_14430,N_14196);
or U14732 (N_14732,N_14368,N_14121);
nor U14733 (N_14733,N_14340,N_14101);
nand U14734 (N_14734,N_14453,N_14239);
nand U14735 (N_14735,N_14244,N_14118);
xor U14736 (N_14736,N_14379,N_14002);
or U14737 (N_14737,N_14074,N_14266);
nand U14738 (N_14738,N_14127,N_14410);
or U14739 (N_14739,N_14259,N_14472);
and U14740 (N_14740,N_14242,N_14427);
nor U14741 (N_14741,N_14435,N_14321);
or U14742 (N_14742,N_14449,N_14312);
xnor U14743 (N_14743,N_14432,N_14219);
and U14744 (N_14744,N_14011,N_14441);
or U14745 (N_14745,N_14152,N_14068);
xnor U14746 (N_14746,N_14004,N_14460);
or U14747 (N_14747,N_14120,N_14429);
nand U14748 (N_14748,N_14421,N_14334);
nor U14749 (N_14749,N_14153,N_14301);
nor U14750 (N_14750,N_14039,N_14346);
or U14751 (N_14751,N_14408,N_14292);
and U14752 (N_14752,N_14317,N_14099);
nor U14753 (N_14753,N_14010,N_14406);
or U14754 (N_14754,N_14144,N_14168);
or U14755 (N_14755,N_14285,N_14257);
nor U14756 (N_14756,N_14431,N_14491);
nor U14757 (N_14757,N_14058,N_14261);
nor U14758 (N_14758,N_14049,N_14395);
or U14759 (N_14759,N_14339,N_14088);
xnor U14760 (N_14760,N_14238,N_14074);
nor U14761 (N_14761,N_14236,N_14153);
nand U14762 (N_14762,N_14070,N_14168);
or U14763 (N_14763,N_14360,N_14251);
nor U14764 (N_14764,N_14377,N_14098);
xnor U14765 (N_14765,N_14420,N_14489);
and U14766 (N_14766,N_14345,N_14188);
nand U14767 (N_14767,N_14358,N_14155);
nand U14768 (N_14768,N_14067,N_14194);
nor U14769 (N_14769,N_14358,N_14431);
nand U14770 (N_14770,N_14464,N_14057);
or U14771 (N_14771,N_14101,N_14089);
xnor U14772 (N_14772,N_14488,N_14076);
xnor U14773 (N_14773,N_14395,N_14414);
xor U14774 (N_14774,N_14290,N_14368);
and U14775 (N_14775,N_14449,N_14297);
or U14776 (N_14776,N_14060,N_14143);
or U14777 (N_14777,N_14126,N_14014);
or U14778 (N_14778,N_14090,N_14248);
nand U14779 (N_14779,N_14300,N_14434);
and U14780 (N_14780,N_14147,N_14005);
xnor U14781 (N_14781,N_14318,N_14384);
and U14782 (N_14782,N_14197,N_14093);
and U14783 (N_14783,N_14207,N_14487);
nor U14784 (N_14784,N_14147,N_14239);
or U14785 (N_14785,N_14121,N_14228);
nor U14786 (N_14786,N_14434,N_14008);
and U14787 (N_14787,N_14275,N_14293);
or U14788 (N_14788,N_14154,N_14497);
or U14789 (N_14789,N_14277,N_14294);
or U14790 (N_14790,N_14230,N_14472);
xor U14791 (N_14791,N_14069,N_14021);
nand U14792 (N_14792,N_14076,N_14405);
or U14793 (N_14793,N_14110,N_14164);
or U14794 (N_14794,N_14166,N_14146);
xor U14795 (N_14795,N_14333,N_14034);
xnor U14796 (N_14796,N_14205,N_14425);
nor U14797 (N_14797,N_14336,N_14179);
xnor U14798 (N_14798,N_14005,N_14046);
nor U14799 (N_14799,N_14419,N_14148);
or U14800 (N_14800,N_14317,N_14200);
or U14801 (N_14801,N_14485,N_14273);
nand U14802 (N_14802,N_14137,N_14330);
xnor U14803 (N_14803,N_14174,N_14143);
xnor U14804 (N_14804,N_14038,N_14360);
xnor U14805 (N_14805,N_14344,N_14335);
and U14806 (N_14806,N_14067,N_14173);
nor U14807 (N_14807,N_14230,N_14131);
nand U14808 (N_14808,N_14282,N_14052);
nor U14809 (N_14809,N_14003,N_14254);
or U14810 (N_14810,N_14314,N_14188);
nor U14811 (N_14811,N_14468,N_14287);
nand U14812 (N_14812,N_14115,N_14459);
nand U14813 (N_14813,N_14376,N_14449);
or U14814 (N_14814,N_14342,N_14155);
nand U14815 (N_14815,N_14125,N_14411);
nor U14816 (N_14816,N_14042,N_14057);
and U14817 (N_14817,N_14114,N_14494);
xor U14818 (N_14818,N_14158,N_14010);
nor U14819 (N_14819,N_14141,N_14114);
nor U14820 (N_14820,N_14291,N_14235);
xnor U14821 (N_14821,N_14268,N_14350);
nor U14822 (N_14822,N_14026,N_14430);
xnor U14823 (N_14823,N_14418,N_14395);
nand U14824 (N_14824,N_14154,N_14141);
nand U14825 (N_14825,N_14152,N_14280);
or U14826 (N_14826,N_14441,N_14070);
nor U14827 (N_14827,N_14364,N_14450);
xnor U14828 (N_14828,N_14413,N_14022);
and U14829 (N_14829,N_14352,N_14312);
nor U14830 (N_14830,N_14218,N_14219);
or U14831 (N_14831,N_14428,N_14425);
xor U14832 (N_14832,N_14355,N_14323);
nand U14833 (N_14833,N_14271,N_14220);
or U14834 (N_14834,N_14450,N_14475);
or U14835 (N_14835,N_14093,N_14435);
and U14836 (N_14836,N_14420,N_14498);
and U14837 (N_14837,N_14248,N_14264);
or U14838 (N_14838,N_14093,N_14283);
nor U14839 (N_14839,N_14128,N_14216);
or U14840 (N_14840,N_14266,N_14076);
xor U14841 (N_14841,N_14376,N_14255);
nand U14842 (N_14842,N_14244,N_14125);
nand U14843 (N_14843,N_14003,N_14328);
and U14844 (N_14844,N_14357,N_14341);
and U14845 (N_14845,N_14083,N_14070);
xnor U14846 (N_14846,N_14128,N_14242);
nor U14847 (N_14847,N_14045,N_14338);
nand U14848 (N_14848,N_14385,N_14362);
nand U14849 (N_14849,N_14408,N_14400);
nand U14850 (N_14850,N_14242,N_14171);
nand U14851 (N_14851,N_14130,N_14418);
or U14852 (N_14852,N_14160,N_14396);
nand U14853 (N_14853,N_14480,N_14489);
or U14854 (N_14854,N_14311,N_14128);
nor U14855 (N_14855,N_14108,N_14177);
nor U14856 (N_14856,N_14327,N_14230);
nor U14857 (N_14857,N_14176,N_14109);
nand U14858 (N_14858,N_14197,N_14392);
nor U14859 (N_14859,N_14244,N_14492);
nand U14860 (N_14860,N_14236,N_14076);
and U14861 (N_14861,N_14167,N_14136);
and U14862 (N_14862,N_14426,N_14100);
nor U14863 (N_14863,N_14426,N_14079);
and U14864 (N_14864,N_14316,N_14268);
nand U14865 (N_14865,N_14441,N_14331);
xnor U14866 (N_14866,N_14224,N_14367);
nand U14867 (N_14867,N_14069,N_14058);
or U14868 (N_14868,N_14380,N_14276);
and U14869 (N_14869,N_14390,N_14468);
nor U14870 (N_14870,N_14466,N_14055);
nand U14871 (N_14871,N_14077,N_14324);
and U14872 (N_14872,N_14426,N_14076);
or U14873 (N_14873,N_14272,N_14235);
nand U14874 (N_14874,N_14468,N_14086);
and U14875 (N_14875,N_14309,N_14060);
nor U14876 (N_14876,N_14065,N_14395);
nor U14877 (N_14877,N_14178,N_14135);
and U14878 (N_14878,N_14003,N_14225);
xnor U14879 (N_14879,N_14090,N_14450);
and U14880 (N_14880,N_14216,N_14186);
or U14881 (N_14881,N_14293,N_14127);
nand U14882 (N_14882,N_14417,N_14434);
nor U14883 (N_14883,N_14381,N_14447);
xnor U14884 (N_14884,N_14138,N_14440);
nor U14885 (N_14885,N_14342,N_14371);
nand U14886 (N_14886,N_14287,N_14417);
or U14887 (N_14887,N_14445,N_14459);
nor U14888 (N_14888,N_14177,N_14201);
nor U14889 (N_14889,N_14499,N_14321);
nand U14890 (N_14890,N_14407,N_14491);
or U14891 (N_14891,N_14274,N_14217);
nor U14892 (N_14892,N_14189,N_14448);
and U14893 (N_14893,N_14182,N_14280);
nand U14894 (N_14894,N_14263,N_14441);
or U14895 (N_14895,N_14485,N_14255);
and U14896 (N_14896,N_14002,N_14356);
nand U14897 (N_14897,N_14447,N_14231);
or U14898 (N_14898,N_14158,N_14021);
nor U14899 (N_14899,N_14164,N_14295);
nor U14900 (N_14900,N_14470,N_14267);
nor U14901 (N_14901,N_14235,N_14288);
nand U14902 (N_14902,N_14335,N_14280);
nand U14903 (N_14903,N_14386,N_14355);
nand U14904 (N_14904,N_14421,N_14418);
xor U14905 (N_14905,N_14295,N_14457);
nand U14906 (N_14906,N_14348,N_14450);
and U14907 (N_14907,N_14417,N_14101);
nand U14908 (N_14908,N_14040,N_14480);
nor U14909 (N_14909,N_14370,N_14169);
xor U14910 (N_14910,N_14395,N_14167);
or U14911 (N_14911,N_14059,N_14405);
xor U14912 (N_14912,N_14443,N_14319);
and U14913 (N_14913,N_14370,N_14403);
nand U14914 (N_14914,N_14282,N_14234);
xor U14915 (N_14915,N_14209,N_14392);
nor U14916 (N_14916,N_14466,N_14286);
xnor U14917 (N_14917,N_14248,N_14407);
and U14918 (N_14918,N_14335,N_14208);
and U14919 (N_14919,N_14121,N_14249);
xor U14920 (N_14920,N_14044,N_14018);
nor U14921 (N_14921,N_14188,N_14102);
nor U14922 (N_14922,N_14288,N_14088);
or U14923 (N_14923,N_14474,N_14387);
nand U14924 (N_14924,N_14323,N_14030);
nand U14925 (N_14925,N_14206,N_14100);
xor U14926 (N_14926,N_14304,N_14394);
nand U14927 (N_14927,N_14092,N_14249);
and U14928 (N_14928,N_14137,N_14173);
and U14929 (N_14929,N_14326,N_14140);
xnor U14930 (N_14930,N_14124,N_14210);
nor U14931 (N_14931,N_14162,N_14074);
or U14932 (N_14932,N_14364,N_14237);
and U14933 (N_14933,N_14207,N_14256);
or U14934 (N_14934,N_14386,N_14441);
xnor U14935 (N_14935,N_14028,N_14486);
nand U14936 (N_14936,N_14377,N_14282);
xor U14937 (N_14937,N_14113,N_14201);
nor U14938 (N_14938,N_14429,N_14223);
and U14939 (N_14939,N_14307,N_14453);
nor U14940 (N_14940,N_14383,N_14265);
nand U14941 (N_14941,N_14061,N_14476);
nor U14942 (N_14942,N_14173,N_14404);
nor U14943 (N_14943,N_14147,N_14462);
nand U14944 (N_14944,N_14387,N_14026);
nand U14945 (N_14945,N_14154,N_14267);
and U14946 (N_14946,N_14279,N_14258);
xnor U14947 (N_14947,N_14020,N_14122);
nor U14948 (N_14948,N_14178,N_14127);
nor U14949 (N_14949,N_14112,N_14358);
nand U14950 (N_14950,N_14456,N_14405);
xnor U14951 (N_14951,N_14239,N_14382);
xor U14952 (N_14952,N_14338,N_14229);
nor U14953 (N_14953,N_14464,N_14424);
xor U14954 (N_14954,N_14193,N_14365);
nor U14955 (N_14955,N_14429,N_14080);
or U14956 (N_14956,N_14490,N_14233);
nand U14957 (N_14957,N_14086,N_14463);
xnor U14958 (N_14958,N_14316,N_14137);
nand U14959 (N_14959,N_14301,N_14150);
or U14960 (N_14960,N_14097,N_14116);
nand U14961 (N_14961,N_14195,N_14203);
nor U14962 (N_14962,N_14395,N_14171);
nand U14963 (N_14963,N_14123,N_14447);
nor U14964 (N_14964,N_14376,N_14284);
nand U14965 (N_14965,N_14099,N_14489);
or U14966 (N_14966,N_14460,N_14287);
nand U14967 (N_14967,N_14194,N_14265);
nand U14968 (N_14968,N_14264,N_14286);
or U14969 (N_14969,N_14047,N_14205);
and U14970 (N_14970,N_14407,N_14328);
and U14971 (N_14971,N_14411,N_14139);
xnor U14972 (N_14972,N_14302,N_14093);
xnor U14973 (N_14973,N_14265,N_14340);
nor U14974 (N_14974,N_14212,N_14409);
and U14975 (N_14975,N_14317,N_14095);
nand U14976 (N_14976,N_14358,N_14369);
nor U14977 (N_14977,N_14089,N_14237);
nor U14978 (N_14978,N_14254,N_14335);
or U14979 (N_14979,N_14330,N_14353);
nor U14980 (N_14980,N_14369,N_14432);
or U14981 (N_14981,N_14409,N_14376);
or U14982 (N_14982,N_14176,N_14475);
nor U14983 (N_14983,N_14165,N_14456);
xnor U14984 (N_14984,N_14301,N_14268);
nand U14985 (N_14985,N_14055,N_14385);
or U14986 (N_14986,N_14186,N_14192);
nor U14987 (N_14987,N_14430,N_14384);
and U14988 (N_14988,N_14248,N_14240);
and U14989 (N_14989,N_14208,N_14479);
nor U14990 (N_14990,N_14473,N_14038);
or U14991 (N_14991,N_14427,N_14172);
or U14992 (N_14992,N_14459,N_14085);
nand U14993 (N_14993,N_14201,N_14065);
and U14994 (N_14994,N_14144,N_14262);
or U14995 (N_14995,N_14495,N_14279);
nor U14996 (N_14996,N_14458,N_14152);
and U14997 (N_14997,N_14181,N_14144);
or U14998 (N_14998,N_14204,N_14445);
xor U14999 (N_14999,N_14356,N_14030);
nand U15000 (N_15000,N_14809,N_14515);
nand U15001 (N_15001,N_14831,N_14876);
nand U15002 (N_15002,N_14897,N_14532);
nand U15003 (N_15003,N_14712,N_14665);
nand U15004 (N_15004,N_14603,N_14577);
nor U15005 (N_15005,N_14600,N_14816);
nand U15006 (N_15006,N_14837,N_14954);
or U15007 (N_15007,N_14738,N_14502);
nor U15008 (N_15008,N_14860,N_14955);
nand U15009 (N_15009,N_14592,N_14854);
xnor U15010 (N_15010,N_14664,N_14678);
or U15011 (N_15011,N_14653,N_14609);
or U15012 (N_15012,N_14898,N_14749);
xnor U15013 (N_15013,N_14740,N_14743);
nor U15014 (N_15014,N_14602,N_14776);
nand U15015 (N_15015,N_14943,N_14588);
nor U15016 (N_15016,N_14680,N_14983);
nor U15017 (N_15017,N_14701,N_14541);
xnor U15018 (N_15018,N_14607,N_14675);
and U15019 (N_15019,N_14704,N_14727);
and U15020 (N_15020,N_14972,N_14919);
nand U15021 (N_15021,N_14579,N_14610);
nand U15022 (N_15022,N_14571,N_14930);
xor U15023 (N_15023,N_14878,N_14873);
nand U15024 (N_15024,N_14666,N_14779);
xnor U15025 (N_15025,N_14732,N_14549);
or U15026 (N_15026,N_14901,N_14881);
nor U15027 (N_15027,N_14775,N_14906);
xnor U15028 (N_15028,N_14889,N_14656);
nor U15029 (N_15029,N_14572,N_14636);
or U15030 (N_15030,N_14514,N_14566);
nand U15031 (N_15031,N_14709,N_14748);
and U15032 (N_15032,N_14542,N_14753);
or U15033 (N_15033,N_14500,N_14751);
and U15034 (N_15034,N_14817,N_14747);
xnor U15035 (N_15035,N_14795,N_14950);
or U15036 (N_15036,N_14679,N_14715);
xnor U15037 (N_15037,N_14564,N_14528);
xor U15038 (N_15038,N_14931,N_14804);
nand U15039 (N_15039,N_14755,N_14843);
nor U15040 (N_15040,N_14540,N_14990);
nor U15041 (N_15041,N_14962,N_14763);
xnor U15042 (N_15042,N_14619,N_14702);
nor U15043 (N_15043,N_14660,N_14924);
and U15044 (N_15044,N_14767,N_14840);
nand U15045 (N_15045,N_14615,N_14956);
or U15046 (N_15046,N_14896,N_14848);
and U15047 (N_15047,N_14829,N_14773);
and U15048 (N_15048,N_14786,N_14605);
nor U15049 (N_15049,N_14811,N_14882);
nand U15050 (N_15050,N_14842,N_14525);
xor U15051 (N_15051,N_14558,N_14714);
and U15052 (N_15052,N_14988,N_14676);
and U15053 (N_15053,N_14511,N_14953);
nor U15054 (N_15054,N_14670,N_14844);
nand U15055 (N_15055,N_14760,N_14830);
or U15056 (N_15056,N_14576,N_14641);
and U15057 (N_15057,N_14698,N_14909);
xnor U15058 (N_15058,N_14874,N_14699);
nand U15059 (N_15059,N_14929,N_14877);
and U15060 (N_15060,N_14810,N_14513);
nand U15061 (N_15061,N_14824,N_14730);
nand U15062 (N_15062,N_14718,N_14964);
nand U15063 (N_15063,N_14958,N_14852);
nor U15064 (N_15064,N_14995,N_14963);
nor U15065 (N_15065,N_14914,N_14923);
nor U15066 (N_15066,N_14681,N_14868);
nand U15067 (N_15067,N_14737,N_14922);
and U15068 (N_15068,N_14569,N_14859);
xnor U15069 (N_15069,N_14543,N_14783);
xnor U15070 (N_15070,N_14517,N_14721);
or U15071 (N_15071,N_14757,N_14875);
xor U15072 (N_15072,N_14947,N_14766);
nand U15073 (N_15073,N_14710,N_14555);
nand U15074 (N_15074,N_14700,N_14774);
or U15075 (N_15075,N_14893,N_14907);
nor U15076 (N_15076,N_14815,N_14601);
nor U15077 (N_15077,N_14890,N_14946);
nand U15078 (N_15078,N_14913,N_14970);
nor U15079 (N_15079,N_14663,N_14677);
nor U15080 (N_15080,N_14512,N_14805);
nor U15081 (N_15081,N_14550,N_14501);
xnor U15082 (N_15082,N_14981,N_14682);
or U15083 (N_15083,N_14520,N_14765);
xor U15084 (N_15084,N_14537,N_14790);
or U15085 (N_15085,N_14904,N_14633);
or U15086 (N_15086,N_14761,N_14966);
and U15087 (N_15087,N_14870,N_14625);
nand U15088 (N_15088,N_14917,N_14888);
nor U15089 (N_15089,N_14937,N_14823);
or U15090 (N_15090,N_14503,N_14582);
and U15091 (N_15091,N_14750,N_14940);
nor U15092 (N_15092,N_14782,N_14869);
or U15093 (N_15093,N_14985,N_14973);
nand U15094 (N_15094,N_14855,N_14960);
xor U15095 (N_15095,N_14819,N_14637);
and U15096 (N_15096,N_14587,N_14705);
or U15097 (N_15097,N_14975,N_14802);
xor U15098 (N_15098,N_14814,N_14581);
nor U15099 (N_15099,N_14711,N_14785);
nand U15100 (N_15100,N_14526,N_14857);
nor U15101 (N_15101,N_14825,N_14616);
nand U15102 (N_15102,N_14647,N_14627);
and U15103 (N_15103,N_14659,N_14735);
xnor U15104 (N_15104,N_14694,N_14912);
xnor U15105 (N_15105,N_14703,N_14872);
or U15106 (N_15106,N_14974,N_14553);
xor U15107 (N_15107,N_14987,N_14768);
xor U15108 (N_15108,N_14936,N_14563);
and U15109 (N_15109,N_14832,N_14803);
nand U15110 (N_15110,N_14865,N_14691);
or U15111 (N_15111,N_14853,N_14724);
or U15112 (N_15112,N_14567,N_14662);
xnor U15113 (N_15113,N_14673,N_14927);
nand U15114 (N_15114,N_14593,N_14591);
and U15115 (N_15115,N_14792,N_14657);
or U15116 (N_15116,N_14826,N_14984);
nand U15117 (N_15117,N_14746,N_14573);
nor U15118 (N_15118,N_14754,N_14903);
or U15119 (N_15119,N_14643,N_14630);
nand U15120 (N_15120,N_14734,N_14575);
xnor U15121 (N_15121,N_14533,N_14851);
xnor U15122 (N_15122,N_14725,N_14612);
nor U15123 (N_15123,N_14871,N_14626);
or U15124 (N_15124,N_14589,N_14764);
and U15125 (N_15125,N_14979,N_14519);
xnor U15126 (N_15126,N_14818,N_14925);
nand U15127 (N_15127,N_14693,N_14733);
or U15128 (N_15128,N_14742,N_14769);
xor U15129 (N_15129,N_14808,N_14892);
nor U15130 (N_15130,N_14684,N_14723);
nor U15131 (N_15131,N_14720,N_14644);
nor U15132 (N_15132,N_14864,N_14863);
or U15133 (N_15133,N_14849,N_14505);
and U15134 (N_15134,N_14989,N_14686);
and U15135 (N_15135,N_14518,N_14726);
xor U15136 (N_15136,N_14507,N_14772);
and U15137 (N_15137,N_14799,N_14687);
and U15138 (N_15138,N_14939,N_14793);
xnor U15139 (N_15139,N_14547,N_14642);
nor U15140 (N_15140,N_14992,N_14902);
and U15141 (N_15141,N_14949,N_14654);
or U15142 (N_15142,N_14690,N_14828);
xor U15143 (N_15143,N_14570,N_14621);
and U15144 (N_15144,N_14697,N_14944);
or U15145 (N_15145,N_14632,N_14778);
nand U15146 (N_15146,N_14961,N_14504);
or U15147 (N_15147,N_14696,N_14640);
nor U15148 (N_15148,N_14586,N_14996);
nand U15149 (N_15149,N_14866,N_14986);
xnor U15150 (N_15150,N_14546,N_14813);
or U15151 (N_15151,N_14821,N_14729);
nor U15152 (N_15152,N_14527,N_14617);
nand U15153 (N_15153,N_14822,N_14980);
xor U15154 (N_15154,N_14516,N_14856);
and U15155 (N_15155,N_14997,N_14834);
nor U15156 (N_15156,N_14941,N_14789);
and U15157 (N_15157,N_14535,N_14999);
xor U15158 (N_15158,N_14798,N_14744);
and U15159 (N_15159,N_14781,N_14736);
xnor U15160 (N_15160,N_14580,N_14771);
or U15161 (N_15161,N_14993,N_14599);
xor U15162 (N_15162,N_14545,N_14523);
and U15163 (N_15163,N_14948,N_14928);
nor U15164 (N_15164,N_14841,N_14672);
nand U15165 (N_15165,N_14652,N_14611);
nor U15166 (N_15166,N_14649,N_14568);
or U15167 (N_15167,N_14982,N_14622);
or U15168 (N_15168,N_14791,N_14595);
nor U15169 (N_15169,N_14536,N_14594);
and U15170 (N_15170,N_14762,N_14935);
nand U15171 (N_15171,N_14574,N_14584);
or U15172 (N_15172,N_14596,N_14638);
nand U15173 (N_15173,N_14971,N_14506);
nor U15174 (N_15174,N_14998,N_14938);
nand U15175 (N_15175,N_14658,N_14634);
or U15176 (N_15176,N_14604,N_14552);
nor U15177 (N_15177,N_14752,N_14692);
xor U15178 (N_15178,N_14784,N_14531);
nand U15179 (N_15179,N_14838,N_14994);
or U15180 (N_15180,N_14548,N_14661);
xnor U15181 (N_15181,N_14777,N_14926);
xor U15182 (N_15182,N_14846,N_14539);
nand U15183 (N_15183,N_14608,N_14707);
and U15184 (N_15184,N_14886,N_14991);
and U15185 (N_15185,N_14880,N_14916);
or U15186 (N_15186,N_14965,N_14648);
nand U15187 (N_15187,N_14780,N_14639);
nand U15188 (N_15188,N_14557,N_14957);
nand U15189 (N_15189,N_14894,N_14806);
or U15190 (N_15190,N_14706,N_14770);
nand U15191 (N_15191,N_14561,N_14969);
xor U15192 (N_15192,N_14529,N_14833);
nand U15193 (N_15193,N_14651,N_14534);
or U15194 (N_15194,N_14835,N_14967);
nor U15195 (N_15195,N_14560,N_14758);
xnor U15196 (N_15196,N_14614,N_14952);
and U15197 (N_15197,N_14884,N_14689);
nor U15198 (N_15198,N_14820,N_14942);
nand U15199 (N_15199,N_14891,N_14508);
xnor U15200 (N_15200,N_14858,N_14669);
nand U15201 (N_15201,N_14847,N_14708);
and U15202 (N_15202,N_14827,N_14900);
nor U15203 (N_15203,N_14812,N_14674);
xor U15204 (N_15204,N_14624,N_14620);
nand U15205 (N_15205,N_14597,N_14731);
xor U15206 (N_15206,N_14728,N_14578);
and U15207 (N_15207,N_14631,N_14861);
or U15208 (N_15208,N_14551,N_14683);
xor U15209 (N_15209,N_14671,N_14667);
xor U15210 (N_15210,N_14976,N_14741);
nor U15211 (N_15211,N_14899,N_14629);
and U15212 (N_15212,N_14745,N_14554);
or U15213 (N_15213,N_14945,N_14717);
nor U15214 (N_15214,N_14668,N_14911);
nor U15215 (N_15215,N_14716,N_14650);
and U15216 (N_15216,N_14583,N_14635);
nand U15217 (N_15217,N_14739,N_14918);
and U15218 (N_15218,N_14606,N_14801);
nand U15219 (N_15219,N_14510,N_14932);
xnor U15220 (N_15220,N_14509,N_14522);
nand U15221 (N_15221,N_14887,N_14977);
and U15222 (N_15222,N_14836,N_14895);
or U15223 (N_15223,N_14951,N_14862);
nor U15224 (N_15224,N_14807,N_14688);
and U15225 (N_15225,N_14565,N_14796);
nor U15226 (N_15226,N_14905,N_14645);
nand U15227 (N_15227,N_14685,N_14559);
xnor U15228 (N_15228,N_14524,N_14885);
nor U15229 (N_15229,N_14756,N_14968);
nand U15230 (N_15230,N_14618,N_14920);
or U15231 (N_15231,N_14713,N_14556);
nor U15232 (N_15232,N_14628,N_14646);
xnor U15233 (N_15233,N_14719,N_14530);
nand U15234 (N_15234,N_14839,N_14585);
and U15235 (N_15235,N_14908,N_14910);
xnor U15236 (N_15236,N_14722,N_14797);
nor U15237 (N_15237,N_14978,N_14613);
xnor U15238 (N_15238,N_14921,N_14934);
nand U15239 (N_15239,N_14800,N_14695);
nand U15240 (N_15240,N_14794,N_14787);
nand U15241 (N_15241,N_14544,N_14590);
nand U15242 (N_15242,N_14598,N_14759);
and U15243 (N_15243,N_14879,N_14788);
nor U15244 (N_15244,N_14538,N_14933);
or U15245 (N_15245,N_14521,N_14655);
xnor U15246 (N_15246,N_14959,N_14850);
nor U15247 (N_15247,N_14623,N_14883);
xnor U15248 (N_15248,N_14562,N_14915);
or U15249 (N_15249,N_14867,N_14845);
nor U15250 (N_15250,N_14506,N_14735);
xnor U15251 (N_15251,N_14536,N_14743);
nand U15252 (N_15252,N_14599,N_14875);
or U15253 (N_15253,N_14595,N_14714);
xnor U15254 (N_15254,N_14663,N_14582);
or U15255 (N_15255,N_14542,N_14892);
or U15256 (N_15256,N_14667,N_14534);
or U15257 (N_15257,N_14793,N_14946);
or U15258 (N_15258,N_14694,N_14587);
xor U15259 (N_15259,N_14815,N_14794);
xnor U15260 (N_15260,N_14694,N_14685);
xnor U15261 (N_15261,N_14555,N_14727);
nand U15262 (N_15262,N_14577,N_14642);
and U15263 (N_15263,N_14654,N_14563);
and U15264 (N_15264,N_14731,N_14591);
nand U15265 (N_15265,N_14577,N_14721);
or U15266 (N_15266,N_14578,N_14992);
nand U15267 (N_15267,N_14995,N_14822);
or U15268 (N_15268,N_14606,N_14641);
xnor U15269 (N_15269,N_14900,N_14548);
nor U15270 (N_15270,N_14844,N_14815);
nor U15271 (N_15271,N_14669,N_14673);
xor U15272 (N_15272,N_14543,N_14729);
and U15273 (N_15273,N_14739,N_14851);
nor U15274 (N_15274,N_14673,N_14792);
or U15275 (N_15275,N_14944,N_14634);
and U15276 (N_15276,N_14757,N_14520);
or U15277 (N_15277,N_14967,N_14834);
or U15278 (N_15278,N_14581,N_14628);
and U15279 (N_15279,N_14517,N_14618);
nand U15280 (N_15280,N_14570,N_14804);
nand U15281 (N_15281,N_14799,N_14537);
or U15282 (N_15282,N_14933,N_14730);
or U15283 (N_15283,N_14578,N_14589);
nor U15284 (N_15284,N_14605,N_14950);
xnor U15285 (N_15285,N_14701,N_14757);
xnor U15286 (N_15286,N_14629,N_14912);
or U15287 (N_15287,N_14815,N_14691);
and U15288 (N_15288,N_14925,N_14970);
xnor U15289 (N_15289,N_14919,N_14530);
nand U15290 (N_15290,N_14635,N_14619);
nand U15291 (N_15291,N_14645,N_14544);
nor U15292 (N_15292,N_14622,N_14729);
or U15293 (N_15293,N_14676,N_14647);
or U15294 (N_15294,N_14720,N_14990);
nand U15295 (N_15295,N_14578,N_14951);
nand U15296 (N_15296,N_14600,N_14808);
nor U15297 (N_15297,N_14658,N_14982);
xor U15298 (N_15298,N_14661,N_14849);
nor U15299 (N_15299,N_14866,N_14772);
nand U15300 (N_15300,N_14861,N_14828);
and U15301 (N_15301,N_14656,N_14801);
and U15302 (N_15302,N_14752,N_14977);
nor U15303 (N_15303,N_14979,N_14717);
nand U15304 (N_15304,N_14814,N_14652);
and U15305 (N_15305,N_14917,N_14687);
or U15306 (N_15306,N_14541,N_14873);
nand U15307 (N_15307,N_14837,N_14752);
and U15308 (N_15308,N_14567,N_14933);
nor U15309 (N_15309,N_14603,N_14997);
and U15310 (N_15310,N_14537,N_14731);
and U15311 (N_15311,N_14726,N_14598);
nand U15312 (N_15312,N_14542,N_14931);
nor U15313 (N_15313,N_14926,N_14659);
nand U15314 (N_15314,N_14748,N_14627);
nor U15315 (N_15315,N_14677,N_14657);
and U15316 (N_15316,N_14544,N_14682);
or U15317 (N_15317,N_14880,N_14800);
nor U15318 (N_15318,N_14601,N_14565);
nor U15319 (N_15319,N_14516,N_14615);
nor U15320 (N_15320,N_14708,N_14519);
nor U15321 (N_15321,N_14708,N_14867);
or U15322 (N_15322,N_14515,N_14503);
xnor U15323 (N_15323,N_14763,N_14588);
or U15324 (N_15324,N_14700,N_14940);
xnor U15325 (N_15325,N_14801,N_14641);
nor U15326 (N_15326,N_14728,N_14894);
nor U15327 (N_15327,N_14892,N_14669);
and U15328 (N_15328,N_14927,N_14668);
nand U15329 (N_15329,N_14511,N_14649);
and U15330 (N_15330,N_14843,N_14507);
nor U15331 (N_15331,N_14993,N_14692);
xnor U15332 (N_15332,N_14838,N_14674);
and U15333 (N_15333,N_14778,N_14638);
and U15334 (N_15334,N_14874,N_14669);
and U15335 (N_15335,N_14709,N_14584);
and U15336 (N_15336,N_14551,N_14748);
xor U15337 (N_15337,N_14709,N_14908);
and U15338 (N_15338,N_14569,N_14899);
and U15339 (N_15339,N_14645,N_14573);
nor U15340 (N_15340,N_14777,N_14709);
nand U15341 (N_15341,N_14670,N_14545);
nand U15342 (N_15342,N_14586,N_14673);
nand U15343 (N_15343,N_14589,N_14716);
or U15344 (N_15344,N_14856,N_14993);
and U15345 (N_15345,N_14724,N_14966);
and U15346 (N_15346,N_14905,N_14798);
xnor U15347 (N_15347,N_14540,N_14784);
or U15348 (N_15348,N_14546,N_14653);
or U15349 (N_15349,N_14800,N_14512);
xor U15350 (N_15350,N_14518,N_14989);
nor U15351 (N_15351,N_14800,N_14839);
or U15352 (N_15352,N_14932,N_14743);
and U15353 (N_15353,N_14868,N_14749);
or U15354 (N_15354,N_14769,N_14676);
xor U15355 (N_15355,N_14587,N_14563);
and U15356 (N_15356,N_14649,N_14693);
xor U15357 (N_15357,N_14921,N_14503);
xor U15358 (N_15358,N_14869,N_14875);
nand U15359 (N_15359,N_14584,N_14852);
or U15360 (N_15360,N_14791,N_14735);
or U15361 (N_15361,N_14676,N_14620);
and U15362 (N_15362,N_14692,N_14884);
xnor U15363 (N_15363,N_14823,N_14528);
nor U15364 (N_15364,N_14886,N_14828);
xor U15365 (N_15365,N_14983,N_14601);
nand U15366 (N_15366,N_14687,N_14785);
nor U15367 (N_15367,N_14691,N_14803);
xor U15368 (N_15368,N_14958,N_14534);
or U15369 (N_15369,N_14928,N_14754);
nand U15370 (N_15370,N_14933,N_14799);
xnor U15371 (N_15371,N_14968,N_14736);
xnor U15372 (N_15372,N_14952,N_14783);
xnor U15373 (N_15373,N_14548,N_14804);
or U15374 (N_15374,N_14615,N_14754);
or U15375 (N_15375,N_14678,N_14753);
xnor U15376 (N_15376,N_14753,N_14613);
or U15377 (N_15377,N_14897,N_14717);
and U15378 (N_15378,N_14815,N_14760);
or U15379 (N_15379,N_14712,N_14990);
nand U15380 (N_15380,N_14705,N_14902);
or U15381 (N_15381,N_14858,N_14654);
xor U15382 (N_15382,N_14812,N_14726);
nand U15383 (N_15383,N_14785,N_14937);
xor U15384 (N_15384,N_14606,N_14809);
nor U15385 (N_15385,N_14527,N_14776);
or U15386 (N_15386,N_14528,N_14755);
nand U15387 (N_15387,N_14872,N_14519);
or U15388 (N_15388,N_14924,N_14684);
nand U15389 (N_15389,N_14746,N_14999);
and U15390 (N_15390,N_14984,N_14924);
nor U15391 (N_15391,N_14676,N_14722);
nor U15392 (N_15392,N_14588,N_14856);
and U15393 (N_15393,N_14718,N_14785);
nor U15394 (N_15394,N_14833,N_14756);
nor U15395 (N_15395,N_14824,N_14956);
nand U15396 (N_15396,N_14891,N_14549);
or U15397 (N_15397,N_14598,N_14584);
or U15398 (N_15398,N_14564,N_14772);
and U15399 (N_15399,N_14957,N_14737);
nand U15400 (N_15400,N_14832,N_14663);
and U15401 (N_15401,N_14655,N_14863);
nor U15402 (N_15402,N_14536,N_14769);
nor U15403 (N_15403,N_14750,N_14925);
nor U15404 (N_15404,N_14792,N_14817);
or U15405 (N_15405,N_14566,N_14651);
xnor U15406 (N_15406,N_14551,N_14949);
or U15407 (N_15407,N_14676,N_14657);
nand U15408 (N_15408,N_14655,N_14805);
xor U15409 (N_15409,N_14907,N_14703);
xor U15410 (N_15410,N_14602,N_14556);
nor U15411 (N_15411,N_14663,N_14554);
nand U15412 (N_15412,N_14762,N_14517);
and U15413 (N_15413,N_14996,N_14674);
nor U15414 (N_15414,N_14519,N_14891);
nor U15415 (N_15415,N_14967,N_14826);
and U15416 (N_15416,N_14990,N_14755);
xor U15417 (N_15417,N_14794,N_14554);
or U15418 (N_15418,N_14674,N_14853);
and U15419 (N_15419,N_14722,N_14987);
xor U15420 (N_15420,N_14638,N_14651);
nor U15421 (N_15421,N_14837,N_14722);
and U15422 (N_15422,N_14645,N_14912);
nand U15423 (N_15423,N_14754,N_14668);
or U15424 (N_15424,N_14681,N_14583);
or U15425 (N_15425,N_14604,N_14883);
nor U15426 (N_15426,N_14642,N_14870);
or U15427 (N_15427,N_14764,N_14717);
or U15428 (N_15428,N_14950,N_14957);
or U15429 (N_15429,N_14944,N_14637);
nor U15430 (N_15430,N_14966,N_14899);
nor U15431 (N_15431,N_14802,N_14941);
xnor U15432 (N_15432,N_14892,N_14911);
or U15433 (N_15433,N_14745,N_14928);
nand U15434 (N_15434,N_14874,N_14695);
or U15435 (N_15435,N_14901,N_14867);
and U15436 (N_15436,N_14507,N_14510);
or U15437 (N_15437,N_14761,N_14743);
xnor U15438 (N_15438,N_14875,N_14634);
nand U15439 (N_15439,N_14773,N_14657);
xor U15440 (N_15440,N_14805,N_14643);
and U15441 (N_15441,N_14867,N_14629);
and U15442 (N_15442,N_14942,N_14643);
xnor U15443 (N_15443,N_14550,N_14798);
nor U15444 (N_15444,N_14647,N_14925);
and U15445 (N_15445,N_14754,N_14979);
nand U15446 (N_15446,N_14872,N_14988);
nand U15447 (N_15447,N_14594,N_14892);
nand U15448 (N_15448,N_14818,N_14908);
nor U15449 (N_15449,N_14771,N_14768);
nor U15450 (N_15450,N_14893,N_14667);
nor U15451 (N_15451,N_14507,N_14574);
and U15452 (N_15452,N_14535,N_14594);
xnor U15453 (N_15453,N_14931,N_14685);
nor U15454 (N_15454,N_14982,N_14940);
nor U15455 (N_15455,N_14614,N_14561);
and U15456 (N_15456,N_14903,N_14721);
nand U15457 (N_15457,N_14782,N_14842);
nand U15458 (N_15458,N_14949,N_14826);
xnor U15459 (N_15459,N_14962,N_14597);
and U15460 (N_15460,N_14976,N_14881);
nand U15461 (N_15461,N_14721,N_14820);
nor U15462 (N_15462,N_14809,N_14921);
nand U15463 (N_15463,N_14687,N_14673);
nand U15464 (N_15464,N_14978,N_14775);
nand U15465 (N_15465,N_14851,N_14751);
nor U15466 (N_15466,N_14501,N_14839);
nand U15467 (N_15467,N_14699,N_14767);
nor U15468 (N_15468,N_14712,N_14976);
and U15469 (N_15469,N_14781,N_14596);
and U15470 (N_15470,N_14582,N_14844);
xnor U15471 (N_15471,N_14970,N_14840);
and U15472 (N_15472,N_14652,N_14563);
and U15473 (N_15473,N_14946,N_14682);
or U15474 (N_15474,N_14646,N_14843);
xnor U15475 (N_15475,N_14884,N_14847);
xor U15476 (N_15476,N_14949,N_14969);
and U15477 (N_15477,N_14922,N_14815);
and U15478 (N_15478,N_14547,N_14935);
or U15479 (N_15479,N_14986,N_14806);
nor U15480 (N_15480,N_14672,N_14957);
and U15481 (N_15481,N_14866,N_14537);
xnor U15482 (N_15482,N_14711,N_14864);
and U15483 (N_15483,N_14607,N_14571);
and U15484 (N_15484,N_14796,N_14709);
xor U15485 (N_15485,N_14817,N_14504);
or U15486 (N_15486,N_14589,N_14617);
xor U15487 (N_15487,N_14599,N_14509);
xor U15488 (N_15488,N_14529,N_14943);
nand U15489 (N_15489,N_14718,N_14960);
or U15490 (N_15490,N_14814,N_14692);
and U15491 (N_15491,N_14765,N_14968);
or U15492 (N_15492,N_14564,N_14925);
nor U15493 (N_15493,N_14638,N_14923);
nor U15494 (N_15494,N_14838,N_14651);
nand U15495 (N_15495,N_14551,N_14974);
nand U15496 (N_15496,N_14576,N_14904);
and U15497 (N_15497,N_14696,N_14985);
nand U15498 (N_15498,N_14714,N_14716);
or U15499 (N_15499,N_14533,N_14875);
or U15500 (N_15500,N_15427,N_15267);
and U15501 (N_15501,N_15373,N_15472);
nand U15502 (N_15502,N_15494,N_15364);
and U15503 (N_15503,N_15159,N_15318);
nand U15504 (N_15504,N_15467,N_15073);
nand U15505 (N_15505,N_15395,N_15014);
nor U15506 (N_15506,N_15123,N_15361);
and U15507 (N_15507,N_15382,N_15431);
xnor U15508 (N_15508,N_15369,N_15356);
and U15509 (N_15509,N_15474,N_15184);
and U15510 (N_15510,N_15259,N_15058);
or U15511 (N_15511,N_15277,N_15186);
or U15512 (N_15512,N_15384,N_15432);
and U15513 (N_15513,N_15232,N_15194);
or U15514 (N_15514,N_15346,N_15397);
nor U15515 (N_15515,N_15291,N_15054);
and U15516 (N_15516,N_15045,N_15111);
and U15517 (N_15517,N_15250,N_15486);
and U15518 (N_15518,N_15377,N_15233);
and U15519 (N_15519,N_15283,N_15446);
or U15520 (N_15520,N_15452,N_15115);
or U15521 (N_15521,N_15362,N_15386);
nand U15522 (N_15522,N_15444,N_15090);
nor U15523 (N_15523,N_15132,N_15400);
nand U15524 (N_15524,N_15198,N_15425);
and U15525 (N_15525,N_15288,N_15099);
xnor U15526 (N_15526,N_15183,N_15448);
nor U15527 (N_15527,N_15281,N_15426);
or U15528 (N_15528,N_15249,N_15398);
and U15529 (N_15529,N_15015,N_15161);
nor U15530 (N_15530,N_15036,N_15342);
or U15531 (N_15531,N_15315,N_15418);
xor U15532 (N_15532,N_15306,N_15326);
nor U15533 (N_15533,N_15244,N_15255);
nand U15534 (N_15534,N_15087,N_15335);
nor U15535 (N_15535,N_15025,N_15088);
or U15536 (N_15536,N_15327,N_15016);
and U15537 (N_15537,N_15145,N_15465);
nand U15538 (N_15538,N_15313,N_15089);
nand U15539 (N_15539,N_15049,N_15236);
nor U15540 (N_15540,N_15153,N_15304);
nor U15541 (N_15541,N_15126,N_15310);
xor U15542 (N_15542,N_15336,N_15443);
xnor U15543 (N_15543,N_15164,N_15032);
and U15544 (N_15544,N_15231,N_15333);
nor U15545 (N_15545,N_15329,N_15018);
xor U15546 (N_15546,N_15389,N_15275);
xor U15547 (N_15547,N_15061,N_15478);
nand U15548 (N_15548,N_15173,N_15119);
xnor U15549 (N_15549,N_15210,N_15404);
or U15550 (N_15550,N_15293,N_15167);
xor U15551 (N_15551,N_15453,N_15043);
nand U15552 (N_15552,N_15168,N_15254);
xnor U15553 (N_15553,N_15357,N_15353);
nor U15554 (N_15554,N_15095,N_15013);
xor U15555 (N_15555,N_15470,N_15358);
nand U15556 (N_15556,N_15050,N_15429);
xnor U15557 (N_15557,N_15227,N_15321);
nand U15558 (N_15558,N_15181,N_15022);
nor U15559 (N_15559,N_15436,N_15039);
xor U15560 (N_15560,N_15270,N_15407);
xor U15561 (N_15561,N_15122,N_15152);
and U15562 (N_15562,N_15038,N_15347);
nor U15563 (N_15563,N_15071,N_15140);
or U15564 (N_15564,N_15121,N_15337);
or U15565 (N_15565,N_15282,N_15187);
xnor U15566 (N_15566,N_15053,N_15157);
nor U15567 (N_15567,N_15352,N_15320);
nor U15568 (N_15568,N_15136,N_15135);
and U15569 (N_15569,N_15492,N_15174);
or U15570 (N_15570,N_15114,N_15219);
nand U15571 (N_15571,N_15031,N_15002);
nand U15572 (N_15572,N_15112,N_15247);
nor U15573 (N_15573,N_15451,N_15480);
nand U15574 (N_15574,N_15142,N_15151);
nand U15575 (N_15575,N_15172,N_15106);
xor U15576 (N_15576,N_15476,N_15417);
nor U15577 (N_15577,N_15348,N_15003);
xnor U15578 (N_15578,N_15411,N_15006);
or U15579 (N_15579,N_15066,N_15276);
or U15580 (N_15580,N_15185,N_15265);
or U15581 (N_15581,N_15289,N_15030);
nor U15582 (N_15582,N_15178,N_15148);
nand U15583 (N_15583,N_15496,N_15208);
nor U15584 (N_15584,N_15332,N_15302);
or U15585 (N_15585,N_15284,N_15158);
nor U15586 (N_15586,N_15242,N_15438);
nand U15587 (N_15587,N_15299,N_15199);
xor U15588 (N_15588,N_15498,N_15027);
nand U15589 (N_15589,N_15440,N_15412);
nand U15590 (N_15590,N_15169,N_15261);
or U15591 (N_15591,N_15056,N_15387);
or U15592 (N_15592,N_15029,N_15359);
nor U15593 (N_15593,N_15235,N_15278);
xnor U15594 (N_15594,N_15221,N_15241);
and U15595 (N_15595,N_15383,N_15256);
or U15596 (N_15596,N_15421,N_15192);
nor U15597 (N_15597,N_15323,N_15298);
or U15598 (N_15598,N_15495,N_15316);
nand U15599 (N_15599,N_15449,N_15442);
or U15600 (N_15600,N_15379,N_15294);
xnor U15601 (N_15601,N_15213,N_15269);
xor U15602 (N_15602,N_15084,N_15092);
and U15603 (N_15603,N_15473,N_15034);
and U15604 (N_15604,N_15351,N_15339);
nand U15605 (N_15605,N_15005,N_15266);
xor U15606 (N_15606,N_15206,N_15487);
nor U15607 (N_15607,N_15202,N_15295);
nor U15608 (N_15608,N_15416,N_15055);
nand U15609 (N_15609,N_15454,N_15120);
or U15610 (N_15610,N_15490,N_15201);
or U15611 (N_15611,N_15380,N_15104);
xor U15612 (N_15612,N_15414,N_15406);
xor U15613 (N_15613,N_15000,N_15493);
and U15614 (N_15614,N_15141,N_15497);
xnor U15615 (N_15615,N_15251,N_15481);
nor U15616 (N_15616,N_15393,N_15220);
and U15617 (N_15617,N_15489,N_15485);
nor U15618 (N_15618,N_15450,N_15190);
and U15619 (N_15619,N_15366,N_15064);
and U15620 (N_15620,N_15154,N_15057);
xnor U15621 (N_15621,N_15238,N_15216);
or U15622 (N_15622,N_15280,N_15457);
xnor U15623 (N_15623,N_15008,N_15130);
xnor U15624 (N_15624,N_15224,N_15410);
and U15625 (N_15625,N_15477,N_15330);
xnor U15626 (N_15626,N_15195,N_15286);
nor U15627 (N_15627,N_15149,N_15100);
nand U15628 (N_15628,N_15466,N_15372);
nor U15629 (N_15629,N_15127,N_15360);
or U15630 (N_15630,N_15047,N_15409);
nand U15631 (N_15631,N_15463,N_15079);
nand U15632 (N_15632,N_15180,N_15239);
xnor U15633 (N_15633,N_15461,N_15097);
and U15634 (N_15634,N_15488,N_15021);
nor U15635 (N_15635,N_15462,N_15033);
nor U15636 (N_15636,N_15285,N_15160);
or U15637 (N_15637,N_15129,N_15143);
nor U15638 (N_15638,N_15307,N_15037);
xnor U15639 (N_15639,N_15253,N_15009);
and U15640 (N_15640,N_15063,N_15207);
and U15641 (N_15641,N_15028,N_15205);
xnor U15642 (N_15642,N_15052,N_15113);
nand U15643 (N_15643,N_15246,N_15203);
nand U15644 (N_15644,N_15471,N_15076);
and U15645 (N_15645,N_15262,N_15072);
nor U15646 (N_15646,N_15434,N_15197);
and U15647 (N_15647,N_15078,N_15370);
or U15648 (N_15648,N_15396,N_15458);
xor U15649 (N_15649,N_15083,N_15222);
xnor U15650 (N_15650,N_15215,N_15441);
nand U15651 (N_15651,N_15096,N_15312);
and U15652 (N_15652,N_15371,N_15223);
and U15653 (N_15653,N_15475,N_15303);
or U15654 (N_15654,N_15101,N_15188);
xor U15655 (N_15655,N_15428,N_15011);
nand U15656 (N_15656,N_15430,N_15040);
and U15657 (N_15657,N_15133,N_15023);
xor U15658 (N_15658,N_15196,N_15290);
xor U15659 (N_15659,N_15062,N_15166);
or U15660 (N_15660,N_15258,N_15212);
or U15661 (N_15661,N_15234,N_15403);
xnor U15662 (N_15662,N_15368,N_15193);
xor U15663 (N_15663,N_15455,N_15138);
nor U15664 (N_15664,N_15399,N_15279);
and U15665 (N_15665,N_15001,N_15060);
nor U15666 (N_15666,N_15182,N_15086);
nand U15667 (N_15667,N_15217,N_15075);
or U15668 (N_15668,N_15109,N_15098);
or U15669 (N_15669,N_15273,N_15419);
and U15670 (N_15670,N_15243,N_15124);
or U15671 (N_15671,N_15110,N_15354);
and U15672 (N_15672,N_15103,N_15211);
xnor U15673 (N_15673,N_15069,N_15317);
and U15674 (N_15674,N_15391,N_15007);
nand U15675 (N_15675,N_15445,N_15345);
or U15676 (N_15676,N_15191,N_15085);
or U15677 (N_15677,N_15435,N_15128);
nor U15678 (N_15678,N_15020,N_15162);
xnor U15679 (N_15679,N_15051,N_15482);
and U15680 (N_15680,N_15413,N_15338);
nand U15681 (N_15681,N_15156,N_15026);
or U15682 (N_15682,N_15204,N_15093);
and U15683 (N_15683,N_15402,N_15245);
nand U15684 (N_15684,N_15107,N_15146);
or U15685 (N_15685,N_15150,N_15340);
or U15686 (N_15686,N_15375,N_15134);
or U15687 (N_15687,N_15248,N_15226);
nand U15688 (N_15688,N_15287,N_15139);
or U15689 (N_15689,N_15237,N_15144);
xor U15690 (N_15690,N_15230,N_15044);
xnor U15691 (N_15691,N_15041,N_15491);
or U15692 (N_15692,N_15456,N_15401);
or U15693 (N_15693,N_15343,N_15171);
or U15694 (N_15694,N_15464,N_15268);
xnor U15695 (N_15695,N_15263,N_15059);
nand U15696 (N_15696,N_15048,N_15314);
or U15697 (N_15697,N_15296,N_15479);
nand U15698 (N_15698,N_15350,N_15300);
nor U15699 (N_15699,N_15272,N_15355);
nor U15700 (N_15700,N_15292,N_15070);
xor U15701 (N_15701,N_15165,N_15468);
xor U15702 (N_15702,N_15175,N_15408);
xnor U15703 (N_15703,N_15271,N_15415);
and U15704 (N_15704,N_15147,N_15209);
nor U15705 (N_15705,N_15170,N_15378);
nand U15706 (N_15706,N_15388,N_15305);
nor U15707 (N_15707,N_15010,N_15424);
and U15708 (N_15708,N_15376,N_15214);
nand U15709 (N_15709,N_15325,N_15125);
nor U15710 (N_15710,N_15200,N_15228);
xnor U15711 (N_15711,N_15082,N_15177);
nor U15712 (N_15712,N_15117,N_15017);
or U15713 (N_15713,N_15484,N_15309);
xor U15714 (N_15714,N_15322,N_15042);
xnor U15715 (N_15715,N_15319,N_15447);
nor U15716 (N_15716,N_15067,N_15324);
nor U15717 (N_15717,N_15301,N_15118);
or U15718 (N_15718,N_15240,N_15394);
nand U15719 (N_15719,N_15341,N_15439);
nor U15720 (N_15720,N_15483,N_15019);
nand U15721 (N_15721,N_15331,N_15163);
nand U15722 (N_15722,N_15229,N_15102);
xor U15723 (N_15723,N_15077,N_15094);
and U15724 (N_15724,N_15499,N_15176);
nand U15725 (N_15725,N_15422,N_15423);
and U15726 (N_15726,N_15367,N_15297);
nand U15727 (N_15727,N_15091,N_15334);
nor U15728 (N_15728,N_15035,N_15080);
nor U15729 (N_15729,N_15252,N_15349);
xor U15730 (N_15730,N_15108,N_15068);
nor U15731 (N_15731,N_15137,N_15257);
nor U15732 (N_15732,N_15024,N_15381);
or U15733 (N_15733,N_15433,N_15328);
or U15734 (N_15734,N_15460,N_15311);
nor U15735 (N_15735,N_15459,N_15074);
nor U15736 (N_15736,N_15469,N_15012);
and U15737 (N_15737,N_15189,N_15390);
nor U15738 (N_15738,N_15308,N_15179);
or U15739 (N_15739,N_15405,N_15420);
and U15740 (N_15740,N_15385,N_15225);
or U15741 (N_15741,N_15274,N_15004);
nand U15742 (N_15742,N_15374,N_15046);
xnor U15743 (N_15743,N_15344,N_15437);
xor U15744 (N_15744,N_15105,N_15081);
and U15745 (N_15745,N_15116,N_15218);
or U15746 (N_15746,N_15065,N_15363);
nor U15747 (N_15747,N_15131,N_15264);
xnor U15748 (N_15748,N_15365,N_15155);
nor U15749 (N_15749,N_15392,N_15260);
nor U15750 (N_15750,N_15101,N_15425);
xor U15751 (N_15751,N_15433,N_15087);
nand U15752 (N_15752,N_15291,N_15090);
xnor U15753 (N_15753,N_15128,N_15266);
or U15754 (N_15754,N_15028,N_15310);
xnor U15755 (N_15755,N_15218,N_15295);
or U15756 (N_15756,N_15487,N_15176);
and U15757 (N_15757,N_15084,N_15366);
or U15758 (N_15758,N_15020,N_15486);
or U15759 (N_15759,N_15023,N_15479);
or U15760 (N_15760,N_15426,N_15280);
nand U15761 (N_15761,N_15309,N_15362);
nor U15762 (N_15762,N_15078,N_15046);
xnor U15763 (N_15763,N_15309,N_15385);
and U15764 (N_15764,N_15058,N_15052);
or U15765 (N_15765,N_15176,N_15271);
and U15766 (N_15766,N_15227,N_15074);
and U15767 (N_15767,N_15329,N_15436);
xor U15768 (N_15768,N_15263,N_15135);
nor U15769 (N_15769,N_15299,N_15233);
nand U15770 (N_15770,N_15464,N_15064);
xnor U15771 (N_15771,N_15315,N_15463);
nand U15772 (N_15772,N_15475,N_15160);
xor U15773 (N_15773,N_15123,N_15279);
or U15774 (N_15774,N_15300,N_15028);
nor U15775 (N_15775,N_15227,N_15047);
xnor U15776 (N_15776,N_15397,N_15143);
nand U15777 (N_15777,N_15388,N_15021);
or U15778 (N_15778,N_15328,N_15030);
nor U15779 (N_15779,N_15246,N_15467);
nand U15780 (N_15780,N_15373,N_15428);
or U15781 (N_15781,N_15071,N_15127);
xnor U15782 (N_15782,N_15284,N_15245);
nor U15783 (N_15783,N_15108,N_15101);
xor U15784 (N_15784,N_15487,N_15108);
and U15785 (N_15785,N_15215,N_15387);
nand U15786 (N_15786,N_15202,N_15462);
nor U15787 (N_15787,N_15355,N_15491);
nand U15788 (N_15788,N_15391,N_15127);
nor U15789 (N_15789,N_15307,N_15186);
or U15790 (N_15790,N_15186,N_15372);
or U15791 (N_15791,N_15042,N_15113);
nor U15792 (N_15792,N_15281,N_15415);
or U15793 (N_15793,N_15082,N_15332);
xor U15794 (N_15794,N_15179,N_15121);
nand U15795 (N_15795,N_15073,N_15228);
nor U15796 (N_15796,N_15246,N_15052);
nor U15797 (N_15797,N_15493,N_15173);
nor U15798 (N_15798,N_15452,N_15143);
and U15799 (N_15799,N_15095,N_15216);
xor U15800 (N_15800,N_15242,N_15166);
and U15801 (N_15801,N_15110,N_15113);
nor U15802 (N_15802,N_15245,N_15471);
nand U15803 (N_15803,N_15000,N_15186);
nor U15804 (N_15804,N_15061,N_15484);
and U15805 (N_15805,N_15292,N_15433);
nor U15806 (N_15806,N_15241,N_15226);
nor U15807 (N_15807,N_15354,N_15480);
and U15808 (N_15808,N_15012,N_15245);
nand U15809 (N_15809,N_15393,N_15209);
and U15810 (N_15810,N_15224,N_15214);
nor U15811 (N_15811,N_15210,N_15242);
or U15812 (N_15812,N_15399,N_15250);
nor U15813 (N_15813,N_15070,N_15442);
xnor U15814 (N_15814,N_15169,N_15354);
xnor U15815 (N_15815,N_15329,N_15017);
or U15816 (N_15816,N_15407,N_15115);
or U15817 (N_15817,N_15408,N_15019);
xnor U15818 (N_15818,N_15057,N_15472);
nand U15819 (N_15819,N_15259,N_15078);
nor U15820 (N_15820,N_15351,N_15034);
nor U15821 (N_15821,N_15073,N_15322);
or U15822 (N_15822,N_15163,N_15358);
xor U15823 (N_15823,N_15236,N_15351);
nor U15824 (N_15824,N_15050,N_15159);
and U15825 (N_15825,N_15464,N_15033);
and U15826 (N_15826,N_15215,N_15055);
nand U15827 (N_15827,N_15457,N_15486);
or U15828 (N_15828,N_15102,N_15452);
or U15829 (N_15829,N_15362,N_15443);
xor U15830 (N_15830,N_15342,N_15441);
nor U15831 (N_15831,N_15159,N_15345);
and U15832 (N_15832,N_15300,N_15256);
and U15833 (N_15833,N_15181,N_15049);
xnor U15834 (N_15834,N_15367,N_15371);
or U15835 (N_15835,N_15233,N_15484);
nor U15836 (N_15836,N_15309,N_15422);
xor U15837 (N_15837,N_15269,N_15454);
or U15838 (N_15838,N_15199,N_15030);
or U15839 (N_15839,N_15055,N_15222);
nor U15840 (N_15840,N_15104,N_15128);
or U15841 (N_15841,N_15296,N_15072);
or U15842 (N_15842,N_15406,N_15204);
and U15843 (N_15843,N_15303,N_15402);
nand U15844 (N_15844,N_15144,N_15100);
or U15845 (N_15845,N_15353,N_15140);
or U15846 (N_15846,N_15238,N_15025);
xnor U15847 (N_15847,N_15487,N_15029);
xnor U15848 (N_15848,N_15144,N_15165);
nand U15849 (N_15849,N_15442,N_15436);
or U15850 (N_15850,N_15028,N_15371);
or U15851 (N_15851,N_15359,N_15457);
nand U15852 (N_15852,N_15409,N_15068);
and U15853 (N_15853,N_15003,N_15315);
or U15854 (N_15854,N_15190,N_15270);
xor U15855 (N_15855,N_15004,N_15266);
xnor U15856 (N_15856,N_15271,N_15290);
nor U15857 (N_15857,N_15126,N_15340);
and U15858 (N_15858,N_15420,N_15101);
nor U15859 (N_15859,N_15323,N_15248);
and U15860 (N_15860,N_15392,N_15413);
xor U15861 (N_15861,N_15192,N_15402);
nor U15862 (N_15862,N_15211,N_15411);
nor U15863 (N_15863,N_15159,N_15436);
nor U15864 (N_15864,N_15470,N_15071);
or U15865 (N_15865,N_15003,N_15243);
or U15866 (N_15866,N_15074,N_15029);
nand U15867 (N_15867,N_15126,N_15141);
nand U15868 (N_15868,N_15346,N_15348);
nor U15869 (N_15869,N_15039,N_15317);
nor U15870 (N_15870,N_15019,N_15329);
and U15871 (N_15871,N_15446,N_15024);
nand U15872 (N_15872,N_15042,N_15055);
xnor U15873 (N_15873,N_15465,N_15230);
xnor U15874 (N_15874,N_15164,N_15442);
or U15875 (N_15875,N_15091,N_15389);
and U15876 (N_15876,N_15081,N_15269);
nor U15877 (N_15877,N_15472,N_15015);
xnor U15878 (N_15878,N_15071,N_15361);
nand U15879 (N_15879,N_15261,N_15385);
xor U15880 (N_15880,N_15169,N_15369);
and U15881 (N_15881,N_15249,N_15446);
nor U15882 (N_15882,N_15271,N_15049);
or U15883 (N_15883,N_15289,N_15178);
xnor U15884 (N_15884,N_15380,N_15224);
nand U15885 (N_15885,N_15131,N_15325);
xnor U15886 (N_15886,N_15263,N_15216);
xnor U15887 (N_15887,N_15020,N_15076);
or U15888 (N_15888,N_15131,N_15275);
or U15889 (N_15889,N_15135,N_15044);
or U15890 (N_15890,N_15343,N_15138);
or U15891 (N_15891,N_15404,N_15183);
or U15892 (N_15892,N_15389,N_15172);
or U15893 (N_15893,N_15113,N_15014);
nor U15894 (N_15894,N_15262,N_15461);
and U15895 (N_15895,N_15078,N_15090);
xor U15896 (N_15896,N_15032,N_15167);
nand U15897 (N_15897,N_15476,N_15100);
nand U15898 (N_15898,N_15072,N_15006);
xnor U15899 (N_15899,N_15494,N_15223);
nand U15900 (N_15900,N_15000,N_15389);
xnor U15901 (N_15901,N_15009,N_15274);
or U15902 (N_15902,N_15366,N_15348);
or U15903 (N_15903,N_15194,N_15411);
xor U15904 (N_15904,N_15021,N_15274);
nand U15905 (N_15905,N_15174,N_15357);
and U15906 (N_15906,N_15189,N_15396);
or U15907 (N_15907,N_15342,N_15278);
and U15908 (N_15908,N_15131,N_15034);
xor U15909 (N_15909,N_15325,N_15477);
and U15910 (N_15910,N_15361,N_15404);
and U15911 (N_15911,N_15410,N_15291);
nand U15912 (N_15912,N_15143,N_15470);
nor U15913 (N_15913,N_15170,N_15004);
and U15914 (N_15914,N_15141,N_15133);
nand U15915 (N_15915,N_15126,N_15210);
nor U15916 (N_15916,N_15375,N_15023);
and U15917 (N_15917,N_15491,N_15223);
xor U15918 (N_15918,N_15417,N_15323);
xor U15919 (N_15919,N_15190,N_15065);
or U15920 (N_15920,N_15491,N_15441);
nor U15921 (N_15921,N_15170,N_15068);
nor U15922 (N_15922,N_15353,N_15137);
nor U15923 (N_15923,N_15216,N_15217);
nor U15924 (N_15924,N_15439,N_15156);
or U15925 (N_15925,N_15359,N_15416);
nand U15926 (N_15926,N_15329,N_15309);
or U15927 (N_15927,N_15221,N_15126);
xor U15928 (N_15928,N_15055,N_15072);
xnor U15929 (N_15929,N_15104,N_15186);
xor U15930 (N_15930,N_15067,N_15412);
or U15931 (N_15931,N_15073,N_15406);
xor U15932 (N_15932,N_15340,N_15268);
nor U15933 (N_15933,N_15433,N_15191);
nor U15934 (N_15934,N_15005,N_15104);
and U15935 (N_15935,N_15066,N_15444);
and U15936 (N_15936,N_15281,N_15223);
nand U15937 (N_15937,N_15268,N_15177);
xor U15938 (N_15938,N_15365,N_15444);
xor U15939 (N_15939,N_15188,N_15349);
or U15940 (N_15940,N_15399,N_15304);
nand U15941 (N_15941,N_15020,N_15059);
nor U15942 (N_15942,N_15456,N_15271);
xnor U15943 (N_15943,N_15059,N_15222);
nand U15944 (N_15944,N_15041,N_15229);
and U15945 (N_15945,N_15022,N_15191);
or U15946 (N_15946,N_15418,N_15357);
nor U15947 (N_15947,N_15189,N_15322);
xor U15948 (N_15948,N_15464,N_15203);
and U15949 (N_15949,N_15286,N_15320);
nor U15950 (N_15950,N_15294,N_15357);
or U15951 (N_15951,N_15108,N_15325);
xor U15952 (N_15952,N_15032,N_15119);
nor U15953 (N_15953,N_15286,N_15206);
xor U15954 (N_15954,N_15271,N_15243);
xnor U15955 (N_15955,N_15164,N_15235);
nand U15956 (N_15956,N_15289,N_15318);
nor U15957 (N_15957,N_15336,N_15062);
or U15958 (N_15958,N_15466,N_15435);
nand U15959 (N_15959,N_15121,N_15254);
and U15960 (N_15960,N_15480,N_15347);
xnor U15961 (N_15961,N_15499,N_15267);
xnor U15962 (N_15962,N_15382,N_15384);
nand U15963 (N_15963,N_15171,N_15017);
or U15964 (N_15964,N_15230,N_15257);
and U15965 (N_15965,N_15052,N_15143);
or U15966 (N_15966,N_15217,N_15054);
or U15967 (N_15967,N_15228,N_15033);
nand U15968 (N_15968,N_15314,N_15363);
or U15969 (N_15969,N_15408,N_15447);
nand U15970 (N_15970,N_15360,N_15082);
nand U15971 (N_15971,N_15170,N_15455);
and U15972 (N_15972,N_15114,N_15259);
nand U15973 (N_15973,N_15273,N_15442);
nor U15974 (N_15974,N_15487,N_15136);
nand U15975 (N_15975,N_15409,N_15168);
xnor U15976 (N_15976,N_15426,N_15473);
xnor U15977 (N_15977,N_15128,N_15021);
xor U15978 (N_15978,N_15020,N_15093);
nor U15979 (N_15979,N_15201,N_15230);
xnor U15980 (N_15980,N_15163,N_15320);
xnor U15981 (N_15981,N_15267,N_15216);
or U15982 (N_15982,N_15232,N_15156);
xor U15983 (N_15983,N_15261,N_15427);
nor U15984 (N_15984,N_15018,N_15096);
nor U15985 (N_15985,N_15099,N_15187);
nor U15986 (N_15986,N_15494,N_15264);
and U15987 (N_15987,N_15405,N_15343);
nor U15988 (N_15988,N_15155,N_15407);
nand U15989 (N_15989,N_15313,N_15182);
and U15990 (N_15990,N_15383,N_15062);
or U15991 (N_15991,N_15479,N_15044);
xor U15992 (N_15992,N_15487,N_15005);
nand U15993 (N_15993,N_15230,N_15075);
nand U15994 (N_15994,N_15199,N_15498);
nor U15995 (N_15995,N_15289,N_15097);
nand U15996 (N_15996,N_15140,N_15087);
nand U15997 (N_15997,N_15325,N_15344);
and U15998 (N_15998,N_15280,N_15469);
or U15999 (N_15999,N_15103,N_15065);
nor U16000 (N_16000,N_15869,N_15662);
nand U16001 (N_16001,N_15649,N_15983);
or U16002 (N_16002,N_15767,N_15504);
xnor U16003 (N_16003,N_15912,N_15924);
nand U16004 (N_16004,N_15974,N_15503);
nand U16005 (N_16005,N_15551,N_15535);
nand U16006 (N_16006,N_15772,N_15773);
nand U16007 (N_16007,N_15698,N_15886);
and U16008 (N_16008,N_15899,N_15600);
and U16009 (N_16009,N_15804,N_15521);
or U16010 (N_16010,N_15618,N_15671);
xor U16011 (N_16011,N_15669,N_15505);
nor U16012 (N_16012,N_15811,N_15839);
or U16013 (N_16013,N_15708,N_15980);
nor U16014 (N_16014,N_15949,N_15776);
xor U16015 (N_16015,N_15881,N_15620);
or U16016 (N_16016,N_15900,N_15780);
nand U16017 (N_16017,N_15583,N_15532);
or U16018 (N_16018,N_15829,N_15511);
or U16019 (N_16019,N_15754,N_15865);
or U16020 (N_16020,N_15691,N_15724);
xor U16021 (N_16021,N_15922,N_15768);
or U16022 (N_16022,N_15760,N_15591);
and U16023 (N_16023,N_15727,N_15947);
and U16024 (N_16024,N_15586,N_15707);
and U16025 (N_16025,N_15634,N_15676);
nand U16026 (N_16026,N_15651,N_15918);
xor U16027 (N_16027,N_15779,N_15571);
or U16028 (N_16028,N_15866,N_15642);
and U16029 (N_16029,N_15904,N_15606);
nand U16030 (N_16030,N_15737,N_15955);
and U16031 (N_16031,N_15952,N_15820);
xnor U16032 (N_16032,N_15761,N_15797);
xnor U16033 (N_16033,N_15850,N_15720);
nand U16034 (N_16034,N_15643,N_15531);
xor U16035 (N_16035,N_15810,N_15885);
nand U16036 (N_16036,N_15646,N_15517);
or U16037 (N_16037,N_15915,N_15515);
and U16038 (N_16038,N_15694,N_15553);
and U16039 (N_16039,N_15965,N_15624);
nor U16040 (N_16040,N_15543,N_15856);
nor U16041 (N_16041,N_15589,N_15700);
xor U16042 (N_16042,N_15680,N_15858);
and U16043 (N_16043,N_15805,N_15750);
nor U16044 (N_16044,N_15587,N_15725);
xnor U16045 (N_16045,N_15681,N_15665);
xnor U16046 (N_16046,N_15911,N_15738);
nor U16047 (N_16047,N_15684,N_15925);
nand U16048 (N_16048,N_15972,N_15635);
xnor U16049 (N_16049,N_15894,N_15860);
nand U16050 (N_16050,N_15568,N_15507);
nor U16051 (N_16051,N_15823,N_15537);
nor U16052 (N_16052,N_15841,N_15909);
or U16053 (N_16053,N_15863,N_15844);
or U16054 (N_16054,N_15943,N_15895);
and U16055 (N_16055,N_15873,N_15978);
xor U16056 (N_16056,N_15514,N_15633);
and U16057 (N_16057,N_15740,N_15661);
xnor U16058 (N_16058,N_15644,N_15993);
xnor U16059 (N_16059,N_15968,N_15812);
xor U16060 (N_16060,N_15647,N_15546);
nor U16061 (N_16061,N_15867,N_15991);
or U16062 (N_16062,N_15948,N_15941);
xor U16063 (N_16063,N_15673,N_15808);
and U16064 (N_16064,N_15963,N_15853);
nand U16065 (N_16065,N_15982,N_15852);
nand U16066 (N_16066,N_15891,N_15574);
and U16067 (N_16067,N_15871,N_15641);
nor U16068 (N_16068,N_15552,N_15913);
xnor U16069 (N_16069,N_15747,N_15752);
or U16070 (N_16070,N_15981,N_15908);
xor U16071 (N_16071,N_15775,N_15687);
xnor U16072 (N_16072,N_15920,N_15778);
and U16073 (N_16073,N_15755,N_15903);
nor U16074 (N_16074,N_15813,N_15715);
nor U16075 (N_16075,N_15872,N_15790);
nor U16076 (N_16076,N_15741,N_15598);
or U16077 (N_16077,N_15988,N_15959);
xnor U16078 (N_16078,N_15544,N_15529);
or U16079 (N_16079,N_15976,N_15857);
nand U16080 (N_16080,N_15622,N_15549);
and U16081 (N_16081,N_15827,N_15842);
nor U16082 (N_16082,N_15845,N_15876);
nand U16083 (N_16083,N_15714,N_15659);
or U16084 (N_16084,N_15621,N_15927);
or U16085 (N_16085,N_15705,N_15601);
xor U16086 (N_16086,N_15854,N_15806);
nand U16087 (N_16087,N_15519,N_15682);
and U16088 (N_16088,N_15807,N_15884);
or U16089 (N_16089,N_15907,N_15935);
nand U16090 (N_16090,N_15558,N_15967);
nor U16091 (N_16091,N_15512,N_15603);
or U16092 (N_16092,N_15625,N_15964);
or U16093 (N_16093,N_15631,N_15992);
nor U16094 (N_16094,N_15939,N_15575);
or U16095 (N_16095,N_15652,N_15926);
or U16096 (N_16096,N_15674,N_15545);
nor U16097 (N_16097,N_15605,N_15914);
xnor U16098 (N_16098,N_15809,N_15655);
nor U16099 (N_16099,N_15999,N_15675);
nor U16100 (N_16100,N_15510,N_15688);
and U16101 (N_16101,N_15679,N_15516);
and U16102 (N_16102,N_15934,N_15580);
nor U16103 (N_16103,N_15716,N_15710);
xor U16104 (N_16104,N_15609,N_15613);
nand U16105 (N_16105,N_15706,N_15821);
nor U16106 (N_16106,N_15728,N_15938);
or U16107 (N_16107,N_15946,N_15771);
nor U16108 (N_16108,N_15759,N_15793);
xnor U16109 (N_16109,N_15763,N_15578);
and U16110 (N_16110,N_15711,N_15629);
nor U16111 (N_16111,N_15801,N_15843);
nand U16112 (N_16112,N_15632,N_15897);
xor U16113 (N_16113,N_15721,N_15880);
xnor U16114 (N_16114,N_15830,N_15803);
or U16115 (N_16115,N_15561,N_15640);
nor U16116 (N_16116,N_15971,N_15685);
and U16117 (N_16117,N_15704,N_15630);
xor U16118 (N_16118,N_15822,N_15798);
and U16119 (N_16119,N_15861,N_15563);
and U16120 (N_16120,N_15937,N_15882);
nor U16121 (N_16121,N_15953,N_15672);
xor U16122 (N_16122,N_15814,N_15743);
nor U16123 (N_16123,N_15757,N_15815);
nor U16124 (N_16124,N_15696,N_15792);
or U16125 (N_16125,N_15910,N_15520);
or U16126 (N_16126,N_15870,N_15732);
xnor U16127 (N_16127,N_15594,N_15559);
or U16128 (N_16128,N_15678,N_15851);
xnor U16129 (N_16129,N_15736,N_15683);
nand U16130 (N_16130,N_15787,N_15539);
nand U16131 (N_16131,N_15824,N_15526);
nor U16132 (N_16132,N_15500,N_15942);
xor U16133 (N_16133,N_15735,N_15612);
or U16134 (N_16134,N_15628,N_15764);
or U16135 (N_16135,N_15686,N_15785);
or U16136 (N_16136,N_15693,N_15921);
or U16137 (N_16137,N_15833,N_15957);
or U16138 (N_16138,N_15931,N_15695);
and U16139 (N_16139,N_15906,N_15523);
nand U16140 (N_16140,N_15566,N_15794);
nand U16141 (N_16141,N_15542,N_15653);
xor U16142 (N_16142,N_15940,N_15670);
nor U16143 (N_16143,N_15874,N_15608);
nand U16144 (N_16144,N_15969,N_15987);
nor U16145 (N_16145,N_15569,N_15723);
nand U16146 (N_16146,N_15834,N_15905);
and U16147 (N_16147,N_15506,N_15994);
nand U16148 (N_16148,N_15555,N_15998);
and U16149 (N_16149,N_15928,N_15799);
or U16150 (N_16150,N_15557,N_15956);
nand U16151 (N_16151,N_15560,N_15954);
or U16152 (N_16152,N_15567,N_15637);
or U16153 (N_16153,N_15595,N_15879);
and U16154 (N_16154,N_15590,N_15883);
and U16155 (N_16155,N_15789,N_15795);
nand U16156 (N_16156,N_15864,N_15958);
xnor U16157 (N_16157,N_15933,N_15565);
nor U16158 (N_16158,N_15547,N_15975);
nor U16159 (N_16159,N_15733,N_15656);
xor U16160 (N_16160,N_15533,N_15770);
and U16161 (N_16161,N_15997,N_15826);
xor U16162 (N_16162,N_15709,N_15689);
xor U16163 (N_16163,N_15611,N_15577);
nor U16164 (N_16164,N_15862,N_15846);
nor U16165 (N_16165,N_15917,N_15731);
nand U16166 (N_16166,N_15753,N_15658);
and U16167 (N_16167,N_15663,N_15745);
nor U16168 (N_16168,N_15849,N_15916);
xnor U16169 (N_16169,N_15848,N_15718);
or U16170 (N_16170,N_15888,N_15627);
nor U16171 (N_16171,N_15588,N_15893);
nand U16172 (N_16172,N_15828,N_15668);
or U16173 (N_16173,N_15751,N_15717);
or U16174 (N_16174,N_15746,N_15945);
xnor U16175 (N_16175,N_15638,N_15832);
nand U16176 (N_16176,N_15701,N_15944);
and U16177 (N_16177,N_15889,N_15734);
xnor U16178 (N_16178,N_15722,N_15744);
xnor U16179 (N_16179,N_15781,N_15599);
nand U16180 (N_16180,N_15703,N_15784);
and U16181 (N_16181,N_15749,N_15576);
nor U16182 (N_16182,N_15616,N_15585);
or U16183 (N_16183,N_15847,N_15530);
nor U16184 (N_16184,N_15648,N_15667);
xnor U16185 (N_16185,N_15742,N_15713);
and U16186 (N_16186,N_15617,N_15645);
nand U16187 (N_16187,N_15766,N_15892);
or U16188 (N_16188,N_15636,N_15730);
or U16189 (N_16189,N_15973,N_15548);
nor U16190 (N_16190,N_15901,N_15786);
nor U16191 (N_16191,N_15825,N_15623);
nand U16192 (N_16192,N_15739,N_15509);
nor U16193 (N_16193,N_15898,N_15769);
or U16194 (N_16194,N_15619,N_15887);
xnor U16195 (N_16195,N_15541,N_15697);
nor U16196 (N_16196,N_15932,N_15783);
nand U16197 (N_16197,N_15877,N_15534);
nand U16198 (N_16198,N_15602,N_15513);
and U16199 (N_16199,N_15719,N_15923);
or U16200 (N_16200,N_15614,N_15582);
nand U16201 (N_16201,N_15748,N_15782);
xnor U16202 (N_16202,N_15584,N_15835);
nand U16203 (N_16203,N_15989,N_15816);
xor U16204 (N_16204,N_15831,N_15536);
or U16205 (N_16205,N_15572,N_15800);
or U16206 (N_16206,N_15984,N_15593);
or U16207 (N_16207,N_15970,N_15607);
nor U16208 (N_16208,N_15936,N_15528);
and U16209 (N_16209,N_15579,N_15657);
xor U16210 (N_16210,N_15859,N_15878);
xnor U16211 (N_16211,N_15837,N_15525);
and U16212 (N_16212,N_15666,N_15996);
xor U16213 (N_16213,N_15985,N_15758);
nand U16214 (N_16214,N_15501,N_15690);
nor U16215 (N_16215,N_15699,N_15977);
and U16216 (N_16216,N_15902,N_15951);
xor U16217 (N_16217,N_15639,N_15610);
nor U16218 (N_16218,N_15819,N_15990);
xor U16219 (N_16219,N_15664,N_15929);
and U16220 (N_16220,N_15960,N_15592);
xor U16221 (N_16221,N_15777,N_15838);
or U16222 (N_16222,N_15524,N_15712);
nor U16223 (N_16223,N_15791,N_15729);
nor U16224 (N_16224,N_15508,N_15660);
nor U16225 (N_16225,N_15527,N_15756);
nand U16226 (N_16226,N_15961,N_15765);
and U16227 (N_16227,N_15522,N_15836);
xor U16228 (N_16228,N_15562,N_15597);
nor U16229 (N_16229,N_15788,N_15995);
nand U16230 (N_16230,N_15919,N_15518);
nand U16231 (N_16231,N_15540,N_15986);
nand U16232 (N_16232,N_15570,N_15502);
or U16233 (N_16233,N_15615,N_15950);
or U16234 (N_16234,N_15604,N_15890);
nor U16235 (N_16235,N_15550,N_15581);
or U16236 (N_16236,N_15868,N_15677);
nand U16237 (N_16237,N_15726,N_15650);
and U16238 (N_16238,N_15692,N_15840);
or U16239 (N_16239,N_15875,N_15979);
nor U16240 (N_16240,N_15564,N_15896);
nand U16241 (N_16241,N_15818,N_15774);
nor U16242 (N_16242,N_15796,N_15702);
xnor U16243 (N_16243,N_15962,N_15573);
nor U16244 (N_16244,N_15930,N_15966);
and U16245 (N_16245,N_15554,N_15855);
and U16246 (N_16246,N_15626,N_15762);
or U16247 (N_16247,N_15817,N_15556);
or U16248 (N_16248,N_15538,N_15596);
nand U16249 (N_16249,N_15654,N_15802);
nand U16250 (N_16250,N_15792,N_15732);
or U16251 (N_16251,N_15988,N_15599);
and U16252 (N_16252,N_15538,N_15669);
or U16253 (N_16253,N_15651,N_15615);
and U16254 (N_16254,N_15935,N_15986);
or U16255 (N_16255,N_15563,N_15993);
nor U16256 (N_16256,N_15875,N_15639);
nor U16257 (N_16257,N_15947,N_15572);
and U16258 (N_16258,N_15539,N_15646);
xor U16259 (N_16259,N_15817,N_15543);
nand U16260 (N_16260,N_15744,N_15827);
nand U16261 (N_16261,N_15581,N_15602);
and U16262 (N_16262,N_15658,N_15533);
and U16263 (N_16263,N_15651,N_15585);
and U16264 (N_16264,N_15633,N_15745);
nor U16265 (N_16265,N_15623,N_15518);
nor U16266 (N_16266,N_15755,N_15757);
nand U16267 (N_16267,N_15912,N_15997);
nand U16268 (N_16268,N_15892,N_15531);
nand U16269 (N_16269,N_15841,N_15662);
xnor U16270 (N_16270,N_15623,N_15754);
and U16271 (N_16271,N_15607,N_15772);
xor U16272 (N_16272,N_15678,N_15813);
nor U16273 (N_16273,N_15891,N_15630);
xnor U16274 (N_16274,N_15917,N_15771);
or U16275 (N_16275,N_15685,N_15625);
nand U16276 (N_16276,N_15749,N_15622);
or U16277 (N_16277,N_15559,N_15789);
or U16278 (N_16278,N_15939,N_15928);
and U16279 (N_16279,N_15671,N_15796);
xnor U16280 (N_16280,N_15982,N_15749);
nor U16281 (N_16281,N_15635,N_15706);
xnor U16282 (N_16282,N_15681,N_15789);
or U16283 (N_16283,N_15780,N_15963);
nor U16284 (N_16284,N_15809,N_15564);
nor U16285 (N_16285,N_15655,N_15824);
or U16286 (N_16286,N_15564,N_15947);
xor U16287 (N_16287,N_15606,N_15727);
nand U16288 (N_16288,N_15788,N_15509);
or U16289 (N_16289,N_15857,N_15949);
xnor U16290 (N_16290,N_15673,N_15524);
and U16291 (N_16291,N_15933,N_15899);
and U16292 (N_16292,N_15572,N_15595);
and U16293 (N_16293,N_15700,N_15934);
or U16294 (N_16294,N_15654,N_15919);
nor U16295 (N_16295,N_15785,N_15629);
or U16296 (N_16296,N_15757,N_15675);
nand U16297 (N_16297,N_15836,N_15852);
xor U16298 (N_16298,N_15865,N_15600);
xnor U16299 (N_16299,N_15672,N_15619);
xnor U16300 (N_16300,N_15988,N_15652);
xnor U16301 (N_16301,N_15979,N_15959);
and U16302 (N_16302,N_15658,N_15661);
xnor U16303 (N_16303,N_15916,N_15999);
and U16304 (N_16304,N_15695,N_15728);
nand U16305 (N_16305,N_15742,N_15543);
nor U16306 (N_16306,N_15541,N_15730);
nand U16307 (N_16307,N_15998,N_15885);
and U16308 (N_16308,N_15942,N_15896);
and U16309 (N_16309,N_15745,N_15520);
xnor U16310 (N_16310,N_15979,N_15600);
and U16311 (N_16311,N_15545,N_15778);
xor U16312 (N_16312,N_15716,N_15685);
or U16313 (N_16313,N_15511,N_15833);
or U16314 (N_16314,N_15884,N_15880);
or U16315 (N_16315,N_15759,N_15828);
and U16316 (N_16316,N_15712,N_15724);
xor U16317 (N_16317,N_15943,N_15633);
nand U16318 (N_16318,N_15739,N_15725);
and U16319 (N_16319,N_15843,N_15965);
or U16320 (N_16320,N_15816,N_15827);
and U16321 (N_16321,N_15785,N_15559);
xor U16322 (N_16322,N_15990,N_15709);
or U16323 (N_16323,N_15915,N_15722);
xor U16324 (N_16324,N_15645,N_15608);
nor U16325 (N_16325,N_15665,N_15853);
nor U16326 (N_16326,N_15887,N_15953);
xor U16327 (N_16327,N_15759,N_15523);
or U16328 (N_16328,N_15732,N_15608);
xor U16329 (N_16329,N_15685,N_15983);
and U16330 (N_16330,N_15717,N_15924);
nor U16331 (N_16331,N_15864,N_15504);
nor U16332 (N_16332,N_15926,N_15895);
xor U16333 (N_16333,N_15611,N_15627);
nand U16334 (N_16334,N_15778,N_15658);
nor U16335 (N_16335,N_15902,N_15868);
or U16336 (N_16336,N_15755,N_15696);
nor U16337 (N_16337,N_15570,N_15731);
and U16338 (N_16338,N_15606,N_15589);
or U16339 (N_16339,N_15801,N_15616);
nor U16340 (N_16340,N_15876,N_15747);
nor U16341 (N_16341,N_15829,N_15925);
and U16342 (N_16342,N_15651,N_15702);
and U16343 (N_16343,N_15754,N_15803);
or U16344 (N_16344,N_15725,N_15855);
nand U16345 (N_16345,N_15878,N_15926);
nor U16346 (N_16346,N_15931,N_15898);
nand U16347 (N_16347,N_15590,N_15839);
nand U16348 (N_16348,N_15555,N_15709);
and U16349 (N_16349,N_15672,N_15642);
xnor U16350 (N_16350,N_15848,N_15574);
and U16351 (N_16351,N_15931,N_15759);
xnor U16352 (N_16352,N_15678,N_15938);
and U16353 (N_16353,N_15576,N_15879);
nor U16354 (N_16354,N_15533,N_15521);
or U16355 (N_16355,N_15585,N_15837);
nand U16356 (N_16356,N_15869,N_15558);
xor U16357 (N_16357,N_15712,N_15541);
or U16358 (N_16358,N_15900,N_15611);
and U16359 (N_16359,N_15952,N_15983);
nor U16360 (N_16360,N_15504,N_15841);
or U16361 (N_16361,N_15989,N_15626);
or U16362 (N_16362,N_15865,N_15707);
nand U16363 (N_16363,N_15762,N_15698);
or U16364 (N_16364,N_15786,N_15921);
nor U16365 (N_16365,N_15848,N_15601);
nor U16366 (N_16366,N_15554,N_15775);
nor U16367 (N_16367,N_15836,N_15658);
or U16368 (N_16368,N_15944,N_15509);
or U16369 (N_16369,N_15774,N_15628);
xnor U16370 (N_16370,N_15695,N_15875);
or U16371 (N_16371,N_15657,N_15692);
or U16372 (N_16372,N_15576,N_15811);
and U16373 (N_16373,N_15512,N_15695);
and U16374 (N_16374,N_15988,N_15860);
xnor U16375 (N_16375,N_15972,N_15930);
nor U16376 (N_16376,N_15855,N_15666);
nand U16377 (N_16377,N_15697,N_15696);
nand U16378 (N_16378,N_15597,N_15674);
nand U16379 (N_16379,N_15786,N_15654);
nor U16380 (N_16380,N_15881,N_15872);
or U16381 (N_16381,N_15838,N_15690);
nor U16382 (N_16382,N_15964,N_15658);
nand U16383 (N_16383,N_15952,N_15778);
nand U16384 (N_16384,N_15876,N_15553);
nor U16385 (N_16385,N_15643,N_15672);
nand U16386 (N_16386,N_15727,N_15880);
or U16387 (N_16387,N_15745,N_15662);
and U16388 (N_16388,N_15626,N_15912);
and U16389 (N_16389,N_15902,N_15869);
nor U16390 (N_16390,N_15983,N_15761);
and U16391 (N_16391,N_15512,N_15639);
xnor U16392 (N_16392,N_15884,N_15669);
and U16393 (N_16393,N_15699,N_15723);
or U16394 (N_16394,N_15728,N_15886);
nand U16395 (N_16395,N_15908,N_15550);
or U16396 (N_16396,N_15821,N_15818);
nand U16397 (N_16397,N_15932,N_15822);
nor U16398 (N_16398,N_15781,N_15963);
or U16399 (N_16399,N_15782,N_15801);
nand U16400 (N_16400,N_15561,N_15715);
or U16401 (N_16401,N_15975,N_15889);
nor U16402 (N_16402,N_15572,N_15868);
nand U16403 (N_16403,N_15785,N_15518);
nor U16404 (N_16404,N_15697,N_15819);
or U16405 (N_16405,N_15881,N_15804);
or U16406 (N_16406,N_15896,N_15686);
or U16407 (N_16407,N_15667,N_15975);
xnor U16408 (N_16408,N_15535,N_15896);
xor U16409 (N_16409,N_15922,N_15798);
xor U16410 (N_16410,N_15555,N_15857);
xor U16411 (N_16411,N_15604,N_15955);
and U16412 (N_16412,N_15886,N_15582);
and U16413 (N_16413,N_15760,N_15667);
and U16414 (N_16414,N_15709,N_15713);
xor U16415 (N_16415,N_15870,N_15736);
nand U16416 (N_16416,N_15682,N_15814);
nor U16417 (N_16417,N_15529,N_15812);
nor U16418 (N_16418,N_15965,N_15635);
and U16419 (N_16419,N_15527,N_15615);
nand U16420 (N_16420,N_15510,N_15685);
xor U16421 (N_16421,N_15912,N_15678);
nor U16422 (N_16422,N_15678,N_15977);
xor U16423 (N_16423,N_15681,N_15510);
and U16424 (N_16424,N_15581,N_15780);
or U16425 (N_16425,N_15922,N_15696);
nor U16426 (N_16426,N_15946,N_15878);
nand U16427 (N_16427,N_15821,N_15683);
and U16428 (N_16428,N_15621,N_15603);
or U16429 (N_16429,N_15976,N_15907);
nor U16430 (N_16430,N_15982,N_15506);
or U16431 (N_16431,N_15984,N_15913);
nand U16432 (N_16432,N_15950,N_15825);
nand U16433 (N_16433,N_15666,N_15934);
or U16434 (N_16434,N_15675,N_15804);
or U16435 (N_16435,N_15940,N_15518);
or U16436 (N_16436,N_15610,N_15579);
xnor U16437 (N_16437,N_15650,N_15910);
xor U16438 (N_16438,N_15740,N_15626);
and U16439 (N_16439,N_15681,N_15586);
nand U16440 (N_16440,N_15518,N_15558);
nand U16441 (N_16441,N_15748,N_15554);
or U16442 (N_16442,N_15801,N_15607);
nand U16443 (N_16443,N_15662,N_15880);
and U16444 (N_16444,N_15996,N_15656);
nand U16445 (N_16445,N_15663,N_15871);
and U16446 (N_16446,N_15852,N_15575);
or U16447 (N_16447,N_15623,N_15920);
xnor U16448 (N_16448,N_15704,N_15564);
xnor U16449 (N_16449,N_15786,N_15570);
or U16450 (N_16450,N_15690,N_15851);
nor U16451 (N_16451,N_15746,N_15604);
nand U16452 (N_16452,N_15999,N_15523);
xor U16453 (N_16453,N_15646,N_15744);
nand U16454 (N_16454,N_15546,N_15753);
nand U16455 (N_16455,N_15849,N_15736);
nand U16456 (N_16456,N_15553,N_15688);
and U16457 (N_16457,N_15754,N_15744);
nand U16458 (N_16458,N_15855,N_15867);
nor U16459 (N_16459,N_15936,N_15751);
or U16460 (N_16460,N_15929,N_15660);
and U16461 (N_16461,N_15779,N_15781);
and U16462 (N_16462,N_15731,N_15921);
or U16463 (N_16463,N_15524,N_15858);
nor U16464 (N_16464,N_15627,N_15884);
xnor U16465 (N_16465,N_15932,N_15988);
or U16466 (N_16466,N_15510,N_15923);
nand U16467 (N_16467,N_15979,N_15914);
xor U16468 (N_16468,N_15790,N_15738);
nand U16469 (N_16469,N_15762,N_15509);
nand U16470 (N_16470,N_15687,N_15826);
nand U16471 (N_16471,N_15934,N_15655);
xnor U16472 (N_16472,N_15579,N_15700);
nand U16473 (N_16473,N_15825,N_15911);
xor U16474 (N_16474,N_15789,N_15913);
xnor U16475 (N_16475,N_15574,N_15899);
and U16476 (N_16476,N_15813,N_15868);
and U16477 (N_16477,N_15520,N_15826);
nor U16478 (N_16478,N_15674,N_15681);
or U16479 (N_16479,N_15716,N_15894);
nand U16480 (N_16480,N_15549,N_15598);
xor U16481 (N_16481,N_15656,N_15523);
nor U16482 (N_16482,N_15738,N_15934);
or U16483 (N_16483,N_15638,N_15542);
or U16484 (N_16484,N_15605,N_15827);
nand U16485 (N_16485,N_15893,N_15676);
xnor U16486 (N_16486,N_15845,N_15662);
or U16487 (N_16487,N_15939,N_15974);
and U16488 (N_16488,N_15984,N_15894);
nand U16489 (N_16489,N_15998,N_15923);
nor U16490 (N_16490,N_15697,N_15949);
or U16491 (N_16491,N_15596,N_15856);
and U16492 (N_16492,N_15811,N_15847);
nor U16493 (N_16493,N_15651,N_15658);
nor U16494 (N_16494,N_15912,N_15547);
xor U16495 (N_16495,N_15857,N_15702);
or U16496 (N_16496,N_15550,N_15763);
nand U16497 (N_16497,N_15787,N_15509);
and U16498 (N_16498,N_15812,N_15575);
and U16499 (N_16499,N_15619,N_15676);
xor U16500 (N_16500,N_16077,N_16394);
or U16501 (N_16501,N_16109,N_16432);
xnor U16502 (N_16502,N_16067,N_16392);
nor U16503 (N_16503,N_16453,N_16466);
or U16504 (N_16504,N_16039,N_16018);
or U16505 (N_16505,N_16162,N_16324);
or U16506 (N_16506,N_16342,N_16002);
nor U16507 (N_16507,N_16448,N_16033);
nor U16508 (N_16508,N_16118,N_16477);
xor U16509 (N_16509,N_16371,N_16104);
or U16510 (N_16510,N_16182,N_16016);
nand U16511 (N_16511,N_16210,N_16485);
xor U16512 (N_16512,N_16377,N_16256);
or U16513 (N_16513,N_16006,N_16278);
and U16514 (N_16514,N_16131,N_16156);
xor U16515 (N_16515,N_16396,N_16232);
nor U16516 (N_16516,N_16456,N_16017);
or U16517 (N_16517,N_16151,N_16034);
nand U16518 (N_16518,N_16395,N_16042);
or U16519 (N_16519,N_16132,N_16273);
nand U16520 (N_16520,N_16025,N_16455);
nand U16521 (N_16521,N_16023,N_16199);
nor U16522 (N_16522,N_16462,N_16242);
xor U16523 (N_16523,N_16435,N_16046);
or U16524 (N_16524,N_16114,N_16476);
xor U16525 (N_16525,N_16133,N_16063);
nand U16526 (N_16526,N_16478,N_16010);
nor U16527 (N_16527,N_16458,N_16145);
and U16528 (N_16528,N_16467,N_16030);
nand U16529 (N_16529,N_16051,N_16292);
xor U16530 (N_16530,N_16386,N_16139);
or U16531 (N_16531,N_16321,N_16027);
nand U16532 (N_16532,N_16106,N_16289);
or U16533 (N_16533,N_16360,N_16098);
xor U16534 (N_16534,N_16147,N_16347);
and U16535 (N_16535,N_16446,N_16438);
nor U16536 (N_16536,N_16004,N_16171);
nor U16537 (N_16537,N_16247,N_16142);
or U16538 (N_16538,N_16208,N_16239);
nor U16539 (N_16539,N_16263,N_16196);
nor U16540 (N_16540,N_16425,N_16172);
nand U16541 (N_16541,N_16301,N_16419);
and U16542 (N_16542,N_16329,N_16452);
xor U16543 (N_16543,N_16358,N_16188);
and U16544 (N_16544,N_16314,N_16400);
and U16545 (N_16545,N_16113,N_16009);
nand U16546 (N_16546,N_16164,N_16416);
nor U16547 (N_16547,N_16097,N_16311);
xnor U16548 (N_16548,N_16473,N_16101);
and U16549 (N_16549,N_16436,N_16262);
nor U16550 (N_16550,N_16045,N_16043);
nand U16551 (N_16551,N_16074,N_16176);
xor U16552 (N_16552,N_16417,N_16235);
or U16553 (N_16553,N_16120,N_16433);
or U16554 (N_16554,N_16424,N_16261);
or U16555 (N_16555,N_16225,N_16241);
nor U16556 (N_16556,N_16308,N_16090);
nor U16557 (N_16557,N_16193,N_16204);
nor U16558 (N_16558,N_16355,N_16335);
nor U16559 (N_16559,N_16079,N_16069);
nor U16560 (N_16560,N_16306,N_16212);
or U16561 (N_16561,N_16330,N_16431);
nand U16562 (N_16562,N_16294,N_16245);
nand U16563 (N_16563,N_16169,N_16073);
or U16564 (N_16564,N_16270,N_16222);
xnor U16565 (N_16565,N_16076,N_16299);
and U16566 (N_16566,N_16056,N_16482);
or U16567 (N_16567,N_16055,N_16460);
nor U16568 (N_16568,N_16237,N_16205);
or U16569 (N_16569,N_16489,N_16298);
or U16570 (N_16570,N_16325,N_16170);
nand U16571 (N_16571,N_16334,N_16108);
nand U16572 (N_16572,N_16402,N_16226);
or U16573 (N_16573,N_16457,N_16344);
xor U16574 (N_16574,N_16154,N_16498);
or U16575 (N_16575,N_16026,N_16326);
and U16576 (N_16576,N_16061,N_16340);
xor U16577 (N_16577,N_16060,N_16373);
or U16578 (N_16578,N_16053,N_16412);
nand U16579 (N_16579,N_16072,N_16385);
nor U16580 (N_16580,N_16008,N_16494);
nand U16581 (N_16581,N_16096,N_16185);
and U16582 (N_16582,N_16336,N_16166);
and U16583 (N_16583,N_16341,N_16014);
nand U16584 (N_16584,N_16338,N_16231);
nor U16585 (N_16585,N_16389,N_16150);
nor U16586 (N_16586,N_16037,N_16024);
nand U16587 (N_16587,N_16062,N_16200);
xnor U16588 (N_16588,N_16219,N_16066);
xor U16589 (N_16589,N_16266,N_16493);
or U16590 (N_16590,N_16442,N_16190);
xor U16591 (N_16591,N_16174,N_16252);
and U16592 (N_16592,N_16345,N_16092);
or U16593 (N_16593,N_16369,N_16091);
nor U16594 (N_16594,N_16243,N_16257);
and U16595 (N_16595,N_16209,N_16071);
xor U16596 (N_16596,N_16420,N_16070);
nand U16597 (N_16597,N_16454,N_16475);
nand U16598 (N_16598,N_16168,N_16192);
xor U16599 (N_16599,N_16286,N_16487);
nand U16600 (N_16600,N_16302,N_16268);
nand U16601 (N_16601,N_16028,N_16313);
xor U16602 (N_16602,N_16418,N_16280);
nand U16603 (N_16603,N_16215,N_16233);
nor U16604 (N_16604,N_16359,N_16496);
nor U16605 (N_16605,N_16491,N_16187);
and U16606 (N_16606,N_16178,N_16000);
nand U16607 (N_16607,N_16474,N_16123);
nor U16608 (N_16608,N_16288,N_16103);
and U16609 (N_16609,N_16372,N_16332);
and U16610 (N_16610,N_16155,N_16181);
or U16611 (N_16611,N_16381,N_16451);
xnor U16612 (N_16612,N_16364,N_16281);
nor U16613 (N_16613,N_16031,N_16144);
nand U16614 (N_16614,N_16349,N_16234);
or U16615 (N_16615,N_16022,N_16001);
nor U16616 (N_16616,N_16309,N_16259);
xor U16617 (N_16617,N_16230,N_16497);
nand U16618 (N_16618,N_16414,N_16366);
xor U16619 (N_16619,N_16320,N_16003);
nand U16620 (N_16620,N_16216,N_16111);
nor U16621 (N_16621,N_16032,N_16152);
nor U16622 (N_16622,N_16180,N_16058);
nand U16623 (N_16623,N_16323,N_16107);
nor U16624 (N_16624,N_16064,N_16253);
nand U16625 (N_16625,N_16175,N_16183);
nor U16626 (N_16626,N_16469,N_16319);
or U16627 (N_16627,N_16422,N_16057);
nor U16628 (N_16628,N_16227,N_16430);
xor U16629 (N_16629,N_16429,N_16282);
or U16630 (N_16630,N_16272,N_16005);
xnor U16631 (N_16631,N_16088,N_16054);
nand U16632 (N_16632,N_16179,N_16129);
nor U16633 (N_16633,N_16439,N_16383);
nand U16634 (N_16634,N_16224,N_16189);
and U16635 (N_16635,N_16084,N_16110);
nor U16636 (N_16636,N_16015,N_16221);
and U16637 (N_16637,N_16038,N_16143);
nand U16638 (N_16638,N_16305,N_16117);
and U16639 (N_16639,N_16102,N_16165);
nand U16640 (N_16640,N_16351,N_16036);
and U16641 (N_16641,N_16040,N_16213);
nand U16642 (N_16642,N_16413,N_16303);
and U16643 (N_16643,N_16246,N_16206);
xor U16644 (N_16644,N_16228,N_16134);
nand U16645 (N_16645,N_16379,N_16406);
nor U16646 (N_16646,N_16408,N_16007);
and U16647 (N_16647,N_16148,N_16285);
or U16648 (N_16648,N_16440,N_16483);
or U16649 (N_16649,N_16094,N_16378);
nand U16650 (N_16650,N_16128,N_16409);
or U16651 (N_16651,N_16295,N_16390);
or U16652 (N_16652,N_16068,N_16130);
xor U16653 (N_16653,N_16201,N_16158);
nand U16654 (N_16654,N_16443,N_16217);
nand U16655 (N_16655,N_16488,N_16307);
nand U16656 (N_16656,N_16121,N_16157);
and U16657 (N_16657,N_16153,N_16059);
or U16658 (N_16658,N_16447,N_16315);
xor U16659 (N_16659,N_16095,N_16141);
and U16660 (N_16660,N_16461,N_16251);
xor U16661 (N_16661,N_16019,N_16397);
and U16662 (N_16662,N_16258,N_16481);
and U16663 (N_16663,N_16391,N_16207);
xor U16664 (N_16664,N_16011,N_16480);
and U16665 (N_16665,N_16177,N_16255);
and U16666 (N_16666,N_16211,N_16124);
or U16667 (N_16667,N_16140,N_16125);
or U16668 (N_16668,N_16099,N_16339);
or U16669 (N_16669,N_16322,N_16353);
nor U16670 (N_16670,N_16052,N_16290);
xnor U16671 (N_16671,N_16279,N_16248);
nor U16672 (N_16672,N_16087,N_16184);
and U16673 (N_16673,N_16472,N_16310);
and U16674 (N_16674,N_16410,N_16161);
nor U16675 (N_16675,N_16387,N_16384);
or U16676 (N_16676,N_16499,N_16044);
nand U16677 (N_16677,N_16049,N_16393);
nand U16678 (N_16678,N_16312,N_16444);
xnor U16679 (N_16679,N_16159,N_16367);
xnor U16680 (N_16680,N_16464,N_16405);
and U16681 (N_16681,N_16013,N_16236);
nor U16682 (N_16682,N_16361,N_16403);
and U16683 (N_16683,N_16267,N_16115);
or U16684 (N_16684,N_16459,N_16283);
or U16685 (N_16685,N_16297,N_16202);
and U16686 (N_16686,N_16160,N_16085);
and U16687 (N_16687,N_16012,N_16250);
nor U16688 (N_16688,N_16375,N_16317);
nor U16689 (N_16689,N_16354,N_16421);
xnor U16690 (N_16690,N_16388,N_16050);
xnor U16691 (N_16691,N_16470,N_16083);
xor U16692 (N_16692,N_16249,N_16362);
nor U16693 (N_16693,N_16214,N_16471);
xnor U16694 (N_16694,N_16137,N_16490);
and U16695 (N_16695,N_16116,N_16437);
nor U16696 (N_16696,N_16407,N_16374);
nor U16697 (N_16697,N_16218,N_16122);
or U16698 (N_16698,N_16275,N_16398);
nor U16699 (N_16699,N_16352,N_16449);
or U16700 (N_16700,N_16434,N_16203);
and U16701 (N_16701,N_16260,N_16086);
nand U16702 (N_16702,N_16399,N_16463);
nand U16703 (N_16703,N_16484,N_16304);
and U16704 (N_16704,N_16357,N_16271);
or U16705 (N_16705,N_16146,N_16426);
and U16706 (N_16706,N_16041,N_16065);
xnor U16707 (N_16707,N_16495,N_16441);
nor U16708 (N_16708,N_16316,N_16277);
nor U16709 (N_16709,N_16195,N_16229);
nor U16710 (N_16710,N_16082,N_16376);
xnor U16711 (N_16711,N_16254,N_16293);
and U16712 (N_16712,N_16479,N_16080);
and U16713 (N_16713,N_16445,N_16328);
nand U16714 (N_16714,N_16138,N_16365);
nor U16715 (N_16715,N_16173,N_16284);
and U16716 (N_16716,N_16136,N_16370);
xnor U16717 (N_16717,N_16105,N_16404);
nand U16718 (N_16718,N_16428,N_16382);
and U16719 (N_16719,N_16331,N_16346);
and U16720 (N_16720,N_16112,N_16135);
and U16721 (N_16721,N_16291,N_16265);
and U16722 (N_16722,N_16198,N_16240);
nor U16723 (N_16723,N_16274,N_16296);
xor U16724 (N_16724,N_16411,N_16380);
xnor U16725 (N_16725,N_16100,N_16167);
and U16726 (N_16726,N_16149,N_16415);
and U16727 (N_16727,N_16075,N_16081);
nor U16728 (N_16728,N_16078,N_16465);
nand U16729 (N_16729,N_16350,N_16029);
or U16730 (N_16730,N_16468,N_16348);
or U16731 (N_16731,N_16423,N_16191);
xnor U16732 (N_16732,N_16450,N_16093);
nor U16733 (N_16733,N_16492,N_16089);
nand U16734 (N_16734,N_16300,N_16337);
or U16735 (N_16735,N_16368,N_16238);
or U16736 (N_16736,N_16269,N_16427);
and U16737 (N_16737,N_16333,N_16035);
nor U16738 (N_16738,N_16048,N_16327);
nand U16739 (N_16739,N_16021,N_16486);
and U16740 (N_16740,N_16194,N_16047);
nand U16741 (N_16741,N_16220,N_16186);
or U16742 (N_16742,N_16223,N_16276);
nand U16743 (N_16743,N_16401,N_16126);
and U16744 (N_16744,N_16244,N_16163);
nand U16745 (N_16745,N_16119,N_16020);
xor U16746 (N_16746,N_16287,N_16363);
nor U16747 (N_16747,N_16318,N_16264);
nor U16748 (N_16748,N_16356,N_16343);
nand U16749 (N_16749,N_16127,N_16197);
and U16750 (N_16750,N_16306,N_16407);
xor U16751 (N_16751,N_16161,N_16279);
nand U16752 (N_16752,N_16113,N_16136);
and U16753 (N_16753,N_16403,N_16150);
nand U16754 (N_16754,N_16207,N_16451);
xnor U16755 (N_16755,N_16142,N_16089);
xor U16756 (N_16756,N_16399,N_16466);
nor U16757 (N_16757,N_16270,N_16183);
nor U16758 (N_16758,N_16381,N_16207);
xor U16759 (N_16759,N_16301,N_16052);
nor U16760 (N_16760,N_16432,N_16317);
nor U16761 (N_16761,N_16433,N_16366);
nor U16762 (N_16762,N_16322,N_16276);
and U16763 (N_16763,N_16397,N_16231);
or U16764 (N_16764,N_16400,N_16309);
xnor U16765 (N_16765,N_16033,N_16350);
or U16766 (N_16766,N_16111,N_16290);
nor U16767 (N_16767,N_16214,N_16094);
xnor U16768 (N_16768,N_16334,N_16430);
or U16769 (N_16769,N_16273,N_16307);
nor U16770 (N_16770,N_16246,N_16437);
nor U16771 (N_16771,N_16196,N_16382);
xnor U16772 (N_16772,N_16233,N_16297);
xor U16773 (N_16773,N_16377,N_16097);
and U16774 (N_16774,N_16210,N_16455);
nor U16775 (N_16775,N_16317,N_16443);
or U16776 (N_16776,N_16191,N_16363);
xor U16777 (N_16777,N_16048,N_16487);
or U16778 (N_16778,N_16207,N_16067);
nand U16779 (N_16779,N_16392,N_16419);
and U16780 (N_16780,N_16342,N_16231);
or U16781 (N_16781,N_16393,N_16050);
xnor U16782 (N_16782,N_16045,N_16055);
or U16783 (N_16783,N_16492,N_16186);
and U16784 (N_16784,N_16112,N_16280);
xnor U16785 (N_16785,N_16485,N_16218);
or U16786 (N_16786,N_16225,N_16417);
xnor U16787 (N_16787,N_16163,N_16452);
or U16788 (N_16788,N_16445,N_16137);
and U16789 (N_16789,N_16321,N_16460);
and U16790 (N_16790,N_16231,N_16138);
or U16791 (N_16791,N_16107,N_16268);
xor U16792 (N_16792,N_16430,N_16456);
xor U16793 (N_16793,N_16468,N_16074);
or U16794 (N_16794,N_16189,N_16219);
and U16795 (N_16795,N_16085,N_16142);
xor U16796 (N_16796,N_16119,N_16428);
xnor U16797 (N_16797,N_16203,N_16101);
nand U16798 (N_16798,N_16022,N_16272);
nand U16799 (N_16799,N_16096,N_16135);
nor U16800 (N_16800,N_16254,N_16379);
xnor U16801 (N_16801,N_16472,N_16443);
nor U16802 (N_16802,N_16483,N_16044);
or U16803 (N_16803,N_16107,N_16074);
nand U16804 (N_16804,N_16086,N_16315);
xnor U16805 (N_16805,N_16381,N_16225);
nand U16806 (N_16806,N_16261,N_16488);
and U16807 (N_16807,N_16202,N_16499);
and U16808 (N_16808,N_16456,N_16296);
or U16809 (N_16809,N_16292,N_16368);
and U16810 (N_16810,N_16114,N_16053);
and U16811 (N_16811,N_16314,N_16331);
and U16812 (N_16812,N_16476,N_16121);
xnor U16813 (N_16813,N_16493,N_16178);
xor U16814 (N_16814,N_16015,N_16037);
or U16815 (N_16815,N_16043,N_16263);
nand U16816 (N_16816,N_16335,N_16320);
or U16817 (N_16817,N_16300,N_16167);
or U16818 (N_16818,N_16419,N_16214);
and U16819 (N_16819,N_16264,N_16295);
nor U16820 (N_16820,N_16329,N_16335);
nor U16821 (N_16821,N_16313,N_16226);
and U16822 (N_16822,N_16148,N_16366);
or U16823 (N_16823,N_16149,N_16445);
and U16824 (N_16824,N_16442,N_16233);
nand U16825 (N_16825,N_16109,N_16368);
nor U16826 (N_16826,N_16042,N_16312);
nor U16827 (N_16827,N_16285,N_16456);
nor U16828 (N_16828,N_16418,N_16090);
nand U16829 (N_16829,N_16245,N_16185);
and U16830 (N_16830,N_16471,N_16279);
xor U16831 (N_16831,N_16303,N_16054);
xnor U16832 (N_16832,N_16098,N_16329);
and U16833 (N_16833,N_16100,N_16393);
xor U16834 (N_16834,N_16364,N_16074);
nor U16835 (N_16835,N_16102,N_16303);
nand U16836 (N_16836,N_16210,N_16057);
xor U16837 (N_16837,N_16424,N_16285);
or U16838 (N_16838,N_16332,N_16091);
and U16839 (N_16839,N_16463,N_16475);
xor U16840 (N_16840,N_16451,N_16230);
or U16841 (N_16841,N_16020,N_16167);
and U16842 (N_16842,N_16437,N_16245);
or U16843 (N_16843,N_16165,N_16209);
and U16844 (N_16844,N_16245,N_16429);
or U16845 (N_16845,N_16069,N_16159);
nor U16846 (N_16846,N_16461,N_16239);
and U16847 (N_16847,N_16109,N_16294);
xor U16848 (N_16848,N_16079,N_16105);
or U16849 (N_16849,N_16060,N_16225);
nor U16850 (N_16850,N_16057,N_16493);
or U16851 (N_16851,N_16459,N_16277);
nor U16852 (N_16852,N_16292,N_16130);
xnor U16853 (N_16853,N_16428,N_16316);
and U16854 (N_16854,N_16363,N_16070);
and U16855 (N_16855,N_16465,N_16379);
and U16856 (N_16856,N_16053,N_16493);
or U16857 (N_16857,N_16046,N_16193);
nand U16858 (N_16858,N_16324,N_16202);
and U16859 (N_16859,N_16212,N_16345);
or U16860 (N_16860,N_16406,N_16092);
and U16861 (N_16861,N_16058,N_16398);
nor U16862 (N_16862,N_16123,N_16389);
xor U16863 (N_16863,N_16240,N_16229);
or U16864 (N_16864,N_16198,N_16491);
nor U16865 (N_16865,N_16454,N_16451);
xor U16866 (N_16866,N_16077,N_16364);
and U16867 (N_16867,N_16287,N_16114);
and U16868 (N_16868,N_16234,N_16486);
nand U16869 (N_16869,N_16277,N_16186);
nor U16870 (N_16870,N_16337,N_16177);
xor U16871 (N_16871,N_16349,N_16169);
xor U16872 (N_16872,N_16061,N_16267);
nand U16873 (N_16873,N_16311,N_16196);
nand U16874 (N_16874,N_16322,N_16131);
nor U16875 (N_16875,N_16428,N_16361);
or U16876 (N_16876,N_16217,N_16380);
nand U16877 (N_16877,N_16033,N_16427);
nand U16878 (N_16878,N_16185,N_16446);
or U16879 (N_16879,N_16161,N_16248);
xnor U16880 (N_16880,N_16285,N_16411);
and U16881 (N_16881,N_16011,N_16411);
and U16882 (N_16882,N_16151,N_16467);
and U16883 (N_16883,N_16283,N_16414);
nand U16884 (N_16884,N_16126,N_16195);
nand U16885 (N_16885,N_16060,N_16140);
xnor U16886 (N_16886,N_16043,N_16315);
xor U16887 (N_16887,N_16107,N_16370);
and U16888 (N_16888,N_16359,N_16125);
nor U16889 (N_16889,N_16350,N_16435);
xnor U16890 (N_16890,N_16131,N_16342);
and U16891 (N_16891,N_16148,N_16486);
or U16892 (N_16892,N_16049,N_16040);
xnor U16893 (N_16893,N_16385,N_16339);
and U16894 (N_16894,N_16221,N_16470);
xnor U16895 (N_16895,N_16335,N_16462);
xor U16896 (N_16896,N_16478,N_16221);
nand U16897 (N_16897,N_16188,N_16380);
and U16898 (N_16898,N_16434,N_16498);
xnor U16899 (N_16899,N_16394,N_16366);
nand U16900 (N_16900,N_16167,N_16290);
nand U16901 (N_16901,N_16464,N_16233);
nor U16902 (N_16902,N_16094,N_16066);
nand U16903 (N_16903,N_16177,N_16409);
or U16904 (N_16904,N_16075,N_16169);
and U16905 (N_16905,N_16175,N_16308);
nand U16906 (N_16906,N_16455,N_16159);
nand U16907 (N_16907,N_16000,N_16076);
nor U16908 (N_16908,N_16171,N_16409);
or U16909 (N_16909,N_16370,N_16132);
and U16910 (N_16910,N_16218,N_16405);
and U16911 (N_16911,N_16161,N_16083);
xnor U16912 (N_16912,N_16117,N_16260);
xnor U16913 (N_16913,N_16061,N_16344);
and U16914 (N_16914,N_16358,N_16466);
or U16915 (N_16915,N_16487,N_16310);
or U16916 (N_16916,N_16052,N_16276);
and U16917 (N_16917,N_16379,N_16069);
or U16918 (N_16918,N_16369,N_16290);
nor U16919 (N_16919,N_16393,N_16070);
nand U16920 (N_16920,N_16317,N_16338);
nor U16921 (N_16921,N_16387,N_16455);
nor U16922 (N_16922,N_16364,N_16098);
xnor U16923 (N_16923,N_16369,N_16039);
or U16924 (N_16924,N_16454,N_16384);
xnor U16925 (N_16925,N_16057,N_16262);
nor U16926 (N_16926,N_16341,N_16016);
nand U16927 (N_16927,N_16386,N_16292);
or U16928 (N_16928,N_16011,N_16203);
and U16929 (N_16929,N_16237,N_16068);
or U16930 (N_16930,N_16376,N_16198);
nor U16931 (N_16931,N_16003,N_16260);
and U16932 (N_16932,N_16048,N_16331);
xor U16933 (N_16933,N_16144,N_16409);
and U16934 (N_16934,N_16469,N_16274);
or U16935 (N_16935,N_16141,N_16300);
or U16936 (N_16936,N_16096,N_16265);
and U16937 (N_16937,N_16207,N_16487);
or U16938 (N_16938,N_16305,N_16329);
or U16939 (N_16939,N_16388,N_16017);
and U16940 (N_16940,N_16441,N_16331);
nor U16941 (N_16941,N_16117,N_16220);
nor U16942 (N_16942,N_16419,N_16220);
xor U16943 (N_16943,N_16161,N_16377);
xnor U16944 (N_16944,N_16193,N_16084);
nor U16945 (N_16945,N_16073,N_16034);
nand U16946 (N_16946,N_16317,N_16391);
and U16947 (N_16947,N_16154,N_16348);
xnor U16948 (N_16948,N_16264,N_16269);
and U16949 (N_16949,N_16370,N_16493);
nor U16950 (N_16950,N_16124,N_16427);
or U16951 (N_16951,N_16358,N_16339);
xor U16952 (N_16952,N_16148,N_16450);
nor U16953 (N_16953,N_16328,N_16270);
xnor U16954 (N_16954,N_16309,N_16192);
xor U16955 (N_16955,N_16327,N_16417);
xor U16956 (N_16956,N_16468,N_16431);
nand U16957 (N_16957,N_16376,N_16462);
or U16958 (N_16958,N_16334,N_16043);
or U16959 (N_16959,N_16497,N_16212);
and U16960 (N_16960,N_16204,N_16053);
and U16961 (N_16961,N_16197,N_16318);
and U16962 (N_16962,N_16196,N_16318);
or U16963 (N_16963,N_16201,N_16430);
nor U16964 (N_16964,N_16282,N_16121);
nand U16965 (N_16965,N_16480,N_16090);
xor U16966 (N_16966,N_16286,N_16351);
nand U16967 (N_16967,N_16432,N_16256);
xor U16968 (N_16968,N_16490,N_16476);
or U16969 (N_16969,N_16381,N_16232);
nor U16970 (N_16970,N_16022,N_16104);
nand U16971 (N_16971,N_16460,N_16497);
and U16972 (N_16972,N_16084,N_16231);
or U16973 (N_16973,N_16252,N_16375);
xnor U16974 (N_16974,N_16442,N_16012);
nand U16975 (N_16975,N_16311,N_16150);
nand U16976 (N_16976,N_16163,N_16286);
or U16977 (N_16977,N_16332,N_16405);
nor U16978 (N_16978,N_16473,N_16180);
or U16979 (N_16979,N_16063,N_16311);
or U16980 (N_16980,N_16474,N_16403);
or U16981 (N_16981,N_16051,N_16066);
or U16982 (N_16982,N_16123,N_16467);
and U16983 (N_16983,N_16424,N_16128);
xnor U16984 (N_16984,N_16069,N_16498);
and U16985 (N_16985,N_16276,N_16264);
nor U16986 (N_16986,N_16306,N_16315);
or U16987 (N_16987,N_16024,N_16010);
and U16988 (N_16988,N_16362,N_16303);
or U16989 (N_16989,N_16393,N_16319);
nand U16990 (N_16990,N_16037,N_16459);
nand U16991 (N_16991,N_16117,N_16318);
nand U16992 (N_16992,N_16170,N_16009);
nor U16993 (N_16993,N_16203,N_16342);
or U16994 (N_16994,N_16412,N_16131);
nand U16995 (N_16995,N_16067,N_16034);
or U16996 (N_16996,N_16387,N_16222);
xor U16997 (N_16997,N_16263,N_16176);
or U16998 (N_16998,N_16425,N_16003);
nor U16999 (N_16999,N_16271,N_16074);
nor U17000 (N_17000,N_16790,N_16849);
or U17001 (N_17001,N_16766,N_16716);
and U17002 (N_17002,N_16811,N_16813);
and U17003 (N_17003,N_16703,N_16587);
or U17004 (N_17004,N_16659,N_16707);
nand U17005 (N_17005,N_16529,N_16897);
nor U17006 (N_17006,N_16691,N_16988);
or U17007 (N_17007,N_16743,N_16965);
or U17008 (N_17008,N_16568,N_16604);
nor U17009 (N_17009,N_16748,N_16530);
and U17010 (N_17010,N_16692,N_16741);
or U17011 (N_17011,N_16963,N_16526);
nand U17012 (N_17012,N_16954,N_16945);
nand U17013 (N_17013,N_16927,N_16991);
nand U17014 (N_17014,N_16599,N_16627);
nand U17015 (N_17015,N_16773,N_16961);
nand U17016 (N_17016,N_16505,N_16630);
or U17017 (N_17017,N_16739,N_16933);
nand U17018 (N_17018,N_16794,N_16888);
nor U17019 (N_17019,N_16767,N_16534);
nor U17020 (N_17020,N_16839,N_16914);
and U17021 (N_17021,N_16779,N_16872);
xnor U17022 (N_17022,N_16871,N_16580);
or U17023 (N_17023,N_16569,N_16738);
nand U17024 (N_17024,N_16972,N_16728);
or U17025 (N_17025,N_16926,N_16996);
nand U17026 (N_17026,N_16917,N_16605);
nand U17027 (N_17027,N_16626,N_16772);
xnor U17028 (N_17028,N_16806,N_16786);
nand U17029 (N_17029,N_16870,N_16575);
or U17030 (N_17030,N_16524,N_16665);
nand U17031 (N_17031,N_16643,N_16859);
or U17032 (N_17032,N_16899,N_16522);
and U17033 (N_17033,N_16845,N_16631);
or U17034 (N_17034,N_16733,N_16782);
nand U17035 (N_17035,N_16902,N_16803);
xor U17036 (N_17036,N_16907,N_16876);
nand U17037 (N_17037,N_16544,N_16590);
or U17038 (N_17038,N_16805,N_16893);
nor U17039 (N_17039,N_16612,N_16636);
nand U17040 (N_17040,N_16969,N_16921);
nor U17041 (N_17041,N_16552,N_16559);
and U17042 (N_17042,N_16622,N_16750);
xor U17043 (N_17043,N_16567,N_16618);
xor U17044 (N_17044,N_16900,N_16621);
nor U17045 (N_17045,N_16638,N_16516);
xor U17046 (N_17046,N_16712,N_16701);
and U17047 (N_17047,N_16539,N_16702);
nand U17048 (N_17048,N_16873,N_16810);
or U17049 (N_17049,N_16573,N_16925);
nor U17050 (N_17050,N_16520,N_16936);
nor U17051 (N_17051,N_16637,N_16721);
nor U17052 (N_17052,N_16841,N_16932);
nand U17053 (N_17053,N_16710,N_16668);
xnor U17054 (N_17054,N_16912,N_16864);
nand U17055 (N_17055,N_16800,N_16856);
nor U17056 (N_17056,N_16950,N_16753);
nand U17057 (N_17057,N_16827,N_16549);
xnor U17058 (N_17058,N_16862,N_16960);
nand U17059 (N_17059,N_16765,N_16828);
nand U17060 (N_17060,N_16832,N_16635);
xnor U17061 (N_17061,N_16910,N_16880);
and U17062 (N_17062,N_16584,N_16746);
or U17063 (N_17063,N_16901,N_16656);
and U17064 (N_17064,N_16601,N_16628);
xor U17065 (N_17065,N_16595,N_16589);
nor U17066 (N_17066,N_16690,N_16672);
nor U17067 (N_17067,N_16970,N_16787);
nor U17068 (N_17068,N_16578,N_16648);
xnor U17069 (N_17069,N_16642,N_16557);
and U17070 (N_17070,N_16756,N_16998);
or U17071 (N_17071,N_16586,N_16629);
or U17072 (N_17072,N_16987,N_16905);
and U17073 (N_17073,N_16726,N_16514);
nor U17074 (N_17074,N_16562,N_16858);
xnor U17075 (N_17075,N_16755,N_16531);
nand U17076 (N_17076,N_16744,N_16757);
and U17077 (N_17077,N_16688,N_16942);
xor U17078 (N_17078,N_16594,N_16609);
or U17079 (N_17079,N_16918,N_16644);
xnor U17080 (N_17080,N_16650,N_16980);
and U17081 (N_17081,N_16713,N_16973);
or U17082 (N_17082,N_16639,N_16669);
or U17083 (N_17083,N_16745,N_16546);
nor U17084 (N_17084,N_16503,N_16930);
nor U17085 (N_17085,N_16935,N_16734);
or U17086 (N_17086,N_16831,N_16597);
or U17087 (N_17087,N_16585,N_16985);
xnor U17088 (N_17088,N_16857,N_16896);
nor U17089 (N_17089,N_16764,N_16671);
xnor U17090 (N_17090,N_16820,N_16882);
and U17091 (N_17091,N_16795,N_16684);
and U17092 (N_17092,N_16566,N_16596);
or U17093 (N_17093,N_16508,N_16572);
and U17094 (N_17094,N_16667,N_16598);
or U17095 (N_17095,N_16956,N_16678);
or U17096 (N_17096,N_16550,N_16898);
or U17097 (N_17097,N_16780,N_16708);
nand U17098 (N_17098,N_16797,N_16962);
or U17099 (N_17099,N_16588,N_16694);
or U17100 (N_17100,N_16606,N_16920);
xor U17101 (N_17101,N_16735,N_16545);
xnor U17102 (N_17102,N_16666,N_16682);
nand U17103 (N_17103,N_16679,N_16697);
xor U17104 (N_17104,N_16830,N_16775);
nand U17105 (N_17105,N_16819,N_16561);
xor U17106 (N_17106,N_16681,N_16556);
nand U17107 (N_17107,N_16719,N_16967);
nand U17108 (N_17108,N_16974,N_16885);
or U17109 (N_17109,N_16940,N_16994);
nand U17110 (N_17110,N_16615,N_16822);
xor U17111 (N_17111,N_16928,N_16647);
or U17112 (N_17112,N_16730,N_16789);
nand U17113 (N_17113,N_16953,N_16990);
and U17114 (N_17114,N_16641,N_16513);
nand U17115 (N_17115,N_16592,N_16658);
and U17116 (N_17116,N_16722,N_16661);
nand U17117 (N_17117,N_16651,N_16836);
or U17118 (N_17118,N_16603,N_16814);
xor U17119 (N_17119,N_16868,N_16706);
nand U17120 (N_17120,N_16776,N_16555);
xor U17121 (N_17121,N_16619,N_16720);
xor U17122 (N_17122,N_16982,N_16946);
nor U17123 (N_17123,N_16815,N_16564);
or U17124 (N_17124,N_16506,N_16653);
nor U17125 (N_17125,N_16616,N_16848);
and U17126 (N_17126,N_16760,N_16784);
nand U17127 (N_17127,N_16511,N_16817);
and U17128 (N_17128,N_16812,N_16818);
nand U17129 (N_17129,N_16976,N_16664);
and U17130 (N_17130,N_16754,N_16751);
nand U17131 (N_17131,N_16971,N_16892);
or U17132 (N_17132,N_16521,N_16610);
and U17133 (N_17133,N_16923,N_16560);
or U17134 (N_17134,N_16769,N_16986);
nor U17135 (N_17135,N_16816,N_16951);
and U17136 (N_17136,N_16574,N_16889);
or U17137 (N_17137,N_16995,N_16948);
nor U17138 (N_17138,N_16582,N_16821);
xor U17139 (N_17139,N_16645,N_16649);
nand U17140 (N_17140,N_16542,N_16686);
and U17141 (N_17141,N_16652,N_16724);
or U17142 (N_17142,N_16977,N_16532);
or U17143 (N_17143,N_16717,N_16558);
and U17144 (N_17144,N_16931,N_16854);
and U17145 (N_17145,N_16640,N_16939);
nand U17146 (N_17146,N_16975,N_16838);
and U17147 (N_17147,N_16657,N_16676);
xor U17148 (N_17148,N_16993,N_16509);
or U17149 (N_17149,N_16607,N_16736);
nor U17150 (N_17150,N_16519,N_16887);
nand U17151 (N_17151,N_16891,N_16727);
or U17152 (N_17152,N_16504,N_16533);
or U17153 (N_17153,N_16808,N_16673);
nor U17154 (N_17154,N_16909,N_16731);
or U17155 (N_17155,N_16835,N_16979);
xor U17156 (N_17156,N_16583,N_16711);
nand U17157 (N_17157,N_16632,N_16538);
nor U17158 (N_17158,N_16623,N_16823);
or U17159 (N_17159,N_16911,N_16916);
xnor U17160 (N_17160,N_16781,N_16747);
and U17161 (N_17161,N_16861,N_16807);
and U17162 (N_17162,N_16949,N_16624);
nand U17163 (N_17163,N_16978,N_16715);
or U17164 (N_17164,N_16762,N_16759);
xor U17165 (N_17165,N_16829,N_16613);
xor U17166 (N_17166,N_16725,N_16551);
xor U17167 (N_17167,N_16934,N_16709);
nor U17168 (N_17168,N_16548,N_16704);
xnor U17169 (N_17169,N_16771,N_16846);
nand U17170 (N_17170,N_16737,N_16525);
or U17171 (N_17171,N_16984,N_16698);
and U17172 (N_17172,N_16693,N_16802);
and U17173 (N_17173,N_16523,N_16884);
and U17174 (N_17174,N_16913,N_16774);
and U17175 (N_17175,N_16675,N_16879);
and U17176 (N_17176,N_16763,N_16791);
xnor U17177 (N_17177,N_16502,N_16783);
nand U17178 (N_17178,N_16959,N_16768);
nor U17179 (N_17179,N_16799,N_16788);
and U17180 (N_17180,N_16579,N_16528);
or U17181 (N_17181,N_16517,N_16761);
or U17182 (N_17182,N_16906,N_16536);
xor U17183 (N_17183,N_16705,N_16571);
xor U17184 (N_17184,N_16518,N_16860);
or U17185 (N_17185,N_16924,N_16674);
and U17186 (N_17186,N_16537,N_16500);
or U17187 (N_17187,N_16554,N_16894);
or U17188 (N_17188,N_16922,N_16853);
nor U17189 (N_17189,N_16919,N_16680);
xnor U17190 (N_17190,N_16777,N_16999);
nand U17191 (N_17191,N_16947,N_16826);
and U17192 (N_17192,N_16625,N_16577);
nor U17193 (N_17193,N_16798,N_16843);
and U17194 (N_17194,N_16563,N_16565);
xor U17195 (N_17195,N_16850,N_16833);
xnor U17196 (N_17196,N_16878,N_16540);
or U17197 (N_17197,N_16989,N_16867);
or U17198 (N_17198,N_16929,N_16983);
nand U17199 (N_17199,N_16581,N_16654);
xnor U17200 (N_17200,N_16655,N_16877);
nand U17201 (N_17201,N_16943,N_16723);
nand U17202 (N_17202,N_16883,N_16700);
or U17203 (N_17203,N_16512,N_16685);
xor U17204 (N_17204,N_16591,N_16793);
nand U17205 (N_17205,N_16507,N_16714);
and U17206 (N_17206,N_16614,N_16718);
nor U17207 (N_17207,N_16992,N_16968);
xor U17208 (N_17208,N_16608,N_16915);
xnor U17209 (N_17209,N_16593,N_16869);
nand U17210 (N_17210,N_16809,N_16699);
nand U17211 (N_17211,N_16981,N_16958);
xnor U17212 (N_17212,N_16851,N_16997);
nand U17213 (N_17213,N_16801,N_16908);
xor U17214 (N_17214,N_16842,N_16740);
or U17215 (N_17215,N_16729,N_16875);
xor U17216 (N_17216,N_16964,N_16844);
or U17217 (N_17217,N_16874,N_16570);
nand U17218 (N_17218,N_16855,N_16938);
or U17219 (N_17219,N_16903,N_16952);
nand U17220 (N_17220,N_16510,N_16600);
and U17221 (N_17221,N_16941,N_16695);
nand U17222 (N_17222,N_16677,N_16670);
nor U17223 (N_17223,N_16660,N_16834);
xor U17224 (N_17224,N_16683,N_16770);
nand U17225 (N_17225,N_16904,N_16541);
xnor U17226 (N_17226,N_16785,N_16535);
xnor U17227 (N_17227,N_16742,N_16752);
or U17228 (N_17228,N_16758,N_16646);
nor U17229 (N_17229,N_16547,N_16944);
and U17230 (N_17230,N_16847,N_16663);
or U17231 (N_17231,N_16515,N_16527);
nor U17232 (N_17232,N_16865,N_16732);
and U17233 (N_17233,N_16696,N_16620);
nor U17234 (N_17234,N_16501,N_16937);
and U17235 (N_17235,N_16895,N_16824);
and U17236 (N_17236,N_16840,N_16866);
nor U17237 (N_17237,N_16837,N_16804);
and U17238 (N_17238,N_16553,N_16689);
xor U17239 (N_17239,N_16633,N_16966);
nor U17240 (N_17240,N_16863,N_16792);
or U17241 (N_17241,N_16687,N_16886);
nor U17242 (N_17242,N_16602,N_16881);
xor U17243 (N_17243,N_16890,N_16543);
nand U17244 (N_17244,N_16634,N_16611);
xnor U17245 (N_17245,N_16617,N_16778);
xnor U17246 (N_17246,N_16576,N_16955);
and U17247 (N_17247,N_16749,N_16662);
and U17248 (N_17248,N_16957,N_16825);
and U17249 (N_17249,N_16852,N_16796);
nand U17250 (N_17250,N_16648,N_16984);
xnor U17251 (N_17251,N_16872,N_16637);
xor U17252 (N_17252,N_16536,N_16919);
xor U17253 (N_17253,N_16939,N_16693);
xor U17254 (N_17254,N_16912,N_16860);
nor U17255 (N_17255,N_16876,N_16654);
xnor U17256 (N_17256,N_16662,N_16952);
or U17257 (N_17257,N_16570,N_16784);
or U17258 (N_17258,N_16812,N_16711);
or U17259 (N_17259,N_16507,N_16637);
nor U17260 (N_17260,N_16914,N_16769);
nand U17261 (N_17261,N_16762,N_16681);
nand U17262 (N_17262,N_16981,N_16903);
nand U17263 (N_17263,N_16658,N_16704);
and U17264 (N_17264,N_16621,N_16797);
and U17265 (N_17265,N_16754,N_16877);
nand U17266 (N_17266,N_16938,N_16645);
xnor U17267 (N_17267,N_16546,N_16948);
or U17268 (N_17268,N_16503,N_16729);
and U17269 (N_17269,N_16512,N_16873);
or U17270 (N_17270,N_16979,N_16892);
xor U17271 (N_17271,N_16532,N_16531);
or U17272 (N_17272,N_16609,N_16883);
nand U17273 (N_17273,N_16983,N_16700);
and U17274 (N_17274,N_16999,N_16948);
nand U17275 (N_17275,N_16657,N_16839);
or U17276 (N_17276,N_16681,N_16522);
nand U17277 (N_17277,N_16879,N_16537);
nor U17278 (N_17278,N_16888,N_16557);
nor U17279 (N_17279,N_16926,N_16681);
and U17280 (N_17280,N_16837,N_16746);
or U17281 (N_17281,N_16520,N_16565);
and U17282 (N_17282,N_16629,N_16853);
nor U17283 (N_17283,N_16810,N_16749);
or U17284 (N_17284,N_16611,N_16785);
xnor U17285 (N_17285,N_16936,N_16769);
or U17286 (N_17286,N_16648,N_16520);
nor U17287 (N_17287,N_16560,N_16697);
nor U17288 (N_17288,N_16869,N_16850);
nor U17289 (N_17289,N_16750,N_16611);
or U17290 (N_17290,N_16570,N_16709);
nand U17291 (N_17291,N_16531,N_16927);
nand U17292 (N_17292,N_16853,N_16697);
nor U17293 (N_17293,N_16948,N_16778);
xnor U17294 (N_17294,N_16859,N_16910);
nand U17295 (N_17295,N_16500,N_16693);
or U17296 (N_17296,N_16984,N_16764);
or U17297 (N_17297,N_16805,N_16708);
or U17298 (N_17298,N_16851,N_16823);
xor U17299 (N_17299,N_16940,N_16645);
xor U17300 (N_17300,N_16712,N_16992);
xor U17301 (N_17301,N_16901,N_16950);
xor U17302 (N_17302,N_16837,N_16782);
or U17303 (N_17303,N_16867,N_16527);
xor U17304 (N_17304,N_16879,N_16679);
nand U17305 (N_17305,N_16835,N_16941);
nor U17306 (N_17306,N_16912,N_16576);
and U17307 (N_17307,N_16981,N_16768);
nor U17308 (N_17308,N_16984,N_16568);
nor U17309 (N_17309,N_16906,N_16901);
or U17310 (N_17310,N_16916,N_16937);
nor U17311 (N_17311,N_16653,N_16533);
and U17312 (N_17312,N_16588,N_16751);
nand U17313 (N_17313,N_16855,N_16969);
or U17314 (N_17314,N_16972,N_16988);
and U17315 (N_17315,N_16731,N_16527);
nand U17316 (N_17316,N_16592,N_16637);
or U17317 (N_17317,N_16681,N_16713);
nor U17318 (N_17318,N_16750,N_16914);
nor U17319 (N_17319,N_16986,N_16832);
nor U17320 (N_17320,N_16898,N_16798);
or U17321 (N_17321,N_16677,N_16623);
xnor U17322 (N_17322,N_16670,N_16637);
xor U17323 (N_17323,N_16727,N_16964);
nor U17324 (N_17324,N_16805,N_16974);
xnor U17325 (N_17325,N_16779,N_16675);
nor U17326 (N_17326,N_16744,N_16921);
or U17327 (N_17327,N_16765,N_16742);
nor U17328 (N_17328,N_16701,N_16950);
and U17329 (N_17329,N_16753,N_16956);
nand U17330 (N_17330,N_16622,N_16797);
xnor U17331 (N_17331,N_16557,N_16813);
and U17332 (N_17332,N_16850,N_16555);
nand U17333 (N_17333,N_16841,N_16919);
nand U17334 (N_17334,N_16659,N_16896);
xnor U17335 (N_17335,N_16624,N_16662);
or U17336 (N_17336,N_16562,N_16641);
and U17337 (N_17337,N_16689,N_16637);
and U17338 (N_17338,N_16931,N_16751);
nor U17339 (N_17339,N_16840,N_16518);
nand U17340 (N_17340,N_16664,N_16947);
or U17341 (N_17341,N_16627,N_16610);
nor U17342 (N_17342,N_16750,N_16759);
nor U17343 (N_17343,N_16683,N_16955);
or U17344 (N_17344,N_16847,N_16653);
nor U17345 (N_17345,N_16792,N_16512);
nand U17346 (N_17346,N_16752,N_16512);
nand U17347 (N_17347,N_16561,N_16659);
and U17348 (N_17348,N_16987,N_16538);
nand U17349 (N_17349,N_16839,N_16554);
xor U17350 (N_17350,N_16562,N_16966);
and U17351 (N_17351,N_16746,N_16606);
nand U17352 (N_17352,N_16734,N_16962);
nor U17353 (N_17353,N_16777,N_16780);
nor U17354 (N_17354,N_16538,N_16624);
and U17355 (N_17355,N_16749,N_16581);
or U17356 (N_17356,N_16625,N_16823);
and U17357 (N_17357,N_16967,N_16899);
or U17358 (N_17358,N_16600,N_16881);
nor U17359 (N_17359,N_16870,N_16736);
nor U17360 (N_17360,N_16832,N_16969);
and U17361 (N_17361,N_16570,N_16893);
xnor U17362 (N_17362,N_16943,N_16942);
xor U17363 (N_17363,N_16529,N_16785);
and U17364 (N_17364,N_16763,N_16979);
nor U17365 (N_17365,N_16597,N_16915);
xnor U17366 (N_17366,N_16875,N_16989);
xnor U17367 (N_17367,N_16942,N_16770);
nor U17368 (N_17368,N_16634,N_16599);
nand U17369 (N_17369,N_16752,N_16741);
and U17370 (N_17370,N_16759,N_16985);
nand U17371 (N_17371,N_16830,N_16689);
nand U17372 (N_17372,N_16917,N_16829);
and U17373 (N_17373,N_16618,N_16790);
nor U17374 (N_17374,N_16735,N_16710);
xor U17375 (N_17375,N_16628,N_16796);
and U17376 (N_17376,N_16632,N_16536);
xnor U17377 (N_17377,N_16602,N_16526);
nand U17378 (N_17378,N_16902,N_16769);
xnor U17379 (N_17379,N_16633,N_16894);
nand U17380 (N_17380,N_16636,N_16678);
xor U17381 (N_17381,N_16580,N_16815);
nand U17382 (N_17382,N_16805,N_16989);
nand U17383 (N_17383,N_16938,N_16528);
nand U17384 (N_17384,N_16539,N_16689);
or U17385 (N_17385,N_16867,N_16552);
and U17386 (N_17386,N_16621,N_16809);
nand U17387 (N_17387,N_16603,N_16591);
nand U17388 (N_17388,N_16996,N_16649);
nor U17389 (N_17389,N_16508,N_16568);
nor U17390 (N_17390,N_16808,N_16661);
and U17391 (N_17391,N_16728,N_16768);
xor U17392 (N_17392,N_16822,N_16590);
and U17393 (N_17393,N_16893,N_16574);
nand U17394 (N_17394,N_16687,N_16664);
or U17395 (N_17395,N_16830,N_16999);
nand U17396 (N_17396,N_16767,N_16947);
xnor U17397 (N_17397,N_16527,N_16864);
or U17398 (N_17398,N_16855,N_16724);
nand U17399 (N_17399,N_16554,N_16543);
or U17400 (N_17400,N_16722,N_16886);
nand U17401 (N_17401,N_16862,N_16698);
nor U17402 (N_17402,N_16719,N_16553);
xor U17403 (N_17403,N_16597,N_16596);
nor U17404 (N_17404,N_16738,N_16901);
nand U17405 (N_17405,N_16823,N_16958);
and U17406 (N_17406,N_16512,N_16785);
nor U17407 (N_17407,N_16608,N_16857);
and U17408 (N_17408,N_16601,N_16543);
and U17409 (N_17409,N_16672,N_16812);
or U17410 (N_17410,N_16606,N_16600);
xor U17411 (N_17411,N_16928,N_16970);
xor U17412 (N_17412,N_16789,N_16567);
nor U17413 (N_17413,N_16731,N_16640);
nor U17414 (N_17414,N_16843,N_16730);
and U17415 (N_17415,N_16911,N_16584);
nor U17416 (N_17416,N_16692,N_16985);
nor U17417 (N_17417,N_16733,N_16714);
nand U17418 (N_17418,N_16711,N_16601);
nor U17419 (N_17419,N_16726,N_16568);
and U17420 (N_17420,N_16923,N_16972);
nand U17421 (N_17421,N_16720,N_16875);
nand U17422 (N_17422,N_16936,N_16818);
nor U17423 (N_17423,N_16851,N_16938);
or U17424 (N_17424,N_16676,N_16561);
nor U17425 (N_17425,N_16852,N_16776);
and U17426 (N_17426,N_16915,N_16585);
nor U17427 (N_17427,N_16927,N_16587);
xor U17428 (N_17428,N_16998,N_16916);
and U17429 (N_17429,N_16558,N_16822);
nand U17430 (N_17430,N_16949,N_16510);
nor U17431 (N_17431,N_16621,N_16822);
or U17432 (N_17432,N_16881,N_16884);
and U17433 (N_17433,N_16601,N_16598);
and U17434 (N_17434,N_16872,N_16672);
xnor U17435 (N_17435,N_16924,N_16618);
or U17436 (N_17436,N_16907,N_16585);
or U17437 (N_17437,N_16634,N_16754);
nand U17438 (N_17438,N_16942,N_16836);
and U17439 (N_17439,N_16533,N_16683);
nor U17440 (N_17440,N_16859,N_16593);
xnor U17441 (N_17441,N_16802,N_16591);
or U17442 (N_17442,N_16627,N_16825);
nand U17443 (N_17443,N_16831,N_16666);
nand U17444 (N_17444,N_16793,N_16548);
or U17445 (N_17445,N_16539,N_16570);
nor U17446 (N_17446,N_16717,N_16615);
xnor U17447 (N_17447,N_16906,N_16726);
or U17448 (N_17448,N_16829,N_16959);
nor U17449 (N_17449,N_16597,N_16606);
nor U17450 (N_17450,N_16628,N_16704);
nor U17451 (N_17451,N_16990,N_16992);
or U17452 (N_17452,N_16528,N_16692);
and U17453 (N_17453,N_16588,N_16549);
xor U17454 (N_17454,N_16940,N_16595);
nand U17455 (N_17455,N_16949,N_16621);
nand U17456 (N_17456,N_16971,N_16870);
xor U17457 (N_17457,N_16644,N_16755);
nand U17458 (N_17458,N_16708,N_16692);
xor U17459 (N_17459,N_16852,N_16631);
xnor U17460 (N_17460,N_16698,N_16619);
and U17461 (N_17461,N_16690,N_16823);
and U17462 (N_17462,N_16711,N_16929);
or U17463 (N_17463,N_16997,N_16665);
or U17464 (N_17464,N_16888,N_16546);
and U17465 (N_17465,N_16839,N_16802);
nor U17466 (N_17466,N_16780,N_16962);
nor U17467 (N_17467,N_16650,N_16946);
nand U17468 (N_17468,N_16815,N_16694);
and U17469 (N_17469,N_16571,N_16657);
and U17470 (N_17470,N_16640,N_16811);
nor U17471 (N_17471,N_16699,N_16649);
or U17472 (N_17472,N_16749,N_16972);
nor U17473 (N_17473,N_16596,N_16706);
and U17474 (N_17474,N_16732,N_16503);
nand U17475 (N_17475,N_16646,N_16721);
nand U17476 (N_17476,N_16965,N_16740);
xnor U17477 (N_17477,N_16730,N_16578);
or U17478 (N_17478,N_16589,N_16604);
xnor U17479 (N_17479,N_16555,N_16751);
and U17480 (N_17480,N_16518,N_16937);
and U17481 (N_17481,N_16842,N_16899);
nand U17482 (N_17482,N_16953,N_16902);
and U17483 (N_17483,N_16632,N_16503);
nor U17484 (N_17484,N_16705,N_16534);
xor U17485 (N_17485,N_16566,N_16934);
nor U17486 (N_17486,N_16524,N_16809);
and U17487 (N_17487,N_16922,N_16560);
nor U17488 (N_17488,N_16693,N_16743);
and U17489 (N_17489,N_16847,N_16934);
nor U17490 (N_17490,N_16998,N_16844);
nor U17491 (N_17491,N_16818,N_16530);
and U17492 (N_17492,N_16831,N_16796);
nand U17493 (N_17493,N_16663,N_16732);
and U17494 (N_17494,N_16931,N_16802);
nor U17495 (N_17495,N_16906,N_16888);
nand U17496 (N_17496,N_16947,N_16835);
nor U17497 (N_17497,N_16737,N_16704);
or U17498 (N_17498,N_16691,N_16622);
xnor U17499 (N_17499,N_16718,N_16987);
or U17500 (N_17500,N_17475,N_17497);
and U17501 (N_17501,N_17439,N_17239);
nor U17502 (N_17502,N_17402,N_17216);
and U17503 (N_17503,N_17010,N_17045);
nand U17504 (N_17504,N_17449,N_17370);
nor U17505 (N_17505,N_17009,N_17396);
or U17506 (N_17506,N_17426,N_17037);
and U17507 (N_17507,N_17338,N_17485);
or U17508 (N_17508,N_17266,N_17321);
nor U17509 (N_17509,N_17435,N_17339);
nor U17510 (N_17510,N_17210,N_17020);
xnor U17511 (N_17511,N_17131,N_17021);
and U17512 (N_17512,N_17223,N_17265);
nand U17513 (N_17513,N_17227,N_17109);
nand U17514 (N_17514,N_17005,N_17200);
or U17515 (N_17515,N_17376,N_17208);
xnor U17516 (N_17516,N_17305,N_17440);
and U17517 (N_17517,N_17060,N_17425);
xnor U17518 (N_17518,N_17309,N_17405);
nand U17519 (N_17519,N_17457,N_17167);
and U17520 (N_17520,N_17031,N_17065);
nor U17521 (N_17521,N_17384,N_17052);
nand U17522 (N_17522,N_17261,N_17282);
or U17523 (N_17523,N_17471,N_17203);
or U17524 (N_17524,N_17178,N_17313);
xor U17525 (N_17525,N_17142,N_17491);
nor U17526 (N_17526,N_17311,N_17241);
and U17527 (N_17527,N_17111,N_17036);
nor U17528 (N_17528,N_17272,N_17455);
or U17529 (N_17529,N_17296,N_17377);
or U17530 (N_17530,N_17168,N_17018);
nor U17531 (N_17531,N_17153,N_17026);
xor U17532 (N_17532,N_17038,N_17127);
nor U17533 (N_17533,N_17089,N_17304);
nand U17534 (N_17534,N_17161,N_17092);
xnor U17535 (N_17535,N_17137,N_17195);
and U17536 (N_17536,N_17225,N_17229);
nand U17537 (N_17537,N_17199,N_17141);
xor U17538 (N_17538,N_17248,N_17289);
nand U17539 (N_17539,N_17076,N_17262);
nor U17540 (N_17540,N_17243,N_17140);
nand U17541 (N_17541,N_17003,N_17416);
nor U17542 (N_17542,N_17270,N_17401);
nor U17543 (N_17543,N_17107,N_17443);
or U17544 (N_17544,N_17252,N_17119);
nand U17545 (N_17545,N_17333,N_17336);
nor U17546 (N_17546,N_17205,N_17108);
and U17547 (N_17547,N_17410,N_17447);
xor U17548 (N_17548,N_17367,N_17334);
or U17549 (N_17549,N_17156,N_17007);
nand U17550 (N_17550,N_17024,N_17068);
xor U17551 (N_17551,N_17433,N_17351);
xnor U17552 (N_17552,N_17383,N_17035);
and U17553 (N_17553,N_17171,N_17206);
nand U17554 (N_17554,N_17352,N_17335);
or U17555 (N_17555,N_17030,N_17423);
nand U17556 (N_17556,N_17049,N_17464);
or U17557 (N_17557,N_17274,N_17209);
or U17558 (N_17558,N_17436,N_17326);
and U17559 (N_17559,N_17247,N_17152);
nor U17560 (N_17560,N_17215,N_17213);
and U17561 (N_17561,N_17102,N_17197);
xnor U17562 (N_17562,N_17479,N_17498);
nand U17563 (N_17563,N_17177,N_17059);
nand U17564 (N_17564,N_17421,N_17337);
or U17565 (N_17565,N_17079,N_17063);
nor U17566 (N_17566,N_17044,N_17245);
nand U17567 (N_17567,N_17353,N_17364);
xor U17568 (N_17568,N_17162,N_17157);
nor U17569 (N_17569,N_17409,N_17269);
xor U17570 (N_17570,N_17072,N_17032);
nor U17571 (N_17571,N_17285,N_17190);
or U17572 (N_17572,N_17347,N_17175);
xnor U17573 (N_17573,N_17123,N_17230);
xor U17574 (N_17574,N_17244,N_17417);
nand U17575 (N_17575,N_17254,N_17332);
nor U17576 (N_17576,N_17414,N_17323);
nor U17577 (N_17577,N_17104,N_17488);
nor U17578 (N_17578,N_17438,N_17188);
nor U17579 (N_17579,N_17138,N_17412);
xnor U17580 (N_17580,N_17105,N_17481);
xnor U17581 (N_17581,N_17187,N_17070);
nor U17582 (N_17582,N_17120,N_17317);
and U17583 (N_17583,N_17166,N_17028);
nor U17584 (N_17584,N_17389,N_17374);
nand U17585 (N_17585,N_17379,N_17150);
and U17586 (N_17586,N_17180,N_17048);
and U17587 (N_17587,N_17484,N_17135);
nand U17588 (N_17588,N_17429,N_17487);
xnor U17589 (N_17589,N_17495,N_17240);
or U17590 (N_17590,N_17098,N_17226);
nor U17591 (N_17591,N_17399,N_17341);
and U17592 (N_17592,N_17477,N_17053);
nand U17593 (N_17593,N_17090,N_17378);
or U17594 (N_17594,N_17329,N_17393);
or U17595 (N_17595,N_17027,N_17486);
nand U17596 (N_17596,N_17354,N_17281);
and U17597 (N_17597,N_17386,N_17173);
and U17598 (N_17598,N_17460,N_17290);
xnor U17599 (N_17599,N_17307,N_17058);
xnor U17600 (N_17600,N_17413,N_17375);
xnor U17601 (N_17601,N_17418,N_17381);
nor U17602 (N_17602,N_17343,N_17218);
xor U17603 (N_17603,N_17144,N_17012);
nand U17604 (N_17604,N_17004,N_17118);
or U17605 (N_17605,N_17441,N_17047);
nor U17606 (N_17606,N_17453,N_17350);
nor U17607 (N_17607,N_17330,N_17204);
nor U17608 (N_17608,N_17328,N_17291);
or U17609 (N_17609,N_17061,N_17366);
nor U17610 (N_17610,N_17451,N_17346);
nor U17611 (N_17611,N_17388,N_17077);
and U17612 (N_17612,N_17404,N_17469);
nand U17613 (N_17613,N_17255,N_17126);
xor U17614 (N_17614,N_17181,N_17277);
nor U17615 (N_17615,N_17392,N_17081);
nand U17616 (N_17616,N_17106,N_17428);
nand U17617 (N_17617,N_17033,N_17349);
nand U17618 (N_17618,N_17198,N_17094);
or U17619 (N_17619,N_17182,N_17437);
or U17620 (N_17620,N_17236,N_17160);
xor U17621 (N_17621,N_17422,N_17019);
xor U17622 (N_17622,N_17459,N_17006);
xnor U17623 (N_17623,N_17041,N_17001);
nand U17624 (N_17624,N_17040,N_17263);
and U17625 (N_17625,N_17008,N_17297);
or U17626 (N_17626,N_17348,N_17125);
nor U17627 (N_17627,N_17163,N_17043);
nor U17628 (N_17628,N_17278,N_17325);
or U17629 (N_17629,N_17113,N_17258);
xor U17630 (N_17630,N_17000,N_17080);
xor U17631 (N_17631,N_17073,N_17315);
nand U17632 (N_17632,N_17302,N_17222);
nand U17633 (N_17633,N_17452,N_17232);
nor U17634 (N_17634,N_17042,N_17463);
nor U17635 (N_17635,N_17124,N_17286);
xnor U17636 (N_17636,N_17221,N_17115);
and U17637 (N_17637,N_17264,N_17308);
xnor U17638 (N_17638,N_17234,N_17238);
nand U17639 (N_17639,N_17318,N_17380);
nor U17640 (N_17640,N_17039,N_17114);
nand U17641 (N_17641,N_17331,N_17155);
nand U17642 (N_17642,N_17319,N_17298);
xor U17643 (N_17643,N_17088,N_17112);
and U17644 (N_17644,N_17470,N_17116);
xnor U17645 (N_17645,N_17496,N_17276);
and U17646 (N_17646,N_17397,N_17476);
and U17647 (N_17647,N_17093,N_17344);
xor U17648 (N_17648,N_17097,N_17251);
nor U17649 (N_17649,N_17085,N_17034);
nor U17650 (N_17650,N_17253,N_17283);
nor U17651 (N_17651,N_17300,N_17246);
or U17652 (N_17652,N_17029,N_17450);
nand U17653 (N_17653,N_17342,N_17117);
and U17654 (N_17654,N_17489,N_17267);
nor U17655 (N_17655,N_17231,N_17235);
or U17656 (N_17656,N_17151,N_17084);
nand U17657 (N_17657,N_17363,N_17202);
nand U17658 (N_17658,N_17014,N_17301);
xnor U17659 (N_17659,N_17165,N_17442);
and U17660 (N_17660,N_17327,N_17303);
nand U17661 (N_17661,N_17445,N_17492);
xnor U17662 (N_17662,N_17419,N_17154);
xor U17663 (N_17663,N_17023,N_17299);
nor U17664 (N_17664,N_17273,N_17083);
nor U17665 (N_17665,N_17170,N_17193);
nor U17666 (N_17666,N_17082,N_17212);
or U17667 (N_17667,N_17186,N_17087);
nor U17668 (N_17668,N_17294,N_17067);
nor U17669 (N_17669,N_17217,N_17207);
or U17670 (N_17670,N_17444,N_17016);
xor U17671 (N_17671,N_17340,N_17145);
and U17672 (N_17672,N_17288,N_17249);
nand U17673 (N_17673,N_17385,N_17196);
and U17674 (N_17674,N_17483,N_17136);
nand U17675 (N_17675,N_17172,N_17293);
nor U17676 (N_17676,N_17257,N_17357);
nor U17677 (N_17677,N_17233,N_17179);
xnor U17678 (N_17678,N_17075,N_17101);
nand U17679 (N_17679,N_17482,N_17250);
or U17680 (N_17680,N_17415,N_17129);
xnor U17681 (N_17681,N_17295,N_17345);
or U17682 (N_17682,N_17499,N_17134);
nor U17683 (N_17683,N_17406,N_17174);
nor U17684 (N_17684,N_17260,N_17054);
and U17685 (N_17685,N_17066,N_17096);
xor U17686 (N_17686,N_17395,N_17362);
xor U17687 (N_17687,N_17280,N_17176);
nand U17688 (N_17688,N_17224,N_17394);
and U17689 (N_17689,N_17462,N_17259);
or U17690 (N_17690,N_17391,N_17320);
nor U17691 (N_17691,N_17078,N_17184);
nand U17692 (N_17692,N_17312,N_17086);
and U17693 (N_17693,N_17474,N_17403);
xor U17694 (N_17694,N_17424,N_17368);
nor U17695 (N_17695,N_17159,N_17103);
nor U17696 (N_17696,N_17011,N_17057);
and U17697 (N_17697,N_17373,N_17387);
xor U17698 (N_17698,N_17022,N_17110);
nor U17699 (N_17699,N_17133,N_17466);
nand U17700 (N_17700,N_17369,N_17015);
and U17701 (N_17701,N_17356,N_17478);
xnor U17702 (N_17702,N_17493,N_17411);
xnor U17703 (N_17703,N_17316,N_17132);
or U17704 (N_17704,N_17467,N_17494);
nor U17705 (N_17705,N_17310,N_17201);
or U17706 (N_17706,N_17279,N_17446);
nand U17707 (N_17707,N_17458,N_17192);
and U17708 (N_17708,N_17139,N_17191);
nand U17709 (N_17709,N_17324,N_17149);
nor U17710 (N_17710,N_17062,N_17372);
and U17711 (N_17711,N_17284,N_17268);
and U17712 (N_17712,N_17013,N_17434);
nor U17713 (N_17713,N_17448,N_17194);
or U17714 (N_17714,N_17322,N_17220);
xor U17715 (N_17715,N_17055,N_17400);
and U17716 (N_17716,N_17128,N_17473);
xnor U17717 (N_17717,N_17358,N_17256);
and U17718 (N_17718,N_17100,N_17025);
xnor U17719 (N_17719,N_17390,N_17214);
or U17720 (N_17720,N_17355,N_17095);
nor U17721 (N_17721,N_17069,N_17122);
or U17722 (N_17722,N_17360,N_17465);
nand U17723 (N_17723,N_17398,N_17228);
and U17724 (N_17724,N_17468,N_17430);
and U17725 (N_17725,N_17183,N_17472);
xor U17726 (N_17726,N_17432,N_17091);
nor U17727 (N_17727,N_17454,N_17017);
xor U17728 (N_17728,N_17121,N_17051);
nand U17729 (N_17729,N_17292,N_17046);
and U17730 (N_17730,N_17287,N_17056);
xor U17731 (N_17731,N_17158,N_17148);
xnor U17732 (N_17732,N_17382,N_17143);
nand U17733 (N_17733,N_17456,N_17219);
xnor U17734 (N_17734,N_17147,N_17461);
xnor U17735 (N_17735,N_17237,N_17242);
or U17736 (N_17736,N_17146,N_17271);
or U17737 (N_17737,N_17490,N_17002);
or U17738 (N_17738,N_17371,N_17314);
nand U17739 (N_17739,N_17169,N_17050);
nor U17740 (N_17740,N_17185,N_17306);
and U17741 (N_17741,N_17071,N_17427);
or U17742 (N_17742,N_17407,N_17211);
nor U17743 (N_17743,N_17408,N_17480);
nand U17744 (N_17744,N_17099,N_17164);
xor U17745 (N_17745,N_17189,N_17275);
xnor U17746 (N_17746,N_17431,N_17130);
nor U17747 (N_17747,N_17359,N_17361);
nor U17748 (N_17748,N_17074,N_17064);
or U17749 (N_17749,N_17420,N_17365);
and U17750 (N_17750,N_17303,N_17126);
nand U17751 (N_17751,N_17480,N_17137);
and U17752 (N_17752,N_17345,N_17037);
nor U17753 (N_17753,N_17399,N_17266);
and U17754 (N_17754,N_17212,N_17435);
xor U17755 (N_17755,N_17387,N_17461);
nor U17756 (N_17756,N_17355,N_17394);
xor U17757 (N_17757,N_17144,N_17467);
or U17758 (N_17758,N_17088,N_17174);
and U17759 (N_17759,N_17187,N_17113);
xor U17760 (N_17760,N_17464,N_17409);
xnor U17761 (N_17761,N_17412,N_17475);
nor U17762 (N_17762,N_17076,N_17078);
or U17763 (N_17763,N_17348,N_17160);
nand U17764 (N_17764,N_17351,N_17153);
xor U17765 (N_17765,N_17423,N_17495);
or U17766 (N_17766,N_17486,N_17399);
nand U17767 (N_17767,N_17142,N_17045);
and U17768 (N_17768,N_17135,N_17329);
xnor U17769 (N_17769,N_17009,N_17470);
and U17770 (N_17770,N_17497,N_17165);
and U17771 (N_17771,N_17368,N_17404);
nor U17772 (N_17772,N_17246,N_17449);
or U17773 (N_17773,N_17303,N_17395);
nand U17774 (N_17774,N_17248,N_17417);
nand U17775 (N_17775,N_17274,N_17486);
nor U17776 (N_17776,N_17032,N_17297);
nand U17777 (N_17777,N_17418,N_17280);
and U17778 (N_17778,N_17375,N_17419);
or U17779 (N_17779,N_17268,N_17425);
nor U17780 (N_17780,N_17203,N_17450);
nand U17781 (N_17781,N_17176,N_17348);
xnor U17782 (N_17782,N_17063,N_17372);
nor U17783 (N_17783,N_17147,N_17226);
xor U17784 (N_17784,N_17215,N_17240);
and U17785 (N_17785,N_17373,N_17087);
or U17786 (N_17786,N_17430,N_17319);
nand U17787 (N_17787,N_17238,N_17295);
nand U17788 (N_17788,N_17143,N_17116);
xnor U17789 (N_17789,N_17105,N_17426);
nand U17790 (N_17790,N_17196,N_17203);
or U17791 (N_17791,N_17147,N_17441);
nand U17792 (N_17792,N_17324,N_17265);
nand U17793 (N_17793,N_17233,N_17365);
nor U17794 (N_17794,N_17131,N_17203);
nor U17795 (N_17795,N_17040,N_17167);
nand U17796 (N_17796,N_17138,N_17128);
xnor U17797 (N_17797,N_17482,N_17189);
and U17798 (N_17798,N_17491,N_17162);
nand U17799 (N_17799,N_17398,N_17058);
nand U17800 (N_17800,N_17222,N_17216);
xnor U17801 (N_17801,N_17079,N_17173);
or U17802 (N_17802,N_17208,N_17085);
or U17803 (N_17803,N_17295,N_17368);
and U17804 (N_17804,N_17019,N_17221);
nor U17805 (N_17805,N_17190,N_17386);
and U17806 (N_17806,N_17465,N_17363);
nand U17807 (N_17807,N_17169,N_17486);
xnor U17808 (N_17808,N_17191,N_17307);
nor U17809 (N_17809,N_17033,N_17237);
xor U17810 (N_17810,N_17162,N_17398);
and U17811 (N_17811,N_17110,N_17075);
and U17812 (N_17812,N_17381,N_17453);
or U17813 (N_17813,N_17474,N_17464);
and U17814 (N_17814,N_17349,N_17406);
nor U17815 (N_17815,N_17142,N_17087);
and U17816 (N_17816,N_17011,N_17311);
and U17817 (N_17817,N_17244,N_17423);
or U17818 (N_17818,N_17471,N_17357);
nand U17819 (N_17819,N_17479,N_17246);
or U17820 (N_17820,N_17274,N_17419);
xor U17821 (N_17821,N_17126,N_17033);
nand U17822 (N_17822,N_17064,N_17411);
nand U17823 (N_17823,N_17085,N_17293);
and U17824 (N_17824,N_17187,N_17221);
nor U17825 (N_17825,N_17485,N_17491);
and U17826 (N_17826,N_17417,N_17254);
or U17827 (N_17827,N_17253,N_17274);
nand U17828 (N_17828,N_17494,N_17391);
xnor U17829 (N_17829,N_17230,N_17092);
nor U17830 (N_17830,N_17399,N_17462);
xor U17831 (N_17831,N_17083,N_17250);
and U17832 (N_17832,N_17445,N_17405);
xor U17833 (N_17833,N_17115,N_17196);
nor U17834 (N_17834,N_17089,N_17418);
or U17835 (N_17835,N_17461,N_17261);
xnor U17836 (N_17836,N_17084,N_17087);
xor U17837 (N_17837,N_17338,N_17478);
and U17838 (N_17838,N_17115,N_17348);
nor U17839 (N_17839,N_17288,N_17427);
or U17840 (N_17840,N_17372,N_17052);
and U17841 (N_17841,N_17183,N_17253);
and U17842 (N_17842,N_17249,N_17159);
or U17843 (N_17843,N_17482,N_17079);
nor U17844 (N_17844,N_17340,N_17497);
xnor U17845 (N_17845,N_17280,N_17133);
xnor U17846 (N_17846,N_17017,N_17260);
nor U17847 (N_17847,N_17307,N_17079);
or U17848 (N_17848,N_17059,N_17016);
or U17849 (N_17849,N_17435,N_17424);
xnor U17850 (N_17850,N_17203,N_17301);
xor U17851 (N_17851,N_17096,N_17130);
nand U17852 (N_17852,N_17424,N_17366);
xor U17853 (N_17853,N_17281,N_17259);
nor U17854 (N_17854,N_17152,N_17158);
nor U17855 (N_17855,N_17353,N_17262);
xnor U17856 (N_17856,N_17366,N_17305);
or U17857 (N_17857,N_17410,N_17486);
xor U17858 (N_17858,N_17168,N_17073);
and U17859 (N_17859,N_17009,N_17109);
nor U17860 (N_17860,N_17316,N_17400);
nor U17861 (N_17861,N_17225,N_17231);
nor U17862 (N_17862,N_17191,N_17451);
and U17863 (N_17863,N_17052,N_17483);
and U17864 (N_17864,N_17116,N_17280);
xor U17865 (N_17865,N_17171,N_17303);
and U17866 (N_17866,N_17043,N_17167);
nand U17867 (N_17867,N_17415,N_17012);
or U17868 (N_17868,N_17244,N_17095);
nand U17869 (N_17869,N_17478,N_17462);
or U17870 (N_17870,N_17033,N_17013);
xnor U17871 (N_17871,N_17369,N_17054);
or U17872 (N_17872,N_17113,N_17017);
and U17873 (N_17873,N_17059,N_17393);
nor U17874 (N_17874,N_17216,N_17491);
nor U17875 (N_17875,N_17024,N_17116);
xnor U17876 (N_17876,N_17494,N_17121);
xor U17877 (N_17877,N_17414,N_17438);
and U17878 (N_17878,N_17001,N_17446);
nor U17879 (N_17879,N_17290,N_17170);
xor U17880 (N_17880,N_17248,N_17264);
and U17881 (N_17881,N_17224,N_17111);
xnor U17882 (N_17882,N_17487,N_17393);
and U17883 (N_17883,N_17496,N_17024);
or U17884 (N_17884,N_17238,N_17301);
xor U17885 (N_17885,N_17418,N_17296);
xor U17886 (N_17886,N_17195,N_17404);
nand U17887 (N_17887,N_17342,N_17280);
nand U17888 (N_17888,N_17197,N_17172);
nand U17889 (N_17889,N_17174,N_17267);
or U17890 (N_17890,N_17298,N_17106);
nor U17891 (N_17891,N_17321,N_17273);
and U17892 (N_17892,N_17357,N_17490);
and U17893 (N_17893,N_17384,N_17342);
nor U17894 (N_17894,N_17186,N_17072);
and U17895 (N_17895,N_17194,N_17004);
nor U17896 (N_17896,N_17313,N_17328);
xnor U17897 (N_17897,N_17253,N_17298);
or U17898 (N_17898,N_17474,N_17273);
or U17899 (N_17899,N_17139,N_17028);
xor U17900 (N_17900,N_17124,N_17233);
nor U17901 (N_17901,N_17148,N_17332);
xnor U17902 (N_17902,N_17092,N_17052);
nor U17903 (N_17903,N_17414,N_17024);
xnor U17904 (N_17904,N_17013,N_17157);
nand U17905 (N_17905,N_17360,N_17298);
nand U17906 (N_17906,N_17491,N_17279);
nor U17907 (N_17907,N_17138,N_17041);
nor U17908 (N_17908,N_17498,N_17284);
xnor U17909 (N_17909,N_17269,N_17368);
xor U17910 (N_17910,N_17124,N_17062);
and U17911 (N_17911,N_17201,N_17176);
or U17912 (N_17912,N_17470,N_17128);
xnor U17913 (N_17913,N_17147,N_17196);
xnor U17914 (N_17914,N_17024,N_17325);
nor U17915 (N_17915,N_17346,N_17010);
and U17916 (N_17916,N_17170,N_17350);
or U17917 (N_17917,N_17216,N_17125);
nand U17918 (N_17918,N_17393,N_17018);
nor U17919 (N_17919,N_17154,N_17257);
xor U17920 (N_17920,N_17315,N_17358);
or U17921 (N_17921,N_17038,N_17124);
nand U17922 (N_17922,N_17455,N_17004);
or U17923 (N_17923,N_17374,N_17324);
and U17924 (N_17924,N_17048,N_17060);
xor U17925 (N_17925,N_17215,N_17203);
nor U17926 (N_17926,N_17462,N_17448);
or U17927 (N_17927,N_17029,N_17315);
xor U17928 (N_17928,N_17260,N_17460);
xnor U17929 (N_17929,N_17207,N_17456);
xor U17930 (N_17930,N_17297,N_17349);
and U17931 (N_17931,N_17016,N_17152);
and U17932 (N_17932,N_17074,N_17058);
nor U17933 (N_17933,N_17013,N_17488);
and U17934 (N_17934,N_17350,N_17058);
and U17935 (N_17935,N_17159,N_17056);
nand U17936 (N_17936,N_17058,N_17123);
nand U17937 (N_17937,N_17111,N_17062);
or U17938 (N_17938,N_17284,N_17319);
xnor U17939 (N_17939,N_17378,N_17390);
xor U17940 (N_17940,N_17437,N_17322);
or U17941 (N_17941,N_17388,N_17015);
nor U17942 (N_17942,N_17254,N_17028);
nand U17943 (N_17943,N_17245,N_17433);
or U17944 (N_17944,N_17407,N_17372);
nor U17945 (N_17945,N_17176,N_17496);
xnor U17946 (N_17946,N_17296,N_17156);
nor U17947 (N_17947,N_17103,N_17131);
nor U17948 (N_17948,N_17077,N_17119);
or U17949 (N_17949,N_17337,N_17248);
nand U17950 (N_17950,N_17376,N_17238);
nor U17951 (N_17951,N_17206,N_17415);
or U17952 (N_17952,N_17326,N_17259);
nand U17953 (N_17953,N_17399,N_17209);
and U17954 (N_17954,N_17034,N_17366);
nor U17955 (N_17955,N_17062,N_17465);
nor U17956 (N_17956,N_17389,N_17475);
nand U17957 (N_17957,N_17431,N_17232);
xor U17958 (N_17958,N_17228,N_17423);
xnor U17959 (N_17959,N_17363,N_17194);
xnor U17960 (N_17960,N_17420,N_17252);
nand U17961 (N_17961,N_17001,N_17368);
or U17962 (N_17962,N_17204,N_17357);
nor U17963 (N_17963,N_17179,N_17186);
and U17964 (N_17964,N_17490,N_17342);
and U17965 (N_17965,N_17152,N_17217);
or U17966 (N_17966,N_17196,N_17306);
xor U17967 (N_17967,N_17407,N_17236);
nand U17968 (N_17968,N_17249,N_17219);
nand U17969 (N_17969,N_17016,N_17012);
and U17970 (N_17970,N_17135,N_17153);
or U17971 (N_17971,N_17300,N_17035);
nand U17972 (N_17972,N_17363,N_17395);
nand U17973 (N_17973,N_17278,N_17013);
nand U17974 (N_17974,N_17369,N_17253);
nand U17975 (N_17975,N_17176,N_17305);
nor U17976 (N_17976,N_17451,N_17153);
nor U17977 (N_17977,N_17331,N_17409);
xor U17978 (N_17978,N_17401,N_17400);
nand U17979 (N_17979,N_17120,N_17310);
nand U17980 (N_17980,N_17427,N_17078);
nor U17981 (N_17981,N_17084,N_17052);
nor U17982 (N_17982,N_17167,N_17085);
xnor U17983 (N_17983,N_17477,N_17175);
and U17984 (N_17984,N_17194,N_17324);
nand U17985 (N_17985,N_17016,N_17335);
or U17986 (N_17986,N_17493,N_17211);
xnor U17987 (N_17987,N_17252,N_17049);
nor U17988 (N_17988,N_17026,N_17190);
xnor U17989 (N_17989,N_17394,N_17323);
xnor U17990 (N_17990,N_17230,N_17026);
nand U17991 (N_17991,N_17187,N_17401);
xnor U17992 (N_17992,N_17212,N_17402);
and U17993 (N_17993,N_17426,N_17235);
and U17994 (N_17994,N_17187,N_17045);
nor U17995 (N_17995,N_17002,N_17111);
nand U17996 (N_17996,N_17195,N_17139);
nand U17997 (N_17997,N_17196,N_17042);
and U17998 (N_17998,N_17262,N_17217);
xor U17999 (N_17999,N_17039,N_17004);
nand U18000 (N_18000,N_17609,N_17598);
nor U18001 (N_18001,N_17631,N_17887);
nor U18002 (N_18002,N_17641,N_17828);
nand U18003 (N_18003,N_17614,N_17522);
nor U18004 (N_18004,N_17584,N_17506);
and U18005 (N_18005,N_17503,N_17940);
nor U18006 (N_18006,N_17585,N_17814);
nor U18007 (N_18007,N_17694,N_17508);
xnor U18008 (N_18008,N_17956,N_17693);
xor U18009 (N_18009,N_17580,N_17864);
nand U18010 (N_18010,N_17821,N_17516);
or U18011 (N_18011,N_17966,N_17946);
and U18012 (N_18012,N_17568,N_17911);
xnor U18013 (N_18013,N_17791,N_17768);
nand U18014 (N_18014,N_17850,N_17872);
xor U18015 (N_18015,N_17504,N_17812);
nor U18016 (N_18016,N_17686,N_17615);
or U18017 (N_18017,N_17889,N_17852);
or U18018 (N_18018,N_17886,N_17752);
or U18019 (N_18019,N_17639,N_17514);
and U18020 (N_18020,N_17663,N_17566);
nor U18021 (N_18021,N_17803,N_17815);
xor U18022 (N_18022,N_17804,N_17955);
and U18023 (N_18023,N_17715,N_17826);
and U18024 (N_18024,N_17511,N_17685);
and U18025 (N_18025,N_17684,N_17860);
and U18026 (N_18026,N_17729,N_17848);
xor U18027 (N_18027,N_17755,N_17648);
or U18028 (N_18028,N_17865,N_17710);
nor U18029 (N_18029,N_17595,N_17957);
xnor U18030 (N_18030,N_17664,N_17737);
and U18031 (N_18031,N_17870,N_17934);
nor U18032 (N_18032,N_17780,N_17976);
xnor U18033 (N_18033,N_17843,N_17625);
and U18034 (N_18034,N_17820,N_17844);
nor U18035 (N_18035,N_17905,N_17990);
or U18036 (N_18036,N_17787,N_17696);
xor U18037 (N_18037,N_17569,N_17670);
or U18038 (N_18038,N_17851,N_17888);
or U18039 (N_18039,N_17903,N_17611);
nand U18040 (N_18040,N_17853,N_17979);
nand U18041 (N_18041,N_17950,N_17662);
and U18042 (N_18042,N_17770,N_17939);
nand U18043 (N_18043,N_17588,N_17512);
xor U18044 (N_18044,N_17739,N_17970);
or U18045 (N_18045,N_17721,N_17777);
or U18046 (N_18046,N_17863,N_17666);
nand U18047 (N_18047,N_17628,N_17859);
or U18048 (N_18048,N_17608,N_17700);
and U18049 (N_18049,N_17834,N_17753);
xnor U18050 (N_18050,N_17786,N_17640);
xor U18051 (N_18051,N_17682,N_17873);
and U18052 (N_18052,N_17871,N_17731);
or U18053 (N_18053,N_17788,N_17652);
nand U18054 (N_18054,N_17881,N_17965);
or U18055 (N_18055,N_17936,N_17758);
xor U18056 (N_18056,N_17540,N_17901);
nand U18057 (N_18057,N_17691,N_17894);
nor U18058 (N_18058,N_17885,N_17722);
xor U18059 (N_18059,N_17784,N_17633);
nand U18060 (N_18060,N_17725,N_17751);
nor U18061 (N_18061,N_17763,N_17654);
nand U18062 (N_18062,N_17741,N_17717);
or U18063 (N_18063,N_17525,N_17973);
or U18064 (N_18064,N_17938,N_17866);
xor U18065 (N_18065,N_17782,N_17712);
nand U18066 (N_18066,N_17714,N_17656);
or U18067 (N_18067,N_17541,N_17773);
and U18068 (N_18068,N_17879,N_17621);
or U18069 (N_18069,N_17984,N_17981);
xnor U18070 (N_18070,N_17718,N_17573);
nor U18071 (N_18071,N_17762,N_17749);
xnor U18072 (N_18072,N_17944,N_17507);
nor U18073 (N_18073,N_17623,N_17515);
and U18074 (N_18074,N_17775,N_17672);
and U18075 (N_18075,N_17612,N_17627);
and U18076 (N_18076,N_17618,N_17993);
or U18077 (N_18077,N_17530,N_17500);
nand U18078 (N_18078,N_17501,N_17519);
or U18079 (N_18079,N_17747,N_17667);
and U18080 (N_18080,N_17575,N_17605);
nor U18081 (N_18081,N_17964,N_17730);
nor U18082 (N_18082,N_17931,N_17977);
and U18083 (N_18083,N_17690,N_17744);
xor U18084 (N_18084,N_17898,N_17838);
or U18085 (N_18085,N_17526,N_17858);
xnor U18086 (N_18086,N_17698,N_17831);
and U18087 (N_18087,N_17902,N_17527);
or U18088 (N_18088,N_17620,N_17520);
or U18089 (N_18089,N_17555,N_17942);
nand U18090 (N_18090,N_17660,N_17937);
nand U18091 (N_18091,N_17671,N_17510);
nand U18092 (N_18092,N_17845,N_17706);
nor U18093 (N_18093,N_17783,N_17759);
or U18094 (N_18094,N_17592,N_17819);
xor U18095 (N_18095,N_17825,N_17891);
nor U18096 (N_18096,N_17792,N_17842);
nor U18097 (N_18097,N_17771,N_17896);
nor U18098 (N_18098,N_17743,N_17805);
or U18099 (N_18099,N_17920,N_17883);
and U18100 (N_18100,N_17547,N_17810);
xor U18101 (N_18101,N_17807,N_17968);
nand U18102 (N_18102,N_17897,N_17932);
xor U18103 (N_18103,N_17914,N_17745);
nor U18104 (N_18104,N_17818,N_17912);
and U18105 (N_18105,N_17997,N_17794);
and U18106 (N_18106,N_17553,N_17742);
and U18107 (N_18107,N_17567,N_17680);
nor U18108 (N_18108,N_17960,N_17558);
nand U18109 (N_18109,N_17638,N_17796);
xor U18110 (N_18110,N_17972,N_17740);
xor U18111 (N_18111,N_17548,N_17816);
nand U18112 (N_18112,N_17980,N_17996);
xnor U18113 (N_18113,N_17849,N_17907);
nor U18114 (N_18114,N_17673,N_17554);
xnor U18115 (N_18115,N_17665,N_17550);
or U18116 (N_18116,N_17579,N_17534);
nand U18117 (N_18117,N_17529,N_17653);
nand U18118 (N_18118,N_17702,N_17687);
nand U18119 (N_18119,N_17813,N_17716);
nand U18120 (N_18120,N_17929,N_17969);
or U18121 (N_18121,N_17925,N_17982);
and U18122 (N_18122,N_17890,N_17589);
and U18123 (N_18123,N_17926,N_17798);
nor U18124 (N_18124,N_17531,N_17622);
nand U18125 (N_18125,N_17836,N_17817);
nand U18126 (N_18126,N_17617,N_17538);
nand U18127 (N_18127,N_17750,N_17989);
nor U18128 (N_18128,N_17757,N_17785);
and U18129 (N_18129,N_17587,N_17586);
and U18130 (N_18130,N_17822,N_17732);
nand U18131 (N_18131,N_17657,N_17776);
nand U18132 (N_18132,N_17711,N_17795);
nor U18133 (N_18133,N_17635,N_17809);
nand U18134 (N_18134,N_17829,N_17992);
or U18135 (N_18135,N_17913,N_17591);
nor U18136 (N_18136,N_17517,N_17724);
or U18137 (N_18137,N_17854,N_17606);
xnor U18138 (N_18138,N_17923,N_17847);
nor U18139 (N_18139,N_17629,N_17998);
or U18140 (N_18140,N_17532,N_17578);
nor U18141 (N_18141,N_17918,N_17893);
or U18142 (N_18142,N_17613,N_17659);
or U18143 (N_18143,N_17941,N_17833);
and U18144 (N_18144,N_17823,N_17616);
and U18145 (N_18145,N_17882,N_17876);
and U18146 (N_18146,N_17708,N_17692);
nor U18147 (N_18147,N_17600,N_17935);
or U18148 (N_18148,N_17953,N_17774);
xor U18149 (N_18149,N_17542,N_17945);
and U18150 (N_18150,N_17811,N_17899);
nor U18151 (N_18151,N_17720,N_17764);
xnor U18152 (N_18152,N_17701,N_17769);
and U18153 (N_18153,N_17727,N_17832);
nor U18154 (N_18154,N_17719,N_17557);
xnor U18155 (N_18155,N_17695,N_17892);
and U18156 (N_18156,N_17726,N_17961);
xnor U18157 (N_18157,N_17760,N_17857);
xor U18158 (N_18158,N_17921,N_17528);
nand U18159 (N_18159,N_17571,N_17723);
or U18160 (N_18160,N_17778,N_17746);
nor U18161 (N_18161,N_17827,N_17999);
and U18162 (N_18162,N_17539,N_17874);
or U18163 (N_18163,N_17521,N_17669);
or U18164 (N_18164,N_17602,N_17904);
or U18165 (N_18165,N_17703,N_17734);
or U18166 (N_18166,N_17781,N_17975);
nor U18167 (N_18167,N_17802,N_17658);
or U18168 (N_18168,N_17846,N_17869);
nand U18169 (N_18169,N_17593,N_17645);
nor U18170 (N_18170,N_17546,N_17552);
and U18171 (N_18171,N_17962,N_17910);
xnor U18172 (N_18172,N_17748,N_17971);
and U18173 (N_18173,N_17689,N_17556);
or U18174 (N_18174,N_17766,N_17661);
nand U18175 (N_18175,N_17841,N_17933);
nor U18176 (N_18176,N_17943,N_17705);
xor U18177 (N_18177,N_17668,N_17988);
nor U18178 (N_18178,N_17524,N_17675);
and U18179 (N_18179,N_17767,N_17643);
nor U18180 (N_18180,N_17927,N_17544);
nand U18181 (N_18181,N_17909,N_17549);
nor U18182 (N_18182,N_17919,N_17952);
nor U18183 (N_18183,N_17789,N_17924);
nor U18184 (N_18184,N_17806,N_17601);
nor U18185 (N_18185,N_17596,N_17634);
or U18186 (N_18186,N_17908,N_17824);
nand U18187 (N_18187,N_17572,N_17735);
and U18188 (N_18188,N_17676,N_17974);
xor U18189 (N_18189,N_17728,N_17505);
nand U18190 (N_18190,N_17867,N_17683);
nor U18191 (N_18191,N_17835,N_17799);
and U18192 (N_18192,N_17754,N_17800);
xor U18193 (N_18193,N_17576,N_17878);
or U18194 (N_18194,N_17626,N_17709);
nor U18195 (N_18195,N_17991,N_17978);
nor U18196 (N_18196,N_17947,N_17699);
or U18197 (N_18197,N_17537,N_17916);
or U18198 (N_18198,N_17837,N_17681);
nand U18199 (N_18199,N_17808,N_17906);
or U18200 (N_18200,N_17679,N_17562);
nand U18201 (N_18201,N_17958,N_17756);
and U18202 (N_18202,N_17875,N_17985);
and U18203 (N_18203,N_17523,N_17518);
or U18204 (N_18204,N_17880,N_17551);
xnor U18205 (N_18205,N_17688,N_17949);
and U18206 (N_18206,N_17545,N_17861);
nor U18207 (N_18207,N_17513,N_17599);
or U18208 (N_18208,N_17738,N_17765);
or U18209 (N_18209,N_17563,N_17637);
nor U18210 (N_18210,N_17535,N_17793);
xnor U18211 (N_18211,N_17895,N_17594);
nand U18212 (N_18212,N_17536,N_17590);
nand U18213 (N_18213,N_17644,N_17772);
nor U18214 (N_18214,N_17951,N_17603);
xor U18215 (N_18215,N_17677,N_17582);
xor U18216 (N_18216,N_17651,N_17862);
nand U18217 (N_18217,N_17983,N_17650);
xnor U18218 (N_18218,N_17502,N_17877);
and U18219 (N_18219,N_17570,N_17581);
and U18220 (N_18220,N_17632,N_17607);
nand U18221 (N_18221,N_17915,N_17987);
xnor U18222 (N_18222,N_17561,N_17610);
nand U18223 (N_18223,N_17994,N_17830);
or U18224 (N_18224,N_17559,N_17604);
or U18225 (N_18225,N_17543,N_17779);
xnor U18226 (N_18226,N_17560,N_17713);
and U18227 (N_18227,N_17533,N_17884);
nor U18228 (N_18228,N_17963,N_17930);
xor U18229 (N_18229,N_17509,N_17790);
xor U18230 (N_18230,N_17564,N_17840);
xnor U18231 (N_18231,N_17922,N_17917);
nor U18232 (N_18232,N_17928,N_17900);
nand U18233 (N_18233,N_17948,N_17577);
or U18234 (N_18234,N_17801,N_17733);
or U18235 (N_18235,N_17868,N_17697);
xnor U18236 (N_18236,N_17624,N_17967);
or U18237 (N_18237,N_17954,N_17630);
xnor U18238 (N_18238,N_17704,N_17619);
nor U18239 (N_18239,N_17647,N_17856);
and U18240 (N_18240,N_17565,N_17642);
nor U18241 (N_18241,N_17707,N_17636);
xnor U18242 (N_18242,N_17736,N_17855);
nor U18243 (N_18243,N_17839,N_17674);
and U18244 (N_18244,N_17583,N_17574);
nand U18245 (N_18245,N_17678,N_17986);
or U18246 (N_18246,N_17597,N_17797);
nor U18247 (N_18247,N_17959,N_17995);
or U18248 (N_18248,N_17655,N_17649);
and U18249 (N_18249,N_17646,N_17761);
or U18250 (N_18250,N_17509,N_17624);
nor U18251 (N_18251,N_17615,N_17944);
and U18252 (N_18252,N_17653,N_17867);
and U18253 (N_18253,N_17910,N_17967);
nor U18254 (N_18254,N_17636,N_17831);
xnor U18255 (N_18255,N_17502,N_17803);
and U18256 (N_18256,N_17553,N_17797);
nand U18257 (N_18257,N_17524,N_17561);
nor U18258 (N_18258,N_17659,N_17816);
nand U18259 (N_18259,N_17884,N_17506);
xor U18260 (N_18260,N_17538,N_17924);
or U18261 (N_18261,N_17729,N_17747);
or U18262 (N_18262,N_17908,N_17960);
nor U18263 (N_18263,N_17786,N_17997);
or U18264 (N_18264,N_17592,N_17967);
or U18265 (N_18265,N_17968,N_17529);
nand U18266 (N_18266,N_17988,N_17706);
or U18267 (N_18267,N_17848,N_17506);
nand U18268 (N_18268,N_17885,N_17653);
and U18269 (N_18269,N_17763,N_17630);
or U18270 (N_18270,N_17757,N_17650);
nor U18271 (N_18271,N_17756,N_17633);
nor U18272 (N_18272,N_17881,N_17933);
xnor U18273 (N_18273,N_17869,N_17977);
nand U18274 (N_18274,N_17533,N_17774);
nor U18275 (N_18275,N_17708,N_17966);
nand U18276 (N_18276,N_17586,N_17942);
nand U18277 (N_18277,N_17547,N_17774);
nand U18278 (N_18278,N_17508,N_17793);
and U18279 (N_18279,N_17774,N_17609);
xnor U18280 (N_18280,N_17937,N_17539);
and U18281 (N_18281,N_17596,N_17548);
and U18282 (N_18282,N_17518,N_17862);
nor U18283 (N_18283,N_17905,N_17606);
xor U18284 (N_18284,N_17717,N_17797);
or U18285 (N_18285,N_17593,N_17561);
xnor U18286 (N_18286,N_17961,N_17755);
and U18287 (N_18287,N_17960,N_17618);
or U18288 (N_18288,N_17981,N_17775);
or U18289 (N_18289,N_17778,N_17844);
or U18290 (N_18290,N_17906,N_17731);
nand U18291 (N_18291,N_17587,N_17872);
nand U18292 (N_18292,N_17566,N_17828);
nor U18293 (N_18293,N_17866,N_17899);
nor U18294 (N_18294,N_17632,N_17711);
nand U18295 (N_18295,N_17503,N_17755);
nand U18296 (N_18296,N_17955,N_17524);
nor U18297 (N_18297,N_17999,N_17768);
nor U18298 (N_18298,N_17932,N_17759);
nor U18299 (N_18299,N_17659,N_17982);
xor U18300 (N_18300,N_17991,N_17553);
xor U18301 (N_18301,N_17987,N_17893);
xor U18302 (N_18302,N_17851,N_17774);
or U18303 (N_18303,N_17915,N_17779);
xnor U18304 (N_18304,N_17935,N_17809);
nand U18305 (N_18305,N_17729,N_17598);
and U18306 (N_18306,N_17631,N_17712);
or U18307 (N_18307,N_17746,N_17523);
xnor U18308 (N_18308,N_17558,N_17935);
or U18309 (N_18309,N_17969,N_17541);
xnor U18310 (N_18310,N_17877,N_17571);
or U18311 (N_18311,N_17753,N_17554);
nand U18312 (N_18312,N_17658,N_17796);
nor U18313 (N_18313,N_17554,N_17687);
xnor U18314 (N_18314,N_17881,N_17914);
xnor U18315 (N_18315,N_17760,N_17599);
nor U18316 (N_18316,N_17921,N_17690);
or U18317 (N_18317,N_17562,N_17641);
xnor U18318 (N_18318,N_17884,N_17538);
or U18319 (N_18319,N_17520,N_17703);
nand U18320 (N_18320,N_17551,N_17745);
xor U18321 (N_18321,N_17659,N_17892);
or U18322 (N_18322,N_17646,N_17689);
and U18323 (N_18323,N_17971,N_17616);
nand U18324 (N_18324,N_17914,N_17538);
nand U18325 (N_18325,N_17665,N_17627);
nor U18326 (N_18326,N_17946,N_17616);
nor U18327 (N_18327,N_17592,N_17952);
xor U18328 (N_18328,N_17870,N_17880);
and U18329 (N_18329,N_17991,N_17819);
nor U18330 (N_18330,N_17985,N_17607);
or U18331 (N_18331,N_17887,N_17681);
and U18332 (N_18332,N_17954,N_17930);
and U18333 (N_18333,N_17750,N_17540);
or U18334 (N_18334,N_17966,N_17927);
nand U18335 (N_18335,N_17904,N_17538);
and U18336 (N_18336,N_17815,N_17968);
and U18337 (N_18337,N_17926,N_17828);
nor U18338 (N_18338,N_17801,N_17803);
nor U18339 (N_18339,N_17819,N_17596);
xor U18340 (N_18340,N_17979,N_17512);
xor U18341 (N_18341,N_17902,N_17962);
xor U18342 (N_18342,N_17913,N_17699);
nand U18343 (N_18343,N_17820,N_17803);
or U18344 (N_18344,N_17962,N_17824);
xnor U18345 (N_18345,N_17942,N_17910);
xnor U18346 (N_18346,N_17523,N_17866);
nor U18347 (N_18347,N_17599,N_17680);
and U18348 (N_18348,N_17751,N_17829);
or U18349 (N_18349,N_17810,N_17725);
nor U18350 (N_18350,N_17511,N_17789);
xnor U18351 (N_18351,N_17662,N_17561);
nor U18352 (N_18352,N_17513,N_17878);
xnor U18353 (N_18353,N_17975,N_17942);
nand U18354 (N_18354,N_17779,N_17937);
xnor U18355 (N_18355,N_17626,N_17900);
nand U18356 (N_18356,N_17549,N_17706);
nand U18357 (N_18357,N_17873,N_17804);
nor U18358 (N_18358,N_17531,N_17768);
nor U18359 (N_18359,N_17711,N_17824);
or U18360 (N_18360,N_17541,N_17781);
and U18361 (N_18361,N_17955,N_17958);
xnor U18362 (N_18362,N_17737,N_17930);
nand U18363 (N_18363,N_17563,N_17667);
nor U18364 (N_18364,N_17622,N_17682);
or U18365 (N_18365,N_17600,N_17999);
and U18366 (N_18366,N_17658,N_17806);
or U18367 (N_18367,N_17529,N_17696);
nor U18368 (N_18368,N_17651,N_17609);
or U18369 (N_18369,N_17739,N_17690);
and U18370 (N_18370,N_17742,N_17728);
or U18371 (N_18371,N_17637,N_17576);
nand U18372 (N_18372,N_17710,N_17569);
nand U18373 (N_18373,N_17841,N_17668);
nor U18374 (N_18374,N_17729,N_17615);
or U18375 (N_18375,N_17684,N_17513);
and U18376 (N_18376,N_17833,N_17903);
and U18377 (N_18377,N_17569,N_17552);
and U18378 (N_18378,N_17558,N_17972);
nor U18379 (N_18379,N_17603,N_17580);
or U18380 (N_18380,N_17977,N_17590);
nand U18381 (N_18381,N_17792,N_17685);
nor U18382 (N_18382,N_17686,N_17936);
xnor U18383 (N_18383,N_17561,N_17570);
nand U18384 (N_18384,N_17980,N_17821);
and U18385 (N_18385,N_17992,N_17746);
nand U18386 (N_18386,N_17931,N_17863);
and U18387 (N_18387,N_17601,N_17817);
nand U18388 (N_18388,N_17911,N_17932);
nand U18389 (N_18389,N_17761,N_17684);
or U18390 (N_18390,N_17699,N_17925);
nand U18391 (N_18391,N_17835,N_17514);
or U18392 (N_18392,N_17943,N_17678);
and U18393 (N_18393,N_17717,N_17649);
and U18394 (N_18394,N_17886,N_17709);
and U18395 (N_18395,N_17915,N_17830);
and U18396 (N_18396,N_17961,N_17910);
nor U18397 (N_18397,N_17543,N_17561);
nand U18398 (N_18398,N_17986,N_17731);
or U18399 (N_18399,N_17971,N_17833);
nor U18400 (N_18400,N_17548,N_17952);
nor U18401 (N_18401,N_17875,N_17789);
or U18402 (N_18402,N_17598,N_17695);
nor U18403 (N_18403,N_17650,N_17747);
and U18404 (N_18404,N_17768,N_17799);
nand U18405 (N_18405,N_17660,N_17508);
xor U18406 (N_18406,N_17841,N_17920);
and U18407 (N_18407,N_17600,N_17549);
nor U18408 (N_18408,N_17512,N_17893);
or U18409 (N_18409,N_17843,N_17618);
and U18410 (N_18410,N_17791,N_17550);
and U18411 (N_18411,N_17872,N_17557);
or U18412 (N_18412,N_17998,N_17939);
nand U18413 (N_18413,N_17802,N_17765);
nand U18414 (N_18414,N_17672,N_17852);
and U18415 (N_18415,N_17577,N_17835);
and U18416 (N_18416,N_17650,N_17715);
and U18417 (N_18417,N_17812,N_17741);
or U18418 (N_18418,N_17704,N_17887);
xor U18419 (N_18419,N_17929,N_17665);
nor U18420 (N_18420,N_17895,N_17827);
xor U18421 (N_18421,N_17501,N_17747);
and U18422 (N_18422,N_17671,N_17924);
nand U18423 (N_18423,N_17677,N_17835);
xnor U18424 (N_18424,N_17564,N_17999);
xor U18425 (N_18425,N_17700,N_17967);
xnor U18426 (N_18426,N_17541,N_17718);
nor U18427 (N_18427,N_17532,N_17512);
and U18428 (N_18428,N_17818,N_17916);
or U18429 (N_18429,N_17963,N_17571);
nand U18430 (N_18430,N_17879,N_17782);
xor U18431 (N_18431,N_17528,N_17750);
nand U18432 (N_18432,N_17501,N_17697);
xor U18433 (N_18433,N_17765,N_17526);
and U18434 (N_18434,N_17623,N_17924);
xnor U18435 (N_18435,N_17869,N_17830);
xor U18436 (N_18436,N_17563,N_17721);
and U18437 (N_18437,N_17508,N_17713);
nor U18438 (N_18438,N_17888,N_17662);
and U18439 (N_18439,N_17939,N_17520);
or U18440 (N_18440,N_17501,N_17996);
xnor U18441 (N_18441,N_17905,N_17662);
and U18442 (N_18442,N_17834,N_17711);
nand U18443 (N_18443,N_17662,N_17656);
nor U18444 (N_18444,N_17767,N_17618);
xnor U18445 (N_18445,N_17715,N_17996);
nand U18446 (N_18446,N_17642,N_17585);
nor U18447 (N_18447,N_17819,N_17544);
nand U18448 (N_18448,N_17794,N_17588);
or U18449 (N_18449,N_17780,N_17657);
nand U18450 (N_18450,N_17879,N_17527);
nor U18451 (N_18451,N_17969,N_17834);
nand U18452 (N_18452,N_17596,N_17861);
xor U18453 (N_18453,N_17672,N_17906);
nor U18454 (N_18454,N_17973,N_17955);
and U18455 (N_18455,N_17756,N_17801);
or U18456 (N_18456,N_17864,N_17704);
and U18457 (N_18457,N_17869,N_17539);
nand U18458 (N_18458,N_17548,N_17911);
nor U18459 (N_18459,N_17572,N_17882);
nand U18460 (N_18460,N_17800,N_17648);
nor U18461 (N_18461,N_17581,N_17885);
nand U18462 (N_18462,N_17505,N_17868);
and U18463 (N_18463,N_17823,N_17958);
nor U18464 (N_18464,N_17979,N_17948);
nand U18465 (N_18465,N_17801,N_17938);
nor U18466 (N_18466,N_17960,N_17503);
and U18467 (N_18467,N_17707,N_17824);
nor U18468 (N_18468,N_17752,N_17785);
and U18469 (N_18469,N_17597,N_17971);
and U18470 (N_18470,N_17982,N_17712);
and U18471 (N_18471,N_17550,N_17565);
nand U18472 (N_18472,N_17697,N_17576);
nand U18473 (N_18473,N_17997,N_17668);
nand U18474 (N_18474,N_17870,N_17855);
nand U18475 (N_18475,N_17585,N_17639);
nor U18476 (N_18476,N_17752,N_17695);
nor U18477 (N_18477,N_17618,N_17628);
and U18478 (N_18478,N_17819,N_17821);
xor U18479 (N_18479,N_17605,N_17791);
nor U18480 (N_18480,N_17653,N_17604);
nor U18481 (N_18481,N_17593,N_17508);
xnor U18482 (N_18482,N_17965,N_17836);
and U18483 (N_18483,N_17654,N_17893);
xor U18484 (N_18484,N_17543,N_17694);
nor U18485 (N_18485,N_17862,N_17726);
nand U18486 (N_18486,N_17677,N_17509);
and U18487 (N_18487,N_17859,N_17914);
xor U18488 (N_18488,N_17768,N_17729);
or U18489 (N_18489,N_17713,N_17826);
and U18490 (N_18490,N_17834,N_17550);
and U18491 (N_18491,N_17676,N_17755);
xor U18492 (N_18492,N_17615,N_17913);
nand U18493 (N_18493,N_17998,N_17559);
xnor U18494 (N_18494,N_17727,N_17918);
xnor U18495 (N_18495,N_17783,N_17918);
xor U18496 (N_18496,N_17784,N_17560);
nor U18497 (N_18497,N_17782,N_17871);
xor U18498 (N_18498,N_17512,N_17770);
nor U18499 (N_18499,N_17804,N_17823);
or U18500 (N_18500,N_18457,N_18177);
nand U18501 (N_18501,N_18057,N_18107);
and U18502 (N_18502,N_18391,N_18454);
nand U18503 (N_18503,N_18449,N_18331);
or U18504 (N_18504,N_18366,N_18039);
and U18505 (N_18505,N_18142,N_18014);
xnor U18506 (N_18506,N_18049,N_18059);
nand U18507 (N_18507,N_18072,N_18225);
and U18508 (N_18508,N_18179,N_18293);
nor U18509 (N_18509,N_18055,N_18117);
and U18510 (N_18510,N_18223,N_18497);
nand U18511 (N_18511,N_18483,N_18378);
or U18512 (N_18512,N_18489,N_18283);
xnor U18513 (N_18513,N_18292,N_18173);
xnor U18514 (N_18514,N_18328,N_18314);
or U18515 (N_18515,N_18376,N_18315);
xor U18516 (N_18516,N_18008,N_18433);
nor U18517 (N_18517,N_18069,N_18487);
xnor U18518 (N_18518,N_18037,N_18329);
or U18519 (N_18519,N_18090,N_18175);
and U18520 (N_18520,N_18320,N_18254);
xor U18521 (N_18521,N_18273,N_18446);
or U18522 (N_18522,N_18015,N_18036);
nor U18523 (N_18523,N_18056,N_18070);
nor U18524 (N_18524,N_18143,N_18369);
nor U18525 (N_18525,N_18379,N_18438);
or U18526 (N_18526,N_18176,N_18333);
and U18527 (N_18527,N_18421,N_18345);
and U18528 (N_18528,N_18127,N_18406);
or U18529 (N_18529,N_18389,N_18306);
or U18530 (N_18530,N_18208,N_18271);
or U18531 (N_18531,N_18052,N_18181);
nand U18532 (N_18532,N_18066,N_18099);
xor U18533 (N_18533,N_18250,N_18459);
and U18534 (N_18534,N_18004,N_18134);
and U18535 (N_18535,N_18397,N_18441);
and U18536 (N_18536,N_18160,N_18237);
xnor U18537 (N_18537,N_18131,N_18150);
xor U18538 (N_18538,N_18246,N_18129);
xnor U18539 (N_18539,N_18398,N_18390);
nor U18540 (N_18540,N_18182,N_18122);
or U18541 (N_18541,N_18195,N_18124);
xor U18542 (N_18542,N_18047,N_18490);
xor U18543 (N_18543,N_18388,N_18262);
and U18544 (N_18544,N_18365,N_18247);
nor U18545 (N_18545,N_18276,N_18197);
and U18546 (N_18546,N_18217,N_18227);
and U18547 (N_18547,N_18322,N_18383);
xor U18548 (N_18548,N_18432,N_18263);
xor U18549 (N_18549,N_18229,N_18327);
or U18550 (N_18550,N_18347,N_18463);
nand U18551 (N_18551,N_18111,N_18380);
nand U18552 (N_18552,N_18155,N_18042);
and U18553 (N_18553,N_18285,N_18017);
or U18554 (N_18554,N_18209,N_18447);
nor U18555 (N_18555,N_18086,N_18377);
and U18556 (N_18556,N_18058,N_18310);
and U18557 (N_18557,N_18443,N_18244);
and U18558 (N_18558,N_18470,N_18112);
or U18559 (N_18559,N_18394,N_18309);
xor U18560 (N_18560,N_18106,N_18191);
nor U18561 (N_18561,N_18005,N_18288);
xor U18562 (N_18562,N_18157,N_18230);
or U18563 (N_18563,N_18201,N_18451);
nor U18564 (N_18564,N_18027,N_18295);
xnor U18565 (N_18565,N_18499,N_18339);
nand U18566 (N_18566,N_18113,N_18171);
nand U18567 (N_18567,N_18243,N_18346);
nor U18568 (N_18568,N_18408,N_18220);
and U18569 (N_18569,N_18026,N_18105);
nor U18570 (N_18570,N_18486,N_18165);
nand U18571 (N_18571,N_18256,N_18304);
nor U18572 (N_18572,N_18172,N_18275);
or U18573 (N_18573,N_18340,N_18458);
nand U18574 (N_18574,N_18420,N_18016);
and U18575 (N_18575,N_18469,N_18030);
nand U18576 (N_18576,N_18202,N_18317);
and U18577 (N_18577,N_18279,N_18402);
nand U18578 (N_18578,N_18411,N_18481);
nand U18579 (N_18579,N_18257,N_18278);
nor U18580 (N_18580,N_18050,N_18423);
nor U18581 (N_18581,N_18401,N_18342);
xnor U18582 (N_18582,N_18405,N_18348);
nor U18583 (N_18583,N_18218,N_18410);
and U18584 (N_18584,N_18448,N_18073);
nor U18585 (N_18585,N_18232,N_18149);
and U18586 (N_18586,N_18418,N_18214);
xnor U18587 (N_18587,N_18350,N_18011);
xor U18588 (N_18588,N_18434,N_18185);
nand U18589 (N_18589,N_18084,N_18029);
nand U18590 (N_18590,N_18419,N_18159);
and U18591 (N_18591,N_18436,N_18097);
or U18592 (N_18592,N_18357,N_18137);
nand U18593 (N_18593,N_18094,N_18139);
nand U18594 (N_18594,N_18424,N_18088);
nand U18595 (N_18595,N_18362,N_18178);
and U18596 (N_18596,N_18409,N_18428);
and U18597 (N_18597,N_18242,N_18269);
xor U18598 (N_18598,N_18368,N_18071);
and U18599 (N_18599,N_18162,N_18152);
xnor U18600 (N_18600,N_18038,N_18392);
nand U18601 (N_18601,N_18248,N_18240);
and U18602 (N_18602,N_18453,N_18087);
nor U18603 (N_18603,N_18210,N_18393);
and U18604 (N_18604,N_18425,N_18298);
or U18605 (N_18605,N_18018,N_18110);
and U18606 (N_18606,N_18167,N_18450);
nor U18607 (N_18607,N_18216,N_18114);
xnor U18608 (N_18608,N_18205,N_18465);
xnor U18609 (N_18609,N_18082,N_18300);
nand U18610 (N_18610,N_18455,N_18207);
nand U18611 (N_18611,N_18341,N_18174);
nand U18612 (N_18612,N_18003,N_18031);
and U18613 (N_18613,N_18138,N_18133);
nor U18614 (N_18614,N_18062,N_18168);
nand U18615 (N_18615,N_18330,N_18277);
xnor U18616 (N_18616,N_18187,N_18266);
or U18617 (N_18617,N_18480,N_18482);
or U18618 (N_18618,N_18194,N_18102);
xnor U18619 (N_18619,N_18265,N_18060);
or U18620 (N_18620,N_18075,N_18104);
xnor U18621 (N_18621,N_18079,N_18080);
or U18622 (N_18622,N_18221,N_18032);
xor U18623 (N_18623,N_18477,N_18287);
nand U18624 (N_18624,N_18145,N_18386);
or U18625 (N_18625,N_18461,N_18065);
or U18626 (N_18626,N_18100,N_18204);
xnor U18627 (N_18627,N_18158,N_18337);
xor U18628 (N_18628,N_18170,N_18089);
xor U18629 (N_18629,N_18078,N_18395);
and U18630 (N_18630,N_18372,N_18325);
or U18631 (N_18631,N_18353,N_18198);
xnor U18632 (N_18632,N_18466,N_18123);
xnor U18633 (N_18633,N_18312,N_18280);
nand U18634 (N_18634,N_18381,N_18028);
xnor U18635 (N_18635,N_18096,N_18442);
nand U18636 (N_18636,N_18120,N_18444);
or U18637 (N_18637,N_18101,N_18282);
xnor U18638 (N_18638,N_18332,N_18196);
and U18639 (N_18639,N_18493,N_18061);
nand U18640 (N_18640,N_18146,N_18316);
or U18641 (N_18641,N_18002,N_18249);
nand U18642 (N_18642,N_18422,N_18460);
or U18643 (N_18643,N_18053,N_18296);
nor U18644 (N_18644,N_18021,N_18498);
and U18645 (N_18645,N_18313,N_18399);
nand U18646 (N_18646,N_18259,N_18351);
xor U18647 (N_18647,N_18302,N_18268);
nand U18648 (N_18648,N_18108,N_18299);
xor U18649 (N_18649,N_18374,N_18164);
nand U18650 (N_18650,N_18235,N_18251);
nor U18651 (N_18651,N_18206,N_18148);
nor U18652 (N_18652,N_18437,N_18343);
nor U18653 (N_18653,N_18462,N_18141);
xor U18654 (N_18654,N_18414,N_18153);
xor U18655 (N_18655,N_18189,N_18488);
xor U18656 (N_18656,N_18367,N_18355);
nand U18657 (N_18657,N_18128,N_18006);
nor U18658 (N_18658,N_18464,N_18404);
nor U18659 (N_18659,N_18338,N_18245);
or U18660 (N_18660,N_18478,N_18212);
or U18661 (N_18661,N_18290,N_18035);
or U18662 (N_18662,N_18067,N_18496);
nor U18663 (N_18663,N_18349,N_18126);
nand U18664 (N_18664,N_18294,N_18023);
or U18665 (N_18665,N_18334,N_18260);
and U18666 (N_18666,N_18413,N_18307);
xor U18667 (N_18667,N_18132,N_18430);
or U18668 (N_18668,N_18211,N_18284);
nor U18669 (N_18669,N_18119,N_18236);
and U18670 (N_18670,N_18479,N_18324);
xor U18671 (N_18671,N_18387,N_18321);
or U18672 (N_18672,N_18064,N_18429);
xnor U18673 (N_18673,N_18431,N_18475);
xnor U18674 (N_18674,N_18456,N_18241);
and U18675 (N_18675,N_18092,N_18311);
nor U18676 (N_18676,N_18068,N_18228);
or U18677 (N_18677,N_18103,N_18136);
nand U18678 (N_18678,N_18161,N_18001);
nor U18679 (N_18679,N_18115,N_18258);
and U18680 (N_18680,N_18130,N_18382);
xor U18681 (N_18681,N_18095,N_18024);
or U18682 (N_18682,N_18473,N_18358);
nand U18683 (N_18683,N_18091,N_18190);
and U18684 (N_18684,N_18396,N_18468);
or U18685 (N_18685,N_18233,N_18156);
xor U18686 (N_18686,N_18239,N_18494);
or U18687 (N_18687,N_18151,N_18224);
and U18688 (N_18688,N_18048,N_18435);
nand U18689 (N_18689,N_18040,N_18440);
nor U18690 (N_18690,N_18472,N_18264);
and U18691 (N_18691,N_18289,N_18360);
and U18692 (N_18692,N_18231,N_18000);
and U18693 (N_18693,N_18484,N_18354);
and U18694 (N_18694,N_18416,N_18125);
or U18695 (N_18695,N_18200,N_18274);
nand U18696 (N_18696,N_18281,N_18359);
and U18697 (N_18697,N_18012,N_18025);
or U18698 (N_18698,N_18272,N_18199);
xor U18699 (N_18699,N_18384,N_18188);
xnor U18700 (N_18700,N_18166,N_18303);
and U18701 (N_18701,N_18226,N_18184);
and U18702 (N_18702,N_18471,N_18041);
nor U18703 (N_18703,N_18163,N_18253);
nor U18704 (N_18704,N_18375,N_18118);
nor U18705 (N_18705,N_18193,N_18020);
and U18706 (N_18706,N_18407,N_18007);
xor U18707 (N_18707,N_18085,N_18043);
xor U18708 (N_18708,N_18445,N_18467);
nand U18709 (N_18709,N_18297,N_18412);
nor U18710 (N_18710,N_18252,N_18474);
nand U18711 (N_18711,N_18076,N_18364);
nand U18712 (N_18712,N_18135,N_18335);
nand U18713 (N_18713,N_18439,N_18169);
nand U18714 (N_18714,N_18051,N_18270);
and U18715 (N_18715,N_18077,N_18081);
nand U18716 (N_18716,N_18491,N_18045);
nor U18717 (N_18717,N_18054,N_18318);
or U18718 (N_18718,N_18183,N_18323);
or U18719 (N_18719,N_18009,N_18452);
or U18720 (N_18720,N_18180,N_18370);
nand U18721 (N_18721,N_18013,N_18022);
xor U18722 (N_18722,N_18385,N_18371);
nand U18723 (N_18723,N_18301,N_18033);
and U18724 (N_18724,N_18010,N_18192);
xor U18725 (N_18725,N_18234,N_18121);
xor U18726 (N_18726,N_18098,N_18485);
and U18727 (N_18727,N_18186,N_18083);
or U18728 (N_18728,N_18427,N_18109);
nand U18729 (N_18729,N_18222,N_18361);
nor U18730 (N_18730,N_18144,N_18476);
and U18731 (N_18731,N_18415,N_18019);
nand U18732 (N_18732,N_18203,N_18352);
nor U18733 (N_18733,N_18308,N_18344);
and U18734 (N_18734,N_18426,N_18215);
nand U18735 (N_18735,N_18213,N_18154);
nor U18736 (N_18736,N_18147,N_18403);
nand U18737 (N_18737,N_18116,N_18291);
or U18738 (N_18738,N_18305,N_18326);
nor U18739 (N_18739,N_18074,N_18356);
nor U18740 (N_18740,N_18363,N_18400);
nand U18741 (N_18741,N_18255,N_18373);
nand U18742 (N_18742,N_18336,N_18093);
or U18743 (N_18743,N_18495,N_18063);
or U18744 (N_18744,N_18417,N_18238);
and U18745 (N_18745,N_18492,N_18044);
nand U18746 (N_18746,N_18319,N_18034);
and U18747 (N_18747,N_18219,N_18046);
and U18748 (N_18748,N_18261,N_18286);
or U18749 (N_18749,N_18140,N_18267);
and U18750 (N_18750,N_18306,N_18310);
nand U18751 (N_18751,N_18015,N_18157);
or U18752 (N_18752,N_18007,N_18067);
or U18753 (N_18753,N_18194,N_18398);
nor U18754 (N_18754,N_18343,N_18220);
or U18755 (N_18755,N_18365,N_18232);
and U18756 (N_18756,N_18360,N_18141);
xnor U18757 (N_18757,N_18439,N_18227);
nand U18758 (N_18758,N_18402,N_18254);
or U18759 (N_18759,N_18011,N_18305);
nand U18760 (N_18760,N_18450,N_18295);
and U18761 (N_18761,N_18396,N_18435);
or U18762 (N_18762,N_18395,N_18396);
or U18763 (N_18763,N_18055,N_18405);
or U18764 (N_18764,N_18186,N_18203);
nand U18765 (N_18765,N_18477,N_18183);
and U18766 (N_18766,N_18051,N_18010);
xor U18767 (N_18767,N_18282,N_18170);
and U18768 (N_18768,N_18322,N_18292);
or U18769 (N_18769,N_18088,N_18091);
and U18770 (N_18770,N_18406,N_18335);
or U18771 (N_18771,N_18449,N_18248);
xnor U18772 (N_18772,N_18006,N_18236);
or U18773 (N_18773,N_18444,N_18427);
and U18774 (N_18774,N_18325,N_18071);
nor U18775 (N_18775,N_18471,N_18472);
xor U18776 (N_18776,N_18472,N_18035);
xnor U18777 (N_18777,N_18294,N_18481);
xnor U18778 (N_18778,N_18442,N_18220);
and U18779 (N_18779,N_18206,N_18408);
nand U18780 (N_18780,N_18089,N_18217);
nor U18781 (N_18781,N_18334,N_18348);
xor U18782 (N_18782,N_18270,N_18335);
nor U18783 (N_18783,N_18200,N_18048);
nor U18784 (N_18784,N_18223,N_18093);
nor U18785 (N_18785,N_18225,N_18456);
and U18786 (N_18786,N_18140,N_18437);
xor U18787 (N_18787,N_18406,N_18255);
xnor U18788 (N_18788,N_18136,N_18389);
nor U18789 (N_18789,N_18073,N_18278);
nand U18790 (N_18790,N_18288,N_18396);
xor U18791 (N_18791,N_18320,N_18446);
and U18792 (N_18792,N_18155,N_18114);
nand U18793 (N_18793,N_18468,N_18205);
xnor U18794 (N_18794,N_18479,N_18168);
nand U18795 (N_18795,N_18134,N_18053);
or U18796 (N_18796,N_18147,N_18065);
nor U18797 (N_18797,N_18033,N_18436);
nand U18798 (N_18798,N_18490,N_18233);
xor U18799 (N_18799,N_18301,N_18232);
xor U18800 (N_18800,N_18112,N_18171);
or U18801 (N_18801,N_18369,N_18399);
and U18802 (N_18802,N_18221,N_18182);
xnor U18803 (N_18803,N_18446,N_18248);
or U18804 (N_18804,N_18232,N_18399);
nand U18805 (N_18805,N_18283,N_18119);
or U18806 (N_18806,N_18449,N_18083);
and U18807 (N_18807,N_18119,N_18128);
nand U18808 (N_18808,N_18090,N_18068);
and U18809 (N_18809,N_18157,N_18364);
nor U18810 (N_18810,N_18109,N_18443);
and U18811 (N_18811,N_18460,N_18434);
xor U18812 (N_18812,N_18368,N_18053);
nor U18813 (N_18813,N_18272,N_18205);
nand U18814 (N_18814,N_18438,N_18156);
or U18815 (N_18815,N_18268,N_18479);
nor U18816 (N_18816,N_18303,N_18175);
nor U18817 (N_18817,N_18247,N_18452);
or U18818 (N_18818,N_18150,N_18200);
nor U18819 (N_18819,N_18007,N_18009);
or U18820 (N_18820,N_18027,N_18170);
and U18821 (N_18821,N_18394,N_18027);
or U18822 (N_18822,N_18036,N_18208);
or U18823 (N_18823,N_18200,N_18080);
nor U18824 (N_18824,N_18451,N_18157);
nor U18825 (N_18825,N_18222,N_18483);
and U18826 (N_18826,N_18109,N_18083);
nor U18827 (N_18827,N_18385,N_18357);
or U18828 (N_18828,N_18143,N_18471);
nand U18829 (N_18829,N_18451,N_18228);
nand U18830 (N_18830,N_18150,N_18002);
xor U18831 (N_18831,N_18469,N_18032);
nand U18832 (N_18832,N_18174,N_18232);
or U18833 (N_18833,N_18445,N_18176);
nor U18834 (N_18834,N_18316,N_18220);
xnor U18835 (N_18835,N_18150,N_18327);
nand U18836 (N_18836,N_18228,N_18157);
and U18837 (N_18837,N_18157,N_18327);
or U18838 (N_18838,N_18389,N_18202);
and U18839 (N_18839,N_18324,N_18041);
nor U18840 (N_18840,N_18384,N_18074);
xor U18841 (N_18841,N_18217,N_18282);
nand U18842 (N_18842,N_18354,N_18365);
xnor U18843 (N_18843,N_18100,N_18395);
nor U18844 (N_18844,N_18317,N_18248);
nor U18845 (N_18845,N_18115,N_18279);
or U18846 (N_18846,N_18152,N_18372);
xnor U18847 (N_18847,N_18364,N_18349);
nor U18848 (N_18848,N_18398,N_18097);
and U18849 (N_18849,N_18397,N_18303);
xor U18850 (N_18850,N_18479,N_18258);
and U18851 (N_18851,N_18207,N_18337);
and U18852 (N_18852,N_18419,N_18070);
nand U18853 (N_18853,N_18407,N_18278);
nor U18854 (N_18854,N_18045,N_18425);
xnor U18855 (N_18855,N_18241,N_18167);
nand U18856 (N_18856,N_18246,N_18023);
nor U18857 (N_18857,N_18036,N_18266);
and U18858 (N_18858,N_18435,N_18205);
and U18859 (N_18859,N_18297,N_18488);
nand U18860 (N_18860,N_18035,N_18234);
and U18861 (N_18861,N_18023,N_18351);
or U18862 (N_18862,N_18114,N_18275);
or U18863 (N_18863,N_18026,N_18318);
or U18864 (N_18864,N_18389,N_18011);
nand U18865 (N_18865,N_18051,N_18096);
nand U18866 (N_18866,N_18064,N_18078);
xor U18867 (N_18867,N_18476,N_18034);
xor U18868 (N_18868,N_18045,N_18415);
and U18869 (N_18869,N_18322,N_18277);
nand U18870 (N_18870,N_18023,N_18149);
xor U18871 (N_18871,N_18448,N_18419);
nor U18872 (N_18872,N_18190,N_18314);
or U18873 (N_18873,N_18301,N_18357);
and U18874 (N_18874,N_18142,N_18486);
nor U18875 (N_18875,N_18113,N_18291);
nand U18876 (N_18876,N_18203,N_18300);
nor U18877 (N_18877,N_18350,N_18050);
xor U18878 (N_18878,N_18419,N_18350);
xnor U18879 (N_18879,N_18124,N_18203);
nand U18880 (N_18880,N_18232,N_18454);
or U18881 (N_18881,N_18330,N_18347);
nand U18882 (N_18882,N_18318,N_18316);
and U18883 (N_18883,N_18385,N_18024);
nand U18884 (N_18884,N_18286,N_18119);
xor U18885 (N_18885,N_18431,N_18330);
and U18886 (N_18886,N_18094,N_18182);
and U18887 (N_18887,N_18135,N_18307);
xnor U18888 (N_18888,N_18112,N_18323);
nand U18889 (N_18889,N_18385,N_18044);
xor U18890 (N_18890,N_18374,N_18025);
and U18891 (N_18891,N_18325,N_18176);
or U18892 (N_18892,N_18228,N_18414);
nand U18893 (N_18893,N_18048,N_18275);
and U18894 (N_18894,N_18135,N_18244);
xnor U18895 (N_18895,N_18088,N_18142);
nand U18896 (N_18896,N_18435,N_18433);
xor U18897 (N_18897,N_18169,N_18409);
and U18898 (N_18898,N_18370,N_18230);
xnor U18899 (N_18899,N_18474,N_18205);
nor U18900 (N_18900,N_18166,N_18410);
nand U18901 (N_18901,N_18437,N_18019);
and U18902 (N_18902,N_18381,N_18230);
xnor U18903 (N_18903,N_18191,N_18116);
nor U18904 (N_18904,N_18170,N_18254);
and U18905 (N_18905,N_18104,N_18229);
nand U18906 (N_18906,N_18288,N_18246);
or U18907 (N_18907,N_18422,N_18329);
or U18908 (N_18908,N_18012,N_18252);
and U18909 (N_18909,N_18218,N_18244);
nand U18910 (N_18910,N_18119,N_18322);
nand U18911 (N_18911,N_18268,N_18297);
or U18912 (N_18912,N_18413,N_18473);
and U18913 (N_18913,N_18042,N_18425);
nand U18914 (N_18914,N_18390,N_18322);
nor U18915 (N_18915,N_18183,N_18321);
nor U18916 (N_18916,N_18351,N_18158);
nand U18917 (N_18917,N_18293,N_18370);
nor U18918 (N_18918,N_18296,N_18225);
xnor U18919 (N_18919,N_18395,N_18176);
nor U18920 (N_18920,N_18459,N_18219);
xnor U18921 (N_18921,N_18324,N_18480);
or U18922 (N_18922,N_18121,N_18357);
xor U18923 (N_18923,N_18162,N_18058);
and U18924 (N_18924,N_18272,N_18421);
nand U18925 (N_18925,N_18221,N_18372);
nand U18926 (N_18926,N_18360,N_18045);
nand U18927 (N_18927,N_18312,N_18250);
and U18928 (N_18928,N_18467,N_18184);
nor U18929 (N_18929,N_18400,N_18040);
nor U18930 (N_18930,N_18456,N_18434);
nand U18931 (N_18931,N_18057,N_18348);
nand U18932 (N_18932,N_18458,N_18317);
nand U18933 (N_18933,N_18197,N_18155);
or U18934 (N_18934,N_18241,N_18199);
or U18935 (N_18935,N_18405,N_18154);
and U18936 (N_18936,N_18266,N_18082);
or U18937 (N_18937,N_18130,N_18018);
nand U18938 (N_18938,N_18012,N_18042);
xnor U18939 (N_18939,N_18055,N_18113);
nor U18940 (N_18940,N_18291,N_18243);
xnor U18941 (N_18941,N_18471,N_18128);
nor U18942 (N_18942,N_18107,N_18009);
nand U18943 (N_18943,N_18374,N_18487);
nand U18944 (N_18944,N_18236,N_18027);
xnor U18945 (N_18945,N_18037,N_18306);
and U18946 (N_18946,N_18083,N_18056);
nand U18947 (N_18947,N_18094,N_18194);
and U18948 (N_18948,N_18037,N_18454);
xnor U18949 (N_18949,N_18438,N_18175);
and U18950 (N_18950,N_18216,N_18243);
nor U18951 (N_18951,N_18183,N_18232);
xor U18952 (N_18952,N_18438,N_18055);
xor U18953 (N_18953,N_18492,N_18159);
nand U18954 (N_18954,N_18280,N_18030);
and U18955 (N_18955,N_18256,N_18143);
or U18956 (N_18956,N_18257,N_18455);
xor U18957 (N_18957,N_18436,N_18157);
and U18958 (N_18958,N_18199,N_18098);
and U18959 (N_18959,N_18421,N_18338);
xnor U18960 (N_18960,N_18480,N_18367);
xnor U18961 (N_18961,N_18185,N_18000);
nor U18962 (N_18962,N_18133,N_18303);
xnor U18963 (N_18963,N_18028,N_18151);
or U18964 (N_18964,N_18205,N_18240);
nor U18965 (N_18965,N_18230,N_18403);
nand U18966 (N_18966,N_18133,N_18051);
nand U18967 (N_18967,N_18384,N_18417);
nand U18968 (N_18968,N_18240,N_18099);
nand U18969 (N_18969,N_18311,N_18025);
or U18970 (N_18970,N_18074,N_18176);
nand U18971 (N_18971,N_18456,N_18271);
nor U18972 (N_18972,N_18028,N_18497);
or U18973 (N_18973,N_18460,N_18306);
nor U18974 (N_18974,N_18013,N_18209);
xnor U18975 (N_18975,N_18248,N_18265);
nor U18976 (N_18976,N_18103,N_18222);
or U18977 (N_18977,N_18087,N_18076);
and U18978 (N_18978,N_18139,N_18192);
nor U18979 (N_18979,N_18190,N_18150);
xor U18980 (N_18980,N_18092,N_18016);
xnor U18981 (N_18981,N_18003,N_18365);
or U18982 (N_18982,N_18090,N_18127);
xor U18983 (N_18983,N_18184,N_18203);
and U18984 (N_18984,N_18059,N_18053);
or U18985 (N_18985,N_18271,N_18127);
xor U18986 (N_18986,N_18457,N_18218);
or U18987 (N_18987,N_18396,N_18187);
nor U18988 (N_18988,N_18051,N_18258);
and U18989 (N_18989,N_18159,N_18223);
nor U18990 (N_18990,N_18416,N_18481);
nand U18991 (N_18991,N_18330,N_18474);
or U18992 (N_18992,N_18359,N_18168);
xor U18993 (N_18993,N_18094,N_18465);
and U18994 (N_18994,N_18362,N_18383);
xnor U18995 (N_18995,N_18008,N_18005);
and U18996 (N_18996,N_18087,N_18221);
or U18997 (N_18997,N_18172,N_18199);
xor U18998 (N_18998,N_18234,N_18230);
and U18999 (N_18999,N_18387,N_18032);
and U19000 (N_19000,N_18913,N_18647);
nand U19001 (N_19001,N_18563,N_18974);
or U19002 (N_19002,N_18654,N_18622);
and U19003 (N_19003,N_18823,N_18729);
xnor U19004 (N_19004,N_18648,N_18676);
nand U19005 (N_19005,N_18741,N_18507);
xor U19006 (N_19006,N_18668,N_18540);
or U19007 (N_19007,N_18952,N_18776);
xor U19008 (N_19008,N_18801,N_18773);
or U19009 (N_19009,N_18617,N_18956);
xor U19010 (N_19010,N_18783,N_18626);
nand U19011 (N_19011,N_18827,N_18670);
xor U19012 (N_19012,N_18531,N_18895);
nor U19013 (N_19013,N_18559,N_18873);
nand U19014 (N_19014,N_18808,N_18708);
nand U19015 (N_19015,N_18953,N_18949);
nand U19016 (N_19016,N_18853,N_18569);
nor U19017 (N_19017,N_18565,N_18607);
nand U19018 (N_19018,N_18968,N_18574);
and U19019 (N_19019,N_18532,N_18929);
and U19020 (N_19020,N_18738,N_18810);
nand U19021 (N_19021,N_18983,N_18696);
xor U19022 (N_19022,N_18642,N_18671);
xnor U19023 (N_19023,N_18730,N_18639);
and U19024 (N_19024,N_18864,N_18751);
nand U19025 (N_19025,N_18589,N_18562);
or U19026 (N_19026,N_18637,N_18862);
nor U19027 (N_19027,N_18723,N_18971);
nand U19028 (N_19028,N_18760,N_18796);
xor U19029 (N_19029,N_18609,N_18852);
nand U19030 (N_19030,N_18807,N_18888);
nor U19031 (N_19031,N_18934,N_18917);
and U19032 (N_19032,N_18980,N_18948);
nor U19033 (N_19033,N_18533,N_18877);
and U19034 (N_19034,N_18814,N_18608);
xnor U19035 (N_19035,N_18542,N_18868);
nand U19036 (N_19036,N_18833,N_18889);
xor U19037 (N_19037,N_18904,N_18893);
nor U19038 (N_19038,N_18761,N_18580);
or U19039 (N_19039,N_18887,N_18892);
xor U19040 (N_19040,N_18746,N_18941);
xor U19041 (N_19041,N_18597,N_18970);
nor U19042 (N_19042,N_18602,N_18994);
nand U19043 (N_19043,N_18510,N_18718);
or U19044 (N_19044,N_18902,N_18899);
or U19045 (N_19045,N_18973,N_18906);
or U19046 (N_19046,N_18950,N_18963);
nand U19047 (N_19047,N_18679,N_18525);
nand U19048 (N_19048,N_18838,N_18651);
nor U19049 (N_19049,N_18727,N_18811);
and U19050 (N_19050,N_18713,N_18716);
and U19051 (N_19051,N_18988,N_18936);
nor U19052 (N_19052,N_18944,N_18615);
and U19053 (N_19053,N_18728,N_18739);
or U19054 (N_19054,N_18560,N_18744);
and U19055 (N_19055,N_18859,N_18610);
and U19056 (N_19056,N_18534,N_18969);
nor U19057 (N_19057,N_18511,N_18915);
or U19058 (N_19058,N_18835,N_18524);
xnor U19059 (N_19059,N_18619,N_18703);
and U19060 (N_19060,N_18839,N_18733);
xnor U19061 (N_19061,N_18631,N_18896);
nor U19062 (N_19062,N_18571,N_18981);
nor U19063 (N_19063,N_18630,N_18866);
nand U19064 (N_19064,N_18762,N_18914);
or U19065 (N_19065,N_18998,N_18707);
nor U19066 (N_19066,N_18678,N_18752);
and U19067 (N_19067,N_18598,N_18794);
nor U19068 (N_19068,N_18770,N_18551);
xnor U19069 (N_19069,N_18919,N_18517);
or U19070 (N_19070,N_18515,N_18684);
or U19071 (N_19071,N_18656,N_18884);
nor U19072 (N_19072,N_18621,N_18584);
xnor U19073 (N_19073,N_18557,N_18669);
or U19074 (N_19074,N_18790,N_18688);
or U19075 (N_19075,N_18771,N_18674);
nand U19076 (N_19076,N_18828,N_18965);
xnor U19077 (N_19077,N_18832,N_18673);
nand U19078 (N_19078,N_18735,N_18754);
nand U19079 (N_19079,N_18942,N_18901);
nor U19080 (N_19080,N_18659,N_18847);
nor U19081 (N_19081,N_18699,N_18529);
xor U19082 (N_19082,N_18725,N_18961);
nor U19083 (N_19083,N_18781,N_18989);
and U19084 (N_19084,N_18694,N_18613);
or U19085 (N_19085,N_18911,N_18516);
or U19086 (N_19086,N_18675,N_18795);
nand U19087 (N_19087,N_18691,N_18820);
nor U19088 (N_19088,N_18742,N_18695);
or U19089 (N_19089,N_18854,N_18863);
or U19090 (N_19090,N_18860,N_18819);
nor U19091 (N_19091,N_18528,N_18840);
and U19092 (N_19092,N_18977,N_18975);
nand U19093 (N_19093,N_18588,N_18611);
and U19094 (N_19094,N_18697,N_18652);
and U19095 (N_19095,N_18928,N_18745);
nand U19096 (N_19096,N_18653,N_18541);
and U19097 (N_19097,N_18805,N_18509);
and U19098 (N_19098,N_18712,N_18502);
and U19099 (N_19099,N_18701,N_18951);
xnor U19100 (N_19100,N_18966,N_18698);
nand U19101 (N_19101,N_18931,N_18550);
and U19102 (N_19102,N_18849,N_18851);
or U19103 (N_19103,N_18612,N_18867);
and U19104 (N_19104,N_18779,N_18908);
nor U19105 (N_19105,N_18909,N_18905);
or U19106 (N_19106,N_18797,N_18791);
or U19107 (N_19107,N_18857,N_18638);
nor U19108 (N_19108,N_18537,N_18635);
xnor U19109 (N_19109,N_18978,N_18960);
and U19110 (N_19110,N_18686,N_18883);
nor U19111 (N_19111,N_18641,N_18768);
or U19112 (N_19112,N_18806,N_18705);
and U19113 (N_19113,N_18544,N_18620);
nand U19114 (N_19114,N_18596,N_18865);
nor U19115 (N_19115,N_18690,N_18818);
xor U19116 (N_19116,N_18891,N_18660);
xor U19117 (N_19117,N_18552,N_18798);
or U19118 (N_19118,N_18880,N_18958);
and U19119 (N_19119,N_18564,N_18784);
or U19120 (N_19120,N_18848,N_18743);
or U19121 (N_19121,N_18843,N_18759);
nand U19122 (N_19122,N_18943,N_18792);
xnor U19123 (N_19123,N_18924,N_18907);
nand U19124 (N_19124,N_18526,N_18955);
nor U19125 (N_19125,N_18967,N_18603);
or U19126 (N_19126,N_18817,N_18523);
or U19127 (N_19127,N_18554,N_18527);
or U19128 (N_19128,N_18519,N_18765);
xor U19129 (N_19129,N_18926,N_18755);
nand U19130 (N_19130,N_18570,N_18549);
or U19131 (N_19131,N_18583,N_18632);
xnor U19132 (N_19132,N_18855,N_18935);
nand U19133 (N_19133,N_18578,N_18581);
and U19134 (N_19134,N_18547,N_18939);
nand U19135 (N_19135,N_18561,N_18940);
or U19136 (N_19136,N_18986,N_18719);
or U19137 (N_19137,N_18748,N_18979);
nor U19138 (N_19138,N_18772,N_18869);
xnor U19139 (N_19139,N_18655,N_18976);
and U19140 (N_19140,N_18545,N_18825);
nand U19141 (N_19141,N_18870,N_18957);
nor U19142 (N_19142,N_18558,N_18898);
nand U19143 (N_19143,N_18740,N_18831);
nor U19144 (N_19144,N_18845,N_18627);
nor U19145 (N_19145,N_18782,N_18885);
xor U19146 (N_19146,N_18769,N_18604);
and U19147 (N_19147,N_18576,N_18945);
or U19148 (N_19148,N_18645,N_18594);
or U19149 (N_19149,N_18824,N_18984);
xor U19150 (N_19150,N_18664,N_18758);
or U19151 (N_19151,N_18923,N_18927);
xor U19152 (N_19152,N_18995,N_18520);
and U19153 (N_19153,N_18681,N_18894);
or U19154 (N_19154,N_18996,N_18625);
nor U19155 (N_19155,N_18882,N_18757);
or U19156 (N_19156,N_18793,N_18658);
nand U19157 (N_19157,N_18714,N_18846);
xor U19158 (N_19158,N_18513,N_18692);
nor U19159 (N_19159,N_18592,N_18572);
and U19160 (N_19160,N_18775,N_18922);
or U19161 (N_19161,N_18937,N_18766);
nand U19162 (N_19162,N_18643,N_18932);
xnor U19163 (N_19163,N_18813,N_18579);
nand U19164 (N_19164,N_18680,N_18663);
nand U19165 (N_19165,N_18841,N_18535);
or U19166 (N_19166,N_18732,N_18590);
and U19167 (N_19167,N_18665,N_18842);
xor U19168 (N_19168,N_18777,N_18662);
or U19169 (N_19169,N_18591,N_18925);
nand U19170 (N_19170,N_18875,N_18804);
xnor U19171 (N_19171,N_18938,N_18667);
nand U19172 (N_19172,N_18556,N_18518);
xor U19173 (N_19173,N_18724,N_18717);
and U19174 (N_19174,N_18972,N_18815);
and U19175 (N_19175,N_18753,N_18715);
nor U19176 (N_19176,N_18710,N_18506);
and U19177 (N_19177,N_18990,N_18997);
or U19178 (N_19178,N_18720,N_18821);
nand U19179 (N_19179,N_18921,N_18577);
xor U19180 (N_19180,N_18543,N_18700);
xnor U19181 (N_19181,N_18872,N_18763);
nand U19182 (N_19182,N_18566,N_18644);
or U19183 (N_19183,N_18844,N_18858);
or U19184 (N_19184,N_18623,N_18897);
nand U19185 (N_19185,N_18573,N_18586);
xnor U19186 (N_19186,N_18521,N_18881);
or U19187 (N_19187,N_18764,N_18683);
and U19188 (N_19188,N_18582,N_18514);
nand U19189 (N_19189,N_18829,N_18991);
nand U19190 (N_19190,N_18685,N_18987);
nor U19191 (N_19191,N_18747,N_18546);
nor U19192 (N_19192,N_18536,N_18706);
nand U19193 (N_19193,N_18508,N_18856);
or U19194 (N_19194,N_18749,N_18780);
nor U19195 (N_19195,N_18505,N_18778);
and U19196 (N_19196,N_18916,N_18787);
or U19197 (N_19197,N_18874,N_18954);
xnor U19198 (N_19198,N_18946,N_18666);
nor U19199 (N_19199,N_18789,N_18861);
and U19200 (N_19200,N_18606,N_18734);
xnor U19201 (N_19201,N_18538,N_18910);
nor U19202 (N_19202,N_18879,N_18822);
or U19203 (N_19203,N_18830,N_18786);
nor U19204 (N_19204,N_18501,N_18585);
or U19205 (N_19205,N_18522,N_18593);
or U19206 (N_19206,N_18614,N_18568);
and U19207 (N_19207,N_18657,N_18530);
or U19208 (N_19208,N_18756,N_18918);
and U19209 (N_19209,N_18890,N_18618);
xor U19210 (N_19210,N_18736,N_18567);
and U19211 (N_19211,N_18737,N_18785);
nor U19212 (N_19212,N_18876,N_18834);
and U19213 (N_19213,N_18964,N_18687);
xnor U19214 (N_19214,N_18555,N_18799);
nor U19215 (N_19215,N_18920,N_18600);
xor U19216 (N_19216,N_18812,N_18837);
nand U19217 (N_19217,N_18702,N_18616);
or U19218 (N_19218,N_18722,N_18767);
nor U19219 (N_19219,N_18871,N_18553);
nand U19220 (N_19220,N_18512,N_18999);
xor U19221 (N_19221,N_18539,N_18504);
nand U19222 (N_19222,N_18628,N_18587);
xor U19223 (N_19223,N_18629,N_18633);
xnor U19224 (N_19224,N_18682,N_18689);
and U19225 (N_19225,N_18947,N_18634);
nor U19226 (N_19226,N_18774,N_18802);
nand U19227 (N_19227,N_18800,N_18624);
and U19228 (N_19228,N_18672,N_18646);
or U19229 (N_19229,N_18959,N_18595);
xnor U19230 (N_19230,N_18993,N_18599);
nand U19231 (N_19231,N_18982,N_18788);
nand U19232 (N_19232,N_18711,N_18601);
and U19233 (N_19233,N_18661,N_18693);
or U19234 (N_19234,N_18649,N_18677);
xor U19235 (N_19235,N_18809,N_18704);
and U19236 (N_19236,N_18850,N_18878);
xor U19237 (N_19237,N_18503,N_18650);
xnor U19238 (N_19238,N_18912,N_18962);
nor U19239 (N_19239,N_18750,N_18640);
nand U19240 (N_19240,N_18709,N_18933);
xnor U19241 (N_19241,N_18826,N_18803);
and U19242 (N_19242,N_18548,N_18605);
nor U19243 (N_19243,N_18930,N_18886);
nor U19244 (N_19244,N_18992,N_18726);
nor U19245 (N_19245,N_18985,N_18903);
nand U19246 (N_19246,N_18816,N_18575);
and U19247 (N_19247,N_18636,N_18731);
or U19248 (N_19248,N_18500,N_18900);
nor U19249 (N_19249,N_18721,N_18836);
nand U19250 (N_19250,N_18875,N_18763);
nor U19251 (N_19251,N_18982,N_18506);
and U19252 (N_19252,N_18964,N_18559);
nand U19253 (N_19253,N_18894,N_18864);
nor U19254 (N_19254,N_18934,N_18853);
nor U19255 (N_19255,N_18563,N_18512);
or U19256 (N_19256,N_18669,N_18597);
nor U19257 (N_19257,N_18505,N_18649);
nor U19258 (N_19258,N_18830,N_18516);
xnor U19259 (N_19259,N_18909,N_18613);
nor U19260 (N_19260,N_18701,N_18949);
nor U19261 (N_19261,N_18558,N_18886);
nor U19262 (N_19262,N_18804,N_18881);
xor U19263 (N_19263,N_18837,N_18889);
nand U19264 (N_19264,N_18687,N_18794);
nor U19265 (N_19265,N_18749,N_18529);
or U19266 (N_19266,N_18545,N_18866);
nor U19267 (N_19267,N_18523,N_18527);
nor U19268 (N_19268,N_18904,N_18634);
nor U19269 (N_19269,N_18940,N_18810);
and U19270 (N_19270,N_18942,N_18728);
nand U19271 (N_19271,N_18697,N_18915);
nor U19272 (N_19272,N_18518,N_18994);
nor U19273 (N_19273,N_18996,N_18785);
and U19274 (N_19274,N_18552,N_18781);
and U19275 (N_19275,N_18835,N_18617);
or U19276 (N_19276,N_18507,N_18644);
nor U19277 (N_19277,N_18766,N_18908);
or U19278 (N_19278,N_18845,N_18857);
or U19279 (N_19279,N_18649,N_18689);
or U19280 (N_19280,N_18557,N_18941);
nor U19281 (N_19281,N_18669,N_18741);
nand U19282 (N_19282,N_18554,N_18754);
and U19283 (N_19283,N_18697,N_18967);
xnor U19284 (N_19284,N_18959,N_18659);
or U19285 (N_19285,N_18597,N_18675);
or U19286 (N_19286,N_18930,N_18688);
nor U19287 (N_19287,N_18970,N_18863);
and U19288 (N_19288,N_18507,N_18613);
nand U19289 (N_19289,N_18583,N_18671);
and U19290 (N_19290,N_18558,N_18546);
xor U19291 (N_19291,N_18556,N_18683);
xor U19292 (N_19292,N_18791,N_18518);
xnor U19293 (N_19293,N_18971,N_18863);
or U19294 (N_19294,N_18514,N_18700);
xnor U19295 (N_19295,N_18841,N_18710);
or U19296 (N_19296,N_18873,N_18862);
nor U19297 (N_19297,N_18834,N_18669);
nor U19298 (N_19298,N_18950,N_18787);
nand U19299 (N_19299,N_18754,N_18771);
nand U19300 (N_19300,N_18651,N_18807);
and U19301 (N_19301,N_18844,N_18862);
nor U19302 (N_19302,N_18549,N_18785);
and U19303 (N_19303,N_18789,N_18675);
or U19304 (N_19304,N_18510,N_18838);
or U19305 (N_19305,N_18728,N_18577);
and U19306 (N_19306,N_18753,N_18956);
or U19307 (N_19307,N_18974,N_18938);
xnor U19308 (N_19308,N_18773,N_18708);
nor U19309 (N_19309,N_18870,N_18871);
or U19310 (N_19310,N_18524,N_18896);
xor U19311 (N_19311,N_18680,N_18575);
xnor U19312 (N_19312,N_18933,N_18811);
xor U19313 (N_19313,N_18819,N_18800);
nor U19314 (N_19314,N_18848,N_18870);
xnor U19315 (N_19315,N_18991,N_18811);
nand U19316 (N_19316,N_18715,N_18572);
and U19317 (N_19317,N_18555,N_18971);
nor U19318 (N_19318,N_18688,N_18523);
nand U19319 (N_19319,N_18603,N_18906);
nand U19320 (N_19320,N_18587,N_18942);
xnor U19321 (N_19321,N_18842,N_18989);
nand U19322 (N_19322,N_18689,N_18602);
nor U19323 (N_19323,N_18561,N_18982);
nand U19324 (N_19324,N_18923,N_18811);
and U19325 (N_19325,N_18839,N_18706);
nor U19326 (N_19326,N_18703,N_18689);
and U19327 (N_19327,N_18541,N_18740);
nor U19328 (N_19328,N_18850,N_18941);
nand U19329 (N_19329,N_18571,N_18591);
and U19330 (N_19330,N_18760,N_18950);
and U19331 (N_19331,N_18674,N_18538);
nand U19332 (N_19332,N_18768,N_18819);
and U19333 (N_19333,N_18761,N_18733);
or U19334 (N_19334,N_18876,N_18897);
xnor U19335 (N_19335,N_18548,N_18619);
or U19336 (N_19336,N_18713,N_18746);
xnor U19337 (N_19337,N_18736,N_18524);
and U19338 (N_19338,N_18942,N_18877);
xnor U19339 (N_19339,N_18661,N_18594);
xor U19340 (N_19340,N_18569,N_18735);
and U19341 (N_19341,N_18645,N_18903);
or U19342 (N_19342,N_18643,N_18799);
xnor U19343 (N_19343,N_18985,N_18679);
or U19344 (N_19344,N_18573,N_18589);
nor U19345 (N_19345,N_18962,N_18852);
and U19346 (N_19346,N_18993,N_18514);
or U19347 (N_19347,N_18936,N_18981);
or U19348 (N_19348,N_18623,N_18598);
xor U19349 (N_19349,N_18632,N_18699);
nor U19350 (N_19350,N_18675,N_18677);
nor U19351 (N_19351,N_18704,N_18565);
and U19352 (N_19352,N_18860,N_18955);
nand U19353 (N_19353,N_18754,N_18975);
nand U19354 (N_19354,N_18657,N_18734);
nand U19355 (N_19355,N_18611,N_18857);
xor U19356 (N_19356,N_18602,N_18738);
nand U19357 (N_19357,N_18871,N_18650);
or U19358 (N_19358,N_18761,N_18592);
nand U19359 (N_19359,N_18728,N_18641);
and U19360 (N_19360,N_18539,N_18815);
xor U19361 (N_19361,N_18904,N_18629);
xnor U19362 (N_19362,N_18627,N_18760);
or U19363 (N_19363,N_18658,N_18903);
nor U19364 (N_19364,N_18522,N_18783);
and U19365 (N_19365,N_18708,N_18850);
nor U19366 (N_19366,N_18890,N_18832);
or U19367 (N_19367,N_18514,N_18526);
xnor U19368 (N_19368,N_18714,N_18952);
or U19369 (N_19369,N_18505,N_18978);
nand U19370 (N_19370,N_18774,N_18825);
nand U19371 (N_19371,N_18563,N_18747);
or U19372 (N_19372,N_18894,N_18581);
nor U19373 (N_19373,N_18620,N_18961);
or U19374 (N_19374,N_18918,N_18815);
and U19375 (N_19375,N_18918,N_18823);
xor U19376 (N_19376,N_18515,N_18958);
and U19377 (N_19377,N_18892,N_18605);
and U19378 (N_19378,N_18503,N_18513);
or U19379 (N_19379,N_18676,N_18799);
or U19380 (N_19380,N_18673,N_18703);
or U19381 (N_19381,N_18573,N_18851);
or U19382 (N_19382,N_18958,N_18569);
xnor U19383 (N_19383,N_18638,N_18800);
nor U19384 (N_19384,N_18584,N_18934);
xor U19385 (N_19385,N_18960,N_18756);
xor U19386 (N_19386,N_18601,N_18878);
nor U19387 (N_19387,N_18515,N_18694);
nor U19388 (N_19388,N_18955,N_18986);
nor U19389 (N_19389,N_18902,N_18533);
nand U19390 (N_19390,N_18538,N_18886);
nand U19391 (N_19391,N_18570,N_18868);
nand U19392 (N_19392,N_18984,N_18843);
nor U19393 (N_19393,N_18696,N_18519);
xnor U19394 (N_19394,N_18731,N_18550);
xor U19395 (N_19395,N_18727,N_18951);
or U19396 (N_19396,N_18594,N_18665);
or U19397 (N_19397,N_18618,N_18915);
nand U19398 (N_19398,N_18603,N_18755);
and U19399 (N_19399,N_18856,N_18539);
nor U19400 (N_19400,N_18667,N_18820);
or U19401 (N_19401,N_18875,N_18635);
xor U19402 (N_19402,N_18758,N_18824);
xnor U19403 (N_19403,N_18769,N_18541);
nand U19404 (N_19404,N_18626,N_18536);
and U19405 (N_19405,N_18695,N_18711);
or U19406 (N_19406,N_18882,N_18835);
xor U19407 (N_19407,N_18741,N_18671);
or U19408 (N_19408,N_18751,N_18558);
or U19409 (N_19409,N_18944,N_18701);
nand U19410 (N_19410,N_18576,N_18517);
nand U19411 (N_19411,N_18814,N_18605);
or U19412 (N_19412,N_18969,N_18732);
nand U19413 (N_19413,N_18673,N_18914);
nand U19414 (N_19414,N_18765,N_18686);
or U19415 (N_19415,N_18694,N_18505);
nor U19416 (N_19416,N_18750,N_18889);
and U19417 (N_19417,N_18850,N_18533);
or U19418 (N_19418,N_18658,N_18921);
nor U19419 (N_19419,N_18648,N_18820);
or U19420 (N_19420,N_18516,N_18921);
nand U19421 (N_19421,N_18956,N_18588);
or U19422 (N_19422,N_18559,N_18560);
or U19423 (N_19423,N_18786,N_18939);
or U19424 (N_19424,N_18695,N_18571);
or U19425 (N_19425,N_18539,N_18831);
nor U19426 (N_19426,N_18740,N_18659);
or U19427 (N_19427,N_18956,N_18538);
nor U19428 (N_19428,N_18840,N_18595);
xnor U19429 (N_19429,N_18694,N_18684);
xor U19430 (N_19430,N_18852,N_18780);
nor U19431 (N_19431,N_18554,N_18755);
and U19432 (N_19432,N_18906,N_18843);
and U19433 (N_19433,N_18515,N_18755);
and U19434 (N_19434,N_18510,N_18921);
and U19435 (N_19435,N_18647,N_18933);
or U19436 (N_19436,N_18737,N_18534);
or U19437 (N_19437,N_18837,N_18869);
nand U19438 (N_19438,N_18978,N_18732);
xor U19439 (N_19439,N_18819,N_18745);
nor U19440 (N_19440,N_18968,N_18678);
nor U19441 (N_19441,N_18813,N_18966);
xor U19442 (N_19442,N_18748,N_18635);
and U19443 (N_19443,N_18630,N_18893);
or U19444 (N_19444,N_18701,N_18539);
xnor U19445 (N_19445,N_18614,N_18683);
xnor U19446 (N_19446,N_18517,N_18755);
or U19447 (N_19447,N_18579,N_18752);
and U19448 (N_19448,N_18579,N_18552);
nand U19449 (N_19449,N_18976,N_18703);
xor U19450 (N_19450,N_18763,N_18877);
xnor U19451 (N_19451,N_18923,N_18640);
and U19452 (N_19452,N_18765,N_18522);
nand U19453 (N_19453,N_18641,N_18628);
and U19454 (N_19454,N_18665,N_18584);
nor U19455 (N_19455,N_18787,N_18576);
xor U19456 (N_19456,N_18745,N_18622);
nor U19457 (N_19457,N_18943,N_18922);
nand U19458 (N_19458,N_18708,N_18863);
and U19459 (N_19459,N_18788,N_18817);
and U19460 (N_19460,N_18830,N_18963);
and U19461 (N_19461,N_18997,N_18994);
xnor U19462 (N_19462,N_18888,N_18728);
or U19463 (N_19463,N_18949,N_18833);
and U19464 (N_19464,N_18700,N_18866);
nand U19465 (N_19465,N_18841,N_18572);
nand U19466 (N_19466,N_18743,N_18628);
or U19467 (N_19467,N_18647,N_18636);
nor U19468 (N_19468,N_18728,N_18657);
nor U19469 (N_19469,N_18766,N_18869);
xnor U19470 (N_19470,N_18533,N_18934);
nand U19471 (N_19471,N_18624,N_18573);
or U19472 (N_19472,N_18502,N_18854);
nor U19473 (N_19473,N_18949,N_18561);
or U19474 (N_19474,N_18555,N_18731);
or U19475 (N_19475,N_18934,N_18619);
nand U19476 (N_19476,N_18637,N_18921);
nand U19477 (N_19477,N_18524,N_18621);
nand U19478 (N_19478,N_18945,N_18985);
or U19479 (N_19479,N_18643,N_18508);
and U19480 (N_19480,N_18706,N_18682);
nor U19481 (N_19481,N_18667,N_18530);
xnor U19482 (N_19482,N_18581,N_18538);
or U19483 (N_19483,N_18633,N_18638);
nand U19484 (N_19484,N_18744,N_18618);
xnor U19485 (N_19485,N_18543,N_18788);
xor U19486 (N_19486,N_18849,N_18836);
nor U19487 (N_19487,N_18803,N_18689);
or U19488 (N_19488,N_18609,N_18879);
nand U19489 (N_19489,N_18815,N_18717);
nor U19490 (N_19490,N_18623,N_18647);
nand U19491 (N_19491,N_18893,N_18770);
xor U19492 (N_19492,N_18834,N_18895);
nor U19493 (N_19493,N_18899,N_18657);
nor U19494 (N_19494,N_18961,N_18721);
xor U19495 (N_19495,N_18987,N_18863);
xor U19496 (N_19496,N_18632,N_18861);
nand U19497 (N_19497,N_18970,N_18601);
or U19498 (N_19498,N_18774,N_18980);
xnor U19499 (N_19499,N_18502,N_18764);
nand U19500 (N_19500,N_19318,N_19267);
nand U19501 (N_19501,N_19413,N_19356);
nand U19502 (N_19502,N_19423,N_19253);
nand U19503 (N_19503,N_19002,N_19308);
and U19504 (N_19504,N_19192,N_19128);
or U19505 (N_19505,N_19179,N_19204);
and U19506 (N_19506,N_19397,N_19132);
nand U19507 (N_19507,N_19355,N_19010);
and U19508 (N_19508,N_19060,N_19429);
or U19509 (N_19509,N_19035,N_19415);
nand U19510 (N_19510,N_19435,N_19233);
or U19511 (N_19511,N_19240,N_19114);
and U19512 (N_19512,N_19215,N_19218);
or U19513 (N_19513,N_19438,N_19419);
nor U19514 (N_19514,N_19069,N_19021);
nand U19515 (N_19515,N_19191,N_19012);
nand U19516 (N_19516,N_19393,N_19291);
xor U19517 (N_19517,N_19183,N_19292);
nor U19518 (N_19518,N_19156,N_19321);
or U19519 (N_19519,N_19352,N_19015);
xnor U19520 (N_19520,N_19273,N_19162);
and U19521 (N_19521,N_19259,N_19351);
xor U19522 (N_19522,N_19299,N_19470);
or U19523 (N_19523,N_19258,N_19108);
xnor U19524 (N_19524,N_19490,N_19363);
and U19525 (N_19525,N_19476,N_19357);
xor U19526 (N_19526,N_19484,N_19322);
and U19527 (N_19527,N_19123,N_19074);
or U19528 (N_19528,N_19234,N_19450);
or U19529 (N_19529,N_19383,N_19445);
and U19530 (N_19530,N_19182,N_19211);
xnor U19531 (N_19531,N_19049,N_19485);
xnor U19532 (N_19532,N_19054,N_19073);
or U19533 (N_19533,N_19288,N_19460);
nor U19534 (N_19534,N_19120,N_19311);
nor U19535 (N_19535,N_19326,N_19327);
and U19536 (N_19536,N_19214,N_19305);
or U19537 (N_19537,N_19029,N_19366);
xnor U19538 (N_19538,N_19339,N_19085);
xor U19539 (N_19539,N_19473,N_19283);
xnor U19540 (N_19540,N_19334,N_19464);
or U19541 (N_19541,N_19081,N_19125);
nor U19542 (N_19542,N_19055,N_19064);
nand U19543 (N_19543,N_19061,N_19409);
nor U19544 (N_19544,N_19011,N_19263);
or U19545 (N_19545,N_19471,N_19222);
or U19546 (N_19546,N_19377,N_19301);
or U19547 (N_19547,N_19312,N_19494);
nor U19548 (N_19548,N_19197,N_19037);
nor U19549 (N_19549,N_19406,N_19353);
and U19550 (N_19550,N_19426,N_19195);
and U19551 (N_19551,N_19082,N_19001);
or U19552 (N_19552,N_19167,N_19019);
xnor U19553 (N_19553,N_19497,N_19129);
nand U19554 (N_19554,N_19070,N_19431);
nand U19555 (N_19555,N_19480,N_19389);
nor U19556 (N_19556,N_19396,N_19294);
nor U19557 (N_19557,N_19076,N_19041);
and U19558 (N_19558,N_19401,N_19400);
and U19559 (N_19559,N_19428,N_19407);
xnor U19560 (N_19560,N_19287,N_19360);
nand U19561 (N_19561,N_19342,N_19439);
or U19562 (N_19562,N_19220,N_19372);
or U19563 (N_19563,N_19155,N_19039);
xnor U19564 (N_19564,N_19236,N_19024);
and U19565 (N_19565,N_19379,N_19455);
xor U19566 (N_19566,N_19091,N_19395);
xnor U19567 (N_19567,N_19194,N_19331);
nand U19568 (N_19568,N_19138,N_19229);
nand U19569 (N_19569,N_19141,N_19424);
and U19570 (N_19570,N_19048,N_19316);
nand U19571 (N_19571,N_19408,N_19140);
or U19572 (N_19572,N_19034,N_19149);
and U19573 (N_19573,N_19142,N_19042);
or U19574 (N_19574,N_19185,N_19254);
and U19575 (N_19575,N_19063,N_19018);
nor U19576 (N_19576,N_19340,N_19105);
xor U19577 (N_19577,N_19089,N_19119);
nor U19578 (N_19578,N_19136,N_19205);
or U19579 (N_19579,N_19153,N_19232);
nor U19580 (N_19580,N_19244,N_19038);
nor U19581 (N_19581,N_19434,N_19067);
nor U19582 (N_19582,N_19219,N_19314);
xnor U19583 (N_19583,N_19201,N_19269);
xnor U19584 (N_19584,N_19482,N_19491);
and U19585 (N_19585,N_19453,N_19371);
nand U19586 (N_19586,N_19341,N_19022);
nor U19587 (N_19587,N_19152,N_19178);
or U19588 (N_19588,N_19370,N_19184);
xnor U19589 (N_19589,N_19248,N_19096);
nand U19590 (N_19590,N_19422,N_19092);
or U19591 (N_19591,N_19157,N_19378);
xnor U19592 (N_19592,N_19416,N_19242);
or U19593 (N_19593,N_19007,N_19225);
xor U19594 (N_19594,N_19499,N_19040);
and U19595 (N_19595,N_19104,N_19452);
and U19596 (N_19596,N_19264,N_19032);
nor U19597 (N_19597,N_19079,N_19087);
nor U19598 (N_19598,N_19297,N_19093);
xor U19599 (N_19599,N_19243,N_19000);
xor U19600 (N_19600,N_19386,N_19295);
nand U19601 (N_19601,N_19112,N_19493);
nor U19602 (N_19602,N_19097,N_19320);
nor U19603 (N_19603,N_19373,N_19062);
and U19604 (N_19604,N_19255,N_19090);
or U19605 (N_19605,N_19492,N_19375);
nand U19606 (N_19606,N_19210,N_19025);
or U19607 (N_19607,N_19173,N_19381);
xnor U19608 (N_19608,N_19053,N_19442);
xnor U19609 (N_19609,N_19465,N_19349);
nor U19610 (N_19610,N_19056,N_19005);
nand U19611 (N_19611,N_19071,N_19475);
nand U19612 (N_19612,N_19279,N_19262);
xnor U19613 (N_19613,N_19190,N_19080);
nand U19614 (N_19614,N_19016,N_19148);
nor U19615 (N_19615,N_19134,N_19151);
and U19616 (N_19616,N_19221,N_19425);
nand U19617 (N_19617,N_19083,N_19354);
nor U19618 (N_19618,N_19247,N_19391);
xnor U19619 (N_19619,N_19365,N_19177);
nand U19620 (N_19620,N_19402,N_19223);
xor U19621 (N_19621,N_19382,N_19325);
xnor U19622 (N_19622,N_19266,N_19059);
nand U19623 (N_19623,N_19137,N_19293);
nand U19624 (N_19624,N_19447,N_19224);
nor U19625 (N_19625,N_19454,N_19043);
and U19626 (N_19626,N_19216,N_19446);
nor U19627 (N_19627,N_19203,N_19186);
nor U19628 (N_19628,N_19239,N_19282);
nand U19629 (N_19629,N_19394,N_19169);
or U19630 (N_19630,N_19489,N_19324);
xor U19631 (N_19631,N_19147,N_19417);
nand U19632 (N_19632,N_19472,N_19033);
nand U19633 (N_19633,N_19166,N_19066);
or U19634 (N_19634,N_19433,N_19376);
or U19635 (N_19635,N_19346,N_19461);
and U19636 (N_19636,N_19335,N_19101);
and U19637 (N_19637,N_19020,N_19006);
nand U19638 (N_19638,N_19348,N_19468);
and U19639 (N_19639,N_19296,N_19458);
and U19640 (N_19640,N_19046,N_19130);
nor U19641 (N_19641,N_19367,N_19388);
or U19642 (N_19642,N_19026,N_19380);
nor U19643 (N_19643,N_19171,N_19337);
and U19644 (N_19644,N_19170,N_19483);
nand U19645 (N_19645,N_19250,N_19462);
and U19646 (N_19646,N_19289,N_19168);
nor U19647 (N_19647,N_19004,N_19017);
nand U19648 (N_19648,N_19014,N_19068);
and U19649 (N_19649,N_19304,N_19481);
or U19650 (N_19650,N_19095,N_19106);
or U19651 (N_19651,N_19237,N_19044);
nor U19652 (N_19652,N_19172,N_19256);
nand U19653 (N_19653,N_19030,N_19414);
or U19654 (N_19654,N_19281,N_19023);
nand U19655 (N_19655,N_19418,N_19175);
and U19656 (N_19656,N_19109,N_19474);
or U19657 (N_19657,N_19338,N_19193);
nor U19658 (N_19658,N_19495,N_19051);
nand U19659 (N_19659,N_19487,N_19084);
and U19660 (N_19660,N_19275,N_19350);
nand U19661 (N_19661,N_19217,N_19440);
xnor U19662 (N_19662,N_19159,N_19078);
and U19663 (N_19663,N_19163,N_19496);
xnor U19664 (N_19664,N_19075,N_19052);
xnor U19665 (N_19665,N_19072,N_19412);
and U19666 (N_19666,N_19143,N_19031);
xnor U19667 (N_19667,N_19276,N_19261);
and U19668 (N_19668,N_19241,N_19303);
nand U19669 (N_19669,N_19045,N_19307);
xnor U19670 (N_19670,N_19477,N_19430);
nand U19671 (N_19671,N_19306,N_19404);
and U19672 (N_19672,N_19459,N_19336);
or U19673 (N_19673,N_19027,N_19405);
nand U19674 (N_19674,N_19399,N_19479);
xnor U19675 (N_19675,N_19347,N_19116);
and U19676 (N_19676,N_19124,N_19309);
nor U19677 (N_19677,N_19113,N_19420);
nand U19678 (N_19678,N_19364,N_19121);
nor U19679 (N_19679,N_19209,N_19328);
nor U19680 (N_19680,N_19368,N_19126);
xnor U19681 (N_19681,N_19131,N_19207);
nor U19682 (N_19682,N_19392,N_19107);
or U19683 (N_19683,N_19127,N_19238);
and U19684 (N_19684,N_19013,N_19317);
and U19685 (N_19685,N_19421,N_19290);
and U19686 (N_19686,N_19286,N_19298);
or U19687 (N_19687,N_19199,N_19047);
nor U19688 (N_19688,N_19160,N_19036);
nand U19689 (N_19689,N_19135,N_19174);
or U19690 (N_19690,N_19231,N_19161);
nand U19691 (N_19691,N_19164,N_19427);
xor U19692 (N_19692,N_19362,N_19226);
nor U19693 (N_19693,N_19150,N_19154);
nand U19694 (N_19694,N_19227,N_19385);
and U19695 (N_19695,N_19246,N_19486);
xnor U19696 (N_19696,N_19181,N_19488);
nand U19697 (N_19697,N_19330,N_19088);
nand U19698 (N_19698,N_19198,N_19272);
and U19699 (N_19699,N_19323,N_19249);
xor U19700 (N_19700,N_19099,N_19274);
or U19701 (N_19701,N_19103,N_19384);
and U19702 (N_19702,N_19189,N_19111);
nand U19703 (N_19703,N_19457,N_19102);
and U19704 (N_19704,N_19456,N_19300);
nor U19705 (N_19705,N_19268,N_19009);
and U19706 (N_19706,N_19100,N_19230);
and U19707 (N_19707,N_19165,N_19398);
nand U19708 (N_19708,N_19333,N_19110);
nand U19709 (N_19709,N_19315,N_19098);
or U19710 (N_19710,N_19122,N_19369);
nand U19711 (N_19711,N_19278,N_19213);
nand U19712 (N_19712,N_19478,N_19358);
or U19713 (N_19713,N_19146,N_19065);
nor U19714 (N_19714,N_19390,N_19361);
or U19715 (N_19715,N_19228,N_19245);
or U19716 (N_19716,N_19271,N_19437);
xnor U19717 (N_19717,N_19319,N_19374);
nand U19718 (N_19718,N_19188,N_19432);
or U19719 (N_19719,N_19206,N_19345);
or U19720 (N_19720,N_19008,N_19212);
nor U19721 (N_19721,N_19094,N_19077);
xor U19722 (N_19722,N_19410,N_19448);
nand U19723 (N_19723,N_19118,N_19176);
nand U19724 (N_19724,N_19202,N_19252);
nor U19725 (N_19725,N_19436,N_19028);
xor U19726 (N_19726,N_19050,N_19277);
nand U19727 (N_19727,N_19313,N_19449);
and U19728 (N_19728,N_19145,N_19251);
nand U19729 (N_19729,N_19208,N_19284);
and U19730 (N_19730,N_19003,N_19411);
xor U19731 (N_19731,N_19498,N_19344);
nand U19732 (N_19732,N_19463,N_19466);
xor U19733 (N_19733,N_19467,N_19444);
xnor U19734 (N_19734,N_19196,N_19115);
and U19735 (N_19735,N_19187,N_19270);
xnor U19736 (N_19736,N_19280,N_19200);
nand U19737 (N_19737,N_19260,N_19285);
xor U19738 (N_19738,N_19469,N_19343);
nor U19739 (N_19739,N_19387,N_19158);
nand U19740 (N_19740,N_19057,N_19332);
nand U19741 (N_19741,N_19403,N_19329);
xor U19742 (N_19742,N_19302,N_19139);
xnor U19743 (N_19743,N_19441,N_19359);
nand U19744 (N_19744,N_19117,N_19086);
xor U19745 (N_19745,N_19443,N_19235);
nand U19746 (N_19746,N_19180,N_19451);
nand U19747 (N_19747,N_19133,N_19058);
or U19748 (N_19748,N_19144,N_19310);
and U19749 (N_19749,N_19265,N_19257);
or U19750 (N_19750,N_19445,N_19432);
xor U19751 (N_19751,N_19121,N_19040);
and U19752 (N_19752,N_19144,N_19120);
nor U19753 (N_19753,N_19483,N_19435);
xnor U19754 (N_19754,N_19251,N_19174);
nand U19755 (N_19755,N_19239,N_19140);
xnor U19756 (N_19756,N_19457,N_19402);
nor U19757 (N_19757,N_19214,N_19401);
nor U19758 (N_19758,N_19431,N_19039);
and U19759 (N_19759,N_19288,N_19046);
nand U19760 (N_19760,N_19268,N_19465);
nand U19761 (N_19761,N_19023,N_19325);
nand U19762 (N_19762,N_19005,N_19425);
xnor U19763 (N_19763,N_19135,N_19185);
or U19764 (N_19764,N_19025,N_19440);
nor U19765 (N_19765,N_19202,N_19400);
and U19766 (N_19766,N_19265,N_19078);
xnor U19767 (N_19767,N_19442,N_19014);
and U19768 (N_19768,N_19031,N_19430);
or U19769 (N_19769,N_19090,N_19295);
nor U19770 (N_19770,N_19379,N_19063);
nand U19771 (N_19771,N_19335,N_19209);
nand U19772 (N_19772,N_19061,N_19439);
xnor U19773 (N_19773,N_19007,N_19314);
nor U19774 (N_19774,N_19189,N_19411);
xor U19775 (N_19775,N_19000,N_19117);
or U19776 (N_19776,N_19076,N_19281);
xor U19777 (N_19777,N_19397,N_19416);
xor U19778 (N_19778,N_19060,N_19349);
or U19779 (N_19779,N_19293,N_19263);
nand U19780 (N_19780,N_19026,N_19303);
and U19781 (N_19781,N_19330,N_19161);
or U19782 (N_19782,N_19187,N_19366);
xnor U19783 (N_19783,N_19260,N_19272);
and U19784 (N_19784,N_19038,N_19075);
xor U19785 (N_19785,N_19115,N_19420);
nor U19786 (N_19786,N_19327,N_19021);
xnor U19787 (N_19787,N_19034,N_19297);
xnor U19788 (N_19788,N_19057,N_19211);
or U19789 (N_19789,N_19474,N_19399);
nand U19790 (N_19790,N_19395,N_19185);
xnor U19791 (N_19791,N_19193,N_19452);
xor U19792 (N_19792,N_19028,N_19279);
nor U19793 (N_19793,N_19273,N_19262);
nand U19794 (N_19794,N_19496,N_19345);
or U19795 (N_19795,N_19211,N_19126);
and U19796 (N_19796,N_19305,N_19210);
xnor U19797 (N_19797,N_19430,N_19484);
and U19798 (N_19798,N_19295,N_19424);
nor U19799 (N_19799,N_19227,N_19414);
xor U19800 (N_19800,N_19254,N_19335);
or U19801 (N_19801,N_19156,N_19043);
nor U19802 (N_19802,N_19489,N_19199);
and U19803 (N_19803,N_19240,N_19061);
and U19804 (N_19804,N_19415,N_19258);
nor U19805 (N_19805,N_19150,N_19219);
or U19806 (N_19806,N_19161,N_19062);
nand U19807 (N_19807,N_19021,N_19355);
nand U19808 (N_19808,N_19039,N_19269);
nand U19809 (N_19809,N_19188,N_19184);
xnor U19810 (N_19810,N_19103,N_19327);
and U19811 (N_19811,N_19438,N_19110);
nor U19812 (N_19812,N_19320,N_19494);
or U19813 (N_19813,N_19313,N_19128);
nor U19814 (N_19814,N_19474,N_19460);
nand U19815 (N_19815,N_19239,N_19129);
nand U19816 (N_19816,N_19371,N_19173);
and U19817 (N_19817,N_19253,N_19490);
or U19818 (N_19818,N_19372,N_19213);
nand U19819 (N_19819,N_19067,N_19002);
nand U19820 (N_19820,N_19451,N_19329);
or U19821 (N_19821,N_19277,N_19080);
nand U19822 (N_19822,N_19427,N_19373);
xnor U19823 (N_19823,N_19095,N_19468);
nand U19824 (N_19824,N_19090,N_19187);
nor U19825 (N_19825,N_19059,N_19464);
and U19826 (N_19826,N_19498,N_19401);
xor U19827 (N_19827,N_19167,N_19356);
nand U19828 (N_19828,N_19477,N_19262);
and U19829 (N_19829,N_19352,N_19451);
xnor U19830 (N_19830,N_19009,N_19156);
nand U19831 (N_19831,N_19154,N_19119);
xnor U19832 (N_19832,N_19289,N_19181);
nor U19833 (N_19833,N_19480,N_19269);
and U19834 (N_19834,N_19244,N_19227);
or U19835 (N_19835,N_19221,N_19412);
nor U19836 (N_19836,N_19272,N_19347);
and U19837 (N_19837,N_19462,N_19252);
or U19838 (N_19838,N_19444,N_19107);
or U19839 (N_19839,N_19333,N_19395);
or U19840 (N_19840,N_19486,N_19361);
nor U19841 (N_19841,N_19160,N_19349);
nor U19842 (N_19842,N_19315,N_19429);
xor U19843 (N_19843,N_19275,N_19115);
nand U19844 (N_19844,N_19005,N_19488);
nor U19845 (N_19845,N_19337,N_19008);
or U19846 (N_19846,N_19167,N_19164);
and U19847 (N_19847,N_19035,N_19379);
xor U19848 (N_19848,N_19252,N_19017);
and U19849 (N_19849,N_19396,N_19430);
xnor U19850 (N_19850,N_19492,N_19388);
and U19851 (N_19851,N_19119,N_19366);
nand U19852 (N_19852,N_19105,N_19241);
or U19853 (N_19853,N_19086,N_19284);
nand U19854 (N_19854,N_19344,N_19483);
nor U19855 (N_19855,N_19411,N_19359);
or U19856 (N_19856,N_19257,N_19014);
xor U19857 (N_19857,N_19080,N_19027);
or U19858 (N_19858,N_19289,N_19308);
or U19859 (N_19859,N_19135,N_19117);
and U19860 (N_19860,N_19174,N_19499);
nor U19861 (N_19861,N_19489,N_19354);
or U19862 (N_19862,N_19097,N_19178);
and U19863 (N_19863,N_19216,N_19135);
nor U19864 (N_19864,N_19236,N_19015);
nor U19865 (N_19865,N_19150,N_19273);
and U19866 (N_19866,N_19337,N_19382);
or U19867 (N_19867,N_19127,N_19336);
nor U19868 (N_19868,N_19169,N_19485);
nand U19869 (N_19869,N_19199,N_19480);
and U19870 (N_19870,N_19226,N_19407);
and U19871 (N_19871,N_19382,N_19131);
and U19872 (N_19872,N_19005,N_19131);
nor U19873 (N_19873,N_19281,N_19354);
and U19874 (N_19874,N_19222,N_19091);
or U19875 (N_19875,N_19497,N_19398);
and U19876 (N_19876,N_19282,N_19336);
nand U19877 (N_19877,N_19320,N_19086);
nor U19878 (N_19878,N_19146,N_19148);
xnor U19879 (N_19879,N_19355,N_19221);
nor U19880 (N_19880,N_19155,N_19032);
nand U19881 (N_19881,N_19429,N_19412);
and U19882 (N_19882,N_19399,N_19252);
or U19883 (N_19883,N_19120,N_19471);
xor U19884 (N_19884,N_19215,N_19235);
or U19885 (N_19885,N_19208,N_19191);
or U19886 (N_19886,N_19348,N_19260);
nor U19887 (N_19887,N_19445,N_19007);
nor U19888 (N_19888,N_19113,N_19018);
nand U19889 (N_19889,N_19132,N_19067);
and U19890 (N_19890,N_19494,N_19399);
nor U19891 (N_19891,N_19374,N_19465);
xnor U19892 (N_19892,N_19481,N_19037);
nand U19893 (N_19893,N_19017,N_19450);
nor U19894 (N_19894,N_19142,N_19215);
or U19895 (N_19895,N_19021,N_19247);
nand U19896 (N_19896,N_19324,N_19025);
nand U19897 (N_19897,N_19457,N_19465);
or U19898 (N_19898,N_19269,N_19261);
and U19899 (N_19899,N_19262,N_19019);
nor U19900 (N_19900,N_19430,N_19482);
and U19901 (N_19901,N_19196,N_19328);
nand U19902 (N_19902,N_19155,N_19161);
xnor U19903 (N_19903,N_19382,N_19355);
nor U19904 (N_19904,N_19122,N_19415);
xor U19905 (N_19905,N_19329,N_19254);
xor U19906 (N_19906,N_19307,N_19180);
or U19907 (N_19907,N_19495,N_19289);
or U19908 (N_19908,N_19241,N_19115);
or U19909 (N_19909,N_19471,N_19445);
nor U19910 (N_19910,N_19199,N_19152);
or U19911 (N_19911,N_19291,N_19363);
nand U19912 (N_19912,N_19159,N_19089);
nand U19913 (N_19913,N_19125,N_19498);
nand U19914 (N_19914,N_19150,N_19485);
nand U19915 (N_19915,N_19403,N_19474);
nor U19916 (N_19916,N_19368,N_19333);
nor U19917 (N_19917,N_19400,N_19148);
and U19918 (N_19918,N_19199,N_19053);
nor U19919 (N_19919,N_19163,N_19018);
or U19920 (N_19920,N_19051,N_19187);
nand U19921 (N_19921,N_19199,N_19419);
and U19922 (N_19922,N_19228,N_19213);
or U19923 (N_19923,N_19183,N_19443);
and U19924 (N_19924,N_19307,N_19016);
or U19925 (N_19925,N_19384,N_19362);
or U19926 (N_19926,N_19422,N_19022);
and U19927 (N_19927,N_19106,N_19207);
or U19928 (N_19928,N_19271,N_19047);
nand U19929 (N_19929,N_19319,N_19000);
nor U19930 (N_19930,N_19256,N_19116);
xor U19931 (N_19931,N_19004,N_19062);
or U19932 (N_19932,N_19253,N_19159);
or U19933 (N_19933,N_19168,N_19255);
xor U19934 (N_19934,N_19260,N_19028);
and U19935 (N_19935,N_19233,N_19227);
nor U19936 (N_19936,N_19088,N_19129);
and U19937 (N_19937,N_19002,N_19309);
nor U19938 (N_19938,N_19275,N_19243);
and U19939 (N_19939,N_19437,N_19467);
and U19940 (N_19940,N_19348,N_19433);
and U19941 (N_19941,N_19229,N_19266);
or U19942 (N_19942,N_19157,N_19054);
xnor U19943 (N_19943,N_19058,N_19266);
or U19944 (N_19944,N_19175,N_19327);
xnor U19945 (N_19945,N_19180,N_19175);
xnor U19946 (N_19946,N_19478,N_19104);
and U19947 (N_19947,N_19291,N_19064);
and U19948 (N_19948,N_19311,N_19245);
or U19949 (N_19949,N_19499,N_19279);
xnor U19950 (N_19950,N_19280,N_19318);
and U19951 (N_19951,N_19156,N_19174);
or U19952 (N_19952,N_19069,N_19390);
and U19953 (N_19953,N_19009,N_19173);
xor U19954 (N_19954,N_19030,N_19184);
and U19955 (N_19955,N_19054,N_19245);
nor U19956 (N_19956,N_19109,N_19169);
and U19957 (N_19957,N_19053,N_19111);
nand U19958 (N_19958,N_19396,N_19076);
or U19959 (N_19959,N_19212,N_19477);
and U19960 (N_19960,N_19225,N_19132);
nand U19961 (N_19961,N_19399,N_19012);
or U19962 (N_19962,N_19227,N_19327);
xnor U19963 (N_19963,N_19055,N_19292);
xor U19964 (N_19964,N_19270,N_19028);
and U19965 (N_19965,N_19348,N_19301);
nand U19966 (N_19966,N_19337,N_19329);
nor U19967 (N_19967,N_19362,N_19461);
and U19968 (N_19968,N_19188,N_19394);
xor U19969 (N_19969,N_19274,N_19235);
xor U19970 (N_19970,N_19145,N_19027);
nand U19971 (N_19971,N_19142,N_19127);
xor U19972 (N_19972,N_19307,N_19370);
nor U19973 (N_19973,N_19014,N_19071);
nor U19974 (N_19974,N_19084,N_19154);
or U19975 (N_19975,N_19457,N_19291);
nand U19976 (N_19976,N_19186,N_19000);
and U19977 (N_19977,N_19027,N_19221);
or U19978 (N_19978,N_19252,N_19080);
xor U19979 (N_19979,N_19210,N_19218);
or U19980 (N_19980,N_19064,N_19306);
and U19981 (N_19981,N_19449,N_19061);
nand U19982 (N_19982,N_19112,N_19161);
nor U19983 (N_19983,N_19319,N_19444);
xnor U19984 (N_19984,N_19148,N_19272);
nor U19985 (N_19985,N_19017,N_19388);
nand U19986 (N_19986,N_19251,N_19086);
or U19987 (N_19987,N_19027,N_19092);
xnor U19988 (N_19988,N_19334,N_19243);
or U19989 (N_19989,N_19264,N_19164);
nand U19990 (N_19990,N_19121,N_19105);
nor U19991 (N_19991,N_19475,N_19168);
nor U19992 (N_19992,N_19256,N_19399);
or U19993 (N_19993,N_19263,N_19326);
or U19994 (N_19994,N_19446,N_19082);
and U19995 (N_19995,N_19142,N_19436);
or U19996 (N_19996,N_19040,N_19443);
and U19997 (N_19997,N_19024,N_19336);
nor U19998 (N_19998,N_19230,N_19232);
xor U19999 (N_19999,N_19443,N_19456);
nand U20000 (N_20000,N_19667,N_19977);
nor U20001 (N_20001,N_19980,N_19922);
and U20002 (N_20002,N_19966,N_19801);
nand U20003 (N_20003,N_19893,N_19989);
xnor U20004 (N_20004,N_19639,N_19759);
nor U20005 (N_20005,N_19779,N_19994);
and U20006 (N_20006,N_19552,N_19656);
and U20007 (N_20007,N_19988,N_19903);
xnor U20008 (N_20008,N_19682,N_19769);
or U20009 (N_20009,N_19685,N_19756);
xnor U20010 (N_20010,N_19723,N_19590);
nand U20011 (N_20011,N_19679,N_19666);
nor U20012 (N_20012,N_19613,N_19974);
and U20013 (N_20013,N_19939,N_19703);
nor U20014 (N_20014,N_19500,N_19617);
and U20015 (N_20015,N_19586,N_19529);
or U20016 (N_20016,N_19565,N_19564);
xnor U20017 (N_20017,N_19884,N_19715);
nor U20018 (N_20018,N_19580,N_19844);
and U20019 (N_20019,N_19936,N_19768);
xor U20020 (N_20020,N_19686,N_19897);
xor U20021 (N_20021,N_19864,N_19584);
xnor U20022 (N_20022,N_19751,N_19694);
xnor U20023 (N_20023,N_19971,N_19691);
or U20024 (N_20024,N_19985,N_19910);
xor U20025 (N_20025,N_19585,N_19662);
nand U20026 (N_20026,N_19536,N_19889);
or U20027 (N_20027,N_19963,N_19752);
and U20028 (N_20028,N_19891,N_19876);
nor U20029 (N_20029,N_19962,N_19815);
xnor U20030 (N_20030,N_19938,N_19842);
or U20031 (N_20031,N_19803,N_19986);
or U20032 (N_20032,N_19537,N_19885);
and U20033 (N_20033,N_19643,N_19792);
or U20034 (N_20034,N_19758,N_19961);
and U20035 (N_20035,N_19736,N_19941);
nor U20036 (N_20036,N_19784,N_19557);
or U20037 (N_20037,N_19507,N_19787);
xnor U20038 (N_20038,N_19550,N_19589);
nor U20039 (N_20039,N_19735,N_19840);
xnor U20040 (N_20040,N_19834,N_19932);
or U20041 (N_20041,N_19942,N_19785);
xnor U20042 (N_20042,N_19622,N_19970);
or U20043 (N_20043,N_19947,N_19604);
or U20044 (N_20044,N_19503,N_19722);
nor U20045 (N_20045,N_19850,N_19919);
or U20046 (N_20046,N_19866,N_19553);
nand U20047 (N_20047,N_19821,N_19531);
or U20048 (N_20048,N_19514,N_19915);
or U20049 (N_20049,N_19773,N_19510);
and U20050 (N_20050,N_19664,N_19865);
nand U20051 (N_20051,N_19807,N_19581);
or U20052 (N_20052,N_19601,N_19765);
and U20053 (N_20053,N_19778,N_19771);
nand U20054 (N_20054,N_19518,N_19506);
and U20055 (N_20055,N_19804,N_19766);
and U20056 (N_20056,N_19798,N_19599);
xnor U20057 (N_20057,N_19588,N_19653);
and U20058 (N_20058,N_19764,N_19859);
nand U20059 (N_20059,N_19567,N_19505);
xor U20060 (N_20060,N_19946,N_19772);
nand U20061 (N_20061,N_19857,N_19576);
or U20062 (N_20062,N_19502,N_19517);
nand U20063 (N_20063,N_19727,N_19888);
nand U20064 (N_20064,N_19848,N_19992);
nor U20065 (N_20065,N_19657,N_19862);
nor U20066 (N_20066,N_19949,N_19647);
xor U20067 (N_20067,N_19923,N_19693);
and U20068 (N_20068,N_19627,N_19526);
or U20069 (N_20069,N_19561,N_19654);
and U20070 (N_20070,N_19563,N_19539);
xor U20071 (N_20071,N_19912,N_19650);
or U20072 (N_20072,N_19943,N_19770);
and U20073 (N_20073,N_19721,N_19661);
or U20074 (N_20074,N_19595,N_19515);
or U20075 (N_20075,N_19849,N_19806);
or U20076 (N_20076,N_19976,N_19959);
nand U20077 (N_20077,N_19556,N_19729);
or U20078 (N_20078,N_19763,N_19958);
or U20079 (N_20079,N_19991,N_19794);
nor U20080 (N_20080,N_19838,N_19695);
and U20081 (N_20081,N_19819,N_19973);
or U20082 (N_20082,N_19737,N_19892);
and U20083 (N_20083,N_19718,N_19600);
nor U20084 (N_20084,N_19810,N_19609);
nor U20085 (N_20085,N_19931,N_19578);
and U20086 (N_20086,N_19641,N_19835);
xnor U20087 (N_20087,N_19987,N_19545);
nand U20088 (N_20088,N_19908,N_19605);
or U20089 (N_20089,N_19720,N_19619);
nor U20090 (N_20090,N_19624,N_19504);
or U20091 (N_20091,N_19603,N_19791);
nor U20092 (N_20092,N_19559,N_19937);
xnor U20093 (N_20093,N_19646,N_19786);
or U20094 (N_20094,N_19861,N_19684);
xnor U20095 (N_20095,N_19816,N_19548);
and U20096 (N_20096,N_19955,N_19725);
nand U20097 (N_20097,N_19614,N_19841);
xnor U20098 (N_20098,N_19978,N_19879);
nand U20099 (N_20099,N_19696,N_19761);
xor U20100 (N_20100,N_19640,N_19520);
and U20101 (N_20101,N_19812,N_19793);
or U20102 (N_20102,N_19890,N_19728);
xnor U20103 (N_20103,N_19621,N_19530);
and U20104 (N_20104,N_19633,N_19607);
xnor U20105 (N_20105,N_19521,N_19512);
nor U20106 (N_20106,N_19832,N_19523);
nand U20107 (N_20107,N_19555,N_19571);
and U20108 (N_20108,N_19837,N_19524);
xor U20109 (N_20109,N_19707,N_19940);
nor U20110 (N_20110,N_19975,N_19896);
or U20111 (N_20111,N_19540,N_19683);
nor U20112 (N_20112,N_19809,N_19926);
xnor U20113 (N_20113,N_19511,N_19533);
nor U20114 (N_20114,N_19928,N_19655);
or U20115 (N_20115,N_19914,N_19620);
xor U20116 (N_20116,N_19731,N_19598);
xnor U20117 (N_20117,N_19984,N_19541);
or U20118 (N_20118,N_19706,N_19566);
and U20119 (N_20119,N_19826,N_19870);
nand U20120 (N_20120,N_19636,N_19847);
and U20121 (N_20121,N_19558,N_19519);
or U20122 (N_20122,N_19960,N_19630);
or U20123 (N_20123,N_19795,N_19573);
nand U20124 (N_20124,N_19920,N_19790);
or U20125 (N_20125,N_19674,N_19574);
and U20126 (N_20126,N_19659,N_19734);
nand U20127 (N_20127,N_19783,N_19909);
xor U20128 (N_20128,N_19999,N_19594);
and U20129 (N_20129,N_19749,N_19508);
or U20130 (N_20130,N_19916,N_19501);
nor U20131 (N_20131,N_19899,N_19587);
xor U20132 (N_20132,N_19957,N_19907);
nor U20133 (N_20133,N_19775,N_19660);
nor U20134 (N_20134,N_19927,N_19740);
and U20135 (N_20135,N_19719,N_19592);
nor U20136 (N_20136,N_19813,N_19995);
or U20137 (N_20137,N_19782,N_19542);
and U20138 (N_20138,N_19670,N_19611);
nand U20139 (N_20139,N_19591,N_19827);
or U20140 (N_20140,N_19945,N_19753);
or U20141 (N_20141,N_19699,N_19711);
and U20142 (N_20142,N_19712,N_19917);
xor U20143 (N_20143,N_19799,N_19547);
and U20144 (N_20144,N_19615,N_19532);
or U20145 (N_20145,N_19534,N_19606);
xor U20146 (N_20146,N_19616,N_19602);
nand U20147 (N_20147,N_19669,N_19886);
nand U20148 (N_20148,N_19814,N_19797);
or U20149 (N_20149,N_19948,N_19672);
nor U20150 (N_20150,N_19733,N_19527);
xnor U20151 (N_20151,N_19709,N_19516);
xor U20152 (N_20152,N_19638,N_19538);
or U20153 (N_20153,N_19741,N_19853);
nor U20154 (N_20154,N_19743,N_19716);
nor U20155 (N_20155,N_19950,N_19811);
nor U20156 (N_20156,N_19549,N_19668);
nor U20157 (N_20157,N_19967,N_19996);
nor U20158 (N_20158,N_19637,N_19568);
and U20159 (N_20159,N_19855,N_19757);
and U20160 (N_20160,N_19867,N_19911);
xor U20161 (N_20161,N_19675,N_19644);
or U20162 (N_20162,N_19872,N_19881);
xnor U20163 (N_20163,N_19700,N_19868);
or U20164 (N_20164,N_19535,N_19651);
or U20165 (N_20165,N_19902,N_19680);
and U20166 (N_20166,N_19569,N_19746);
and U20167 (N_20167,N_19596,N_19788);
xnor U20168 (N_20168,N_19969,N_19845);
xor U20169 (N_20169,N_19856,N_19895);
nor U20170 (N_20170,N_19968,N_19780);
or U20171 (N_20171,N_19953,N_19635);
xnor U20172 (N_20172,N_19972,N_19951);
nand U20173 (N_20173,N_19688,N_19701);
and U20174 (N_20174,N_19705,N_19874);
xnor U20175 (N_20175,N_19748,N_19632);
xnor U20176 (N_20176,N_19828,N_19717);
xnor U20177 (N_20177,N_19577,N_19575);
nand U20178 (N_20178,N_19933,N_19805);
nor U20179 (N_20179,N_19572,N_19993);
and U20180 (N_20180,N_19871,N_19687);
xnor U20181 (N_20181,N_19829,N_19882);
or U20182 (N_20182,N_19839,N_19822);
nand U20183 (N_20183,N_19634,N_19901);
nand U20184 (N_20184,N_19789,N_19658);
nor U20185 (N_20185,N_19702,N_19554);
nor U20186 (N_20186,N_19597,N_19860);
nand U20187 (N_20187,N_19671,N_19509);
and U20188 (N_20188,N_19551,N_19808);
and U20189 (N_20189,N_19628,N_19513);
xnor U20190 (N_20190,N_19665,N_19593);
nand U20191 (N_20191,N_19796,N_19983);
nor U20192 (N_20192,N_19877,N_19851);
and U20193 (N_20193,N_19645,N_19823);
and U20194 (N_20194,N_19935,N_19649);
and U20195 (N_20195,N_19710,N_19964);
nand U20196 (N_20196,N_19979,N_19579);
and U20197 (N_20197,N_19677,N_19863);
xor U20198 (N_20198,N_19726,N_19998);
xnor U20199 (N_20199,N_19676,N_19618);
xnor U20200 (N_20200,N_19883,N_19982);
and U20201 (N_20201,N_19824,N_19704);
nor U20202 (N_20202,N_19652,N_19754);
nor U20203 (N_20203,N_19678,N_19781);
nand U20204 (N_20204,N_19918,N_19742);
xnor U20205 (N_20205,N_19755,N_19732);
nor U20206 (N_20206,N_19854,N_19528);
nand U20207 (N_20207,N_19689,N_19543);
or U20208 (N_20208,N_19544,N_19562);
xor U20209 (N_20209,N_19981,N_19852);
or U20210 (N_20210,N_19738,N_19724);
nor U20211 (N_20211,N_19760,N_19990);
xnor U20212 (N_20212,N_19843,N_19817);
xor U20213 (N_20213,N_19629,N_19648);
and U20214 (N_20214,N_19583,N_19713);
nand U20215 (N_20215,N_19730,N_19612);
xnor U20216 (N_20216,N_19608,N_19623);
nand U20217 (N_20217,N_19776,N_19610);
or U20218 (N_20218,N_19913,N_19869);
nand U20219 (N_20219,N_19930,N_19924);
xnor U20220 (N_20220,N_19929,N_19582);
nand U20221 (N_20221,N_19663,N_19546);
and U20222 (N_20222,N_19626,N_19681);
nor U20223 (N_20223,N_19750,N_19925);
and U20224 (N_20224,N_19825,N_19697);
or U20225 (N_20225,N_19745,N_19570);
xor U20226 (N_20226,N_19820,N_19858);
or U20227 (N_20227,N_19956,N_19906);
and U20228 (N_20228,N_19954,N_19965);
or U20229 (N_20229,N_19875,N_19673);
nand U20230 (N_20230,N_19747,N_19631);
and U20231 (N_20231,N_19800,N_19831);
and U20232 (N_20232,N_19698,N_19904);
nand U20233 (N_20233,N_19818,N_19522);
nor U20234 (N_20234,N_19880,N_19830);
or U20235 (N_20235,N_19774,N_19642);
nor U20236 (N_20236,N_19887,N_19560);
xor U20237 (N_20237,N_19625,N_19934);
xnor U20238 (N_20238,N_19836,N_19690);
nand U20239 (N_20239,N_19525,N_19714);
xor U20240 (N_20240,N_19921,N_19777);
nor U20241 (N_20241,N_19894,N_19905);
or U20242 (N_20242,N_19878,N_19692);
xnor U20243 (N_20243,N_19900,N_19873);
nor U20244 (N_20244,N_19846,N_19767);
and U20245 (N_20245,N_19944,N_19744);
nor U20246 (N_20246,N_19739,N_19997);
nor U20247 (N_20247,N_19708,N_19952);
and U20248 (N_20248,N_19833,N_19802);
xnor U20249 (N_20249,N_19762,N_19898);
nor U20250 (N_20250,N_19966,N_19787);
nand U20251 (N_20251,N_19572,N_19580);
nand U20252 (N_20252,N_19954,N_19708);
and U20253 (N_20253,N_19613,N_19657);
nor U20254 (N_20254,N_19850,N_19667);
and U20255 (N_20255,N_19825,N_19779);
nor U20256 (N_20256,N_19852,N_19751);
and U20257 (N_20257,N_19532,N_19668);
xor U20258 (N_20258,N_19701,N_19983);
nand U20259 (N_20259,N_19875,N_19612);
nand U20260 (N_20260,N_19870,N_19782);
or U20261 (N_20261,N_19593,N_19574);
xor U20262 (N_20262,N_19677,N_19712);
and U20263 (N_20263,N_19564,N_19901);
nor U20264 (N_20264,N_19663,N_19712);
nand U20265 (N_20265,N_19683,N_19821);
xnor U20266 (N_20266,N_19927,N_19973);
xnor U20267 (N_20267,N_19680,N_19987);
nand U20268 (N_20268,N_19529,N_19590);
nand U20269 (N_20269,N_19753,N_19637);
xnor U20270 (N_20270,N_19587,N_19562);
xnor U20271 (N_20271,N_19645,N_19961);
and U20272 (N_20272,N_19754,N_19849);
xnor U20273 (N_20273,N_19640,N_19533);
or U20274 (N_20274,N_19778,N_19953);
xor U20275 (N_20275,N_19985,N_19884);
nand U20276 (N_20276,N_19514,N_19796);
or U20277 (N_20277,N_19864,N_19747);
nor U20278 (N_20278,N_19849,N_19889);
xor U20279 (N_20279,N_19756,N_19873);
nor U20280 (N_20280,N_19834,N_19885);
nor U20281 (N_20281,N_19593,N_19533);
nand U20282 (N_20282,N_19502,N_19957);
xnor U20283 (N_20283,N_19781,N_19896);
and U20284 (N_20284,N_19661,N_19643);
nor U20285 (N_20285,N_19967,N_19872);
nor U20286 (N_20286,N_19959,N_19938);
and U20287 (N_20287,N_19803,N_19819);
xnor U20288 (N_20288,N_19689,N_19866);
nand U20289 (N_20289,N_19893,N_19714);
nand U20290 (N_20290,N_19857,N_19503);
nor U20291 (N_20291,N_19798,N_19512);
nor U20292 (N_20292,N_19855,N_19944);
and U20293 (N_20293,N_19823,N_19597);
nand U20294 (N_20294,N_19837,N_19917);
or U20295 (N_20295,N_19715,N_19587);
nand U20296 (N_20296,N_19828,N_19598);
xor U20297 (N_20297,N_19504,N_19689);
xor U20298 (N_20298,N_19607,N_19954);
or U20299 (N_20299,N_19657,N_19844);
xor U20300 (N_20300,N_19983,N_19850);
nand U20301 (N_20301,N_19787,N_19744);
nand U20302 (N_20302,N_19696,N_19733);
xor U20303 (N_20303,N_19736,N_19624);
nor U20304 (N_20304,N_19774,N_19974);
and U20305 (N_20305,N_19717,N_19584);
and U20306 (N_20306,N_19546,N_19739);
nand U20307 (N_20307,N_19825,N_19937);
and U20308 (N_20308,N_19641,N_19745);
and U20309 (N_20309,N_19863,N_19654);
nand U20310 (N_20310,N_19994,N_19753);
nor U20311 (N_20311,N_19688,N_19629);
xor U20312 (N_20312,N_19787,N_19751);
xor U20313 (N_20313,N_19634,N_19511);
xnor U20314 (N_20314,N_19867,N_19972);
xor U20315 (N_20315,N_19567,N_19772);
or U20316 (N_20316,N_19584,N_19821);
xnor U20317 (N_20317,N_19506,N_19927);
nand U20318 (N_20318,N_19535,N_19623);
or U20319 (N_20319,N_19758,N_19912);
nand U20320 (N_20320,N_19798,N_19976);
or U20321 (N_20321,N_19709,N_19799);
and U20322 (N_20322,N_19551,N_19753);
nand U20323 (N_20323,N_19731,N_19686);
nand U20324 (N_20324,N_19888,N_19937);
or U20325 (N_20325,N_19962,N_19646);
or U20326 (N_20326,N_19912,N_19629);
nand U20327 (N_20327,N_19596,N_19723);
nor U20328 (N_20328,N_19942,N_19668);
nand U20329 (N_20329,N_19853,N_19950);
xnor U20330 (N_20330,N_19618,N_19757);
or U20331 (N_20331,N_19952,N_19697);
or U20332 (N_20332,N_19760,N_19913);
nand U20333 (N_20333,N_19892,N_19619);
nor U20334 (N_20334,N_19633,N_19726);
xor U20335 (N_20335,N_19772,N_19858);
nand U20336 (N_20336,N_19847,N_19663);
nor U20337 (N_20337,N_19943,N_19505);
nand U20338 (N_20338,N_19860,N_19613);
nand U20339 (N_20339,N_19760,N_19610);
and U20340 (N_20340,N_19556,N_19958);
xnor U20341 (N_20341,N_19820,N_19700);
or U20342 (N_20342,N_19672,N_19647);
nor U20343 (N_20343,N_19931,N_19547);
nand U20344 (N_20344,N_19639,N_19727);
and U20345 (N_20345,N_19572,N_19883);
nor U20346 (N_20346,N_19759,N_19882);
xnor U20347 (N_20347,N_19832,N_19749);
xor U20348 (N_20348,N_19962,N_19757);
and U20349 (N_20349,N_19677,N_19761);
nand U20350 (N_20350,N_19675,N_19735);
nor U20351 (N_20351,N_19609,N_19826);
xnor U20352 (N_20352,N_19867,N_19535);
nand U20353 (N_20353,N_19866,N_19781);
and U20354 (N_20354,N_19852,N_19908);
xor U20355 (N_20355,N_19523,N_19712);
and U20356 (N_20356,N_19807,N_19961);
nand U20357 (N_20357,N_19961,N_19914);
or U20358 (N_20358,N_19997,N_19611);
nor U20359 (N_20359,N_19510,N_19624);
nand U20360 (N_20360,N_19910,N_19560);
xor U20361 (N_20361,N_19748,N_19668);
or U20362 (N_20362,N_19654,N_19763);
xor U20363 (N_20363,N_19754,N_19646);
and U20364 (N_20364,N_19604,N_19974);
and U20365 (N_20365,N_19855,N_19514);
xnor U20366 (N_20366,N_19574,N_19790);
or U20367 (N_20367,N_19884,N_19598);
and U20368 (N_20368,N_19673,N_19625);
xor U20369 (N_20369,N_19954,N_19754);
and U20370 (N_20370,N_19743,N_19631);
xnor U20371 (N_20371,N_19511,N_19789);
nand U20372 (N_20372,N_19725,N_19573);
nor U20373 (N_20373,N_19629,N_19544);
xnor U20374 (N_20374,N_19764,N_19927);
nand U20375 (N_20375,N_19916,N_19528);
nand U20376 (N_20376,N_19767,N_19762);
or U20377 (N_20377,N_19775,N_19619);
nor U20378 (N_20378,N_19792,N_19921);
and U20379 (N_20379,N_19634,N_19839);
xnor U20380 (N_20380,N_19690,N_19798);
and U20381 (N_20381,N_19681,N_19951);
and U20382 (N_20382,N_19583,N_19699);
xnor U20383 (N_20383,N_19883,N_19727);
or U20384 (N_20384,N_19903,N_19859);
or U20385 (N_20385,N_19588,N_19531);
xor U20386 (N_20386,N_19705,N_19687);
xnor U20387 (N_20387,N_19918,N_19645);
nand U20388 (N_20388,N_19596,N_19738);
nor U20389 (N_20389,N_19779,N_19877);
xnor U20390 (N_20390,N_19744,N_19581);
nor U20391 (N_20391,N_19647,N_19859);
or U20392 (N_20392,N_19503,N_19650);
xnor U20393 (N_20393,N_19918,N_19663);
and U20394 (N_20394,N_19697,N_19939);
nor U20395 (N_20395,N_19702,N_19649);
or U20396 (N_20396,N_19708,N_19943);
nor U20397 (N_20397,N_19926,N_19573);
nand U20398 (N_20398,N_19856,N_19805);
and U20399 (N_20399,N_19603,N_19562);
nor U20400 (N_20400,N_19665,N_19541);
nor U20401 (N_20401,N_19870,N_19872);
or U20402 (N_20402,N_19897,N_19888);
nor U20403 (N_20403,N_19752,N_19639);
and U20404 (N_20404,N_19535,N_19803);
or U20405 (N_20405,N_19861,N_19881);
and U20406 (N_20406,N_19715,N_19868);
and U20407 (N_20407,N_19542,N_19533);
nor U20408 (N_20408,N_19517,N_19811);
nand U20409 (N_20409,N_19638,N_19751);
nor U20410 (N_20410,N_19927,N_19614);
nand U20411 (N_20411,N_19717,N_19698);
and U20412 (N_20412,N_19986,N_19555);
xnor U20413 (N_20413,N_19824,N_19887);
or U20414 (N_20414,N_19907,N_19777);
nand U20415 (N_20415,N_19993,N_19603);
nand U20416 (N_20416,N_19967,N_19870);
nor U20417 (N_20417,N_19930,N_19925);
and U20418 (N_20418,N_19921,N_19580);
nor U20419 (N_20419,N_19572,N_19814);
or U20420 (N_20420,N_19506,N_19664);
nor U20421 (N_20421,N_19997,N_19684);
nor U20422 (N_20422,N_19551,N_19814);
and U20423 (N_20423,N_19748,N_19779);
xnor U20424 (N_20424,N_19556,N_19886);
nor U20425 (N_20425,N_19797,N_19806);
or U20426 (N_20426,N_19802,N_19962);
xor U20427 (N_20427,N_19650,N_19888);
or U20428 (N_20428,N_19884,N_19831);
or U20429 (N_20429,N_19805,N_19675);
nor U20430 (N_20430,N_19514,N_19944);
nor U20431 (N_20431,N_19970,N_19789);
nor U20432 (N_20432,N_19735,N_19509);
nor U20433 (N_20433,N_19656,N_19637);
nand U20434 (N_20434,N_19766,N_19594);
nor U20435 (N_20435,N_19574,N_19771);
or U20436 (N_20436,N_19615,N_19916);
or U20437 (N_20437,N_19809,N_19504);
or U20438 (N_20438,N_19614,N_19532);
xnor U20439 (N_20439,N_19890,N_19893);
nand U20440 (N_20440,N_19869,N_19898);
nor U20441 (N_20441,N_19797,N_19616);
nand U20442 (N_20442,N_19998,N_19507);
and U20443 (N_20443,N_19768,N_19746);
and U20444 (N_20444,N_19787,N_19819);
and U20445 (N_20445,N_19546,N_19620);
and U20446 (N_20446,N_19793,N_19895);
nand U20447 (N_20447,N_19620,N_19645);
xor U20448 (N_20448,N_19906,N_19830);
nor U20449 (N_20449,N_19837,N_19783);
and U20450 (N_20450,N_19705,N_19696);
nor U20451 (N_20451,N_19901,N_19628);
nor U20452 (N_20452,N_19719,N_19938);
nor U20453 (N_20453,N_19982,N_19718);
nand U20454 (N_20454,N_19646,N_19828);
and U20455 (N_20455,N_19811,N_19571);
xnor U20456 (N_20456,N_19860,N_19966);
xor U20457 (N_20457,N_19794,N_19909);
and U20458 (N_20458,N_19993,N_19695);
nand U20459 (N_20459,N_19758,N_19772);
nand U20460 (N_20460,N_19787,N_19871);
xor U20461 (N_20461,N_19794,N_19650);
nand U20462 (N_20462,N_19726,N_19896);
or U20463 (N_20463,N_19947,N_19738);
nand U20464 (N_20464,N_19600,N_19609);
and U20465 (N_20465,N_19837,N_19631);
nor U20466 (N_20466,N_19981,N_19727);
and U20467 (N_20467,N_19940,N_19538);
nor U20468 (N_20468,N_19587,N_19769);
or U20469 (N_20469,N_19979,N_19913);
nand U20470 (N_20470,N_19542,N_19872);
xor U20471 (N_20471,N_19853,N_19675);
and U20472 (N_20472,N_19766,N_19732);
or U20473 (N_20473,N_19572,N_19578);
or U20474 (N_20474,N_19849,N_19631);
xor U20475 (N_20475,N_19637,N_19520);
and U20476 (N_20476,N_19723,N_19550);
nand U20477 (N_20477,N_19924,N_19615);
nand U20478 (N_20478,N_19856,N_19504);
and U20479 (N_20479,N_19774,N_19648);
nor U20480 (N_20480,N_19658,N_19817);
xor U20481 (N_20481,N_19780,N_19617);
and U20482 (N_20482,N_19888,N_19614);
nor U20483 (N_20483,N_19660,N_19688);
xnor U20484 (N_20484,N_19750,N_19542);
nand U20485 (N_20485,N_19777,N_19715);
or U20486 (N_20486,N_19953,N_19692);
nand U20487 (N_20487,N_19622,N_19800);
or U20488 (N_20488,N_19688,N_19866);
or U20489 (N_20489,N_19818,N_19830);
and U20490 (N_20490,N_19985,N_19852);
or U20491 (N_20491,N_19583,N_19806);
or U20492 (N_20492,N_19856,N_19563);
and U20493 (N_20493,N_19967,N_19822);
or U20494 (N_20494,N_19724,N_19913);
or U20495 (N_20495,N_19962,N_19836);
or U20496 (N_20496,N_19942,N_19569);
nor U20497 (N_20497,N_19808,N_19674);
xor U20498 (N_20498,N_19736,N_19802);
xor U20499 (N_20499,N_19947,N_19529);
nand U20500 (N_20500,N_20302,N_20132);
xnor U20501 (N_20501,N_20474,N_20164);
nor U20502 (N_20502,N_20410,N_20133);
xor U20503 (N_20503,N_20021,N_20108);
or U20504 (N_20504,N_20285,N_20489);
nor U20505 (N_20505,N_20230,N_20432);
nand U20506 (N_20506,N_20388,N_20239);
and U20507 (N_20507,N_20014,N_20318);
and U20508 (N_20508,N_20217,N_20494);
xor U20509 (N_20509,N_20436,N_20391);
nor U20510 (N_20510,N_20402,N_20060);
or U20511 (N_20511,N_20315,N_20268);
and U20512 (N_20512,N_20360,N_20481);
nand U20513 (N_20513,N_20333,N_20303);
nor U20514 (N_20514,N_20219,N_20387);
nor U20515 (N_20515,N_20054,N_20176);
nor U20516 (N_20516,N_20479,N_20447);
xnor U20517 (N_20517,N_20063,N_20148);
xor U20518 (N_20518,N_20496,N_20144);
nor U20519 (N_20519,N_20135,N_20320);
xor U20520 (N_20520,N_20109,N_20362);
nand U20521 (N_20521,N_20450,N_20162);
xor U20522 (N_20522,N_20131,N_20119);
xor U20523 (N_20523,N_20346,N_20192);
xor U20524 (N_20524,N_20294,N_20233);
and U20525 (N_20525,N_20195,N_20273);
nand U20526 (N_20526,N_20039,N_20062);
or U20527 (N_20527,N_20311,N_20331);
or U20528 (N_20528,N_20100,N_20035);
xnor U20529 (N_20529,N_20417,N_20401);
and U20530 (N_20530,N_20161,N_20099);
nand U20531 (N_20531,N_20258,N_20016);
or U20532 (N_20532,N_20407,N_20006);
and U20533 (N_20533,N_20288,N_20202);
xor U20534 (N_20534,N_20399,N_20363);
nor U20535 (N_20535,N_20462,N_20000);
nand U20536 (N_20536,N_20348,N_20439);
or U20537 (N_20537,N_20057,N_20389);
and U20538 (N_20538,N_20174,N_20361);
nor U20539 (N_20539,N_20068,N_20046);
nand U20540 (N_20540,N_20143,N_20456);
nand U20541 (N_20541,N_20177,N_20498);
nor U20542 (N_20542,N_20246,N_20169);
nor U20543 (N_20543,N_20327,N_20368);
nand U20544 (N_20544,N_20122,N_20326);
nand U20545 (N_20545,N_20491,N_20075);
nor U20546 (N_20546,N_20266,N_20280);
nand U20547 (N_20547,N_20422,N_20191);
nor U20548 (N_20548,N_20061,N_20465);
or U20549 (N_20549,N_20194,N_20136);
nor U20550 (N_20550,N_20305,N_20340);
or U20551 (N_20551,N_20188,N_20138);
nor U20552 (N_20552,N_20356,N_20338);
nand U20553 (N_20553,N_20015,N_20008);
and U20554 (N_20554,N_20382,N_20329);
xnor U20555 (N_20555,N_20291,N_20224);
and U20556 (N_20556,N_20196,N_20409);
nor U20557 (N_20557,N_20189,N_20145);
or U20558 (N_20558,N_20421,N_20254);
or U20559 (N_20559,N_20209,N_20220);
and U20560 (N_20560,N_20396,N_20055);
or U20561 (N_20561,N_20437,N_20012);
nor U20562 (N_20562,N_20293,N_20257);
nor U20563 (N_20563,N_20250,N_20415);
nor U20564 (N_20564,N_20232,N_20124);
xnor U20565 (N_20565,N_20264,N_20026);
xor U20566 (N_20566,N_20449,N_20301);
xnor U20567 (N_20567,N_20113,N_20282);
nand U20568 (N_20568,N_20078,N_20277);
or U20569 (N_20569,N_20354,N_20065);
and U20570 (N_20570,N_20337,N_20056);
or U20571 (N_20571,N_20395,N_20272);
or U20572 (N_20572,N_20339,N_20335);
xor U20573 (N_20573,N_20098,N_20229);
xor U20574 (N_20574,N_20115,N_20438);
and U20575 (N_20575,N_20096,N_20183);
xnor U20576 (N_20576,N_20107,N_20097);
and U20577 (N_20577,N_20137,N_20134);
and U20578 (N_20578,N_20234,N_20087);
and U20579 (N_20579,N_20235,N_20070);
xnor U20580 (N_20580,N_20269,N_20466);
nand U20581 (N_20581,N_20385,N_20393);
and U20582 (N_20582,N_20166,N_20170);
nand U20583 (N_20583,N_20165,N_20412);
nand U20584 (N_20584,N_20029,N_20306);
nand U20585 (N_20585,N_20041,N_20238);
nor U20586 (N_20586,N_20158,N_20084);
xor U20587 (N_20587,N_20228,N_20022);
nor U20588 (N_20588,N_20076,N_20441);
and U20589 (N_20589,N_20429,N_20405);
and U20590 (N_20590,N_20427,N_20111);
nor U20591 (N_20591,N_20168,N_20353);
or U20592 (N_20592,N_20081,N_20398);
nor U20593 (N_20593,N_20470,N_20497);
nand U20594 (N_20594,N_20446,N_20094);
nor U20595 (N_20595,N_20178,N_20343);
xnor U20596 (N_20596,N_20430,N_20112);
nor U20597 (N_20597,N_20307,N_20355);
and U20598 (N_20598,N_20344,N_20106);
or U20599 (N_20599,N_20324,N_20197);
or U20600 (N_20600,N_20027,N_20444);
or U20601 (N_20601,N_20295,N_20198);
xnor U20602 (N_20602,N_20005,N_20478);
nor U20603 (N_20603,N_20480,N_20187);
nand U20604 (N_20604,N_20067,N_20286);
xnor U20605 (N_20605,N_20211,N_20275);
and U20606 (N_20606,N_20236,N_20036);
nand U20607 (N_20607,N_20154,N_20386);
nand U20608 (N_20608,N_20488,N_20364);
or U20609 (N_20609,N_20079,N_20180);
xnor U20610 (N_20610,N_20040,N_20179);
nor U20611 (N_20611,N_20184,N_20101);
nor U20612 (N_20612,N_20359,N_20271);
nor U20613 (N_20613,N_20117,N_20156);
and U20614 (N_20614,N_20216,N_20045);
or U20615 (N_20615,N_20038,N_20019);
and U20616 (N_20616,N_20349,N_20414);
xor U20617 (N_20617,N_20043,N_20074);
or U20618 (N_20618,N_20181,N_20457);
and U20619 (N_20619,N_20086,N_20247);
and U20620 (N_20620,N_20284,N_20123);
nor U20621 (N_20621,N_20102,N_20406);
nor U20622 (N_20622,N_20126,N_20292);
nand U20623 (N_20623,N_20423,N_20077);
nor U20624 (N_20624,N_20426,N_20376);
nand U20625 (N_20625,N_20051,N_20314);
nor U20626 (N_20626,N_20296,N_20492);
nand U20627 (N_20627,N_20153,N_20066);
and U20628 (N_20628,N_20428,N_20475);
nor U20629 (N_20629,N_20256,N_20218);
nor U20630 (N_20630,N_20118,N_20142);
nor U20631 (N_20631,N_20297,N_20241);
and U20632 (N_20632,N_20011,N_20298);
xnor U20633 (N_20633,N_20226,N_20253);
xor U20634 (N_20634,N_20050,N_20003);
nor U20635 (N_20635,N_20010,N_20009);
and U20636 (N_20636,N_20468,N_20167);
and U20637 (N_20637,N_20400,N_20274);
nor U20638 (N_20638,N_20372,N_20304);
nor U20639 (N_20639,N_20073,N_20433);
xnor U20640 (N_20640,N_20321,N_20201);
nor U20641 (N_20641,N_20317,N_20199);
or U20642 (N_20642,N_20152,N_20370);
nor U20643 (N_20643,N_20203,N_20095);
nand U20644 (N_20644,N_20049,N_20418);
and U20645 (N_20645,N_20267,N_20495);
xor U20646 (N_20646,N_20215,N_20004);
nor U20647 (N_20647,N_20416,N_20037);
nor U20648 (N_20648,N_20350,N_20411);
and U20649 (N_20649,N_20313,N_20160);
nand U20650 (N_20650,N_20259,N_20443);
xor U20651 (N_20651,N_20249,N_20044);
or U20652 (N_20652,N_20064,N_20319);
xnor U20653 (N_20653,N_20129,N_20287);
nor U20654 (N_20654,N_20227,N_20172);
or U20655 (N_20655,N_20213,N_20082);
nor U20656 (N_20656,N_20330,N_20289);
nand U20657 (N_20657,N_20461,N_20173);
and U20658 (N_20658,N_20093,N_20379);
xnor U20659 (N_20659,N_20394,N_20310);
nand U20660 (N_20660,N_20459,N_20408);
nor U20661 (N_20661,N_20323,N_20140);
and U20662 (N_20662,N_20210,N_20467);
or U20663 (N_20663,N_20089,N_20283);
nand U20664 (N_20664,N_20445,N_20033);
and U20665 (N_20665,N_20476,N_20493);
and U20666 (N_20666,N_20185,N_20141);
or U20667 (N_20667,N_20300,N_20245);
xnor U20668 (N_20668,N_20263,N_20031);
or U20669 (N_20669,N_20130,N_20251);
and U20670 (N_20670,N_20440,N_20345);
xor U20671 (N_20671,N_20223,N_20424);
or U20672 (N_20672,N_20403,N_20128);
or U20673 (N_20673,N_20384,N_20347);
or U20674 (N_20674,N_20278,N_20206);
xnor U20675 (N_20675,N_20455,N_20454);
nand U20676 (N_20676,N_20352,N_20463);
xor U20677 (N_20677,N_20052,N_20371);
or U20678 (N_20678,N_20200,N_20255);
xor U20679 (N_20679,N_20042,N_20369);
xor U20680 (N_20680,N_20451,N_20242);
and U20681 (N_20681,N_20204,N_20413);
xor U20682 (N_20682,N_20390,N_20182);
xnor U20683 (N_20683,N_20281,N_20342);
or U20684 (N_20684,N_20483,N_20002);
xnor U20685 (N_20685,N_20085,N_20435);
xnor U20686 (N_20686,N_20208,N_20090);
or U20687 (N_20687,N_20237,N_20262);
and U20688 (N_20688,N_20442,N_20155);
or U20689 (N_20689,N_20265,N_20270);
xor U20690 (N_20690,N_20469,N_20448);
and U20691 (N_20691,N_20114,N_20116);
nand U20692 (N_20692,N_20103,N_20207);
nor U20693 (N_20693,N_20023,N_20121);
xor U20694 (N_20694,N_20030,N_20299);
or U20695 (N_20695,N_20471,N_20221);
and U20696 (N_20696,N_20244,N_20452);
nand U20697 (N_20697,N_20334,N_20377);
nand U20698 (N_20698,N_20071,N_20477);
xor U20699 (N_20699,N_20147,N_20120);
xor U20700 (N_20700,N_20308,N_20425);
nand U20701 (N_20701,N_20088,N_20490);
or U20702 (N_20702,N_20186,N_20336);
or U20703 (N_20703,N_20499,N_20225);
nand U20704 (N_20704,N_20028,N_20072);
xor U20705 (N_20705,N_20316,N_20205);
xor U20706 (N_20706,N_20351,N_20397);
and U20707 (N_20707,N_20110,N_20290);
nor U20708 (N_20708,N_20240,N_20458);
xnor U20709 (N_20709,N_20034,N_20163);
or U20710 (N_20710,N_20378,N_20024);
nor U20711 (N_20711,N_20139,N_20175);
nor U20712 (N_20712,N_20366,N_20150);
or U20713 (N_20713,N_20243,N_20171);
nor U20714 (N_20714,N_20059,N_20214);
nand U20715 (N_20715,N_20001,N_20069);
xnor U20716 (N_20716,N_20260,N_20127);
or U20717 (N_20717,N_20261,N_20125);
xnor U20718 (N_20718,N_20190,N_20248);
or U20719 (N_20719,N_20309,N_20193);
or U20720 (N_20720,N_20312,N_20322);
and U20721 (N_20721,N_20212,N_20020);
and U20722 (N_20722,N_20083,N_20104);
xor U20723 (N_20723,N_20013,N_20222);
nor U20724 (N_20724,N_20404,N_20018);
or U20725 (N_20725,N_20007,N_20383);
nand U20726 (N_20726,N_20341,N_20328);
nor U20727 (N_20727,N_20105,N_20048);
nor U20728 (N_20728,N_20453,N_20357);
or U20729 (N_20729,N_20151,N_20159);
xnor U20730 (N_20730,N_20380,N_20149);
or U20731 (N_20731,N_20473,N_20092);
xnor U20732 (N_20732,N_20047,N_20080);
xnor U20733 (N_20733,N_20431,N_20486);
nor U20734 (N_20734,N_20472,N_20091);
xor U20735 (N_20735,N_20392,N_20252);
nand U20736 (N_20736,N_20146,N_20434);
or U20737 (N_20737,N_20053,N_20157);
and U20738 (N_20738,N_20325,N_20419);
and U20739 (N_20739,N_20420,N_20231);
xor U20740 (N_20740,N_20358,N_20025);
xor U20741 (N_20741,N_20485,N_20374);
xnor U20742 (N_20742,N_20365,N_20460);
xor U20743 (N_20743,N_20375,N_20464);
nor U20744 (N_20744,N_20367,N_20487);
or U20745 (N_20745,N_20373,N_20032);
nand U20746 (N_20746,N_20484,N_20332);
nand U20747 (N_20747,N_20058,N_20276);
nand U20748 (N_20748,N_20279,N_20482);
xnor U20749 (N_20749,N_20381,N_20017);
and U20750 (N_20750,N_20161,N_20246);
nor U20751 (N_20751,N_20305,N_20139);
and U20752 (N_20752,N_20159,N_20404);
and U20753 (N_20753,N_20431,N_20004);
or U20754 (N_20754,N_20140,N_20336);
or U20755 (N_20755,N_20168,N_20111);
xnor U20756 (N_20756,N_20130,N_20055);
or U20757 (N_20757,N_20241,N_20074);
xor U20758 (N_20758,N_20041,N_20151);
nor U20759 (N_20759,N_20026,N_20108);
xnor U20760 (N_20760,N_20057,N_20098);
or U20761 (N_20761,N_20366,N_20106);
xor U20762 (N_20762,N_20150,N_20220);
xor U20763 (N_20763,N_20088,N_20456);
or U20764 (N_20764,N_20347,N_20210);
nand U20765 (N_20765,N_20149,N_20345);
and U20766 (N_20766,N_20383,N_20262);
nor U20767 (N_20767,N_20461,N_20482);
xor U20768 (N_20768,N_20121,N_20193);
or U20769 (N_20769,N_20301,N_20467);
nor U20770 (N_20770,N_20482,N_20224);
or U20771 (N_20771,N_20249,N_20233);
and U20772 (N_20772,N_20045,N_20382);
and U20773 (N_20773,N_20011,N_20132);
nand U20774 (N_20774,N_20307,N_20055);
or U20775 (N_20775,N_20214,N_20493);
xnor U20776 (N_20776,N_20418,N_20048);
and U20777 (N_20777,N_20487,N_20376);
xnor U20778 (N_20778,N_20189,N_20207);
nand U20779 (N_20779,N_20322,N_20205);
xor U20780 (N_20780,N_20125,N_20113);
and U20781 (N_20781,N_20182,N_20449);
or U20782 (N_20782,N_20051,N_20177);
and U20783 (N_20783,N_20472,N_20258);
or U20784 (N_20784,N_20493,N_20010);
xnor U20785 (N_20785,N_20436,N_20022);
or U20786 (N_20786,N_20253,N_20259);
and U20787 (N_20787,N_20204,N_20116);
nand U20788 (N_20788,N_20452,N_20242);
nand U20789 (N_20789,N_20393,N_20381);
or U20790 (N_20790,N_20145,N_20456);
xor U20791 (N_20791,N_20147,N_20491);
nand U20792 (N_20792,N_20049,N_20470);
xor U20793 (N_20793,N_20051,N_20432);
or U20794 (N_20794,N_20101,N_20318);
and U20795 (N_20795,N_20464,N_20372);
nand U20796 (N_20796,N_20461,N_20395);
nand U20797 (N_20797,N_20220,N_20084);
xor U20798 (N_20798,N_20489,N_20137);
nand U20799 (N_20799,N_20114,N_20004);
or U20800 (N_20800,N_20209,N_20031);
or U20801 (N_20801,N_20369,N_20024);
nand U20802 (N_20802,N_20060,N_20478);
or U20803 (N_20803,N_20212,N_20049);
nand U20804 (N_20804,N_20021,N_20242);
nor U20805 (N_20805,N_20426,N_20308);
and U20806 (N_20806,N_20457,N_20182);
xor U20807 (N_20807,N_20313,N_20345);
or U20808 (N_20808,N_20105,N_20102);
xor U20809 (N_20809,N_20416,N_20175);
nor U20810 (N_20810,N_20468,N_20464);
nand U20811 (N_20811,N_20341,N_20131);
nor U20812 (N_20812,N_20325,N_20192);
xor U20813 (N_20813,N_20380,N_20315);
xnor U20814 (N_20814,N_20450,N_20196);
or U20815 (N_20815,N_20180,N_20418);
and U20816 (N_20816,N_20391,N_20336);
and U20817 (N_20817,N_20164,N_20317);
nor U20818 (N_20818,N_20496,N_20423);
xnor U20819 (N_20819,N_20221,N_20040);
and U20820 (N_20820,N_20431,N_20121);
xor U20821 (N_20821,N_20446,N_20313);
and U20822 (N_20822,N_20348,N_20357);
nor U20823 (N_20823,N_20313,N_20088);
nand U20824 (N_20824,N_20439,N_20486);
or U20825 (N_20825,N_20093,N_20249);
nor U20826 (N_20826,N_20253,N_20234);
nand U20827 (N_20827,N_20143,N_20065);
xnor U20828 (N_20828,N_20470,N_20226);
and U20829 (N_20829,N_20227,N_20074);
nand U20830 (N_20830,N_20270,N_20063);
or U20831 (N_20831,N_20455,N_20195);
xor U20832 (N_20832,N_20422,N_20239);
xnor U20833 (N_20833,N_20058,N_20389);
and U20834 (N_20834,N_20341,N_20308);
nor U20835 (N_20835,N_20058,N_20046);
xnor U20836 (N_20836,N_20225,N_20021);
or U20837 (N_20837,N_20281,N_20283);
nor U20838 (N_20838,N_20126,N_20488);
xnor U20839 (N_20839,N_20309,N_20000);
nand U20840 (N_20840,N_20121,N_20185);
nand U20841 (N_20841,N_20162,N_20103);
or U20842 (N_20842,N_20027,N_20016);
xnor U20843 (N_20843,N_20213,N_20266);
and U20844 (N_20844,N_20153,N_20266);
nand U20845 (N_20845,N_20382,N_20114);
or U20846 (N_20846,N_20284,N_20231);
xor U20847 (N_20847,N_20258,N_20239);
nor U20848 (N_20848,N_20175,N_20103);
and U20849 (N_20849,N_20411,N_20075);
nor U20850 (N_20850,N_20455,N_20291);
nand U20851 (N_20851,N_20279,N_20425);
nand U20852 (N_20852,N_20461,N_20265);
nand U20853 (N_20853,N_20188,N_20345);
or U20854 (N_20854,N_20494,N_20439);
nand U20855 (N_20855,N_20189,N_20362);
nor U20856 (N_20856,N_20420,N_20143);
and U20857 (N_20857,N_20198,N_20413);
and U20858 (N_20858,N_20144,N_20449);
nor U20859 (N_20859,N_20263,N_20455);
and U20860 (N_20860,N_20267,N_20145);
nor U20861 (N_20861,N_20298,N_20379);
or U20862 (N_20862,N_20384,N_20329);
nor U20863 (N_20863,N_20016,N_20263);
nor U20864 (N_20864,N_20151,N_20292);
xnor U20865 (N_20865,N_20431,N_20492);
nor U20866 (N_20866,N_20006,N_20338);
or U20867 (N_20867,N_20305,N_20470);
nor U20868 (N_20868,N_20112,N_20061);
or U20869 (N_20869,N_20001,N_20284);
and U20870 (N_20870,N_20207,N_20098);
nor U20871 (N_20871,N_20047,N_20087);
xnor U20872 (N_20872,N_20479,N_20243);
or U20873 (N_20873,N_20134,N_20232);
and U20874 (N_20874,N_20274,N_20385);
xnor U20875 (N_20875,N_20030,N_20208);
nand U20876 (N_20876,N_20025,N_20109);
and U20877 (N_20877,N_20140,N_20281);
nor U20878 (N_20878,N_20185,N_20337);
and U20879 (N_20879,N_20439,N_20286);
or U20880 (N_20880,N_20037,N_20480);
and U20881 (N_20881,N_20236,N_20078);
nor U20882 (N_20882,N_20463,N_20142);
nor U20883 (N_20883,N_20104,N_20097);
or U20884 (N_20884,N_20324,N_20317);
nor U20885 (N_20885,N_20316,N_20446);
and U20886 (N_20886,N_20065,N_20323);
nand U20887 (N_20887,N_20358,N_20194);
or U20888 (N_20888,N_20431,N_20183);
nor U20889 (N_20889,N_20270,N_20233);
and U20890 (N_20890,N_20238,N_20266);
nand U20891 (N_20891,N_20333,N_20239);
xnor U20892 (N_20892,N_20166,N_20254);
xor U20893 (N_20893,N_20032,N_20168);
and U20894 (N_20894,N_20196,N_20065);
and U20895 (N_20895,N_20125,N_20145);
xnor U20896 (N_20896,N_20137,N_20405);
or U20897 (N_20897,N_20321,N_20356);
xnor U20898 (N_20898,N_20487,N_20093);
nor U20899 (N_20899,N_20094,N_20023);
nand U20900 (N_20900,N_20402,N_20382);
nor U20901 (N_20901,N_20153,N_20123);
xnor U20902 (N_20902,N_20378,N_20350);
xnor U20903 (N_20903,N_20095,N_20077);
and U20904 (N_20904,N_20182,N_20098);
nor U20905 (N_20905,N_20046,N_20334);
and U20906 (N_20906,N_20185,N_20264);
or U20907 (N_20907,N_20032,N_20332);
or U20908 (N_20908,N_20485,N_20484);
and U20909 (N_20909,N_20423,N_20171);
or U20910 (N_20910,N_20478,N_20275);
nor U20911 (N_20911,N_20288,N_20388);
or U20912 (N_20912,N_20489,N_20445);
and U20913 (N_20913,N_20191,N_20108);
nand U20914 (N_20914,N_20236,N_20093);
nor U20915 (N_20915,N_20341,N_20076);
nor U20916 (N_20916,N_20214,N_20254);
or U20917 (N_20917,N_20151,N_20224);
xnor U20918 (N_20918,N_20192,N_20377);
xnor U20919 (N_20919,N_20499,N_20099);
and U20920 (N_20920,N_20493,N_20150);
and U20921 (N_20921,N_20397,N_20346);
nor U20922 (N_20922,N_20312,N_20464);
and U20923 (N_20923,N_20312,N_20211);
nor U20924 (N_20924,N_20026,N_20368);
xnor U20925 (N_20925,N_20295,N_20102);
nor U20926 (N_20926,N_20140,N_20419);
xor U20927 (N_20927,N_20344,N_20073);
xor U20928 (N_20928,N_20265,N_20463);
and U20929 (N_20929,N_20123,N_20043);
or U20930 (N_20930,N_20068,N_20384);
or U20931 (N_20931,N_20496,N_20414);
xor U20932 (N_20932,N_20246,N_20261);
xnor U20933 (N_20933,N_20224,N_20312);
and U20934 (N_20934,N_20233,N_20222);
and U20935 (N_20935,N_20234,N_20294);
nor U20936 (N_20936,N_20261,N_20358);
or U20937 (N_20937,N_20078,N_20406);
nor U20938 (N_20938,N_20416,N_20385);
or U20939 (N_20939,N_20202,N_20371);
nand U20940 (N_20940,N_20172,N_20032);
or U20941 (N_20941,N_20480,N_20299);
nor U20942 (N_20942,N_20389,N_20331);
xnor U20943 (N_20943,N_20200,N_20466);
and U20944 (N_20944,N_20359,N_20259);
or U20945 (N_20945,N_20045,N_20472);
nor U20946 (N_20946,N_20182,N_20283);
or U20947 (N_20947,N_20041,N_20301);
and U20948 (N_20948,N_20296,N_20078);
nor U20949 (N_20949,N_20161,N_20327);
nand U20950 (N_20950,N_20005,N_20408);
xnor U20951 (N_20951,N_20475,N_20348);
nand U20952 (N_20952,N_20467,N_20431);
nor U20953 (N_20953,N_20262,N_20197);
xnor U20954 (N_20954,N_20031,N_20452);
nand U20955 (N_20955,N_20239,N_20278);
nand U20956 (N_20956,N_20355,N_20087);
xnor U20957 (N_20957,N_20153,N_20028);
xnor U20958 (N_20958,N_20333,N_20245);
or U20959 (N_20959,N_20190,N_20435);
or U20960 (N_20960,N_20396,N_20059);
or U20961 (N_20961,N_20110,N_20482);
and U20962 (N_20962,N_20289,N_20131);
and U20963 (N_20963,N_20307,N_20492);
nand U20964 (N_20964,N_20329,N_20074);
xor U20965 (N_20965,N_20041,N_20258);
xnor U20966 (N_20966,N_20471,N_20495);
nor U20967 (N_20967,N_20371,N_20125);
xnor U20968 (N_20968,N_20115,N_20284);
xor U20969 (N_20969,N_20232,N_20288);
nor U20970 (N_20970,N_20093,N_20380);
nand U20971 (N_20971,N_20213,N_20456);
xnor U20972 (N_20972,N_20378,N_20495);
nor U20973 (N_20973,N_20143,N_20010);
and U20974 (N_20974,N_20272,N_20309);
xor U20975 (N_20975,N_20460,N_20204);
nand U20976 (N_20976,N_20004,N_20462);
xnor U20977 (N_20977,N_20325,N_20002);
nor U20978 (N_20978,N_20430,N_20250);
nand U20979 (N_20979,N_20043,N_20023);
and U20980 (N_20980,N_20125,N_20185);
nor U20981 (N_20981,N_20132,N_20376);
or U20982 (N_20982,N_20054,N_20442);
and U20983 (N_20983,N_20406,N_20456);
nand U20984 (N_20984,N_20370,N_20494);
xnor U20985 (N_20985,N_20381,N_20246);
and U20986 (N_20986,N_20273,N_20099);
xor U20987 (N_20987,N_20381,N_20050);
xnor U20988 (N_20988,N_20216,N_20083);
nor U20989 (N_20989,N_20126,N_20473);
or U20990 (N_20990,N_20343,N_20421);
nand U20991 (N_20991,N_20238,N_20090);
nor U20992 (N_20992,N_20056,N_20369);
nor U20993 (N_20993,N_20318,N_20082);
and U20994 (N_20994,N_20250,N_20378);
xnor U20995 (N_20995,N_20012,N_20157);
xnor U20996 (N_20996,N_20264,N_20365);
or U20997 (N_20997,N_20283,N_20362);
and U20998 (N_20998,N_20049,N_20425);
nor U20999 (N_20999,N_20307,N_20187);
or U21000 (N_21000,N_20865,N_20836);
nor U21001 (N_21001,N_20973,N_20977);
and U21002 (N_21002,N_20926,N_20538);
and U21003 (N_21003,N_20953,N_20637);
nand U21004 (N_21004,N_20942,N_20888);
nand U21005 (N_21005,N_20666,N_20545);
or U21006 (N_21006,N_20726,N_20842);
nor U21007 (N_21007,N_20630,N_20718);
nor U21008 (N_21008,N_20745,N_20732);
nand U21009 (N_21009,N_20959,N_20510);
or U21010 (N_21010,N_20871,N_20565);
xnor U21011 (N_21011,N_20777,N_20742);
or U21012 (N_21012,N_20567,N_20548);
nor U21013 (N_21013,N_20863,N_20859);
and U21014 (N_21014,N_20883,N_20508);
xor U21015 (N_21015,N_20828,N_20585);
xnor U21016 (N_21016,N_20833,N_20829);
or U21017 (N_21017,N_20982,N_20825);
xor U21018 (N_21018,N_20712,N_20930);
xnor U21019 (N_21019,N_20678,N_20932);
nor U21020 (N_21020,N_20940,N_20586);
nor U21021 (N_21021,N_20866,N_20700);
and U21022 (N_21022,N_20664,N_20612);
xnor U21023 (N_21023,N_20936,N_20544);
and U21024 (N_21024,N_20787,N_20920);
xnor U21025 (N_21025,N_20806,N_20980);
and U21026 (N_21026,N_20507,N_20872);
and U21027 (N_21027,N_20750,N_20788);
xor U21028 (N_21028,N_20546,N_20658);
xnor U21029 (N_21029,N_20796,N_20600);
and U21030 (N_21030,N_20961,N_20790);
xor U21031 (N_21031,N_20646,N_20801);
and U21032 (N_21032,N_20967,N_20903);
nor U21033 (N_21033,N_20992,N_20906);
or U21034 (N_21034,N_20537,N_20744);
xor U21035 (N_21035,N_20584,N_20618);
xor U21036 (N_21036,N_20627,N_20861);
xor U21037 (N_21037,N_20847,N_20519);
and U21038 (N_21038,N_20784,N_20945);
and U21039 (N_21039,N_20730,N_20955);
xnor U21040 (N_21040,N_20756,N_20993);
or U21041 (N_21041,N_20900,N_20832);
nand U21042 (N_21042,N_20530,N_20831);
or U21043 (N_21043,N_20764,N_20938);
nor U21044 (N_21044,N_20765,N_20540);
xor U21045 (N_21045,N_20799,N_20740);
or U21046 (N_21046,N_20970,N_20608);
nand U21047 (N_21047,N_20766,N_20757);
nand U21048 (N_21048,N_20746,N_20975);
xnor U21049 (N_21049,N_20710,N_20909);
nand U21050 (N_21050,N_20759,N_20918);
nand U21051 (N_21051,N_20613,N_20533);
nor U21052 (N_21052,N_20772,N_20615);
nand U21053 (N_21053,N_20556,N_20725);
xor U21054 (N_21054,N_20824,N_20962);
or U21055 (N_21055,N_20514,N_20723);
nor U21056 (N_21056,N_20914,N_20502);
or U21057 (N_21057,N_20602,N_20948);
nor U21058 (N_21058,N_20879,N_20703);
xor U21059 (N_21059,N_20793,N_20748);
and U21060 (N_21060,N_20823,N_20775);
nand U21061 (N_21061,N_20885,N_20693);
nor U21062 (N_21062,N_20997,N_20868);
and U21063 (N_21063,N_20601,N_20937);
nand U21064 (N_21064,N_20620,N_20820);
xor U21065 (N_21065,N_20672,N_20682);
xnor U21066 (N_21066,N_20968,N_20752);
or U21067 (N_21067,N_20786,N_20684);
xor U21068 (N_21068,N_20532,N_20683);
and U21069 (N_21069,N_20887,N_20628);
nor U21070 (N_21070,N_20578,N_20986);
or U21071 (N_21071,N_20529,N_20513);
xnor U21072 (N_21072,N_20943,N_20990);
nor U21073 (N_21073,N_20884,N_20898);
or U21074 (N_21074,N_20649,N_20606);
nor U21075 (N_21075,N_20535,N_20522);
xor U21076 (N_21076,N_20645,N_20941);
or U21077 (N_21077,N_20669,N_20598);
xnor U21078 (N_21078,N_20654,N_20837);
or U21079 (N_21079,N_20518,N_20735);
xnor U21080 (N_21080,N_20713,N_20983);
nor U21081 (N_21081,N_20706,N_20919);
xor U21082 (N_21082,N_20599,N_20902);
or U21083 (N_21083,N_20631,N_20794);
or U21084 (N_21084,N_20852,N_20624);
nand U21085 (N_21085,N_20721,N_20695);
nand U21086 (N_21086,N_20526,N_20517);
and U21087 (N_21087,N_20509,N_20792);
and U21088 (N_21088,N_20512,N_20560);
xor U21089 (N_21089,N_20581,N_20737);
or U21090 (N_21090,N_20877,N_20743);
xor U21091 (N_21091,N_20674,N_20729);
or U21092 (N_21092,N_20768,N_20774);
xnor U21093 (N_21093,N_20570,N_20839);
nand U21094 (N_21094,N_20952,N_20773);
nor U21095 (N_21095,N_20960,N_20855);
or U21096 (N_21096,N_20857,N_20890);
or U21097 (N_21097,N_20935,N_20853);
nor U21098 (N_21098,N_20922,N_20549);
xor U21099 (N_21099,N_20660,N_20605);
nor U21100 (N_21100,N_20886,N_20636);
nor U21101 (N_21101,N_20964,N_20619);
nand U21102 (N_21102,N_20629,N_20848);
nand U21103 (N_21103,N_20841,N_20503);
nand U21104 (N_21104,N_20617,N_20657);
and U21105 (N_21105,N_20644,N_20821);
nand U21106 (N_21106,N_20779,N_20690);
nor U21107 (N_21107,N_20681,N_20551);
and U21108 (N_21108,N_20873,N_20840);
or U21109 (N_21109,N_20838,N_20826);
nor U21110 (N_21110,N_20607,N_20651);
xor U21111 (N_21111,N_20623,N_20907);
xor U21112 (N_21112,N_20604,N_20642);
nand U21113 (N_21113,N_20711,N_20870);
nor U21114 (N_21114,N_20878,N_20500);
xnor U21115 (N_21115,N_20754,N_20845);
nand U21116 (N_21116,N_20528,N_20876);
xnor U21117 (N_21117,N_20568,N_20719);
xnor U21118 (N_21118,N_20812,N_20692);
and U21119 (N_21119,N_20609,N_20661);
nand U21120 (N_21120,N_20950,N_20553);
and U21121 (N_21121,N_20846,N_20869);
and U21122 (N_21122,N_20969,N_20778);
nor U21123 (N_21123,N_20724,N_20667);
nand U21124 (N_21124,N_20771,N_20668);
nand U21125 (N_21125,N_20554,N_20817);
or U21126 (N_21126,N_20717,N_20807);
or U21127 (N_21127,N_20734,N_20506);
nand U21128 (N_21128,N_20632,N_20834);
and U21129 (N_21129,N_20596,N_20641);
nor U21130 (N_21130,N_20856,N_20781);
and U21131 (N_21131,N_20699,N_20755);
nor U21132 (N_21132,N_20647,N_20727);
nand U21133 (N_21133,N_20648,N_20689);
nand U21134 (N_21134,N_20753,N_20827);
nor U21135 (N_21135,N_20558,N_20946);
or U21136 (N_21136,N_20951,N_20675);
nor U21137 (N_21137,N_20639,N_20763);
and U21138 (N_21138,N_20972,N_20738);
nor U21139 (N_21139,N_20927,N_20552);
nand U21140 (N_21140,N_20989,N_20761);
nand U21141 (N_21141,N_20923,N_20679);
or U21142 (N_21142,N_20731,N_20574);
nand U21143 (N_21143,N_20963,N_20999);
or U21144 (N_21144,N_20728,N_20802);
xnor U21145 (N_21145,N_20767,N_20687);
and U21146 (N_21146,N_20874,N_20944);
nor U21147 (N_21147,N_20789,N_20697);
and U21148 (N_21148,N_20653,N_20671);
or U21149 (N_21149,N_20860,N_20776);
xnor U21150 (N_21150,N_20576,N_20611);
xnor U21151 (N_21151,N_20656,N_20908);
and U21152 (N_21152,N_20715,N_20901);
nand U21153 (N_21153,N_20803,N_20722);
nand U21154 (N_21154,N_20896,N_20531);
xnor U21155 (N_21155,N_20956,N_20939);
or U21156 (N_21156,N_20593,N_20928);
or U21157 (N_21157,N_20921,N_20714);
nand U21158 (N_21158,N_20614,N_20652);
or U21159 (N_21159,N_20813,N_20539);
nand U21160 (N_21160,N_20736,N_20580);
xnor U21161 (N_21161,N_20931,N_20751);
nand U21162 (N_21162,N_20835,N_20591);
nor U21163 (N_21163,N_20979,N_20917);
xnor U21164 (N_21164,N_20588,N_20851);
or U21165 (N_21165,N_20573,N_20889);
or U21166 (N_21166,N_20701,N_20633);
and U21167 (N_21167,N_20741,N_20662);
and U21168 (N_21168,N_20676,N_20843);
nand U21169 (N_21169,N_20892,N_20696);
and U21170 (N_21170,N_20911,N_20893);
nand U21171 (N_21171,N_20563,N_20650);
nor U21172 (N_21172,N_20978,N_20910);
nor U21173 (N_21173,N_20541,N_20809);
xor U21174 (N_21174,N_20536,N_20597);
nand U21175 (N_21175,N_20610,N_20858);
xnor U21176 (N_21176,N_20670,N_20579);
and U21177 (N_21177,N_20515,N_20844);
nor U21178 (N_21178,N_20822,N_20716);
and U21179 (N_21179,N_20543,N_20557);
nor U21180 (N_21180,N_20673,N_20733);
nand U21181 (N_21181,N_20643,N_20720);
or U21182 (N_21182,N_20569,N_20704);
and U21183 (N_21183,N_20665,N_20561);
or U21184 (N_21184,N_20698,N_20805);
and U21185 (N_21185,N_20791,N_20905);
nand U21186 (N_21186,N_20795,N_20572);
xnor U21187 (N_21187,N_20957,N_20897);
or U21188 (N_21188,N_20808,N_20542);
or U21189 (N_21189,N_20622,N_20677);
and U21190 (N_21190,N_20797,N_20640);
xnor U21191 (N_21191,N_20505,N_20988);
and U21192 (N_21192,N_20815,N_20635);
and U21193 (N_21193,N_20864,N_20769);
or U21194 (N_21194,N_20929,N_20819);
nand U21195 (N_21195,N_20747,N_20810);
nand U21196 (N_21196,N_20867,N_20991);
nor U21197 (N_21197,N_20782,N_20760);
nor U21198 (N_21198,N_20739,N_20749);
nor U21199 (N_21199,N_20987,N_20984);
xnor U21200 (N_21200,N_20849,N_20616);
and U21201 (N_21201,N_20934,N_20981);
xnor U21202 (N_21202,N_20811,N_20912);
or U21203 (N_21203,N_20830,N_20996);
nor U21204 (N_21204,N_20995,N_20709);
or U21205 (N_21205,N_20916,N_20501);
xnor U21206 (N_21206,N_20949,N_20555);
nand U21207 (N_21207,N_20954,N_20958);
and U21208 (N_21208,N_20862,N_20785);
or U21209 (N_21209,N_20655,N_20881);
nor U21210 (N_21210,N_20998,N_20592);
nand U21211 (N_21211,N_20594,N_20566);
and U21212 (N_21212,N_20974,N_20895);
nor U21213 (N_21213,N_20547,N_20691);
or U21214 (N_21214,N_20504,N_20663);
or U21215 (N_21215,N_20688,N_20798);
nand U21216 (N_21216,N_20634,N_20702);
nor U21217 (N_21217,N_20523,N_20933);
and U21218 (N_21218,N_20818,N_20595);
xnor U21219 (N_21219,N_20971,N_20758);
or U21220 (N_21220,N_20659,N_20783);
nand U21221 (N_21221,N_20707,N_20525);
xor U21222 (N_21222,N_20559,N_20626);
xnor U21223 (N_21223,N_20577,N_20780);
or U21224 (N_21224,N_20854,N_20587);
and U21225 (N_21225,N_20686,N_20524);
xor U21226 (N_21226,N_20520,N_20708);
nand U21227 (N_21227,N_20534,N_20804);
or U21228 (N_21228,N_20925,N_20583);
or U21229 (N_21229,N_20965,N_20571);
nor U21230 (N_21230,N_20976,N_20564);
nand U21231 (N_21231,N_20850,N_20899);
nand U21232 (N_21232,N_20621,N_20590);
and U21233 (N_21233,N_20575,N_20516);
and U21234 (N_21234,N_20685,N_20924);
and U21235 (N_21235,N_20880,N_20891);
nor U21236 (N_21236,N_20527,N_20770);
nor U21237 (N_21237,N_20589,N_20947);
or U21238 (N_21238,N_20762,N_20875);
or U21239 (N_21239,N_20582,N_20638);
nor U21240 (N_21240,N_20966,N_20816);
or U21241 (N_21241,N_20915,N_20882);
or U21242 (N_21242,N_20913,N_20814);
nand U21243 (N_21243,N_20894,N_20603);
and U21244 (N_21244,N_20694,N_20904);
nor U21245 (N_21245,N_20800,N_20625);
and U21246 (N_21246,N_20985,N_20521);
and U21247 (N_21247,N_20511,N_20562);
nor U21248 (N_21248,N_20705,N_20994);
and U21249 (N_21249,N_20550,N_20680);
and U21250 (N_21250,N_20869,N_20690);
nor U21251 (N_21251,N_20904,N_20707);
and U21252 (N_21252,N_20885,N_20665);
xnor U21253 (N_21253,N_20668,N_20514);
xor U21254 (N_21254,N_20921,N_20910);
nand U21255 (N_21255,N_20547,N_20502);
nand U21256 (N_21256,N_20813,N_20787);
or U21257 (N_21257,N_20527,N_20588);
and U21258 (N_21258,N_20965,N_20892);
or U21259 (N_21259,N_20925,N_20869);
or U21260 (N_21260,N_20649,N_20816);
nand U21261 (N_21261,N_20527,N_20642);
nand U21262 (N_21262,N_20767,N_20664);
or U21263 (N_21263,N_20530,N_20898);
and U21264 (N_21264,N_20550,N_20788);
and U21265 (N_21265,N_20741,N_20857);
or U21266 (N_21266,N_20796,N_20643);
and U21267 (N_21267,N_20748,N_20716);
nand U21268 (N_21268,N_20601,N_20538);
xor U21269 (N_21269,N_20892,N_20611);
and U21270 (N_21270,N_20759,N_20852);
or U21271 (N_21271,N_20657,N_20816);
and U21272 (N_21272,N_20631,N_20836);
and U21273 (N_21273,N_20703,N_20808);
nor U21274 (N_21274,N_20899,N_20846);
xor U21275 (N_21275,N_20795,N_20785);
and U21276 (N_21276,N_20574,N_20518);
xor U21277 (N_21277,N_20658,N_20760);
and U21278 (N_21278,N_20952,N_20996);
or U21279 (N_21279,N_20661,N_20888);
xnor U21280 (N_21280,N_20949,N_20835);
nor U21281 (N_21281,N_20605,N_20960);
nor U21282 (N_21282,N_20834,N_20525);
and U21283 (N_21283,N_20822,N_20501);
and U21284 (N_21284,N_20673,N_20633);
xnor U21285 (N_21285,N_20724,N_20660);
and U21286 (N_21286,N_20892,N_20713);
nand U21287 (N_21287,N_20948,N_20971);
xor U21288 (N_21288,N_20826,N_20920);
and U21289 (N_21289,N_20574,N_20964);
and U21290 (N_21290,N_20873,N_20828);
nor U21291 (N_21291,N_20550,N_20921);
xor U21292 (N_21292,N_20591,N_20613);
nor U21293 (N_21293,N_20823,N_20980);
and U21294 (N_21294,N_20915,N_20783);
and U21295 (N_21295,N_20737,N_20763);
nand U21296 (N_21296,N_20636,N_20711);
and U21297 (N_21297,N_20943,N_20571);
or U21298 (N_21298,N_20917,N_20593);
nand U21299 (N_21299,N_20698,N_20777);
and U21300 (N_21300,N_20867,N_20578);
xnor U21301 (N_21301,N_20624,N_20616);
or U21302 (N_21302,N_20517,N_20556);
nor U21303 (N_21303,N_20838,N_20558);
or U21304 (N_21304,N_20616,N_20528);
and U21305 (N_21305,N_20928,N_20973);
nor U21306 (N_21306,N_20613,N_20667);
xor U21307 (N_21307,N_20633,N_20709);
nand U21308 (N_21308,N_20657,N_20574);
nand U21309 (N_21309,N_20623,N_20754);
nor U21310 (N_21310,N_20595,N_20915);
xnor U21311 (N_21311,N_20946,N_20912);
or U21312 (N_21312,N_20850,N_20648);
nand U21313 (N_21313,N_20575,N_20507);
xor U21314 (N_21314,N_20520,N_20690);
nand U21315 (N_21315,N_20539,N_20543);
nor U21316 (N_21316,N_20863,N_20885);
and U21317 (N_21317,N_20729,N_20943);
xnor U21318 (N_21318,N_20908,N_20664);
nand U21319 (N_21319,N_20534,N_20786);
nand U21320 (N_21320,N_20633,N_20878);
and U21321 (N_21321,N_20878,N_20662);
nor U21322 (N_21322,N_20567,N_20551);
nand U21323 (N_21323,N_20932,N_20808);
nand U21324 (N_21324,N_20729,N_20817);
and U21325 (N_21325,N_20869,N_20790);
xor U21326 (N_21326,N_20729,N_20824);
or U21327 (N_21327,N_20773,N_20860);
and U21328 (N_21328,N_20567,N_20793);
nor U21329 (N_21329,N_20882,N_20870);
or U21330 (N_21330,N_20805,N_20572);
nor U21331 (N_21331,N_20927,N_20722);
or U21332 (N_21332,N_20575,N_20882);
and U21333 (N_21333,N_20982,N_20678);
nand U21334 (N_21334,N_20635,N_20756);
xor U21335 (N_21335,N_20848,N_20575);
xor U21336 (N_21336,N_20689,N_20808);
nor U21337 (N_21337,N_20651,N_20678);
and U21338 (N_21338,N_20864,N_20992);
nor U21339 (N_21339,N_20505,N_20836);
nor U21340 (N_21340,N_20852,N_20848);
nand U21341 (N_21341,N_20945,N_20691);
or U21342 (N_21342,N_20763,N_20611);
xor U21343 (N_21343,N_20631,N_20867);
or U21344 (N_21344,N_20842,N_20705);
and U21345 (N_21345,N_20770,N_20971);
nand U21346 (N_21346,N_20615,N_20878);
and U21347 (N_21347,N_20671,N_20658);
xnor U21348 (N_21348,N_20812,N_20973);
xor U21349 (N_21349,N_20625,N_20834);
nand U21350 (N_21350,N_20817,N_20820);
or U21351 (N_21351,N_20933,N_20669);
or U21352 (N_21352,N_20593,N_20611);
nand U21353 (N_21353,N_20663,N_20597);
or U21354 (N_21354,N_20948,N_20911);
xnor U21355 (N_21355,N_20608,N_20633);
or U21356 (N_21356,N_20568,N_20744);
xnor U21357 (N_21357,N_20948,N_20678);
xor U21358 (N_21358,N_20859,N_20547);
and U21359 (N_21359,N_20572,N_20969);
nand U21360 (N_21360,N_20556,N_20918);
nand U21361 (N_21361,N_20850,N_20582);
or U21362 (N_21362,N_20821,N_20762);
nand U21363 (N_21363,N_20946,N_20903);
xnor U21364 (N_21364,N_20784,N_20843);
nand U21365 (N_21365,N_20985,N_20814);
and U21366 (N_21366,N_20633,N_20540);
nor U21367 (N_21367,N_20632,N_20974);
and U21368 (N_21368,N_20525,N_20637);
xor U21369 (N_21369,N_20958,N_20868);
nand U21370 (N_21370,N_20540,N_20594);
or U21371 (N_21371,N_20874,N_20684);
and U21372 (N_21372,N_20748,N_20569);
nand U21373 (N_21373,N_20953,N_20764);
and U21374 (N_21374,N_20719,N_20899);
nor U21375 (N_21375,N_20980,N_20770);
or U21376 (N_21376,N_20694,N_20733);
xor U21377 (N_21377,N_20646,N_20587);
nand U21378 (N_21378,N_20847,N_20792);
or U21379 (N_21379,N_20625,N_20541);
nor U21380 (N_21380,N_20593,N_20779);
and U21381 (N_21381,N_20743,N_20607);
nand U21382 (N_21382,N_20783,N_20943);
nor U21383 (N_21383,N_20657,N_20976);
xor U21384 (N_21384,N_20866,N_20900);
xor U21385 (N_21385,N_20973,N_20890);
or U21386 (N_21386,N_20790,N_20614);
nand U21387 (N_21387,N_20845,N_20954);
and U21388 (N_21388,N_20826,N_20669);
or U21389 (N_21389,N_20678,N_20794);
xnor U21390 (N_21390,N_20851,N_20962);
or U21391 (N_21391,N_20582,N_20879);
and U21392 (N_21392,N_20631,N_20770);
nor U21393 (N_21393,N_20998,N_20838);
nor U21394 (N_21394,N_20526,N_20798);
xor U21395 (N_21395,N_20775,N_20700);
or U21396 (N_21396,N_20941,N_20953);
or U21397 (N_21397,N_20938,N_20832);
nand U21398 (N_21398,N_20699,N_20873);
and U21399 (N_21399,N_20544,N_20864);
and U21400 (N_21400,N_20733,N_20857);
xnor U21401 (N_21401,N_20544,N_20623);
nand U21402 (N_21402,N_20875,N_20605);
or U21403 (N_21403,N_20631,N_20545);
nand U21404 (N_21404,N_20760,N_20890);
xnor U21405 (N_21405,N_20963,N_20899);
nand U21406 (N_21406,N_20648,N_20754);
nand U21407 (N_21407,N_20929,N_20705);
or U21408 (N_21408,N_20729,N_20897);
or U21409 (N_21409,N_20804,N_20975);
and U21410 (N_21410,N_20547,N_20723);
xnor U21411 (N_21411,N_20725,N_20537);
xnor U21412 (N_21412,N_20611,N_20946);
or U21413 (N_21413,N_20746,N_20732);
and U21414 (N_21414,N_20741,N_20614);
xor U21415 (N_21415,N_20527,N_20650);
xnor U21416 (N_21416,N_20727,N_20952);
xnor U21417 (N_21417,N_20920,N_20885);
nor U21418 (N_21418,N_20521,N_20572);
nand U21419 (N_21419,N_20860,N_20557);
and U21420 (N_21420,N_20599,N_20642);
xnor U21421 (N_21421,N_20771,N_20738);
and U21422 (N_21422,N_20893,N_20724);
and U21423 (N_21423,N_20539,N_20838);
or U21424 (N_21424,N_20966,N_20529);
or U21425 (N_21425,N_20812,N_20935);
and U21426 (N_21426,N_20807,N_20708);
and U21427 (N_21427,N_20758,N_20683);
xor U21428 (N_21428,N_20813,N_20807);
nand U21429 (N_21429,N_20710,N_20543);
xnor U21430 (N_21430,N_20849,N_20853);
nor U21431 (N_21431,N_20645,N_20595);
xnor U21432 (N_21432,N_20839,N_20726);
and U21433 (N_21433,N_20687,N_20879);
nor U21434 (N_21434,N_20507,N_20887);
or U21435 (N_21435,N_20959,N_20837);
or U21436 (N_21436,N_20907,N_20669);
nand U21437 (N_21437,N_20647,N_20981);
or U21438 (N_21438,N_20916,N_20514);
or U21439 (N_21439,N_20860,N_20502);
nor U21440 (N_21440,N_20828,N_20770);
xnor U21441 (N_21441,N_20656,N_20748);
nand U21442 (N_21442,N_20678,N_20795);
and U21443 (N_21443,N_20577,N_20588);
nor U21444 (N_21444,N_20574,N_20801);
nor U21445 (N_21445,N_20750,N_20957);
and U21446 (N_21446,N_20910,N_20789);
nand U21447 (N_21447,N_20592,N_20953);
and U21448 (N_21448,N_20905,N_20547);
and U21449 (N_21449,N_20833,N_20627);
and U21450 (N_21450,N_20835,N_20886);
nor U21451 (N_21451,N_20922,N_20951);
or U21452 (N_21452,N_20788,N_20723);
and U21453 (N_21453,N_20598,N_20560);
and U21454 (N_21454,N_20750,N_20581);
nand U21455 (N_21455,N_20957,N_20523);
nand U21456 (N_21456,N_20850,N_20876);
or U21457 (N_21457,N_20925,N_20845);
or U21458 (N_21458,N_20503,N_20918);
nand U21459 (N_21459,N_20500,N_20660);
nor U21460 (N_21460,N_20650,N_20707);
or U21461 (N_21461,N_20651,N_20571);
nand U21462 (N_21462,N_20945,N_20552);
xor U21463 (N_21463,N_20520,N_20760);
nand U21464 (N_21464,N_20852,N_20646);
and U21465 (N_21465,N_20813,N_20829);
nand U21466 (N_21466,N_20634,N_20751);
nor U21467 (N_21467,N_20688,N_20974);
xor U21468 (N_21468,N_20520,N_20545);
and U21469 (N_21469,N_20833,N_20898);
xor U21470 (N_21470,N_20512,N_20952);
nand U21471 (N_21471,N_20553,N_20935);
or U21472 (N_21472,N_20844,N_20826);
nor U21473 (N_21473,N_20995,N_20922);
xnor U21474 (N_21474,N_20595,N_20709);
or U21475 (N_21475,N_20662,N_20574);
xor U21476 (N_21476,N_20717,N_20887);
or U21477 (N_21477,N_20718,N_20551);
and U21478 (N_21478,N_20943,N_20603);
xor U21479 (N_21479,N_20821,N_20546);
and U21480 (N_21480,N_20611,N_20919);
and U21481 (N_21481,N_20940,N_20924);
nor U21482 (N_21482,N_20674,N_20575);
or U21483 (N_21483,N_20964,N_20626);
and U21484 (N_21484,N_20696,N_20978);
and U21485 (N_21485,N_20786,N_20607);
nand U21486 (N_21486,N_20787,N_20994);
or U21487 (N_21487,N_20917,N_20501);
nor U21488 (N_21488,N_20702,N_20503);
and U21489 (N_21489,N_20908,N_20922);
and U21490 (N_21490,N_20522,N_20764);
xnor U21491 (N_21491,N_20787,N_20770);
nor U21492 (N_21492,N_20970,N_20862);
xnor U21493 (N_21493,N_20561,N_20756);
or U21494 (N_21494,N_20894,N_20786);
nand U21495 (N_21495,N_20520,N_20670);
xnor U21496 (N_21496,N_20513,N_20638);
xor U21497 (N_21497,N_20676,N_20641);
xnor U21498 (N_21498,N_20556,N_20693);
and U21499 (N_21499,N_20789,N_20681);
nand U21500 (N_21500,N_21427,N_21276);
xor U21501 (N_21501,N_21486,N_21212);
nor U21502 (N_21502,N_21431,N_21408);
nor U21503 (N_21503,N_21102,N_21006);
nor U21504 (N_21504,N_21121,N_21363);
nand U21505 (N_21505,N_21269,N_21459);
nor U21506 (N_21506,N_21166,N_21345);
nor U21507 (N_21507,N_21359,N_21259);
nor U21508 (N_21508,N_21044,N_21379);
nor U21509 (N_21509,N_21018,N_21133);
and U21510 (N_21510,N_21029,N_21234);
and U21511 (N_21511,N_21442,N_21441);
or U21512 (N_21512,N_21423,N_21150);
nor U21513 (N_21513,N_21065,N_21344);
xnor U21514 (N_21514,N_21098,N_21145);
nand U21515 (N_21515,N_21267,N_21484);
nor U21516 (N_21516,N_21074,N_21451);
or U21517 (N_21517,N_21456,N_21156);
xnor U21518 (N_21518,N_21348,N_21125);
nand U21519 (N_21519,N_21017,N_21289);
and U21520 (N_21520,N_21055,N_21089);
and U21521 (N_21521,N_21462,N_21090);
and U21522 (N_21522,N_21415,N_21438);
or U21523 (N_21523,N_21199,N_21368);
nand U21524 (N_21524,N_21262,N_21346);
or U21525 (N_21525,N_21132,N_21097);
and U21526 (N_21526,N_21163,N_21308);
and U21527 (N_21527,N_21436,N_21034);
xor U21528 (N_21528,N_21306,N_21180);
xnor U21529 (N_21529,N_21024,N_21015);
and U21530 (N_21530,N_21053,N_21331);
or U21531 (N_21531,N_21045,N_21179);
nor U21532 (N_21532,N_21161,N_21086);
or U21533 (N_21533,N_21092,N_21112);
and U21534 (N_21534,N_21047,N_21305);
xor U21535 (N_21535,N_21338,N_21186);
nor U21536 (N_21536,N_21190,N_21217);
nor U21537 (N_21537,N_21387,N_21005);
and U21538 (N_21538,N_21321,N_21116);
and U21539 (N_21539,N_21296,N_21059);
and U21540 (N_21540,N_21214,N_21035);
nand U21541 (N_21541,N_21274,N_21482);
and U21542 (N_21542,N_21072,N_21030);
xor U21543 (N_21543,N_21286,N_21008);
or U21544 (N_21544,N_21302,N_21081);
xnor U21545 (N_21545,N_21114,N_21494);
or U21546 (N_21546,N_21106,N_21070);
nor U21547 (N_21547,N_21432,N_21463);
xnor U21548 (N_21548,N_21380,N_21157);
xnor U21549 (N_21549,N_21389,N_21160);
or U21550 (N_21550,N_21253,N_21388);
nand U21551 (N_21551,N_21196,N_21007);
nand U21552 (N_21552,N_21202,N_21236);
nand U21553 (N_21553,N_21319,N_21069);
xor U21554 (N_21554,N_21333,N_21271);
xor U21555 (N_21555,N_21407,N_21096);
nor U21556 (N_21556,N_21002,N_21499);
and U21557 (N_21557,N_21022,N_21192);
nand U21558 (N_21558,N_21085,N_21362);
nor U21559 (N_21559,N_21291,N_21210);
nand U21560 (N_21560,N_21310,N_21122);
nand U21561 (N_21561,N_21144,N_21447);
nor U21562 (N_21562,N_21245,N_21094);
nand U21563 (N_21563,N_21266,N_21315);
nand U21564 (N_21564,N_21257,N_21168);
and U21565 (N_21565,N_21252,N_21304);
xor U21566 (N_21566,N_21365,N_21128);
nor U21567 (N_21567,N_21275,N_21317);
or U21568 (N_21568,N_21285,N_21301);
nor U21569 (N_21569,N_21011,N_21298);
nand U21570 (N_21570,N_21413,N_21324);
nor U21571 (N_21571,N_21187,N_21063);
nand U21572 (N_21572,N_21421,N_21420);
and U21573 (N_21573,N_21038,N_21323);
and U21574 (N_21574,N_21472,N_21207);
nor U21575 (N_21575,N_21205,N_21327);
xor U21576 (N_21576,N_21312,N_21171);
nor U21577 (N_21577,N_21470,N_21467);
or U21578 (N_21578,N_21107,N_21231);
or U21579 (N_21579,N_21240,N_21131);
and U21580 (N_21580,N_21314,N_21465);
or U21581 (N_21581,N_21292,N_21352);
nand U21582 (N_21582,N_21215,N_21078);
nand U21583 (N_21583,N_21454,N_21490);
and U21584 (N_21584,N_21062,N_21433);
xor U21585 (N_21585,N_21258,N_21211);
xor U21586 (N_21586,N_21221,N_21256);
xnor U21587 (N_21587,N_21417,N_21109);
xnor U21588 (N_21588,N_21382,N_21347);
and U21589 (N_21589,N_21040,N_21140);
and U21590 (N_21590,N_21246,N_21049);
nand U21591 (N_21591,N_21410,N_21371);
nand U21592 (N_21592,N_21084,N_21158);
and U21593 (N_21593,N_21129,N_21228);
nand U21594 (N_21594,N_21309,N_21143);
nor U21595 (N_21595,N_21142,N_21360);
nand U21596 (N_21596,N_21381,N_21087);
nand U21597 (N_21597,N_21244,N_21077);
nor U21598 (N_21598,N_21137,N_21100);
and U21599 (N_21599,N_21169,N_21066);
xnor U21600 (N_21600,N_21043,N_21076);
xnor U21601 (N_21601,N_21393,N_21439);
nor U21602 (N_21602,N_21282,N_21225);
nor U21603 (N_21603,N_21091,N_21457);
nor U21604 (N_21604,N_21430,N_21437);
nand U21605 (N_21605,N_21127,N_21229);
nor U21606 (N_21606,N_21399,N_21342);
and U21607 (N_21607,N_21284,N_21108);
nand U21608 (N_21608,N_21406,N_21334);
or U21609 (N_21609,N_21395,N_21003);
or U21610 (N_21610,N_21268,N_21479);
nand U21611 (N_21611,N_21343,N_21119);
nor U21612 (N_21612,N_21281,N_21031);
xnor U21613 (N_21613,N_21364,N_21481);
nor U21614 (N_21614,N_21216,N_21135);
or U21615 (N_21615,N_21016,N_21004);
and U21616 (N_21616,N_21466,N_21455);
xnor U21617 (N_21617,N_21260,N_21445);
or U21618 (N_21618,N_21195,N_21299);
and U21619 (N_21619,N_21188,N_21372);
and U21620 (N_21620,N_21435,N_21358);
or U21621 (N_21621,N_21104,N_21279);
xnor U21622 (N_21622,N_21021,N_21464);
nor U21623 (N_21623,N_21079,N_21083);
and U21624 (N_21624,N_21067,N_21394);
nand U21625 (N_21625,N_21148,N_21111);
and U21626 (N_21626,N_21340,N_21329);
or U21627 (N_21627,N_21193,N_21110);
and U21628 (N_21628,N_21287,N_21283);
nand U21629 (N_21629,N_21165,N_21453);
nand U21630 (N_21630,N_21398,N_21429);
nand U21631 (N_21631,N_21009,N_21058);
or U21632 (N_21632,N_21012,N_21336);
nor U21633 (N_21633,N_21028,N_21369);
or U21634 (N_21634,N_21238,N_21496);
or U21635 (N_21635,N_21224,N_21383);
or U21636 (N_21636,N_21164,N_21474);
nand U21637 (N_21637,N_21095,N_21023);
nor U21638 (N_21638,N_21060,N_21316);
nor U21639 (N_21639,N_21130,N_21449);
and U21640 (N_21640,N_21469,N_21220);
or U21641 (N_21641,N_21219,N_21170);
and U21642 (N_21642,N_21042,N_21026);
xnor U21643 (N_21643,N_21458,N_21390);
nand U21644 (N_21644,N_21411,N_21476);
xor U21645 (N_21645,N_21303,N_21139);
nand U21646 (N_21646,N_21071,N_21014);
and U21647 (N_21647,N_21376,N_21088);
or U21648 (N_21648,N_21239,N_21332);
or U21649 (N_21649,N_21318,N_21233);
nand U21650 (N_21650,N_21374,N_21354);
xnor U21651 (N_21651,N_21434,N_21183);
and U21652 (N_21652,N_21073,N_21254);
nand U21653 (N_21653,N_21136,N_21123);
xnor U21654 (N_21654,N_21475,N_21209);
nand U21655 (N_21655,N_21293,N_21057);
nand U21656 (N_21656,N_21370,N_21033);
nor U21657 (N_21657,N_21471,N_21339);
xnor U21658 (N_21658,N_21487,N_21495);
nor U21659 (N_21659,N_21206,N_21322);
xnor U21660 (N_21660,N_21162,N_21392);
or U21661 (N_21661,N_21001,N_21311);
nand U21662 (N_21662,N_21201,N_21222);
and U21663 (N_21663,N_21175,N_21232);
xor U21664 (N_21664,N_21056,N_21356);
or U21665 (N_21665,N_21230,N_21051);
or U21666 (N_21666,N_21341,N_21046);
nand U21667 (N_21667,N_21147,N_21326);
xnor U21668 (N_21668,N_21159,N_21235);
nor U21669 (N_21669,N_21019,N_21138);
nand U21670 (N_21670,N_21172,N_21082);
and U21671 (N_21671,N_21272,N_21227);
or U21672 (N_21672,N_21270,N_21337);
nor U21673 (N_21673,N_21277,N_21025);
nor U21674 (N_21674,N_21353,N_21204);
and U21675 (N_21675,N_21404,N_21264);
nor U21676 (N_21676,N_21013,N_21386);
or U21677 (N_21677,N_21416,N_21443);
nand U21678 (N_21678,N_21054,N_21307);
nor U21679 (N_21679,N_21378,N_21151);
nor U21680 (N_21680,N_21294,N_21134);
xor U21681 (N_21681,N_21027,N_21099);
xnor U21682 (N_21682,N_21419,N_21237);
nor U21683 (N_21683,N_21010,N_21320);
nor U21684 (N_21684,N_21243,N_21313);
or U21685 (N_21685,N_21335,N_21428);
and U21686 (N_21686,N_21498,N_21497);
nand U21687 (N_21687,N_21101,N_21241);
nor U21688 (N_21688,N_21349,N_21203);
xnor U21689 (N_21689,N_21037,N_21426);
and U21690 (N_21690,N_21032,N_21414);
and U21691 (N_21691,N_21153,N_21126);
or U21692 (N_21692,N_21146,N_21351);
xnor U21693 (N_21693,N_21152,N_21249);
nand U21694 (N_21694,N_21493,N_21167);
xnor U21695 (N_21695,N_21113,N_21020);
nand U21696 (N_21696,N_21248,N_21105);
nor U21697 (N_21697,N_21048,N_21173);
nand U21698 (N_21698,N_21182,N_21491);
nor U21699 (N_21699,N_21357,N_21280);
or U21700 (N_21700,N_21141,N_21273);
and U21701 (N_21701,N_21460,N_21355);
and U21702 (N_21702,N_21242,N_21295);
xnor U21703 (N_21703,N_21485,N_21174);
or U21704 (N_21704,N_21093,N_21440);
nor U21705 (N_21705,N_21424,N_21223);
nor U21706 (N_21706,N_21461,N_21080);
nand U21707 (N_21707,N_21178,N_21297);
nor U21708 (N_21708,N_21117,N_21412);
nand U21709 (N_21709,N_21367,N_21185);
or U21710 (N_21710,N_21103,N_21120);
or U21711 (N_21711,N_21373,N_21400);
nor U21712 (N_21712,N_21492,N_21265);
and U21713 (N_21713,N_21366,N_21483);
or U21714 (N_21714,N_21052,N_21444);
xor U21715 (N_21715,N_21405,N_21488);
nand U21716 (N_21716,N_21377,N_21154);
nor U21717 (N_21717,N_21477,N_21115);
and U21718 (N_21718,N_21064,N_21480);
nand U21719 (N_21719,N_21361,N_21418);
nor U21720 (N_21720,N_21385,N_21300);
nor U21721 (N_21721,N_21036,N_21208);
or U21722 (N_21722,N_21213,N_21226);
xnor U21723 (N_21723,N_21384,N_21402);
nand U21724 (N_21724,N_21325,N_21261);
xor U21725 (N_21725,N_21290,N_21450);
and U21726 (N_21726,N_21288,N_21478);
or U21727 (N_21727,N_21448,N_21401);
nor U21728 (N_21728,N_21039,N_21191);
and U21729 (N_21729,N_21263,N_21041);
and U21730 (N_21730,N_21118,N_21255);
nand U21731 (N_21731,N_21422,N_21061);
or U21732 (N_21732,N_21247,N_21198);
and U21733 (N_21733,N_21473,N_21396);
and U21734 (N_21734,N_21200,N_21124);
nand U21735 (N_21735,N_21075,N_21425);
nand U21736 (N_21736,N_21189,N_21468);
nand U21737 (N_21737,N_21177,N_21050);
xor U21738 (N_21738,N_21184,N_21409);
nor U21739 (N_21739,N_21181,N_21251);
xnor U21740 (N_21740,N_21330,N_21391);
nor U21741 (N_21741,N_21197,N_21218);
nand U21742 (N_21742,N_21350,N_21489);
nor U21743 (N_21743,N_21403,N_21397);
xnor U21744 (N_21744,N_21194,N_21155);
and U21745 (N_21745,N_21328,N_21452);
nor U21746 (N_21746,N_21250,N_21000);
nor U21747 (N_21747,N_21278,N_21176);
nor U21748 (N_21748,N_21149,N_21446);
xor U21749 (N_21749,N_21375,N_21068);
and U21750 (N_21750,N_21234,N_21351);
and U21751 (N_21751,N_21173,N_21026);
nor U21752 (N_21752,N_21189,N_21226);
xor U21753 (N_21753,N_21441,N_21123);
nor U21754 (N_21754,N_21076,N_21187);
and U21755 (N_21755,N_21330,N_21265);
or U21756 (N_21756,N_21426,N_21113);
nor U21757 (N_21757,N_21494,N_21361);
xor U21758 (N_21758,N_21499,N_21419);
and U21759 (N_21759,N_21030,N_21457);
nor U21760 (N_21760,N_21439,N_21254);
nand U21761 (N_21761,N_21036,N_21136);
and U21762 (N_21762,N_21036,N_21436);
or U21763 (N_21763,N_21396,N_21407);
nand U21764 (N_21764,N_21376,N_21065);
nand U21765 (N_21765,N_21184,N_21010);
xnor U21766 (N_21766,N_21373,N_21162);
xor U21767 (N_21767,N_21081,N_21142);
xor U21768 (N_21768,N_21354,N_21224);
xor U21769 (N_21769,N_21370,N_21179);
nand U21770 (N_21770,N_21046,N_21294);
nor U21771 (N_21771,N_21279,N_21487);
nor U21772 (N_21772,N_21183,N_21131);
and U21773 (N_21773,N_21197,N_21371);
xnor U21774 (N_21774,N_21118,N_21105);
or U21775 (N_21775,N_21416,N_21180);
nor U21776 (N_21776,N_21473,N_21108);
nor U21777 (N_21777,N_21227,N_21105);
xnor U21778 (N_21778,N_21192,N_21062);
xnor U21779 (N_21779,N_21392,N_21444);
nor U21780 (N_21780,N_21190,N_21474);
nor U21781 (N_21781,N_21324,N_21292);
xor U21782 (N_21782,N_21458,N_21276);
nor U21783 (N_21783,N_21000,N_21358);
xnor U21784 (N_21784,N_21173,N_21205);
or U21785 (N_21785,N_21064,N_21353);
and U21786 (N_21786,N_21402,N_21221);
nand U21787 (N_21787,N_21366,N_21119);
and U21788 (N_21788,N_21154,N_21112);
and U21789 (N_21789,N_21050,N_21235);
nand U21790 (N_21790,N_21258,N_21141);
or U21791 (N_21791,N_21167,N_21217);
nor U21792 (N_21792,N_21168,N_21192);
and U21793 (N_21793,N_21486,N_21497);
nor U21794 (N_21794,N_21235,N_21348);
or U21795 (N_21795,N_21300,N_21005);
nand U21796 (N_21796,N_21168,N_21283);
and U21797 (N_21797,N_21222,N_21402);
nor U21798 (N_21798,N_21314,N_21332);
or U21799 (N_21799,N_21187,N_21466);
xor U21800 (N_21800,N_21093,N_21279);
xnor U21801 (N_21801,N_21112,N_21062);
nand U21802 (N_21802,N_21414,N_21462);
xnor U21803 (N_21803,N_21091,N_21160);
nand U21804 (N_21804,N_21499,N_21278);
and U21805 (N_21805,N_21202,N_21168);
nor U21806 (N_21806,N_21107,N_21037);
nand U21807 (N_21807,N_21239,N_21013);
nor U21808 (N_21808,N_21017,N_21034);
or U21809 (N_21809,N_21040,N_21110);
and U21810 (N_21810,N_21246,N_21358);
nand U21811 (N_21811,N_21379,N_21357);
and U21812 (N_21812,N_21077,N_21479);
xor U21813 (N_21813,N_21221,N_21206);
xnor U21814 (N_21814,N_21105,N_21318);
and U21815 (N_21815,N_21292,N_21203);
xor U21816 (N_21816,N_21281,N_21175);
and U21817 (N_21817,N_21463,N_21107);
or U21818 (N_21818,N_21328,N_21236);
nand U21819 (N_21819,N_21160,N_21182);
or U21820 (N_21820,N_21177,N_21025);
nand U21821 (N_21821,N_21096,N_21451);
or U21822 (N_21822,N_21049,N_21172);
or U21823 (N_21823,N_21336,N_21128);
or U21824 (N_21824,N_21491,N_21016);
or U21825 (N_21825,N_21255,N_21288);
nand U21826 (N_21826,N_21211,N_21162);
nand U21827 (N_21827,N_21420,N_21280);
xor U21828 (N_21828,N_21087,N_21408);
xnor U21829 (N_21829,N_21130,N_21069);
xnor U21830 (N_21830,N_21357,N_21203);
or U21831 (N_21831,N_21166,N_21453);
or U21832 (N_21832,N_21139,N_21438);
and U21833 (N_21833,N_21245,N_21255);
or U21834 (N_21834,N_21086,N_21301);
and U21835 (N_21835,N_21276,N_21069);
or U21836 (N_21836,N_21254,N_21311);
and U21837 (N_21837,N_21399,N_21483);
or U21838 (N_21838,N_21231,N_21150);
nor U21839 (N_21839,N_21321,N_21238);
and U21840 (N_21840,N_21189,N_21248);
and U21841 (N_21841,N_21050,N_21169);
nand U21842 (N_21842,N_21128,N_21072);
or U21843 (N_21843,N_21187,N_21495);
nand U21844 (N_21844,N_21322,N_21463);
xor U21845 (N_21845,N_21030,N_21173);
xnor U21846 (N_21846,N_21494,N_21475);
and U21847 (N_21847,N_21499,N_21250);
and U21848 (N_21848,N_21262,N_21223);
and U21849 (N_21849,N_21072,N_21289);
nand U21850 (N_21850,N_21069,N_21320);
xor U21851 (N_21851,N_21391,N_21338);
and U21852 (N_21852,N_21255,N_21027);
nor U21853 (N_21853,N_21434,N_21090);
xor U21854 (N_21854,N_21439,N_21169);
and U21855 (N_21855,N_21482,N_21348);
or U21856 (N_21856,N_21033,N_21389);
xnor U21857 (N_21857,N_21396,N_21431);
or U21858 (N_21858,N_21032,N_21040);
nor U21859 (N_21859,N_21073,N_21064);
xnor U21860 (N_21860,N_21002,N_21280);
or U21861 (N_21861,N_21414,N_21469);
nand U21862 (N_21862,N_21293,N_21080);
nand U21863 (N_21863,N_21041,N_21490);
and U21864 (N_21864,N_21498,N_21041);
xor U21865 (N_21865,N_21057,N_21012);
and U21866 (N_21866,N_21394,N_21102);
and U21867 (N_21867,N_21038,N_21380);
or U21868 (N_21868,N_21311,N_21138);
nand U21869 (N_21869,N_21394,N_21294);
and U21870 (N_21870,N_21274,N_21026);
and U21871 (N_21871,N_21282,N_21028);
xor U21872 (N_21872,N_21223,N_21067);
nor U21873 (N_21873,N_21474,N_21260);
and U21874 (N_21874,N_21087,N_21079);
or U21875 (N_21875,N_21193,N_21430);
nor U21876 (N_21876,N_21486,N_21341);
or U21877 (N_21877,N_21010,N_21012);
nor U21878 (N_21878,N_21029,N_21053);
nand U21879 (N_21879,N_21368,N_21484);
nor U21880 (N_21880,N_21122,N_21253);
and U21881 (N_21881,N_21451,N_21360);
or U21882 (N_21882,N_21338,N_21412);
nand U21883 (N_21883,N_21203,N_21034);
xor U21884 (N_21884,N_21439,N_21110);
nand U21885 (N_21885,N_21031,N_21214);
or U21886 (N_21886,N_21149,N_21386);
xnor U21887 (N_21887,N_21443,N_21295);
and U21888 (N_21888,N_21161,N_21476);
and U21889 (N_21889,N_21108,N_21283);
xnor U21890 (N_21890,N_21471,N_21352);
nor U21891 (N_21891,N_21399,N_21025);
and U21892 (N_21892,N_21306,N_21375);
xor U21893 (N_21893,N_21133,N_21296);
xnor U21894 (N_21894,N_21170,N_21136);
nor U21895 (N_21895,N_21260,N_21142);
xor U21896 (N_21896,N_21338,N_21189);
or U21897 (N_21897,N_21043,N_21323);
nor U21898 (N_21898,N_21395,N_21270);
and U21899 (N_21899,N_21211,N_21346);
and U21900 (N_21900,N_21441,N_21230);
nand U21901 (N_21901,N_21279,N_21271);
nand U21902 (N_21902,N_21240,N_21077);
or U21903 (N_21903,N_21265,N_21043);
xnor U21904 (N_21904,N_21435,N_21332);
or U21905 (N_21905,N_21174,N_21360);
nor U21906 (N_21906,N_21270,N_21152);
nand U21907 (N_21907,N_21108,N_21031);
or U21908 (N_21908,N_21325,N_21435);
xor U21909 (N_21909,N_21330,N_21034);
and U21910 (N_21910,N_21074,N_21131);
xor U21911 (N_21911,N_21173,N_21406);
and U21912 (N_21912,N_21153,N_21383);
xnor U21913 (N_21913,N_21201,N_21157);
and U21914 (N_21914,N_21350,N_21079);
and U21915 (N_21915,N_21107,N_21328);
or U21916 (N_21916,N_21067,N_21041);
and U21917 (N_21917,N_21382,N_21268);
nor U21918 (N_21918,N_21363,N_21253);
nand U21919 (N_21919,N_21329,N_21162);
nand U21920 (N_21920,N_21061,N_21416);
nand U21921 (N_21921,N_21421,N_21300);
xor U21922 (N_21922,N_21109,N_21303);
nor U21923 (N_21923,N_21078,N_21102);
xnor U21924 (N_21924,N_21315,N_21083);
or U21925 (N_21925,N_21466,N_21306);
nor U21926 (N_21926,N_21172,N_21080);
nand U21927 (N_21927,N_21073,N_21116);
or U21928 (N_21928,N_21335,N_21010);
and U21929 (N_21929,N_21195,N_21368);
nand U21930 (N_21930,N_21114,N_21447);
xor U21931 (N_21931,N_21405,N_21412);
xnor U21932 (N_21932,N_21205,N_21281);
or U21933 (N_21933,N_21388,N_21441);
xnor U21934 (N_21934,N_21302,N_21070);
nor U21935 (N_21935,N_21385,N_21387);
nor U21936 (N_21936,N_21319,N_21496);
and U21937 (N_21937,N_21286,N_21259);
nor U21938 (N_21938,N_21097,N_21110);
and U21939 (N_21939,N_21131,N_21471);
or U21940 (N_21940,N_21286,N_21451);
xor U21941 (N_21941,N_21188,N_21369);
and U21942 (N_21942,N_21137,N_21119);
nor U21943 (N_21943,N_21492,N_21303);
and U21944 (N_21944,N_21457,N_21323);
and U21945 (N_21945,N_21096,N_21153);
xnor U21946 (N_21946,N_21191,N_21238);
or U21947 (N_21947,N_21080,N_21236);
xnor U21948 (N_21948,N_21196,N_21189);
nor U21949 (N_21949,N_21002,N_21496);
or U21950 (N_21950,N_21175,N_21136);
and U21951 (N_21951,N_21411,N_21439);
and U21952 (N_21952,N_21482,N_21431);
or U21953 (N_21953,N_21467,N_21026);
and U21954 (N_21954,N_21249,N_21433);
nand U21955 (N_21955,N_21443,N_21174);
nor U21956 (N_21956,N_21379,N_21004);
nand U21957 (N_21957,N_21286,N_21025);
nor U21958 (N_21958,N_21277,N_21186);
nand U21959 (N_21959,N_21078,N_21158);
and U21960 (N_21960,N_21069,N_21119);
or U21961 (N_21961,N_21439,N_21170);
xnor U21962 (N_21962,N_21211,N_21135);
xor U21963 (N_21963,N_21400,N_21003);
and U21964 (N_21964,N_21376,N_21187);
nand U21965 (N_21965,N_21432,N_21024);
nand U21966 (N_21966,N_21204,N_21457);
and U21967 (N_21967,N_21090,N_21032);
nand U21968 (N_21968,N_21384,N_21076);
nor U21969 (N_21969,N_21017,N_21267);
nand U21970 (N_21970,N_21026,N_21352);
nor U21971 (N_21971,N_21277,N_21040);
or U21972 (N_21972,N_21248,N_21169);
nor U21973 (N_21973,N_21292,N_21327);
nand U21974 (N_21974,N_21361,N_21120);
and U21975 (N_21975,N_21169,N_21302);
nor U21976 (N_21976,N_21322,N_21359);
and U21977 (N_21977,N_21027,N_21167);
nor U21978 (N_21978,N_21412,N_21000);
or U21979 (N_21979,N_21318,N_21460);
nor U21980 (N_21980,N_21431,N_21038);
or U21981 (N_21981,N_21134,N_21050);
xnor U21982 (N_21982,N_21418,N_21282);
nor U21983 (N_21983,N_21365,N_21211);
nor U21984 (N_21984,N_21354,N_21155);
and U21985 (N_21985,N_21345,N_21150);
nand U21986 (N_21986,N_21108,N_21012);
and U21987 (N_21987,N_21102,N_21169);
nand U21988 (N_21988,N_21115,N_21225);
and U21989 (N_21989,N_21297,N_21226);
or U21990 (N_21990,N_21093,N_21392);
or U21991 (N_21991,N_21033,N_21138);
and U21992 (N_21992,N_21161,N_21229);
nand U21993 (N_21993,N_21275,N_21230);
or U21994 (N_21994,N_21323,N_21400);
xnor U21995 (N_21995,N_21112,N_21131);
nand U21996 (N_21996,N_21250,N_21366);
xor U21997 (N_21997,N_21019,N_21453);
nand U21998 (N_21998,N_21163,N_21250);
and U21999 (N_21999,N_21225,N_21070);
nand U22000 (N_22000,N_21963,N_21637);
or U22001 (N_22001,N_21842,N_21614);
or U22002 (N_22002,N_21778,N_21839);
or U22003 (N_22003,N_21663,N_21611);
and U22004 (N_22004,N_21796,N_21516);
nor U22005 (N_22005,N_21782,N_21832);
nand U22006 (N_22006,N_21632,N_21831);
nor U22007 (N_22007,N_21819,N_21922);
nor U22008 (N_22008,N_21514,N_21952);
nand U22009 (N_22009,N_21977,N_21931);
xor U22010 (N_22010,N_21609,N_21723);
nor U22011 (N_22011,N_21915,N_21949);
xor U22012 (N_22012,N_21884,N_21508);
nor U22013 (N_22013,N_21648,N_21826);
nand U22014 (N_22014,N_21942,N_21934);
or U22015 (N_22015,N_21652,N_21850);
nor U22016 (N_22016,N_21994,N_21789);
nor U22017 (N_22017,N_21909,N_21947);
xnor U22018 (N_22018,N_21792,N_21580);
or U22019 (N_22019,N_21904,N_21858);
xnor U22020 (N_22020,N_21622,N_21866);
nor U22021 (N_22021,N_21917,N_21607);
nor U22022 (N_22022,N_21657,N_21533);
nor U22023 (N_22023,N_21720,N_21555);
xnor U22024 (N_22024,N_21523,N_21847);
and U22025 (N_22025,N_21820,N_21989);
nor U22026 (N_22026,N_21667,N_21939);
and U22027 (N_22027,N_21608,N_21996);
and U22028 (N_22028,N_21550,N_21581);
nand U22029 (N_22029,N_21874,N_21927);
xor U22030 (N_22030,N_21623,N_21865);
xnor U22031 (N_22031,N_21510,N_21505);
xnor U22032 (N_22032,N_21702,N_21746);
or U22033 (N_22033,N_21728,N_21762);
and U22034 (N_22034,N_21861,N_21993);
nand U22035 (N_22035,N_21734,N_21871);
xor U22036 (N_22036,N_21737,N_21597);
or U22037 (N_22037,N_21846,N_21683);
nand U22038 (N_22038,N_21818,N_21857);
or U22039 (N_22039,N_21668,N_21578);
nand U22040 (N_22040,N_21670,N_21973);
or U22041 (N_22041,N_21690,N_21735);
nand U22042 (N_22042,N_21816,N_21827);
or U22043 (N_22043,N_21935,N_21719);
nand U22044 (N_22044,N_21671,N_21946);
xor U22045 (N_22045,N_21836,N_21659);
and U22046 (N_22046,N_21802,N_21674);
nand U22047 (N_22047,N_21914,N_21798);
nor U22048 (N_22048,N_21686,N_21713);
and U22049 (N_22049,N_21665,N_21599);
nor U22050 (N_22050,N_21743,N_21525);
xor U22051 (N_22051,N_21638,N_21888);
nand U22052 (N_22052,N_21862,N_21684);
nor U22053 (N_22053,N_21968,N_21695);
nand U22054 (N_22054,N_21639,N_21691);
xnor U22055 (N_22055,N_21716,N_21509);
nor U22056 (N_22056,N_21651,N_21751);
nor U22057 (N_22057,N_21618,N_21504);
xor U22058 (N_22058,N_21741,N_21901);
or U22059 (N_22059,N_21572,N_21642);
xor U22060 (N_22060,N_21726,N_21679);
nand U22061 (N_22061,N_21678,N_21520);
or U22062 (N_22062,N_21784,N_21824);
xor U22063 (N_22063,N_21813,N_21664);
and U22064 (N_22064,N_21913,N_21795);
and U22065 (N_22065,N_21945,N_21604);
and U22066 (N_22066,N_21879,N_21529);
nor U22067 (N_22067,N_21635,N_21545);
nand U22068 (N_22068,N_21907,N_21967);
and U22069 (N_22069,N_21768,N_21808);
nand U22070 (N_22070,N_21985,N_21958);
or U22071 (N_22071,N_21605,N_21929);
nand U22072 (N_22072,N_21785,N_21969);
nand U22073 (N_22073,N_21714,N_21835);
nand U22074 (N_22074,N_21972,N_21588);
nor U22075 (N_22075,N_21892,N_21752);
xor U22076 (N_22076,N_21771,N_21717);
or U22077 (N_22077,N_21528,N_21673);
or U22078 (N_22078,N_21849,N_21693);
nor U22079 (N_22079,N_21616,N_21838);
nand U22080 (N_22080,N_21910,N_21675);
nor U22081 (N_22081,N_21513,N_21692);
nand U22082 (N_22082,N_21507,N_21527);
and U22083 (N_22083,N_21805,N_21598);
and U22084 (N_22084,N_21983,N_21841);
nor U22085 (N_22085,N_21754,N_21769);
nand U22086 (N_22086,N_21562,N_21755);
xor U22087 (N_22087,N_21571,N_21577);
nor U22088 (N_22088,N_21617,N_21930);
or U22089 (N_22089,N_21556,N_21794);
or U22090 (N_22090,N_21924,N_21797);
xnor U22091 (N_22091,N_21987,N_21627);
nand U22092 (N_22092,N_21955,N_21700);
nor U22093 (N_22093,N_21512,N_21626);
nor U22094 (N_22094,N_21911,N_21902);
or U22095 (N_22095,N_21783,N_21640);
xnor U22096 (N_22096,N_21740,N_21919);
or U22097 (N_22097,N_21536,N_21685);
or U22098 (N_22098,N_21870,N_21653);
or U22099 (N_22099,N_21666,N_21926);
and U22100 (N_22100,N_21965,N_21610);
and U22101 (N_22101,N_21722,N_21697);
nand U22102 (N_22102,N_21887,N_21918);
xnor U22103 (N_22103,N_21551,N_21933);
xor U22104 (N_22104,N_21759,N_21511);
and U22105 (N_22105,N_21656,N_21753);
xnor U22106 (N_22106,N_21654,N_21767);
and U22107 (N_22107,N_21823,N_21645);
xnor U22108 (N_22108,N_21522,N_21547);
or U22109 (N_22109,N_21756,N_21982);
nor U22110 (N_22110,N_21957,N_21875);
and U22111 (N_22111,N_21567,N_21817);
or U22112 (N_22112,N_21636,N_21594);
or U22113 (N_22113,N_21701,N_21843);
nor U22114 (N_22114,N_21786,N_21574);
or U22115 (N_22115,N_21791,N_21699);
nor U22116 (N_22116,N_21526,N_21764);
xnor U22117 (N_22117,N_21540,N_21810);
nor U22118 (N_22118,N_21809,N_21583);
or U22119 (N_22119,N_21732,N_21852);
nor U22120 (N_22120,N_21559,N_21573);
and U22121 (N_22121,N_21951,N_21601);
xnor U22122 (N_22122,N_21906,N_21564);
and U22123 (N_22123,N_21706,N_21956);
nand U22124 (N_22124,N_21541,N_21979);
xnor U22125 (N_22125,N_21705,N_21585);
or U22126 (N_22126,N_21530,N_21897);
and U22127 (N_22127,N_21848,N_21660);
nor U22128 (N_22128,N_21502,N_21694);
or U22129 (N_22129,N_21672,N_21962);
nand U22130 (N_22130,N_21689,N_21576);
nor U22131 (N_22131,N_21730,N_21586);
nand U22132 (N_22132,N_21855,N_21960);
nand U22133 (N_22133,N_21736,N_21643);
xor U22134 (N_22134,N_21613,N_21634);
xnor U22135 (N_22135,N_21943,N_21553);
and U22136 (N_22136,N_21971,N_21908);
xor U22137 (N_22137,N_21709,N_21851);
or U22138 (N_22138,N_21537,N_21602);
or U22139 (N_22139,N_21758,N_21704);
nand U22140 (N_22140,N_21591,N_21825);
and U22141 (N_22141,N_21811,N_21775);
nor U22142 (N_22142,N_21621,N_21787);
and U22143 (N_22143,N_21711,N_21921);
nor U22144 (N_22144,N_21538,N_21707);
and U22145 (N_22145,N_21806,N_21696);
or U22146 (N_22146,N_21974,N_21822);
nand U22147 (N_22147,N_21928,N_21834);
and U22148 (N_22148,N_21524,N_21765);
and U22149 (N_22149,N_21669,N_21761);
nand U22150 (N_22150,N_21773,N_21940);
or U22151 (N_22151,N_21501,N_21641);
xor U22152 (N_22152,N_21568,N_21944);
and U22153 (N_22153,N_21725,N_21912);
or U22154 (N_22154,N_21676,N_21582);
or U22155 (N_22155,N_21649,N_21548);
and U22156 (N_22156,N_21544,N_21620);
xor U22157 (N_22157,N_21763,N_21860);
nor U22158 (N_22158,N_21998,N_21747);
or U22159 (N_22159,N_21631,N_21629);
or U22160 (N_22160,N_21774,N_21655);
xor U22161 (N_22161,N_21886,N_21923);
xor U22162 (N_22162,N_21590,N_21964);
nor U22163 (N_22163,N_21549,N_21814);
xor U22164 (N_22164,N_21885,N_21995);
xor U22165 (N_22165,N_21543,N_21587);
xnor U22166 (N_22166,N_21698,N_21727);
or U22167 (N_22167,N_21845,N_21615);
and U22168 (N_22168,N_21953,N_21519);
nand U22169 (N_22169,N_21646,N_21938);
and U22170 (N_22170,N_21625,N_21812);
and U22171 (N_22171,N_21745,N_21724);
nand U22172 (N_22172,N_21619,N_21954);
nand U22173 (N_22173,N_21876,N_21715);
nand U22174 (N_22174,N_21970,N_21868);
or U22175 (N_22175,N_21554,N_21677);
or U22176 (N_22176,N_21630,N_21733);
and U22177 (N_22177,N_21790,N_21920);
nor U22178 (N_22178,N_21560,N_21595);
or U22179 (N_22179,N_21566,N_21731);
nor U22180 (N_22180,N_21712,N_21729);
xor U22181 (N_22181,N_21503,N_21833);
nand U22182 (N_22182,N_21889,N_21718);
xnor U22183 (N_22183,N_21606,N_21986);
or U22184 (N_22184,N_21558,N_21772);
and U22185 (N_22185,N_21854,N_21932);
nand U22186 (N_22186,N_21807,N_21988);
nand U22187 (N_22187,N_21542,N_21760);
xnor U22188 (N_22188,N_21603,N_21781);
nor U22189 (N_22189,N_21644,N_21688);
xor U22190 (N_22190,N_21661,N_21966);
nor U22191 (N_22191,N_21779,N_21900);
nand U22192 (N_22192,N_21867,N_21890);
nand U22193 (N_22193,N_21518,N_21650);
and U22194 (N_22194,N_21600,N_21877);
and U22195 (N_22195,N_21873,N_21681);
nand U22196 (N_22196,N_21708,N_21557);
nand U22197 (N_22197,N_21905,N_21863);
nand U22198 (N_22198,N_21570,N_21575);
or U22199 (N_22199,N_21828,N_21894);
and U22200 (N_22200,N_21788,N_21853);
xor U22201 (N_22201,N_21766,N_21658);
nand U22202 (N_22202,N_21780,N_21830);
xor U22203 (N_22203,N_21898,N_21687);
xnor U22204 (N_22204,N_21565,N_21976);
nand U22205 (N_22205,N_21800,N_21978);
nand U22206 (N_22206,N_21804,N_21552);
nand U22207 (N_22207,N_21896,N_21984);
and U22208 (N_22208,N_21647,N_21959);
nand U22209 (N_22209,N_21532,N_21829);
xor U22210 (N_22210,N_21721,N_21742);
nor U22211 (N_22211,N_21992,N_21750);
nor U22212 (N_22212,N_21883,N_21776);
and U22213 (N_22213,N_21937,N_21856);
or U22214 (N_22214,N_21903,N_21997);
or U22215 (N_22215,N_21624,N_21981);
or U22216 (N_22216,N_21869,N_21878);
and U22217 (N_22217,N_21500,N_21749);
or U22218 (N_22218,N_21534,N_21569);
nor U22219 (N_22219,N_21799,N_21563);
nor U22220 (N_22220,N_21561,N_21579);
and U22221 (N_22221,N_21859,N_21837);
nand U22222 (N_22222,N_21801,N_21991);
nor U22223 (N_22223,N_21757,N_21593);
nor U22224 (N_22224,N_21770,N_21710);
or U22225 (N_22225,N_21680,N_21872);
or U22226 (N_22226,N_21531,N_21916);
or U22227 (N_22227,N_21793,N_21975);
or U22228 (N_22228,N_21891,N_21882);
nor U22229 (N_22229,N_21703,N_21682);
xor U22230 (N_22230,N_21948,N_21592);
or U22231 (N_22231,N_21589,N_21744);
nand U22232 (N_22232,N_21803,N_21739);
or U22233 (N_22233,N_21880,N_21899);
nand U22234 (N_22234,N_21515,N_21925);
or U22235 (N_22235,N_21893,N_21815);
nand U22236 (N_22236,N_21999,N_21895);
xnor U22237 (N_22237,N_21517,N_21506);
nand U22238 (N_22238,N_21612,N_21596);
or U22239 (N_22239,N_21546,N_21535);
xnor U22240 (N_22240,N_21840,N_21941);
nor U22241 (N_22241,N_21864,N_21662);
xor U22242 (N_22242,N_21777,N_21584);
nand U22243 (N_22243,N_21980,N_21539);
nand U22244 (N_22244,N_21961,N_21844);
or U22245 (N_22245,N_21748,N_21521);
and U22246 (N_22246,N_21950,N_21990);
and U22247 (N_22247,N_21821,N_21881);
nand U22248 (N_22248,N_21936,N_21738);
nand U22249 (N_22249,N_21628,N_21633);
or U22250 (N_22250,N_21826,N_21924);
nor U22251 (N_22251,N_21643,N_21612);
and U22252 (N_22252,N_21705,N_21593);
nor U22253 (N_22253,N_21550,N_21896);
or U22254 (N_22254,N_21713,N_21505);
or U22255 (N_22255,N_21735,N_21533);
nor U22256 (N_22256,N_21576,N_21638);
xor U22257 (N_22257,N_21882,N_21937);
nor U22258 (N_22258,N_21694,N_21889);
nand U22259 (N_22259,N_21680,N_21619);
nor U22260 (N_22260,N_21671,N_21965);
or U22261 (N_22261,N_21620,N_21971);
nor U22262 (N_22262,N_21855,N_21507);
xor U22263 (N_22263,N_21993,N_21723);
xor U22264 (N_22264,N_21686,N_21688);
nor U22265 (N_22265,N_21903,N_21610);
or U22266 (N_22266,N_21702,N_21866);
nand U22267 (N_22267,N_21549,N_21654);
or U22268 (N_22268,N_21954,N_21841);
or U22269 (N_22269,N_21615,N_21922);
xnor U22270 (N_22270,N_21916,N_21504);
nor U22271 (N_22271,N_21689,N_21721);
and U22272 (N_22272,N_21774,N_21917);
or U22273 (N_22273,N_21732,N_21720);
nand U22274 (N_22274,N_21730,N_21905);
and U22275 (N_22275,N_21540,N_21670);
nand U22276 (N_22276,N_21820,N_21806);
xnor U22277 (N_22277,N_21963,N_21790);
nor U22278 (N_22278,N_21898,N_21573);
or U22279 (N_22279,N_21888,N_21902);
nand U22280 (N_22280,N_21818,N_21572);
nand U22281 (N_22281,N_21707,N_21617);
nand U22282 (N_22282,N_21744,N_21934);
nor U22283 (N_22283,N_21622,N_21773);
or U22284 (N_22284,N_21796,N_21946);
nand U22285 (N_22285,N_21627,N_21762);
nand U22286 (N_22286,N_21932,N_21504);
xor U22287 (N_22287,N_21798,N_21789);
or U22288 (N_22288,N_21534,N_21653);
and U22289 (N_22289,N_21898,N_21956);
nor U22290 (N_22290,N_21624,N_21596);
nor U22291 (N_22291,N_21915,N_21859);
nor U22292 (N_22292,N_21554,N_21607);
and U22293 (N_22293,N_21863,N_21787);
nand U22294 (N_22294,N_21622,N_21903);
or U22295 (N_22295,N_21685,N_21853);
nor U22296 (N_22296,N_21528,N_21840);
or U22297 (N_22297,N_21839,N_21904);
nor U22298 (N_22298,N_21836,N_21820);
xor U22299 (N_22299,N_21869,N_21560);
or U22300 (N_22300,N_21699,N_21957);
and U22301 (N_22301,N_21856,N_21717);
nand U22302 (N_22302,N_21530,N_21640);
and U22303 (N_22303,N_21510,N_21983);
xnor U22304 (N_22304,N_21857,N_21776);
nand U22305 (N_22305,N_21801,N_21665);
nand U22306 (N_22306,N_21808,N_21556);
nor U22307 (N_22307,N_21710,N_21532);
and U22308 (N_22308,N_21697,N_21529);
nor U22309 (N_22309,N_21753,N_21818);
xnor U22310 (N_22310,N_21508,N_21845);
nand U22311 (N_22311,N_21678,N_21591);
xnor U22312 (N_22312,N_21546,N_21685);
nand U22313 (N_22313,N_21753,N_21740);
xnor U22314 (N_22314,N_21784,N_21899);
nor U22315 (N_22315,N_21682,N_21642);
xor U22316 (N_22316,N_21827,N_21634);
nor U22317 (N_22317,N_21913,N_21650);
or U22318 (N_22318,N_21969,N_21911);
nor U22319 (N_22319,N_21596,N_21830);
and U22320 (N_22320,N_21623,N_21611);
nand U22321 (N_22321,N_21775,N_21614);
xor U22322 (N_22322,N_21963,N_21852);
xor U22323 (N_22323,N_21574,N_21826);
and U22324 (N_22324,N_21525,N_21584);
nand U22325 (N_22325,N_21622,N_21700);
and U22326 (N_22326,N_21879,N_21860);
xor U22327 (N_22327,N_21947,N_21616);
nand U22328 (N_22328,N_21575,N_21801);
nor U22329 (N_22329,N_21704,N_21632);
xnor U22330 (N_22330,N_21655,N_21611);
nand U22331 (N_22331,N_21575,N_21780);
and U22332 (N_22332,N_21515,N_21637);
or U22333 (N_22333,N_21789,N_21526);
nor U22334 (N_22334,N_21631,N_21792);
xor U22335 (N_22335,N_21996,N_21835);
xnor U22336 (N_22336,N_21565,N_21728);
xnor U22337 (N_22337,N_21761,N_21744);
xor U22338 (N_22338,N_21757,N_21647);
xor U22339 (N_22339,N_21745,N_21515);
or U22340 (N_22340,N_21568,N_21772);
and U22341 (N_22341,N_21994,N_21594);
and U22342 (N_22342,N_21640,N_21789);
xor U22343 (N_22343,N_21788,N_21678);
nor U22344 (N_22344,N_21517,N_21694);
or U22345 (N_22345,N_21786,N_21972);
nand U22346 (N_22346,N_21925,N_21531);
or U22347 (N_22347,N_21905,N_21768);
and U22348 (N_22348,N_21804,N_21734);
xnor U22349 (N_22349,N_21682,N_21699);
and U22350 (N_22350,N_21585,N_21897);
or U22351 (N_22351,N_21934,N_21631);
xnor U22352 (N_22352,N_21811,N_21701);
nor U22353 (N_22353,N_21623,N_21613);
xnor U22354 (N_22354,N_21928,N_21860);
nor U22355 (N_22355,N_21607,N_21652);
nand U22356 (N_22356,N_21609,N_21502);
xor U22357 (N_22357,N_21708,N_21738);
xor U22358 (N_22358,N_21741,N_21815);
nand U22359 (N_22359,N_21617,N_21546);
and U22360 (N_22360,N_21619,N_21663);
and U22361 (N_22361,N_21649,N_21570);
xnor U22362 (N_22362,N_21893,N_21651);
xnor U22363 (N_22363,N_21532,N_21716);
nor U22364 (N_22364,N_21989,N_21941);
nor U22365 (N_22365,N_21544,N_21929);
and U22366 (N_22366,N_21712,N_21718);
nor U22367 (N_22367,N_21756,N_21661);
nor U22368 (N_22368,N_21813,N_21775);
xor U22369 (N_22369,N_21989,N_21630);
nor U22370 (N_22370,N_21585,N_21778);
nand U22371 (N_22371,N_21802,N_21730);
and U22372 (N_22372,N_21510,N_21875);
xnor U22373 (N_22373,N_21722,N_21881);
xnor U22374 (N_22374,N_21872,N_21724);
or U22375 (N_22375,N_21655,N_21622);
or U22376 (N_22376,N_21556,N_21821);
nor U22377 (N_22377,N_21544,N_21961);
xnor U22378 (N_22378,N_21906,N_21965);
and U22379 (N_22379,N_21646,N_21837);
nor U22380 (N_22380,N_21793,N_21799);
and U22381 (N_22381,N_21987,N_21935);
nand U22382 (N_22382,N_21933,N_21659);
nor U22383 (N_22383,N_21869,N_21804);
and U22384 (N_22384,N_21769,N_21674);
nand U22385 (N_22385,N_21769,N_21743);
or U22386 (N_22386,N_21691,N_21676);
or U22387 (N_22387,N_21853,N_21556);
or U22388 (N_22388,N_21803,N_21919);
xor U22389 (N_22389,N_21941,N_21551);
nand U22390 (N_22390,N_21846,N_21554);
or U22391 (N_22391,N_21959,N_21716);
nor U22392 (N_22392,N_21869,N_21523);
and U22393 (N_22393,N_21684,N_21544);
and U22394 (N_22394,N_21960,N_21844);
or U22395 (N_22395,N_21783,N_21534);
and U22396 (N_22396,N_21573,N_21990);
and U22397 (N_22397,N_21823,N_21888);
nand U22398 (N_22398,N_21614,N_21547);
xor U22399 (N_22399,N_21778,N_21526);
nor U22400 (N_22400,N_21591,N_21894);
nor U22401 (N_22401,N_21789,N_21542);
nand U22402 (N_22402,N_21757,N_21956);
and U22403 (N_22403,N_21656,N_21523);
and U22404 (N_22404,N_21941,N_21971);
and U22405 (N_22405,N_21902,N_21500);
xnor U22406 (N_22406,N_21652,N_21548);
or U22407 (N_22407,N_21566,N_21668);
and U22408 (N_22408,N_21563,N_21642);
nor U22409 (N_22409,N_21950,N_21608);
or U22410 (N_22410,N_21540,N_21552);
xor U22411 (N_22411,N_21657,N_21772);
nor U22412 (N_22412,N_21787,N_21724);
or U22413 (N_22413,N_21555,N_21871);
nor U22414 (N_22414,N_21887,N_21536);
nor U22415 (N_22415,N_21960,N_21604);
and U22416 (N_22416,N_21891,N_21687);
xnor U22417 (N_22417,N_21577,N_21966);
and U22418 (N_22418,N_21800,N_21821);
or U22419 (N_22419,N_21657,N_21761);
xor U22420 (N_22420,N_21861,N_21673);
xnor U22421 (N_22421,N_21932,N_21714);
or U22422 (N_22422,N_21961,N_21527);
or U22423 (N_22423,N_21828,N_21981);
xor U22424 (N_22424,N_21672,N_21580);
nor U22425 (N_22425,N_21721,N_21703);
or U22426 (N_22426,N_21973,N_21843);
and U22427 (N_22427,N_21839,N_21876);
or U22428 (N_22428,N_21555,N_21686);
nand U22429 (N_22429,N_21743,N_21716);
xnor U22430 (N_22430,N_21671,N_21820);
nand U22431 (N_22431,N_21679,N_21759);
nor U22432 (N_22432,N_21643,N_21526);
or U22433 (N_22433,N_21546,N_21792);
nor U22434 (N_22434,N_21925,N_21852);
nand U22435 (N_22435,N_21705,N_21902);
nand U22436 (N_22436,N_21552,N_21926);
nor U22437 (N_22437,N_21858,N_21814);
xor U22438 (N_22438,N_21971,N_21636);
xor U22439 (N_22439,N_21782,N_21887);
or U22440 (N_22440,N_21655,N_21554);
or U22441 (N_22441,N_21914,N_21764);
nor U22442 (N_22442,N_21545,N_21783);
and U22443 (N_22443,N_21879,N_21825);
nor U22444 (N_22444,N_21521,N_21876);
nand U22445 (N_22445,N_21935,N_21970);
or U22446 (N_22446,N_21942,N_21677);
xnor U22447 (N_22447,N_21641,N_21803);
and U22448 (N_22448,N_21908,N_21590);
or U22449 (N_22449,N_21793,N_21672);
xor U22450 (N_22450,N_21680,N_21991);
or U22451 (N_22451,N_21842,N_21881);
xor U22452 (N_22452,N_21875,N_21534);
nor U22453 (N_22453,N_21566,N_21697);
nor U22454 (N_22454,N_21847,N_21996);
xnor U22455 (N_22455,N_21668,N_21839);
nand U22456 (N_22456,N_21916,N_21533);
nand U22457 (N_22457,N_21742,N_21593);
or U22458 (N_22458,N_21628,N_21595);
xor U22459 (N_22459,N_21923,N_21587);
xnor U22460 (N_22460,N_21595,N_21991);
nand U22461 (N_22461,N_21942,N_21602);
xor U22462 (N_22462,N_21842,N_21910);
and U22463 (N_22463,N_21558,N_21999);
and U22464 (N_22464,N_21625,N_21504);
nand U22465 (N_22465,N_21624,N_21829);
nor U22466 (N_22466,N_21646,N_21666);
nand U22467 (N_22467,N_21866,N_21973);
and U22468 (N_22468,N_21976,N_21650);
xnor U22469 (N_22469,N_21887,N_21706);
nor U22470 (N_22470,N_21885,N_21597);
nor U22471 (N_22471,N_21696,N_21839);
nand U22472 (N_22472,N_21592,N_21809);
nor U22473 (N_22473,N_21749,N_21541);
nand U22474 (N_22474,N_21528,N_21677);
nor U22475 (N_22475,N_21877,N_21886);
xnor U22476 (N_22476,N_21760,N_21560);
xnor U22477 (N_22477,N_21956,N_21593);
and U22478 (N_22478,N_21715,N_21735);
and U22479 (N_22479,N_21604,N_21704);
nand U22480 (N_22480,N_21570,N_21665);
or U22481 (N_22481,N_21742,N_21887);
and U22482 (N_22482,N_21609,N_21689);
nand U22483 (N_22483,N_21697,N_21875);
xor U22484 (N_22484,N_21879,N_21867);
nand U22485 (N_22485,N_21810,N_21913);
nor U22486 (N_22486,N_21625,N_21867);
and U22487 (N_22487,N_21907,N_21761);
xnor U22488 (N_22488,N_21959,N_21834);
and U22489 (N_22489,N_21532,N_21780);
and U22490 (N_22490,N_21628,N_21812);
nor U22491 (N_22491,N_21884,N_21778);
xor U22492 (N_22492,N_21530,N_21844);
nor U22493 (N_22493,N_21693,N_21893);
nor U22494 (N_22494,N_21604,N_21539);
or U22495 (N_22495,N_21780,N_21601);
nand U22496 (N_22496,N_21932,N_21973);
or U22497 (N_22497,N_21967,N_21758);
xnor U22498 (N_22498,N_21730,N_21696);
and U22499 (N_22499,N_21742,N_21863);
or U22500 (N_22500,N_22443,N_22334);
nor U22501 (N_22501,N_22196,N_22450);
or U22502 (N_22502,N_22139,N_22438);
nand U22503 (N_22503,N_22027,N_22363);
nand U22504 (N_22504,N_22041,N_22067);
nand U22505 (N_22505,N_22049,N_22128);
and U22506 (N_22506,N_22216,N_22491);
and U22507 (N_22507,N_22335,N_22458);
or U22508 (N_22508,N_22129,N_22276);
xnor U22509 (N_22509,N_22286,N_22215);
or U22510 (N_22510,N_22386,N_22315);
xnor U22511 (N_22511,N_22384,N_22451);
xor U22512 (N_22512,N_22261,N_22298);
nand U22513 (N_22513,N_22475,N_22273);
or U22514 (N_22514,N_22252,N_22373);
nor U22515 (N_22515,N_22417,N_22225);
nand U22516 (N_22516,N_22006,N_22357);
nand U22517 (N_22517,N_22400,N_22448);
nand U22518 (N_22518,N_22299,N_22415);
nand U22519 (N_22519,N_22105,N_22060);
nand U22520 (N_22520,N_22176,N_22122);
or U22521 (N_22521,N_22178,N_22078);
and U22522 (N_22522,N_22388,N_22038);
nor U22523 (N_22523,N_22396,N_22358);
nand U22524 (N_22524,N_22277,N_22249);
xnor U22525 (N_22525,N_22248,N_22020);
and U22526 (N_22526,N_22354,N_22211);
xor U22527 (N_22527,N_22452,N_22399);
or U22528 (N_22528,N_22093,N_22408);
or U22529 (N_22529,N_22200,N_22203);
and U22530 (N_22530,N_22403,N_22307);
nand U22531 (N_22531,N_22207,N_22444);
and U22532 (N_22532,N_22285,N_22103);
nor U22533 (N_22533,N_22181,N_22247);
xnor U22534 (N_22534,N_22425,N_22441);
nand U22535 (N_22535,N_22472,N_22222);
and U22536 (N_22536,N_22208,N_22017);
and U22537 (N_22537,N_22025,N_22231);
nand U22538 (N_22538,N_22187,N_22494);
xor U22539 (N_22539,N_22063,N_22083);
nor U22540 (N_22540,N_22087,N_22137);
nor U22541 (N_22541,N_22412,N_22381);
and U22542 (N_22542,N_22165,N_22221);
nor U22543 (N_22543,N_22056,N_22242);
nor U22544 (N_22544,N_22317,N_22353);
nand U22545 (N_22545,N_22086,N_22439);
or U22546 (N_22546,N_22497,N_22360);
nor U22547 (N_22547,N_22449,N_22162);
or U22548 (N_22548,N_22202,N_22119);
or U22549 (N_22549,N_22191,N_22468);
or U22550 (N_22550,N_22008,N_22486);
or U22551 (N_22551,N_22218,N_22346);
nand U22552 (N_22552,N_22467,N_22471);
xor U22553 (N_22553,N_22167,N_22465);
nor U22554 (N_22554,N_22433,N_22032);
nor U22555 (N_22555,N_22136,N_22376);
nor U22556 (N_22556,N_22320,N_22104);
or U22557 (N_22557,N_22096,N_22095);
xnor U22558 (N_22558,N_22295,N_22476);
nand U22559 (N_22559,N_22340,N_22350);
and U22560 (N_22560,N_22427,N_22309);
or U22561 (N_22561,N_22151,N_22253);
or U22562 (N_22562,N_22397,N_22291);
nor U22563 (N_22563,N_22237,N_22062);
or U22564 (N_22564,N_22485,N_22199);
or U22565 (N_22565,N_22344,N_22143);
nor U22566 (N_22566,N_22304,N_22430);
nor U22567 (N_22567,N_22023,N_22488);
or U22568 (N_22568,N_22455,N_22132);
xor U22569 (N_22569,N_22287,N_22058);
and U22570 (N_22570,N_22398,N_22311);
nor U22571 (N_22571,N_22493,N_22442);
and U22572 (N_22572,N_22016,N_22289);
xor U22573 (N_22573,N_22153,N_22057);
and U22574 (N_22574,N_22303,N_22026);
and U22575 (N_22575,N_22102,N_22134);
nand U22576 (N_22576,N_22391,N_22414);
and U22577 (N_22577,N_22004,N_22257);
nor U22578 (N_22578,N_22238,N_22292);
xor U22579 (N_22579,N_22477,N_22126);
and U22580 (N_22580,N_22009,N_22039);
nor U22581 (N_22581,N_22219,N_22305);
nand U22582 (N_22582,N_22308,N_22213);
or U22583 (N_22583,N_22243,N_22319);
nand U22584 (N_22584,N_22115,N_22157);
or U22585 (N_22585,N_22375,N_22236);
nand U22586 (N_22586,N_22380,N_22499);
or U22587 (N_22587,N_22082,N_22091);
nor U22588 (N_22588,N_22436,N_22330);
xor U22589 (N_22589,N_22015,N_22445);
or U22590 (N_22590,N_22053,N_22235);
or U22591 (N_22591,N_22367,N_22045);
xnor U22592 (N_22592,N_22158,N_22481);
nor U22593 (N_22593,N_22492,N_22431);
nand U22594 (N_22594,N_22434,N_22270);
or U22595 (N_22595,N_22055,N_22068);
and U22596 (N_22596,N_22021,N_22379);
and U22597 (N_22597,N_22409,N_22478);
nand U22598 (N_22598,N_22395,N_22401);
and U22599 (N_22599,N_22495,N_22003);
nand U22600 (N_22600,N_22031,N_22271);
nand U22601 (N_22601,N_22234,N_22141);
or U22602 (N_22602,N_22229,N_22254);
xnor U22603 (N_22603,N_22002,N_22099);
xnor U22604 (N_22604,N_22177,N_22239);
nor U22605 (N_22605,N_22364,N_22327);
nor U22606 (N_22606,N_22185,N_22352);
or U22607 (N_22607,N_22255,N_22097);
nor U22608 (N_22608,N_22496,N_22163);
nor U22609 (N_22609,N_22269,N_22101);
nand U22610 (N_22610,N_22005,N_22259);
nor U22611 (N_22611,N_22462,N_22265);
and U22612 (N_22612,N_22047,N_22461);
xor U22613 (N_22613,N_22166,N_22175);
xor U22614 (N_22614,N_22404,N_22012);
nor U22615 (N_22615,N_22470,N_22085);
nor U22616 (N_22616,N_22189,N_22090);
and U22617 (N_22617,N_22283,N_22326);
xor U22618 (N_22618,N_22356,N_22226);
nand U22619 (N_22619,N_22392,N_22416);
and U22620 (N_22620,N_22161,N_22256);
and U22621 (N_22621,N_22378,N_22370);
xnor U22622 (N_22622,N_22170,N_22127);
nand U22623 (N_22623,N_22028,N_22297);
nand U22624 (N_22624,N_22150,N_22424);
xnor U22625 (N_22625,N_22421,N_22098);
or U22626 (N_22626,N_22114,N_22355);
nor U22627 (N_22627,N_22044,N_22263);
or U22628 (N_22628,N_22473,N_22149);
or U22629 (N_22629,N_22490,N_22147);
xor U22630 (N_22630,N_22301,N_22343);
nor U22631 (N_22631,N_22197,N_22065);
and U22632 (N_22632,N_22437,N_22489);
xor U22633 (N_22633,N_22368,N_22071);
xor U22634 (N_22634,N_22423,N_22156);
nor U22635 (N_22635,N_22075,N_22076);
and U22636 (N_22636,N_22447,N_22107);
or U22637 (N_22637,N_22389,N_22281);
and U22638 (N_22638,N_22074,N_22453);
or U22639 (N_22639,N_22328,N_22073);
nor U22640 (N_22640,N_22100,N_22474);
and U22641 (N_22641,N_22325,N_22125);
and U22642 (N_22642,N_22106,N_22140);
and U22643 (N_22643,N_22131,N_22174);
or U22644 (N_22644,N_22419,N_22413);
nand U22645 (N_22645,N_22172,N_22007);
nand U22646 (N_22646,N_22022,N_22275);
nor U22647 (N_22647,N_22169,N_22069);
and U22648 (N_22648,N_22418,N_22011);
or U22649 (N_22649,N_22498,N_22332);
xnor U22650 (N_22650,N_22300,N_22124);
nor U22651 (N_22651,N_22195,N_22064);
and U22652 (N_22652,N_22179,N_22456);
xor U22653 (N_22653,N_22422,N_22435);
nor U22654 (N_22654,N_22382,N_22460);
nand U22655 (N_22655,N_22037,N_22402);
and U22656 (N_22656,N_22324,N_22142);
and U22657 (N_22657,N_22469,N_22390);
or U22658 (N_22658,N_22089,N_22043);
or U22659 (N_22659,N_22018,N_22144);
and U22660 (N_22660,N_22410,N_22168);
or U22661 (N_22661,N_22333,N_22341);
nor U22662 (N_22662,N_22224,N_22278);
nor U22663 (N_22663,N_22204,N_22145);
or U22664 (N_22664,N_22429,N_22371);
or U22665 (N_22665,N_22072,N_22088);
xnor U22666 (N_22666,N_22080,N_22446);
or U22667 (N_22667,N_22267,N_22426);
nor U22668 (N_22668,N_22116,N_22407);
or U22669 (N_22669,N_22383,N_22362);
and U22670 (N_22670,N_22194,N_22316);
or U22671 (N_22671,N_22323,N_22306);
and U22672 (N_22672,N_22280,N_22349);
or U22673 (N_22673,N_22464,N_22123);
xnor U22674 (N_22674,N_22066,N_22318);
nand U22675 (N_22675,N_22251,N_22040);
and U22676 (N_22676,N_22394,N_22454);
and U22677 (N_22677,N_22138,N_22113);
or U22678 (N_22678,N_22024,N_22385);
or U22679 (N_22679,N_22480,N_22059);
and U22680 (N_22680,N_22393,N_22220);
and U22681 (N_22681,N_22479,N_22345);
xor U22682 (N_22682,N_22209,N_22244);
and U22683 (N_22683,N_22228,N_22361);
or U22684 (N_22684,N_22054,N_22019);
xnor U22685 (N_22685,N_22457,N_22171);
nor U22686 (N_22686,N_22051,N_22154);
xor U22687 (N_22687,N_22035,N_22029);
nor U22688 (N_22688,N_22329,N_22198);
nand U22689 (N_22689,N_22034,N_22013);
or U22690 (N_22690,N_22117,N_22233);
nand U22691 (N_22691,N_22369,N_22109);
xnor U22692 (N_22692,N_22210,N_22201);
nand U22693 (N_22693,N_22250,N_22420);
nor U22694 (N_22694,N_22081,N_22046);
xor U22695 (N_22695,N_22459,N_22406);
nand U22696 (N_22696,N_22206,N_22279);
nand U22697 (N_22697,N_22188,N_22387);
or U22698 (N_22698,N_22314,N_22372);
nor U22699 (N_22699,N_22374,N_22359);
nor U22700 (N_22700,N_22342,N_22014);
and U22701 (N_22701,N_22230,N_22070);
or U22702 (N_22702,N_22217,N_22121);
and U22703 (N_22703,N_22159,N_22205);
nand U22704 (N_22704,N_22042,N_22302);
nor U22705 (N_22705,N_22266,N_22193);
or U22706 (N_22706,N_22282,N_22260);
nor U22707 (N_22707,N_22186,N_22212);
nand U22708 (N_22708,N_22182,N_22284);
or U22709 (N_22709,N_22120,N_22321);
nor U22710 (N_22710,N_22463,N_22312);
or U22711 (N_22711,N_22133,N_22272);
and U22712 (N_22712,N_22050,N_22183);
xor U22713 (N_22713,N_22405,N_22487);
nand U22714 (N_22714,N_22246,N_22148);
xnor U22715 (N_22715,N_22118,N_22036);
or U22716 (N_22716,N_22214,N_22432);
or U22717 (N_22717,N_22366,N_22428);
nand U22718 (N_22718,N_22365,N_22245);
nand U22719 (N_22719,N_22440,N_22466);
xnor U22720 (N_22720,N_22110,N_22092);
or U22721 (N_22721,N_22000,N_22079);
or U22722 (N_22722,N_22347,N_22268);
and U22723 (N_22723,N_22339,N_22152);
nand U22724 (N_22724,N_22160,N_22173);
xor U22725 (N_22725,N_22223,N_22240);
nor U22726 (N_22726,N_22411,N_22377);
xnor U22727 (N_22727,N_22290,N_22108);
xnor U22728 (N_22728,N_22001,N_22111);
or U22729 (N_22729,N_22190,N_22482);
and U22730 (N_22730,N_22155,N_22130);
or U22731 (N_22731,N_22264,N_22258);
nand U22732 (N_22732,N_22184,N_22146);
nand U22733 (N_22733,N_22010,N_22338);
nand U22734 (N_22734,N_22135,N_22313);
nand U22735 (N_22735,N_22296,N_22192);
nand U22736 (N_22736,N_22262,N_22351);
or U22737 (N_22737,N_22112,N_22241);
and U22738 (N_22738,N_22232,N_22293);
or U22739 (N_22739,N_22084,N_22048);
nor U22740 (N_22740,N_22061,N_22331);
and U22741 (N_22741,N_22337,N_22484);
xor U22742 (N_22742,N_22310,N_22077);
and U22743 (N_22743,N_22227,N_22094);
xor U22744 (N_22744,N_22274,N_22030);
nand U22745 (N_22745,N_22052,N_22288);
nand U22746 (N_22746,N_22294,N_22322);
or U22747 (N_22747,N_22336,N_22033);
nor U22748 (N_22748,N_22180,N_22483);
or U22749 (N_22749,N_22164,N_22348);
xor U22750 (N_22750,N_22091,N_22460);
and U22751 (N_22751,N_22133,N_22483);
or U22752 (N_22752,N_22398,N_22187);
xnor U22753 (N_22753,N_22048,N_22182);
nand U22754 (N_22754,N_22409,N_22031);
or U22755 (N_22755,N_22208,N_22200);
and U22756 (N_22756,N_22137,N_22024);
nand U22757 (N_22757,N_22218,N_22413);
xnor U22758 (N_22758,N_22153,N_22011);
and U22759 (N_22759,N_22355,N_22385);
and U22760 (N_22760,N_22063,N_22386);
nand U22761 (N_22761,N_22056,N_22176);
and U22762 (N_22762,N_22262,N_22110);
xnor U22763 (N_22763,N_22111,N_22397);
and U22764 (N_22764,N_22234,N_22002);
nand U22765 (N_22765,N_22396,N_22094);
xor U22766 (N_22766,N_22059,N_22320);
nor U22767 (N_22767,N_22172,N_22038);
and U22768 (N_22768,N_22373,N_22248);
and U22769 (N_22769,N_22213,N_22204);
or U22770 (N_22770,N_22334,N_22173);
or U22771 (N_22771,N_22132,N_22408);
and U22772 (N_22772,N_22006,N_22273);
or U22773 (N_22773,N_22154,N_22055);
nand U22774 (N_22774,N_22345,N_22151);
xnor U22775 (N_22775,N_22106,N_22263);
and U22776 (N_22776,N_22483,N_22126);
nand U22777 (N_22777,N_22057,N_22006);
and U22778 (N_22778,N_22498,N_22226);
or U22779 (N_22779,N_22018,N_22173);
nor U22780 (N_22780,N_22232,N_22473);
xnor U22781 (N_22781,N_22372,N_22219);
nor U22782 (N_22782,N_22354,N_22102);
nand U22783 (N_22783,N_22105,N_22106);
xor U22784 (N_22784,N_22220,N_22478);
or U22785 (N_22785,N_22030,N_22230);
xor U22786 (N_22786,N_22433,N_22301);
and U22787 (N_22787,N_22126,N_22147);
nand U22788 (N_22788,N_22379,N_22432);
xor U22789 (N_22789,N_22057,N_22045);
xnor U22790 (N_22790,N_22140,N_22482);
nor U22791 (N_22791,N_22339,N_22444);
nand U22792 (N_22792,N_22352,N_22465);
and U22793 (N_22793,N_22454,N_22368);
and U22794 (N_22794,N_22263,N_22144);
and U22795 (N_22795,N_22209,N_22418);
nor U22796 (N_22796,N_22373,N_22254);
nand U22797 (N_22797,N_22294,N_22265);
nand U22798 (N_22798,N_22026,N_22482);
and U22799 (N_22799,N_22096,N_22352);
nand U22800 (N_22800,N_22305,N_22380);
nor U22801 (N_22801,N_22131,N_22054);
xnor U22802 (N_22802,N_22276,N_22465);
xnor U22803 (N_22803,N_22078,N_22010);
nand U22804 (N_22804,N_22084,N_22034);
nand U22805 (N_22805,N_22261,N_22107);
or U22806 (N_22806,N_22246,N_22007);
nor U22807 (N_22807,N_22124,N_22022);
or U22808 (N_22808,N_22349,N_22485);
and U22809 (N_22809,N_22333,N_22257);
nand U22810 (N_22810,N_22383,N_22376);
nor U22811 (N_22811,N_22033,N_22309);
and U22812 (N_22812,N_22331,N_22391);
nand U22813 (N_22813,N_22187,N_22372);
and U22814 (N_22814,N_22211,N_22229);
nor U22815 (N_22815,N_22366,N_22317);
and U22816 (N_22816,N_22434,N_22217);
and U22817 (N_22817,N_22009,N_22232);
or U22818 (N_22818,N_22008,N_22370);
or U22819 (N_22819,N_22406,N_22027);
nand U22820 (N_22820,N_22022,N_22224);
nor U22821 (N_22821,N_22489,N_22216);
and U22822 (N_22822,N_22021,N_22394);
xor U22823 (N_22823,N_22447,N_22414);
xnor U22824 (N_22824,N_22047,N_22331);
and U22825 (N_22825,N_22092,N_22108);
or U22826 (N_22826,N_22449,N_22331);
xor U22827 (N_22827,N_22404,N_22301);
or U22828 (N_22828,N_22420,N_22059);
xor U22829 (N_22829,N_22120,N_22457);
nor U22830 (N_22830,N_22222,N_22089);
nand U22831 (N_22831,N_22426,N_22082);
xnor U22832 (N_22832,N_22462,N_22469);
or U22833 (N_22833,N_22442,N_22483);
nand U22834 (N_22834,N_22065,N_22363);
xor U22835 (N_22835,N_22461,N_22170);
and U22836 (N_22836,N_22415,N_22480);
or U22837 (N_22837,N_22239,N_22060);
or U22838 (N_22838,N_22259,N_22407);
xor U22839 (N_22839,N_22246,N_22105);
nor U22840 (N_22840,N_22273,N_22466);
xnor U22841 (N_22841,N_22294,N_22134);
or U22842 (N_22842,N_22372,N_22112);
or U22843 (N_22843,N_22074,N_22270);
nand U22844 (N_22844,N_22464,N_22182);
xnor U22845 (N_22845,N_22424,N_22330);
nand U22846 (N_22846,N_22200,N_22440);
nand U22847 (N_22847,N_22257,N_22457);
or U22848 (N_22848,N_22088,N_22136);
or U22849 (N_22849,N_22255,N_22279);
or U22850 (N_22850,N_22349,N_22169);
xor U22851 (N_22851,N_22247,N_22236);
or U22852 (N_22852,N_22149,N_22032);
nor U22853 (N_22853,N_22157,N_22401);
and U22854 (N_22854,N_22274,N_22369);
nor U22855 (N_22855,N_22303,N_22146);
nor U22856 (N_22856,N_22396,N_22474);
xnor U22857 (N_22857,N_22357,N_22226);
nor U22858 (N_22858,N_22132,N_22001);
nor U22859 (N_22859,N_22014,N_22442);
xor U22860 (N_22860,N_22299,N_22235);
nand U22861 (N_22861,N_22046,N_22301);
or U22862 (N_22862,N_22480,N_22478);
and U22863 (N_22863,N_22176,N_22015);
and U22864 (N_22864,N_22231,N_22086);
and U22865 (N_22865,N_22214,N_22257);
or U22866 (N_22866,N_22251,N_22194);
and U22867 (N_22867,N_22336,N_22107);
nor U22868 (N_22868,N_22418,N_22382);
nand U22869 (N_22869,N_22334,N_22261);
and U22870 (N_22870,N_22293,N_22408);
xnor U22871 (N_22871,N_22089,N_22207);
nor U22872 (N_22872,N_22161,N_22323);
nor U22873 (N_22873,N_22066,N_22225);
or U22874 (N_22874,N_22272,N_22390);
nor U22875 (N_22875,N_22086,N_22471);
and U22876 (N_22876,N_22344,N_22432);
nor U22877 (N_22877,N_22202,N_22326);
or U22878 (N_22878,N_22014,N_22310);
and U22879 (N_22879,N_22386,N_22183);
and U22880 (N_22880,N_22247,N_22435);
nor U22881 (N_22881,N_22238,N_22022);
xor U22882 (N_22882,N_22026,N_22460);
nand U22883 (N_22883,N_22363,N_22345);
or U22884 (N_22884,N_22293,N_22010);
or U22885 (N_22885,N_22016,N_22242);
and U22886 (N_22886,N_22136,N_22446);
or U22887 (N_22887,N_22449,N_22069);
nand U22888 (N_22888,N_22169,N_22414);
nor U22889 (N_22889,N_22075,N_22338);
nor U22890 (N_22890,N_22385,N_22168);
or U22891 (N_22891,N_22350,N_22248);
or U22892 (N_22892,N_22253,N_22262);
xor U22893 (N_22893,N_22094,N_22155);
or U22894 (N_22894,N_22152,N_22199);
xor U22895 (N_22895,N_22099,N_22150);
and U22896 (N_22896,N_22101,N_22032);
nor U22897 (N_22897,N_22036,N_22152);
or U22898 (N_22898,N_22384,N_22009);
and U22899 (N_22899,N_22084,N_22140);
and U22900 (N_22900,N_22138,N_22410);
or U22901 (N_22901,N_22218,N_22335);
and U22902 (N_22902,N_22462,N_22360);
and U22903 (N_22903,N_22402,N_22276);
nor U22904 (N_22904,N_22193,N_22043);
nand U22905 (N_22905,N_22117,N_22335);
nor U22906 (N_22906,N_22127,N_22032);
xnor U22907 (N_22907,N_22306,N_22007);
and U22908 (N_22908,N_22219,N_22095);
nand U22909 (N_22909,N_22185,N_22499);
nor U22910 (N_22910,N_22359,N_22208);
and U22911 (N_22911,N_22092,N_22278);
nand U22912 (N_22912,N_22000,N_22313);
xnor U22913 (N_22913,N_22343,N_22421);
xnor U22914 (N_22914,N_22365,N_22423);
nor U22915 (N_22915,N_22256,N_22174);
and U22916 (N_22916,N_22499,N_22020);
nor U22917 (N_22917,N_22251,N_22162);
and U22918 (N_22918,N_22199,N_22237);
nand U22919 (N_22919,N_22295,N_22242);
nand U22920 (N_22920,N_22385,N_22222);
nor U22921 (N_22921,N_22324,N_22004);
and U22922 (N_22922,N_22138,N_22190);
nand U22923 (N_22923,N_22431,N_22438);
or U22924 (N_22924,N_22106,N_22382);
xor U22925 (N_22925,N_22383,N_22470);
nor U22926 (N_22926,N_22114,N_22020);
nor U22927 (N_22927,N_22445,N_22287);
and U22928 (N_22928,N_22425,N_22108);
and U22929 (N_22929,N_22441,N_22185);
nor U22930 (N_22930,N_22074,N_22063);
or U22931 (N_22931,N_22297,N_22466);
or U22932 (N_22932,N_22035,N_22483);
and U22933 (N_22933,N_22083,N_22033);
nand U22934 (N_22934,N_22362,N_22263);
xnor U22935 (N_22935,N_22106,N_22299);
and U22936 (N_22936,N_22245,N_22437);
and U22937 (N_22937,N_22077,N_22398);
and U22938 (N_22938,N_22352,N_22385);
and U22939 (N_22939,N_22487,N_22077);
nand U22940 (N_22940,N_22175,N_22158);
or U22941 (N_22941,N_22197,N_22478);
nor U22942 (N_22942,N_22036,N_22489);
nor U22943 (N_22943,N_22400,N_22044);
and U22944 (N_22944,N_22482,N_22039);
and U22945 (N_22945,N_22113,N_22439);
and U22946 (N_22946,N_22328,N_22207);
xnor U22947 (N_22947,N_22200,N_22405);
xor U22948 (N_22948,N_22308,N_22112);
or U22949 (N_22949,N_22056,N_22239);
nand U22950 (N_22950,N_22407,N_22398);
and U22951 (N_22951,N_22108,N_22144);
or U22952 (N_22952,N_22274,N_22421);
nand U22953 (N_22953,N_22346,N_22383);
xnor U22954 (N_22954,N_22216,N_22141);
nand U22955 (N_22955,N_22159,N_22495);
xnor U22956 (N_22956,N_22281,N_22370);
or U22957 (N_22957,N_22093,N_22458);
or U22958 (N_22958,N_22248,N_22482);
or U22959 (N_22959,N_22300,N_22354);
or U22960 (N_22960,N_22322,N_22062);
or U22961 (N_22961,N_22335,N_22364);
or U22962 (N_22962,N_22422,N_22091);
xor U22963 (N_22963,N_22102,N_22388);
nor U22964 (N_22964,N_22191,N_22161);
and U22965 (N_22965,N_22093,N_22129);
nor U22966 (N_22966,N_22316,N_22089);
nand U22967 (N_22967,N_22246,N_22058);
and U22968 (N_22968,N_22416,N_22144);
xnor U22969 (N_22969,N_22188,N_22484);
nand U22970 (N_22970,N_22063,N_22010);
nor U22971 (N_22971,N_22055,N_22038);
nor U22972 (N_22972,N_22394,N_22334);
nand U22973 (N_22973,N_22453,N_22292);
and U22974 (N_22974,N_22274,N_22241);
nand U22975 (N_22975,N_22182,N_22108);
or U22976 (N_22976,N_22222,N_22012);
or U22977 (N_22977,N_22166,N_22440);
nor U22978 (N_22978,N_22487,N_22480);
nor U22979 (N_22979,N_22064,N_22116);
or U22980 (N_22980,N_22432,N_22482);
nor U22981 (N_22981,N_22005,N_22450);
xor U22982 (N_22982,N_22034,N_22001);
nor U22983 (N_22983,N_22357,N_22321);
nand U22984 (N_22984,N_22494,N_22437);
nor U22985 (N_22985,N_22166,N_22110);
nor U22986 (N_22986,N_22193,N_22190);
xor U22987 (N_22987,N_22152,N_22013);
and U22988 (N_22988,N_22181,N_22137);
and U22989 (N_22989,N_22368,N_22456);
nand U22990 (N_22990,N_22127,N_22439);
and U22991 (N_22991,N_22045,N_22215);
nand U22992 (N_22992,N_22175,N_22269);
or U22993 (N_22993,N_22340,N_22133);
or U22994 (N_22994,N_22412,N_22273);
and U22995 (N_22995,N_22083,N_22472);
xnor U22996 (N_22996,N_22010,N_22343);
xor U22997 (N_22997,N_22033,N_22069);
xor U22998 (N_22998,N_22275,N_22193);
and U22999 (N_22999,N_22240,N_22039);
or U23000 (N_23000,N_22982,N_22664);
xor U23001 (N_23001,N_22667,N_22783);
and U23002 (N_23002,N_22796,N_22518);
or U23003 (N_23003,N_22539,N_22703);
nand U23004 (N_23004,N_22613,N_22617);
nor U23005 (N_23005,N_22891,N_22719);
and U23006 (N_23006,N_22793,N_22627);
xor U23007 (N_23007,N_22663,N_22780);
or U23008 (N_23008,N_22556,N_22749);
or U23009 (N_23009,N_22750,N_22923);
or U23010 (N_23010,N_22665,N_22880);
nand U23011 (N_23011,N_22771,N_22991);
nor U23012 (N_23012,N_22971,N_22887);
xnor U23013 (N_23013,N_22946,N_22616);
and U23014 (N_23014,N_22961,N_22715);
and U23015 (N_23015,N_22552,N_22945);
nor U23016 (N_23016,N_22547,N_22799);
nand U23017 (N_23017,N_22936,N_22521);
or U23018 (N_23018,N_22953,N_22758);
and U23019 (N_23019,N_22943,N_22563);
or U23020 (N_23020,N_22840,N_22984);
nand U23021 (N_23021,N_22735,N_22754);
nor U23022 (N_23022,N_22713,N_22975);
nand U23023 (N_23023,N_22721,N_22583);
or U23024 (N_23024,N_22965,N_22952);
xnor U23025 (N_23025,N_22841,N_22906);
xor U23026 (N_23026,N_22918,N_22836);
nand U23027 (N_23027,N_22543,N_22890);
xor U23028 (N_23028,N_22960,N_22578);
or U23029 (N_23029,N_22893,N_22531);
xor U23030 (N_23030,N_22888,N_22673);
and U23031 (N_23031,N_22859,N_22768);
nand U23032 (N_23032,N_22761,N_22803);
or U23033 (N_23033,N_22541,N_22509);
nand U23034 (N_23034,N_22620,N_22564);
and U23035 (N_23035,N_22660,N_22827);
nand U23036 (N_23036,N_22698,N_22864);
xnor U23037 (N_23037,N_22897,N_22789);
nand U23038 (N_23038,N_22769,N_22901);
xor U23039 (N_23039,N_22992,N_22561);
and U23040 (N_23040,N_22767,N_22808);
and U23041 (N_23041,N_22656,N_22886);
xnor U23042 (N_23042,N_22516,N_22681);
nor U23043 (N_23043,N_22702,N_22643);
nand U23044 (N_23044,N_22637,N_22668);
xor U23045 (N_23045,N_22559,N_22802);
nor U23046 (N_23046,N_22650,N_22527);
nand U23047 (N_23047,N_22804,N_22981);
or U23048 (N_23048,N_22869,N_22636);
or U23049 (N_23049,N_22874,N_22909);
nand U23050 (N_23050,N_22959,N_22844);
or U23051 (N_23051,N_22582,N_22677);
or U23052 (N_23052,N_22528,N_22845);
and U23053 (N_23053,N_22514,N_22725);
and U23054 (N_23054,N_22565,N_22862);
or U23055 (N_23055,N_22995,N_22898);
nor U23056 (N_23056,N_22977,N_22674);
nor U23057 (N_23057,N_22553,N_22927);
and U23058 (N_23058,N_22608,N_22957);
xor U23059 (N_23059,N_22649,N_22776);
nor U23060 (N_23060,N_22594,N_22996);
xor U23061 (N_23061,N_22655,N_22885);
nand U23062 (N_23062,N_22586,N_22525);
and U23063 (N_23063,N_22630,N_22595);
nand U23064 (N_23064,N_22837,N_22512);
nand U23065 (N_23065,N_22732,N_22700);
nand U23066 (N_23066,N_22603,N_22574);
nand U23067 (N_23067,N_22504,N_22588);
xor U23068 (N_23068,N_22645,N_22612);
nor U23069 (N_23069,N_22666,N_22648);
and U23070 (N_23070,N_22654,N_22904);
nand U23071 (N_23071,N_22724,N_22892);
nor U23072 (N_23072,N_22611,N_22966);
nor U23073 (N_23073,N_22680,N_22598);
nor U23074 (N_23074,N_22640,N_22867);
nor U23075 (N_23075,N_22903,N_22696);
nand U23076 (N_23076,N_22810,N_22711);
xnor U23077 (N_23077,N_22733,N_22591);
xnor U23078 (N_23078,N_22860,N_22765);
xnor U23079 (N_23079,N_22999,N_22872);
nor U23080 (N_23080,N_22832,N_22694);
xor U23081 (N_23081,N_22989,N_22942);
and U23082 (N_23082,N_22917,N_22778);
and U23083 (N_23083,N_22653,N_22670);
nor U23084 (N_23084,N_22753,N_22931);
nor U23085 (N_23085,N_22596,N_22882);
nor U23086 (N_23086,N_22939,N_22729);
nor U23087 (N_23087,N_22642,N_22523);
and U23088 (N_23088,N_22628,N_22838);
nand U23089 (N_23089,N_22795,N_22508);
xor U23090 (N_23090,N_22770,N_22902);
nand U23091 (N_23091,N_22605,N_22562);
nor U23092 (N_23092,N_22911,N_22947);
or U23093 (N_23093,N_22878,N_22671);
xnor U23094 (N_23094,N_22881,N_22817);
nor U23095 (N_23095,N_22772,N_22631);
xor U23096 (N_23096,N_22532,N_22932);
or U23097 (N_23097,N_22956,N_22720);
nand U23098 (N_23098,N_22619,N_22752);
nand U23099 (N_23099,N_22592,N_22730);
and U23100 (N_23100,N_22584,N_22905);
nand U23101 (N_23101,N_22699,N_22658);
nand U23102 (N_23102,N_22820,N_22575);
nand U23103 (N_23103,N_22533,N_22690);
or U23104 (N_23104,N_22922,N_22784);
and U23105 (N_23105,N_22585,N_22756);
or U23106 (N_23106,N_22507,N_22744);
or U23107 (N_23107,N_22950,N_22842);
xor U23108 (N_23108,N_22938,N_22614);
or U23109 (N_23109,N_22983,N_22572);
or U23110 (N_23110,N_22825,N_22590);
nand U23111 (N_23111,N_22566,N_22689);
or U23112 (N_23112,N_22538,N_22863);
nand U23113 (N_23113,N_22958,N_22546);
nand U23114 (N_23114,N_22550,N_22548);
nor U23115 (N_23115,N_22970,N_22624);
nor U23116 (N_23116,N_22933,N_22912);
and U23117 (N_23117,N_22638,N_22745);
and U23118 (N_23118,N_22714,N_22900);
nand U23119 (N_23119,N_22661,N_22914);
nand U23120 (N_23120,N_22625,N_22751);
nand U23121 (N_23121,N_22540,N_22526);
nor U23122 (N_23122,N_22686,N_22928);
nor U23123 (N_23123,N_22641,N_22651);
nor U23124 (N_23124,N_22717,N_22916);
nand U23125 (N_23125,N_22988,N_22895);
and U23126 (N_23126,N_22978,N_22522);
nand U23127 (N_23127,N_22974,N_22899);
xor U23128 (N_23128,N_22763,N_22728);
and U23129 (N_23129,N_22814,N_22779);
and U23130 (N_23130,N_22632,N_22781);
nor U23131 (N_23131,N_22513,N_22894);
xor U23132 (N_23132,N_22519,N_22524);
xor U23133 (N_23133,N_22908,N_22822);
or U23134 (N_23134,N_22697,N_22707);
xnor U23135 (N_23135,N_22774,N_22748);
nand U23136 (N_23136,N_22785,N_22951);
nor U23137 (N_23137,N_22581,N_22934);
xnor U23138 (N_23138,N_22839,N_22693);
nand U23139 (N_23139,N_22811,N_22879);
and U23140 (N_23140,N_22766,N_22791);
nand U23141 (N_23141,N_22558,N_22587);
nor U23142 (N_23142,N_22662,N_22850);
and U23143 (N_23143,N_22722,N_22871);
nand U23144 (N_23144,N_22747,N_22963);
and U23145 (N_23145,N_22821,N_22683);
and U23146 (N_23146,N_22557,N_22705);
and U23147 (N_23147,N_22600,N_22964);
xor U23148 (N_23148,N_22846,N_22618);
xor U23149 (N_23149,N_22503,N_22819);
nand U23150 (N_23150,N_22985,N_22742);
xnor U23151 (N_23151,N_22935,N_22604);
nand U23152 (N_23152,N_22775,N_22551);
xor U23153 (N_23153,N_22968,N_22736);
nand U23154 (N_23154,N_22834,N_22571);
or U23155 (N_23155,N_22855,N_22955);
nand U23156 (N_23156,N_22568,N_22607);
and U23157 (N_23157,N_22716,N_22746);
nand U23158 (N_23158,N_22828,N_22506);
nor U23159 (N_23159,N_22500,N_22907);
nor U23160 (N_23160,N_22994,N_22852);
nand U23161 (N_23161,N_22998,N_22520);
nand U23162 (N_23162,N_22826,N_22738);
nand U23163 (N_23163,N_22569,N_22517);
xnor U23164 (N_23164,N_22921,N_22815);
nand U23165 (N_23165,N_22857,N_22913);
and U23166 (N_23166,N_22812,N_22731);
and U23167 (N_23167,N_22635,N_22997);
nand U23168 (N_23168,N_22669,N_22755);
xor U23169 (N_23169,N_22510,N_22726);
nor U23170 (N_23170,N_22773,N_22876);
xnor U23171 (N_23171,N_22861,N_22829);
nor U23172 (N_23172,N_22831,N_22589);
or U23173 (N_23173,N_22708,N_22823);
and U23174 (N_23174,N_22626,N_22925);
nand U23175 (N_23175,N_22830,N_22739);
or U23176 (N_23176,N_22554,N_22801);
xnor U23177 (N_23177,N_22623,N_22684);
and U23178 (N_23178,N_22601,N_22987);
or U23179 (N_23179,N_22877,N_22807);
or U23180 (N_23180,N_22760,N_22606);
nor U23181 (N_23181,N_22941,N_22579);
nand U23182 (N_23182,N_22549,N_22972);
and U23183 (N_23183,N_22597,N_22743);
xor U23184 (N_23184,N_22816,N_22884);
xor U23185 (N_23185,N_22515,N_22502);
and U23186 (N_23186,N_22639,N_22621);
nor U23187 (N_23187,N_22709,N_22692);
xnor U23188 (N_23188,N_22593,N_22727);
xor U23189 (N_23189,N_22764,N_22809);
nor U23190 (N_23190,N_22759,N_22962);
nand U23191 (N_23191,N_22622,N_22573);
nand U23192 (N_23192,N_22937,N_22602);
and U23193 (N_23193,N_22542,N_22737);
nand U23194 (N_23194,N_22560,N_22915);
nand U23195 (N_23195,N_22870,N_22976);
or U23196 (N_23196,N_22610,N_22954);
xor U23197 (N_23197,N_22687,N_22659);
nand U23198 (N_23198,N_22986,N_22967);
nand U23199 (N_23199,N_22944,N_22723);
or U23200 (N_23200,N_22740,N_22672);
nor U23201 (N_23201,N_22993,N_22536);
nand U23202 (N_23202,N_22940,N_22534);
nor U23203 (N_23203,N_22688,N_22695);
and U23204 (N_23204,N_22919,N_22990);
xnor U23205 (N_23205,N_22644,N_22501);
or U23206 (N_23206,N_22675,N_22949);
nor U23207 (N_23207,N_22741,N_22896);
and U23208 (N_23208,N_22813,N_22576);
or U23209 (N_23209,N_22511,N_22798);
and U23210 (N_23210,N_22875,N_22792);
xnor U23211 (N_23211,N_22777,N_22920);
and U23212 (N_23212,N_22924,N_22570);
and U23213 (N_23213,N_22609,N_22657);
nand U23214 (N_23214,N_22718,N_22847);
xor U23215 (N_23215,N_22567,N_22866);
nand U23216 (N_23216,N_22529,N_22678);
nor U23217 (N_23217,N_22910,N_22926);
xor U23218 (N_23218,N_22646,N_22762);
and U23219 (N_23219,N_22633,N_22979);
nand U23220 (N_23220,N_22599,N_22883);
and U23221 (N_23221,N_22544,N_22757);
or U23222 (N_23222,N_22889,N_22856);
nand U23223 (N_23223,N_22634,N_22858);
nand U23224 (N_23224,N_22704,N_22930);
xor U23225 (N_23225,N_22849,N_22629);
nor U23226 (N_23226,N_22787,N_22682);
nand U23227 (N_23227,N_22853,N_22797);
nor U23228 (N_23228,N_22580,N_22710);
or U23229 (N_23229,N_22685,N_22555);
nor U23230 (N_23230,N_22805,N_22868);
nor U23231 (N_23231,N_22865,N_22833);
nand U23232 (N_23232,N_22577,N_22980);
or U23233 (N_23233,N_22535,N_22691);
nand U23234 (N_23234,N_22782,N_22537);
nand U23235 (N_23235,N_22545,N_22843);
or U23236 (N_23236,N_22676,N_22973);
nor U23237 (N_23237,N_22530,N_22835);
nand U23238 (N_23238,N_22712,N_22854);
nor U23239 (N_23239,N_22615,N_22734);
or U23240 (N_23240,N_22806,N_22848);
and U23241 (N_23241,N_22948,N_22652);
nand U23242 (N_23242,N_22873,N_22794);
or U23243 (N_23243,N_22679,N_22788);
xnor U23244 (N_23244,N_22505,N_22824);
nor U23245 (N_23245,N_22929,N_22706);
and U23246 (N_23246,N_22786,N_22818);
and U23247 (N_23247,N_22647,N_22800);
nand U23248 (N_23248,N_22851,N_22969);
and U23249 (N_23249,N_22701,N_22790);
xor U23250 (N_23250,N_22775,N_22951);
or U23251 (N_23251,N_22958,N_22665);
xor U23252 (N_23252,N_22823,N_22946);
or U23253 (N_23253,N_22815,N_22842);
nand U23254 (N_23254,N_22542,N_22545);
xor U23255 (N_23255,N_22514,N_22940);
and U23256 (N_23256,N_22578,N_22507);
xor U23257 (N_23257,N_22594,N_22727);
xnor U23258 (N_23258,N_22765,N_22658);
nand U23259 (N_23259,N_22923,N_22690);
or U23260 (N_23260,N_22885,N_22614);
or U23261 (N_23261,N_22732,N_22675);
or U23262 (N_23262,N_22605,N_22701);
and U23263 (N_23263,N_22791,N_22687);
xnor U23264 (N_23264,N_22585,N_22711);
nand U23265 (N_23265,N_22882,N_22727);
and U23266 (N_23266,N_22615,N_22579);
nor U23267 (N_23267,N_22952,N_22846);
or U23268 (N_23268,N_22798,N_22941);
and U23269 (N_23269,N_22862,N_22885);
and U23270 (N_23270,N_22953,N_22857);
and U23271 (N_23271,N_22989,N_22727);
nand U23272 (N_23272,N_22695,N_22710);
nand U23273 (N_23273,N_22897,N_22530);
and U23274 (N_23274,N_22858,N_22960);
or U23275 (N_23275,N_22992,N_22606);
nor U23276 (N_23276,N_22622,N_22923);
or U23277 (N_23277,N_22692,N_22984);
xor U23278 (N_23278,N_22541,N_22964);
xnor U23279 (N_23279,N_22984,N_22875);
xor U23280 (N_23280,N_22695,N_22707);
and U23281 (N_23281,N_22552,N_22681);
nor U23282 (N_23282,N_22528,N_22934);
nand U23283 (N_23283,N_22674,N_22577);
nand U23284 (N_23284,N_22873,N_22593);
nor U23285 (N_23285,N_22989,N_22654);
and U23286 (N_23286,N_22700,N_22548);
xnor U23287 (N_23287,N_22795,N_22654);
nor U23288 (N_23288,N_22528,N_22666);
nor U23289 (N_23289,N_22567,N_22532);
xor U23290 (N_23290,N_22555,N_22930);
and U23291 (N_23291,N_22556,N_22854);
nand U23292 (N_23292,N_22505,N_22536);
and U23293 (N_23293,N_22939,N_22525);
and U23294 (N_23294,N_22966,N_22992);
xor U23295 (N_23295,N_22849,N_22604);
or U23296 (N_23296,N_22501,N_22597);
and U23297 (N_23297,N_22670,N_22767);
nor U23298 (N_23298,N_22955,N_22796);
nor U23299 (N_23299,N_22723,N_22503);
nor U23300 (N_23300,N_22514,N_22892);
or U23301 (N_23301,N_22587,N_22930);
nor U23302 (N_23302,N_22551,N_22725);
nor U23303 (N_23303,N_22931,N_22624);
and U23304 (N_23304,N_22670,N_22954);
or U23305 (N_23305,N_22569,N_22989);
or U23306 (N_23306,N_22686,N_22728);
or U23307 (N_23307,N_22835,N_22932);
and U23308 (N_23308,N_22736,N_22807);
and U23309 (N_23309,N_22749,N_22635);
xnor U23310 (N_23310,N_22763,N_22720);
or U23311 (N_23311,N_22901,N_22925);
nand U23312 (N_23312,N_22822,N_22643);
nand U23313 (N_23313,N_22646,N_22994);
or U23314 (N_23314,N_22563,N_22822);
and U23315 (N_23315,N_22888,N_22926);
nand U23316 (N_23316,N_22883,N_22641);
nor U23317 (N_23317,N_22634,N_22874);
xnor U23318 (N_23318,N_22976,N_22711);
and U23319 (N_23319,N_22535,N_22653);
xnor U23320 (N_23320,N_22692,N_22637);
or U23321 (N_23321,N_22505,N_22570);
xnor U23322 (N_23322,N_22815,N_22947);
nor U23323 (N_23323,N_22627,N_22790);
xor U23324 (N_23324,N_22965,N_22637);
xor U23325 (N_23325,N_22606,N_22971);
or U23326 (N_23326,N_22608,N_22995);
and U23327 (N_23327,N_22555,N_22518);
and U23328 (N_23328,N_22915,N_22883);
and U23329 (N_23329,N_22633,N_22728);
nand U23330 (N_23330,N_22779,N_22769);
nand U23331 (N_23331,N_22635,N_22809);
xnor U23332 (N_23332,N_22597,N_22778);
xnor U23333 (N_23333,N_22627,N_22734);
nor U23334 (N_23334,N_22672,N_22915);
and U23335 (N_23335,N_22951,N_22649);
and U23336 (N_23336,N_22893,N_22589);
and U23337 (N_23337,N_22607,N_22882);
nand U23338 (N_23338,N_22725,N_22914);
and U23339 (N_23339,N_22820,N_22902);
and U23340 (N_23340,N_22955,N_22548);
nor U23341 (N_23341,N_22857,N_22589);
xor U23342 (N_23342,N_22703,N_22631);
and U23343 (N_23343,N_22707,N_22846);
or U23344 (N_23344,N_22526,N_22649);
or U23345 (N_23345,N_22964,N_22862);
or U23346 (N_23346,N_22886,N_22754);
nor U23347 (N_23347,N_22663,N_22511);
nand U23348 (N_23348,N_22749,N_22794);
and U23349 (N_23349,N_22960,N_22642);
xnor U23350 (N_23350,N_22680,N_22660);
xnor U23351 (N_23351,N_22719,N_22543);
or U23352 (N_23352,N_22694,N_22917);
xnor U23353 (N_23353,N_22583,N_22930);
or U23354 (N_23354,N_22531,N_22935);
and U23355 (N_23355,N_22558,N_22542);
nor U23356 (N_23356,N_22524,N_22819);
nand U23357 (N_23357,N_22739,N_22580);
xor U23358 (N_23358,N_22832,N_22574);
and U23359 (N_23359,N_22994,N_22712);
xor U23360 (N_23360,N_22951,N_22637);
nand U23361 (N_23361,N_22527,N_22815);
nand U23362 (N_23362,N_22663,N_22702);
or U23363 (N_23363,N_22961,N_22949);
xnor U23364 (N_23364,N_22670,N_22590);
or U23365 (N_23365,N_22939,N_22536);
nor U23366 (N_23366,N_22629,N_22565);
and U23367 (N_23367,N_22993,N_22808);
nand U23368 (N_23368,N_22557,N_22685);
xnor U23369 (N_23369,N_22951,N_22930);
nand U23370 (N_23370,N_22839,N_22780);
nor U23371 (N_23371,N_22659,N_22637);
or U23372 (N_23372,N_22778,N_22649);
nand U23373 (N_23373,N_22758,N_22638);
or U23374 (N_23374,N_22981,N_22823);
nand U23375 (N_23375,N_22838,N_22599);
nor U23376 (N_23376,N_22899,N_22552);
and U23377 (N_23377,N_22858,N_22502);
xor U23378 (N_23378,N_22611,N_22552);
nor U23379 (N_23379,N_22933,N_22880);
and U23380 (N_23380,N_22547,N_22731);
xor U23381 (N_23381,N_22758,N_22797);
nand U23382 (N_23382,N_22974,N_22582);
xnor U23383 (N_23383,N_22927,N_22906);
nor U23384 (N_23384,N_22745,N_22845);
or U23385 (N_23385,N_22752,N_22622);
xor U23386 (N_23386,N_22607,N_22577);
or U23387 (N_23387,N_22585,N_22781);
xor U23388 (N_23388,N_22943,N_22994);
or U23389 (N_23389,N_22938,N_22959);
and U23390 (N_23390,N_22542,N_22654);
nand U23391 (N_23391,N_22669,N_22919);
nor U23392 (N_23392,N_22778,N_22744);
xnor U23393 (N_23393,N_22956,N_22671);
xnor U23394 (N_23394,N_22809,N_22717);
nor U23395 (N_23395,N_22599,N_22834);
and U23396 (N_23396,N_22951,N_22572);
and U23397 (N_23397,N_22718,N_22959);
xor U23398 (N_23398,N_22748,N_22620);
or U23399 (N_23399,N_22968,N_22730);
nand U23400 (N_23400,N_22776,N_22642);
nor U23401 (N_23401,N_22510,N_22889);
xor U23402 (N_23402,N_22575,N_22698);
nor U23403 (N_23403,N_22579,N_22823);
nand U23404 (N_23404,N_22912,N_22735);
xnor U23405 (N_23405,N_22883,N_22970);
and U23406 (N_23406,N_22740,N_22664);
nor U23407 (N_23407,N_22597,N_22810);
or U23408 (N_23408,N_22726,N_22825);
xor U23409 (N_23409,N_22713,N_22654);
and U23410 (N_23410,N_22984,N_22625);
nand U23411 (N_23411,N_22637,N_22826);
and U23412 (N_23412,N_22842,N_22545);
and U23413 (N_23413,N_22582,N_22781);
xnor U23414 (N_23414,N_22654,N_22735);
or U23415 (N_23415,N_22869,N_22735);
or U23416 (N_23416,N_22686,N_22631);
nor U23417 (N_23417,N_22978,N_22546);
xnor U23418 (N_23418,N_22546,N_22579);
nor U23419 (N_23419,N_22756,N_22894);
nand U23420 (N_23420,N_22833,N_22628);
nor U23421 (N_23421,N_22916,N_22831);
xnor U23422 (N_23422,N_22615,N_22865);
and U23423 (N_23423,N_22875,N_22996);
nand U23424 (N_23424,N_22816,N_22579);
nor U23425 (N_23425,N_22579,N_22893);
nand U23426 (N_23426,N_22570,N_22792);
nor U23427 (N_23427,N_22591,N_22661);
and U23428 (N_23428,N_22801,N_22912);
or U23429 (N_23429,N_22656,N_22599);
or U23430 (N_23430,N_22759,N_22914);
nor U23431 (N_23431,N_22873,N_22906);
xor U23432 (N_23432,N_22842,N_22690);
xnor U23433 (N_23433,N_22552,N_22626);
or U23434 (N_23434,N_22870,N_22932);
or U23435 (N_23435,N_22984,N_22798);
xor U23436 (N_23436,N_22565,N_22833);
xor U23437 (N_23437,N_22661,N_22957);
and U23438 (N_23438,N_22948,N_22564);
xor U23439 (N_23439,N_22875,N_22518);
nand U23440 (N_23440,N_22848,N_22987);
or U23441 (N_23441,N_22876,N_22819);
and U23442 (N_23442,N_22609,N_22739);
or U23443 (N_23443,N_22975,N_22922);
nand U23444 (N_23444,N_22573,N_22751);
xnor U23445 (N_23445,N_22610,N_22584);
nor U23446 (N_23446,N_22969,N_22629);
xor U23447 (N_23447,N_22840,N_22512);
or U23448 (N_23448,N_22577,N_22669);
xnor U23449 (N_23449,N_22960,N_22874);
nand U23450 (N_23450,N_22704,N_22557);
and U23451 (N_23451,N_22914,N_22691);
or U23452 (N_23452,N_22801,N_22900);
or U23453 (N_23453,N_22941,N_22785);
and U23454 (N_23454,N_22651,N_22541);
and U23455 (N_23455,N_22638,N_22547);
xnor U23456 (N_23456,N_22552,N_22823);
or U23457 (N_23457,N_22592,N_22722);
xnor U23458 (N_23458,N_22778,N_22994);
nor U23459 (N_23459,N_22706,N_22750);
and U23460 (N_23460,N_22800,N_22510);
nand U23461 (N_23461,N_22685,N_22592);
nand U23462 (N_23462,N_22708,N_22589);
nand U23463 (N_23463,N_22763,N_22963);
and U23464 (N_23464,N_22694,N_22750);
and U23465 (N_23465,N_22872,N_22641);
xor U23466 (N_23466,N_22968,N_22790);
or U23467 (N_23467,N_22775,N_22948);
and U23468 (N_23468,N_22613,N_22577);
xnor U23469 (N_23469,N_22806,N_22970);
or U23470 (N_23470,N_22599,N_22886);
xnor U23471 (N_23471,N_22647,N_22859);
nand U23472 (N_23472,N_22540,N_22634);
or U23473 (N_23473,N_22645,N_22738);
nor U23474 (N_23474,N_22757,N_22503);
nand U23475 (N_23475,N_22674,N_22523);
nor U23476 (N_23476,N_22571,N_22774);
and U23477 (N_23477,N_22788,N_22726);
nand U23478 (N_23478,N_22877,N_22705);
nor U23479 (N_23479,N_22957,N_22931);
and U23480 (N_23480,N_22917,N_22578);
xnor U23481 (N_23481,N_22803,N_22915);
and U23482 (N_23482,N_22781,N_22680);
xnor U23483 (N_23483,N_22700,N_22643);
and U23484 (N_23484,N_22641,N_22501);
nor U23485 (N_23485,N_22513,N_22717);
nor U23486 (N_23486,N_22674,N_22500);
and U23487 (N_23487,N_22615,N_22790);
xnor U23488 (N_23488,N_22612,N_22727);
nor U23489 (N_23489,N_22817,N_22912);
nor U23490 (N_23490,N_22636,N_22756);
and U23491 (N_23491,N_22774,N_22796);
or U23492 (N_23492,N_22671,N_22890);
nor U23493 (N_23493,N_22647,N_22555);
and U23494 (N_23494,N_22739,N_22773);
nor U23495 (N_23495,N_22542,N_22728);
or U23496 (N_23496,N_22780,N_22545);
nand U23497 (N_23497,N_22796,N_22861);
xnor U23498 (N_23498,N_22547,N_22506);
and U23499 (N_23499,N_22912,N_22527);
xnor U23500 (N_23500,N_23156,N_23251);
xor U23501 (N_23501,N_23287,N_23270);
and U23502 (N_23502,N_23348,N_23434);
xor U23503 (N_23503,N_23247,N_23312);
nor U23504 (N_23504,N_23030,N_23412);
nand U23505 (N_23505,N_23281,N_23289);
or U23506 (N_23506,N_23228,N_23387);
or U23507 (N_23507,N_23186,N_23246);
xnor U23508 (N_23508,N_23341,N_23305);
and U23509 (N_23509,N_23410,N_23005);
or U23510 (N_23510,N_23469,N_23211);
nor U23511 (N_23511,N_23429,N_23350);
nand U23512 (N_23512,N_23214,N_23200);
or U23513 (N_23513,N_23315,N_23314);
nor U23514 (N_23514,N_23295,N_23174);
or U23515 (N_23515,N_23282,N_23013);
nor U23516 (N_23516,N_23226,N_23032);
or U23517 (N_23517,N_23206,N_23274);
nand U23518 (N_23518,N_23094,N_23385);
nor U23519 (N_23519,N_23166,N_23450);
nor U23520 (N_23520,N_23235,N_23024);
and U23521 (N_23521,N_23271,N_23140);
or U23522 (N_23522,N_23203,N_23275);
nand U23523 (N_23523,N_23382,N_23327);
nor U23524 (N_23524,N_23239,N_23119);
and U23525 (N_23525,N_23234,N_23273);
nand U23526 (N_23526,N_23151,N_23000);
xnor U23527 (N_23527,N_23378,N_23499);
or U23528 (N_23528,N_23061,N_23218);
nor U23529 (N_23529,N_23019,N_23145);
nand U23530 (N_23530,N_23188,N_23016);
xor U23531 (N_23531,N_23413,N_23456);
nor U23532 (N_23532,N_23321,N_23379);
or U23533 (N_23533,N_23340,N_23080);
nand U23534 (N_23534,N_23031,N_23056);
nor U23535 (N_23535,N_23149,N_23470);
nor U23536 (N_23536,N_23306,N_23109);
nor U23537 (N_23537,N_23054,N_23114);
or U23538 (N_23538,N_23424,N_23224);
nor U23539 (N_23539,N_23048,N_23195);
nor U23540 (N_23540,N_23337,N_23134);
nor U23541 (N_23541,N_23397,N_23343);
nand U23542 (N_23542,N_23349,N_23041);
and U23543 (N_23543,N_23062,N_23053);
or U23544 (N_23544,N_23227,N_23448);
xnor U23545 (N_23545,N_23003,N_23199);
nand U23546 (N_23546,N_23331,N_23285);
or U23547 (N_23547,N_23263,N_23460);
or U23548 (N_23548,N_23357,N_23493);
xor U23549 (N_23549,N_23169,N_23046);
or U23550 (N_23550,N_23344,N_23127);
or U23551 (N_23551,N_23360,N_23394);
xor U23552 (N_23552,N_23478,N_23216);
and U23553 (N_23553,N_23250,N_23447);
and U23554 (N_23554,N_23490,N_23130);
xor U23555 (N_23555,N_23044,N_23428);
xor U23556 (N_23556,N_23143,N_23027);
and U23557 (N_23557,N_23437,N_23123);
nand U23558 (N_23558,N_23418,N_23459);
and U23559 (N_23559,N_23453,N_23088);
nand U23560 (N_23560,N_23242,N_23029);
nor U23561 (N_23561,N_23259,N_23290);
xnor U23562 (N_23562,N_23255,N_23322);
nand U23563 (N_23563,N_23388,N_23171);
xor U23564 (N_23564,N_23391,N_23495);
xor U23565 (N_23565,N_23262,N_23443);
xor U23566 (N_23566,N_23189,N_23162);
nor U23567 (N_23567,N_23345,N_23398);
and U23568 (N_23568,N_23317,N_23323);
nand U23569 (N_23569,N_23198,N_23332);
nor U23570 (N_23570,N_23417,N_23480);
nand U23571 (N_23571,N_23307,N_23192);
nand U23572 (N_23572,N_23297,N_23082);
and U23573 (N_23573,N_23373,N_23135);
or U23574 (N_23574,N_23485,N_23220);
nor U23575 (N_23575,N_23395,N_23219);
and U23576 (N_23576,N_23254,N_23302);
nand U23577 (N_23577,N_23419,N_23291);
nor U23578 (N_23578,N_23187,N_23416);
or U23579 (N_23579,N_23008,N_23426);
or U23580 (N_23580,N_23217,N_23488);
or U23581 (N_23581,N_23052,N_23445);
or U23582 (N_23582,N_23496,N_23083);
or U23583 (N_23583,N_23444,N_23040);
and U23584 (N_23584,N_23090,N_23409);
and U23585 (N_23585,N_23159,N_23095);
nor U23586 (N_23586,N_23209,N_23351);
or U23587 (N_23587,N_23489,N_23280);
nor U23588 (N_23588,N_23414,N_23361);
nand U23589 (N_23589,N_23022,N_23097);
and U23590 (N_23590,N_23284,N_23181);
nand U23591 (N_23591,N_23288,N_23381);
and U23592 (N_23592,N_23363,N_23115);
or U23593 (N_23593,N_23201,N_23472);
nor U23594 (N_23594,N_23436,N_23461);
nor U23595 (N_23595,N_23304,N_23455);
nand U23596 (N_23596,N_23479,N_23276);
nand U23597 (N_23597,N_23197,N_23205);
nand U23598 (N_23598,N_23320,N_23244);
nor U23599 (N_23599,N_23475,N_23474);
nand U23600 (N_23600,N_23012,N_23477);
or U23601 (N_23601,N_23213,N_23069);
nand U23602 (N_23602,N_23215,N_23150);
and U23603 (N_23603,N_23481,N_23085);
xor U23604 (N_23604,N_23325,N_23487);
xnor U23605 (N_23605,N_23384,N_23408);
or U23606 (N_23606,N_23452,N_23014);
nor U23607 (N_23607,N_23374,N_23491);
nand U23608 (N_23608,N_23043,N_23015);
and U23609 (N_23609,N_23463,N_23066);
xnor U23610 (N_23610,N_23256,N_23333);
and U23611 (N_23611,N_23164,N_23347);
and U23612 (N_23612,N_23393,N_23268);
xor U23613 (N_23613,N_23131,N_23035);
nor U23614 (N_23614,N_23006,N_23081);
or U23615 (N_23615,N_23371,N_23180);
or U23616 (N_23616,N_23110,N_23415);
nand U23617 (N_23617,N_23068,N_23104);
or U23618 (N_23618,N_23241,N_23252);
nor U23619 (N_23619,N_23467,N_23039);
xor U23620 (N_23620,N_23208,N_23070);
nand U23621 (N_23621,N_23342,N_23329);
nand U23622 (N_23622,N_23328,N_23036);
and U23623 (N_23623,N_23042,N_23458);
xor U23624 (N_23624,N_23120,N_23111);
xnor U23625 (N_23625,N_23438,N_23258);
or U23626 (N_23626,N_23231,N_23316);
xor U23627 (N_23627,N_23079,N_23101);
nor U23628 (N_23628,N_23072,N_23196);
xnor U23629 (N_23629,N_23355,N_23002);
nand U23630 (N_23630,N_23153,N_23279);
nor U23631 (N_23631,N_23155,N_23264);
and U23632 (N_23632,N_23133,N_23148);
nor U23633 (N_23633,N_23091,N_23126);
xnor U23634 (N_23634,N_23300,N_23406);
xor U23635 (N_23635,N_23034,N_23486);
and U23636 (N_23636,N_23286,N_23383);
or U23637 (N_23637,N_23138,N_23178);
nand U23638 (N_23638,N_23296,N_23191);
nor U23639 (N_23639,N_23009,N_23064);
nor U23640 (N_23640,N_23007,N_23310);
or U23641 (N_23641,N_23167,N_23075);
and U23642 (N_23642,N_23059,N_23099);
xor U23643 (N_23643,N_23377,N_23170);
xnor U23644 (N_23644,N_23179,N_23336);
or U23645 (N_23645,N_23232,N_23172);
nand U23646 (N_23646,N_23098,N_23060);
nand U23647 (N_23647,N_23190,N_23121);
nor U23648 (N_23648,N_23425,N_23432);
nor U23649 (N_23649,N_23175,N_23089);
or U23650 (N_23650,N_23267,N_23045);
xor U23651 (N_23651,N_23492,N_23117);
or U23652 (N_23652,N_23272,N_23364);
nor U23653 (N_23653,N_23466,N_23354);
and U23654 (N_23654,N_23365,N_23222);
xnor U23655 (N_23655,N_23292,N_23165);
nor U23656 (N_23656,N_23464,N_23237);
nor U23657 (N_23657,N_23338,N_23118);
xnor U23658 (N_23658,N_23225,N_23229);
or U23659 (N_23659,N_23071,N_23405);
nand U23660 (N_23660,N_23346,N_23077);
xnor U23661 (N_23661,N_23058,N_23230);
xor U23662 (N_23662,N_23476,N_23400);
or U23663 (N_23663,N_23411,N_23309);
and U23664 (N_23664,N_23396,N_23261);
nor U23665 (N_23665,N_23113,N_23102);
nor U23666 (N_23666,N_23380,N_23497);
nor U23667 (N_23667,N_23154,N_23334);
nor U23668 (N_23668,N_23142,N_23356);
nand U23669 (N_23669,N_23168,N_23294);
nand U23670 (N_23670,N_23207,N_23087);
and U23671 (N_23671,N_23441,N_23245);
xnor U23672 (N_23672,N_23144,N_23366);
nand U23673 (N_23673,N_23137,N_23092);
nor U23674 (N_23674,N_23185,N_23063);
or U23675 (N_23675,N_23362,N_23112);
and U23676 (N_23676,N_23372,N_23482);
xnor U23677 (N_23677,N_23440,N_23402);
xor U23678 (N_23678,N_23240,N_23236);
nor U23679 (N_23679,N_23370,N_23392);
or U23680 (N_23680,N_23407,N_23269);
or U23681 (N_23681,N_23161,N_23301);
xnor U23682 (N_23682,N_23047,N_23389);
or U23683 (N_23683,N_23132,N_23277);
nor U23684 (N_23684,N_23177,N_23146);
and U23685 (N_23685,N_23318,N_23147);
nand U23686 (N_23686,N_23105,N_23033);
nand U23687 (N_23687,N_23116,N_23157);
nor U23688 (N_23688,N_23353,N_23249);
or U23689 (N_23689,N_23427,N_23139);
and U23690 (N_23690,N_23194,N_23093);
nand U23691 (N_23691,N_23358,N_23100);
or U23692 (N_23692,N_23423,N_23293);
and U23693 (N_23693,N_23339,N_23173);
xnor U23694 (N_23694,N_23011,N_23330);
xnor U23695 (N_23695,N_23375,N_23212);
nor U23696 (N_23696,N_23086,N_23433);
and U23697 (N_23697,N_23128,N_23017);
xor U23698 (N_23698,N_23136,N_23324);
and U23699 (N_23699,N_23369,N_23359);
nand U23700 (N_23700,N_23298,N_23451);
xor U23701 (N_23701,N_23023,N_23401);
and U23702 (N_23702,N_23160,N_23078);
nand U23703 (N_23703,N_23404,N_23430);
xnor U23704 (N_23704,N_23390,N_23107);
nor U23705 (N_23705,N_23004,N_23025);
xor U23706 (N_23706,N_23163,N_23182);
and U23707 (N_23707,N_23238,N_23484);
nand U23708 (N_23708,N_23253,N_23454);
xor U23709 (N_23709,N_23001,N_23122);
nor U23710 (N_23710,N_23326,N_23193);
and U23711 (N_23711,N_23257,N_23096);
nor U23712 (N_23712,N_23278,N_23352);
nor U23713 (N_23713,N_23084,N_23158);
nand U23714 (N_23714,N_23442,N_23223);
xor U23715 (N_23715,N_23176,N_23210);
nand U23716 (N_23716,N_23204,N_23457);
nand U23717 (N_23717,N_23125,N_23471);
or U23718 (N_23718,N_23367,N_23422);
or U23719 (N_23719,N_23465,N_23319);
nand U23720 (N_23720,N_23073,N_23028);
nor U23721 (N_23721,N_23446,N_23141);
nand U23722 (N_23722,N_23308,N_23265);
nand U23723 (N_23723,N_23462,N_23335);
nand U23724 (N_23724,N_23184,N_23021);
nor U23725 (N_23725,N_23473,N_23435);
xor U23726 (N_23726,N_23266,N_23233);
xor U23727 (N_23727,N_23183,N_23108);
or U23728 (N_23728,N_23018,N_23124);
nor U23729 (N_23729,N_23303,N_23403);
and U23730 (N_23730,N_23076,N_23050);
xnor U23731 (N_23731,N_23243,N_23439);
nor U23732 (N_23732,N_23106,N_23420);
and U23733 (N_23733,N_23065,N_23152);
nand U23734 (N_23734,N_23399,N_23055);
and U23735 (N_23735,N_23103,N_23202);
and U23736 (N_23736,N_23311,N_23313);
nand U23737 (N_23737,N_23129,N_23421);
xor U23738 (N_23738,N_23051,N_23260);
nor U23739 (N_23739,N_23386,N_23483);
and U23740 (N_23740,N_23376,N_23010);
xnor U23741 (N_23741,N_23067,N_23431);
xor U23742 (N_23742,N_23037,N_23494);
and U23743 (N_23743,N_23057,N_23283);
nor U23744 (N_23744,N_23248,N_23038);
nand U23745 (N_23745,N_23449,N_23299);
nor U23746 (N_23746,N_23026,N_23074);
and U23747 (N_23747,N_23468,N_23498);
or U23748 (N_23748,N_23049,N_23368);
nor U23749 (N_23749,N_23020,N_23221);
or U23750 (N_23750,N_23358,N_23499);
nand U23751 (N_23751,N_23245,N_23289);
or U23752 (N_23752,N_23121,N_23423);
nand U23753 (N_23753,N_23130,N_23401);
xnor U23754 (N_23754,N_23131,N_23065);
nor U23755 (N_23755,N_23003,N_23445);
nand U23756 (N_23756,N_23290,N_23439);
and U23757 (N_23757,N_23272,N_23170);
nand U23758 (N_23758,N_23043,N_23078);
nor U23759 (N_23759,N_23069,N_23482);
or U23760 (N_23760,N_23071,N_23279);
nor U23761 (N_23761,N_23415,N_23077);
nor U23762 (N_23762,N_23235,N_23104);
or U23763 (N_23763,N_23070,N_23105);
and U23764 (N_23764,N_23192,N_23496);
or U23765 (N_23765,N_23396,N_23001);
and U23766 (N_23766,N_23359,N_23194);
nor U23767 (N_23767,N_23337,N_23420);
nor U23768 (N_23768,N_23071,N_23359);
xor U23769 (N_23769,N_23480,N_23013);
or U23770 (N_23770,N_23076,N_23088);
and U23771 (N_23771,N_23462,N_23093);
nand U23772 (N_23772,N_23324,N_23367);
xnor U23773 (N_23773,N_23259,N_23403);
xnor U23774 (N_23774,N_23462,N_23077);
nand U23775 (N_23775,N_23166,N_23396);
nor U23776 (N_23776,N_23276,N_23284);
and U23777 (N_23777,N_23240,N_23360);
nor U23778 (N_23778,N_23214,N_23449);
nor U23779 (N_23779,N_23156,N_23282);
xnor U23780 (N_23780,N_23192,N_23161);
nor U23781 (N_23781,N_23345,N_23279);
or U23782 (N_23782,N_23329,N_23304);
nand U23783 (N_23783,N_23168,N_23477);
nor U23784 (N_23784,N_23015,N_23280);
and U23785 (N_23785,N_23109,N_23212);
xor U23786 (N_23786,N_23429,N_23067);
xnor U23787 (N_23787,N_23039,N_23423);
xor U23788 (N_23788,N_23290,N_23039);
and U23789 (N_23789,N_23436,N_23154);
or U23790 (N_23790,N_23435,N_23479);
and U23791 (N_23791,N_23159,N_23409);
and U23792 (N_23792,N_23425,N_23238);
nor U23793 (N_23793,N_23190,N_23029);
xor U23794 (N_23794,N_23325,N_23190);
xor U23795 (N_23795,N_23155,N_23495);
nor U23796 (N_23796,N_23216,N_23448);
or U23797 (N_23797,N_23214,N_23240);
nand U23798 (N_23798,N_23179,N_23122);
nor U23799 (N_23799,N_23449,N_23451);
or U23800 (N_23800,N_23198,N_23397);
or U23801 (N_23801,N_23016,N_23490);
xor U23802 (N_23802,N_23059,N_23494);
nand U23803 (N_23803,N_23423,N_23294);
nand U23804 (N_23804,N_23159,N_23240);
nand U23805 (N_23805,N_23390,N_23464);
xor U23806 (N_23806,N_23408,N_23358);
xnor U23807 (N_23807,N_23257,N_23366);
or U23808 (N_23808,N_23448,N_23222);
or U23809 (N_23809,N_23492,N_23274);
nand U23810 (N_23810,N_23079,N_23426);
nand U23811 (N_23811,N_23425,N_23458);
and U23812 (N_23812,N_23409,N_23473);
nand U23813 (N_23813,N_23327,N_23063);
nor U23814 (N_23814,N_23161,N_23265);
xor U23815 (N_23815,N_23345,N_23396);
and U23816 (N_23816,N_23196,N_23272);
xnor U23817 (N_23817,N_23070,N_23274);
nor U23818 (N_23818,N_23370,N_23463);
nor U23819 (N_23819,N_23249,N_23364);
nor U23820 (N_23820,N_23239,N_23091);
nor U23821 (N_23821,N_23454,N_23018);
nor U23822 (N_23822,N_23222,N_23117);
and U23823 (N_23823,N_23093,N_23218);
nand U23824 (N_23824,N_23190,N_23062);
nand U23825 (N_23825,N_23235,N_23222);
nor U23826 (N_23826,N_23232,N_23474);
nand U23827 (N_23827,N_23038,N_23364);
nand U23828 (N_23828,N_23326,N_23069);
nor U23829 (N_23829,N_23188,N_23130);
or U23830 (N_23830,N_23471,N_23415);
nand U23831 (N_23831,N_23086,N_23147);
or U23832 (N_23832,N_23389,N_23011);
nand U23833 (N_23833,N_23347,N_23289);
nor U23834 (N_23834,N_23108,N_23158);
xor U23835 (N_23835,N_23068,N_23284);
nor U23836 (N_23836,N_23125,N_23239);
xnor U23837 (N_23837,N_23001,N_23298);
or U23838 (N_23838,N_23230,N_23140);
or U23839 (N_23839,N_23059,N_23485);
xnor U23840 (N_23840,N_23349,N_23253);
and U23841 (N_23841,N_23039,N_23448);
or U23842 (N_23842,N_23347,N_23048);
nand U23843 (N_23843,N_23182,N_23467);
xnor U23844 (N_23844,N_23004,N_23263);
or U23845 (N_23845,N_23335,N_23361);
or U23846 (N_23846,N_23113,N_23297);
and U23847 (N_23847,N_23044,N_23409);
nand U23848 (N_23848,N_23490,N_23058);
or U23849 (N_23849,N_23421,N_23416);
or U23850 (N_23850,N_23027,N_23445);
nand U23851 (N_23851,N_23269,N_23418);
xor U23852 (N_23852,N_23359,N_23292);
and U23853 (N_23853,N_23088,N_23493);
and U23854 (N_23854,N_23474,N_23306);
and U23855 (N_23855,N_23012,N_23356);
nor U23856 (N_23856,N_23220,N_23373);
nand U23857 (N_23857,N_23415,N_23275);
or U23858 (N_23858,N_23454,N_23218);
and U23859 (N_23859,N_23179,N_23057);
and U23860 (N_23860,N_23274,N_23372);
nand U23861 (N_23861,N_23408,N_23238);
and U23862 (N_23862,N_23328,N_23450);
or U23863 (N_23863,N_23111,N_23034);
nor U23864 (N_23864,N_23062,N_23003);
and U23865 (N_23865,N_23457,N_23331);
nand U23866 (N_23866,N_23010,N_23325);
or U23867 (N_23867,N_23440,N_23478);
nand U23868 (N_23868,N_23456,N_23337);
or U23869 (N_23869,N_23006,N_23023);
nor U23870 (N_23870,N_23301,N_23076);
or U23871 (N_23871,N_23024,N_23065);
or U23872 (N_23872,N_23483,N_23435);
nor U23873 (N_23873,N_23489,N_23241);
nor U23874 (N_23874,N_23003,N_23070);
nand U23875 (N_23875,N_23346,N_23171);
or U23876 (N_23876,N_23346,N_23401);
nand U23877 (N_23877,N_23219,N_23209);
xor U23878 (N_23878,N_23088,N_23212);
nand U23879 (N_23879,N_23373,N_23060);
or U23880 (N_23880,N_23129,N_23477);
nand U23881 (N_23881,N_23064,N_23366);
nand U23882 (N_23882,N_23434,N_23496);
and U23883 (N_23883,N_23195,N_23123);
nand U23884 (N_23884,N_23496,N_23307);
and U23885 (N_23885,N_23199,N_23467);
nor U23886 (N_23886,N_23121,N_23424);
xor U23887 (N_23887,N_23010,N_23174);
nand U23888 (N_23888,N_23017,N_23232);
nand U23889 (N_23889,N_23285,N_23308);
or U23890 (N_23890,N_23273,N_23082);
or U23891 (N_23891,N_23347,N_23031);
or U23892 (N_23892,N_23390,N_23261);
or U23893 (N_23893,N_23324,N_23208);
or U23894 (N_23894,N_23249,N_23075);
xnor U23895 (N_23895,N_23253,N_23259);
xnor U23896 (N_23896,N_23364,N_23459);
or U23897 (N_23897,N_23245,N_23495);
or U23898 (N_23898,N_23479,N_23440);
nand U23899 (N_23899,N_23354,N_23056);
nand U23900 (N_23900,N_23094,N_23151);
and U23901 (N_23901,N_23223,N_23075);
or U23902 (N_23902,N_23414,N_23377);
nand U23903 (N_23903,N_23422,N_23157);
nand U23904 (N_23904,N_23161,N_23014);
and U23905 (N_23905,N_23039,N_23311);
xnor U23906 (N_23906,N_23471,N_23192);
and U23907 (N_23907,N_23343,N_23435);
nor U23908 (N_23908,N_23085,N_23296);
nand U23909 (N_23909,N_23217,N_23284);
nor U23910 (N_23910,N_23328,N_23084);
and U23911 (N_23911,N_23407,N_23087);
or U23912 (N_23912,N_23369,N_23033);
nand U23913 (N_23913,N_23231,N_23456);
xnor U23914 (N_23914,N_23175,N_23016);
or U23915 (N_23915,N_23043,N_23285);
nor U23916 (N_23916,N_23119,N_23194);
and U23917 (N_23917,N_23483,N_23153);
nand U23918 (N_23918,N_23093,N_23054);
and U23919 (N_23919,N_23465,N_23192);
nand U23920 (N_23920,N_23212,N_23282);
nand U23921 (N_23921,N_23409,N_23173);
or U23922 (N_23922,N_23129,N_23151);
and U23923 (N_23923,N_23166,N_23221);
nand U23924 (N_23924,N_23148,N_23324);
xor U23925 (N_23925,N_23474,N_23343);
and U23926 (N_23926,N_23114,N_23372);
nor U23927 (N_23927,N_23004,N_23228);
nor U23928 (N_23928,N_23265,N_23277);
nor U23929 (N_23929,N_23094,N_23399);
nor U23930 (N_23930,N_23095,N_23199);
and U23931 (N_23931,N_23463,N_23100);
xor U23932 (N_23932,N_23155,N_23363);
nand U23933 (N_23933,N_23112,N_23340);
nor U23934 (N_23934,N_23112,N_23358);
nand U23935 (N_23935,N_23130,N_23446);
and U23936 (N_23936,N_23356,N_23372);
nor U23937 (N_23937,N_23022,N_23348);
xnor U23938 (N_23938,N_23428,N_23372);
and U23939 (N_23939,N_23006,N_23285);
xnor U23940 (N_23940,N_23056,N_23421);
nand U23941 (N_23941,N_23471,N_23194);
nand U23942 (N_23942,N_23159,N_23330);
nor U23943 (N_23943,N_23209,N_23119);
xor U23944 (N_23944,N_23449,N_23478);
or U23945 (N_23945,N_23259,N_23194);
xor U23946 (N_23946,N_23060,N_23352);
or U23947 (N_23947,N_23227,N_23188);
nand U23948 (N_23948,N_23493,N_23492);
nor U23949 (N_23949,N_23320,N_23012);
nor U23950 (N_23950,N_23378,N_23481);
or U23951 (N_23951,N_23373,N_23490);
nand U23952 (N_23952,N_23348,N_23180);
or U23953 (N_23953,N_23045,N_23398);
nand U23954 (N_23954,N_23259,N_23378);
nor U23955 (N_23955,N_23069,N_23145);
or U23956 (N_23956,N_23261,N_23187);
nand U23957 (N_23957,N_23461,N_23386);
or U23958 (N_23958,N_23315,N_23012);
nor U23959 (N_23959,N_23438,N_23318);
nand U23960 (N_23960,N_23278,N_23496);
nand U23961 (N_23961,N_23332,N_23197);
nor U23962 (N_23962,N_23332,N_23170);
nand U23963 (N_23963,N_23153,N_23315);
and U23964 (N_23964,N_23175,N_23361);
xor U23965 (N_23965,N_23325,N_23470);
and U23966 (N_23966,N_23308,N_23369);
nand U23967 (N_23967,N_23267,N_23088);
and U23968 (N_23968,N_23141,N_23094);
nand U23969 (N_23969,N_23022,N_23287);
nor U23970 (N_23970,N_23458,N_23241);
nor U23971 (N_23971,N_23388,N_23248);
and U23972 (N_23972,N_23171,N_23464);
nor U23973 (N_23973,N_23150,N_23277);
nand U23974 (N_23974,N_23443,N_23216);
and U23975 (N_23975,N_23151,N_23021);
nor U23976 (N_23976,N_23240,N_23067);
nor U23977 (N_23977,N_23141,N_23189);
nor U23978 (N_23978,N_23251,N_23362);
nor U23979 (N_23979,N_23203,N_23078);
or U23980 (N_23980,N_23254,N_23436);
and U23981 (N_23981,N_23474,N_23491);
nor U23982 (N_23982,N_23085,N_23467);
xor U23983 (N_23983,N_23076,N_23425);
and U23984 (N_23984,N_23041,N_23332);
or U23985 (N_23985,N_23360,N_23085);
nand U23986 (N_23986,N_23110,N_23250);
xnor U23987 (N_23987,N_23278,N_23152);
nand U23988 (N_23988,N_23244,N_23117);
nand U23989 (N_23989,N_23171,N_23140);
xnor U23990 (N_23990,N_23050,N_23477);
nor U23991 (N_23991,N_23326,N_23302);
and U23992 (N_23992,N_23115,N_23193);
xor U23993 (N_23993,N_23191,N_23197);
and U23994 (N_23994,N_23253,N_23416);
or U23995 (N_23995,N_23269,N_23188);
nand U23996 (N_23996,N_23432,N_23164);
and U23997 (N_23997,N_23257,N_23046);
xor U23998 (N_23998,N_23413,N_23291);
nor U23999 (N_23999,N_23173,N_23188);
nand U24000 (N_24000,N_23833,N_23981);
nor U24001 (N_24001,N_23542,N_23653);
and U24002 (N_24002,N_23657,N_23968);
nor U24003 (N_24003,N_23672,N_23610);
xor U24004 (N_24004,N_23975,N_23611);
xnor U24005 (N_24005,N_23540,N_23907);
nor U24006 (N_24006,N_23849,N_23505);
nand U24007 (N_24007,N_23738,N_23888);
xnor U24008 (N_24008,N_23662,N_23659);
xor U24009 (N_24009,N_23520,N_23810);
xor U24010 (N_24010,N_23543,N_23934);
and U24011 (N_24011,N_23623,N_23652);
nand U24012 (N_24012,N_23517,N_23928);
xor U24013 (N_24013,N_23523,N_23963);
nor U24014 (N_24014,N_23946,N_23777);
nand U24015 (N_24015,N_23510,N_23728);
xor U24016 (N_24016,N_23801,N_23622);
nand U24017 (N_24017,N_23614,N_23587);
or U24018 (N_24018,N_23966,N_23685);
or U24019 (N_24019,N_23702,N_23912);
nand U24020 (N_24020,N_23769,N_23950);
and U24021 (N_24021,N_23628,N_23835);
or U24022 (N_24022,N_23739,N_23607);
and U24023 (N_24023,N_23964,N_23765);
or U24024 (N_24024,N_23575,N_23632);
or U24025 (N_24025,N_23629,N_23961);
nand U24026 (N_24026,N_23507,N_23548);
nor U24027 (N_24027,N_23902,N_23973);
nor U24028 (N_24028,N_23819,N_23838);
xor U24029 (N_24029,N_23846,N_23640);
nor U24030 (N_24030,N_23820,N_23861);
nor U24031 (N_24031,N_23803,N_23802);
and U24032 (N_24032,N_23730,N_23696);
xor U24033 (N_24033,N_23567,N_23816);
nand U24034 (N_24034,N_23648,N_23668);
xor U24035 (N_24035,N_23650,N_23641);
and U24036 (N_24036,N_23564,N_23868);
nand U24037 (N_24037,N_23938,N_23895);
nor U24038 (N_24038,N_23954,N_23785);
nor U24039 (N_24039,N_23832,N_23624);
xnor U24040 (N_24040,N_23856,N_23951);
nor U24041 (N_24041,N_23501,N_23549);
and U24042 (N_24042,N_23593,N_23609);
or U24043 (N_24043,N_23615,N_23710);
or U24044 (N_24044,N_23750,N_23527);
and U24045 (N_24045,N_23502,N_23732);
or U24046 (N_24046,N_23790,N_23851);
and U24047 (N_24047,N_23974,N_23508);
or U24048 (N_24048,N_23625,N_23960);
nand U24049 (N_24049,N_23660,N_23736);
and U24050 (N_24050,N_23991,N_23970);
nor U24051 (N_24051,N_23681,N_23559);
xor U24052 (N_24052,N_23636,N_23519);
nand U24053 (N_24053,N_23779,N_23689);
xnor U24054 (N_24054,N_23879,N_23828);
and U24055 (N_24055,N_23642,N_23714);
nor U24056 (N_24056,N_23698,N_23942);
nand U24057 (N_24057,N_23591,N_23724);
and U24058 (N_24058,N_23918,N_23705);
nor U24059 (N_24059,N_23515,N_23677);
nand U24060 (N_24060,N_23890,N_23550);
or U24061 (N_24061,N_23786,N_23663);
nor U24062 (N_24062,N_23500,N_23658);
or U24063 (N_24063,N_23572,N_23757);
nor U24064 (N_24064,N_23733,N_23701);
nand U24065 (N_24065,N_23830,N_23644);
nor U24066 (N_24066,N_23923,N_23682);
nor U24067 (N_24067,N_23583,N_23993);
and U24068 (N_24068,N_23512,N_23612);
xor U24069 (N_24069,N_23751,N_23656);
or U24070 (N_24070,N_23949,N_23541);
nor U24071 (N_24071,N_23772,N_23921);
nor U24072 (N_24072,N_23726,N_23885);
xnor U24073 (N_24073,N_23864,N_23684);
nand U24074 (N_24074,N_23620,N_23744);
and U24075 (N_24075,N_23843,N_23845);
nand U24076 (N_24076,N_23944,N_23742);
and U24077 (N_24077,N_23821,N_23576);
xnor U24078 (N_24078,N_23773,N_23734);
xnor U24079 (N_24079,N_23978,N_23678);
nand U24080 (N_24080,N_23870,N_23852);
xnor U24081 (N_24081,N_23920,N_23827);
nor U24082 (N_24082,N_23878,N_23670);
and U24083 (N_24083,N_23976,N_23909);
nand U24084 (N_24084,N_23539,N_23649);
xnor U24085 (N_24085,N_23651,N_23789);
nand U24086 (N_24086,N_23778,N_23796);
nand U24087 (N_24087,N_23910,N_23797);
xnor U24088 (N_24088,N_23618,N_23834);
or U24089 (N_24089,N_23875,N_23688);
xor U24090 (N_24090,N_23631,N_23933);
and U24091 (N_24091,N_23673,N_23917);
and U24092 (N_24092,N_23967,N_23700);
and U24093 (N_24093,N_23535,N_23638);
nor U24094 (N_24094,N_23997,N_23883);
and U24095 (N_24095,N_23899,N_23807);
or U24096 (N_24096,N_23999,N_23518);
nor U24097 (N_24097,N_23514,N_23661);
nor U24098 (N_24098,N_23774,N_23655);
or U24099 (N_24099,N_23783,N_23882);
and U24100 (N_24100,N_23667,N_23545);
nand U24101 (N_24101,N_23729,N_23504);
or U24102 (N_24102,N_23536,N_23747);
nand U24103 (N_24103,N_23630,N_23871);
xor U24104 (N_24104,N_23980,N_23606);
nand U24105 (N_24105,N_23608,N_23905);
nor U24106 (N_24106,N_23605,N_23647);
or U24107 (N_24107,N_23720,N_23903);
xnor U24108 (N_24108,N_23844,N_23537);
xor U24109 (N_24109,N_23697,N_23692);
nor U24110 (N_24110,N_23853,N_23633);
xnor U24111 (N_24111,N_23958,N_23513);
xnor U24112 (N_24112,N_23586,N_23703);
xnor U24113 (N_24113,N_23741,N_23989);
xnor U24114 (N_24114,N_23753,N_23804);
or U24115 (N_24115,N_23982,N_23809);
xor U24116 (N_24116,N_23617,N_23927);
and U24117 (N_24117,N_23686,N_23516);
nand U24118 (N_24118,N_23597,N_23680);
or U24119 (N_24119,N_23547,N_23743);
nand U24120 (N_24120,N_23908,N_23866);
nand U24121 (N_24121,N_23770,N_23764);
nor U24122 (N_24122,N_23948,N_23916);
xor U24123 (N_24123,N_23780,N_23709);
xor U24124 (N_24124,N_23847,N_23619);
and U24125 (N_24125,N_23836,N_23806);
nor U24126 (N_24126,N_23590,N_23898);
nand U24127 (N_24127,N_23880,N_23596);
and U24128 (N_24128,N_23937,N_23767);
or U24129 (N_24129,N_23665,N_23901);
nor U24130 (N_24130,N_23592,N_23931);
nor U24131 (N_24131,N_23737,N_23755);
nor U24132 (N_24132,N_23745,N_23748);
nor U24133 (N_24133,N_23914,N_23805);
or U24134 (N_24134,N_23683,N_23822);
nor U24135 (N_24135,N_23962,N_23872);
nor U24136 (N_24136,N_23639,N_23791);
nand U24137 (N_24137,N_23892,N_23760);
nor U24138 (N_24138,N_23602,N_23675);
nand U24139 (N_24139,N_23585,N_23857);
nand U24140 (N_24140,N_23771,N_23985);
or U24141 (N_24141,N_23761,N_23599);
nand U24142 (N_24142,N_23578,N_23953);
nand U24143 (N_24143,N_23544,N_23793);
xor U24144 (N_24144,N_23509,N_23595);
nand U24145 (N_24145,N_23528,N_23735);
nand U24146 (N_24146,N_23977,N_23842);
xor U24147 (N_24147,N_23848,N_23525);
xnor U24148 (N_24148,N_23531,N_23850);
xnor U24149 (N_24149,N_23814,N_23725);
xnor U24150 (N_24150,N_23913,N_23529);
xnor U24151 (N_24151,N_23815,N_23635);
or U24152 (N_24152,N_23717,N_23723);
nand U24153 (N_24153,N_23788,N_23972);
nand U24154 (N_24154,N_23818,N_23887);
and U24155 (N_24155,N_23929,N_23759);
xor U24156 (N_24156,N_23756,N_23798);
and U24157 (N_24157,N_23711,N_23707);
nand U24158 (N_24158,N_23915,N_23669);
and U24159 (N_24159,N_23579,N_23654);
nor U24160 (N_24160,N_23671,N_23762);
nand U24161 (N_24161,N_23674,N_23926);
or U24162 (N_24162,N_23746,N_23679);
and U24163 (N_24163,N_23566,N_23922);
nand U24164 (N_24164,N_23781,N_23795);
or U24165 (N_24165,N_23699,N_23987);
or U24166 (N_24166,N_23565,N_23824);
nor U24167 (N_24167,N_23560,N_23896);
xnor U24168 (N_24168,N_23563,N_23580);
nand U24169 (N_24169,N_23693,N_23530);
and U24170 (N_24170,N_23940,N_23616);
or U24171 (N_24171,N_23666,N_23690);
xor U24172 (N_24172,N_23534,N_23643);
and U24173 (N_24173,N_23526,N_23800);
or U24174 (N_24174,N_23932,N_23877);
nor U24175 (N_24175,N_23718,N_23704);
and U24176 (N_24176,N_23936,N_23706);
nand U24177 (N_24177,N_23996,N_23749);
xor U24178 (N_24178,N_23957,N_23553);
or U24179 (N_24179,N_23837,N_23521);
or U24180 (N_24180,N_23584,N_23947);
nand U24181 (N_24181,N_23600,N_23691);
nor U24182 (N_24182,N_23721,N_23854);
nor U24183 (N_24183,N_23716,N_23841);
nand U24184 (N_24184,N_23752,N_23998);
nor U24185 (N_24185,N_23522,N_23984);
xor U24186 (N_24186,N_23867,N_23831);
and U24187 (N_24187,N_23604,N_23823);
and U24188 (N_24188,N_23722,N_23897);
nand U24189 (N_24189,N_23556,N_23740);
and U24190 (N_24190,N_23524,N_23613);
nor U24191 (N_24191,N_23969,N_23826);
nor U24192 (N_24192,N_23876,N_23959);
nand U24193 (N_24193,N_23538,N_23784);
xnor U24194 (N_24194,N_23571,N_23562);
or U24195 (N_24195,N_23945,N_23551);
nor U24196 (N_24196,N_23971,N_23992);
nand U24197 (N_24197,N_23889,N_23603);
and U24198 (N_24198,N_23727,N_23782);
and U24199 (N_24199,N_23988,N_23935);
nor U24200 (N_24200,N_23594,N_23862);
or U24201 (N_24201,N_23646,N_23855);
nor U24202 (N_24202,N_23839,N_23874);
nor U24203 (N_24203,N_23569,N_23808);
xnor U24204 (N_24204,N_23694,N_23695);
and U24205 (N_24205,N_23825,N_23943);
nor U24206 (N_24206,N_23768,N_23995);
xor U24207 (N_24207,N_23811,N_23840);
xor U24208 (N_24208,N_23634,N_23891);
and U24209 (N_24209,N_23930,N_23775);
nor U24210 (N_24210,N_23829,N_23924);
nor U24211 (N_24211,N_23581,N_23794);
nand U24212 (N_24212,N_23965,N_23561);
xor U24213 (N_24213,N_23904,N_23865);
nor U24214 (N_24214,N_23754,N_23506);
and U24215 (N_24215,N_23812,N_23858);
and U24216 (N_24216,N_23952,N_23676);
nand U24217 (N_24217,N_23664,N_23555);
and U24218 (N_24218,N_23637,N_23817);
and U24219 (N_24219,N_23588,N_23546);
and U24220 (N_24220,N_23939,N_23919);
or U24221 (N_24221,N_23573,N_23869);
and U24222 (N_24222,N_23503,N_23713);
nand U24223 (N_24223,N_23574,N_23589);
or U24224 (N_24224,N_23787,N_23533);
nand U24225 (N_24225,N_23863,N_23955);
nand U24226 (N_24226,N_23886,N_23601);
and U24227 (N_24227,N_23554,N_23900);
nor U24228 (N_24228,N_23941,N_23687);
or U24229 (N_24229,N_23621,N_23577);
or U24230 (N_24230,N_23582,N_23994);
nor U24231 (N_24231,N_23708,N_23712);
or U24232 (N_24232,N_23986,N_23715);
nand U24233 (N_24233,N_23532,N_23881);
xor U24234 (N_24234,N_23552,N_23511);
or U24235 (N_24235,N_23557,N_23956);
xor U24236 (N_24236,N_23873,N_23894);
xnor U24237 (N_24237,N_23719,N_23645);
xor U24238 (N_24238,N_23906,N_23990);
xor U24239 (N_24239,N_23893,N_23911);
and U24240 (N_24240,N_23860,N_23570);
or U24241 (N_24241,N_23925,N_23983);
xor U24242 (N_24242,N_23558,N_23776);
or U24243 (N_24243,N_23568,N_23598);
xnor U24244 (N_24244,N_23763,N_23884);
nand U24245 (N_24245,N_23627,N_23766);
xnor U24246 (N_24246,N_23979,N_23731);
nand U24247 (N_24247,N_23813,N_23792);
or U24248 (N_24248,N_23859,N_23626);
nand U24249 (N_24249,N_23758,N_23799);
and U24250 (N_24250,N_23502,N_23664);
and U24251 (N_24251,N_23863,N_23597);
xnor U24252 (N_24252,N_23824,N_23564);
xnor U24253 (N_24253,N_23761,N_23605);
xnor U24254 (N_24254,N_23520,N_23568);
xnor U24255 (N_24255,N_23539,N_23765);
nor U24256 (N_24256,N_23842,N_23674);
xor U24257 (N_24257,N_23633,N_23540);
nor U24258 (N_24258,N_23506,N_23763);
xor U24259 (N_24259,N_23589,N_23918);
or U24260 (N_24260,N_23647,N_23823);
or U24261 (N_24261,N_23732,N_23906);
xnor U24262 (N_24262,N_23600,N_23802);
or U24263 (N_24263,N_23785,N_23998);
nor U24264 (N_24264,N_23802,N_23867);
xnor U24265 (N_24265,N_23560,N_23544);
or U24266 (N_24266,N_23789,N_23851);
xnor U24267 (N_24267,N_23557,N_23600);
or U24268 (N_24268,N_23722,N_23807);
or U24269 (N_24269,N_23671,N_23638);
or U24270 (N_24270,N_23609,N_23611);
nand U24271 (N_24271,N_23622,N_23618);
xnor U24272 (N_24272,N_23612,N_23829);
and U24273 (N_24273,N_23682,N_23500);
nor U24274 (N_24274,N_23762,N_23918);
nor U24275 (N_24275,N_23913,N_23679);
and U24276 (N_24276,N_23810,N_23622);
nor U24277 (N_24277,N_23739,N_23546);
or U24278 (N_24278,N_23749,N_23566);
nor U24279 (N_24279,N_23670,N_23601);
and U24280 (N_24280,N_23500,N_23615);
nand U24281 (N_24281,N_23507,N_23614);
and U24282 (N_24282,N_23790,N_23599);
and U24283 (N_24283,N_23598,N_23994);
or U24284 (N_24284,N_23830,N_23948);
nor U24285 (N_24285,N_23835,N_23856);
nor U24286 (N_24286,N_23731,N_23599);
xnor U24287 (N_24287,N_23968,N_23624);
or U24288 (N_24288,N_23961,N_23887);
or U24289 (N_24289,N_23502,N_23900);
nor U24290 (N_24290,N_23985,N_23637);
nand U24291 (N_24291,N_23598,N_23557);
or U24292 (N_24292,N_23526,N_23507);
nor U24293 (N_24293,N_23845,N_23588);
nand U24294 (N_24294,N_23590,N_23722);
nand U24295 (N_24295,N_23649,N_23760);
and U24296 (N_24296,N_23765,N_23547);
nor U24297 (N_24297,N_23787,N_23558);
nor U24298 (N_24298,N_23616,N_23967);
nand U24299 (N_24299,N_23890,N_23810);
or U24300 (N_24300,N_23702,N_23575);
or U24301 (N_24301,N_23967,N_23999);
or U24302 (N_24302,N_23930,N_23998);
nand U24303 (N_24303,N_23906,N_23577);
xnor U24304 (N_24304,N_23586,N_23713);
or U24305 (N_24305,N_23607,N_23722);
nor U24306 (N_24306,N_23773,N_23745);
nand U24307 (N_24307,N_23722,N_23891);
and U24308 (N_24308,N_23662,N_23519);
and U24309 (N_24309,N_23672,N_23823);
or U24310 (N_24310,N_23733,N_23958);
nor U24311 (N_24311,N_23831,N_23503);
and U24312 (N_24312,N_23629,N_23964);
or U24313 (N_24313,N_23599,N_23826);
nor U24314 (N_24314,N_23833,N_23599);
nand U24315 (N_24315,N_23637,N_23529);
nor U24316 (N_24316,N_23530,N_23682);
nor U24317 (N_24317,N_23848,N_23845);
nor U24318 (N_24318,N_23580,N_23752);
nand U24319 (N_24319,N_23851,N_23685);
nand U24320 (N_24320,N_23795,N_23877);
or U24321 (N_24321,N_23642,N_23926);
or U24322 (N_24322,N_23546,N_23693);
nor U24323 (N_24323,N_23960,N_23620);
nor U24324 (N_24324,N_23782,N_23902);
or U24325 (N_24325,N_23576,N_23924);
or U24326 (N_24326,N_23568,N_23990);
nand U24327 (N_24327,N_23517,N_23584);
and U24328 (N_24328,N_23745,N_23982);
nor U24329 (N_24329,N_23744,N_23734);
xor U24330 (N_24330,N_23908,N_23763);
or U24331 (N_24331,N_23921,N_23872);
nand U24332 (N_24332,N_23747,N_23629);
xor U24333 (N_24333,N_23941,N_23540);
or U24334 (N_24334,N_23584,N_23550);
and U24335 (N_24335,N_23822,N_23818);
and U24336 (N_24336,N_23992,N_23557);
nand U24337 (N_24337,N_23679,N_23889);
or U24338 (N_24338,N_23615,N_23549);
nand U24339 (N_24339,N_23689,N_23949);
nand U24340 (N_24340,N_23762,N_23942);
and U24341 (N_24341,N_23722,N_23975);
nor U24342 (N_24342,N_23503,N_23886);
or U24343 (N_24343,N_23904,N_23786);
xor U24344 (N_24344,N_23566,N_23834);
xnor U24345 (N_24345,N_23918,N_23724);
xnor U24346 (N_24346,N_23629,N_23858);
nand U24347 (N_24347,N_23893,N_23566);
or U24348 (N_24348,N_23777,N_23624);
or U24349 (N_24349,N_23861,N_23519);
nor U24350 (N_24350,N_23567,N_23940);
xnor U24351 (N_24351,N_23794,N_23671);
xor U24352 (N_24352,N_23682,N_23827);
and U24353 (N_24353,N_23935,N_23698);
nor U24354 (N_24354,N_23638,N_23708);
and U24355 (N_24355,N_23914,N_23630);
or U24356 (N_24356,N_23513,N_23916);
nand U24357 (N_24357,N_23647,N_23521);
or U24358 (N_24358,N_23648,N_23820);
nor U24359 (N_24359,N_23590,N_23946);
nor U24360 (N_24360,N_23969,N_23749);
nor U24361 (N_24361,N_23999,N_23651);
nand U24362 (N_24362,N_23921,N_23782);
nor U24363 (N_24363,N_23987,N_23743);
xnor U24364 (N_24364,N_23531,N_23990);
and U24365 (N_24365,N_23610,N_23718);
nand U24366 (N_24366,N_23579,N_23875);
or U24367 (N_24367,N_23985,N_23892);
and U24368 (N_24368,N_23901,N_23948);
and U24369 (N_24369,N_23963,N_23664);
xor U24370 (N_24370,N_23737,N_23580);
and U24371 (N_24371,N_23660,N_23609);
nand U24372 (N_24372,N_23678,N_23744);
nand U24373 (N_24373,N_23520,N_23747);
or U24374 (N_24374,N_23861,N_23919);
xnor U24375 (N_24375,N_23808,N_23737);
nor U24376 (N_24376,N_23919,N_23535);
nand U24377 (N_24377,N_23680,N_23955);
nand U24378 (N_24378,N_23969,N_23588);
and U24379 (N_24379,N_23732,N_23527);
nor U24380 (N_24380,N_23830,N_23875);
nor U24381 (N_24381,N_23801,N_23991);
nand U24382 (N_24382,N_23955,N_23810);
nand U24383 (N_24383,N_23545,N_23525);
or U24384 (N_24384,N_23714,N_23591);
or U24385 (N_24385,N_23826,N_23796);
xnor U24386 (N_24386,N_23669,N_23702);
xor U24387 (N_24387,N_23896,N_23657);
xnor U24388 (N_24388,N_23589,N_23643);
xor U24389 (N_24389,N_23811,N_23762);
or U24390 (N_24390,N_23738,N_23580);
nand U24391 (N_24391,N_23589,N_23709);
or U24392 (N_24392,N_23618,N_23617);
xor U24393 (N_24393,N_23914,N_23931);
xor U24394 (N_24394,N_23565,N_23826);
nand U24395 (N_24395,N_23575,N_23998);
nor U24396 (N_24396,N_23954,N_23709);
or U24397 (N_24397,N_23632,N_23942);
nand U24398 (N_24398,N_23514,N_23865);
nor U24399 (N_24399,N_23789,N_23635);
xnor U24400 (N_24400,N_23676,N_23852);
nor U24401 (N_24401,N_23815,N_23502);
xor U24402 (N_24402,N_23867,N_23950);
nand U24403 (N_24403,N_23650,N_23577);
nand U24404 (N_24404,N_23753,N_23812);
nor U24405 (N_24405,N_23666,N_23552);
nand U24406 (N_24406,N_23915,N_23946);
nand U24407 (N_24407,N_23538,N_23685);
nand U24408 (N_24408,N_23680,N_23915);
xor U24409 (N_24409,N_23629,N_23657);
or U24410 (N_24410,N_23653,N_23903);
nand U24411 (N_24411,N_23549,N_23768);
or U24412 (N_24412,N_23981,N_23830);
nand U24413 (N_24413,N_23705,N_23856);
nand U24414 (N_24414,N_23584,N_23572);
nor U24415 (N_24415,N_23510,N_23906);
or U24416 (N_24416,N_23712,N_23936);
xor U24417 (N_24417,N_23838,N_23967);
and U24418 (N_24418,N_23547,N_23984);
xnor U24419 (N_24419,N_23542,N_23867);
and U24420 (N_24420,N_23630,N_23987);
nor U24421 (N_24421,N_23853,N_23656);
nor U24422 (N_24422,N_23762,N_23852);
and U24423 (N_24423,N_23706,N_23955);
and U24424 (N_24424,N_23953,N_23504);
or U24425 (N_24425,N_23637,N_23643);
or U24426 (N_24426,N_23520,N_23932);
xor U24427 (N_24427,N_23572,N_23579);
or U24428 (N_24428,N_23771,N_23761);
nor U24429 (N_24429,N_23974,N_23933);
nand U24430 (N_24430,N_23918,N_23595);
xor U24431 (N_24431,N_23815,N_23754);
nor U24432 (N_24432,N_23636,N_23838);
nand U24433 (N_24433,N_23603,N_23909);
nor U24434 (N_24434,N_23607,N_23956);
nand U24435 (N_24435,N_23808,N_23870);
xnor U24436 (N_24436,N_23783,N_23875);
and U24437 (N_24437,N_23881,N_23592);
and U24438 (N_24438,N_23805,N_23539);
nor U24439 (N_24439,N_23850,N_23892);
nand U24440 (N_24440,N_23774,N_23548);
nand U24441 (N_24441,N_23501,N_23555);
xor U24442 (N_24442,N_23587,N_23557);
and U24443 (N_24443,N_23690,N_23826);
nand U24444 (N_24444,N_23623,N_23514);
and U24445 (N_24445,N_23503,N_23846);
or U24446 (N_24446,N_23784,N_23514);
and U24447 (N_24447,N_23958,N_23523);
nand U24448 (N_24448,N_23585,N_23575);
nand U24449 (N_24449,N_23996,N_23706);
nor U24450 (N_24450,N_23609,N_23837);
or U24451 (N_24451,N_23893,N_23612);
and U24452 (N_24452,N_23790,N_23840);
and U24453 (N_24453,N_23737,N_23931);
xnor U24454 (N_24454,N_23886,N_23992);
nand U24455 (N_24455,N_23712,N_23782);
and U24456 (N_24456,N_23958,N_23850);
and U24457 (N_24457,N_23598,N_23504);
nor U24458 (N_24458,N_23537,N_23944);
nor U24459 (N_24459,N_23754,N_23669);
nand U24460 (N_24460,N_23562,N_23971);
and U24461 (N_24461,N_23804,N_23846);
and U24462 (N_24462,N_23727,N_23717);
nor U24463 (N_24463,N_23543,N_23897);
or U24464 (N_24464,N_23608,N_23767);
and U24465 (N_24465,N_23799,N_23751);
xor U24466 (N_24466,N_23853,N_23608);
xnor U24467 (N_24467,N_23568,N_23711);
nor U24468 (N_24468,N_23559,N_23659);
nor U24469 (N_24469,N_23782,N_23864);
xnor U24470 (N_24470,N_23873,N_23990);
and U24471 (N_24471,N_23914,N_23696);
nand U24472 (N_24472,N_23991,N_23979);
xor U24473 (N_24473,N_23884,N_23778);
nand U24474 (N_24474,N_23817,N_23614);
and U24475 (N_24475,N_23523,N_23943);
nand U24476 (N_24476,N_23842,N_23604);
and U24477 (N_24477,N_23684,N_23999);
nor U24478 (N_24478,N_23965,N_23662);
nor U24479 (N_24479,N_23901,N_23614);
nand U24480 (N_24480,N_23918,N_23601);
xnor U24481 (N_24481,N_23588,N_23785);
and U24482 (N_24482,N_23537,N_23804);
and U24483 (N_24483,N_23559,N_23747);
nand U24484 (N_24484,N_23931,N_23953);
xnor U24485 (N_24485,N_23925,N_23752);
or U24486 (N_24486,N_23844,N_23781);
and U24487 (N_24487,N_23520,N_23752);
or U24488 (N_24488,N_23696,N_23587);
and U24489 (N_24489,N_23812,N_23987);
or U24490 (N_24490,N_23796,N_23575);
and U24491 (N_24491,N_23818,N_23897);
nand U24492 (N_24492,N_23976,N_23772);
or U24493 (N_24493,N_23664,N_23562);
or U24494 (N_24494,N_23718,N_23719);
and U24495 (N_24495,N_23720,N_23884);
or U24496 (N_24496,N_23994,N_23853);
xor U24497 (N_24497,N_23616,N_23953);
nand U24498 (N_24498,N_23585,N_23611);
nor U24499 (N_24499,N_23693,N_23822);
nor U24500 (N_24500,N_24366,N_24408);
xor U24501 (N_24501,N_24139,N_24039);
and U24502 (N_24502,N_24297,N_24467);
or U24503 (N_24503,N_24225,N_24498);
xor U24504 (N_24504,N_24314,N_24047);
nand U24505 (N_24505,N_24472,N_24245);
and U24506 (N_24506,N_24329,N_24360);
nor U24507 (N_24507,N_24392,N_24443);
xor U24508 (N_24508,N_24198,N_24000);
or U24509 (N_24509,N_24110,N_24174);
or U24510 (N_24510,N_24119,N_24013);
and U24511 (N_24511,N_24418,N_24203);
nand U24512 (N_24512,N_24341,N_24221);
nand U24513 (N_24513,N_24493,N_24098);
or U24514 (N_24514,N_24288,N_24157);
and U24515 (N_24515,N_24061,N_24046);
and U24516 (N_24516,N_24137,N_24099);
or U24517 (N_24517,N_24216,N_24454);
nand U24518 (N_24518,N_24295,N_24227);
or U24519 (N_24519,N_24283,N_24315);
xnor U24520 (N_24520,N_24277,N_24450);
nor U24521 (N_24521,N_24171,N_24217);
and U24522 (N_24522,N_24004,N_24187);
nor U24523 (N_24523,N_24343,N_24199);
xnor U24524 (N_24524,N_24460,N_24263);
nor U24525 (N_24525,N_24079,N_24457);
nand U24526 (N_24526,N_24095,N_24432);
or U24527 (N_24527,N_24275,N_24388);
nand U24528 (N_24528,N_24173,N_24369);
or U24529 (N_24529,N_24016,N_24378);
xor U24530 (N_24530,N_24089,N_24237);
nand U24531 (N_24531,N_24011,N_24224);
nor U24532 (N_24532,N_24147,N_24433);
or U24533 (N_24533,N_24400,N_24232);
nand U24534 (N_24534,N_24105,N_24488);
xnor U24535 (N_24535,N_24351,N_24213);
nand U24536 (N_24536,N_24299,N_24274);
or U24537 (N_24537,N_24131,N_24386);
and U24538 (N_24538,N_24406,N_24186);
nor U24539 (N_24539,N_24322,N_24380);
and U24540 (N_24540,N_24142,N_24358);
and U24541 (N_24541,N_24168,N_24185);
or U24542 (N_24542,N_24037,N_24162);
or U24543 (N_24543,N_24051,N_24086);
and U24544 (N_24544,N_24175,N_24354);
xor U24545 (N_24545,N_24293,N_24482);
nand U24546 (N_24546,N_24278,N_24497);
nor U24547 (N_24547,N_24441,N_24396);
or U24548 (N_24548,N_24024,N_24349);
or U24549 (N_24549,N_24003,N_24012);
nor U24550 (N_24550,N_24133,N_24008);
nor U24551 (N_24551,N_24383,N_24347);
nor U24552 (N_24552,N_24026,N_24280);
nand U24553 (N_24553,N_24149,N_24385);
nor U24554 (N_24554,N_24251,N_24136);
and U24555 (N_24555,N_24429,N_24077);
or U24556 (N_24556,N_24248,N_24097);
and U24557 (N_24557,N_24115,N_24474);
or U24558 (N_24558,N_24442,N_24310);
and U24559 (N_24559,N_24065,N_24238);
nand U24560 (N_24560,N_24464,N_24017);
xnor U24561 (N_24561,N_24144,N_24107);
or U24562 (N_24562,N_24326,N_24453);
nor U24563 (N_24563,N_24269,N_24019);
nand U24564 (N_24564,N_24179,N_24313);
or U24565 (N_24565,N_24090,N_24207);
nor U24566 (N_24566,N_24255,N_24172);
nand U24567 (N_24567,N_24356,N_24328);
nor U24568 (N_24568,N_24291,N_24153);
and U24569 (N_24569,N_24176,N_24338);
xnor U24570 (N_24570,N_24091,N_24438);
or U24571 (N_24571,N_24395,N_24368);
and U24572 (N_24572,N_24375,N_24018);
nand U24573 (N_24573,N_24054,N_24020);
xnor U24574 (N_24574,N_24270,N_24308);
nor U24575 (N_24575,N_24449,N_24169);
nand U24576 (N_24576,N_24468,N_24062);
nand U24577 (N_24577,N_24132,N_24233);
nand U24578 (N_24578,N_24240,N_24182);
and U24579 (N_24579,N_24188,N_24028);
or U24580 (N_24580,N_24276,N_24080);
xnor U24581 (N_24581,N_24066,N_24236);
and U24582 (N_24582,N_24284,N_24499);
and U24583 (N_24583,N_24446,N_24150);
and U24584 (N_24584,N_24140,N_24242);
xor U24585 (N_24585,N_24475,N_24370);
nand U24586 (N_24586,N_24158,N_24264);
and U24587 (N_24587,N_24034,N_24391);
nor U24588 (N_24588,N_24415,N_24009);
nor U24589 (N_24589,N_24440,N_24025);
nor U24590 (N_24590,N_24336,N_24362);
nor U24591 (N_24591,N_24285,N_24102);
nand U24592 (N_24592,N_24160,N_24154);
and U24593 (N_24593,N_24471,N_24231);
nor U24594 (N_24594,N_24466,N_24282);
or U24595 (N_24595,N_24412,N_24112);
and U24596 (N_24596,N_24252,N_24022);
or U24597 (N_24597,N_24307,N_24312);
xnor U24598 (N_24598,N_24404,N_24381);
nand U24599 (N_24599,N_24289,N_24072);
nand U24600 (N_24600,N_24267,N_24123);
nand U24601 (N_24601,N_24407,N_24214);
nand U24602 (N_24602,N_24364,N_24439);
or U24603 (N_24603,N_24296,N_24481);
xor U24604 (N_24604,N_24292,N_24032);
and U24605 (N_24605,N_24320,N_24155);
or U24606 (N_24606,N_24094,N_24294);
xnor U24607 (N_24607,N_24410,N_24036);
nor U24608 (N_24608,N_24228,N_24287);
xor U24609 (N_24609,N_24335,N_24124);
nor U24610 (N_24610,N_24161,N_24060);
or U24611 (N_24611,N_24492,N_24363);
xor U24612 (N_24612,N_24053,N_24071);
nor U24613 (N_24613,N_24042,N_24100);
and U24614 (N_24614,N_24254,N_24040);
or U24615 (N_24615,N_24479,N_24134);
nor U24616 (N_24616,N_24290,N_24428);
nand U24617 (N_24617,N_24201,N_24070);
or U24618 (N_24618,N_24082,N_24266);
nor U24619 (N_24619,N_24048,N_24279);
nand U24620 (N_24620,N_24361,N_24325);
or U24621 (N_24621,N_24330,N_24208);
and U24622 (N_24622,N_24067,N_24226);
or U24623 (N_24623,N_24063,N_24081);
nor U24624 (N_24624,N_24430,N_24350);
xor U24625 (N_24625,N_24235,N_24253);
xnor U24626 (N_24626,N_24166,N_24215);
nand U24627 (N_24627,N_24331,N_24027);
nand U24628 (N_24628,N_24163,N_24480);
nand U24629 (N_24629,N_24035,N_24348);
xor U24630 (N_24630,N_24402,N_24257);
and U24631 (N_24631,N_24222,N_24390);
and U24632 (N_24632,N_24210,N_24318);
nor U24633 (N_24633,N_24050,N_24195);
nor U24634 (N_24634,N_24298,N_24494);
nand U24635 (N_24635,N_24268,N_24411);
xnor U24636 (N_24636,N_24118,N_24319);
nand U24637 (N_24637,N_24445,N_24423);
and U24638 (N_24638,N_24377,N_24359);
or U24639 (N_24639,N_24444,N_24247);
and U24640 (N_24640,N_24333,N_24355);
xor U24641 (N_24641,N_24409,N_24064);
xnor U24642 (N_24642,N_24470,N_24109);
and U24643 (N_24643,N_24374,N_24405);
and U24644 (N_24644,N_24151,N_24164);
nand U24645 (N_24645,N_24473,N_24246);
xnor U24646 (N_24646,N_24401,N_24128);
nand U24647 (N_24647,N_24043,N_24068);
nor U24648 (N_24648,N_24194,N_24431);
or U24649 (N_24649,N_24165,N_24399);
nor U24650 (N_24650,N_24317,N_24321);
and U24651 (N_24651,N_24209,N_24286);
xnor U24652 (N_24652,N_24311,N_24014);
xnor U24653 (N_24653,N_24262,N_24465);
xor U24654 (N_24654,N_24126,N_24414);
nand U24655 (N_24655,N_24376,N_24478);
nand U24656 (N_24656,N_24323,N_24249);
nor U24657 (N_24657,N_24434,N_24244);
or U24658 (N_24658,N_24177,N_24491);
or U24659 (N_24659,N_24337,N_24015);
xnor U24660 (N_24660,N_24145,N_24141);
xnor U24661 (N_24661,N_24167,N_24083);
or U24662 (N_24662,N_24273,N_24074);
nand U24663 (N_24663,N_24223,N_24397);
or U24664 (N_24664,N_24170,N_24239);
xor U24665 (N_24665,N_24243,N_24116);
nand U24666 (N_24666,N_24031,N_24372);
nor U24667 (N_24667,N_24485,N_24200);
nand U24668 (N_24668,N_24357,N_24420);
and U24669 (N_24669,N_24146,N_24041);
and U24670 (N_24670,N_24342,N_24191);
or U24671 (N_24671,N_24353,N_24085);
nor U24672 (N_24672,N_24211,N_24129);
or U24673 (N_24673,N_24258,N_24087);
nand U24674 (N_24674,N_24462,N_24059);
and U24675 (N_24675,N_24271,N_24463);
xor U24676 (N_24676,N_24055,N_24426);
nor U24677 (N_24677,N_24413,N_24135);
nor U24678 (N_24678,N_24044,N_24069);
xnor U24679 (N_24679,N_24490,N_24106);
nand U24680 (N_24680,N_24121,N_24309);
nand U24681 (N_24681,N_24416,N_24180);
and U24682 (N_24682,N_24092,N_24148);
nand U24683 (N_24683,N_24384,N_24345);
and U24684 (N_24684,N_24340,N_24447);
and U24685 (N_24685,N_24265,N_24339);
or U24686 (N_24686,N_24389,N_24049);
and U24687 (N_24687,N_24189,N_24477);
xnor U24688 (N_24688,N_24346,N_24250);
and U24689 (N_24689,N_24058,N_24206);
nor U24690 (N_24690,N_24379,N_24192);
nor U24691 (N_24691,N_24334,N_24403);
xnor U24692 (N_24692,N_24204,N_24256);
and U24693 (N_24693,N_24458,N_24056);
xnor U24694 (N_24694,N_24006,N_24425);
nor U24695 (N_24695,N_24030,N_24156);
nand U24696 (N_24696,N_24108,N_24219);
xor U24697 (N_24697,N_24178,N_24382);
nand U24698 (N_24698,N_24005,N_24371);
nor U24699 (N_24699,N_24114,N_24459);
or U24700 (N_24700,N_24029,N_24367);
nand U24701 (N_24701,N_24394,N_24436);
or U24702 (N_24702,N_24435,N_24205);
and U24703 (N_24703,N_24421,N_24111);
xor U24704 (N_24704,N_24127,N_24489);
or U24705 (N_24705,N_24424,N_24096);
nor U24706 (N_24706,N_24152,N_24487);
nand U24707 (N_24707,N_24352,N_24052);
nor U24708 (N_24708,N_24202,N_24220);
nand U24709 (N_24709,N_24365,N_24218);
nand U24710 (N_24710,N_24300,N_24057);
and U24711 (N_24711,N_24084,N_24130);
nand U24712 (N_24712,N_24007,N_24393);
xor U24713 (N_24713,N_24303,N_24302);
and U24714 (N_24714,N_24033,N_24078);
xnor U24715 (N_24715,N_24045,N_24456);
nand U24716 (N_24716,N_24093,N_24259);
and U24717 (N_24717,N_24104,N_24437);
and U24718 (N_24718,N_24197,N_24196);
xnor U24719 (N_24719,N_24332,N_24373);
nor U24720 (N_24720,N_24143,N_24122);
or U24721 (N_24721,N_24138,N_24101);
xor U24722 (N_24722,N_24234,N_24260);
nand U24723 (N_24723,N_24387,N_24398);
xor U24724 (N_24724,N_24281,N_24261);
and U24725 (N_24725,N_24301,N_24427);
xnor U24726 (N_24726,N_24451,N_24327);
nand U24727 (N_24727,N_24073,N_24183);
nor U24728 (N_24728,N_24076,N_24159);
nor U24729 (N_24729,N_24452,N_24212);
and U24730 (N_24730,N_24469,N_24190);
and U24731 (N_24731,N_24021,N_24113);
and U24732 (N_24732,N_24229,N_24304);
and U24733 (N_24733,N_24422,N_24305);
or U24734 (N_24734,N_24272,N_24419);
or U24735 (N_24735,N_24125,N_24495);
nor U24736 (N_24736,N_24230,N_24184);
xor U24737 (N_24737,N_24324,N_24181);
xnor U24738 (N_24738,N_24075,N_24038);
or U24739 (N_24739,N_24103,N_24344);
nor U24740 (N_24740,N_24193,N_24316);
or U24741 (N_24741,N_24241,N_24461);
and U24742 (N_24742,N_24010,N_24088);
nor U24743 (N_24743,N_24306,N_24120);
nor U24744 (N_24744,N_24496,N_24483);
nand U24745 (N_24745,N_24476,N_24448);
xor U24746 (N_24746,N_24486,N_24023);
and U24747 (N_24747,N_24001,N_24484);
and U24748 (N_24748,N_24117,N_24455);
nand U24749 (N_24749,N_24002,N_24417);
nor U24750 (N_24750,N_24217,N_24195);
and U24751 (N_24751,N_24358,N_24207);
nand U24752 (N_24752,N_24344,N_24489);
nor U24753 (N_24753,N_24225,N_24440);
and U24754 (N_24754,N_24327,N_24191);
and U24755 (N_24755,N_24472,N_24253);
and U24756 (N_24756,N_24273,N_24208);
nor U24757 (N_24757,N_24155,N_24277);
nand U24758 (N_24758,N_24295,N_24363);
nand U24759 (N_24759,N_24327,N_24131);
xor U24760 (N_24760,N_24300,N_24464);
xnor U24761 (N_24761,N_24177,N_24211);
nor U24762 (N_24762,N_24406,N_24000);
and U24763 (N_24763,N_24137,N_24470);
and U24764 (N_24764,N_24393,N_24452);
and U24765 (N_24765,N_24347,N_24200);
and U24766 (N_24766,N_24322,N_24193);
and U24767 (N_24767,N_24420,N_24453);
and U24768 (N_24768,N_24250,N_24183);
or U24769 (N_24769,N_24462,N_24362);
nand U24770 (N_24770,N_24000,N_24362);
xnor U24771 (N_24771,N_24408,N_24189);
or U24772 (N_24772,N_24216,N_24411);
or U24773 (N_24773,N_24297,N_24356);
xnor U24774 (N_24774,N_24229,N_24155);
xor U24775 (N_24775,N_24136,N_24333);
nand U24776 (N_24776,N_24199,N_24379);
xnor U24777 (N_24777,N_24341,N_24412);
nand U24778 (N_24778,N_24212,N_24151);
nand U24779 (N_24779,N_24273,N_24234);
and U24780 (N_24780,N_24215,N_24057);
nand U24781 (N_24781,N_24241,N_24380);
xor U24782 (N_24782,N_24483,N_24360);
nor U24783 (N_24783,N_24134,N_24401);
or U24784 (N_24784,N_24441,N_24245);
xnor U24785 (N_24785,N_24284,N_24304);
or U24786 (N_24786,N_24334,N_24180);
xor U24787 (N_24787,N_24369,N_24092);
nor U24788 (N_24788,N_24252,N_24169);
xor U24789 (N_24789,N_24320,N_24300);
or U24790 (N_24790,N_24224,N_24305);
or U24791 (N_24791,N_24484,N_24111);
or U24792 (N_24792,N_24464,N_24116);
nand U24793 (N_24793,N_24483,N_24026);
xor U24794 (N_24794,N_24143,N_24389);
nor U24795 (N_24795,N_24291,N_24282);
and U24796 (N_24796,N_24307,N_24189);
nand U24797 (N_24797,N_24349,N_24169);
nor U24798 (N_24798,N_24222,N_24077);
or U24799 (N_24799,N_24372,N_24393);
and U24800 (N_24800,N_24353,N_24194);
and U24801 (N_24801,N_24493,N_24367);
xnor U24802 (N_24802,N_24470,N_24454);
nand U24803 (N_24803,N_24467,N_24041);
nand U24804 (N_24804,N_24482,N_24036);
xnor U24805 (N_24805,N_24272,N_24428);
xor U24806 (N_24806,N_24295,N_24315);
and U24807 (N_24807,N_24082,N_24390);
or U24808 (N_24808,N_24399,N_24139);
xor U24809 (N_24809,N_24266,N_24360);
nand U24810 (N_24810,N_24215,N_24430);
xnor U24811 (N_24811,N_24358,N_24091);
and U24812 (N_24812,N_24350,N_24246);
nand U24813 (N_24813,N_24005,N_24200);
nor U24814 (N_24814,N_24140,N_24150);
nor U24815 (N_24815,N_24119,N_24411);
xnor U24816 (N_24816,N_24125,N_24147);
nor U24817 (N_24817,N_24128,N_24297);
or U24818 (N_24818,N_24275,N_24119);
and U24819 (N_24819,N_24287,N_24425);
nor U24820 (N_24820,N_24440,N_24314);
nor U24821 (N_24821,N_24294,N_24171);
xor U24822 (N_24822,N_24455,N_24019);
xor U24823 (N_24823,N_24409,N_24154);
nor U24824 (N_24824,N_24074,N_24054);
and U24825 (N_24825,N_24441,N_24420);
and U24826 (N_24826,N_24427,N_24026);
or U24827 (N_24827,N_24077,N_24376);
nor U24828 (N_24828,N_24262,N_24071);
xor U24829 (N_24829,N_24094,N_24170);
or U24830 (N_24830,N_24135,N_24223);
nand U24831 (N_24831,N_24100,N_24271);
nor U24832 (N_24832,N_24258,N_24244);
and U24833 (N_24833,N_24103,N_24202);
and U24834 (N_24834,N_24175,N_24288);
xor U24835 (N_24835,N_24381,N_24197);
xor U24836 (N_24836,N_24281,N_24240);
nor U24837 (N_24837,N_24273,N_24192);
xnor U24838 (N_24838,N_24157,N_24498);
or U24839 (N_24839,N_24097,N_24235);
xnor U24840 (N_24840,N_24025,N_24039);
and U24841 (N_24841,N_24452,N_24000);
nand U24842 (N_24842,N_24345,N_24413);
nor U24843 (N_24843,N_24170,N_24326);
or U24844 (N_24844,N_24111,N_24446);
nand U24845 (N_24845,N_24232,N_24086);
nor U24846 (N_24846,N_24364,N_24495);
or U24847 (N_24847,N_24196,N_24499);
nand U24848 (N_24848,N_24138,N_24468);
nor U24849 (N_24849,N_24373,N_24483);
xor U24850 (N_24850,N_24168,N_24070);
nor U24851 (N_24851,N_24143,N_24060);
or U24852 (N_24852,N_24429,N_24170);
nor U24853 (N_24853,N_24354,N_24346);
or U24854 (N_24854,N_24388,N_24077);
and U24855 (N_24855,N_24122,N_24488);
nand U24856 (N_24856,N_24300,N_24369);
nor U24857 (N_24857,N_24439,N_24117);
nor U24858 (N_24858,N_24268,N_24321);
or U24859 (N_24859,N_24357,N_24080);
xor U24860 (N_24860,N_24400,N_24494);
nand U24861 (N_24861,N_24492,N_24190);
xor U24862 (N_24862,N_24142,N_24070);
nor U24863 (N_24863,N_24145,N_24074);
nor U24864 (N_24864,N_24250,N_24222);
nand U24865 (N_24865,N_24198,N_24024);
nand U24866 (N_24866,N_24399,N_24354);
or U24867 (N_24867,N_24292,N_24141);
xor U24868 (N_24868,N_24185,N_24295);
nor U24869 (N_24869,N_24350,N_24238);
nand U24870 (N_24870,N_24449,N_24399);
nor U24871 (N_24871,N_24027,N_24214);
nand U24872 (N_24872,N_24043,N_24477);
nor U24873 (N_24873,N_24433,N_24093);
and U24874 (N_24874,N_24466,N_24021);
xnor U24875 (N_24875,N_24159,N_24158);
nor U24876 (N_24876,N_24206,N_24143);
xor U24877 (N_24877,N_24468,N_24221);
xnor U24878 (N_24878,N_24212,N_24486);
and U24879 (N_24879,N_24422,N_24402);
nor U24880 (N_24880,N_24493,N_24309);
or U24881 (N_24881,N_24044,N_24379);
or U24882 (N_24882,N_24234,N_24117);
and U24883 (N_24883,N_24486,N_24358);
and U24884 (N_24884,N_24467,N_24364);
and U24885 (N_24885,N_24095,N_24368);
nor U24886 (N_24886,N_24150,N_24025);
and U24887 (N_24887,N_24047,N_24378);
xnor U24888 (N_24888,N_24399,N_24105);
and U24889 (N_24889,N_24105,N_24375);
nand U24890 (N_24890,N_24374,N_24240);
or U24891 (N_24891,N_24182,N_24161);
or U24892 (N_24892,N_24048,N_24342);
and U24893 (N_24893,N_24115,N_24025);
xor U24894 (N_24894,N_24483,N_24103);
nor U24895 (N_24895,N_24388,N_24399);
nand U24896 (N_24896,N_24108,N_24367);
nor U24897 (N_24897,N_24279,N_24261);
xnor U24898 (N_24898,N_24388,N_24125);
and U24899 (N_24899,N_24070,N_24154);
and U24900 (N_24900,N_24005,N_24396);
or U24901 (N_24901,N_24277,N_24337);
and U24902 (N_24902,N_24171,N_24451);
or U24903 (N_24903,N_24017,N_24030);
nand U24904 (N_24904,N_24060,N_24014);
nor U24905 (N_24905,N_24127,N_24219);
and U24906 (N_24906,N_24415,N_24400);
xor U24907 (N_24907,N_24324,N_24414);
and U24908 (N_24908,N_24453,N_24117);
xor U24909 (N_24909,N_24118,N_24033);
xnor U24910 (N_24910,N_24132,N_24093);
nand U24911 (N_24911,N_24441,N_24041);
and U24912 (N_24912,N_24079,N_24023);
nand U24913 (N_24913,N_24370,N_24421);
nand U24914 (N_24914,N_24359,N_24252);
nand U24915 (N_24915,N_24423,N_24224);
nand U24916 (N_24916,N_24254,N_24168);
or U24917 (N_24917,N_24022,N_24320);
nor U24918 (N_24918,N_24009,N_24411);
or U24919 (N_24919,N_24292,N_24348);
nor U24920 (N_24920,N_24378,N_24202);
and U24921 (N_24921,N_24432,N_24223);
xnor U24922 (N_24922,N_24481,N_24429);
nor U24923 (N_24923,N_24239,N_24353);
and U24924 (N_24924,N_24351,N_24293);
and U24925 (N_24925,N_24075,N_24071);
nand U24926 (N_24926,N_24112,N_24396);
or U24927 (N_24927,N_24295,N_24455);
nor U24928 (N_24928,N_24498,N_24286);
or U24929 (N_24929,N_24472,N_24143);
nor U24930 (N_24930,N_24260,N_24139);
xnor U24931 (N_24931,N_24486,N_24060);
or U24932 (N_24932,N_24112,N_24416);
nor U24933 (N_24933,N_24458,N_24150);
or U24934 (N_24934,N_24223,N_24029);
nand U24935 (N_24935,N_24299,N_24085);
nand U24936 (N_24936,N_24441,N_24027);
nor U24937 (N_24937,N_24138,N_24068);
and U24938 (N_24938,N_24336,N_24409);
nand U24939 (N_24939,N_24032,N_24030);
and U24940 (N_24940,N_24183,N_24430);
and U24941 (N_24941,N_24291,N_24287);
xnor U24942 (N_24942,N_24093,N_24381);
nor U24943 (N_24943,N_24083,N_24062);
xor U24944 (N_24944,N_24134,N_24136);
and U24945 (N_24945,N_24383,N_24354);
nor U24946 (N_24946,N_24286,N_24446);
xor U24947 (N_24947,N_24387,N_24040);
nand U24948 (N_24948,N_24164,N_24047);
and U24949 (N_24949,N_24069,N_24400);
nand U24950 (N_24950,N_24323,N_24172);
and U24951 (N_24951,N_24413,N_24218);
nor U24952 (N_24952,N_24174,N_24033);
xnor U24953 (N_24953,N_24241,N_24395);
or U24954 (N_24954,N_24495,N_24006);
xor U24955 (N_24955,N_24348,N_24121);
xnor U24956 (N_24956,N_24167,N_24398);
xor U24957 (N_24957,N_24191,N_24019);
or U24958 (N_24958,N_24384,N_24013);
xor U24959 (N_24959,N_24477,N_24491);
nand U24960 (N_24960,N_24466,N_24109);
nand U24961 (N_24961,N_24121,N_24305);
and U24962 (N_24962,N_24351,N_24445);
nor U24963 (N_24963,N_24456,N_24132);
or U24964 (N_24964,N_24093,N_24434);
nor U24965 (N_24965,N_24363,N_24419);
nand U24966 (N_24966,N_24244,N_24279);
nand U24967 (N_24967,N_24471,N_24303);
nand U24968 (N_24968,N_24091,N_24173);
nor U24969 (N_24969,N_24002,N_24135);
nand U24970 (N_24970,N_24175,N_24326);
nand U24971 (N_24971,N_24054,N_24346);
or U24972 (N_24972,N_24020,N_24133);
and U24973 (N_24973,N_24228,N_24257);
and U24974 (N_24974,N_24241,N_24454);
nand U24975 (N_24975,N_24112,N_24274);
nand U24976 (N_24976,N_24375,N_24337);
xor U24977 (N_24977,N_24460,N_24375);
and U24978 (N_24978,N_24491,N_24423);
nand U24979 (N_24979,N_24112,N_24430);
and U24980 (N_24980,N_24068,N_24321);
xnor U24981 (N_24981,N_24208,N_24298);
and U24982 (N_24982,N_24346,N_24025);
xnor U24983 (N_24983,N_24083,N_24054);
or U24984 (N_24984,N_24124,N_24346);
or U24985 (N_24985,N_24338,N_24123);
and U24986 (N_24986,N_24150,N_24417);
nor U24987 (N_24987,N_24342,N_24087);
nand U24988 (N_24988,N_24397,N_24164);
nor U24989 (N_24989,N_24114,N_24212);
and U24990 (N_24990,N_24325,N_24238);
nor U24991 (N_24991,N_24185,N_24105);
or U24992 (N_24992,N_24106,N_24456);
xnor U24993 (N_24993,N_24178,N_24188);
or U24994 (N_24994,N_24487,N_24280);
nor U24995 (N_24995,N_24252,N_24155);
and U24996 (N_24996,N_24468,N_24380);
and U24997 (N_24997,N_24104,N_24340);
nand U24998 (N_24998,N_24468,N_24323);
xnor U24999 (N_24999,N_24035,N_24140);
or UO_0 (O_0,N_24882,N_24853);
xor UO_1 (O_1,N_24833,N_24883);
xnor UO_2 (O_2,N_24861,N_24566);
xor UO_3 (O_3,N_24845,N_24571);
xnor UO_4 (O_4,N_24758,N_24790);
nand UO_5 (O_5,N_24534,N_24786);
or UO_6 (O_6,N_24726,N_24843);
or UO_7 (O_7,N_24747,N_24776);
xor UO_8 (O_8,N_24946,N_24909);
and UO_9 (O_9,N_24701,N_24766);
nor UO_10 (O_10,N_24818,N_24742);
and UO_11 (O_11,N_24675,N_24737);
nand UO_12 (O_12,N_24616,N_24892);
xnor UO_13 (O_13,N_24867,N_24588);
xor UO_14 (O_14,N_24983,N_24784);
or UO_15 (O_15,N_24942,N_24510);
and UO_16 (O_16,N_24695,N_24585);
nor UO_17 (O_17,N_24556,N_24968);
xnor UO_18 (O_18,N_24783,N_24810);
nor UO_19 (O_19,N_24609,N_24565);
nand UO_20 (O_20,N_24604,N_24620);
or UO_21 (O_21,N_24512,N_24836);
or UO_22 (O_22,N_24638,N_24956);
xnor UO_23 (O_23,N_24513,N_24605);
xor UO_24 (O_24,N_24598,N_24580);
or UO_25 (O_25,N_24645,N_24660);
or UO_26 (O_26,N_24986,N_24944);
nand UO_27 (O_27,N_24862,N_24553);
nand UO_28 (O_28,N_24622,N_24817);
and UO_29 (O_29,N_24757,N_24506);
xnor UO_30 (O_30,N_24997,N_24540);
nand UO_31 (O_31,N_24576,N_24981);
xnor UO_32 (O_32,N_24811,N_24641);
nand UO_33 (O_33,N_24739,N_24711);
or UO_34 (O_34,N_24750,N_24708);
nand UO_35 (O_35,N_24606,N_24679);
nand UO_36 (O_36,N_24802,N_24754);
or UO_37 (O_37,N_24971,N_24644);
nor UO_38 (O_38,N_24772,N_24600);
nand UO_39 (O_39,N_24940,N_24718);
or UO_40 (O_40,N_24891,N_24799);
and UO_41 (O_41,N_24612,N_24814);
and UO_42 (O_42,N_24508,N_24652);
and UO_43 (O_43,N_24621,N_24929);
or UO_44 (O_44,N_24943,N_24670);
or UO_45 (O_45,N_24805,N_24846);
nor UO_46 (O_46,N_24524,N_24694);
nor UO_47 (O_47,N_24586,N_24584);
nor UO_48 (O_48,N_24686,N_24906);
xnor UO_49 (O_49,N_24979,N_24521);
nand UO_50 (O_50,N_24869,N_24775);
or UO_51 (O_51,N_24541,N_24561);
and UO_52 (O_52,N_24982,N_24728);
and UO_53 (O_53,N_24536,N_24665);
xor UO_54 (O_54,N_24629,N_24590);
or UO_55 (O_55,N_24567,N_24730);
and UO_56 (O_56,N_24927,N_24721);
or UO_57 (O_57,N_24562,N_24939);
nor UO_58 (O_58,N_24889,N_24949);
xor UO_59 (O_59,N_24879,N_24859);
or UO_60 (O_60,N_24624,N_24785);
xor UO_61 (O_61,N_24819,N_24863);
nand UO_62 (O_62,N_24597,N_24875);
nor UO_63 (O_63,N_24911,N_24537);
xnor UO_64 (O_64,N_24976,N_24920);
or UO_65 (O_65,N_24837,N_24503);
xor UO_66 (O_66,N_24528,N_24959);
nand UO_67 (O_67,N_24934,N_24895);
xor UO_68 (O_68,N_24936,N_24907);
nor UO_69 (O_69,N_24668,N_24995);
or UO_70 (O_70,N_24866,N_24778);
or UO_71 (O_71,N_24885,N_24824);
or UO_72 (O_72,N_24633,N_24681);
and UO_73 (O_73,N_24820,N_24674);
nor UO_74 (O_74,N_24991,N_24926);
xor UO_75 (O_75,N_24630,N_24552);
or UO_76 (O_76,N_24878,N_24813);
and UO_77 (O_77,N_24910,N_24768);
and UO_78 (O_78,N_24841,N_24693);
and UO_79 (O_79,N_24842,N_24957);
and UO_80 (O_80,N_24557,N_24676);
nand UO_81 (O_81,N_24706,N_24860);
and UO_82 (O_82,N_24608,N_24801);
xnor UO_83 (O_83,N_24912,N_24579);
nand UO_84 (O_84,N_24509,N_24847);
xor UO_85 (O_85,N_24713,N_24854);
or UO_86 (O_86,N_24852,N_24558);
and UO_87 (O_87,N_24947,N_24962);
nand UO_88 (O_88,N_24890,N_24559);
nor UO_89 (O_89,N_24529,N_24539);
or UO_90 (O_90,N_24734,N_24984);
nand UO_91 (O_91,N_24764,N_24823);
xor UO_92 (O_92,N_24632,N_24526);
or UO_93 (O_93,N_24953,N_24733);
xnor UO_94 (O_94,N_24888,N_24967);
or UO_95 (O_95,N_24932,N_24827);
xor UO_96 (O_96,N_24914,N_24654);
and UO_97 (O_97,N_24748,N_24667);
and UO_98 (O_98,N_24871,N_24699);
xnor UO_99 (O_99,N_24792,N_24725);
xor UO_100 (O_100,N_24542,N_24573);
nand UO_101 (O_101,N_24723,N_24808);
and UO_102 (O_102,N_24753,N_24951);
nand UO_103 (O_103,N_24518,N_24822);
and UO_104 (O_104,N_24602,N_24856);
xnor UO_105 (O_105,N_24704,N_24840);
or UO_106 (O_106,N_24803,N_24627);
nor UO_107 (O_107,N_24500,N_24678);
nor UO_108 (O_108,N_24731,N_24831);
or UO_109 (O_109,N_24649,N_24990);
or UO_110 (O_110,N_24570,N_24514);
or UO_111 (O_111,N_24712,N_24583);
and UO_112 (O_112,N_24653,N_24844);
nand UO_113 (O_113,N_24501,N_24886);
and UO_114 (O_114,N_24687,N_24596);
and UO_115 (O_115,N_24999,N_24809);
and UO_116 (O_116,N_24568,N_24646);
nand UO_117 (O_117,N_24851,N_24918);
and UO_118 (O_118,N_24774,N_24782);
xnor UO_119 (O_119,N_24825,N_24787);
nor UO_120 (O_120,N_24755,N_24582);
xnor UO_121 (O_121,N_24515,N_24680);
or UO_122 (O_122,N_24777,N_24835);
xor UO_123 (O_123,N_24575,N_24732);
nor UO_124 (O_124,N_24672,N_24952);
and UO_125 (O_125,N_24839,N_24752);
nand UO_126 (O_126,N_24830,N_24549);
or UO_127 (O_127,N_24517,N_24963);
nand UO_128 (O_128,N_24950,N_24751);
nor UO_129 (O_129,N_24560,N_24707);
or UO_130 (O_130,N_24794,N_24905);
or UO_131 (O_131,N_24966,N_24611);
nor UO_132 (O_132,N_24922,N_24796);
xor UO_133 (O_133,N_24715,N_24525);
xnor UO_134 (O_134,N_24975,N_24930);
nor UO_135 (O_135,N_24662,N_24759);
or UO_136 (O_136,N_24780,N_24603);
nor UO_137 (O_137,N_24625,N_24736);
nand UO_138 (O_138,N_24650,N_24996);
nor UO_139 (O_139,N_24682,N_24807);
or UO_140 (O_140,N_24789,N_24614);
and UO_141 (O_141,N_24970,N_24639);
xnor UO_142 (O_142,N_24569,N_24896);
nand UO_143 (O_143,N_24887,N_24761);
or UO_144 (O_144,N_24941,N_24893);
or UO_145 (O_145,N_24900,N_24945);
nand UO_146 (O_146,N_24987,N_24505);
or UO_147 (O_147,N_24993,N_24709);
or UO_148 (O_148,N_24700,N_24716);
xnor UO_149 (O_149,N_24877,N_24874);
or UO_150 (O_150,N_24741,N_24925);
xor UO_151 (O_151,N_24684,N_24661);
or UO_152 (O_152,N_24659,N_24587);
nor UO_153 (O_153,N_24791,N_24714);
nor UO_154 (O_154,N_24973,N_24550);
xor UO_155 (O_155,N_24771,N_24743);
and UO_156 (O_156,N_24938,N_24548);
nor UO_157 (O_157,N_24692,N_24593);
xnor UO_158 (O_158,N_24523,N_24601);
or UO_159 (O_159,N_24880,N_24677);
and UO_160 (O_160,N_24520,N_24812);
or UO_161 (O_161,N_24535,N_24720);
nand UO_162 (O_162,N_24815,N_24821);
or UO_163 (O_163,N_24980,N_24648);
and UO_164 (O_164,N_24904,N_24798);
xor UO_165 (O_165,N_24795,N_24502);
nand UO_166 (O_166,N_24637,N_24858);
and UO_167 (O_167,N_24873,N_24994);
nand UO_168 (O_168,N_24705,N_24848);
and UO_169 (O_169,N_24933,N_24989);
and UO_170 (O_170,N_24804,N_24635);
nand UO_171 (O_171,N_24702,N_24921);
xnor UO_172 (O_172,N_24626,N_24738);
or UO_173 (O_173,N_24954,N_24769);
and UO_174 (O_174,N_24685,N_24903);
xnor UO_175 (O_175,N_24770,N_24985);
or UO_176 (O_176,N_24865,N_24507);
nor UO_177 (O_177,N_24763,N_24688);
and UO_178 (O_178,N_24901,N_24746);
and UO_179 (O_179,N_24663,N_24683);
xor UO_180 (O_180,N_24894,N_24577);
nor UO_181 (O_181,N_24960,N_24533);
and UO_182 (O_182,N_24913,N_24978);
nand UO_183 (O_183,N_24710,N_24998);
xnor UO_184 (O_184,N_24828,N_24855);
nor UO_185 (O_185,N_24618,N_24592);
and UO_186 (O_186,N_24511,N_24977);
and UO_187 (O_187,N_24628,N_24749);
or UO_188 (O_188,N_24897,N_24826);
nand UO_189 (O_189,N_24972,N_24689);
or UO_190 (O_190,N_24669,N_24902);
nor UO_191 (O_191,N_24727,N_24574);
nand UO_192 (O_192,N_24703,N_24555);
or UO_193 (O_193,N_24834,N_24642);
nand UO_194 (O_194,N_24781,N_24864);
xnor UO_195 (O_195,N_24613,N_24756);
and UO_196 (O_196,N_24546,N_24961);
xor UO_197 (O_197,N_24779,N_24647);
and UO_198 (O_198,N_24717,N_24631);
nand UO_199 (O_199,N_24916,N_24988);
nand UO_200 (O_200,N_24800,N_24917);
nor UO_201 (O_201,N_24543,N_24767);
nand UO_202 (O_202,N_24623,N_24581);
xor UO_203 (O_203,N_24838,N_24617);
nand UO_204 (O_204,N_24530,N_24564);
and UO_205 (O_205,N_24931,N_24698);
nand UO_206 (O_206,N_24958,N_24881);
or UO_207 (O_207,N_24857,N_24696);
xor UO_208 (O_208,N_24643,N_24610);
xor UO_209 (O_209,N_24634,N_24547);
nand UO_210 (O_210,N_24589,N_24671);
nand UO_211 (O_211,N_24832,N_24992);
xnor UO_212 (O_212,N_24544,N_24527);
xor UO_213 (O_213,N_24765,N_24591);
and UO_214 (O_214,N_24563,N_24948);
nor UO_215 (O_215,N_24788,N_24816);
xor UO_216 (O_216,N_24908,N_24915);
and UO_217 (O_217,N_24658,N_24724);
nor UO_218 (O_218,N_24773,N_24884);
or UO_219 (O_219,N_24762,N_24554);
nand UO_220 (O_220,N_24745,N_24923);
and UO_221 (O_221,N_24640,N_24924);
nand UO_222 (O_222,N_24969,N_24868);
xor UO_223 (O_223,N_24964,N_24532);
and UO_224 (O_224,N_24522,N_24551);
and UO_225 (O_225,N_24666,N_24729);
xnor UO_226 (O_226,N_24872,N_24657);
xor UO_227 (O_227,N_24673,N_24607);
xnor UO_228 (O_228,N_24850,N_24516);
or UO_229 (O_229,N_24919,N_24935);
nand UO_230 (O_230,N_24870,N_24735);
xnor UO_231 (O_231,N_24545,N_24619);
and UO_232 (O_232,N_24690,N_24876);
nand UO_233 (O_233,N_24636,N_24719);
or UO_234 (O_234,N_24928,N_24697);
nor UO_235 (O_235,N_24974,N_24797);
and UO_236 (O_236,N_24655,N_24531);
and UO_237 (O_237,N_24955,N_24594);
nor UO_238 (O_238,N_24849,N_24651);
or UO_239 (O_239,N_24898,N_24760);
nand UO_240 (O_240,N_24965,N_24578);
or UO_241 (O_241,N_24664,N_24829);
and UO_242 (O_242,N_24722,N_24656);
and UO_243 (O_243,N_24691,N_24538);
and UO_244 (O_244,N_24595,N_24806);
nand UO_245 (O_245,N_24744,N_24899);
and UO_246 (O_246,N_24740,N_24504);
nor UO_247 (O_247,N_24793,N_24572);
xnor UO_248 (O_248,N_24599,N_24937);
nor UO_249 (O_249,N_24519,N_24615);
nand UO_250 (O_250,N_24727,N_24747);
nor UO_251 (O_251,N_24907,N_24997);
and UO_252 (O_252,N_24511,N_24519);
and UO_253 (O_253,N_24835,N_24718);
xor UO_254 (O_254,N_24684,N_24520);
and UO_255 (O_255,N_24608,N_24947);
nand UO_256 (O_256,N_24606,N_24928);
xor UO_257 (O_257,N_24779,N_24583);
nor UO_258 (O_258,N_24558,N_24784);
or UO_259 (O_259,N_24936,N_24805);
xor UO_260 (O_260,N_24573,N_24719);
or UO_261 (O_261,N_24527,N_24526);
and UO_262 (O_262,N_24692,N_24816);
nand UO_263 (O_263,N_24952,N_24947);
and UO_264 (O_264,N_24595,N_24752);
or UO_265 (O_265,N_24591,N_24561);
nand UO_266 (O_266,N_24846,N_24989);
nor UO_267 (O_267,N_24888,N_24878);
and UO_268 (O_268,N_24783,N_24620);
and UO_269 (O_269,N_24587,N_24529);
or UO_270 (O_270,N_24626,N_24901);
and UO_271 (O_271,N_24675,N_24704);
nand UO_272 (O_272,N_24643,N_24940);
xnor UO_273 (O_273,N_24613,N_24702);
nand UO_274 (O_274,N_24646,N_24971);
nand UO_275 (O_275,N_24512,N_24993);
or UO_276 (O_276,N_24824,N_24925);
nor UO_277 (O_277,N_24865,N_24649);
and UO_278 (O_278,N_24727,N_24807);
nand UO_279 (O_279,N_24800,N_24629);
xor UO_280 (O_280,N_24688,N_24792);
xor UO_281 (O_281,N_24904,N_24679);
and UO_282 (O_282,N_24535,N_24804);
nor UO_283 (O_283,N_24820,N_24500);
nor UO_284 (O_284,N_24698,N_24505);
nand UO_285 (O_285,N_24606,N_24738);
and UO_286 (O_286,N_24608,N_24992);
or UO_287 (O_287,N_24910,N_24820);
xnor UO_288 (O_288,N_24938,N_24714);
and UO_289 (O_289,N_24841,N_24740);
and UO_290 (O_290,N_24551,N_24590);
nor UO_291 (O_291,N_24746,N_24671);
or UO_292 (O_292,N_24684,N_24560);
nor UO_293 (O_293,N_24749,N_24889);
nor UO_294 (O_294,N_24669,N_24501);
and UO_295 (O_295,N_24624,N_24802);
and UO_296 (O_296,N_24965,N_24649);
xor UO_297 (O_297,N_24913,N_24862);
or UO_298 (O_298,N_24553,N_24569);
nor UO_299 (O_299,N_24657,N_24914);
xor UO_300 (O_300,N_24849,N_24988);
nand UO_301 (O_301,N_24904,N_24718);
xnor UO_302 (O_302,N_24903,N_24662);
and UO_303 (O_303,N_24778,N_24503);
or UO_304 (O_304,N_24517,N_24821);
nor UO_305 (O_305,N_24529,N_24971);
or UO_306 (O_306,N_24757,N_24647);
nand UO_307 (O_307,N_24914,N_24864);
nand UO_308 (O_308,N_24540,N_24672);
and UO_309 (O_309,N_24837,N_24734);
and UO_310 (O_310,N_24769,N_24643);
nor UO_311 (O_311,N_24542,N_24868);
xor UO_312 (O_312,N_24795,N_24569);
and UO_313 (O_313,N_24529,N_24533);
xnor UO_314 (O_314,N_24953,N_24537);
xor UO_315 (O_315,N_24809,N_24609);
nor UO_316 (O_316,N_24882,N_24876);
or UO_317 (O_317,N_24726,N_24856);
or UO_318 (O_318,N_24575,N_24981);
xnor UO_319 (O_319,N_24745,N_24592);
nor UO_320 (O_320,N_24914,N_24688);
xor UO_321 (O_321,N_24660,N_24776);
or UO_322 (O_322,N_24723,N_24719);
nor UO_323 (O_323,N_24831,N_24936);
xnor UO_324 (O_324,N_24532,N_24739);
nand UO_325 (O_325,N_24991,N_24732);
nor UO_326 (O_326,N_24578,N_24593);
nand UO_327 (O_327,N_24605,N_24827);
xor UO_328 (O_328,N_24678,N_24875);
xnor UO_329 (O_329,N_24949,N_24716);
nand UO_330 (O_330,N_24952,N_24845);
or UO_331 (O_331,N_24777,N_24938);
xnor UO_332 (O_332,N_24570,N_24636);
xnor UO_333 (O_333,N_24583,N_24756);
nor UO_334 (O_334,N_24880,N_24968);
and UO_335 (O_335,N_24827,N_24666);
nor UO_336 (O_336,N_24845,N_24806);
nor UO_337 (O_337,N_24551,N_24610);
and UO_338 (O_338,N_24957,N_24818);
and UO_339 (O_339,N_24577,N_24640);
and UO_340 (O_340,N_24734,N_24888);
nand UO_341 (O_341,N_24883,N_24547);
or UO_342 (O_342,N_24954,N_24574);
nand UO_343 (O_343,N_24784,N_24665);
or UO_344 (O_344,N_24761,N_24808);
and UO_345 (O_345,N_24726,N_24773);
or UO_346 (O_346,N_24765,N_24915);
xnor UO_347 (O_347,N_24794,N_24834);
or UO_348 (O_348,N_24792,N_24647);
xnor UO_349 (O_349,N_24603,N_24748);
or UO_350 (O_350,N_24982,N_24736);
xnor UO_351 (O_351,N_24512,N_24734);
or UO_352 (O_352,N_24907,N_24974);
or UO_353 (O_353,N_24561,N_24510);
nand UO_354 (O_354,N_24665,N_24848);
xnor UO_355 (O_355,N_24676,N_24970);
xnor UO_356 (O_356,N_24575,N_24978);
nor UO_357 (O_357,N_24757,N_24586);
nor UO_358 (O_358,N_24647,N_24555);
nand UO_359 (O_359,N_24810,N_24886);
nor UO_360 (O_360,N_24669,N_24637);
or UO_361 (O_361,N_24994,N_24796);
nor UO_362 (O_362,N_24800,N_24648);
or UO_363 (O_363,N_24828,N_24674);
xnor UO_364 (O_364,N_24564,N_24999);
and UO_365 (O_365,N_24853,N_24903);
and UO_366 (O_366,N_24865,N_24817);
or UO_367 (O_367,N_24902,N_24879);
or UO_368 (O_368,N_24726,N_24793);
xor UO_369 (O_369,N_24777,N_24703);
xor UO_370 (O_370,N_24605,N_24541);
nand UO_371 (O_371,N_24795,N_24733);
xor UO_372 (O_372,N_24553,N_24730);
and UO_373 (O_373,N_24902,N_24737);
or UO_374 (O_374,N_24524,N_24728);
xnor UO_375 (O_375,N_24546,N_24533);
nand UO_376 (O_376,N_24635,N_24795);
nand UO_377 (O_377,N_24711,N_24807);
and UO_378 (O_378,N_24585,N_24926);
nor UO_379 (O_379,N_24863,N_24669);
nand UO_380 (O_380,N_24949,N_24985);
and UO_381 (O_381,N_24840,N_24925);
or UO_382 (O_382,N_24585,N_24997);
xor UO_383 (O_383,N_24888,N_24512);
xnor UO_384 (O_384,N_24654,N_24845);
xor UO_385 (O_385,N_24659,N_24510);
or UO_386 (O_386,N_24993,N_24686);
and UO_387 (O_387,N_24507,N_24795);
nor UO_388 (O_388,N_24782,N_24865);
and UO_389 (O_389,N_24577,N_24741);
and UO_390 (O_390,N_24818,N_24998);
xor UO_391 (O_391,N_24644,N_24758);
and UO_392 (O_392,N_24941,N_24817);
nor UO_393 (O_393,N_24768,N_24804);
and UO_394 (O_394,N_24583,N_24738);
nor UO_395 (O_395,N_24761,N_24661);
nor UO_396 (O_396,N_24804,N_24597);
nor UO_397 (O_397,N_24975,N_24671);
xnor UO_398 (O_398,N_24936,N_24843);
or UO_399 (O_399,N_24912,N_24865);
nand UO_400 (O_400,N_24579,N_24976);
or UO_401 (O_401,N_24711,N_24521);
nand UO_402 (O_402,N_24632,N_24840);
nor UO_403 (O_403,N_24600,N_24722);
and UO_404 (O_404,N_24592,N_24920);
xor UO_405 (O_405,N_24563,N_24610);
or UO_406 (O_406,N_24795,N_24957);
xnor UO_407 (O_407,N_24800,N_24712);
or UO_408 (O_408,N_24695,N_24520);
or UO_409 (O_409,N_24820,N_24881);
or UO_410 (O_410,N_24696,N_24671);
xor UO_411 (O_411,N_24632,N_24950);
nor UO_412 (O_412,N_24849,N_24650);
xnor UO_413 (O_413,N_24624,N_24564);
nand UO_414 (O_414,N_24686,N_24649);
and UO_415 (O_415,N_24709,N_24908);
or UO_416 (O_416,N_24919,N_24731);
xor UO_417 (O_417,N_24986,N_24521);
nand UO_418 (O_418,N_24903,N_24646);
and UO_419 (O_419,N_24524,N_24610);
xnor UO_420 (O_420,N_24502,N_24670);
or UO_421 (O_421,N_24822,N_24674);
nand UO_422 (O_422,N_24772,N_24752);
nand UO_423 (O_423,N_24506,N_24509);
or UO_424 (O_424,N_24588,N_24644);
xor UO_425 (O_425,N_24718,N_24974);
or UO_426 (O_426,N_24775,N_24996);
or UO_427 (O_427,N_24736,N_24517);
nand UO_428 (O_428,N_24839,N_24589);
or UO_429 (O_429,N_24601,N_24690);
or UO_430 (O_430,N_24653,N_24514);
nand UO_431 (O_431,N_24821,N_24512);
or UO_432 (O_432,N_24556,N_24788);
xnor UO_433 (O_433,N_24775,N_24514);
xor UO_434 (O_434,N_24703,N_24629);
xor UO_435 (O_435,N_24507,N_24514);
and UO_436 (O_436,N_24828,N_24501);
and UO_437 (O_437,N_24579,N_24959);
and UO_438 (O_438,N_24889,N_24711);
or UO_439 (O_439,N_24932,N_24526);
or UO_440 (O_440,N_24991,N_24831);
xor UO_441 (O_441,N_24855,N_24578);
or UO_442 (O_442,N_24693,N_24616);
nor UO_443 (O_443,N_24570,N_24790);
xnor UO_444 (O_444,N_24625,N_24526);
nor UO_445 (O_445,N_24913,N_24804);
xnor UO_446 (O_446,N_24643,N_24831);
and UO_447 (O_447,N_24622,N_24584);
xor UO_448 (O_448,N_24756,N_24833);
nand UO_449 (O_449,N_24861,N_24684);
and UO_450 (O_450,N_24765,N_24861);
or UO_451 (O_451,N_24544,N_24575);
xor UO_452 (O_452,N_24504,N_24640);
or UO_453 (O_453,N_24619,N_24936);
xnor UO_454 (O_454,N_24575,N_24577);
or UO_455 (O_455,N_24890,N_24573);
or UO_456 (O_456,N_24811,N_24534);
or UO_457 (O_457,N_24550,N_24665);
nand UO_458 (O_458,N_24828,N_24716);
or UO_459 (O_459,N_24588,N_24918);
and UO_460 (O_460,N_24617,N_24903);
nand UO_461 (O_461,N_24752,N_24801);
nor UO_462 (O_462,N_24874,N_24780);
and UO_463 (O_463,N_24830,N_24531);
or UO_464 (O_464,N_24545,N_24647);
or UO_465 (O_465,N_24607,N_24951);
or UO_466 (O_466,N_24761,N_24981);
nor UO_467 (O_467,N_24608,N_24582);
nand UO_468 (O_468,N_24712,N_24846);
nand UO_469 (O_469,N_24697,N_24869);
xor UO_470 (O_470,N_24591,N_24596);
and UO_471 (O_471,N_24882,N_24893);
and UO_472 (O_472,N_24878,N_24692);
or UO_473 (O_473,N_24583,N_24696);
nor UO_474 (O_474,N_24712,N_24552);
nor UO_475 (O_475,N_24948,N_24760);
xor UO_476 (O_476,N_24711,N_24771);
nor UO_477 (O_477,N_24838,N_24972);
nand UO_478 (O_478,N_24966,N_24738);
nor UO_479 (O_479,N_24511,N_24716);
or UO_480 (O_480,N_24513,N_24682);
nand UO_481 (O_481,N_24932,N_24716);
nand UO_482 (O_482,N_24667,N_24753);
nor UO_483 (O_483,N_24906,N_24568);
nor UO_484 (O_484,N_24813,N_24604);
or UO_485 (O_485,N_24876,N_24506);
and UO_486 (O_486,N_24928,N_24561);
nand UO_487 (O_487,N_24597,N_24692);
xor UO_488 (O_488,N_24577,N_24664);
nor UO_489 (O_489,N_24548,N_24501);
nand UO_490 (O_490,N_24536,N_24870);
nand UO_491 (O_491,N_24770,N_24653);
or UO_492 (O_492,N_24882,N_24747);
nor UO_493 (O_493,N_24529,N_24935);
and UO_494 (O_494,N_24906,N_24555);
or UO_495 (O_495,N_24711,N_24933);
or UO_496 (O_496,N_24987,N_24569);
or UO_497 (O_497,N_24913,N_24968);
nand UO_498 (O_498,N_24933,N_24818);
nor UO_499 (O_499,N_24939,N_24951);
and UO_500 (O_500,N_24869,N_24653);
nand UO_501 (O_501,N_24865,N_24688);
xor UO_502 (O_502,N_24650,N_24519);
or UO_503 (O_503,N_24557,N_24908);
xnor UO_504 (O_504,N_24999,N_24916);
and UO_505 (O_505,N_24764,N_24685);
or UO_506 (O_506,N_24772,N_24769);
or UO_507 (O_507,N_24682,N_24645);
nor UO_508 (O_508,N_24793,N_24735);
and UO_509 (O_509,N_24942,N_24725);
nor UO_510 (O_510,N_24938,N_24607);
nand UO_511 (O_511,N_24651,N_24932);
nand UO_512 (O_512,N_24914,N_24663);
nor UO_513 (O_513,N_24789,N_24530);
or UO_514 (O_514,N_24864,N_24640);
nand UO_515 (O_515,N_24861,N_24725);
or UO_516 (O_516,N_24814,N_24600);
nor UO_517 (O_517,N_24628,N_24566);
or UO_518 (O_518,N_24963,N_24847);
nand UO_519 (O_519,N_24676,N_24630);
xnor UO_520 (O_520,N_24668,N_24653);
or UO_521 (O_521,N_24847,N_24762);
xor UO_522 (O_522,N_24544,N_24590);
xnor UO_523 (O_523,N_24626,N_24817);
nor UO_524 (O_524,N_24661,N_24949);
and UO_525 (O_525,N_24561,N_24882);
or UO_526 (O_526,N_24617,N_24667);
nor UO_527 (O_527,N_24868,N_24909);
and UO_528 (O_528,N_24963,N_24632);
xor UO_529 (O_529,N_24599,N_24780);
or UO_530 (O_530,N_24943,N_24893);
nor UO_531 (O_531,N_24909,N_24846);
nand UO_532 (O_532,N_24524,N_24540);
nor UO_533 (O_533,N_24603,N_24846);
or UO_534 (O_534,N_24950,N_24918);
or UO_535 (O_535,N_24592,N_24669);
and UO_536 (O_536,N_24942,N_24656);
and UO_537 (O_537,N_24862,N_24857);
nand UO_538 (O_538,N_24610,N_24533);
or UO_539 (O_539,N_24995,N_24537);
and UO_540 (O_540,N_24645,N_24841);
xor UO_541 (O_541,N_24753,N_24852);
nand UO_542 (O_542,N_24873,N_24592);
and UO_543 (O_543,N_24858,N_24846);
and UO_544 (O_544,N_24931,N_24641);
nand UO_545 (O_545,N_24893,N_24834);
or UO_546 (O_546,N_24888,N_24918);
nor UO_547 (O_547,N_24624,N_24857);
nor UO_548 (O_548,N_24708,N_24548);
xnor UO_549 (O_549,N_24685,N_24949);
xor UO_550 (O_550,N_24618,N_24863);
xnor UO_551 (O_551,N_24952,N_24948);
xnor UO_552 (O_552,N_24727,N_24977);
xnor UO_553 (O_553,N_24783,N_24660);
or UO_554 (O_554,N_24860,N_24501);
xnor UO_555 (O_555,N_24794,N_24695);
xnor UO_556 (O_556,N_24601,N_24989);
or UO_557 (O_557,N_24797,N_24767);
nor UO_558 (O_558,N_24606,N_24651);
nor UO_559 (O_559,N_24508,N_24892);
xor UO_560 (O_560,N_24557,N_24570);
and UO_561 (O_561,N_24686,N_24988);
or UO_562 (O_562,N_24813,N_24676);
xnor UO_563 (O_563,N_24634,N_24857);
nand UO_564 (O_564,N_24697,N_24777);
nor UO_565 (O_565,N_24673,N_24591);
or UO_566 (O_566,N_24773,N_24931);
and UO_567 (O_567,N_24508,N_24880);
and UO_568 (O_568,N_24534,N_24971);
xor UO_569 (O_569,N_24550,N_24592);
xor UO_570 (O_570,N_24976,N_24776);
nand UO_571 (O_571,N_24915,N_24948);
nand UO_572 (O_572,N_24645,N_24554);
nand UO_573 (O_573,N_24516,N_24940);
xnor UO_574 (O_574,N_24588,N_24521);
nor UO_575 (O_575,N_24764,N_24911);
nor UO_576 (O_576,N_24814,N_24941);
xnor UO_577 (O_577,N_24682,N_24736);
and UO_578 (O_578,N_24712,N_24724);
xnor UO_579 (O_579,N_24796,N_24833);
or UO_580 (O_580,N_24758,N_24567);
xnor UO_581 (O_581,N_24627,N_24634);
and UO_582 (O_582,N_24574,N_24542);
nor UO_583 (O_583,N_24661,N_24936);
or UO_584 (O_584,N_24902,N_24811);
nand UO_585 (O_585,N_24603,N_24958);
or UO_586 (O_586,N_24567,N_24752);
and UO_587 (O_587,N_24768,N_24752);
nand UO_588 (O_588,N_24731,N_24736);
nand UO_589 (O_589,N_24788,N_24789);
nand UO_590 (O_590,N_24749,N_24699);
or UO_591 (O_591,N_24759,N_24632);
nor UO_592 (O_592,N_24550,N_24538);
nand UO_593 (O_593,N_24990,N_24824);
nand UO_594 (O_594,N_24520,N_24659);
and UO_595 (O_595,N_24848,N_24873);
nand UO_596 (O_596,N_24678,N_24730);
nor UO_597 (O_597,N_24534,N_24659);
or UO_598 (O_598,N_24517,N_24566);
nor UO_599 (O_599,N_24962,N_24697);
xor UO_600 (O_600,N_24916,N_24618);
and UO_601 (O_601,N_24839,N_24556);
nor UO_602 (O_602,N_24566,N_24978);
nand UO_603 (O_603,N_24691,N_24767);
nand UO_604 (O_604,N_24691,N_24625);
or UO_605 (O_605,N_24991,N_24897);
or UO_606 (O_606,N_24587,N_24996);
nor UO_607 (O_607,N_24885,N_24864);
nor UO_608 (O_608,N_24887,N_24538);
nand UO_609 (O_609,N_24633,N_24823);
nand UO_610 (O_610,N_24541,N_24619);
xnor UO_611 (O_611,N_24895,N_24900);
nor UO_612 (O_612,N_24543,N_24660);
or UO_613 (O_613,N_24556,N_24940);
nand UO_614 (O_614,N_24720,N_24728);
and UO_615 (O_615,N_24651,N_24546);
or UO_616 (O_616,N_24943,N_24985);
xnor UO_617 (O_617,N_24978,N_24909);
nor UO_618 (O_618,N_24783,N_24762);
xnor UO_619 (O_619,N_24528,N_24695);
nand UO_620 (O_620,N_24702,N_24552);
xor UO_621 (O_621,N_24938,N_24742);
nor UO_622 (O_622,N_24613,N_24674);
xnor UO_623 (O_623,N_24644,N_24568);
nor UO_624 (O_624,N_24614,N_24510);
nand UO_625 (O_625,N_24647,N_24766);
xor UO_626 (O_626,N_24773,N_24678);
nor UO_627 (O_627,N_24738,N_24595);
and UO_628 (O_628,N_24517,N_24668);
and UO_629 (O_629,N_24711,N_24970);
nor UO_630 (O_630,N_24597,N_24750);
and UO_631 (O_631,N_24623,N_24698);
and UO_632 (O_632,N_24654,N_24717);
nor UO_633 (O_633,N_24708,N_24698);
xnor UO_634 (O_634,N_24992,N_24987);
nand UO_635 (O_635,N_24761,N_24709);
nand UO_636 (O_636,N_24667,N_24940);
nor UO_637 (O_637,N_24719,N_24628);
or UO_638 (O_638,N_24672,N_24592);
or UO_639 (O_639,N_24643,N_24929);
nand UO_640 (O_640,N_24747,N_24751);
nand UO_641 (O_641,N_24526,N_24962);
or UO_642 (O_642,N_24693,N_24698);
or UO_643 (O_643,N_24857,N_24683);
and UO_644 (O_644,N_24838,N_24517);
and UO_645 (O_645,N_24754,N_24718);
nand UO_646 (O_646,N_24997,N_24668);
and UO_647 (O_647,N_24962,N_24509);
xor UO_648 (O_648,N_24545,N_24781);
and UO_649 (O_649,N_24728,N_24576);
nand UO_650 (O_650,N_24544,N_24690);
or UO_651 (O_651,N_24998,N_24808);
nand UO_652 (O_652,N_24851,N_24762);
nor UO_653 (O_653,N_24957,N_24753);
or UO_654 (O_654,N_24542,N_24536);
nand UO_655 (O_655,N_24697,N_24859);
and UO_656 (O_656,N_24655,N_24792);
nor UO_657 (O_657,N_24787,N_24914);
nand UO_658 (O_658,N_24768,N_24684);
nand UO_659 (O_659,N_24525,N_24783);
xnor UO_660 (O_660,N_24763,N_24920);
nor UO_661 (O_661,N_24860,N_24753);
or UO_662 (O_662,N_24815,N_24554);
nor UO_663 (O_663,N_24763,N_24885);
nor UO_664 (O_664,N_24748,N_24996);
xnor UO_665 (O_665,N_24825,N_24920);
xor UO_666 (O_666,N_24863,N_24952);
or UO_667 (O_667,N_24589,N_24502);
and UO_668 (O_668,N_24643,N_24586);
or UO_669 (O_669,N_24784,N_24947);
nand UO_670 (O_670,N_24738,N_24995);
xor UO_671 (O_671,N_24885,N_24568);
nor UO_672 (O_672,N_24523,N_24718);
or UO_673 (O_673,N_24682,N_24932);
nor UO_674 (O_674,N_24514,N_24892);
xor UO_675 (O_675,N_24861,N_24827);
and UO_676 (O_676,N_24938,N_24839);
nand UO_677 (O_677,N_24627,N_24727);
nor UO_678 (O_678,N_24814,N_24537);
and UO_679 (O_679,N_24560,N_24861);
nor UO_680 (O_680,N_24594,N_24627);
xnor UO_681 (O_681,N_24631,N_24972);
or UO_682 (O_682,N_24792,N_24965);
and UO_683 (O_683,N_24703,N_24577);
nor UO_684 (O_684,N_24837,N_24542);
or UO_685 (O_685,N_24683,N_24819);
nand UO_686 (O_686,N_24515,N_24777);
xor UO_687 (O_687,N_24735,N_24943);
nand UO_688 (O_688,N_24797,N_24796);
nor UO_689 (O_689,N_24660,N_24510);
or UO_690 (O_690,N_24762,N_24711);
xor UO_691 (O_691,N_24778,N_24915);
nor UO_692 (O_692,N_24868,N_24691);
nand UO_693 (O_693,N_24738,N_24862);
and UO_694 (O_694,N_24808,N_24672);
and UO_695 (O_695,N_24823,N_24606);
nand UO_696 (O_696,N_24574,N_24570);
and UO_697 (O_697,N_24743,N_24906);
or UO_698 (O_698,N_24964,N_24948);
nand UO_699 (O_699,N_24606,N_24644);
xnor UO_700 (O_700,N_24759,N_24721);
nand UO_701 (O_701,N_24746,N_24868);
nor UO_702 (O_702,N_24930,N_24936);
xor UO_703 (O_703,N_24826,N_24640);
xnor UO_704 (O_704,N_24821,N_24986);
xor UO_705 (O_705,N_24991,N_24623);
or UO_706 (O_706,N_24920,N_24668);
and UO_707 (O_707,N_24826,N_24663);
nand UO_708 (O_708,N_24621,N_24941);
nor UO_709 (O_709,N_24840,N_24575);
nand UO_710 (O_710,N_24767,N_24967);
nor UO_711 (O_711,N_24902,N_24562);
or UO_712 (O_712,N_24884,N_24686);
or UO_713 (O_713,N_24515,N_24943);
and UO_714 (O_714,N_24625,N_24800);
nor UO_715 (O_715,N_24520,N_24800);
xor UO_716 (O_716,N_24552,N_24935);
nor UO_717 (O_717,N_24648,N_24842);
and UO_718 (O_718,N_24704,N_24641);
nor UO_719 (O_719,N_24700,N_24986);
xnor UO_720 (O_720,N_24697,N_24887);
nor UO_721 (O_721,N_24633,N_24936);
nor UO_722 (O_722,N_24999,N_24517);
xor UO_723 (O_723,N_24728,N_24854);
or UO_724 (O_724,N_24692,N_24589);
or UO_725 (O_725,N_24928,N_24640);
nand UO_726 (O_726,N_24908,N_24577);
xnor UO_727 (O_727,N_24547,N_24650);
and UO_728 (O_728,N_24627,N_24650);
xor UO_729 (O_729,N_24906,N_24871);
nor UO_730 (O_730,N_24558,N_24573);
xnor UO_731 (O_731,N_24992,N_24998);
and UO_732 (O_732,N_24567,N_24791);
and UO_733 (O_733,N_24869,N_24559);
and UO_734 (O_734,N_24575,N_24599);
and UO_735 (O_735,N_24882,N_24970);
nand UO_736 (O_736,N_24852,N_24822);
or UO_737 (O_737,N_24692,N_24558);
and UO_738 (O_738,N_24774,N_24815);
nor UO_739 (O_739,N_24667,N_24594);
and UO_740 (O_740,N_24796,N_24897);
nor UO_741 (O_741,N_24727,N_24963);
and UO_742 (O_742,N_24949,N_24849);
nand UO_743 (O_743,N_24975,N_24580);
nor UO_744 (O_744,N_24649,N_24906);
nor UO_745 (O_745,N_24596,N_24500);
or UO_746 (O_746,N_24640,N_24910);
and UO_747 (O_747,N_24849,N_24732);
xor UO_748 (O_748,N_24719,N_24957);
xor UO_749 (O_749,N_24767,N_24880);
nor UO_750 (O_750,N_24728,N_24723);
xnor UO_751 (O_751,N_24786,N_24732);
xor UO_752 (O_752,N_24796,N_24858);
nor UO_753 (O_753,N_24673,N_24650);
or UO_754 (O_754,N_24938,N_24645);
nand UO_755 (O_755,N_24986,N_24773);
nand UO_756 (O_756,N_24695,N_24588);
or UO_757 (O_757,N_24565,N_24804);
nand UO_758 (O_758,N_24860,N_24631);
xnor UO_759 (O_759,N_24597,N_24589);
nor UO_760 (O_760,N_24904,N_24872);
xnor UO_761 (O_761,N_24921,N_24650);
xor UO_762 (O_762,N_24921,N_24882);
or UO_763 (O_763,N_24512,N_24569);
nand UO_764 (O_764,N_24858,N_24975);
and UO_765 (O_765,N_24915,N_24921);
nor UO_766 (O_766,N_24846,N_24722);
and UO_767 (O_767,N_24861,N_24786);
nor UO_768 (O_768,N_24729,N_24782);
xnor UO_769 (O_769,N_24561,N_24980);
or UO_770 (O_770,N_24983,N_24519);
xnor UO_771 (O_771,N_24721,N_24528);
nand UO_772 (O_772,N_24940,N_24674);
xor UO_773 (O_773,N_24655,N_24595);
or UO_774 (O_774,N_24791,N_24580);
and UO_775 (O_775,N_24663,N_24664);
and UO_776 (O_776,N_24896,N_24600);
nor UO_777 (O_777,N_24538,N_24884);
and UO_778 (O_778,N_24566,N_24608);
or UO_779 (O_779,N_24513,N_24711);
or UO_780 (O_780,N_24834,N_24528);
or UO_781 (O_781,N_24977,N_24691);
and UO_782 (O_782,N_24832,N_24852);
nor UO_783 (O_783,N_24665,N_24802);
and UO_784 (O_784,N_24989,N_24887);
xnor UO_785 (O_785,N_24520,N_24545);
nand UO_786 (O_786,N_24867,N_24691);
nor UO_787 (O_787,N_24810,N_24696);
nor UO_788 (O_788,N_24788,N_24876);
nand UO_789 (O_789,N_24810,N_24828);
xor UO_790 (O_790,N_24922,N_24611);
nand UO_791 (O_791,N_24879,N_24602);
xnor UO_792 (O_792,N_24721,N_24902);
and UO_793 (O_793,N_24851,N_24637);
nand UO_794 (O_794,N_24765,N_24918);
xnor UO_795 (O_795,N_24679,N_24763);
or UO_796 (O_796,N_24598,N_24909);
xor UO_797 (O_797,N_24797,N_24623);
nor UO_798 (O_798,N_24668,N_24625);
or UO_799 (O_799,N_24910,N_24802);
nor UO_800 (O_800,N_24799,N_24740);
xnor UO_801 (O_801,N_24940,N_24515);
nor UO_802 (O_802,N_24975,N_24828);
or UO_803 (O_803,N_24625,N_24873);
nand UO_804 (O_804,N_24609,N_24693);
xor UO_805 (O_805,N_24974,N_24518);
and UO_806 (O_806,N_24817,N_24828);
nor UO_807 (O_807,N_24798,N_24803);
nor UO_808 (O_808,N_24978,N_24606);
and UO_809 (O_809,N_24868,N_24878);
nand UO_810 (O_810,N_24827,N_24510);
and UO_811 (O_811,N_24892,N_24894);
xnor UO_812 (O_812,N_24576,N_24730);
nand UO_813 (O_813,N_24511,N_24910);
and UO_814 (O_814,N_24674,N_24675);
nor UO_815 (O_815,N_24885,N_24845);
xor UO_816 (O_816,N_24921,N_24968);
nand UO_817 (O_817,N_24564,N_24679);
xnor UO_818 (O_818,N_24859,N_24572);
xnor UO_819 (O_819,N_24872,N_24552);
nand UO_820 (O_820,N_24616,N_24922);
or UO_821 (O_821,N_24643,N_24544);
xnor UO_822 (O_822,N_24886,N_24715);
xor UO_823 (O_823,N_24873,N_24608);
and UO_824 (O_824,N_24596,N_24676);
and UO_825 (O_825,N_24634,N_24534);
nor UO_826 (O_826,N_24857,N_24789);
xnor UO_827 (O_827,N_24897,N_24778);
nand UO_828 (O_828,N_24682,N_24854);
and UO_829 (O_829,N_24667,N_24603);
nand UO_830 (O_830,N_24644,N_24626);
or UO_831 (O_831,N_24694,N_24635);
nor UO_832 (O_832,N_24868,N_24574);
and UO_833 (O_833,N_24571,N_24876);
nor UO_834 (O_834,N_24888,N_24941);
nand UO_835 (O_835,N_24860,N_24865);
or UO_836 (O_836,N_24540,N_24607);
and UO_837 (O_837,N_24779,N_24991);
xnor UO_838 (O_838,N_24669,N_24559);
and UO_839 (O_839,N_24549,N_24841);
and UO_840 (O_840,N_24927,N_24664);
nor UO_841 (O_841,N_24927,N_24937);
or UO_842 (O_842,N_24789,N_24925);
and UO_843 (O_843,N_24595,N_24944);
nand UO_844 (O_844,N_24546,N_24645);
nor UO_845 (O_845,N_24680,N_24573);
nand UO_846 (O_846,N_24502,N_24891);
nor UO_847 (O_847,N_24646,N_24838);
nor UO_848 (O_848,N_24925,N_24875);
or UO_849 (O_849,N_24600,N_24573);
nor UO_850 (O_850,N_24877,N_24687);
and UO_851 (O_851,N_24865,N_24531);
xor UO_852 (O_852,N_24746,N_24896);
and UO_853 (O_853,N_24613,N_24982);
nand UO_854 (O_854,N_24882,N_24807);
and UO_855 (O_855,N_24953,N_24669);
and UO_856 (O_856,N_24544,N_24934);
xor UO_857 (O_857,N_24555,N_24971);
xor UO_858 (O_858,N_24642,N_24960);
xnor UO_859 (O_859,N_24906,N_24581);
or UO_860 (O_860,N_24612,N_24629);
xnor UO_861 (O_861,N_24976,N_24996);
or UO_862 (O_862,N_24621,N_24550);
nor UO_863 (O_863,N_24562,N_24577);
nor UO_864 (O_864,N_24608,N_24609);
nand UO_865 (O_865,N_24546,N_24844);
or UO_866 (O_866,N_24758,N_24638);
nor UO_867 (O_867,N_24712,N_24662);
nand UO_868 (O_868,N_24963,N_24633);
nor UO_869 (O_869,N_24561,N_24650);
and UO_870 (O_870,N_24632,N_24908);
and UO_871 (O_871,N_24682,N_24993);
nand UO_872 (O_872,N_24839,N_24977);
nor UO_873 (O_873,N_24675,N_24908);
nand UO_874 (O_874,N_24946,N_24978);
or UO_875 (O_875,N_24919,N_24551);
nor UO_876 (O_876,N_24606,N_24616);
xnor UO_877 (O_877,N_24522,N_24517);
xor UO_878 (O_878,N_24603,N_24889);
nand UO_879 (O_879,N_24802,N_24827);
and UO_880 (O_880,N_24514,N_24989);
and UO_881 (O_881,N_24673,N_24963);
xnor UO_882 (O_882,N_24855,N_24754);
nor UO_883 (O_883,N_24883,N_24943);
xor UO_884 (O_884,N_24743,N_24953);
nand UO_885 (O_885,N_24646,N_24538);
and UO_886 (O_886,N_24696,N_24628);
xnor UO_887 (O_887,N_24811,N_24716);
nor UO_888 (O_888,N_24887,N_24897);
nand UO_889 (O_889,N_24844,N_24782);
or UO_890 (O_890,N_24949,N_24916);
nand UO_891 (O_891,N_24635,N_24833);
and UO_892 (O_892,N_24673,N_24555);
or UO_893 (O_893,N_24697,N_24518);
nor UO_894 (O_894,N_24868,N_24709);
or UO_895 (O_895,N_24921,N_24955);
xor UO_896 (O_896,N_24804,N_24802);
xnor UO_897 (O_897,N_24759,N_24580);
nand UO_898 (O_898,N_24774,N_24888);
xor UO_899 (O_899,N_24552,N_24742);
or UO_900 (O_900,N_24577,N_24995);
and UO_901 (O_901,N_24534,N_24938);
and UO_902 (O_902,N_24954,N_24697);
nand UO_903 (O_903,N_24826,N_24535);
xnor UO_904 (O_904,N_24606,N_24655);
and UO_905 (O_905,N_24745,N_24877);
nand UO_906 (O_906,N_24772,N_24943);
nand UO_907 (O_907,N_24514,N_24597);
and UO_908 (O_908,N_24617,N_24728);
nand UO_909 (O_909,N_24627,N_24996);
xnor UO_910 (O_910,N_24911,N_24742);
xnor UO_911 (O_911,N_24948,N_24635);
and UO_912 (O_912,N_24744,N_24978);
nor UO_913 (O_913,N_24672,N_24941);
or UO_914 (O_914,N_24881,N_24667);
xor UO_915 (O_915,N_24654,N_24906);
nor UO_916 (O_916,N_24782,N_24563);
nand UO_917 (O_917,N_24826,N_24680);
xor UO_918 (O_918,N_24872,N_24763);
nand UO_919 (O_919,N_24593,N_24925);
nand UO_920 (O_920,N_24927,N_24700);
nor UO_921 (O_921,N_24561,N_24831);
xnor UO_922 (O_922,N_24919,N_24850);
nor UO_923 (O_923,N_24961,N_24769);
nand UO_924 (O_924,N_24506,N_24818);
or UO_925 (O_925,N_24635,N_24523);
nor UO_926 (O_926,N_24713,N_24878);
nand UO_927 (O_927,N_24892,N_24742);
nand UO_928 (O_928,N_24678,N_24857);
and UO_929 (O_929,N_24561,N_24627);
nor UO_930 (O_930,N_24991,N_24532);
nand UO_931 (O_931,N_24883,N_24896);
or UO_932 (O_932,N_24743,N_24653);
nor UO_933 (O_933,N_24916,N_24964);
nand UO_934 (O_934,N_24859,N_24860);
and UO_935 (O_935,N_24907,N_24714);
and UO_936 (O_936,N_24832,N_24985);
nand UO_937 (O_937,N_24722,N_24795);
nor UO_938 (O_938,N_24657,N_24995);
and UO_939 (O_939,N_24765,N_24959);
nand UO_940 (O_940,N_24981,N_24701);
xor UO_941 (O_941,N_24533,N_24954);
or UO_942 (O_942,N_24919,N_24849);
or UO_943 (O_943,N_24983,N_24656);
xor UO_944 (O_944,N_24928,N_24655);
nor UO_945 (O_945,N_24656,N_24766);
and UO_946 (O_946,N_24971,N_24531);
or UO_947 (O_947,N_24917,N_24715);
nor UO_948 (O_948,N_24543,N_24795);
xor UO_949 (O_949,N_24532,N_24868);
or UO_950 (O_950,N_24935,N_24651);
and UO_951 (O_951,N_24672,N_24671);
or UO_952 (O_952,N_24854,N_24669);
nand UO_953 (O_953,N_24751,N_24856);
and UO_954 (O_954,N_24985,N_24544);
and UO_955 (O_955,N_24545,N_24929);
xnor UO_956 (O_956,N_24869,N_24891);
nor UO_957 (O_957,N_24598,N_24697);
nor UO_958 (O_958,N_24916,N_24635);
nor UO_959 (O_959,N_24680,N_24654);
nand UO_960 (O_960,N_24523,N_24994);
or UO_961 (O_961,N_24849,N_24709);
and UO_962 (O_962,N_24749,N_24781);
nor UO_963 (O_963,N_24586,N_24896);
and UO_964 (O_964,N_24502,N_24839);
nand UO_965 (O_965,N_24889,N_24742);
xor UO_966 (O_966,N_24555,N_24782);
nand UO_967 (O_967,N_24669,N_24623);
nand UO_968 (O_968,N_24742,N_24569);
nand UO_969 (O_969,N_24652,N_24821);
and UO_970 (O_970,N_24885,N_24806);
or UO_971 (O_971,N_24588,N_24510);
and UO_972 (O_972,N_24928,N_24730);
nand UO_973 (O_973,N_24979,N_24995);
xnor UO_974 (O_974,N_24705,N_24943);
nor UO_975 (O_975,N_24504,N_24586);
xnor UO_976 (O_976,N_24511,N_24912);
or UO_977 (O_977,N_24916,N_24577);
xor UO_978 (O_978,N_24919,N_24880);
xnor UO_979 (O_979,N_24602,N_24711);
nand UO_980 (O_980,N_24612,N_24521);
nand UO_981 (O_981,N_24838,N_24726);
and UO_982 (O_982,N_24771,N_24547);
or UO_983 (O_983,N_24662,N_24631);
nand UO_984 (O_984,N_24518,N_24577);
nand UO_985 (O_985,N_24803,N_24996);
or UO_986 (O_986,N_24609,N_24607);
and UO_987 (O_987,N_24849,N_24713);
and UO_988 (O_988,N_24790,N_24719);
and UO_989 (O_989,N_24599,N_24850);
and UO_990 (O_990,N_24518,N_24570);
nor UO_991 (O_991,N_24783,N_24781);
or UO_992 (O_992,N_24960,N_24651);
nor UO_993 (O_993,N_24803,N_24648);
or UO_994 (O_994,N_24564,N_24946);
nand UO_995 (O_995,N_24891,N_24940);
and UO_996 (O_996,N_24530,N_24535);
or UO_997 (O_997,N_24917,N_24707);
and UO_998 (O_998,N_24712,N_24883);
and UO_999 (O_999,N_24704,N_24639);
or UO_1000 (O_1000,N_24959,N_24591);
nor UO_1001 (O_1001,N_24604,N_24711);
or UO_1002 (O_1002,N_24837,N_24553);
or UO_1003 (O_1003,N_24812,N_24731);
nor UO_1004 (O_1004,N_24824,N_24776);
nor UO_1005 (O_1005,N_24759,N_24780);
or UO_1006 (O_1006,N_24873,N_24585);
or UO_1007 (O_1007,N_24639,N_24667);
nand UO_1008 (O_1008,N_24945,N_24854);
and UO_1009 (O_1009,N_24725,N_24732);
nor UO_1010 (O_1010,N_24884,N_24952);
nor UO_1011 (O_1011,N_24692,N_24508);
or UO_1012 (O_1012,N_24995,N_24799);
xor UO_1013 (O_1013,N_24790,N_24500);
xor UO_1014 (O_1014,N_24901,N_24934);
xor UO_1015 (O_1015,N_24721,N_24932);
and UO_1016 (O_1016,N_24784,N_24800);
or UO_1017 (O_1017,N_24577,N_24925);
xor UO_1018 (O_1018,N_24622,N_24948);
xor UO_1019 (O_1019,N_24609,N_24660);
or UO_1020 (O_1020,N_24787,N_24999);
or UO_1021 (O_1021,N_24581,N_24596);
nor UO_1022 (O_1022,N_24663,N_24912);
xnor UO_1023 (O_1023,N_24631,N_24884);
nand UO_1024 (O_1024,N_24589,N_24778);
xnor UO_1025 (O_1025,N_24581,N_24788);
xor UO_1026 (O_1026,N_24855,N_24587);
xor UO_1027 (O_1027,N_24538,N_24941);
nand UO_1028 (O_1028,N_24707,N_24912);
xnor UO_1029 (O_1029,N_24739,N_24713);
nor UO_1030 (O_1030,N_24923,N_24634);
nor UO_1031 (O_1031,N_24831,N_24832);
or UO_1032 (O_1032,N_24825,N_24664);
nand UO_1033 (O_1033,N_24923,N_24637);
xor UO_1034 (O_1034,N_24703,N_24895);
or UO_1035 (O_1035,N_24650,N_24587);
nor UO_1036 (O_1036,N_24882,N_24540);
xor UO_1037 (O_1037,N_24548,N_24558);
nor UO_1038 (O_1038,N_24940,N_24731);
or UO_1039 (O_1039,N_24932,N_24839);
and UO_1040 (O_1040,N_24766,N_24597);
and UO_1041 (O_1041,N_24826,N_24706);
xnor UO_1042 (O_1042,N_24520,N_24979);
nor UO_1043 (O_1043,N_24788,N_24804);
nor UO_1044 (O_1044,N_24500,N_24689);
or UO_1045 (O_1045,N_24836,N_24901);
nor UO_1046 (O_1046,N_24753,N_24626);
or UO_1047 (O_1047,N_24843,N_24559);
nor UO_1048 (O_1048,N_24842,N_24672);
xnor UO_1049 (O_1049,N_24638,N_24728);
or UO_1050 (O_1050,N_24699,N_24709);
xor UO_1051 (O_1051,N_24595,N_24797);
nand UO_1052 (O_1052,N_24817,N_24585);
and UO_1053 (O_1053,N_24864,N_24675);
nor UO_1054 (O_1054,N_24811,N_24894);
or UO_1055 (O_1055,N_24506,N_24955);
xor UO_1056 (O_1056,N_24828,N_24963);
nand UO_1057 (O_1057,N_24766,N_24933);
and UO_1058 (O_1058,N_24873,N_24850);
nor UO_1059 (O_1059,N_24627,N_24841);
or UO_1060 (O_1060,N_24628,N_24806);
xnor UO_1061 (O_1061,N_24630,N_24679);
and UO_1062 (O_1062,N_24908,N_24689);
or UO_1063 (O_1063,N_24929,N_24546);
xor UO_1064 (O_1064,N_24694,N_24902);
or UO_1065 (O_1065,N_24690,N_24710);
and UO_1066 (O_1066,N_24596,N_24507);
and UO_1067 (O_1067,N_24960,N_24564);
nor UO_1068 (O_1068,N_24745,N_24670);
or UO_1069 (O_1069,N_24783,N_24673);
nand UO_1070 (O_1070,N_24670,N_24529);
xor UO_1071 (O_1071,N_24699,N_24671);
and UO_1072 (O_1072,N_24926,N_24692);
or UO_1073 (O_1073,N_24569,N_24888);
xnor UO_1074 (O_1074,N_24743,N_24615);
and UO_1075 (O_1075,N_24647,N_24643);
or UO_1076 (O_1076,N_24876,N_24931);
nand UO_1077 (O_1077,N_24754,N_24936);
nor UO_1078 (O_1078,N_24908,N_24973);
or UO_1079 (O_1079,N_24775,N_24527);
and UO_1080 (O_1080,N_24882,N_24766);
and UO_1081 (O_1081,N_24776,N_24749);
xnor UO_1082 (O_1082,N_24530,N_24936);
xor UO_1083 (O_1083,N_24673,N_24960);
or UO_1084 (O_1084,N_24654,N_24693);
or UO_1085 (O_1085,N_24518,N_24892);
xor UO_1086 (O_1086,N_24757,N_24627);
or UO_1087 (O_1087,N_24693,N_24803);
nor UO_1088 (O_1088,N_24882,N_24505);
xor UO_1089 (O_1089,N_24683,N_24739);
nor UO_1090 (O_1090,N_24522,N_24907);
and UO_1091 (O_1091,N_24901,N_24679);
nor UO_1092 (O_1092,N_24998,N_24761);
nor UO_1093 (O_1093,N_24666,N_24761);
nand UO_1094 (O_1094,N_24771,N_24872);
xnor UO_1095 (O_1095,N_24553,N_24976);
nor UO_1096 (O_1096,N_24762,N_24959);
nand UO_1097 (O_1097,N_24715,N_24584);
or UO_1098 (O_1098,N_24553,N_24622);
and UO_1099 (O_1099,N_24818,N_24703);
or UO_1100 (O_1100,N_24566,N_24815);
nand UO_1101 (O_1101,N_24645,N_24866);
and UO_1102 (O_1102,N_24695,N_24844);
nand UO_1103 (O_1103,N_24841,N_24643);
nor UO_1104 (O_1104,N_24843,N_24829);
and UO_1105 (O_1105,N_24948,N_24692);
xnor UO_1106 (O_1106,N_24822,N_24932);
nand UO_1107 (O_1107,N_24509,N_24992);
xor UO_1108 (O_1108,N_24677,N_24812);
or UO_1109 (O_1109,N_24561,N_24982);
or UO_1110 (O_1110,N_24520,N_24954);
nor UO_1111 (O_1111,N_24766,N_24851);
nor UO_1112 (O_1112,N_24681,N_24934);
xor UO_1113 (O_1113,N_24582,N_24939);
xnor UO_1114 (O_1114,N_24583,N_24880);
and UO_1115 (O_1115,N_24905,N_24964);
nor UO_1116 (O_1116,N_24632,N_24644);
nand UO_1117 (O_1117,N_24571,N_24926);
or UO_1118 (O_1118,N_24918,N_24758);
xnor UO_1119 (O_1119,N_24756,N_24709);
nand UO_1120 (O_1120,N_24966,N_24706);
and UO_1121 (O_1121,N_24960,N_24627);
nor UO_1122 (O_1122,N_24501,N_24932);
nand UO_1123 (O_1123,N_24766,N_24887);
nor UO_1124 (O_1124,N_24786,N_24936);
or UO_1125 (O_1125,N_24786,N_24632);
nor UO_1126 (O_1126,N_24835,N_24902);
and UO_1127 (O_1127,N_24908,N_24540);
nor UO_1128 (O_1128,N_24512,N_24642);
xnor UO_1129 (O_1129,N_24523,N_24773);
nor UO_1130 (O_1130,N_24691,N_24748);
or UO_1131 (O_1131,N_24745,N_24907);
nor UO_1132 (O_1132,N_24551,N_24647);
or UO_1133 (O_1133,N_24893,N_24942);
and UO_1134 (O_1134,N_24759,N_24874);
nand UO_1135 (O_1135,N_24756,N_24683);
nor UO_1136 (O_1136,N_24610,N_24706);
and UO_1137 (O_1137,N_24777,N_24665);
or UO_1138 (O_1138,N_24610,N_24938);
nor UO_1139 (O_1139,N_24948,N_24598);
xnor UO_1140 (O_1140,N_24565,N_24928);
and UO_1141 (O_1141,N_24622,N_24903);
or UO_1142 (O_1142,N_24713,N_24856);
nor UO_1143 (O_1143,N_24612,N_24891);
or UO_1144 (O_1144,N_24543,N_24916);
xor UO_1145 (O_1145,N_24663,N_24813);
nor UO_1146 (O_1146,N_24776,N_24877);
and UO_1147 (O_1147,N_24743,N_24622);
and UO_1148 (O_1148,N_24614,N_24613);
and UO_1149 (O_1149,N_24901,N_24785);
nor UO_1150 (O_1150,N_24880,N_24646);
and UO_1151 (O_1151,N_24574,N_24551);
nand UO_1152 (O_1152,N_24920,N_24533);
or UO_1153 (O_1153,N_24962,N_24943);
or UO_1154 (O_1154,N_24780,N_24528);
xor UO_1155 (O_1155,N_24611,N_24941);
or UO_1156 (O_1156,N_24867,N_24800);
and UO_1157 (O_1157,N_24800,N_24519);
and UO_1158 (O_1158,N_24682,N_24658);
xnor UO_1159 (O_1159,N_24618,N_24529);
nand UO_1160 (O_1160,N_24699,N_24833);
nor UO_1161 (O_1161,N_24752,N_24530);
nand UO_1162 (O_1162,N_24523,N_24701);
and UO_1163 (O_1163,N_24995,N_24866);
nor UO_1164 (O_1164,N_24886,N_24944);
or UO_1165 (O_1165,N_24617,N_24915);
nand UO_1166 (O_1166,N_24836,N_24650);
nor UO_1167 (O_1167,N_24709,N_24812);
xnor UO_1168 (O_1168,N_24753,N_24675);
xnor UO_1169 (O_1169,N_24692,N_24522);
and UO_1170 (O_1170,N_24694,N_24929);
xor UO_1171 (O_1171,N_24561,N_24934);
or UO_1172 (O_1172,N_24816,N_24962);
nand UO_1173 (O_1173,N_24850,N_24781);
and UO_1174 (O_1174,N_24594,N_24911);
and UO_1175 (O_1175,N_24654,N_24585);
xor UO_1176 (O_1176,N_24535,N_24806);
and UO_1177 (O_1177,N_24668,N_24700);
nand UO_1178 (O_1178,N_24642,N_24764);
nand UO_1179 (O_1179,N_24585,N_24692);
or UO_1180 (O_1180,N_24694,N_24698);
nor UO_1181 (O_1181,N_24566,N_24814);
and UO_1182 (O_1182,N_24553,N_24705);
nor UO_1183 (O_1183,N_24711,N_24890);
xor UO_1184 (O_1184,N_24991,N_24879);
xor UO_1185 (O_1185,N_24911,N_24673);
and UO_1186 (O_1186,N_24665,N_24684);
and UO_1187 (O_1187,N_24570,N_24979);
xnor UO_1188 (O_1188,N_24963,N_24881);
or UO_1189 (O_1189,N_24537,N_24810);
nor UO_1190 (O_1190,N_24624,N_24543);
or UO_1191 (O_1191,N_24543,N_24500);
nor UO_1192 (O_1192,N_24701,N_24824);
and UO_1193 (O_1193,N_24712,N_24803);
and UO_1194 (O_1194,N_24541,N_24891);
or UO_1195 (O_1195,N_24623,N_24810);
or UO_1196 (O_1196,N_24701,N_24717);
or UO_1197 (O_1197,N_24511,N_24734);
nor UO_1198 (O_1198,N_24677,N_24895);
nor UO_1199 (O_1199,N_24868,N_24857);
nand UO_1200 (O_1200,N_24768,N_24593);
and UO_1201 (O_1201,N_24997,N_24857);
or UO_1202 (O_1202,N_24974,N_24856);
or UO_1203 (O_1203,N_24821,N_24529);
xnor UO_1204 (O_1204,N_24866,N_24826);
and UO_1205 (O_1205,N_24756,N_24991);
nor UO_1206 (O_1206,N_24657,N_24770);
nand UO_1207 (O_1207,N_24741,N_24576);
or UO_1208 (O_1208,N_24526,N_24923);
nor UO_1209 (O_1209,N_24974,N_24996);
nor UO_1210 (O_1210,N_24885,N_24833);
and UO_1211 (O_1211,N_24734,N_24910);
and UO_1212 (O_1212,N_24986,N_24988);
nand UO_1213 (O_1213,N_24974,N_24873);
nor UO_1214 (O_1214,N_24947,N_24935);
and UO_1215 (O_1215,N_24566,N_24811);
xnor UO_1216 (O_1216,N_24941,N_24899);
nand UO_1217 (O_1217,N_24515,N_24826);
and UO_1218 (O_1218,N_24855,N_24747);
nor UO_1219 (O_1219,N_24971,N_24791);
and UO_1220 (O_1220,N_24559,N_24608);
and UO_1221 (O_1221,N_24954,N_24591);
nand UO_1222 (O_1222,N_24674,N_24855);
nand UO_1223 (O_1223,N_24758,N_24826);
xnor UO_1224 (O_1224,N_24928,N_24504);
xor UO_1225 (O_1225,N_24559,N_24688);
xor UO_1226 (O_1226,N_24808,N_24830);
nand UO_1227 (O_1227,N_24768,N_24780);
xor UO_1228 (O_1228,N_24514,N_24696);
nor UO_1229 (O_1229,N_24866,N_24766);
xor UO_1230 (O_1230,N_24763,N_24890);
nand UO_1231 (O_1231,N_24769,N_24668);
nor UO_1232 (O_1232,N_24626,N_24939);
or UO_1233 (O_1233,N_24532,N_24811);
xnor UO_1234 (O_1234,N_24812,N_24601);
and UO_1235 (O_1235,N_24727,N_24504);
nand UO_1236 (O_1236,N_24948,N_24645);
and UO_1237 (O_1237,N_24713,N_24670);
and UO_1238 (O_1238,N_24537,N_24869);
nand UO_1239 (O_1239,N_24559,N_24753);
and UO_1240 (O_1240,N_24824,N_24612);
or UO_1241 (O_1241,N_24707,N_24943);
and UO_1242 (O_1242,N_24786,N_24528);
and UO_1243 (O_1243,N_24928,N_24834);
or UO_1244 (O_1244,N_24995,N_24509);
and UO_1245 (O_1245,N_24837,N_24913);
xnor UO_1246 (O_1246,N_24723,N_24565);
or UO_1247 (O_1247,N_24961,N_24832);
nand UO_1248 (O_1248,N_24668,N_24779);
nor UO_1249 (O_1249,N_24509,N_24858);
nand UO_1250 (O_1250,N_24771,N_24572);
and UO_1251 (O_1251,N_24976,N_24616);
xnor UO_1252 (O_1252,N_24816,N_24951);
and UO_1253 (O_1253,N_24878,N_24651);
xnor UO_1254 (O_1254,N_24995,N_24927);
nand UO_1255 (O_1255,N_24891,N_24561);
xor UO_1256 (O_1256,N_24916,N_24898);
nand UO_1257 (O_1257,N_24700,N_24852);
nor UO_1258 (O_1258,N_24934,N_24811);
nor UO_1259 (O_1259,N_24739,N_24949);
and UO_1260 (O_1260,N_24885,N_24571);
xor UO_1261 (O_1261,N_24815,N_24567);
or UO_1262 (O_1262,N_24637,N_24906);
xnor UO_1263 (O_1263,N_24737,N_24580);
nor UO_1264 (O_1264,N_24864,N_24584);
nand UO_1265 (O_1265,N_24867,N_24733);
xor UO_1266 (O_1266,N_24630,N_24705);
nand UO_1267 (O_1267,N_24691,N_24777);
nor UO_1268 (O_1268,N_24520,N_24784);
xor UO_1269 (O_1269,N_24794,N_24783);
nand UO_1270 (O_1270,N_24509,N_24705);
nand UO_1271 (O_1271,N_24857,N_24915);
xor UO_1272 (O_1272,N_24594,N_24641);
or UO_1273 (O_1273,N_24856,N_24521);
xor UO_1274 (O_1274,N_24913,N_24598);
nor UO_1275 (O_1275,N_24991,N_24562);
nor UO_1276 (O_1276,N_24545,N_24847);
nand UO_1277 (O_1277,N_24911,N_24517);
and UO_1278 (O_1278,N_24647,N_24518);
and UO_1279 (O_1279,N_24813,N_24598);
and UO_1280 (O_1280,N_24846,N_24527);
or UO_1281 (O_1281,N_24898,N_24654);
nand UO_1282 (O_1282,N_24620,N_24875);
xnor UO_1283 (O_1283,N_24760,N_24715);
and UO_1284 (O_1284,N_24950,N_24650);
or UO_1285 (O_1285,N_24666,N_24676);
or UO_1286 (O_1286,N_24995,N_24980);
and UO_1287 (O_1287,N_24667,N_24535);
and UO_1288 (O_1288,N_24925,N_24643);
and UO_1289 (O_1289,N_24906,N_24768);
nand UO_1290 (O_1290,N_24809,N_24652);
xor UO_1291 (O_1291,N_24607,N_24526);
and UO_1292 (O_1292,N_24982,N_24847);
nor UO_1293 (O_1293,N_24562,N_24820);
xnor UO_1294 (O_1294,N_24988,N_24894);
nor UO_1295 (O_1295,N_24601,N_24879);
nand UO_1296 (O_1296,N_24753,N_24765);
and UO_1297 (O_1297,N_24855,N_24916);
nand UO_1298 (O_1298,N_24883,N_24899);
nand UO_1299 (O_1299,N_24718,N_24694);
xnor UO_1300 (O_1300,N_24727,N_24912);
and UO_1301 (O_1301,N_24938,N_24852);
nor UO_1302 (O_1302,N_24769,N_24832);
nand UO_1303 (O_1303,N_24647,N_24595);
xor UO_1304 (O_1304,N_24789,N_24669);
or UO_1305 (O_1305,N_24928,N_24747);
or UO_1306 (O_1306,N_24696,N_24954);
nor UO_1307 (O_1307,N_24621,N_24644);
xnor UO_1308 (O_1308,N_24776,N_24912);
nor UO_1309 (O_1309,N_24872,N_24703);
and UO_1310 (O_1310,N_24589,N_24981);
nor UO_1311 (O_1311,N_24918,N_24834);
or UO_1312 (O_1312,N_24708,N_24899);
or UO_1313 (O_1313,N_24557,N_24948);
xnor UO_1314 (O_1314,N_24878,N_24743);
or UO_1315 (O_1315,N_24831,N_24715);
and UO_1316 (O_1316,N_24867,N_24965);
nand UO_1317 (O_1317,N_24516,N_24763);
nor UO_1318 (O_1318,N_24753,N_24550);
and UO_1319 (O_1319,N_24813,N_24526);
nand UO_1320 (O_1320,N_24989,N_24967);
nor UO_1321 (O_1321,N_24983,N_24638);
and UO_1322 (O_1322,N_24538,N_24620);
and UO_1323 (O_1323,N_24569,N_24717);
nor UO_1324 (O_1324,N_24564,N_24975);
nor UO_1325 (O_1325,N_24840,N_24693);
xnor UO_1326 (O_1326,N_24572,N_24838);
nand UO_1327 (O_1327,N_24532,N_24956);
nor UO_1328 (O_1328,N_24844,N_24615);
or UO_1329 (O_1329,N_24861,N_24963);
nand UO_1330 (O_1330,N_24545,N_24882);
xor UO_1331 (O_1331,N_24523,N_24895);
xnor UO_1332 (O_1332,N_24506,N_24693);
xor UO_1333 (O_1333,N_24830,N_24716);
or UO_1334 (O_1334,N_24540,N_24968);
xor UO_1335 (O_1335,N_24926,N_24672);
nand UO_1336 (O_1336,N_24826,N_24598);
nor UO_1337 (O_1337,N_24783,N_24791);
and UO_1338 (O_1338,N_24779,N_24603);
nand UO_1339 (O_1339,N_24540,N_24745);
nor UO_1340 (O_1340,N_24944,N_24619);
xor UO_1341 (O_1341,N_24790,N_24965);
nor UO_1342 (O_1342,N_24824,N_24934);
nand UO_1343 (O_1343,N_24712,N_24579);
and UO_1344 (O_1344,N_24645,N_24905);
nor UO_1345 (O_1345,N_24731,N_24931);
and UO_1346 (O_1346,N_24774,N_24865);
nand UO_1347 (O_1347,N_24763,N_24772);
xor UO_1348 (O_1348,N_24874,N_24743);
nor UO_1349 (O_1349,N_24676,N_24716);
and UO_1350 (O_1350,N_24535,N_24653);
xnor UO_1351 (O_1351,N_24556,N_24579);
or UO_1352 (O_1352,N_24652,N_24831);
or UO_1353 (O_1353,N_24570,N_24880);
or UO_1354 (O_1354,N_24774,N_24941);
xnor UO_1355 (O_1355,N_24615,N_24868);
xor UO_1356 (O_1356,N_24724,N_24845);
nor UO_1357 (O_1357,N_24728,N_24900);
or UO_1358 (O_1358,N_24649,N_24729);
or UO_1359 (O_1359,N_24725,N_24652);
or UO_1360 (O_1360,N_24517,N_24516);
or UO_1361 (O_1361,N_24907,N_24918);
nand UO_1362 (O_1362,N_24524,N_24504);
or UO_1363 (O_1363,N_24504,N_24667);
xnor UO_1364 (O_1364,N_24517,N_24750);
and UO_1365 (O_1365,N_24965,N_24683);
nand UO_1366 (O_1366,N_24723,N_24978);
nor UO_1367 (O_1367,N_24787,N_24774);
xnor UO_1368 (O_1368,N_24894,N_24579);
or UO_1369 (O_1369,N_24985,N_24876);
xnor UO_1370 (O_1370,N_24614,N_24549);
and UO_1371 (O_1371,N_24737,N_24707);
or UO_1372 (O_1372,N_24696,N_24833);
xor UO_1373 (O_1373,N_24589,N_24569);
or UO_1374 (O_1374,N_24939,N_24632);
and UO_1375 (O_1375,N_24538,N_24571);
nand UO_1376 (O_1376,N_24901,N_24782);
nand UO_1377 (O_1377,N_24506,N_24844);
and UO_1378 (O_1378,N_24579,N_24549);
nor UO_1379 (O_1379,N_24646,N_24936);
xor UO_1380 (O_1380,N_24970,N_24935);
nor UO_1381 (O_1381,N_24719,N_24806);
nand UO_1382 (O_1382,N_24943,N_24543);
and UO_1383 (O_1383,N_24665,N_24983);
nand UO_1384 (O_1384,N_24980,N_24812);
nand UO_1385 (O_1385,N_24630,N_24678);
nand UO_1386 (O_1386,N_24914,N_24907);
or UO_1387 (O_1387,N_24587,N_24773);
nor UO_1388 (O_1388,N_24918,N_24730);
and UO_1389 (O_1389,N_24591,N_24640);
and UO_1390 (O_1390,N_24971,N_24506);
nand UO_1391 (O_1391,N_24844,N_24953);
nand UO_1392 (O_1392,N_24744,N_24541);
xor UO_1393 (O_1393,N_24511,N_24845);
xor UO_1394 (O_1394,N_24668,N_24865);
nand UO_1395 (O_1395,N_24990,N_24854);
nor UO_1396 (O_1396,N_24672,N_24795);
xnor UO_1397 (O_1397,N_24576,N_24940);
or UO_1398 (O_1398,N_24797,N_24651);
and UO_1399 (O_1399,N_24541,N_24822);
or UO_1400 (O_1400,N_24844,N_24889);
and UO_1401 (O_1401,N_24779,N_24766);
nand UO_1402 (O_1402,N_24967,N_24931);
xnor UO_1403 (O_1403,N_24526,N_24685);
nor UO_1404 (O_1404,N_24557,N_24754);
nor UO_1405 (O_1405,N_24701,N_24885);
or UO_1406 (O_1406,N_24735,N_24796);
and UO_1407 (O_1407,N_24715,N_24693);
or UO_1408 (O_1408,N_24608,N_24728);
or UO_1409 (O_1409,N_24829,N_24502);
nor UO_1410 (O_1410,N_24775,N_24545);
nor UO_1411 (O_1411,N_24836,N_24556);
xor UO_1412 (O_1412,N_24844,N_24921);
and UO_1413 (O_1413,N_24743,N_24633);
nor UO_1414 (O_1414,N_24652,N_24844);
or UO_1415 (O_1415,N_24711,N_24549);
or UO_1416 (O_1416,N_24725,N_24676);
nor UO_1417 (O_1417,N_24570,N_24824);
nand UO_1418 (O_1418,N_24903,N_24750);
nor UO_1419 (O_1419,N_24889,N_24782);
nand UO_1420 (O_1420,N_24665,N_24538);
or UO_1421 (O_1421,N_24610,N_24741);
nor UO_1422 (O_1422,N_24683,N_24823);
or UO_1423 (O_1423,N_24722,N_24664);
nor UO_1424 (O_1424,N_24680,N_24910);
xor UO_1425 (O_1425,N_24809,N_24559);
and UO_1426 (O_1426,N_24835,N_24794);
nor UO_1427 (O_1427,N_24914,N_24866);
xnor UO_1428 (O_1428,N_24742,N_24627);
nand UO_1429 (O_1429,N_24883,N_24965);
or UO_1430 (O_1430,N_24681,N_24664);
or UO_1431 (O_1431,N_24590,N_24934);
and UO_1432 (O_1432,N_24640,N_24947);
nor UO_1433 (O_1433,N_24522,N_24730);
and UO_1434 (O_1434,N_24790,N_24539);
xnor UO_1435 (O_1435,N_24821,N_24502);
xor UO_1436 (O_1436,N_24994,N_24842);
xor UO_1437 (O_1437,N_24552,N_24614);
or UO_1438 (O_1438,N_24972,N_24559);
nand UO_1439 (O_1439,N_24531,N_24573);
nand UO_1440 (O_1440,N_24508,N_24870);
and UO_1441 (O_1441,N_24609,N_24537);
and UO_1442 (O_1442,N_24686,N_24747);
and UO_1443 (O_1443,N_24574,N_24913);
nor UO_1444 (O_1444,N_24822,N_24747);
and UO_1445 (O_1445,N_24805,N_24851);
and UO_1446 (O_1446,N_24675,N_24634);
xor UO_1447 (O_1447,N_24602,N_24808);
nand UO_1448 (O_1448,N_24756,N_24817);
nand UO_1449 (O_1449,N_24854,N_24840);
or UO_1450 (O_1450,N_24893,N_24783);
xnor UO_1451 (O_1451,N_24886,N_24744);
xnor UO_1452 (O_1452,N_24647,N_24707);
nor UO_1453 (O_1453,N_24995,N_24789);
xor UO_1454 (O_1454,N_24794,N_24614);
or UO_1455 (O_1455,N_24939,N_24915);
xor UO_1456 (O_1456,N_24880,N_24766);
or UO_1457 (O_1457,N_24902,N_24828);
xnor UO_1458 (O_1458,N_24836,N_24879);
nand UO_1459 (O_1459,N_24772,N_24567);
or UO_1460 (O_1460,N_24902,N_24786);
or UO_1461 (O_1461,N_24624,N_24648);
nand UO_1462 (O_1462,N_24980,N_24572);
or UO_1463 (O_1463,N_24604,N_24522);
nand UO_1464 (O_1464,N_24997,N_24736);
nor UO_1465 (O_1465,N_24628,N_24861);
xnor UO_1466 (O_1466,N_24977,N_24568);
nand UO_1467 (O_1467,N_24780,N_24833);
or UO_1468 (O_1468,N_24887,N_24722);
and UO_1469 (O_1469,N_24964,N_24834);
nand UO_1470 (O_1470,N_24530,N_24709);
nor UO_1471 (O_1471,N_24853,N_24514);
xnor UO_1472 (O_1472,N_24933,N_24941);
or UO_1473 (O_1473,N_24714,N_24642);
xor UO_1474 (O_1474,N_24605,N_24608);
nor UO_1475 (O_1475,N_24811,N_24743);
xor UO_1476 (O_1476,N_24950,N_24661);
xor UO_1477 (O_1477,N_24755,N_24507);
or UO_1478 (O_1478,N_24764,N_24980);
and UO_1479 (O_1479,N_24709,N_24649);
or UO_1480 (O_1480,N_24929,N_24960);
nor UO_1481 (O_1481,N_24811,N_24655);
nand UO_1482 (O_1482,N_24655,N_24567);
nand UO_1483 (O_1483,N_24571,N_24502);
nand UO_1484 (O_1484,N_24710,N_24658);
and UO_1485 (O_1485,N_24527,N_24843);
nand UO_1486 (O_1486,N_24649,N_24678);
and UO_1487 (O_1487,N_24525,N_24739);
nor UO_1488 (O_1488,N_24950,N_24999);
xnor UO_1489 (O_1489,N_24886,N_24506);
xor UO_1490 (O_1490,N_24640,N_24605);
and UO_1491 (O_1491,N_24816,N_24954);
and UO_1492 (O_1492,N_24986,N_24963);
xnor UO_1493 (O_1493,N_24615,N_24576);
or UO_1494 (O_1494,N_24554,N_24716);
and UO_1495 (O_1495,N_24507,N_24971);
and UO_1496 (O_1496,N_24931,N_24964);
xnor UO_1497 (O_1497,N_24741,N_24785);
or UO_1498 (O_1498,N_24669,N_24586);
or UO_1499 (O_1499,N_24592,N_24844);
or UO_1500 (O_1500,N_24975,N_24552);
and UO_1501 (O_1501,N_24650,N_24804);
nand UO_1502 (O_1502,N_24845,N_24510);
and UO_1503 (O_1503,N_24814,N_24790);
nor UO_1504 (O_1504,N_24774,N_24818);
or UO_1505 (O_1505,N_24968,N_24764);
nor UO_1506 (O_1506,N_24790,N_24816);
and UO_1507 (O_1507,N_24896,N_24525);
and UO_1508 (O_1508,N_24615,N_24943);
and UO_1509 (O_1509,N_24602,N_24730);
xor UO_1510 (O_1510,N_24783,N_24775);
xor UO_1511 (O_1511,N_24720,N_24939);
and UO_1512 (O_1512,N_24694,N_24952);
xor UO_1513 (O_1513,N_24704,N_24522);
and UO_1514 (O_1514,N_24678,N_24883);
nor UO_1515 (O_1515,N_24730,N_24873);
xor UO_1516 (O_1516,N_24966,N_24952);
and UO_1517 (O_1517,N_24848,N_24869);
nand UO_1518 (O_1518,N_24874,N_24939);
nand UO_1519 (O_1519,N_24533,N_24792);
nor UO_1520 (O_1520,N_24861,N_24897);
nor UO_1521 (O_1521,N_24602,N_24663);
xor UO_1522 (O_1522,N_24776,N_24816);
and UO_1523 (O_1523,N_24976,N_24546);
or UO_1524 (O_1524,N_24544,N_24713);
nor UO_1525 (O_1525,N_24638,N_24862);
or UO_1526 (O_1526,N_24519,N_24645);
nor UO_1527 (O_1527,N_24541,N_24749);
nand UO_1528 (O_1528,N_24524,N_24992);
xnor UO_1529 (O_1529,N_24740,N_24582);
nand UO_1530 (O_1530,N_24983,N_24952);
nor UO_1531 (O_1531,N_24744,N_24730);
nand UO_1532 (O_1532,N_24522,N_24880);
or UO_1533 (O_1533,N_24986,N_24906);
xnor UO_1534 (O_1534,N_24702,N_24899);
nand UO_1535 (O_1535,N_24672,N_24989);
nand UO_1536 (O_1536,N_24838,N_24693);
and UO_1537 (O_1537,N_24776,N_24626);
nor UO_1538 (O_1538,N_24821,N_24938);
nand UO_1539 (O_1539,N_24829,N_24838);
and UO_1540 (O_1540,N_24598,N_24806);
xnor UO_1541 (O_1541,N_24587,N_24807);
nor UO_1542 (O_1542,N_24731,N_24781);
xnor UO_1543 (O_1543,N_24719,N_24669);
or UO_1544 (O_1544,N_24588,N_24673);
or UO_1545 (O_1545,N_24977,N_24713);
nor UO_1546 (O_1546,N_24668,N_24830);
nand UO_1547 (O_1547,N_24537,N_24687);
or UO_1548 (O_1548,N_24954,N_24922);
and UO_1549 (O_1549,N_24682,N_24701);
and UO_1550 (O_1550,N_24542,N_24860);
nand UO_1551 (O_1551,N_24850,N_24786);
nor UO_1552 (O_1552,N_24752,N_24855);
nand UO_1553 (O_1553,N_24908,N_24816);
nand UO_1554 (O_1554,N_24768,N_24712);
or UO_1555 (O_1555,N_24633,N_24955);
nor UO_1556 (O_1556,N_24914,N_24594);
nor UO_1557 (O_1557,N_24839,N_24798);
and UO_1558 (O_1558,N_24834,N_24617);
and UO_1559 (O_1559,N_24727,N_24841);
xnor UO_1560 (O_1560,N_24517,N_24791);
and UO_1561 (O_1561,N_24934,N_24713);
or UO_1562 (O_1562,N_24727,N_24742);
nor UO_1563 (O_1563,N_24585,N_24629);
and UO_1564 (O_1564,N_24761,N_24851);
and UO_1565 (O_1565,N_24586,N_24857);
nand UO_1566 (O_1566,N_24937,N_24765);
nand UO_1567 (O_1567,N_24744,N_24963);
xnor UO_1568 (O_1568,N_24689,N_24593);
xnor UO_1569 (O_1569,N_24769,N_24812);
nand UO_1570 (O_1570,N_24978,N_24950);
xor UO_1571 (O_1571,N_24911,N_24639);
and UO_1572 (O_1572,N_24618,N_24634);
xnor UO_1573 (O_1573,N_24998,N_24529);
nor UO_1574 (O_1574,N_24712,N_24997);
nand UO_1575 (O_1575,N_24598,N_24952);
and UO_1576 (O_1576,N_24674,N_24788);
and UO_1577 (O_1577,N_24699,N_24916);
nand UO_1578 (O_1578,N_24620,N_24546);
or UO_1579 (O_1579,N_24597,N_24716);
xnor UO_1580 (O_1580,N_24790,N_24735);
xnor UO_1581 (O_1581,N_24649,N_24655);
xnor UO_1582 (O_1582,N_24987,N_24582);
nand UO_1583 (O_1583,N_24603,N_24810);
xor UO_1584 (O_1584,N_24693,N_24966);
xor UO_1585 (O_1585,N_24922,N_24863);
or UO_1586 (O_1586,N_24746,N_24616);
and UO_1587 (O_1587,N_24925,N_24566);
nor UO_1588 (O_1588,N_24833,N_24864);
nand UO_1589 (O_1589,N_24662,N_24598);
nand UO_1590 (O_1590,N_24702,N_24903);
and UO_1591 (O_1591,N_24666,N_24532);
or UO_1592 (O_1592,N_24639,N_24921);
and UO_1593 (O_1593,N_24572,N_24758);
nand UO_1594 (O_1594,N_24686,N_24964);
and UO_1595 (O_1595,N_24645,N_24708);
nand UO_1596 (O_1596,N_24719,N_24584);
nor UO_1597 (O_1597,N_24527,N_24998);
xnor UO_1598 (O_1598,N_24832,N_24642);
nand UO_1599 (O_1599,N_24732,N_24561);
and UO_1600 (O_1600,N_24708,N_24814);
or UO_1601 (O_1601,N_24606,N_24973);
and UO_1602 (O_1602,N_24623,N_24986);
nand UO_1603 (O_1603,N_24596,N_24795);
nor UO_1604 (O_1604,N_24699,N_24626);
and UO_1605 (O_1605,N_24635,N_24626);
and UO_1606 (O_1606,N_24763,N_24739);
nor UO_1607 (O_1607,N_24939,N_24863);
or UO_1608 (O_1608,N_24957,N_24905);
nor UO_1609 (O_1609,N_24961,N_24906);
nand UO_1610 (O_1610,N_24914,N_24579);
xnor UO_1611 (O_1611,N_24540,N_24612);
xor UO_1612 (O_1612,N_24759,N_24833);
nor UO_1613 (O_1613,N_24916,N_24773);
and UO_1614 (O_1614,N_24603,N_24581);
and UO_1615 (O_1615,N_24908,N_24708);
and UO_1616 (O_1616,N_24894,N_24621);
nand UO_1617 (O_1617,N_24791,N_24898);
and UO_1618 (O_1618,N_24990,N_24582);
and UO_1619 (O_1619,N_24720,N_24936);
and UO_1620 (O_1620,N_24710,N_24627);
nor UO_1621 (O_1621,N_24836,N_24861);
and UO_1622 (O_1622,N_24949,N_24829);
and UO_1623 (O_1623,N_24581,N_24597);
xnor UO_1624 (O_1624,N_24667,N_24953);
nor UO_1625 (O_1625,N_24732,N_24787);
xor UO_1626 (O_1626,N_24770,N_24522);
nor UO_1627 (O_1627,N_24659,N_24666);
and UO_1628 (O_1628,N_24943,N_24589);
xnor UO_1629 (O_1629,N_24960,N_24645);
xor UO_1630 (O_1630,N_24941,N_24795);
xnor UO_1631 (O_1631,N_24822,N_24868);
or UO_1632 (O_1632,N_24504,N_24962);
and UO_1633 (O_1633,N_24772,N_24877);
nor UO_1634 (O_1634,N_24564,N_24708);
xor UO_1635 (O_1635,N_24988,N_24813);
xor UO_1636 (O_1636,N_24595,N_24690);
and UO_1637 (O_1637,N_24759,N_24523);
xnor UO_1638 (O_1638,N_24592,N_24718);
nor UO_1639 (O_1639,N_24913,N_24831);
and UO_1640 (O_1640,N_24903,N_24972);
nor UO_1641 (O_1641,N_24621,N_24578);
or UO_1642 (O_1642,N_24739,N_24783);
or UO_1643 (O_1643,N_24707,N_24675);
or UO_1644 (O_1644,N_24738,N_24941);
or UO_1645 (O_1645,N_24587,N_24719);
or UO_1646 (O_1646,N_24517,N_24501);
nand UO_1647 (O_1647,N_24731,N_24543);
nand UO_1648 (O_1648,N_24739,N_24964);
nor UO_1649 (O_1649,N_24541,N_24637);
and UO_1650 (O_1650,N_24938,N_24683);
or UO_1651 (O_1651,N_24642,N_24578);
nand UO_1652 (O_1652,N_24747,N_24679);
and UO_1653 (O_1653,N_24667,N_24532);
and UO_1654 (O_1654,N_24973,N_24855);
and UO_1655 (O_1655,N_24508,N_24602);
xnor UO_1656 (O_1656,N_24901,N_24683);
nor UO_1657 (O_1657,N_24723,N_24548);
or UO_1658 (O_1658,N_24672,N_24739);
or UO_1659 (O_1659,N_24526,N_24698);
xnor UO_1660 (O_1660,N_24635,N_24627);
nand UO_1661 (O_1661,N_24896,N_24584);
nor UO_1662 (O_1662,N_24756,N_24509);
and UO_1663 (O_1663,N_24978,N_24620);
xor UO_1664 (O_1664,N_24994,N_24684);
nor UO_1665 (O_1665,N_24569,N_24665);
and UO_1666 (O_1666,N_24564,N_24615);
nor UO_1667 (O_1667,N_24866,N_24994);
and UO_1668 (O_1668,N_24779,N_24821);
xor UO_1669 (O_1669,N_24703,N_24919);
nand UO_1670 (O_1670,N_24524,N_24715);
or UO_1671 (O_1671,N_24818,N_24712);
and UO_1672 (O_1672,N_24823,N_24836);
nand UO_1673 (O_1673,N_24661,N_24609);
xnor UO_1674 (O_1674,N_24874,N_24876);
nor UO_1675 (O_1675,N_24574,N_24860);
or UO_1676 (O_1676,N_24978,N_24510);
nand UO_1677 (O_1677,N_24949,N_24955);
or UO_1678 (O_1678,N_24804,N_24860);
or UO_1679 (O_1679,N_24756,N_24812);
xor UO_1680 (O_1680,N_24946,N_24620);
nand UO_1681 (O_1681,N_24908,N_24761);
or UO_1682 (O_1682,N_24727,N_24802);
nand UO_1683 (O_1683,N_24719,N_24639);
nand UO_1684 (O_1684,N_24531,N_24620);
nor UO_1685 (O_1685,N_24537,N_24730);
or UO_1686 (O_1686,N_24958,N_24509);
nor UO_1687 (O_1687,N_24905,N_24658);
and UO_1688 (O_1688,N_24763,N_24565);
or UO_1689 (O_1689,N_24798,N_24699);
and UO_1690 (O_1690,N_24573,N_24615);
nor UO_1691 (O_1691,N_24653,N_24912);
and UO_1692 (O_1692,N_24655,N_24696);
or UO_1693 (O_1693,N_24507,N_24941);
or UO_1694 (O_1694,N_24764,N_24860);
and UO_1695 (O_1695,N_24879,N_24729);
and UO_1696 (O_1696,N_24731,N_24673);
and UO_1697 (O_1697,N_24987,N_24747);
xor UO_1698 (O_1698,N_24616,N_24510);
or UO_1699 (O_1699,N_24517,N_24988);
xor UO_1700 (O_1700,N_24973,N_24812);
or UO_1701 (O_1701,N_24915,N_24871);
or UO_1702 (O_1702,N_24961,N_24903);
nand UO_1703 (O_1703,N_24850,N_24920);
or UO_1704 (O_1704,N_24750,N_24738);
nand UO_1705 (O_1705,N_24788,N_24727);
xor UO_1706 (O_1706,N_24988,N_24790);
xor UO_1707 (O_1707,N_24948,N_24920);
nand UO_1708 (O_1708,N_24713,N_24540);
and UO_1709 (O_1709,N_24706,N_24626);
and UO_1710 (O_1710,N_24908,N_24576);
nor UO_1711 (O_1711,N_24853,N_24986);
or UO_1712 (O_1712,N_24829,N_24605);
xor UO_1713 (O_1713,N_24704,N_24624);
xnor UO_1714 (O_1714,N_24608,N_24938);
nand UO_1715 (O_1715,N_24846,N_24841);
xnor UO_1716 (O_1716,N_24832,N_24709);
or UO_1717 (O_1717,N_24503,N_24683);
or UO_1718 (O_1718,N_24872,N_24949);
nand UO_1719 (O_1719,N_24932,N_24786);
and UO_1720 (O_1720,N_24857,N_24758);
nand UO_1721 (O_1721,N_24771,N_24951);
or UO_1722 (O_1722,N_24936,N_24932);
nand UO_1723 (O_1723,N_24812,N_24945);
nor UO_1724 (O_1724,N_24754,N_24740);
xnor UO_1725 (O_1725,N_24946,N_24681);
and UO_1726 (O_1726,N_24701,N_24950);
nor UO_1727 (O_1727,N_24670,N_24839);
or UO_1728 (O_1728,N_24640,N_24595);
nor UO_1729 (O_1729,N_24505,N_24633);
or UO_1730 (O_1730,N_24933,N_24810);
nand UO_1731 (O_1731,N_24778,N_24521);
or UO_1732 (O_1732,N_24504,N_24583);
and UO_1733 (O_1733,N_24761,N_24781);
xnor UO_1734 (O_1734,N_24815,N_24760);
nand UO_1735 (O_1735,N_24697,N_24742);
nor UO_1736 (O_1736,N_24747,N_24639);
xnor UO_1737 (O_1737,N_24905,N_24845);
or UO_1738 (O_1738,N_24956,N_24502);
and UO_1739 (O_1739,N_24678,N_24702);
xnor UO_1740 (O_1740,N_24917,N_24789);
nor UO_1741 (O_1741,N_24622,N_24783);
nand UO_1742 (O_1742,N_24568,N_24719);
or UO_1743 (O_1743,N_24667,N_24707);
or UO_1744 (O_1744,N_24551,N_24514);
and UO_1745 (O_1745,N_24509,N_24781);
nor UO_1746 (O_1746,N_24939,N_24843);
or UO_1747 (O_1747,N_24510,N_24789);
and UO_1748 (O_1748,N_24888,N_24651);
and UO_1749 (O_1749,N_24615,N_24962);
xor UO_1750 (O_1750,N_24971,N_24564);
and UO_1751 (O_1751,N_24811,N_24972);
nor UO_1752 (O_1752,N_24548,N_24705);
xor UO_1753 (O_1753,N_24839,N_24563);
and UO_1754 (O_1754,N_24530,N_24661);
nand UO_1755 (O_1755,N_24802,N_24931);
nor UO_1756 (O_1756,N_24566,N_24561);
nor UO_1757 (O_1757,N_24744,N_24650);
nor UO_1758 (O_1758,N_24629,N_24813);
nor UO_1759 (O_1759,N_24962,N_24827);
xor UO_1760 (O_1760,N_24755,N_24738);
nand UO_1761 (O_1761,N_24899,N_24786);
nor UO_1762 (O_1762,N_24615,N_24612);
xor UO_1763 (O_1763,N_24624,N_24990);
xnor UO_1764 (O_1764,N_24860,N_24880);
or UO_1765 (O_1765,N_24563,N_24975);
nand UO_1766 (O_1766,N_24675,N_24672);
and UO_1767 (O_1767,N_24874,N_24562);
and UO_1768 (O_1768,N_24922,N_24978);
or UO_1769 (O_1769,N_24807,N_24908);
nor UO_1770 (O_1770,N_24916,N_24915);
xnor UO_1771 (O_1771,N_24933,N_24567);
xor UO_1772 (O_1772,N_24727,N_24855);
xor UO_1773 (O_1773,N_24585,N_24666);
nor UO_1774 (O_1774,N_24665,N_24742);
and UO_1775 (O_1775,N_24725,N_24604);
nor UO_1776 (O_1776,N_24652,N_24860);
and UO_1777 (O_1777,N_24569,N_24900);
nor UO_1778 (O_1778,N_24634,N_24924);
nand UO_1779 (O_1779,N_24928,N_24638);
xnor UO_1780 (O_1780,N_24686,N_24607);
or UO_1781 (O_1781,N_24659,N_24544);
nand UO_1782 (O_1782,N_24762,N_24665);
xnor UO_1783 (O_1783,N_24919,N_24560);
nor UO_1784 (O_1784,N_24928,N_24543);
nand UO_1785 (O_1785,N_24898,N_24846);
nand UO_1786 (O_1786,N_24675,N_24617);
xor UO_1787 (O_1787,N_24975,N_24645);
or UO_1788 (O_1788,N_24752,N_24970);
or UO_1789 (O_1789,N_24785,N_24636);
nand UO_1790 (O_1790,N_24594,N_24512);
xor UO_1791 (O_1791,N_24675,N_24798);
nand UO_1792 (O_1792,N_24604,N_24526);
or UO_1793 (O_1793,N_24920,N_24985);
nand UO_1794 (O_1794,N_24760,N_24692);
xnor UO_1795 (O_1795,N_24606,N_24698);
and UO_1796 (O_1796,N_24768,N_24848);
and UO_1797 (O_1797,N_24571,N_24936);
nand UO_1798 (O_1798,N_24623,N_24717);
or UO_1799 (O_1799,N_24580,N_24850);
or UO_1800 (O_1800,N_24559,N_24584);
xor UO_1801 (O_1801,N_24512,N_24824);
or UO_1802 (O_1802,N_24567,N_24901);
xnor UO_1803 (O_1803,N_24953,N_24590);
nand UO_1804 (O_1804,N_24748,N_24798);
nor UO_1805 (O_1805,N_24912,N_24881);
or UO_1806 (O_1806,N_24747,N_24929);
nand UO_1807 (O_1807,N_24502,N_24805);
or UO_1808 (O_1808,N_24820,N_24594);
and UO_1809 (O_1809,N_24777,N_24587);
xnor UO_1810 (O_1810,N_24904,N_24791);
and UO_1811 (O_1811,N_24872,N_24746);
nand UO_1812 (O_1812,N_24732,N_24703);
or UO_1813 (O_1813,N_24674,N_24965);
and UO_1814 (O_1814,N_24868,N_24806);
nor UO_1815 (O_1815,N_24650,N_24845);
nor UO_1816 (O_1816,N_24753,N_24859);
nor UO_1817 (O_1817,N_24774,N_24965);
nand UO_1818 (O_1818,N_24923,N_24513);
nand UO_1819 (O_1819,N_24929,N_24812);
nor UO_1820 (O_1820,N_24553,N_24771);
and UO_1821 (O_1821,N_24619,N_24826);
or UO_1822 (O_1822,N_24977,N_24567);
nor UO_1823 (O_1823,N_24980,N_24880);
xnor UO_1824 (O_1824,N_24584,N_24952);
nor UO_1825 (O_1825,N_24750,N_24739);
or UO_1826 (O_1826,N_24801,N_24650);
nor UO_1827 (O_1827,N_24500,N_24999);
and UO_1828 (O_1828,N_24956,N_24639);
nor UO_1829 (O_1829,N_24725,N_24549);
or UO_1830 (O_1830,N_24722,N_24708);
and UO_1831 (O_1831,N_24742,N_24920);
nand UO_1832 (O_1832,N_24822,N_24552);
nor UO_1833 (O_1833,N_24716,N_24937);
xnor UO_1834 (O_1834,N_24770,N_24937);
or UO_1835 (O_1835,N_24995,N_24872);
and UO_1836 (O_1836,N_24839,N_24638);
or UO_1837 (O_1837,N_24933,N_24577);
nor UO_1838 (O_1838,N_24935,N_24885);
or UO_1839 (O_1839,N_24947,N_24585);
or UO_1840 (O_1840,N_24557,N_24577);
nand UO_1841 (O_1841,N_24975,N_24983);
or UO_1842 (O_1842,N_24972,N_24635);
nor UO_1843 (O_1843,N_24901,N_24896);
nand UO_1844 (O_1844,N_24787,N_24673);
and UO_1845 (O_1845,N_24700,N_24528);
xor UO_1846 (O_1846,N_24915,N_24555);
nor UO_1847 (O_1847,N_24737,N_24787);
or UO_1848 (O_1848,N_24968,N_24607);
or UO_1849 (O_1849,N_24842,N_24745);
xor UO_1850 (O_1850,N_24789,N_24644);
or UO_1851 (O_1851,N_24621,N_24646);
and UO_1852 (O_1852,N_24762,N_24999);
xor UO_1853 (O_1853,N_24637,N_24708);
and UO_1854 (O_1854,N_24981,N_24860);
or UO_1855 (O_1855,N_24659,N_24914);
or UO_1856 (O_1856,N_24707,N_24635);
or UO_1857 (O_1857,N_24582,N_24800);
nor UO_1858 (O_1858,N_24573,N_24830);
xor UO_1859 (O_1859,N_24897,N_24775);
or UO_1860 (O_1860,N_24556,N_24672);
nor UO_1861 (O_1861,N_24576,N_24892);
and UO_1862 (O_1862,N_24635,N_24930);
or UO_1863 (O_1863,N_24628,N_24649);
and UO_1864 (O_1864,N_24682,N_24684);
and UO_1865 (O_1865,N_24916,N_24680);
and UO_1866 (O_1866,N_24591,N_24672);
xnor UO_1867 (O_1867,N_24915,N_24786);
and UO_1868 (O_1868,N_24798,N_24880);
nor UO_1869 (O_1869,N_24938,N_24720);
nor UO_1870 (O_1870,N_24625,N_24887);
or UO_1871 (O_1871,N_24753,N_24589);
nand UO_1872 (O_1872,N_24952,N_24678);
or UO_1873 (O_1873,N_24637,N_24611);
and UO_1874 (O_1874,N_24601,N_24689);
nand UO_1875 (O_1875,N_24809,N_24718);
nor UO_1876 (O_1876,N_24912,N_24771);
nand UO_1877 (O_1877,N_24946,N_24831);
xnor UO_1878 (O_1878,N_24519,N_24915);
xor UO_1879 (O_1879,N_24669,N_24799);
nor UO_1880 (O_1880,N_24566,N_24524);
nor UO_1881 (O_1881,N_24653,N_24839);
or UO_1882 (O_1882,N_24988,N_24648);
nor UO_1883 (O_1883,N_24549,N_24939);
nand UO_1884 (O_1884,N_24583,N_24802);
or UO_1885 (O_1885,N_24967,N_24702);
nor UO_1886 (O_1886,N_24723,N_24636);
and UO_1887 (O_1887,N_24649,N_24706);
nand UO_1888 (O_1888,N_24819,N_24980);
nor UO_1889 (O_1889,N_24906,N_24909);
xor UO_1890 (O_1890,N_24707,N_24751);
and UO_1891 (O_1891,N_24610,N_24775);
and UO_1892 (O_1892,N_24544,N_24598);
and UO_1893 (O_1893,N_24629,N_24889);
nand UO_1894 (O_1894,N_24971,N_24923);
and UO_1895 (O_1895,N_24904,N_24895);
nand UO_1896 (O_1896,N_24824,N_24846);
nor UO_1897 (O_1897,N_24961,N_24672);
xor UO_1898 (O_1898,N_24750,N_24582);
xor UO_1899 (O_1899,N_24988,N_24617);
xnor UO_1900 (O_1900,N_24611,N_24933);
nand UO_1901 (O_1901,N_24702,N_24754);
xor UO_1902 (O_1902,N_24922,N_24755);
or UO_1903 (O_1903,N_24832,N_24695);
nand UO_1904 (O_1904,N_24889,N_24530);
and UO_1905 (O_1905,N_24517,N_24877);
nand UO_1906 (O_1906,N_24735,N_24741);
or UO_1907 (O_1907,N_24693,N_24771);
and UO_1908 (O_1908,N_24828,N_24812);
and UO_1909 (O_1909,N_24737,N_24581);
or UO_1910 (O_1910,N_24778,N_24592);
xor UO_1911 (O_1911,N_24956,N_24513);
or UO_1912 (O_1912,N_24894,N_24977);
nand UO_1913 (O_1913,N_24659,N_24837);
or UO_1914 (O_1914,N_24749,N_24813);
or UO_1915 (O_1915,N_24851,N_24881);
or UO_1916 (O_1916,N_24848,N_24884);
nor UO_1917 (O_1917,N_24873,N_24965);
xnor UO_1918 (O_1918,N_24821,N_24775);
nor UO_1919 (O_1919,N_24752,N_24540);
xor UO_1920 (O_1920,N_24864,N_24960);
and UO_1921 (O_1921,N_24548,N_24845);
xnor UO_1922 (O_1922,N_24813,N_24880);
xor UO_1923 (O_1923,N_24726,N_24511);
nand UO_1924 (O_1924,N_24876,N_24734);
nand UO_1925 (O_1925,N_24612,N_24942);
nor UO_1926 (O_1926,N_24502,N_24580);
nor UO_1927 (O_1927,N_24782,N_24771);
or UO_1928 (O_1928,N_24514,N_24854);
or UO_1929 (O_1929,N_24905,N_24972);
xor UO_1930 (O_1930,N_24847,N_24531);
and UO_1931 (O_1931,N_24672,N_24716);
nand UO_1932 (O_1932,N_24805,N_24838);
and UO_1933 (O_1933,N_24843,N_24638);
or UO_1934 (O_1934,N_24610,N_24875);
nor UO_1935 (O_1935,N_24926,N_24813);
or UO_1936 (O_1936,N_24543,N_24604);
nand UO_1937 (O_1937,N_24602,N_24529);
and UO_1938 (O_1938,N_24935,N_24525);
or UO_1939 (O_1939,N_24962,N_24807);
nor UO_1940 (O_1940,N_24642,N_24825);
and UO_1941 (O_1941,N_24854,N_24927);
xnor UO_1942 (O_1942,N_24997,N_24778);
and UO_1943 (O_1943,N_24680,N_24600);
nand UO_1944 (O_1944,N_24875,N_24707);
xnor UO_1945 (O_1945,N_24803,N_24767);
nand UO_1946 (O_1946,N_24892,N_24500);
xor UO_1947 (O_1947,N_24572,N_24684);
xnor UO_1948 (O_1948,N_24916,N_24956);
or UO_1949 (O_1949,N_24957,N_24883);
and UO_1950 (O_1950,N_24918,N_24655);
nand UO_1951 (O_1951,N_24600,N_24916);
and UO_1952 (O_1952,N_24524,N_24884);
or UO_1953 (O_1953,N_24937,N_24500);
nor UO_1954 (O_1954,N_24694,N_24803);
and UO_1955 (O_1955,N_24903,N_24960);
nand UO_1956 (O_1956,N_24940,N_24650);
or UO_1957 (O_1957,N_24811,N_24806);
or UO_1958 (O_1958,N_24912,N_24699);
xnor UO_1959 (O_1959,N_24689,N_24873);
nor UO_1960 (O_1960,N_24943,N_24671);
nand UO_1961 (O_1961,N_24507,N_24857);
nand UO_1962 (O_1962,N_24686,N_24780);
and UO_1963 (O_1963,N_24786,N_24586);
or UO_1964 (O_1964,N_24507,N_24529);
nor UO_1965 (O_1965,N_24935,N_24730);
and UO_1966 (O_1966,N_24617,N_24794);
nand UO_1967 (O_1967,N_24957,N_24626);
or UO_1968 (O_1968,N_24686,N_24583);
xor UO_1969 (O_1969,N_24502,N_24534);
nor UO_1970 (O_1970,N_24684,N_24952);
xor UO_1971 (O_1971,N_24915,N_24762);
nand UO_1972 (O_1972,N_24830,N_24951);
and UO_1973 (O_1973,N_24885,N_24844);
or UO_1974 (O_1974,N_24877,N_24534);
nand UO_1975 (O_1975,N_24662,N_24907);
or UO_1976 (O_1976,N_24655,N_24965);
and UO_1977 (O_1977,N_24951,N_24859);
and UO_1978 (O_1978,N_24957,N_24951);
nand UO_1979 (O_1979,N_24713,N_24805);
xnor UO_1980 (O_1980,N_24722,N_24500);
and UO_1981 (O_1981,N_24989,N_24983);
or UO_1982 (O_1982,N_24819,N_24830);
nand UO_1983 (O_1983,N_24918,N_24555);
xor UO_1984 (O_1984,N_24967,N_24778);
and UO_1985 (O_1985,N_24511,N_24851);
nand UO_1986 (O_1986,N_24885,N_24988);
and UO_1987 (O_1987,N_24659,N_24623);
or UO_1988 (O_1988,N_24952,N_24529);
and UO_1989 (O_1989,N_24689,N_24811);
or UO_1990 (O_1990,N_24981,N_24587);
xor UO_1991 (O_1991,N_24941,N_24528);
nor UO_1992 (O_1992,N_24947,N_24566);
or UO_1993 (O_1993,N_24745,N_24530);
xnor UO_1994 (O_1994,N_24694,N_24615);
and UO_1995 (O_1995,N_24714,N_24877);
or UO_1996 (O_1996,N_24802,N_24574);
and UO_1997 (O_1997,N_24625,N_24838);
nor UO_1998 (O_1998,N_24924,N_24632);
nand UO_1999 (O_1999,N_24553,N_24662);
or UO_2000 (O_2000,N_24895,N_24514);
xnor UO_2001 (O_2001,N_24752,N_24621);
nand UO_2002 (O_2002,N_24994,N_24903);
nor UO_2003 (O_2003,N_24961,N_24907);
nor UO_2004 (O_2004,N_24573,N_24878);
xnor UO_2005 (O_2005,N_24524,N_24875);
nand UO_2006 (O_2006,N_24857,N_24572);
nand UO_2007 (O_2007,N_24996,N_24777);
or UO_2008 (O_2008,N_24966,N_24901);
or UO_2009 (O_2009,N_24660,N_24766);
xor UO_2010 (O_2010,N_24860,N_24986);
xnor UO_2011 (O_2011,N_24629,N_24683);
xor UO_2012 (O_2012,N_24597,N_24513);
and UO_2013 (O_2013,N_24979,N_24973);
xor UO_2014 (O_2014,N_24829,N_24660);
nand UO_2015 (O_2015,N_24600,N_24701);
xnor UO_2016 (O_2016,N_24819,N_24907);
nand UO_2017 (O_2017,N_24503,N_24671);
or UO_2018 (O_2018,N_24955,N_24536);
or UO_2019 (O_2019,N_24968,N_24621);
and UO_2020 (O_2020,N_24552,N_24937);
and UO_2021 (O_2021,N_24847,N_24687);
or UO_2022 (O_2022,N_24629,N_24681);
nor UO_2023 (O_2023,N_24675,N_24795);
or UO_2024 (O_2024,N_24844,N_24719);
xor UO_2025 (O_2025,N_24656,N_24847);
and UO_2026 (O_2026,N_24986,N_24512);
nor UO_2027 (O_2027,N_24614,N_24829);
xnor UO_2028 (O_2028,N_24560,N_24742);
xor UO_2029 (O_2029,N_24929,N_24797);
and UO_2030 (O_2030,N_24583,N_24752);
and UO_2031 (O_2031,N_24686,N_24613);
or UO_2032 (O_2032,N_24569,N_24614);
or UO_2033 (O_2033,N_24796,N_24885);
xor UO_2034 (O_2034,N_24982,N_24941);
and UO_2035 (O_2035,N_24788,N_24573);
or UO_2036 (O_2036,N_24963,N_24840);
and UO_2037 (O_2037,N_24507,N_24655);
and UO_2038 (O_2038,N_24699,N_24598);
or UO_2039 (O_2039,N_24997,N_24553);
and UO_2040 (O_2040,N_24979,N_24926);
nand UO_2041 (O_2041,N_24850,N_24691);
and UO_2042 (O_2042,N_24610,N_24721);
nand UO_2043 (O_2043,N_24546,N_24615);
and UO_2044 (O_2044,N_24677,N_24754);
nor UO_2045 (O_2045,N_24597,N_24909);
or UO_2046 (O_2046,N_24830,N_24529);
xor UO_2047 (O_2047,N_24967,N_24732);
xnor UO_2048 (O_2048,N_24634,N_24598);
xor UO_2049 (O_2049,N_24764,N_24778);
xor UO_2050 (O_2050,N_24767,N_24824);
nand UO_2051 (O_2051,N_24695,N_24839);
nor UO_2052 (O_2052,N_24820,N_24994);
nand UO_2053 (O_2053,N_24712,N_24532);
nor UO_2054 (O_2054,N_24595,N_24530);
or UO_2055 (O_2055,N_24538,N_24701);
xor UO_2056 (O_2056,N_24880,N_24782);
or UO_2057 (O_2057,N_24676,N_24697);
nor UO_2058 (O_2058,N_24715,N_24888);
nand UO_2059 (O_2059,N_24606,N_24971);
nor UO_2060 (O_2060,N_24601,N_24836);
nand UO_2061 (O_2061,N_24660,N_24657);
xor UO_2062 (O_2062,N_24978,N_24873);
nand UO_2063 (O_2063,N_24552,N_24885);
nand UO_2064 (O_2064,N_24586,N_24847);
nor UO_2065 (O_2065,N_24539,N_24766);
or UO_2066 (O_2066,N_24955,N_24523);
nand UO_2067 (O_2067,N_24944,N_24692);
nor UO_2068 (O_2068,N_24790,N_24653);
nor UO_2069 (O_2069,N_24810,N_24860);
or UO_2070 (O_2070,N_24656,N_24814);
nor UO_2071 (O_2071,N_24791,N_24533);
or UO_2072 (O_2072,N_24688,N_24778);
or UO_2073 (O_2073,N_24832,N_24811);
nor UO_2074 (O_2074,N_24638,N_24630);
nand UO_2075 (O_2075,N_24769,N_24562);
or UO_2076 (O_2076,N_24824,N_24658);
or UO_2077 (O_2077,N_24799,N_24736);
and UO_2078 (O_2078,N_24589,N_24714);
nor UO_2079 (O_2079,N_24754,N_24611);
nor UO_2080 (O_2080,N_24666,N_24777);
or UO_2081 (O_2081,N_24699,N_24731);
nor UO_2082 (O_2082,N_24981,N_24522);
and UO_2083 (O_2083,N_24551,N_24708);
nand UO_2084 (O_2084,N_24771,N_24689);
xor UO_2085 (O_2085,N_24953,N_24712);
or UO_2086 (O_2086,N_24682,N_24748);
and UO_2087 (O_2087,N_24725,N_24921);
or UO_2088 (O_2088,N_24966,N_24977);
or UO_2089 (O_2089,N_24543,N_24634);
xor UO_2090 (O_2090,N_24546,N_24622);
xnor UO_2091 (O_2091,N_24632,N_24662);
nor UO_2092 (O_2092,N_24861,N_24525);
nor UO_2093 (O_2093,N_24880,N_24585);
and UO_2094 (O_2094,N_24999,N_24970);
and UO_2095 (O_2095,N_24508,N_24920);
nand UO_2096 (O_2096,N_24512,N_24853);
xor UO_2097 (O_2097,N_24933,N_24952);
nand UO_2098 (O_2098,N_24871,N_24557);
nor UO_2099 (O_2099,N_24962,N_24571);
nor UO_2100 (O_2100,N_24712,N_24694);
or UO_2101 (O_2101,N_24737,N_24507);
xnor UO_2102 (O_2102,N_24783,N_24905);
nor UO_2103 (O_2103,N_24720,N_24547);
or UO_2104 (O_2104,N_24901,N_24599);
and UO_2105 (O_2105,N_24681,N_24545);
and UO_2106 (O_2106,N_24542,N_24749);
xor UO_2107 (O_2107,N_24833,N_24874);
and UO_2108 (O_2108,N_24659,N_24644);
xor UO_2109 (O_2109,N_24566,N_24516);
xnor UO_2110 (O_2110,N_24973,N_24913);
and UO_2111 (O_2111,N_24679,N_24988);
xnor UO_2112 (O_2112,N_24634,N_24960);
and UO_2113 (O_2113,N_24644,N_24858);
or UO_2114 (O_2114,N_24849,N_24534);
xor UO_2115 (O_2115,N_24815,N_24977);
nand UO_2116 (O_2116,N_24965,N_24559);
or UO_2117 (O_2117,N_24689,N_24540);
and UO_2118 (O_2118,N_24967,N_24555);
nand UO_2119 (O_2119,N_24606,N_24650);
and UO_2120 (O_2120,N_24703,N_24841);
nor UO_2121 (O_2121,N_24844,N_24715);
or UO_2122 (O_2122,N_24858,N_24995);
nor UO_2123 (O_2123,N_24581,N_24513);
nor UO_2124 (O_2124,N_24540,N_24632);
nor UO_2125 (O_2125,N_24873,N_24976);
nand UO_2126 (O_2126,N_24704,N_24538);
and UO_2127 (O_2127,N_24801,N_24566);
and UO_2128 (O_2128,N_24546,N_24599);
xor UO_2129 (O_2129,N_24501,N_24881);
nor UO_2130 (O_2130,N_24683,N_24630);
nor UO_2131 (O_2131,N_24950,N_24896);
nand UO_2132 (O_2132,N_24853,N_24786);
and UO_2133 (O_2133,N_24807,N_24877);
or UO_2134 (O_2134,N_24611,N_24642);
or UO_2135 (O_2135,N_24874,N_24544);
nand UO_2136 (O_2136,N_24564,N_24643);
or UO_2137 (O_2137,N_24859,N_24660);
and UO_2138 (O_2138,N_24784,N_24644);
or UO_2139 (O_2139,N_24766,N_24975);
nand UO_2140 (O_2140,N_24839,N_24762);
nand UO_2141 (O_2141,N_24728,N_24983);
and UO_2142 (O_2142,N_24706,N_24672);
nor UO_2143 (O_2143,N_24529,N_24593);
and UO_2144 (O_2144,N_24883,N_24510);
xnor UO_2145 (O_2145,N_24893,N_24527);
nor UO_2146 (O_2146,N_24525,N_24877);
and UO_2147 (O_2147,N_24917,N_24742);
and UO_2148 (O_2148,N_24557,N_24520);
nor UO_2149 (O_2149,N_24596,N_24957);
or UO_2150 (O_2150,N_24689,N_24657);
and UO_2151 (O_2151,N_24979,N_24982);
xnor UO_2152 (O_2152,N_24962,N_24502);
or UO_2153 (O_2153,N_24863,N_24931);
nor UO_2154 (O_2154,N_24516,N_24800);
nor UO_2155 (O_2155,N_24902,N_24975);
xnor UO_2156 (O_2156,N_24850,N_24627);
or UO_2157 (O_2157,N_24783,N_24966);
and UO_2158 (O_2158,N_24564,N_24850);
nor UO_2159 (O_2159,N_24725,N_24724);
nor UO_2160 (O_2160,N_24868,N_24592);
or UO_2161 (O_2161,N_24938,N_24998);
or UO_2162 (O_2162,N_24552,N_24832);
xnor UO_2163 (O_2163,N_24875,N_24683);
nor UO_2164 (O_2164,N_24849,N_24958);
xnor UO_2165 (O_2165,N_24961,N_24896);
and UO_2166 (O_2166,N_24805,N_24735);
and UO_2167 (O_2167,N_24790,N_24608);
and UO_2168 (O_2168,N_24546,N_24872);
xnor UO_2169 (O_2169,N_24963,N_24522);
xnor UO_2170 (O_2170,N_24632,N_24824);
xor UO_2171 (O_2171,N_24594,N_24804);
nand UO_2172 (O_2172,N_24897,N_24667);
or UO_2173 (O_2173,N_24578,N_24771);
nand UO_2174 (O_2174,N_24978,N_24617);
xnor UO_2175 (O_2175,N_24967,N_24817);
nor UO_2176 (O_2176,N_24906,N_24500);
nor UO_2177 (O_2177,N_24616,N_24968);
and UO_2178 (O_2178,N_24564,N_24634);
and UO_2179 (O_2179,N_24843,N_24879);
and UO_2180 (O_2180,N_24646,N_24596);
nand UO_2181 (O_2181,N_24748,N_24672);
or UO_2182 (O_2182,N_24927,N_24925);
or UO_2183 (O_2183,N_24994,N_24768);
nor UO_2184 (O_2184,N_24507,N_24911);
and UO_2185 (O_2185,N_24566,N_24682);
nor UO_2186 (O_2186,N_24912,N_24895);
nand UO_2187 (O_2187,N_24699,N_24736);
nand UO_2188 (O_2188,N_24764,N_24784);
xnor UO_2189 (O_2189,N_24519,N_24813);
nand UO_2190 (O_2190,N_24740,N_24711);
nor UO_2191 (O_2191,N_24879,N_24611);
xnor UO_2192 (O_2192,N_24689,N_24984);
xnor UO_2193 (O_2193,N_24840,N_24568);
or UO_2194 (O_2194,N_24834,N_24955);
xnor UO_2195 (O_2195,N_24962,N_24762);
nand UO_2196 (O_2196,N_24718,N_24698);
xor UO_2197 (O_2197,N_24772,N_24784);
xnor UO_2198 (O_2198,N_24621,N_24978);
and UO_2199 (O_2199,N_24586,N_24585);
and UO_2200 (O_2200,N_24573,N_24976);
nand UO_2201 (O_2201,N_24834,N_24892);
nor UO_2202 (O_2202,N_24684,N_24975);
nor UO_2203 (O_2203,N_24783,N_24943);
or UO_2204 (O_2204,N_24955,N_24527);
xor UO_2205 (O_2205,N_24710,N_24760);
xor UO_2206 (O_2206,N_24775,N_24680);
nor UO_2207 (O_2207,N_24776,N_24613);
or UO_2208 (O_2208,N_24592,N_24830);
nor UO_2209 (O_2209,N_24855,N_24988);
and UO_2210 (O_2210,N_24844,N_24555);
or UO_2211 (O_2211,N_24765,N_24917);
xnor UO_2212 (O_2212,N_24989,N_24633);
nor UO_2213 (O_2213,N_24652,N_24793);
or UO_2214 (O_2214,N_24687,N_24915);
nor UO_2215 (O_2215,N_24740,N_24871);
nor UO_2216 (O_2216,N_24916,N_24986);
nor UO_2217 (O_2217,N_24594,N_24913);
or UO_2218 (O_2218,N_24940,N_24538);
and UO_2219 (O_2219,N_24657,N_24900);
or UO_2220 (O_2220,N_24614,N_24636);
nor UO_2221 (O_2221,N_24949,N_24564);
and UO_2222 (O_2222,N_24740,N_24771);
nand UO_2223 (O_2223,N_24764,N_24766);
or UO_2224 (O_2224,N_24992,N_24740);
nor UO_2225 (O_2225,N_24732,N_24539);
and UO_2226 (O_2226,N_24919,N_24591);
nand UO_2227 (O_2227,N_24901,N_24831);
nor UO_2228 (O_2228,N_24902,N_24552);
and UO_2229 (O_2229,N_24968,N_24790);
nand UO_2230 (O_2230,N_24826,N_24835);
nand UO_2231 (O_2231,N_24818,N_24531);
and UO_2232 (O_2232,N_24750,N_24941);
xor UO_2233 (O_2233,N_24885,N_24560);
nor UO_2234 (O_2234,N_24571,N_24952);
xor UO_2235 (O_2235,N_24917,N_24721);
xor UO_2236 (O_2236,N_24779,N_24924);
or UO_2237 (O_2237,N_24861,N_24826);
xor UO_2238 (O_2238,N_24880,N_24687);
nor UO_2239 (O_2239,N_24771,N_24908);
nor UO_2240 (O_2240,N_24816,N_24647);
nand UO_2241 (O_2241,N_24669,N_24968);
and UO_2242 (O_2242,N_24770,N_24714);
and UO_2243 (O_2243,N_24847,N_24953);
nor UO_2244 (O_2244,N_24937,N_24865);
nor UO_2245 (O_2245,N_24615,N_24744);
nor UO_2246 (O_2246,N_24574,N_24866);
nand UO_2247 (O_2247,N_24974,N_24627);
and UO_2248 (O_2248,N_24745,N_24978);
xnor UO_2249 (O_2249,N_24762,N_24946);
and UO_2250 (O_2250,N_24669,N_24986);
xnor UO_2251 (O_2251,N_24997,N_24886);
xnor UO_2252 (O_2252,N_24968,N_24776);
xnor UO_2253 (O_2253,N_24908,N_24945);
nor UO_2254 (O_2254,N_24571,N_24799);
or UO_2255 (O_2255,N_24825,N_24820);
or UO_2256 (O_2256,N_24828,N_24610);
xnor UO_2257 (O_2257,N_24842,N_24758);
nor UO_2258 (O_2258,N_24525,N_24835);
nor UO_2259 (O_2259,N_24991,N_24588);
nand UO_2260 (O_2260,N_24547,N_24557);
xor UO_2261 (O_2261,N_24695,N_24824);
nand UO_2262 (O_2262,N_24825,N_24599);
and UO_2263 (O_2263,N_24602,N_24672);
nor UO_2264 (O_2264,N_24724,N_24810);
and UO_2265 (O_2265,N_24792,N_24796);
and UO_2266 (O_2266,N_24861,N_24533);
or UO_2267 (O_2267,N_24616,N_24614);
nand UO_2268 (O_2268,N_24682,N_24713);
and UO_2269 (O_2269,N_24952,N_24946);
nand UO_2270 (O_2270,N_24913,N_24777);
nand UO_2271 (O_2271,N_24865,N_24862);
and UO_2272 (O_2272,N_24667,N_24758);
xor UO_2273 (O_2273,N_24755,N_24977);
xor UO_2274 (O_2274,N_24607,N_24646);
xnor UO_2275 (O_2275,N_24870,N_24607);
xnor UO_2276 (O_2276,N_24843,N_24636);
or UO_2277 (O_2277,N_24916,N_24862);
nor UO_2278 (O_2278,N_24787,N_24759);
nand UO_2279 (O_2279,N_24752,N_24698);
nand UO_2280 (O_2280,N_24892,N_24995);
nor UO_2281 (O_2281,N_24672,N_24571);
xnor UO_2282 (O_2282,N_24946,N_24898);
nor UO_2283 (O_2283,N_24547,N_24822);
nor UO_2284 (O_2284,N_24937,N_24999);
nand UO_2285 (O_2285,N_24505,N_24706);
xnor UO_2286 (O_2286,N_24745,N_24736);
nand UO_2287 (O_2287,N_24886,N_24923);
and UO_2288 (O_2288,N_24938,N_24929);
nand UO_2289 (O_2289,N_24552,N_24645);
or UO_2290 (O_2290,N_24656,N_24562);
nor UO_2291 (O_2291,N_24781,N_24892);
and UO_2292 (O_2292,N_24773,N_24963);
and UO_2293 (O_2293,N_24892,N_24592);
nand UO_2294 (O_2294,N_24835,N_24962);
xor UO_2295 (O_2295,N_24988,N_24999);
and UO_2296 (O_2296,N_24627,N_24806);
or UO_2297 (O_2297,N_24544,N_24501);
nand UO_2298 (O_2298,N_24603,N_24526);
nor UO_2299 (O_2299,N_24597,N_24760);
and UO_2300 (O_2300,N_24801,N_24685);
nor UO_2301 (O_2301,N_24927,N_24891);
and UO_2302 (O_2302,N_24954,N_24891);
nor UO_2303 (O_2303,N_24961,N_24517);
nor UO_2304 (O_2304,N_24558,N_24567);
nor UO_2305 (O_2305,N_24742,N_24829);
or UO_2306 (O_2306,N_24742,N_24551);
nor UO_2307 (O_2307,N_24606,N_24667);
or UO_2308 (O_2308,N_24859,N_24942);
nor UO_2309 (O_2309,N_24887,N_24568);
nand UO_2310 (O_2310,N_24812,N_24840);
xnor UO_2311 (O_2311,N_24579,N_24907);
nand UO_2312 (O_2312,N_24640,N_24995);
and UO_2313 (O_2313,N_24948,N_24617);
or UO_2314 (O_2314,N_24576,N_24678);
or UO_2315 (O_2315,N_24978,N_24892);
or UO_2316 (O_2316,N_24745,N_24847);
and UO_2317 (O_2317,N_24557,N_24760);
and UO_2318 (O_2318,N_24905,N_24526);
or UO_2319 (O_2319,N_24526,N_24988);
nor UO_2320 (O_2320,N_24547,N_24941);
and UO_2321 (O_2321,N_24571,N_24776);
nor UO_2322 (O_2322,N_24844,N_24828);
or UO_2323 (O_2323,N_24688,N_24917);
and UO_2324 (O_2324,N_24798,N_24565);
or UO_2325 (O_2325,N_24582,N_24922);
xnor UO_2326 (O_2326,N_24536,N_24825);
nor UO_2327 (O_2327,N_24944,N_24587);
or UO_2328 (O_2328,N_24783,N_24765);
nor UO_2329 (O_2329,N_24728,N_24518);
or UO_2330 (O_2330,N_24517,N_24928);
xnor UO_2331 (O_2331,N_24893,N_24914);
or UO_2332 (O_2332,N_24975,N_24923);
nor UO_2333 (O_2333,N_24767,N_24553);
and UO_2334 (O_2334,N_24590,N_24990);
xnor UO_2335 (O_2335,N_24701,N_24837);
or UO_2336 (O_2336,N_24535,N_24899);
and UO_2337 (O_2337,N_24686,N_24880);
nor UO_2338 (O_2338,N_24836,N_24544);
nand UO_2339 (O_2339,N_24955,N_24766);
nand UO_2340 (O_2340,N_24561,N_24801);
nor UO_2341 (O_2341,N_24661,N_24748);
or UO_2342 (O_2342,N_24612,N_24912);
or UO_2343 (O_2343,N_24932,N_24752);
or UO_2344 (O_2344,N_24699,N_24730);
and UO_2345 (O_2345,N_24553,N_24541);
and UO_2346 (O_2346,N_24602,N_24820);
nor UO_2347 (O_2347,N_24652,N_24861);
nor UO_2348 (O_2348,N_24976,N_24775);
xor UO_2349 (O_2349,N_24864,N_24875);
and UO_2350 (O_2350,N_24972,N_24657);
nor UO_2351 (O_2351,N_24756,N_24596);
or UO_2352 (O_2352,N_24756,N_24998);
nor UO_2353 (O_2353,N_24575,N_24921);
or UO_2354 (O_2354,N_24934,N_24592);
nor UO_2355 (O_2355,N_24820,N_24930);
nand UO_2356 (O_2356,N_24788,N_24586);
or UO_2357 (O_2357,N_24571,N_24622);
and UO_2358 (O_2358,N_24925,N_24505);
or UO_2359 (O_2359,N_24646,N_24744);
and UO_2360 (O_2360,N_24709,N_24826);
nor UO_2361 (O_2361,N_24524,N_24990);
nand UO_2362 (O_2362,N_24511,N_24873);
nand UO_2363 (O_2363,N_24679,N_24695);
nor UO_2364 (O_2364,N_24711,N_24929);
nor UO_2365 (O_2365,N_24813,N_24809);
nand UO_2366 (O_2366,N_24588,N_24605);
nand UO_2367 (O_2367,N_24865,N_24541);
nand UO_2368 (O_2368,N_24959,N_24698);
xor UO_2369 (O_2369,N_24750,N_24619);
nor UO_2370 (O_2370,N_24630,N_24926);
nand UO_2371 (O_2371,N_24636,N_24768);
and UO_2372 (O_2372,N_24630,N_24579);
and UO_2373 (O_2373,N_24735,N_24718);
xnor UO_2374 (O_2374,N_24520,N_24780);
or UO_2375 (O_2375,N_24581,N_24642);
or UO_2376 (O_2376,N_24729,N_24969);
and UO_2377 (O_2377,N_24732,N_24536);
or UO_2378 (O_2378,N_24847,N_24699);
or UO_2379 (O_2379,N_24865,N_24716);
nand UO_2380 (O_2380,N_24796,N_24719);
nand UO_2381 (O_2381,N_24537,N_24755);
or UO_2382 (O_2382,N_24677,N_24648);
nand UO_2383 (O_2383,N_24792,N_24625);
and UO_2384 (O_2384,N_24558,N_24847);
nand UO_2385 (O_2385,N_24606,N_24562);
xnor UO_2386 (O_2386,N_24700,N_24824);
nor UO_2387 (O_2387,N_24760,N_24962);
and UO_2388 (O_2388,N_24754,N_24596);
and UO_2389 (O_2389,N_24626,N_24900);
or UO_2390 (O_2390,N_24524,N_24887);
xor UO_2391 (O_2391,N_24997,N_24779);
nand UO_2392 (O_2392,N_24560,N_24877);
xor UO_2393 (O_2393,N_24851,N_24779);
and UO_2394 (O_2394,N_24578,N_24963);
nand UO_2395 (O_2395,N_24693,N_24657);
and UO_2396 (O_2396,N_24864,N_24665);
xor UO_2397 (O_2397,N_24583,N_24788);
nor UO_2398 (O_2398,N_24618,N_24573);
xnor UO_2399 (O_2399,N_24531,N_24511);
nand UO_2400 (O_2400,N_24596,N_24889);
xnor UO_2401 (O_2401,N_24837,N_24869);
nand UO_2402 (O_2402,N_24947,N_24773);
nor UO_2403 (O_2403,N_24841,N_24509);
nand UO_2404 (O_2404,N_24961,N_24810);
xnor UO_2405 (O_2405,N_24637,N_24533);
or UO_2406 (O_2406,N_24723,N_24825);
or UO_2407 (O_2407,N_24770,N_24735);
or UO_2408 (O_2408,N_24842,N_24875);
nand UO_2409 (O_2409,N_24710,N_24639);
and UO_2410 (O_2410,N_24628,N_24560);
and UO_2411 (O_2411,N_24581,N_24815);
and UO_2412 (O_2412,N_24962,N_24577);
nand UO_2413 (O_2413,N_24987,N_24574);
nand UO_2414 (O_2414,N_24547,N_24577);
and UO_2415 (O_2415,N_24820,N_24520);
nand UO_2416 (O_2416,N_24864,N_24717);
nor UO_2417 (O_2417,N_24758,N_24676);
nand UO_2418 (O_2418,N_24516,N_24998);
and UO_2419 (O_2419,N_24546,N_24841);
nand UO_2420 (O_2420,N_24501,N_24560);
or UO_2421 (O_2421,N_24546,N_24953);
and UO_2422 (O_2422,N_24636,N_24904);
nand UO_2423 (O_2423,N_24522,N_24771);
and UO_2424 (O_2424,N_24675,N_24578);
nor UO_2425 (O_2425,N_24916,N_24882);
or UO_2426 (O_2426,N_24580,N_24588);
nand UO_2427 (O_2427,N_24944,N_24772);
and UO_2428 (O_2428,N_24611,N_24963);
and UO_2429 (O_2429,N_24629,N_24950);
nand UO_2430 (O_2430,N_24711,N_24798);
and UO_2431 (O_2431,N_24730,N_24644);
and UO_2432 (O_2432,N_24574,N_24799);
xnor UO_2433 (O_2433,N_24962,N_24928);
xnor UO_2434 (O_2434,N_24757,N_24649);
nand UO_2435 (O_2435,N_24809,N_24954);
nand UO_2436 (O_2436,N_24554,N_24881);
or UO_2437 (O_2437,N_24972,N_24508);
or UO_2438 (O_2438,N_24805,N_24861);
and UO_2439 (O_2439,N_24926,N_24614);
or UO_2440 (O_2440,N_24915,N_24798);
xnor UO_2441 (O_2441,N_24587,N_24679);
or UO_2442 (O_2442,N_24573,N_24599);
nand UO_2443 (O_2443,N_24583,N_24807);
nor UO_2444 (O_2444,N_24583,N_24801);
nand UO_2445 (O_2445,N_24738,N_24979);
and UO_2446 (O_2446,N_24617,N_24946);
and UO_2447 (O_2447,N_24505,N_24888);
nand UO_2448 (O_2448,N_24927,N_24572);
nand UO_2449 (O_2449,N_24874,N_24936);
and UO_2450 (O_2450,N_24933,N_24697);
nand UO_2451 (O_2451,N_24503,N_24685);
nand UO_2452 (O_2452,N_24972,N_24910);
and UO_2453 (O_2453,N_24812,N_24800);
xnor UO_2454 (O_2454,N_24847,N_24911);
nand UO_2455 (O_2455,N_24792,N_24986);
nand UO_2456 (O_2456,N_24677,N_24675);
and UO_2457 (O_2457,N_24719,N_24569);
nand UO_2458 (O_2458,N_24558,N_24798);
xnor UO_2459 (O_2459,N_24679,N_24756);
nand UO_2460 (O_2460,N_24572,N_24633);
and UO_2461 (O_2461,N_24959,N_24780);
or UO_2462 (O_2462,N_24760,N_24755);
xor UO_2463 (O_2463,N_24802,N_24596);
nor UO_2464 (O_2464,N_24750,N_24650);
xnor UO_2465 (O_2465,N_24623,N_24675);
and UO_2466 (O_2466,N_24573,N_24574);
and UO_2467 (O_2467,N_24667,N_24933);
or UO_2468 (O_2468,N_24630,N_24892);
and UO_2469 (O_2469,N_24688,N_24586);
nand UO_2470 (O_2470,N_24717,N_24861);
xor UO_2471 (O_2471,N_24621,N_24566);
xnor UO_2472 (O_2472,N_24606,N_24569);
and UO_2473 (O_2473,N_24964,N_24744);
xnor UO_2474 (O_2474,N_24900,N_24683);
nor UO_2475 (O_2475,N_24706,N_24632);
or UO_2476 (O_2476,N_24843,N_24589);
nand UO_2477 (O_2477,N_24649,N_24872);
and UO_2478 (O_2478,N_24739,N_24940);
and UO_2479 (O_2479,N_24966,N_24517);
and UO_2480 (O_2480,N_24651,N_24589);
nand UO_2481 (O_2481,N_24694,N_24962);
nand UO_2482 (O_2482,N_24994,N_24853);
or UO_2483 (O_2483,N_24562,N_24640);
nand UO_2484 (O_2484,N_24506,N_24813);
nor UO_2485 (O_2485,N_24783,N_24593);
xor UO_2486 (O_2486,N_24546,N_24978);
xnor UO_2487 (O_2487,N_24610,N_24827);
nor UO_2488 (O_2488,N_24548,N_24919);
nor UO_2489 (O_2489,N_24905,N_24916);
and UO_2490 (O_2490,N_24661,N_24820);
or UO_2491 (O_2491,N_24742,N_24653);
nand UO_2492 (O_2492,N_24897,N_24747);
and UO_2493 (O_2493,N_24919,N_24564);
xor UO_2494 (O_2494,N_24521,N_24720);
xor UO_2495 (O_2495,N_24768,N_24912);
and UO_2496 (O_2496,N_24525,N_24727);
nor UO_2497 (O_2497,N_24718,N_24559);
xnor UO_2498 (O_2498,N_24866,N_24582);
nand UO_2499 (O_2499,N_24946,N_24595);
xor UO_2500 (O_2500,N_24526,N_24585);
and UO_2501 (O_2501,N_24825,N_24813);
and UO_2502 (O_2502,N_24692,N_24889);
nand UO_2503 (O_2503,N_24866,N_24516);
and UO_2504 (O_2504,N_24909,N_24919);
nand UO_2505 (O_2505,N_24576,N_24548);
nand UO_2506 (O_2506,N_24833,N_24557);
nor UO_2507 (O_2507,N_24878,N_24535);
nand UO_2508 (O_2508,N_24558,N_24892);
or UO_2509 (O_2509,N_24658,N_24730);
and UO_2510 (O_2510,N_24641,N_24587);
and UO_2511 (O_2511,N_24830,N_24753);
nor UO_2512 (O_2512,N_24708,N_24542);
nor UO_2513 (O_2513,N_24774,N_24740);
xor UO_2514 (O_2514,N_24733,N_24720);
nand UO_2515 (O_2515,N_24979,N_24726);
nand UO_2516 (O_2516,N_24820,N_24560);
and UO_2517 (O_2517,N_24644,N_24771);
nand UO_2518 (O_2518,N_24651,N_24535);
nand UO_2519 (O_2519,N_24689,N_24846);
nor UO_2520 (O_2520,N_24908,N_24987);
xnor UO_2521 (O_2521,N_24544,N_24507);
nand UO_2522 (O_2522,N_24882,N_24780);
or UO_2523 (O_2523,N_24893,N_24854);
nand UO_2524 (O_2524,N_24634,N_24867);
or UO_2525 (O_2525,N_24762,N_24861);
nor UO_2526 (O_2526,N_24922,N_24690);
or UO_2527 (O_2527,N_24696,N_24991);
xor UO_2528 (O_2528,N_24860,N_24765);
nand UO_2529 (O_2529,N_24599,N_24526);
nand UO_2530 (O_2530,N_24864,N_24842);
or UO_2531 (O_2531,N_24558,N_24622);
and UO_2532 (O_2532,N_24897,N_24657);
and UO_2533 (O_2533,N_24619,N_24558);
or UO_2534 (O_2534,N_24589,N_24706);
nor UO_2535 (O_2535,N_24871,N_24698);
nand UO_2536 (O_2536,N_24855,N_24623);
nor UO_2537 (O_2537,N_24912,N_24659);
and UO_2538 (O_2538,N_24513,N_24511);
or UO_2539 (O_2539,N_24661,N_24699);
or UO_2540 (O_2540,N_24631,N_24615);
xnor UO_2541 (O_2541,N_24671,N_24868);
xor UO_2542 (O_2542,N_24900,N_24732);
and UO_2543 (O_2543,N_24652,N_24963);
nand UO_2544 (O_2544,N_24923,N_24701);
xnor UO_2545 (O_2545,N_24873,N_24954);
xor UO_2546 (O_2546,N_24911,N_24868);
nor UO_2547 (O_2547,N_24775,N_24711);
and UO_2548 (O_2548,N_24828,N_24984);
and UO_2549 (O_2549,N_24982,N_24608);
and UO_2550 (O_2550,N_24983,N_24949);
nand UO_2551 (O_2551,N_24762,N_24880);
or UO_2552 (O_2552,N_24878,N_24797);
or UO_2553 (O_2553,N_24609,N_24615);
nor UO_2554 (O_2554,N_24640,N_24969);
nand UO_2555 (O_2555,N_24929,N_24830);
and UO_2556 (O_2556,N_24876,N_24728);
or UO_2557 (O_2557,N_24547,N_24649);
or UO_2558 (O_2558,N_24543,N_24775);
xnor UO_2559 (O_2559,N_24899,N_24987);
or UO_2560 (O_2560,N_24694,N_24935);
nor UO_2561 (O_2561,N_24552,N_24592);
nand UO_2562 (O_2562,N_24815,N_24646);
nor UO_2563 (O_2563,N_24720,N_24965);
nand UO_2564 (O_2564,N_24577,N_24972);
nand UO_2565 (O_2565,N_24501,N_24758);
nor UO_2566 (O_2566,N_24782,N_24524);
nand UO_2567 (O_2567,N_24744,N_24552);
xnor UO_2568 (O_2568,N_24980,N_24686);
and UO_2569 (O_2569,N_24997,N_24991);
nor UO_2570 (O_2570,N_24636,N_24613);
xor UO_2571 (O_2571,N_24688,N_24892);
xor UO_2572 (O_2572,N_24852,N_24750);
nor UO_2573 (O_2573,N_24561,N_24742);
nand UO_2574 (O_2574,N_24963,N_24651);
nor UO_2575 (O_2575,N_24804,N_24771);
nand UO_2576 (O_2576,N_24646,N_24884);
and UO_2577 (O_2577,N_24660,N_24512);
nor UO_2578 (O_2578,N_24815,N_24551);
xor UO_2579 (O_2579,N_24976,N_24941);
or UO_2580 (O_2580,N_24573,N_24846);
and UO_2581 (O_2581,N_24528,N_24844);
nor UO_2582 (O_2582,N_24700,N_24975);
and UO_2583 (O_2583,N_24942,N_24934);
xnor UO_2584 (O_2584,N_24833,N_24545);
nand UO_2585 (O_2585,N_24756,N_24741);
or UO_2586 (O_2586,N_24933,N_24652);
and UO_2587 (O_2587,N_24750,N_24555);
nor UO_2588 (O_2588,N_24751,N_24894);
xnor UO_2589 (O_2589,N_24707,N_24822);
and UO_2590 (O_2590,N_24699,N_24885);
and UO_2591 (O_2591,N_24992,N_24852);
and UO_2592 (O_2592,N_24810,N_24627);
and UO_2593 (O_2593,N_24737,N_24812);
nor UO_2594 (O_2594,N_24726,N_24927);
xor UO_2595 (O_2595,N_24832,N_24872);
and UO_2596 (O_2596,N_24709,N_24631);
nor UO_2597 (O_2597,N_24655,N_24794);
or UO_2598 (O_2598,N_24853,N_24715);
nor UO_2599 (O_2599,N_24996,N_24567);
xnor UO_2600 (O_2600,N_24801,N_24820);
or UO_2601 (O_2601,N_24700,N_24857);
and UO_2602 (O_2602,N_24569,N_24963);
or UO_2603 (O_2603,N_24757,N_24715);
and UO_2604 (O_2604,N_24781,N_24923);
xor UO_2605 (O_2605,N_24927,N_24655);
nor UO_2606 (O_2606,N_24769,N_24655);
or UO_2607 (O_2607,N_24623,N_24670);
and UO_2608 (O_2608,N_24697,N_24578);
and UO_2609 (O_2609,N_24547,N_24505);
nor UO_2610 (O_2610,N_24553,N_24907);
or UO_2611 (O_2611,N_24626,N_24613);
nand UO_2612 (O_2612,N_24645,N_24859);
or UO_2613 (O_2613,N_24987,N_24694);
nor UO_2614 (O_2614,N_24813,N_24959);
or UO_2615 (O_2615,N_24822,N_24927);
nand UO_2616 (O_2616,N_24542,N_24674);
or UO_2617 (O_2617,N_24741,N_24569);
nand UO_2618 (O_2618,N_24954,N_24702);
nor UO_2619 (O_2619,N_24529,N_24548);
and UO_2620 (O_2620,N_24568,N_24682);
nand UO_2621 (O_2621,N_24667,N_24848);
xor UO_2622 (O_2622,N_24504,N_24512);
xor UO_2623 (O_2623,N_24526,N_24985);
nor UO_2624 (O_2624,N_24584,N_24606);
or UO_2625 (O_2625,N_24731,N_24942);
xor UO_2626 (O_2626,N_24811,N_24583);
xnor UO_2627 (O_2627,N_24921,N_24757);
nand UO_2628 (O_2628,N_24694,N_24616);
nand UO_2629 (O_2629,N_24611,N_24574);
or UO_2630 (O_2630,N_24702,N_24599);
nand UO_2631 (O_2631,N_24705,N_24653);
or UO_2632 (O_2632,N_24773,N_24799);
xor UO_2633 (O_2633,N_24953,N_24630);
and UO_2634 (O_2634,N_24889,N_24761);
nor UO_2635 (O_2635,N_24733,N_24666);
xor UO_2636 (O_2636,N_24703,N_24893);
or UO_2637 (O_2637,N_24690,N_24727);
nand UO_2638 (O_2638,N_24644,N_24509);
xor UO_2639 (O_2639,N_24628,N_24776);
nor UO_2640 (O_2640,N_24501,N_24651);
xnor UO_2641 (O_2641,N_24909,N_24704);
and UO_2642 (O_2642,N_24797,N_24545);
or UO_2643 (O_2643,N_24600,N_24815);
and UO_2644 (O_2644,N_24900,N_24944);
or UO_2645 (O_2645,N_24646,N_24891);
and UO_2646 (O_2646,N_24542,N_24971);
xor UO_2647 (O_2647,N_24766,N_24809);
nand UO_2648 (O_2648,N_24783,N_24637);
nand UO_2649 (O_2649,N_24629,N_24772);
or UO_2650 (O_2650,N_24754,N_24536);
xor UO_2651 (O_2651,N_24617,N_24820);
and UO_2652 (O_2652,N_24950,N_24857);
and UO_2653 (O_2653,N_24883,N_24724);
xor UO_2654 (O_2654,N_24556,N_24769);
xnor UO_2655 (O_2655,N_24629,N_24799);
nor UO_2656 (O_2656,N_24880,N_24707);
nand UO_2657 (O_2657,N_24635,N_24604);
nor UO_2658 (O_2658,N_24726,N_24834);
or UO_2659 (O_2659,N_24859,N_24519);
and UO_2660 (O_2660,N_24846,N_24531);
nand UO_2661 (O_2661,N_24713,N_24533);
or UO_2662 (O_2662,N_24997,N_24704);
xor UO_2663 (O_2663,N_24856,N_24554);
nor UO_2664 (O_2664,N_24536,N_24565);
nand UO_2665 (O_2665,N_24618,N_24953);
nand UO_2666 (O_2666,N_24610,N_24888);
and UO_2667 (O_2667,N_24708,N_24622);
nand UO_2668 (O_2668,N_24637,N_24529);
nor UO_2669 (O_2669,N_24506,N_24616);
nand UO_2670 (O_2670,N_24860,N_24665);
and UO_2671 (O_2671,N_24728,N_24644);
xor UO_2672 (O_2672,N_24771,N_24968);
xor UO_2673 (O_2673,N_24776,N_24960);
and UO_2674 (O_2674,N_24659,N_24872);
and UO_2675 (O_2675,N_24523,N_24795);
or UO_2676 (O_2676,N_24607,N_24608);
or UO_2677 (O_2677,N_24598,N_24502);
nor UO_2678 (O_2678,N_24588,N_24711);
nand UO_2679 (O_2679,N_24722,N_24707);
xnor UO_2680 (O_2680,N_24523,N_24684);
and UO_2681 (O_2681,N_24805,N_24856);
nand UO_2682 (O_2682,N_24628,N_24503);
xnor UO_2683 (O_2683,N_24885,N_24936);
or UO_2684 (O_2684,N_24561,N_24987);
nor UO_2685 (O_2685,N_24870,N_24638);
xor UO_2686 (O_2686,N_24522,N_24891);
nand UO_2687 (O_2687,N_24930,N_24655);
nor UO_2688 (O_2688,N_24524,N_24506);
and UO_2689 (O_2689,N_24923,N_24905);
xnor UO_2690 (O_2690,N_24768,N_24505);
nand UO_2691 (O_2691,N_24833,N_24556);
xor UO_2692 (O_2692,N_24637,N_24842);
or UO_2693 (O_2693,N_24953,N_24930);
or UO_2694 (O_2694,N_24540,N_24556);
and UO_2695 (O_2695,N_24593,N_24982);
nor UO_2696 (O_2696,N_24627,N_24919);
nand UO_2697 (O_2697,N_24568,N_24642);
or UO_2698 (O_2698,N_24840,N_24595);
nand UO_2699 (O_2699,N_24922,N_24987);
nor UO_2700 (O_2700,N_24898,N_24900);
or UO_2701 (O_2701,N_24543,N_24532);
or UO_2702 (O_2702,N_24544,N_24664);
or UO_2703 (O_2703,N_24715,N_24502);
nand UO_2704 (O_2704,N_24557,N_24902);
xor UO_2705 (O_2705,N_24719,N_24777);
or UO_2706 (O_2706,N_24512,N_24531);
nor UO_2707 (O_2707,N_24594,N_24501);
nand UO_2708 (O_2708,N_24774,N_24509);
and UO_2709 (O_2709,N_24538,N_24903);
xnor UO_2710 (O_2710,N_24970,N_24875);
xnor UO_2711 (O_2711,N_24511,N_24666);
xor UO_2712 (O_2712,N_24891,N_24594);
nand UO_2713 (O_2713,N_24753,N_24874);
or UO_2714 (O_2714,N_24629,N_24580);
or UO_2715 (O_2715,N_24850,N_24971);
nor UO_2716 (O_2716,N_24835,N_24951);
or UO_2717 (O_2717,N_24730,N_24677);
nand UO_2718 (O_2718,N_24898,N_24605);
nor UO_2719 (O_2719,N_24634,N_24699);
nand UO_2720 (O_2720,N_24529,N_24657);
nand UO_2721 (O_2721,N_24520,N_24631);
nand UO_2722 (O_2722,N_24807,N_24566);
nor UO_2723 (O_2723,N_24836,N_24507);
nor UO_2724 (O_2724,N_24942,N_24642);
nand UO_2725 (O_2725,N_24720,N_24878);
nor UO_2726 (O_2726,N_24909,N_24700);
nor UO_2727 (O_2727,N_24606,N_24697);
nor UO_2728 (O_2728,N_24792,N_24648);
and UO_2729 (O_2729,N_24621,N_24591);
nand UO_2730 (O_2730,N_24610,N_24924);
nand UO_2731 (O_2731,N_24668,N_24569);
xor UO_2732 (O_2732,N_24783,N_24559);
and UO_2733 (O_2733,N_24641,N_24957);
nand UO_2734 (O_2734,N_24662,N_24867);
xor UO_2735 (O_2735,N_24664,N_24557);
xor UO_2736 (O_2736,N_24710,N_24962);
nand UO_2737 (O_2737,N_24711,N_24926);
or UO_2738 (O_2738,N_24659,N_24739);
nor UO_2739 (O_2739,N_24933,N_24680);
nor UO_2740 (O_2740,N_24643,N_24681);
nor UO_2741 (O_2741,N_24679,N_24806);
xnor UO_2742 (O_2742,N_24760,N_24961);
nand UO_2743 (O_2743,N_24957,N_24726);
or UO_2744 (O_2744,N_24569,N_24803);
nand UO_2745 (O_2745,N_24794,N_24598);
and UO_2746 (O_2746,N_24629,N_24571);
nor UO_2747 (O_2747,N_24617,N_24989);
nor UO_2748 (O_2748,N_24830,N_24847);
xnor UO_2749 (O_2749,N_24758,N_24526);
or UO_2750 (O_2750,N_24862,N_24760);
xor UO_2751 (O_2751,N_24985,N_24798);
nand UO_2752 (O_2752,N_24694,N_24791);
nand UO_2753 (O_2753,N_24845,N_24758);
nand UO_2754 (O_2754,N_24717,N_24560);
and UO_2755 (O_2755,N_24666,N_24957);
nor UO_2756 (O_2756,N_24695,N_24999);
nor UO_2757 (O_2757,N_24898,N_24553);
xor UO_2758 (O_2758,N_24645,N_24919);
nand UO_2759 (O_2759,N_24527,N_24756);
nand UO_2760 (O_2760,N_24695,N_24881);
xor UO_2761 (O_2761,N_24843,N_24746);
nand UO_2762 (O_2762,N_24817,N_24625);
nor UO_2763 (O_2763,N_24920,N_24642);
xor UO_2764 (O_2764,N_24923,N_24581);
nor UO_2765 (O_2765,N_24527,N_24836);
xor UO_2766 (O_2766,N_24836,N_24501);
and UO_2767 (O_2767,N_24744,N_24750);
xnor UO_2768 (O_2768,N_24613,N_24844);
or UO_2769 (O_2769,N_24808,N_24549);
or UO_2770 (O_2770,N_24859,N_24839);
or UO_2771 (O_2771,N_24520,N_24925);
and UO_2772 (O_2772,N_24504,N_24818);
or UO_2773 (O_2773,N_24929,N_24930);
nor UO_2774 (O_2774,N_24637,N_24854);
and UO_2775 (O_2775,N_24688,N_24582);
nand UO_2776 (O_2776,N_24799,N_24707);
nor UO_2777 (O_2777,N_24588,N_24757);
nand UO_2778 (O_2778,N_24666,N_24664);
or UO_2779 (O_2779,N_24872,N_24962);
nor UO_2780 (O_2780,N_24513,N_24596);
or UO_2781 (O_2781,N_24984,N_24853);
nor UO_2782 (O_2782,N_24572,N_24531);
xor UO_2783 (O_2783,N_24654,N_24750);
xor UO_2784 (O_2784,N_24993,N_24663);
nand UO_2785 (O_2785,N_24539,N_24597);
nand UO_2786 (O_2786,N_24831,N_24959);
or UO_2787 (O_2787,N_24777,N_24630);
nand UO_2788 (O_2788,N_24506,N_24863);
xor UO_2789 (O_2789,N_24709,N_24857);
or UO_2790 (O_2790,N_24704,N_24824);
or UO_2791 (O_2791,N_24631,N_24536);
nand UO_2792 (O_2792,N_24503,N_24936);
nor UO_2793 (O_2793,N_24763,N_24858);
nand UO_2794 (O_2794,N_24590,N_24870);
nand UO_2795 (O_2795,N_24788,N_24670);
and UO_2796 (O_2796,N_24708,N_24647);
nand UO_2797 (O_2797,N_24952,N_24733);
nand UO_2798 (O_2798,N_24809,N_24507);
or UO_2799 (O_2799,N_24577,N_24804);
xnor UO_2800 (O_2800,N_24956,N_24906);
or UO_2801 (O_2801,N_24674,N_24712);
and UO_2802 (O_2802,N_24646,N_24692);
and UO_2803 (O_2803,N_24647,N_24590);
or UO_2804 (O_2804,N_24770,N_24992);
or UO_2805 (O_2805,N_24663,N_24755);
and UO_2806 (O_2806,N_24842,N_24588);
nand UO_2807 (O_2807,N_24547,N_24872);
or UO_2808 (O_2808,N_24738,N_24977);
or UO_2809 (O_2809,N_24993,N_24789);
or UO_2810 (O_2810,N_24740,N_24640);
nand UO_2811 (O_2811,N_24765,N_24954);
nand UO_2812 (O_2812,N_24554,N_24578);
nor UO_2813 (O_2813,N_24922,N_24536);
nor UO_2814 (O_2814,N_24679,N_24980);
nor UO_2815 (O_2815,N_24552,N_24838);
nand UO_2816 (O_2816,N_24858,N_24711);
xnor UO_2817 (O_2817,N_24915,N_24638);
nor UO_2818 (O_2818,N_24645,N_24517);
xor UO_2819 (O_2819,N_24535,N_24763);
and UO_2820 (O_2820,N_24846,N_24509);
nand UO_2821 (O_2821,N_24781,N_24870);
nand UO_2822 (O_2822,N_24892,N_24843);
or UO_2823 (O_2823,N_24740,N_24666);
nand UO_2824 (O_2824,N_24672,N_24919);
nand UO_2825 (O_2825,N_24729,N_24708);
xor UO_2826 (O_2826,N_24815,N_24926);
nor UO_2827 (O_2827,N_24826,N_24695);
nand UO_2828 (O_2828,N_24797,N_24505);
nor UO_2829 (O_2829,N_24731,N_24799);
and UO_2830 (O_2830,N_24775,N_24927);
xnor UO_2831 (O_2831,N_24854,N_24718);
nor UO_2832 (O_2832,N_24976,N_24849);
and UO_2833 (O_2833,N_24836,N_24643);
nor UO_2834 (O_2834,N_24727,N_24782);
nand UO_2835 (O_2835,N_24681,N_24574);
and UO_2836 (O_2836,N_24932,N_24621);
and UO_2837 (O_2837,N_24610,N_24866);
nor UO_2838 (O_2838,N_24941,N_24838);
and UO_2839 (O_2839,N_24916,N_24560);
nor UO_2840 (O_2840,N_24534,N_24850);
or UO_2841 (O_2841,N_24568,N_24825);
xnor UO_2842 (O_2842,N_24891,N_24973);
and UO_2843 (O_2843,N_24507,N_24843);
and UO_2844 (O_2844,N_24894,N_24974);
and UO_2845 (O_2845,N_24930,N_24759);
xnor UO_2846 (O_2846,N_24609,N_24953);
or UO_2847 (O_2847,N_24708,N_24717);
or UO_2848 (O_2848,N_24526,N_24661);
nor UO_2849 (O_2849,N_24826,N_24831);
nor UO_2850 (O_2850,N_24832,N_24822);
nor UO_2851 (O_2851,N_24854,N_24583);
and UO_2852 (O_2852,N_24595,N_24566);
nand UO_2853 (O_2853,N_24601,N_24969);
and UO_2854 (O_2854,N_24800,N_24885);
and UO_2855 (O_2855,N_24849,N_24536);
and UO_2856 (O_2856,N_24831,N_24774);
nand UO_2857 (O_2857,N_24807,N_24548);
or UO_2858 (O_2858,N_24509,N_24744);
xor UO_2859 (O_2859,N_24594,N_24969);
and UO_2860 (O_2860,N_24701,N_24577);
nand UO_2861 (O_2861,N_24505,N_24609);
and UO_2862 (O_2862,N_24863,N_24927);
xnor UO_2863 (O_2863,N_24996,N_24834);
xor UO_2864 (O_2864,N_24528,N_24910);
nor UO_2865 (O_2865,N_24583,N_24963);
and UO_2866 (O_2866,N_24596,N_24781);
nand UO_2867 (O_2867,N_24767,N_24884);
nor UO_2868 (O_2868,N_24886,N_24798);
nand UO_2869 (O_2869,N_24814,N_24933);
nor UO_2870 (O_2870,N_24872,N_24794);
and UO_2871 (O_2871,N_24758,N_24733);
xor UO_2872 (O_2872,N_24883,N_24612);
nor UO_2873 (O_2873,N_24596,N_24798);
and UO_2874 (O_2874,N_24818,N_24733);
or UO_2875 (O_2875,N_24668,N_24954);
nand UO_2876 (O_2876,N_24722,N_24779);
and UO_2877 (O_2877,N_24789,N_24936);
nor UO_2878 (O_2878,N_24731,N_24578);
xor UO_2879 (O_2879,N_24685,N_24734);
nor UO_2880 (O_2880,N_24846,N_24646);
or UO_2881 (O_2881,N_24843,N_24938);
nor UO_2882 (O_2882,N_24740,N_24679);
nand UO_2883 (O_2883,N_24509,N_24957);
nand UO_2884 (O_2884,N_24558,N_24909);
nand UO_2885 (O_2885,N_24516,N_24535);
nor UO_2886 (O_2886,N_24783,N_24898);
or UO_2887 (O_2887,N_24520,N_24885);
nor UO_2888 (O_2888,N_24562,N_24525);
xor UO_2889 (O_2889,N_24781,N_24554);
nor UO_2890 (O_2890,N_24572,N_24507);
or UO_2891 (O_2891,N_24859,N_24540);
nand UO_2892 (O_2892,N_24833,N_24728);
nand UO_2893 (O_2893,N_24690,N_24606);
nand UO_2894 (O_2894,N_24758,N_24898);
or UO_2895 (O_2895,N_24757,N_24982);
or UO_2896 (O_2896,N_24611,N_24764);
nor UO_2897 (O_2897,N_24830,N_24848);
and UO_2898 (O_2898,N_24678,N_24592);
xor UO_2899 (O_2899,N_24916,N_24518);
and UO_2900 (O_2900,N_24937,N_24724);
and UO_2901 (O_2901,N_24679,N_24972);
xnor UO_2902 (O_2902,N_24772,N_24854);
and UO_2903 (O_2903,N_24886,N_24570);
nand UO_2904 (O_2904,N_24510,N_24671);
nor UO_2905 (O_2905,N_24863,N_24690);
xnor UO_2906 (O_2906,N_24764,N_24722);
nand UO_2907 (O_2907,N_24959,N_24867);
or UO_2908 (O_2908,N_24703,N_24988);
xor UO_2909 (O_2909,N_24832,N_24759);
or UO_2910 (O_2910,N_24629,N_24591);
xnor UO_2911 (O_2911,N_24625,N_24834);
nor UO_2912 (O_2912,N_24869,N_24724);
xor UO_2913 (O_2913,N_24716,N_24843);
nor UO_2914 (O_2914,N_24934,N_24962);
xnor UO_2915 (O_2915,N_24704,N_24638);
xnor UO_2916 (O_2916,N_24654,N_24956);
and UO_2917 (O_2917,N_24787,N_24647);
nor UO_2918 (O_2918,N_24992,N_24633);
or UO_2919 (O_2919,N_24876,N_24805);
nor UO_2920 (O_2920,N_24801,N_24821);
nor UO_2921 (O_2921,N_24756,N_24751);
nand UO_2922 (O_2922,N_24544,N_24761);
xnor UO_2923 (O_2923,N_24675,N_24565);
nand UO_2924 (O_2924,N_24867,N_24539);
xnor UO_2925 (O_2925,N_24662,N_24793);
and UO_2926 (O_2926,N_24527,N_24917);
nor UO_2927 (O_2927,N_24590,N_24969);
or UO_2928 (O_2928,N_24834,N_24957);
nand UO_2929 (O_2929,N_24757,N_24841);
nor UO_2930 (O_2930,N_24671,N_24798);
nor UO_2931 (O_2931,N_24779,N_24884);
xor UO_2932 (O_2932,N_24796,N_24920);
nor UO_2933 (O_2933,N_24842,N_24530);
nor UO_2934 (O_2934,N_24794,N_24994);
nand UO_2935 (O_2935,N_24648,N_24877);
and UO_2936 (O_2936,N_24982,N_24639);
nand UO_2937 (O_2937,N_24613,N_24792);
xnor UO_2938 (O_2938,N_24922,N_24539);
and UO_2939 (O_2939,N_24922,N_24721);
xor UO_2940 (O_2940,N_24997,N_24821);
or UO_2941 (O_2941,N_24513,N_24727);
nand UO_2942 (O_2942,N_24829,N_24789);
or UO_2943 (O_2943,N_24897,N_24905);
and UO_2944 (O_2944,N_24933,N_24969);
or UO_2945 (O_2945,N_24553,N_24995);
or UO_2946 (O_2946,N_24840,N_24798);
nand UO_2947 (O_2947,N_24955,N_24867);
xnor UO_2948 (O_2948,N_24816,N_24894);
or UO_2949 (O_2949,N_24748,N_24635);
nor UO_2950 (O_2950,N_24730,N_24957);
or UO_2951 (O_2951,N_24865,N_24720);
nor UO_2952 (O_2952,N_24551,N_24898);
nand UO_2953 (O_2953,N_24656,N_24746);
nand UO_2954 (O_2954,N_24742,N_24512);
and UO_2955 (O_2955,N_24971,N_24968);
xnor UO_2956 (O_2956,N_24911,N_24786);
nand UO_2957 (O_2957,N_24526,N_24544);
or UO_2958 (O_2958,N_24558,N_24741);
nor UO_2959 (O_2959,N_24575,N_24908);
nor UO_2960 (O_2960,N_24703,N_24542);
or UO_2961 (O_2961,N_24671,N_24703);
and UO_2962 (O_2962,N_24820,N_24525);
or UO_2963 (O_2963,N_24913,N_24781);
and UO_2964 (O_2964,N_24632,N_24857);
or UO_2965 (O_2965,N_24919,N_24556);
and UO_2966 (O_2966,N_24564,N_24790);
or UO_2967 (O_2967,N_24877,N_24999);
nand UO_2968 (O_2968,N_24737,N_24605);
nor UO_2969 (O_2969,N_24984,N_24704);
and UO_2970 (O_2970,N_24974,N_24582);
or UO_2971 (O_2971,N_24717,N_24645);
nor UO_2972 (O_2972,N_24671,N_24532);
nor UO_2973 (O_2973,N_24614,N_24825);
or UO_2974 (O_2974,N_24585,N_24812);
nand UO_2975 (O_2975,N_24637,N_24523);
and UO_2976 (O_2976,N_24664,N_24788);
xor UO_2977 (O_2977,N_24755,N_24960);
xnor UO_2978 (O_2978,N_24943,N_24521);
or UO_2979 (O_2979,N_24760,N_24917);
nor UO_2980 (O_2980,N_24667,N_24642);
and UO_2981 (O_2981,N_24611,N_24795);
nor UO_2982 (O_2982,N_24805,N_24819);
nand UO_2983 (O_2983,N_24908,N_24940);
nand UO_2984 (O_2984,N_24636,N_24539);
nand UO_2985 (O_2985,N_24649,N_24814);
and UO_2986 (O_2986,N_24617,N_24876);
xor UO_2987 (O_2987,N_24962,N_24936);
or UO_2988 (O_2988,N_24690,N_24926);
nor UO_2989 (O_2989,N_24508,N_24565);
xor UO_2990 (O_2990,N_24763,N_24717);
nand UO_2991 (O_2991,N_24587,N_24708);
xor UO_2992 (O_2992,N_24500,N_24919);
xnor UO_2993 (O_2993,N_24521,N_24939);
nand UO_2994 (O_2994,N_24575,N_24749);
and UO_2995 (O_2995,N_24620,N_24745);
and UO_2996 (O_2996,N_24873,N_24582);
nor UO_2997 (O_2997,N_24517,N_24576);
nand UO_2998 (O_2998,N_24742,N_24833);
xnor UO_2999 (O_2999,N_24706,N_24965);
endmodule