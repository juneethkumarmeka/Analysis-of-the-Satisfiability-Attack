module basic_3000_30000_3500_100_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1059,In_1026);
nand U1 (N_1,In_644,In_2445);
xor U2 (N_2,In_2267,In_2051);
and U3 (N_3,In_2028,In_1961);
nand U4 (N_4,In_2969,In_2586);
nor U5 (N_5,In_123,In_1948);
nand U6 (N_6,In_938,In_2964);
nor U7 (N_7,In_1137,In_2661);
nand U8 (N_8,In_1247,In_422);
or U9 (N_9,In_1772,In_1104);
or U10 (N_10,In_794,In_2485);
nor U11 (N_11,In_710,In_2551);
nor U12 (N_12,In_197,In_858);
and U13 (N_13,In_2546,In_444);
or U14 (N_14,In_1211,In_2321);
and U15 (N_15,In_745,In_1887);
and U16 (N_16,In_1487,In_364);
or U17 (N_17,In_902,In_1447);
or U18 (N_18,In_2867,In_1387);
or U19 (N_19,In_985,In_2789);
xnor U20 (N_20,In_1505,In_564);
or U21 (N_21,In_1644,In_1987);
and U22 (N_22,In_2709,In_115);
or U23 (N_23,In_2058,In_1375);
and U24 (N_24,In_1632,In_660);
nor U25 (N_25,In_2752,In_2802);
and U26 (N_26,In_2647,In_1965);
nor U27 (N_27,In_1468,In_1103);
xnor U28 (N_28,In_1662,In_1429);
xnor U29 (N_29,In_1646,In_1759);
nor U30 (N_30,In_128,In_683);
nand U31 (N_31,In_299,In_2944);
and U32 (N_32,In_1833,In_697);
nand U33 (N_33,In_2530,In_2140);
xor U34 (N_34,In_201,In_318);
nand U35 (N_35,In_1883,In_2615);
xor U36 (N_36,In_484,In_1284);
and U37 (N_37,In_2383,In_1265);
and U38 (N_38,In_735,In_1074);
nor U39 (N_39,In_1194,In_1323);
nor U40 (N_40,In_350,In_28);
or U41 (N_41,In_175,In_1183);
nand U42 (N_42,In_1845,In_1155);
nor U43 (N_43,In_2759,In_44);
and U44 (N_44,In_1193,In_1302);
or U45 (N_45,In_2504,In_2295);
nor U46 (N_46,In_2856,In_709);
nand U47 (N_47,In_2508,In_502);
or U48 (N_48,In_1495,In_2772);
xor U49 (N_49,In_675,In_692);
nand U50 (N_50,In_2141,In_2325);
nand U51 (N_51,In_574,In_2132);
nand U52 (N_52,In_2370,In_1304);
nand U53 (N_53,In_483,In_248);
and U54 (N_54,In_2701,In_1233);
and U55 (N_55,In_1364,In_1145);
nand U56 (N_56,In_2510,In_698);
or U57 (N_57,In_2719,In_2932);
nor U58 (N_58,In_593,In_649);
xor U59 (N_59,In_2452,In_2684);
xnor U60 (N_60,In_650,In_152);
nor U61 (N_61,In_1869,In_839);
or U62 (N_62,In_1854,In_1692);
or U63 (N_63,In_525,In_1085);
and U64 (N_64,In_846,In_2844);
xor U65 (N_65,In_630,In_1782);
xor U66 (N_66,In_277,In_1484);
or U67 (N_67,In_1035,In_1492);
nand U68 (N_68,In_2150,In_2);
nand U69 (N_69,In_2162,In_951);
nor U70 (N_70,In_2158,In_897);
xnor U71 (N_71,In_2562,In_92);
and U72 (N_72,In_757,In_2946);
and U73 (N_73,In_640,In_1036);
xor U74 (N_74,In_2721,In_2027);
xnor U75 (N_75,In_958,In_2939);
or U76 (N_76,In_1688,In_273);
and U77 (N_77,In_1067,In_2926);
or U78 (N_78,In_2798,In_2423);
nor U79 (N_79,In_2715,In_2520);
and U80 (N_80,In_2481,In_312);
nand U81 (N_81,In_2446,In_2251);
nor U82 (N_82,In_2283,In_1723);
or U83 (N_83,In_1693,In_1175);
or U84 (N_84,In_1628,In_1123);
and U85 (N_85,In_1722,In_1620);
nand U86 (N_86,In_2912,In_1844);
nand U87 (N_87,In_1824,In_1432);
and U88 (N_88,In_1684,In_1301);
nand U89 (N_89,In_2476,In_311);
nand U90 (N_90,In_1511,In_2369);
nand U91 (N_91,In_789,In_2529);
nor U92 (N_92,In_740,In_1865);
or U93 (N_93,In_2927,In_2978);
or U94 (N_94,In_852,In_1139);
and U95 (N_95,In_1762,In_1376);
nor U96 (N_96,In_2489,In_2455);
xnor U97 (N_97,In_379,In_82);
nor U98 (N_98,In_721,In_1368);
or U99 (N_99,In_1130,In_96);
or U100 (N_100,In_2870,In_2623);
nand U101 (N_101,In_2247,In_118);
and U102 (N_102,In_2070,In_2148);
and U103 (N_103,In_2514,In_1070);
or U104 (N_104,In_158,In_2724);
nor U105 (N_105,In_1452,In_2749);
nor U106 (N_106,In_2359,In_278);
nand U107 (N_107,In_1581,In_1348);
nand U108 (N_108,In_2386,In_1899);
xnor U109 (N_109,In_101,In_1399);
nor U110 (N_110,In_1731,In_548);
nand U111 (N_111,In_1148,In_963);
or U112 (N_112,In_908,In_2608);
xor U113 (N_113,In_1951,In_2449);
xnor U114 (N_114,In_1486,In_2518);
or U115 (N_115,In_2794,In_1808);
nand U116 (N_116,In_1326,In_287);
or U117 (N_117,In_2406,In_861);
or U118 (N_118,In_2891,In_2061);
nand U119 (N_119,In_2305,In_134);
xnor U120 (N_120,In_217,In_1702);
nand U121 (N_121,In_409,In_1790);
nor U122 (N_122,In_2569,In_790);
and U123 (N_123,In_406,In_2670);
xnor U124 (N_124,In_301,In_1397);
and U125 (N_125,In_2253,In_1989);
nor U126 (N_126,In_2490,In_2974);
xor U127 (N_127,In_2293,In_1793);
or U128 (N_128,In_1150,In_1340);
xor U129 (N_129,In_2484,In_1236);
and U130 (N_130,In_2071,In_1794);
nor U131 (N_131,In_38,In_2923);
xor U132 (N_132,In_718,In_1332);
or U133 (N_133,In_2373,In_2971);
xor U134 (N_134,In_5,In_270);
nor U135 (N_135,In_1330,In_2074);
or U136 (N_136,In_1999,In_339);
or U137 (N_137,In_2091,In_727);
nor U138 (N_138,In_2788,In_1400);
xnor U139 (N_139,In_453,In_1312);
or U140 (N_140,In_2634,In_2713);
or U141 (N_141,In_1874,In_1079);
nor U142 (N_142,In_1125,In_1599);
xnor U143 (N_143,In_2558,In_202);
nor U144 (N_144,In_1280,In_605);
or U145 (N_145,In_2742,In_1699);
and U146 (N_146,In_666,In_2756);
nand U147 (N_147,In_1333,In_360);
or U148 (N_148,In_863,In_944);
nand U149 (N_149,In_988,In_2109);
nand U150 (N_150,In_1966,In_2873);
nor U151 (N_151,In_2164,In_2997);
and U152 (N_152,In_1308,In_2911);
nand U153 (N_153,In_2747,In_754);
xor U154 (N_154,In_1479,In_2255);
and U155 (N_155,In_983,In_1653);
nor U156 (N_156,In_346,In_1499);
xnor U157 (N_157,In_1296,In_836);
nand U158 (N_158,In_89,In_616);
nor U159 (N_159,In_2730,In_2838);
xor U160 (N_160,In_1954,In_1357);
xor U161 (N_161,In_2221,In_2108);
or U162 (N_162,In_1923,In_271);
nor U163 (N_163,In_1893,In_1658);
and U164 (N_164,In_2516,In_2081);
xnor U165 (N_165,In_116,In_2983);
nor U166 (N_166,In_1473,In_2231);
xor U167 (N_167,In_1876,In_1890);
xor U168 (N_168,In_1045,In_2881);
and U169 (N_169,In_1564,In_763);
or U170 (N_170,In_1986,In_1570);
xnor U171 (N_171,In_143,In_1713);
xor U172 (N_172,In_357,In_1889);
nor U173 (N_173,In_1621,In_1920);
and U174 (N_174,In_2956,In_1633);
and U175 (N_175,In_2063,In_2901);
and U176 (N_176,In_1536,In_2531);
or U177 (N_177,In_1114,In_141);
xor U178 (N_178,In_1389,In_747);
or U179 (N_179,In_1988,In_374);
and U180 (N_180,In_2850,In_682);
or U181 (N_181,In_600,In_471);
xnor U182 (N_182,In_2821,In_40);
nand U183 (N_183,In_1540,In_2130);
nand U184 (N_184,In_1521,In_2338);
nor U185 (N_185,In_451,In_594);
and U186 (N_186,In_1083,In_377);
or U187 (N_187,In_1975,In_722);
nor U188 (N_188,In_359,In_2826);
or U189 (N_189,In_1803,In_730);
and U190 (N_190,In_2493,In_2152);
or U191 (N_191,In_1984,In_1320);
xor U192 (N_192,In_1545,In_1047);
and U193 (N_193,In_284,In_263);
xnor U194 (N_194,In_2843,In_2994);
xnor U195 (N_195,In_2839,In_2077);
xnor U196 (N_196,In_2420,In_1027);
and U197 (N_197,In_1503,In_2167);
or U198 (N_198,In_170,In_1622);
xnor U199 (N_199,In_333,In_1697);
nor U200 (N_200,In_1502,In_2575);
nand U201 (N_201,In_962,In_1610);
xor U202 (N_202,In_862,In_2085);
and U203 (N_203,In_1601,In_769);
nor U204 (N_204,In_1289,In_191);
and U205 (N_205,In_1063,In_883);
xnor U206 (N_206,In_2212,In_2194);
and U207 (N_207,In_407,In_824);
or U208 (N_208,In_955,In_2111);
xor U209 (N_209,In_876,In_2793);
and U210 (N_210,In_2315,In_1940);
nor U211 (N_211,In_35,In_651);
and U212 (N_212,In_1664,In_1917);
or U213 (N_213,In_419,In_245);
nor U214 (N_214,In_2755,In_2536);
and U215 (N_215,In_1480,In_635);
and U216 (N_216,In_937,In_2435);
or U217 (N_217,In_652,In_386);
xor U218 (N_218,In_1600,In_620);
nor U219 (N_219,In_1491,In_654);
nor U220 (N_220,In_545,In_336);
or U221 (N_221,In_2306,In_183);
and U222 (N_222,In_1677,In_2662);
nand U223 (N_223,In_1356,In_2215);
and U224 (N_224,In_1629,In_719);
and U225 (N_225,In_2522,In_822);
and U226 (N_226,In_2534,In_1154);
and U227 (N_227,In_1956,In_93);
and U228 (N_228,In_1317,In_1182);
and U229 (N_229,In_739,In_1441);
nor U230 (N_230,In_2754,In_375);
xnor U231 (N_231,In_353,In_2774);
and U232 (N_232,In_172,In_1345);
and U233 (N_233,In_2426,In_2953);
or U234 (N_234,In_2013,In_2419);
or U235 (N_235,In_2779,In_2790);
xnor U236 (N_236,In_954,In_592);
nand U237 (N_237,In_1589,In_1748);
and U238 (N_238,In_1926,In_1823);
nand U239 (N_239,In_493,In_2578);
nand U240 (N_240,In_680,In_1466);
and U241 (N_241,In_1025,In_16);
nor U242 (N_242,In_410,In_971);
and U243 (N_243,In_2210,In_1678);
or U244 (N_244,In_1347,In_1980);
nor U245 (N_245,In_2133,In_1741);
xor U246 (N_246,In_2765,In_1209);
xnor U247 (N_247,In_1555,In_1377);
and U248 (N_248,In_693,In_1766);
nand U249 (N_249,In_1373,In_1995);
nand U250 (N_250,In_1592,In_2598);
xor U251 (N_251,In_2422,In_2332);
xor U252 (N_252,In_1017,In_588);
nor U253 (N_253,In_2631,In_750);
nor U254 (N_254,In_687,In_546);
nand U255 (N_255,In_1634,In_2766);
nand U256 (N_256,In_1138,In_286);
nor U257 (N_257,In_927,In_2640);
nand U258 (N_258,In_2521,In_1005);
nand U259 (N_259,In_1162,In_845);
or U260 (N_260,In_925,In_214);
nand U261 (N_261,In_61,In_2003);
nor U262 (N_262,In_1242,In_2000);
nand U263 (N_263,In_1590,In_404);
xor U264 (N_264,In_1635,In_1949);
nand U265 (N_265,In_2596,In_1094);
or U266 (N_266,In_665,In_372);
nor U267 (N_267,In_1173,In_1616);
nand U268 (N_268,In_2907,In_80);
and U269 (N_269,In_521,In_1215);
nand U270 (N_270,In_1469,In_1444);
nand U271 (N_271,In_1735,In_992);
or U272 (N_272,In_2031,In_1573);
or U273 (N_273,In_2635,In_2418);
xnor U274 (N_274,In_633,In_2101);
nor U275 (N_275,In_1857,In_2552);
nor U276 (N_276,In_2023,In_999);
nand U277 (N_277,In_1060,In_434);
xnor U278 (N_278,In_511,In_1812);
xor U279 (N_279,In_124,In_1538);
xor U280 (N_280,In_2363,In_1720);
nor U281 (N_281,In_322,In_2758);
or U282 (N_282,In_2541,In_2094);
xor U283 (N_283,In_1195,In_1128);
nand U284 (N_284,In_1146,In_1755);
nor U285 (N_285,In_2260,In_1813);
and U286 (N_286,In_877,In_52);
xnor U287 (N_287,In_950,In_1371);
xor U288 (N_288,In_2625,In_2716);
nor U289 (N_289,In_2746,In_309);
nor U290 (N_290,In_343,In_2833);
or U291 (N_291,In_1134,In_1033);
nor U292 (N_292,In_2436,In_1321);
nand U293 (N_293,In_1497,In_2135);
nor U294 (N_294,In_1732,In_889);
nand U295 (N_295,In_1843,In_2344);
nor U296 (N_296,In_974,In_597);
or U297 (N_297,In_2110,In_1351);
or U298 (N_298,In_2218,In_1181);
nand U299 (N_299,In_2544,In_1878);
xor U300 (N_300,In_1597,In_2859);
xor U301 (N_301,In_1197,In_1614);
or U302 (N_302,In_2041,In_2375);
and U303 (N_303,N_265,In_753);
or U304 (N_304,In_85,In_536);
xor U305 (N_305,In_1271,In_94);
xnor U306 (N_306,In_986,In_543);
and U307 (N_307,In_473,In_972);
or U308 (N_308,In_32,In_1513);
nor U309 (N_309,In_569,In_2156);
nor U310 (N_310,In_1553,In_2066);
or U311 (N_311,In_1850,In_2112);
or U312 (N_312,In_2036,In_2813);
nand U313 (N_313,In_2734,In_1086);
xor U314 (N_314,In_1073,In_1485);
nor U315 (N_315,In_667,In_1645);
xor U316 (N_316,In_788,In_1219);
nor U317 (N_317,In_976,In_420);
or U318 (N_318,In_2176,In_1303);
and U319 (N_319,In_373,In_157);
and U320 (N_320,In_2024,In_1336);
xnor U321 (N_321,In_1087,In_1695);
and U322 (N_322,In_1042,In_2834);
xnor U323 (N_323,In_1216,In_1230);
xnor U324 (N_324,N_224,In_2264);
xor U325 (N_325,In_800,In_1038);
or U326 (N_326,In_480,N_294);
and U327 (N_327,In_923,In_837);
nand U328 (N_328,In_1,In_2035);
xnor U329 (N_329,In_1488,In_2918);
nor U330 (N_330,In_2378,In_2361);
and U331 (N_331,In_487,In_2694);
and U332 (N_332,In_2962,In_261);
or U333 (N_333,In_1529,In_1274);
and U334 (N_334,In_1167,In_1249);
xnor U335 (N_335,N_100,In_2052);
nand U336 (N_336,In_209,In_1819);
and U337 (N_337,In_1921,In_2669);
xor U338 (N_338,In_812,In_2224);
and U339 (N_339,In_155,In_2188);
nor U340 (N_340,In_538,In_1817);
xnor U341 (N_341,In_964,In_1548);
and U342 (N_342,In_1652,In_1269);
or U343 (N_343,In_577,In_1825);
xor U344 (N_344,In_669,In_84);
nand U345 (N_345,In_1852,N_218);
xnor U346 (N_346,In_10,In_2966);
or U347 (N_347,In_423,In_475);
xor U348 (N_348,In_1178,N_213);
xnor U349 (N_349,In_668,In_1171);
and U350 (N_350,N_138,In_413);
or U351 (N_351,N_76,N_28);
and U352 (N_352,In_1919,In_1868);
or U353 (N_353,In_1111,In_922);
xnor U354 (N_354,In_2161,In_2915);
nand U355 (N_355,In_1907,N_246);
nand U356 (N_356,In_2401,In_1282);
or U357 (N_357,In_1405,In_2480);
xnor U358 (N_358,In_1751,In_1906);
nand U359 (N_359,In_868,In_1580);
nand U360 (N_360,In_507,In_2745);
nor U361 (N_361,In_2589,In_2233);
xor U362 (N_362,In_441,In_2393);
xor U363 (N_363,In_1252,In_2987);
or U364 (N_364,In_2689,In_1524);
nor U365 (N_365,In_1300,In_1065);
or U366 (N_366,In_399,N_119);
nor U367 (N_367,In_833,In_2654);
or U368 (N_368,In_2054,In_2909);
or U369 (N_369,In_2460,In_168);
nor U370 (N_370,In_1403,N_98);
nor U371 (N_371,In_2645,In_637);
nand U372 (N_372,In_2883,In_989);
nand U373 (N_373,N_171,In_859);
nand U374 (N_374,In_1796,In_2650);
or U375 (N_375,In_899,In_997);
nor U376 (N_376,N_105,In_458);
and U377 (N_377,In_791,N_285);
or U378 (N_378,In_1957,In_2441);
nor U379 (N_379,In_2137,In_2098);
xor U380 (N_380,N_131,In_356);
nand U381 (N_381,In_57,In_1700);
and U382 (N_382,In_1354,In_1932);
nand U383 (N_383,In_2938,In_390);
nor U384 (N_384,In_695,N_149);
nand U385 (N_385,In_1864,In_2415);
nand U386 (N_386,In_793,In_1659);
nand U387 (N_387,N_217,In_2830);
nand U388 (N_388,In_1971,In_884);
or U389 (N_389,In_2026,In_1390);
xnor U390 (N_390,In_746,In_2319);
nor U391 (N_391,In_1305,N_216);
or U392 (N_392,In_2718,In_1562);
and U393 (N_393,In_498,In_1650);
or U394 (N_394,In_2169,In_756);
xnor U395 (N_395,In_940,In_811);
nand U396 (N_396,In_2588,In_365);
nand U397 (N_397,In_932,N_253);
and U398 (N_398,In_1341,In_2679);
or U399 (N_399,In_2620,In_2065);
and U400 (N_400,In_803,In_1711);
nand U401 (N_401,In_2506,In_392);
and U402 (N_402,In_557,In_266);
xor U403 (N_403,In_1947,In_1343);
or U404 (N_404,In_2868,In_1775);
and U405 (N_405,N_200,In_1196);
nor U406 (N_406,In_25,In_2576);
xor U407 (N_407,In_1836,N_175);
or U408 (N_408,In_907,In_1566);
nor U409 (N_409,In_2958,In_2903);
nand U410 (N_410,In_795,In_1584);
or U411 (N_411,In_1232,In_771);
nand U412 (N_412,In_1572,In_2428);
nor U413 (N_413,In_1648,In_260);
nor U414 (N_414,In_2560,In_1651);
xor U415 (N_415,In_2651,In_2889);
nand U416 (N_416,In_221,N_234);
or U417 (N_417,In_1152,In_247);
nand U418 (N_418,In_2667,In_1034);
nand U419 (N_419,In_780,In_2257);
or U420 (N_420,In_1806,N_29);
nand U421 (N_421,In_924,In_296);
nor U422 (N_422,In_1783,In_784);
or U423 (N_423,In_2600,In_2686);
nor U424 (N_424,In_2822,In_2092);
xnor U425 (N_425,In_2784,In_2427);
nor U426 (N_426,In_1728,N_183);
xor U427 (N_427,In_1832,In_2049);
and U428 (N_428,In_1792,In_1554);
or U429 (N_429,In_53,In_1929);
nand U430 (N_430,In_2463,In_2124);
nor U431 (N_431,In_2871,In_1007);
nor U432 (N_432,N_97,In_68);
nor U433 (N_433,In_2301,In_2314);
nand U434 (N_434,N_273,In_145);
nand U435 (N_435,In_1810,In_672);
xnor U436 (N_436,In_886,In_1112);
nor U437 (N_437,In_2440,In_547);
nor U438 (N_438,In_69,In_2878);
nor U439 (N_439,In_1334,In_184);
or U440 (N_440,In_1799,In_856);
nor U441 (N_441,In_2593,In_1604);
nand U442 (N_442,N_259,N_299);
nand U443 (N_443,In_809,In_2329);
nand U444 (N_444,N_147,In_1105);
and U445 (N_445,In_1443,In_655);
or U446 (N_446,In_1841,In_1478);
and U447 (N_447,In_1258,In_153);
nand U448 (N_448,In_2355,In_2285);
nand U449 (N_449,In_2835,In_349);
xor U450 (N_450,In_2913,In_2614);
xor U451 (N_451,N_108,In_1672);
and U452 (N_452,In_211,In_537);
nand U453 (N_453,In_323,In_321);
and U454 (N_454,In_1754,In_2324);
xor U455 (N_455,In_1424,In_2892);
xor U456 (N_456,In_1089,In_1270);
xor U457 (N_457,In_1264,In_2259);
or U458 (N_458,In_1743,In_2185);
and U459 (N_459,In_1024,In_2331);
and U460 (N_460,In_2992,In_2030);
or U461 (N_461,In_1546,In_1243);
xnor U462 (N_462,In_2131,In_1602);
and U463 (N_463,In_1950,In_738);
xor U464 (N_464,In_1307,In_2665);
or U465 (N_465,In_892,In_2043);
or U466 (N_466,In_1385,In_563);
xnor U467 (N_467,N_257,In_1346);
nand U468 (N_468,In_1687,In_775);
nor U469 (N_469,In_2919,In_2165);
xor U470 (N_470,In_1829,In_1626);
nor U471 (N_471,In_1338,In_2350);
xor U472 (N_472,In_393,In_1605);
xnor U473 (N_473,In_1180,In_1201);
and U474 (N_474,In_977,N_186);
nand U475 (N_475,In_41,In_1942);
nand U476 (N_476,In_2706,In_2323);
nor U477 (N_477,In_1462,In_2478);
and U478 (N_478,In_2523,In_2906);
and U479 (N_479,In_2115,In_678);
and U480 (N_480,In_131,In_1442);
xor U481 (N_481,In_580,In_1260);
and U482 (N_482,In_2948,In_361);
xor U483 (N_483,In_2767,In_2982);
or U484 (N_484,In_2975,In_384);
xor U485 (N_485,In_1608,N_47);
or U486 (N_486,In_1625,In_2379);
and U487 (N_487,In_969,N_248);
nor U488 (N_488,In_246,In_2543);
nor U489 (N_489,In_768,In_2567);
nand U490 (N_490,N_52,N_40);
and U491 (N_491,In_2688,In_774);
nor U492 (N_492,In_2290,In_2687);
nor U493 (N_493,In_820,In_2310);
nand U494 (N_494,In_711,In_1176);
or U495 (N_495,In_147,In_2413);
or U496 (N_496,In_2016,In_1023);
or U497 (N_497,In_2488,In_2151);
and U498 (N_498,In_2246,In_623);
xnor U499 (N_499,In_565,In_389);
and U500 (N_500,In_2082,In_734);
and U501 (N_501,In_250,In_2226);
nor U502 (N_502,In_2696,In_195);
xor U503 (N_503,In_1943,In_2429);
xor U504 (N_504,In_759,In_26);
or U505 (N_505,In_1217,In_2387);
nor U506 (N_506,In_1335,In_2568);
xnor U507 (N_507,In_1858,In_48);
or U508 (N_508,In_2791,In_1031);
or U509 (N_509,N_222,In_766);
and U510 (N_510,In_1863,In_1455);
xor U511 (N_511,In_1891,In_1483);
xor U512 (N_512,In_2638,In_2037);
xnor U513 (N_513,In_2437,In_1177);
and U514 (N_514,In_533,In_2197);
or U515 (N_515,In_2897,In_1828);
or U516 (N_516,N_11,In_455);
and U517 (N_517,In_2641,In_1250);
or U518 (N_518,In_1434,In_395);
xor U519 (N_519,N_112,In_160);
nor U520 (N_520,In_130,In_1707);
nand U521 (N_521,In_1962,In_149);
or U522 (N_522,In_8,In_2557);
xnor U523 (N_523,N_154,In_305);
or U524 (N_524,In_2357,N_107);
or U525 (N_525,In_2502,In_2581);
nand U526 (N_526,In_1192,In_2068);
and U527 (N_527,In_2258,In_2307);
xor U528 (N_528,In_584,In_2599);
and U529 (N_529,In_1670,In_77);
nor U530 (N_530,In_2412,In_2740);
nor U531 (N_531,N_13,In_1506);
xor U532 (N_532,In_2229,In_2492);
and U533 (N_533,N_288,In_340);
nand U534 (N_534,In_2243,In_36);
or U535 (N_535,In_1770,In_2064);
xor U536 (N_536,In_1309,In_1386);
nor U537 (N_537,In_496,In_501);
nor U538 (N_538,In_1682,In_258);
or U539 (N_539,In_1117,In_628);
xnor U540 (N_540,In_807,In_2632);
nand U541 (N_541,In_2764,In_67);
nor U542 (N_542,In_1337,In_2347);
or U543 (N_543,In_2034,In_939);
nor U544 (N_544,In_182,In_2914);
and U545 (N_545,In_618,In_1419);
nand U546 (N_546,In_2820,In_1556);
nor U547 (N_547,In_2252,In_657);
nor U548 (N_548,In_456,In_847);
xnor U549 (N_549,In_744,In_135);
or U550 (N_550,In_2876,In_300);
nor U551 (N_551,In_1905,In_1591);
and U552 (N_552,In_478,In_2245);
xor U553 (N_553,In_933,In_1147);
nand U554 (N_554,N_261,In_1623);
xnor U555 (N_555,In_166,In_2770);
xor U556 (N_556,In_17,In_2875);
nor U557 (N_557,In_1904,In_2621);
nand U558 (N_558,In_1493,In_659);
nor U559 (N_559,In_405,In_1958);
and U560 (N_560,In_930,In_1522);
xor U561 (N_561,In_2168,In_2979);
nor U562 (N_562,In_617,In_2607);
and U563 (N_563,In_2360,In_1287);
xor U564 (N_564,In_1624,In_1785);
or U565 (N_565,In_1719,In_325);
nor U566 (N_566,In_647,In_2814);
and U567 (N_567,In_850,In_1636);
nand U568 (N_568,In_1436,In_1068);
nor U569 (N_569,In_509,In_2592);
or U570 (N_570,In_728,In_2072);
nand U571 (N_571,In_518,N_93);
and U572 (N_572,In_73,In_439);
nor U573 (N_573,In_120,In_1352);
and U574 (N_574,In_2855,N_295);
nand U575 (N_575,N_134,In_779);
or U576 (N_576,In_317,In_674);
and U577 (N_577,In_275,In_1191);
or U578 (N_578,N_181,In_380);
xnor U579 (N_579,In_1246,In_190);
nor U580 (N_580,In_2405,In_489);
or U581 (N_581,In_2410,In_1220);
xnor U582 (N_582,In_237,N_223);
xor U583 (N_583,In_1091,In_1814);
nor U584 (N_584,In_2874,In_2128);
nor U585 (N_585,In_2811,In_1681);
nand U586 (N_586,In_54,In_1272);
xor U587 (N_587,In_2960,In_2047);
xor U588 (N_588,In_1886,In_1019);
xor U589 (N_589,N_63,In_2249);
nor U590 (N_590,In_797,In_676);
and U591 (N_591,In_2515,In_338);
xnor U592 (N_592,In_2173,In_786);
xnor U593 (N_593,In_508,In_531);
nand U594 (N_594,In_90,In_59);
or U595 (N_595,In_1310,N_251);
nor U596 (N_596,N_4,In_1314);
nor U597 (N_597,In_1101,In_1934);
and U598 (N_598,N_197,N_38);
and U599 (N_599,In_1223,In_2271);
and U600 (N_600,N_384,In_45);
nor U601 (N_601,In_1206,In_2976);
nor U602 (N_602,In_1124,In_2846);
nor U603 (N_603,N_151,In_225);
or U604 (N_604,In_532,N_426);
or U605 (N_605,In_1449,N_594);
and U606 (N_606,In_430,In_2566);
nor U607 (N_607,In_2254,In_366);
or U608 (N_608,N_549,In_1795);
or U609 (N_609,N_6,In_1369);
nor U610 (N_610,In_2866,In_1856);
nand U611 (N_611,In_1315,In_1532);
nand U612 (N_612,In_1514,N_231);
xnor U613 (N_613,N_416,In_345);
nor U614 (N_614,In_427,In_2120);
or U615 (N_615,In_2390,N_465);
or U616 (N_616,In_2244,N_593);
or U617 (N_617,In_2928,In_1084);
nor U618 (N_618,In_1185,In_125);
or U619 (N_619,In_1218,In_2198);
nor U620 (N_620,In_188,In_586);
and U621 (N_621,In_885,In_342);
nor U622 (N_622,In_703,In_2494);
nand U623 (N_623,In_352,In_2699);
or U624 (N_624,In_2451,In_2712);
or U625 (N_625,In_1278,In_1041);
nand U626 (N_626,N_320,N_588);
xnor U627 (N_627,In_961,In_351);
nor U628 (N_628,In_2146,In_2382);
and U629 (N_629,In_2084,In_909);
nor U630 (N_630,In_1800,In_2287);
and U631 (N_631,N_399,N_250);
nand U632 (N_632,N_130,In_2465);
nor U633 (N_633,In_156,In_2609);
nor U634 (N_634,In_1225,In_1253);
and U635 (N_635,In_1257,In_2275);
nand U636 (N_636,N_144,N_488);
or U637 (N_637,In_27,In_598);
xor U638 (N_638,In_1238,In_1186);
or U639 (N_639,In_1952,N_538);
nand U640 (N_640,In_749,In_2924);
nand U641 (N_641,In_234,In_446);
xnor U642 (N_642,In_2006,In_798);
xnor U643 (N_643,N_221,In_109);
xor U644 (N_644,In_2273,In_716);
nand U645 (N_645,In_13,N_210);
and U646 (N_646,In_2526,In_705);
nand U647 (N_647,N_192,N_95);
nor U648 (N_648,N_341,N_3);
and U649 (N_649,In_2497,N_227);
xor U650 (N_650,In_1255,In_2622);
nand U651 (N_651,N_481,In_66);
nand U652 (N_652,In_1465,In_2411);
and U653 (N_653,In_1188,In_2582);
nand U654 (N_654,In_1052,In_1595);
and U655 (N_655,N_373,In_1938);
and U656 (N_656,In_622,N_390);
xor U657 (N_657,In_2806,In_348);
or U658 (N_658,In_2346,In_888);
and U659 (N_659,In_1022,In_461);
and U660 (N_660,N_453,In_1767);
or U661 (N_661,In_1383,In_2602);
or U662 (N_662,In_2893,In_2685);
or U663 (N_663,In_2619,N_311);
or U664 (N_664,In_398,In_1577);
or U665 (N_665,In_230,In_213);
xor U666 (N_666,N_271,N_551);
or U667 (N_667,In_302,N_240);
xor U668 (N_668,In_280,N_425);
nand U669 (N_669,In_2134,In_1014);
and U670 (N_670,N_196,N_77);
or U671 (N_671,N_45,In_2311);
nand U672 (N_672,N_307,In_1667);
and U673 (N_673,N_287,N_432);
nand U674 (N_674,In_890,In_47);
nor U675 (N_675,In_2957,In_579);
nor U676 (N_676,In_1897,N_563);
xor U677 (N_677,N_126,In_1204);
nor U678 (N_678,N_595,In_129);
nand U679 (N_679,In_514,In_1050);
nor U680 (N_680,N_44,In_1411);
and U681 (N_681,In_1259,In_236);
xnor U682 (N_682,In_540,N_88);
nand U683 (N_683,In_935,In_1501);
or U684 (N_684,N_326,In_2660);
xnor U685 (N_685,In_1286,N_511);
or U686 (N_686,In_371,In_2786);
xnor U687 (N_687,In_200,In_310);
xnor U688 (N_688,In_556,In_432);
nand U689 (N_689,In_1379,In_2381);
or U690 (N_690,In_470,In_1516);
or U691 (N_691,N_449,In_1727);
or U692 (N_692,In_1712,N_565);
nand U693 (N_693,In_100,In_2643);
nor U694 (N_694,N_532,In_2636);
nand U695 (N_695,In_596,In_840);
or U696 (N_696,N_214,In_495);
xnor U697 (N_697,In_2711,In_2572);
xnor U698 (N_698,N_239,In_813);
nor U699 (N_699,In_878,In_23);
or U700 (N_700,In_1811,In_2727);
nor U701 (N_701,In_1753,In_1910);
xnor U702 (N_702,N_584,In_1088);
xor U703 (N_703,N_276,In_2612);
xnor U704 (N_704,In_2908,In_1902);
nor U705 (N_705,In_2832,In_292);
or U706 (N_706,In_2181,In_1691);
xnor U707 (N_707,In_513,In_144);
nand U708 (N_708,N_215,In_2841);
nor U709 (N_709,In_1241,In_2125);
nor U710 (N_710,In_1165,In_2595);
nand U711 (N_711,In_965,In_1903);
nor U712 (N_712,In_818,In_701);
or U713 (N_713,In_1881,In_515);
or U714 (N_714,In_2937,In_1640);
or U715 (N_715,In_401,In_492);
xor U716 (N_716,In_2276,In_1587);
or U717 (N_717,N_372,In_1421);
nor U718 (N_718,In_102,In_1579);
or U719 (N_719,N_51,N_118);
or U720 (N_720,N_370,N_212);
or U721 (N_721,In_2555,In_1380);
nor U722 (N_722,In_736,In_1184);
xor U723 (N_723,In_1213,In_591);
nor U724 (N_724,In_2471,In_512);
xor U725 (N_725,In_2237,In_2761);
xnor U726 (N_726,In_1072,N_201);
or U727 (N_727,In_2810,In_2781);
nand U728 (N_728,In_2886,In_656);
xor U729 (N_729,In_2200,In_1203);
nand U730 (N_730,In_671,In_2809);
or U731 (N_731,N_555,In_2570);
or U732 (N_732,In_1293,In_117);
nand U733 (N_733,In_1418,In_1888);
and U734 (N_734,In_37,In_855);
and U735 (N_735,In_1029,In_1179);
nor U736 (N_736,In_2050,In_449);
nor U737 (N_737,In_1092,In_1979);
xor U738 (N_738,N_472,In_2121);
nand U739 (N_739,N_79,In_1372);
nor U740 (N_740,N_466,In_638);
or U741 (N_741,N_21,N_577);
nor U742 (N_742,In_1730,In_1657);
xnor U743 (N_743,In_341,In_272);
or U744 (N_744,In_1032,In_1523);
nor U745 (N_745,In_136,In_679);
and U746 (N_746,In_1668,N_494);
nand U747 (N_747,In_70,In_2320);
nand U748 (N_748,In_2209,In_1119);
and U749 (N_749,N_195,In_113);
nand U750 (N_750,In_463,In_2199);
nand U751 (N_751,In_1163,N_429);
and U752 (N_752,In_337,In_2263);
nand U753 (N_753,In_2961,N_172);
and U754 (N_754,In_906,In_585);
and U755 (N_755,In_870,N_312);
or U756 (N_756,N_403,In_2644);
and U757 (N_757,In_499,In_560);
and U758 (N_758,In_328,In_2943);
nand U759 (N_759,In_520,In_1543);
nor U760 (N_760,In_1704,In_2744);
xnor U761 (N_761,In_2728,N_208);
xnor U762 (N_762,In_662,N_393);
nor U763 (N_763,In_2652,N_237);
nand U764 (N_764,In_733,In_1004);
xnor U765 (N_765,In_979,In_1451);
nand U766 (N_766,In_1896,N_139);
or U767 (N_767,In_1430,In_553);
nor U768 (N_768,In_2288,N_585);
xnor U769 (N_769,In_2127,In_1153);
and U770 (N_770,In_1519,In_2626);
or U771 (N_771,N_394,N_166);
or U772 (N_772,In_2507,N_281);
nor U773 (N_773,N_342,N_193);
xor U774 (N_774,In_1724,In_2055);
nand U775 (N_775,N_280,N_484);
nor U776 (N_776,In_1311,In_104);
and U777 (N_777,In_2093,In_2187);
or U778 (N_778,In_193,In_396);
xor U779 (N_779,N_184,In_604);
nand U780 (N_780,In_2941,In_1736);
nand U781 (N_781,In_1396,In_522);
nor U782 (N_782,In_2038,In_2803);
nor U783 (N_783,In_1374,In_2389);
nor U784 (N_784,In_1533,In_866);
nor U785 (N_785,In_895,In_1404);
nand U786 (N_786,In_2751,In_2456);
or U787 (N_787,In_2549,In_1565);
or U788 (N_788,N_527,N_116);
and U789 (N_789,In_1143,N_185);
xor U790 (N_790,In_2099,In_1507);
nor U791 (N_791,In_119,In_1820);
and U792 (N_792,In_2542,N_87);
nand U793 (N_793,In_500,In_2470);
nand U794 (N_794,In_2664,In_1407);
nand U795 (N_795,N_135,In_1784);
nand U796 (N_796,In_1534,N_376);
nor U797 (N_797,N_43,In_1040);
and U798 (N_798,N_148,In_1078);
or U799 (N_799,In_1936,In_2858);
and U800 (N_800,In_1190,N_80);
nand U801 (N_801,In_2104,In_2046);
or U802 (N_802,In_2571,In_437);
xor U803 (N_803,In_1098,N_170);
nand U804 (N_804,In_799,In_2545);
and U805 (N_805,In_1106,In_2467);
or U806 (N_806,In_2469,In_2261);
and U807 (N_807,In_1518,In_743);
and U808 (N_808,In_2801,In_802);
xor U809 (N_809,In_911,In_607);
xnor U810 (N_810,In_304,In_956);
and U811 (N_811,In_122,In_2624);
and U812 (N_812,N_559,In_1457);
and U813 (N_813,N_380,N_22);
nor U814 (N_814,N_508,In_2787);
and U815 (N_815,In_1169,In_1638);
xor U816 (N_816,In_2448,In_2673);
nand U817 (N_817,In_108,In_2947);
or U818 (N_818,In_758,In_1361);
or U819 (N_819,In_1666,In_2434);
nor U820 (N_820,In_460,In_1426);
or U821 (N_821,In_2348,N_92);
xnor U822 (N_822,In_2219,In_1170);
or U823 (N_823,In_79,In_2663);
nand U824 (N_824,In_2377,In_1935);
and U825 (N_825,In_468,N_344);
and U826 (N_826,In_1830,N_7);
nor U827 (N_827,In_2089,In_2512);
or U828 (N_828,In_539,In_2637);
nor U829 (N_829,In_58,In_762);
and U830 (N_830,In_894,In_2505);
or U831 (N_831,In_2391,N_378);
or U832 (N_832,In_1603,In_1663);
xor U833 (N_833,N_454,In_689);
xnor U834 (N_834,In_1136,In_529);
nand U835 (N_835,In_921,N_113);
or U836 (N_836,N_293,In_2933);
xnor U837 (N_837,In_1777,In_2297);
or U838 (N_838,In_215,In_1077);
and U839 (N_839,In_2242,In_1749);
and U840 (N_840,In_1416,N_572);
xnor U841 (N_841,In_2483,N_228);
and U842 (N_842,In_2905,In_1993);
nor U843 (N_843,N_89,In_2163);
nor U844 (N_844,N_15,In_2565);
nand U845 (N_845,In_1141,N_114);
nor U846 (N_846,In_2998,In_142);
or U847 (N_847,In_1496,In_571);
xnor U848 (N_848,In_1585,In_1750);
xnor U849 (N_849,N_8,In_519);
xor U850 (N_850,In_425,N_296);
nand U851 (N_851,In_645,In_853);
nand U852 (N_852,N_554,In_1737);
nand U853 (N_853,In_159,In_2885);
nor U854 (N_854,In_2666,N_446);
nor U855 (N_855,In_1705,In_1882);
xnor U856 (N_856,In_2425,In_1930);
xnor U857 (N_857,In_2895,N_479);
or U858 (N_858,In_2225,In_232);
nand U859 (N_859,In_1472,In_2648);
and U860 (N_860,In_2468,In_684);
nand U861 (N_861,In_551,In_1151);
nor U862 (N_862,In_1413,In_1422);
nand U863 (N_863,In_1370,In_1588);
xor U864 (N_864,In_2725,In_1619);
nand U865 (N_865,In_1508,In_838);
nand U866 (N_866,N_450,In_1156);
nand U867 (N_867,N_60,N_485);
nand U868 (N_868,In_1107,In_761);
or U869 (N_869,N_127,N_561);
or U870 (N_870,In_1701,In_162);
nand U871 (N_871,In_1135,In_99);
xor U872 (N_872,N_56,In_864);
nand U873 (N_873,N_27,In_2585);
xnor U874 (N_874,In_308,In_411);
or U875 (N_875,In_1853,N_169);
nand U876 (N_876,In_576,In_355);
and U877 (N_877,In_814,N_225);
nor U878 (N_878,In_1671,In_893);
nand U879 (N_879,In_1273,In_830);
nor U880 (N_880,In_2537,In_1381);
or U881 (N_881,N_121,In_834);
xor U882 (N_882,In_2353,In_1500);
nand U883 (N_883,In_1964,In_2009);
and U884 (N_884,In_2106,In_2732);
or U885 (N_885,In_2849,In_2863);
or U886 (N_886,In_1214,In_1937);
xnor U887 (N_887,In_2087,In_1051);
and U888 (N_888,N_156,N_343);
or U889 (N_889,In_72,In_998);
nor U890 (N_890,In_331,N_1);
nor U891 (N_891,In_1873,In_1018);
nand U892 (N_892,In_1916,In_1016);
xnor U893 (N_893,In_1827,N_305);
and U894 (N_894,In_2279,In_1675);
or U895 (N_895,In_2559,In_742);
xor U896 (N_896,In_2817,N_573);
nor U897 (N_897,In_466,In_1012);
xor U898 (N_898,In_1734,In_1291);
nor U899 (N_899,In_1263,In_589);
or U900 (N_900,In_2808,In_1747);
or U901 (N_901,In_2230,N_304);
or U902 (N_902,In_1991,In_1706);
nand U903 (N_903,In_957,N_822);
or U904 (N_904,N_413,N_626);
nor U905 (N_905,N_207,In_619);
nand U906 (N_906,N_747,In_2032);
nor U907 (N_907,In_1859,In_2692);
xor U908 (N_908,In_1709,In_2367);
nor U909 (N_909,N_233,N_760);
and U910 (N_910,In_1694,In_127);
xnor U911 (N_911,N_464,In_1425);
or U912 (N_912,In_2334,N_490);
xor U913 (N_913,In_2519,In_835);
or U914 (N_914,In_1515,In_2326);
xor U915 (N_915,N_182,In_1676);
or U916 (N_916,In_2083,In_196);
and U917 (N_917,N_109,N_310);
or U918 (N_918,N_583,In_572);
nor U919 (N_919,N_634,In_1367);
xor U920 (N_920,In_265,In_1530);
and U921 (N_921,In_1366,N_638);
nor U922 (N_922,N_269,N_846);
xor U923 (N_923,In_2079,In_1968);
nor U924 (N_924,N_150,In_1102);
or U925 (N_925,In_1900,In_107);
and U926 (N_926,In_704,In_138);
or U927 (N_927,In_2366,In_1630);
nand U928 (N_928,In_2327,In_2160);
xnor U929 (N_929,In_1837,In_996);
xor U930 (N_930,In_1110,N_252);
nand U931 (N_931,In_448,In_87);
nor U932 (N_932,In_288,In_2217);
nand U933 (N_933,In_1764,N_50);
or U934 (N_934,N_278,In_629);
xnor U935 (N_935,N_365,In_1673);
and U936 (N_936,N_478,N_421);
xnor U937 (N_937,N_898,In_504);
and U938 (N_938,N_434,In_1537);
or U939 (N_939,In_851,In_49);
xnor U940 (N_940,In_1797,In_450);
or U941 (N_941,N_805,In_1778);
and U942 (N_942,In_2376,In_2818);
nor U943 (N_943,In_465,In_126);
or U944 (N_944,In_2107,In_239);
xnor U945 (N_945,In_1821,N_292);
or U946 (N_946,In_717,In_2528);
nand U947 (N_947,In_658,N_661);
nand U948 (N_948,In_764,In_968);
nor U949 (N_949,N_600,In_2008);
nand U950 (N_950,N_820,N_665);
nor U951 (N_951,In_1985,N_290);
xnor U952 (N_952,In_2807,N_540);
xor U953 (N_953,N_862,In_7);
xnor U954 (N_954,In_2205,In_42);
nor U955 (N_955,In_2851,N_145);
nand U956 (N_956,In_1851,N_685);
xor U957 (N_957,N_406,N_386);
or U958 (N_958,In_1649,In_2416);
nor U959 (N_959,In_891,In_1011);
xor U960 (N_960,N_845,N_666);
nand U961 (N_961,N_882,In_1661);
and U962 (N_962,In_2525,In_1685);
nor U963 (N_963,In_2795,In_2342);
xor U964 (N_964,In_1596,In_2473);
or U965 (N_965,In_792,N_423);
or U966 (N_966,In_382,In_2780);
nor U967 (N_967,In_2113,In_1758);
or U968 (N_968,In_2479,In_1870);
nor U969 (N_969,In_615,In_2887);
nor U970 (N_970,In_2384,In_1867);
xnor U971 (N_971,In_915,In_2603);
xnor U972 (N_972,N_438,N_750);
and U973 (N_973,In_2714,In_55);
nor U974 (N_974,In_2836,N_701);
and U975 (N_975,N_190,In_2304);
nor U976 (N_976,N_391,N_712);
and U977 (N_977,N_767,In_1160);
and U978 (N_978,In_2018,In_2763);
and U979 (N_979,N_653,N_348);
xor U980 (N_980,In_559,N_646);
xor U981 (N_981,N_629,In_2656);
xor U982 (N_982,N_606,In_2697);
nor U983 (N_983,N_864,In_708);
or U984 (N_984,In_725,N_684);
or U985 (N_985,In_95,In_1809);
or U986 (N_986,In_1409,N_123);
xnor U987 (N_987,In_315,In_2117);
or U988 (N_988,In_1714,N_831);
nor U989 (N_989,N_533,In_2819);
or U990 (N_990,N_440,In_242);
and U991 (N_991,In_1593,In_1129);
nand U992 (N_992,In_2005,In_2681);
or U993 (N_993,In_2812,N_336);
and U994 (N_994,In_2371,N_576);
or U995 (N_995,N_229,N_179);
or U996 (N_996,In_2404,In_2554);
and U997 (N_997,In_12,In_982);
or U998 (N_998,In_609,N_837);
nand U999 (N_999,N_832,In_1763);
nor U1000 (N_1000,In_477,In_857);
nor U1001 (N_1001,In_2990,In_2823);
and U1002 (N_1002,In_2248,In_447);
or U1003 (N_1003,N_821,In_880);
or U1004 (N_1004,N_632,In_1433);
and U1005 (N_1005,In_1690,In_19);
and U1006 (N_1006,In_397,N_641);
xnor U1007 (N_1007,In_575,N_443);
nand U1008 (N_1008,N_128,In_1318);
nor U1009 (N_1009,In_1807,In_2827);
xor U1010 (N_1010,N_23,N_205);
nor U1011 (N_1011,N_473,In_2020);
nor U1012 (N_1012,N_73,In_2421);
nor U1013 (N_1013,In_1393,In_2223);
or U1014 (N_1014,In_2538,N_762);
and U1015 (N_1015,In_1494,N_39);
nand U1016 (N_1016,N_807,In_602);
nand U1017 (N_1017,In_2616,In_1015);
nand U1018 (N_1018,In_912,N_517);
and U1019 (N_1019,N_887,N_878);
nor U1020 (N_1020,N_753,N_408);
xor U1021 (N_1021,In_403,In_2289);
nor U1022 (N_1022,In_613,In_1277);
or U1023 (N_1023,In_929,In_378);
or U1024 (N_1024,In_984,In_1798);
and U1025 (N_1025,In_960,In_1066);
nor U1026 (N_1026,In_2312,In_1606);
xnor U1027 (N_1027,In_2208,N_655);
and U1028 (N_1028,N_796,In_388);
nand U1029 (N_1029,In_210,N_794);
nor U1030 (N_1030,In_1276,In_530);
nor U1031 (N_1031,In_240,N_748);
xor U1032 (N_1032,In_2831,In_2869);
nand U1033 (N_1033,In_2129,N_681);
nor U1034 (N_1034,N_592,In_685);
nand U1035 (N_1035,N_441,In_781);
and U1036 (N_1036,In_2004,N_671);
or U1037 (N_1037,N_35,N_596);
nor U1038 (N_1038,N_741,In_1226);
and U1039 (N_1039,In_819,In_2816);
or U1040 (N_1040,N_546,N_614);
and U1041 (N_1041,In_187,N_451);
nor U1042 (N_1042,N_853,In_2509);
and U1043 (N_1043,N_718,N_842);
or U1044 (N_1044,In_1861,In_1761);
nand U1045 (N_1045,N_689,In_91);
and U1046 (N_1046,N_766,N_125);
nor U1047 (N_1047,In_2340,In_1000);
or U1048 (N_1048,In_244,In_603);
xor U1049 (N_1049,In_199,N_784);
nand U1050 (N_1050,In_34,N_26);
nor U1051 (N_1051,In_2888,In_2284);
xor U1052 (N_1052,In_2491,N_176);
nor U1053 (N_1053,In_1862,In_2238);
xnor U1054 (N_1054,N_844,In_1008);
nor U1055 (N_1055,N_812,In_1787);
nand U1056 (N_1056,In_279,In_467);
nand U1057 (N_1057,In_2080,N_803);
and U1058 (N_1058,In_462,N_698);
nand U1059 (N_1059,N_682,In_550);
or U1060 (N_1060,In_472,In_995);
or U1061 (N_1061,In_114,N_649);
nand U1062 (N_1062,N_792,In_231);
nor U1063 (N_1063,In_2157,N_793);
xor U1064 (N_1064,In_424,In_334);
xnor U1065 (N_1065,In_429,In_1420);
nand U1066 (N_1066,In_2179,In_50);
nand U1067 (N_1067,N_279,N_867);
nor U1068 (N_1068,In_295,In_2829);
nand U1069 (N_1069,N_436,N_662);
nand U1070 (N_1070,N_469,N_136);
xnor U1071 (N_1071,In_1757,N_660);
nor U1072 (N_1072,N_679,N_849);
or U1073 (N_1073,N_447,In_1578);
nor U1074 (N_1074,In_1262,In_1885);
xnor U1075 (N_1075,In_1164,In_1715);
xnor U1076 (N_1076,N_506,N_830);
xor U1077 (N_1077,In_542,In_2299);
or U1078 (N_1078,In_391,In_1275);
and U1079 (N_1079,N_860,N_571);
xnor U1080 (N_1080,In_1781,N_770);
xor U1081 (N_1081,In_1445,N_337);
nand U1082 (N_1082,In_2671,In_2604);
nor U1083 (N_1083,In_178,N_786);
nand U1084 (N_1084,N_10,In_2296);
and U1085 (N_1085,In_2308,N_18);
nand U1086 (N_1086,In_714,In_1544);
or U1087 (N_1087,In_631,N_360);
nor U1088 (N_1088,In_416,In_253);
xnor U1089 (N_1089,In_1846,In_2042);
nand U1090 (N_1090,In_2433,N_69);
and U1091 (N_1091,N_325,In_2272);
or U1092 (N_1092,In_648,N_165);
nand U1093 (N_1093,In_1131,In_2676);
and U1094 (N_1094,In_510,In_691);
and U1095 (N_1095,In_1261,In_105);
xnor U1096 (N_1096,In_632,In_2535);
xnor U1097 (N_1097,In_2374,In_1122);
xor U1098 (N_1098,In_1319,In_1776);
nand U1099 (N_1099,In_826,N_350);
nor U1100 (N_1100,N_496,N_258);
nand U1101 (N_1101,In_481,N_309);
xnor U1102 (N_1102,N_818,N_605);
nand U1103 (N_1103,In_770,In_583);
and U1104 (N_1104,In_760,In_1994);
xor U1105 (N_1105,N_695,In_243);
and U1106 (N_1106,N_761,In_282);
nor U1107 (N_1107,In_86,In_63);
xnor U1108 (N_1108,In_438,In_2845);
and U1109 (N_1109,N_871,N_407);
and U1110 (N_1110,In_1298,In_2894);
or U1111 (N_1111,N_888,N_514);
xnor U1112 (N_1112,In_2805,In_2356);
nand U1113 (N_1113,In_2122,N_275);
and U1114 (N_1114,In_51,In_1159);
nand U1115 (N_1115,N_580,In_528);
and U1116 (N_1116,N_659,In_2902);
nand U1117 (N_1117,N_619,In_2012);
nand U1118 (N_1118,In_2343,In_2461);
nand U1119 (N_1119,In_1069,In_227);
nor U1120 (N_1120,N_351,In_723);
or U1121 (N_1121,In_1627,In_2500);
and U1122 (N_1122,In_975,In_220);
nor U1123 (N_1123,N_881,N_819);
xnor U1124 (N_1124,In_2337,N_765);
xor U1125 (N_1125,N_392,In_2154);
and U1126 (N_1126,In_1729,In_2019);
xnor U1127 (N_1127,In_2981,In_1997);
nor U1128 (N_1128,In_1974,In_2857);
or U1129 (N_1129,In_443,In_2235);
xor U1130 (N_1130,In_993,N_298);
xor U1131 (N_1131,N_847,In_587);
xnor U1132 (N_1132,In_2882,N_83);
and U1133 (N_1133,N_528,N_230);
nand U1134 (N_1134,In_2166,In_2601);
and U1135 (N_1135,N_72,In_934);
nor U1136 (N_1136,In_2657,N_115);
and U1137 (N_1137,In_2700,In_732);
nor U1138 (N_1138,N_104,N_198);
or U1139 (N_1139,In_2743,In_2653);
and U1140 (N_1140,In_2105,N_520);
nand U1141 (N_1141,N_875,In_1716);
or U1142 (N_1142,N_168,In_2277);
or U1143 (N_1143,In_2533,In_56);
xnor U1144 (N_1144,N_34,In_1414);
nand U1145 (N_1145,In_1235,N_498);
nor U1146 (N_1146,In_1350,In_2103);
xor U1147 (N_1147,In_2116,In_2069);
or U1148 (N_1148,N_338,N_601);
nand U1149 (N_1149,N_470,In_2710);
nor U1150 (N_1150,N_289,In_1100);
or U1151 (N_1151,In_139,In_2680);
nor U1152 (N_1152,In_2618,N_510);
or U1153 (N_1153,In_773,In_715);
xnor U1154 (N_1154,In_681,In_1471);
nand U1155 (N_1155,In_2139,N_759);
nor U1156 (N_1156,N_140,N_705);
xor U1157 (N_1157,In_2587,N_564);
nor U1158 (N_1158,In_1212,In_313);
or U1159 (N_1159,N_331,In_1391);
xor U1160 (N_1160,In_106,In_2733);
and U1161 (N_1161,N_110,In_1290);
nor U1162 (N_1162,N_611,In_2265);
and U1163 (N_1163,N_188,In_2322);
or U1164 (N_1164,In_555,In_1725);
xnor U1165 (N_1165,N_455,In_2580);
and U1166 (N_1166,In_2825,N_841);
nand U1167 (N_1167,In_1095,In_1849);
and U1168 (N_1168,N_433,In_2193);
nor U1169 (N_1169,In_31,In_2591);
nand U1170 (N_1170,In_137,In_2707);
nor U1171 (N_1171,N_835,In_290);
nand U1172 (N_1172,N_226,In_2291);
nor U1173 (N_1173,N_547,In_2486);
xor U1174 (N_1174,N_333,In_1438);
or U1175 (N_1175,In_1567,In_2153);
or U1176 (N_1176,In_2250,In_2935);
or U1177 (N_1177,In_2145,In_823);
nor U1178 (N_1178,In_1327,In_610);
and U1179 (N_1179,In_1847,In_1316);
and U1180 (N_1180,In_293,In_1838);
xnor U1181 (N_1181,N_893,In_1527);
xor U1182 (N_1182,In_910,In_387);
and U1183 (N_1183,In_1509,In_2815);
nand U1184 (N_1184,In_2317,In_2143);
xor U1185 (N_1185,N_356,N_180);
or U1186 (N_1186,In_817,N_17);
and U1187 (N_1187,N_9,In_1969);
or U1188 (N_1188,In_192,In_1525);
xnor U1189 (N_1189,In_1482,N_531);
nor U1190 (N_1190,N_861,N_534);
nand U1191 (N_1191,In_2861,In_1972);
and U1192 (N_1192,In_2227,In_777);
nand U1193 (N_1193,N_872,In_625);
or U1194 (N_1194,In_2495,In_226);
nand U1195 (N_1195,In_1549,In_2503);
xnor U1196 (N_1196,In_421,In_1655);
xor U1197 (N_1197,In_2800,In_65);
nor U1198 (N_1198,N_850,In_608);
nand U1199 (N_1199,In_2262,N_270);
xnor U1200 (N_1200,In_2278,In_2010);
nor U1201 (N_1201,In_1561,N_238);
or U1202 (N_1202,N_243,N_961);
nand U1203 (N_1203,In_2114,N_776);
nor U1204 (N_1204,N_1035,N_313);
xnor U1205 (N_1205,N_994,In_1860);
or U1206 (N_1206,N_636,N_460);
xnor U1207 (N_1207,N_667,In_2457);
nand U1208 (N_1208,N_918,In_1559);
xnor U1209 (N_1209,In_2213,In_1654);
and U1210 (N_1210,N_418,In_1013);
and U1211 (N_1211,In_1835,In_731);
or U1212 (N_1212,N_1171,In_946);
and U1213 (N_1213,In_1166,In_150);
or U1214 (N_1214,In_2900,In_1769);
and U1215 (N_1215,N_755,In_281);
nand U1216 (N_1216,In_2292,N_515);
and U1217 (N_1217,N_787,In_1894);
or U1218 (N_1218,In_148,N_86);
and U1219 (N_1219,N_503,In_233);
nand U1220 (N_1220,N_771,In_2796);
xor U1221 (N_1221,N_799,N_155);
nand U1222 (N_1222,N_633,In_611);
nor U1223 (N_1223,N_463,In_517);
xor U1224 (N_1224,In_1976,N_146);
or U1225 (N_1225,In_1550,In_2368);
nor U1226 (N_1226,In_875,N_315);
and U1227 (N_1227,In_959,N_749);
nand U1228 (N_1228,N_412,In_2417);
xor U1229 (N_1229,In_319,In_928);
nor U1230 (N_1230,N_541,N_1118);
or U1231 (N_1231,N_152,N_657);
and U1232 (N_1232,N_1170,In_1406);
or U1233 (N_1233,N_651,In_256);
nor U1234 (N_1234,N_589,N_1056);
nand U1235 (N_1235,In_1285,In_1450);
nor U1236 (N_1236,N_1120,N_991);
nor U1237 (N_1237,In_1789,N_725);
or U1238 (N_1238,N_903,In_485);
xor U1239 (N_1239,In_11,In_1639);
xor U1240 (N_1240,In_896,N_42);
xnor U1241 (N_1241,In_1046,In_1780);
nand U1242 (N_1242,In_1328,In_1476);
nand U1243 (N_1243,N_431,N_1136);
nand U1244 (N_1244,N_358,In_426);
xnor U1245 (N_1245,In_2936,N_590);
nand U1246 (N_1246,In_901,In_606);
or U1247 (N_1247,N_1043,In_255);
nand U1248 (N_1248,N_1014,N_430);
nand U1249 (N_1249,In_1395,N_1048);
nand U1250 (N_1250,N_33,N_979);
nand U1251 (N_1251,In_2548,N_703);
or U1252 (N_1252,N_947,N_1154);
xnor U1253 (N_1253,In_1892,In_2303);
nand U1254 (N_1254,In_2723,N_1030);
and U1255 (N_1255,N_945,In_2785);
and U1256 (N_1256,In_1057,N_427);
nor U1257 (N_1257,N_1132,In_414);
nand U1258 (N_1258,In_2414,In_2407);
xnor U1259 (N_1259,In_212,In_865);
nand U1260 (N_1260,N_291,N_91);
xor U1261 (N_1261,N_752,In_917);
nor U1262 (N_1262,In_2967,N_938);
nor U1263 (N_1263,N_401,N_768);
xnor U1264 (N_1264,In_2316,N_411);
nand U1265 (N_1265,In_936,N_509);
nand U1266 (N_1266,N_111,N_442);
nor U1267 (N_1267,In_1456,N_1108);
xor U1268 (N_1268,N_568,N_900);
nor U1269 (N_1269,In_1295,N_998);
and U1270 (N_1270,In_1410,In_1679);
and U1271 (N_1271,In_1140,N_1080);
and U1272 (N_1272,N_683,In_2294);
nor U1273 (N_1273,N_1070,In_2339);
xnor U1274 (N_1274,In_2524,In_2917);
xor U1275 (N_1275,N_492,N_163);
nor U1276 (N_1276,N_458,N_1112);
and U1277 (N_1277,N_567,In_2395);
nor U1278 (N_1278,N_1157,In_442);
and U1279 (N_1279,In_737,N_260);
and U1280 (N_1280,In_1044,In_2513);
nor U1281 (N_1281,In_2828,In_1582);
and U1282 (N_1282,In_2351,In_1786);
nand U1283 (N_1283,In_2180,In_169);
or U1284 (N_1284,In_2726,In_2771);
or U1285 (N_1285,In_948,In_2776);
nand U1286 (N_1286,N_1188,In_1826);
nand U1287 (N_1287,In_2556,In_2345);
nor U1288 (N_1288,N_167,N_199);
xor U1289 (N_1289,N_824,In_2364);
xnor U1290 (N_1290,N_1152,In_663);
or U1291 (N_1291,N_797,In_435);
nand U1292 (N_1292,In_844,N_396);
and U1293 (N_1293,In_1840,In_241);
nor U1294 (N_1294,N_117,N_1077);
and U1295 (N_1295,N_728,N_714);
nor U1296 (N_1296,In_2879,In_174);
xnor U1297 (N_1297,In_18,In_573);
and U1298 (N_1298,N_461,N_645);
nor U1299 (N_1299,In_1708,In_9);
nand U1300 (N_1300,N_644,N_328);
and U1301 (N_1301,N_1151,In_415);
and U1302 (N_1302,N_65,In_1912);
and U1303 (N_1303,N_424,N_631);
or U1304 (N_1304,In_1071,In_1563);
or U1305 (N_1305,N_874,In_860);
xor U1306 (N_1306,In_2708,In_1768);
nor U1307 (N_1307,In_1010,In_412);
xor U1308 (N_1308,N_353,In_566);
nand U1309 (N_1309,In_707,N_1069);
nor U1310 (N_1310,N_866,N_1006);
or U1311 (N_1311,N_46,N_920);
or U1312 (N_1312,N_675,In_433);
nor U1313 (N_1313,N_734,In_2737);
or U1314 (N_1314,N_731,N_814);
or U1315 (N_1315,In_1925,N_813);
xnor U1316 (N_1316,N_630,In_370);
or U1317 (N_1317,In_1398,In_776);
or U1318 (N_1318,N_255,In_1076);
or U1319 (N_1319,N_1004,N_263);
xor U1320 (N_1320,N_164,In_2691);
and U1321 (N_1321,In_2682,In_1576);
nand U1322 (N_1322,In_2144,N_857);
nand U1323 (N_1323,In_2496,In_2313);
nor U1324 (N_1324,In_2931,In_482);
nor U1325 (N_1325,N_61,N_1082);
nor U1326 (N_1326,N_1173,In_2649);
xnor U1327 (N_1327,In_713,In_1061);
xnor U1328 (N_1328,N_859,N_483);
xor U1329 (N_1329,N_949,In_1617);
nor U1330 (N_1330,In_78,In_1108);
xnor U1331 (N_1331,In_316,In_2256);
and U1332 (N_1332,In_882,N_204);
xor U1333 (N_1333,N_723,In_2610);
or U1334 (N_1334,In_2220,In_1363);
nand U1335 (N_1335,In_2400,N_791);
or U1336 (N_1336,In_132,N_668);
nor U1337 (N_1337,N_476,In_561);
or U1338 (N_1338,In_2954,N_673);
nand U1339 (N_1339,N_740,In_1299);
or U1340 (N_1340,N_856,In_1520);
and U1341 (N_1341,In_2403,In_1967);
nor U1342 (N_1342,In_614,In_1200);
or U1343 (N_1343,In_64,N_1052);
and U1344 (N_1344,N_628,N_598);
xor U1345 (N_1345,In_383,N_377);
nand U1346 (N_1346,N_301,In_1539);
xor U1347 (N_1347,N_1057,In_653);
xnor U1348 (N_1348,In_229,In_1660);
nand U1349 (N_1349,N_1127,In_2904);
and U1350 (N_1350,In_2472,N_877);
and U1351 (N_1351,In_981,In_2172);
nand U1352 (N_1352,N_996,In_2086);
nor U1353 (N_1353,In_1552,In_842);
nor U1354 (N_1354,In_2397,In_164);
xnor U1355 (N_1355,In_2090,In_1339);
nor U1356 (N_1356,N_1002,N_773);
nor U1357 (N_1357,In_1267,N_268);
xor U1358 (N_1358,In_805,N_948);
xor U1359 (N_1359,In_1149,N_566);
and U1360 (N_1360,N_1113,N_1102);
and U1361 (N_1361,In_2236,N_910);
nor U1362 (N_1362,N_1149,N_53);
nor U1363 (N_1363,N_924,In_1586);
xnor U1364 (N_1364,In_1053,In_1583);
nand U1365 (N_1365,N_400,In_2266);
nor U1366 (N_1366,In_670,In_2149);
and U1367 (N_1367,N_1083,N_395);
and U1368 (N_1368,In_2959,N_574);
and U1369 (N_1369,In_2783,N_708);
or U1370 (N_1370,In_748,N_978);
and U1371 (N_1371,N_62,In_1382);
and U1372 (N_1372,In_1680,N_702);
xnor U1373 (N_1373,N_1047,N_318);
xor U1374 (N_1374,N_375,N_680);
xor U1375 (N_1375,In_778,In_767);
or U1376 (N_1376,In_931,In_1933);
or U1377 (N_1377,In_2234,N_1100);
nand U1378 (N_1378,N_914,In_1237);
nor U1379 (N_1379,N_811,In_2011);
nand U1380 (N_1380,N_935,N_627);
and U1381 (N_1381,N_1003,In_2349);
nor U1382 (N_1382,In_2196,N_727);
and U1383 (N_1383,N_1040,In_2717);
nor U1384 (N_1384,N_779,In_1594);
nand U1385 (N_1385,In_1779,N_330);
nand U1386 (N_1386,N_674,N_20);
or U1387 (N_1387,In_2698,N_757);
or U1388 (N_1388,In_2877,N_522);
nand U1389 (N_1389,In_335,In_2078);
nor U1390 (N_1390,In_30,In_1187);
or U1391 (N_1391,In_2605,N_624);
and U1392 (N_1392,In_1818,In_1459);
or U1393 (N_1393,In_726,N_357);
and U1394 (N_1394,N_1064,In_741);
nor U1395 (N_1395,N_75,In_62);
nor U1396 (N_1396,In_1189,In_1911);
nor U1397 (N_1397,In_2750,In_816);
nor U1398 (N_1398,N_622,In_2358);
xnor U1399 (N_1399,N_367,N_980);
nor U1400 (N_1400,In_2668,In_1222);
xor U1401 (N_1401,In_1244,N_1199);
and U1402 (N_1402,N_362,N_984);
or U1403 (N_1403,In_1609,N_892);
nor U1404 (N_1404,In_1791,In_2842);
nand U1405 (N_1405,N_550,In_2968);
and U1406 (N_1406,N_670,In_2748);
nand U1407 (N_1407,In_1294,N_863);
nor U1408 (N_1408,In_1266,N_68);
nor U1409 (N_1409,N_435,In_1528);
nor U1410 (N_1410,In_810,In_1927);
or U1411 (N_1411,In_590,N_1065);
nor U1412 (N_1412,In_228,In_712);
nand U1413 (N_1413,N_1041,In_720);
nor U1414 (N_1414,N_347,In_459);
nor U1415 (N_1415,In_599,In_1816);
xor U1416 (N_1416,In_544,In_2211);
xor U1417 (N_1417,N_474,N_1097);
xnor U1418 (N_1418,N_1187,In_1558);
and U1419 (N_1419,N_781,N_891);
and U1420 (N_1420,In_2949,In_2002);
nand U1421 (N_1421,In_952,N_942);
or U1422 (N_1422,N_70,N_963);
or U1423 (N_1423,N_102,In_46);
and U1424 (N_1424,In_869,In_2837);
or U1425 (N_1425,N_1092,In_2693);
and U1426 (N_1426,In_1121,In_2118);
and U1427 (N_1427,In_903,N_487);
xor U1428 (N_1428,N_658,N_954);
nand U1429 (N_1429,N_272,N_722);
nor U1430 (N_1430,In_664,In_2584);
xnor U1431 (N_1431,N_1139,N_699);
or U1432 (N_1432,N_962,In_661);
or U1433 (N_1433,In_1402,In_1717);
and U1434 (N_1434,N_398,N_1051);
or U1435 (N_1435,N_505,In_2239);
xor U1436 (N_1436,N_816,N_922);
nand U1437 (N_1437,In_872,N_804);
or U1438 (N_1438,In_621,In_1009);
or U1439 (N_1439,In_696,In_2443);
and U1440 (N_1440,N_828,In_249);
nor U1441 (N_1441,In_2970,N_579);
xnor U1442 (N_1442,In_2738,N_1160);
and U1443 (N_1443,In_2773,N_415);
or U1444 (N_1444,N_886,N_81);
nand U1445 (N_1445,In_785,In_751);
xnor U1446 (N_1446,In_476,N_241);
xor U1447 (N_1447,In_1168,N_521);
and U1448 (N_1448,In_1428,N_973);
xor U1449 (N_1449,In_2155,In_829);
and U1450 (N_1450,In_1618,In_1210);
and U1451 (N_1451,In_2942,N_129);
and U1452 (N_1452,In_1417,In_264);
nor U1453 (N_1453,In_2182,N_927);
or U1454 (N_1454,N_1078,In_2007);
xor U1455 (N_1455,In_1686,N_529);
nor U1456 (N_1456,In_2675,In_1703);
nand U1457 (N_1457,In_2862,In_2022);
nand U1458 (N_1458,In_2617,N_194);
nand U1459 (N_1459,In_1760,N_507);
xor U1460 (N_1460,N_697,In_1963);
or U1461 (N_1461,N_1045,In_881);
nor U1462 (N_1462,N_1142,N_1074);
or U1463 (N_1463,N_1125,In_1613);
xnor U1464 (N_1464,In_2952,N_704);
xnor U1465 (N_1465,N_613,N_720);
nor U1466 (N_1466,In_831,N_933);
xnor U1467 (N_1467,In_146,In_2768);
nand U1468 (N_1468,In_2852,In_1002);
xnor U1469 (N_1469,In_2561,N_445);
xnor U1470 (N_1470,N_967,N_810);
nand U1471 (N_1471,N_716,N_59);
or U1472 (N_1472,N_202,In_1470);
nor U1473 (N_1473,N_1179,In_1547);
xnor U1474 (N_1474,In_297,N_843);
xor U1475 (N_1475,N_1079,In_2462);
and U1476 (N_1476,N_960,In_1251);
nor U1477 (N_1477,N_1198,N_67);
and U1478 (N_1478,N_1185,In_2482);
nor U1479 (N_1479,N_726,N_48);
nand U1480 (N_1480,In_1510,In_1064);
nand U1481 (N_1481,N_777,N_314);
nor U1482 (N_1482,N_1090,In_1970);
nand U1483 (N_1483,In_534,In_700);
xnor U1484 (N_1484,In_2300,In_2639);
or U1485 (N_1485,In_2916,N_1099);
or U1486 (N_1486,N_480,In_1349);
nand U1487 (N_1487,N_277,N_1038);
xor U1488 (N_1488,In_1358,N_587);
nor U1489 (N_1489,In_1855,In_806);
nor U1490 (N_1490,In_1504,N_772);
and U1491 (N_1491,In_2126,N_1022);
nand U1492 (N_1492,In_2925,N_1053);
nor U1493 (N_1493,N_1146,N_371);
or U1494 (N_1494,In_918,N_717);
nand U1495 (N_1495,In_469,In_1474);
nor U1496 (N_1496,N_1095,N_1049);
nand U1497 (N_1497,N_743,In_1075);
nand U1498 (N_1498,In_570,In_1109);
nor U1499 (N_1499,In_2088,N_1091);
nor U1500 (N_1500,N_1168,N_719);
or U1501 (N_1501,N_1362,In_1458);
xnor U1502 (N_1502,In_1641,In_677);
nor U1503 (N_1503,In_2447,In_1918);
xor U1504 (N_1504,In_251,N_1075);
xor U1505 (N_1505,In_1740,N_955);
and U1506 (N_1506,In_254,N_647);
and U1507 (N_1507,In_320,In_2929);
and U1508 (N_1508,N_1332,N_1156);
nor U1509 (N_1509,In_369,N_939);
and U1510 (N_1510,In_394,N_1184);
nand U1511 (N_1511,In_1435,N_739);
nor U1512 (N_1512,In_2984,N_688);
nand U1513 (N_1513,In_1446,In_1440);
nor U1514 (N_1514,N_1042,In_2517);
nand U1515 (N_1515,N_383,In_185);
nor U1516 (N_1516,N_316,In_1978);
or U1517 (N_1517,In_900,In_2431);
and U1518 (N_1518,N_1318,In_2799);
nand U1519 (N_1519,N_247,N_1265);
or U1520 (N_1520,N_55,In_1461);
and U1521 (N_1521,In_1431,N_1394);
and U1522 (N_1522,N_1238,In_1093);
and U1523 (N_1523,N_908,In_873);
nand U1524 (N_1524,In_1467,In_2695);
and U1525 (N_1525,In_690,N_956);
nor U1526 (N_1526,N_1479,In_2318);
nand U1527 (N_1527,N_1480,N_873);
or U1528 (N_1528,N_1195,N_1458);
nand U1529 (N_1529,In_1773,In_562);
nand U1530 (N_1530,N_452,In_2001);
nand U1531 (N_1531,In_1498,In_2920);
nor U1532 (N_1532,N_1388,In_624);
xnor U1533 (N_1533,N_160,N_1435);
or U1534 (N_1534,N_907,N_737);
or U1535 (N_1535,N_345,In_825);
or U1536 (N_1536,In_2527,N_623);
or U1537 (N_1537,N_1135,In_330);
and U1538 (N_1538,In_235,N_894);
xnor U1539 (N_1539,In_285,In_2985);
and U1540 (N_1540,In_1815,In_2309);
nor U1541 (N_1541,N_1444,N_642);
nor U1542 (N_1542,In_140,In_2408);
or U1543 (N_1543,In_2178,N_1443);
nand U1544 (N_1544,N_1340,N_1291);
or U1545 (N_1545,N_1401,In_1901);
nor U1546 (N_1546,In_2097,In_454);
and U1547 (N_1547,N_1115,In_75);
nand U1548 (N_1548,In_2100,N_902);
nand U1549 (N_1549,In_1157,N_944);
and U1550 (N_1550,N_815,In_1946);
xnor U1551 (N_1551,In_2475,In_2102);
and U1552 (N_1552,N_1147,N_359);
or U1553 (N_1553,N_756,In_724);
nand U1554 (N_1554,In_121,In_2594);
xor U1555 (N_1555,In_2175,N_556);
or U1556 (N_1556,In_1207,N_500);
or U1557 (N_1557,In_1647,N_1417);
or U1558 (N_1558,In_269,N_444);
xor U1559 (N_1559,N_1266,N_1236);
nor U1560 (N_1560,N_928,N_1104);
nand U1561 (N_1561,N_795,In_2611);
nand U1562 (N_1562,N_122,In_755);
xor U1563 (N_1563,N_1144,In_1689);
xor U1564 (N_1564,N_1162,N_1071);
or U1565 (N_1565,In_2477,In_238);
xor U1566 (N_1566,N_535,In_1928);
or U1567 (N_1567,In_39,N_560);
or U1568 (N_1568,In_2095,In_2898);
nor U1569 (N_1569,N_300,In_1221);
and U1570 (N_1570,N_1126,N_1111);
nor U1571 (N_1571,N_557,In_2579);
xor U1572 (N_1572,In_283,In_1924);
nor U1573 (N_1573,N_189,In_43);
and U1574 (N_1574,N_1379,In_1279);
nand U1575 (N_1575,In_2945,In_2282);
and U1576 (N_1576,N_518,In_2950);
or U1577 (N_1577,In_216,N_419);
nand U1578 (N_1578,N_1381,In_464);
nor U1579 (N_1579,In_2286,In_1454);
xnor U1580 (N_1580,N_1203,N_1096);
and U1581 (N_1581,N_1153,N_1334);
and U1582 (N_1582,In_2778,N_974);
and U1583 (N_1583,N_1084,N_459);
nand U1584 (N_1584,In_2864,In_1490);
nor U1585 (N_1585,N_782,N_324);
nor U1586 (N_1586,N_1143,In_595);
nand U1587 (N_1587,N_1450,In_2999);
and U1588 (N_1588,N_1211,N_780);
nand U1589 (N_1589,N_729,In_978);
xnor U1590 (N_1590,N_74,In_1388);
and U1591 (N_1591,N_1009,In_1116);
or U1592 (N_1592,N_1487,N_1032);
xnor U1593 (N_1593,In_966,N_1013);
nor U1594 (N_1594,N_951,N_1421);
xnor U1595 (N_1595,N_389,In_2392);
and U1596 (N_1596,N_929,In_1427);
nand U1597 (N_1597,N_1399,N_575);
nor U1598 (N_1598,N_746,In_821);
nor U1599 (N_1599,In_1489,N_410);
nor U1600 (N_1600,N_1208,In_1642);
and U1601 (N_1601,N_789,N_14);
or U1602 (N_1602,N_1346,N_1445);
and U1603 (N_1603,In_702,In_2973);
xor U1604 (N_1604,In_2430,N_764);
xnor U1605 (N_1605,In_2385,N_1296);
or U1606 (N_1606,In_1099,In_29);
nor U1607 (N_1607,In_1224,N_1129);
or U1608 (N_1608,N_976,N_1233);
and U1609 (N_1609,N_1192,In_1021);
or U1610 (N_1610,In_526,In_568);
and U1611 (N_1611,N_952,In_1464);
xor U1612 (N_1612,In_2683,In_2453);
xnor U1613 (N_1613,In_2216,N_1110);
or U1614 (N_1614,N_943,N_1380);
or U1615 (N_1615,N_1018,In_327);
xnor U1616 (N_1616,N_329,In_2201);
nor U1617 (N_1617,N_1121,In_2762);
xor U1618 (N_1618,In_1631,N_696);
nand U1619 (N_1619,In_2232,In_1842);
nand U1620 (N_1620,N_1365,In_368);
nor U1621 (N_1621,In_81,In_1439);
nand U1622 (N_1622,N_1465,N_24);
and U1623 (N_1623,In_2045,In_21);
xor U1624 (N_1624,In_1080,N_82);
or U1625 (N_1625,N_620,N_1437);
or U1626 (N_1626,N_209,N_525);
xnor U1627 (N_1627,In_2777,N_1495);
and U1628 (N_1628,N_1363,In_2206);
xor U1629 (N_1629,In_74,In_1199);
xnor U1630 (N_1630,N_249,In_1256);
nand U1631 (N_1631,In_554,N_387);
xor U1632 (N_1632,In_2501,N_203);
xnor U1633 (N_1633,N_1088,N_678);
xor U1634 (N_1634,In_306,In_967);
nor U1635 (N_1635,In_418,N_99);
nor U1636 (N_1636,N_1345,N_1400);
nor U1637 (N_1637,N_1473,N_1007);
xor U1638 (N_1638,In_1656,In_2757);
nor U1639 (N_1639,N_468,N_1410);
xor U1640 (N_1640,In_2075,In_867);
nand U1641 (N_1641,In_1698,N_1485);
xor U1642 (N_1642,N_1423,N_1271);
nor U1643 (N_1643,In_2195,N_1449);
nand U1644 (N_1644,N_790,N_162);
or U1645 (N_1645,N_340,In_1898);
nor U1646 (N_1646,N_1315,In_1202);
or U1647 (N_1647,N_1408,In_1615);
nand U1648 (N_1648,In_524,In_1996);
nand U1649 (N_1649,N_972,In_1922);
xnor U1650 (N_1650,In_627,In_1415);
nand U1651 (N_1651,N_693,In_2189);
or U1652 (N_1652,N_1277,N_334);
nor U1653 (N_1653,In_942,In_1822);
and U1654 (N_1654,N_895,In_1281);
nor U1655 (N_1655,N_1248,N_1189);
nand U1656 (N_1656,N_1264,In_1283);
or U1657 (N_1657,N_1251,N_1060);
nor U1658 (N_1658,In_167,N_1062);
xnor U1659 (N_1659,In_2540,N_1481);
nor U1660 (N_1660,N_404,In_1535);
xor U1661 (N_1661,In_1738,N_694);
nor U1662 (N_1662,In_1048,N_153);
or U1663 (N_1663,N_1493,In_552);
or U1664 (N_1664,In_549,N_1462);
xor U1665 (N_1665,N_1178,In_535);
or U1666 (N_1666,In_2865,In_987);
xor U1667 (N_1667,N_1194,In_332);
and U1668 (N_1668,N_552,N_1158);
nor U1669 (N_1669,N_1159,In_111);
nor U1670 (N_1670,In_20,N_840);
nor U1671 (N_1671,In_1113,N_41);
and U1672 (N_1672,N_1137,N_103);
xnor U1673 (N_1673,In_1408,In_1322);
nand U1674 (N_1674,N_1260,In_2977);
and U1675 (N_1675,In_133,N_1311);
nand U1676 (N_1676,N_1175,N_742);
xor U1677 (N_1677,In_2539,N_523);
nor U1678 (N_1678,N_855,N_462);
nor U1679 (N_1679,N_1411,N_1464);
nor U1680 (N_1680,N_1010,In_1908);
or U1681 (N_1681,N_1374,In_2583);
nand U1682 (N_1682,In_970,N_1275);
and U1683 (N_1683,In_2989,In_2880);
xnor U1684 (N_1684,N_1256,N_267);
and U1685 (N_1685,In_1718,N_1310);
and U1686 (N_1686,N_495,In_1158);
nand U1687 (N_1687,N_220,N_582);
nor U1688 (N_1688,In_1771,N_1098);
nand U1689 (N_1689,N_603,In_772);
or U1690 (N_1690,In_2067,In_990);
nor U1691 (N_1691,N_911,N_486);
nor U1692 (N_1692,N_178,N_707);
nand U1693 (N_1693,In_941,In_76);
and U1694 (N_1694,In_347,In_2553);
or U1695 (N_1695,N_1258,N_971);
nand U1696 (N_1696,N_992,In_163);
xnor U1697 (N_1697,N_926,In_874);
xor U1698 (N_1698,N_817,In_1423);
nand U1699 (N_1699,N_124,In_2590);
or U1700 (N_1700,N_798,N_827);
xor U1701 (N_1701,N_1491,N_1230);
nor U1702 (N_1702,In_363,In_920);
nor U1703 (N_1703,In_1126,N_896);
and U1704 (N_1704,In_646,N_1180);
nor U1705 (N_1705,In_2017,N_1312);
nand U1706 (N_1706,N_368,N_889);
xor U1707 (N_1707,N_1214,In_497);
and U1708 (N_1708,N_1299,In_2183);
or U1709 (N_1709,In_2399,N_437);
nand U1710 (N_1710,N_1382,N_800);
nand U1711 (N_1711,In_307,In_1977);
xnor U1712 (N_1712,N_236,N_157);
and U1713 (N_1713,N_516,N_1044);
nand U1714 (N_1714,N_1246,N_751);
and U1715 (N_1715,In_294,In_2703);
or U1716 (N_1716,In_2458,N_369);
or U1717 (N_1717,N_783,In_1765);
nor U1718 (N_1718,In_324,N_132);
or U1719 (N_1719,In_2993,In_1001);
or U1720 (N_1720,In_2464,In_2138);
or U1721 (N_1721,In_180,N_235);
nor U1722 (N_1722,N_1046,N_1244);
or U1723 (N_1723,N_1351,N_1089);
nand U1724 (N_1724,N_709,N_501);
or U1725 (N_1725,N_1122,N_1434);
or U1726 (N_1726,In_203,In_2268);
nor U1727 (N_1727,In_1805,N_870);
nand U1728 (N_1728,In_688,In_2659);
and U1729 (N_1729,N_1323,In_2328);
or U1730 (N_1730,In_516,N_852);
or U1731 (N_1731,In_1983,In_2731);
nor U1732 (N_1732,N_999,In_2741);
xor U1733 (N_1733,In_2056,In_1475);
nand U1734 (N_1734,In_1941,N_322);
nor U1735 (N_1735,N_1300,N_1331);
xnor U1736 (N_1736,N_1397,N_1361);
or U1737 (N_1737,In_636,N_402);
and U1738 (N_1738,N_1221,N_519);
nor U1739 (N_1739,N_489,In_578);
nand U1740 (N_1740,N_283,N_968);
xor U1741 (N_1741,In_2705,N_1008);
and U1742 (N_1742,In_362,N_1404);
and U1743 (N_1743,In_110,In_268);
and U1744 (N_1744,In_1953,N_1215);
xnor U1745 (N_1745,In_2204,N_953);
or U1746 (N_1746,N_512,N_303);
nand U1747 (N_1747,In_2222,N_1050);
or U1748 (N_1748,In_171,N_1317);
xnor U1749 (N_1749,N_1241,In_2672);
xor U1750 (N_1750,N_745,In_161);
nor U1751 (N_1751,In_24,N_921);
nand U1752 (N_1752,In_98,N_366);
and U1753 (N_1753,N_1255,N_925);
nand U1754 (N_1754,N_536,In_1665);
nand U1755 (N_1755,In_1460,In_1915);
xnor U1756 (N_1756,In_181,In_2934);
nand U1757 (N_1757,In_581,N_1359);
xnor U1758 (N_1758,N_981,In_1006);
nand U1759 (N_1759,N_58,In_2190);
nand U1760 (N_1760,N_1304,N_323);
nor U1761 (N_1761,N_965,In_2025);
nand U1762 (N_1762,N_656,N_652);
nor U1763 (N_1763,N_5,In_2986);
nand U1764 (N_1764,N_1140,In_2015);
or U1765 (N_1765,N_721,N_1366);
and U1766 (N_1766,In_2438,N_885);
xor U1767 (N_1767,In_1331,N_1287);
and U1768 (N_1768,N_1376,N_420);
xor U1769 (N_1769,N_785,N_1368);
nor U1770 (N_1770,N_1204,In_2372);
and U1771 (N_1771,N_12,In_1056);
nand U1772 (N_1772,N_1000,In_1234);
and U1773 (N_1773,In_1292,N_989);
and U1774 (N_1774,N_332,N_733);
nor U1775 (N_1775,N_936,In_1568);
or U1776 (N_1776,N_941,N_381);
or U1777 (N_1777,In_879,N_621);
and U1778 (N_1778,N_868,In_488);
nand U1779 (N_1779,N_608,In_2658);
nor U1780 (N_1780,In_2170,N_66);
nor U1781 (N_1781,In_97,N_1349);
or U1782 (N_1782,In_2972,N_1252);
and U1783 (N_1783,N_57,N_1355);
xor U1784 (N_1784,In_2630,In_1127);
xnor U1785 (N_1785,In_1268,In_2174);
nor U1786 (N_1786,In_2511,In_1161);
xor U1787 (N_1787,N_1273,In_1895);
nand U1788 (N_1788,In_1118,N_1305);
nand U1789 (N_1789,In_1598,N_1133);
xnor U1790 (N_1790,N_1109,N_958);
nand U1791 (N_1791,N_1459,N_1026);
or U1792 (N_1792,N_1395,In_2996);
nand U1793 (N_1793,N_865,In_523);
or U1794 (N_1794,N_700,In_2048);
and U1795 (N_1795,N_1213,In_2330);
nand U1796 (N_1796,N_1322,N_302);
nor U1797 (N_1797,In_2910,N_1232);
xnor U1798 (N_1798,In_1463,In_2872);
or U1799 (N_1799,In_2940,N_985);
xnor U1800 (N_1800,N_1703,N_1072);
nor U1801 (N_1801,N_839,N_1741);
nand U1802 (N_1802,N_599,N_1665);
and U1803 (N_1803,N_1519,N_1250);
or U1804 (N_1804,N_1760,N_1711);
nor U1805 (N_1805,In_2988,N_558);
or U1806 (N_1806,N_1117,In_1288);
nand U1807 (N_1807,N_1292,N_1516);
or U1808 (N_1808,N_1313,In_289);
or U1809 (N_1809,N_1015,In_179);
nor U1810 (N_1810,N_1306,N_1294);
xor U1811 (N_1811,N_919,N_1319);
nor U1812 (N_1812,In_2792,N_1378);
xor U1813 (N_1813,In_1955,N_1796);
and U1814 (N_1814,N_825,N_1579);
xor U1815 (N_1815,N_1403,N_1533);
nand U1816 (N_1816,In_887,In_2739);
nand U1817 (N_1817,N_977,In_1437);
and U1818 (N_1818,N_1377,In_257);
and U1819 (N_1819,N_1023,N_1783);
nand U1820 (N_1820,In_259,In_224);
nor U1821 (N_1821,N_1201,N_32);
xnor U1822 (N_1822,N_1353,In_2354);
nand U1823 (N_1823,In_2424,N_1222);
or U1824 (N_1824,N_1581,N_219);
or U1825 (N_1825,N_677,N_1688);
nor U1826 (N_1826,N_1540,N_931);
nor U1827 (N_1827,In_22,N_1792);
nand U1828 (N_1828,N_1593,In_1909);
nor U1829 (N_1829,N_1059,N_1216);
nor U1830 (N_1830,N_1768,In_1028);
or U1831 (N_1831,N_1607,N_471);
nor U1832 (N_1832,In_1726,N_1297);
and U1833 (N_1833,In_506,N_754);
or U1834 (N_1834,N_732,In_641);
and U1835 (N_1835,In_601,N_1398);
and U1836 (N_1836,In_3,N_543);
nor U1837 (N_1837,N_1526,N_916);
nor U1838 (N_1838,N_1573,N_1604);
nand U1839 (N_1839,N_1024,N_422);
and U1840 (N_1840,N_1691,In_381);
nand U1841 (N_1841,N_414,In_2442);
xnor U1842 (N_1842,In_1834,N_1652);
nor U1843 (N_1843,In_699,In_804);
xor U1844 (N_1844,N_1514,N_1348);
or U1845 (N_1845,N_1301,In_2333);
xnor U1846 (N_1846,In_626,In_848);
or U1847 (N_1847,In_1557,In_1054);
nand U1848 (N_1848,In_1362,N_1290);
nor U1849 (N_1849,In_474,N_1571);
nand U1850 (N_1850,In_2394,N_1448);
nand U1851 (N_1851,N_711,N_986);
and U1852 (N_1852,N_1228,N_1746);
or U1853 (N_1853,In_2191,N_1501);
xor U1854 (N_1854,In_1560,N_1654);
or U1855 (N_1855,In_2444,N_1350);
xnor U1856 (N_1856,N_467,N_1165);
and U1857 (N_1857,In_1871,N_1585);
xnor U1858 (N_1858,N_917,N_1527);
xor U1859 (N_1859,In_2577,N_542);
nor U1860 (N_1860,In_112,N_101);
nand U1861 (N_1861,N_1314,In_2147);
nor U1862 (N_1862,N_1586,In_801);
xor U1863 (N_1863,N_1620,N_493);
nor U1864 (N_1864,In_60,N_869);
nor U1865 (N_1865,N_1645,In_1003);
xor U1866 (N_1866,N_1343,In_582);
and U1867 (N_1867,N_581,In_913);
or U1868 (N_1868,N_851,N_1774);
nand U1869 (N_1869,N_1436,In_1401);
and U1870 (N_1870,In_1733,In_1208);
xor U1871 (N_1871,N_1280,In_1998);
nand U1872 (N_1872,N_1695,In_1392);
nor U1873 (N_1873,N_1114,N_25);
and U1874 (N_1874,N_1547,N_1663);
and U1875 (N_1875,In_385,N_1321);
and U1876 (N_1876,N_1200,N_1025);
or U1877 (N_1877,N_1326,N_142);
xnor U1878 (N_1878,N_1727,In_1030);
xor U1879 (N_1879,N_1623,N_1548);
or U1880 (N_1880,N_906,In_841);
and U1881 (N_1881,In_808,In_1324);
nor U1882 (N_1882,N_987,In_849);
and U1883 (N_1883,N_806,N_1502);
nor U1884 (N_1884,N_1649,N_1601);
xnor U1885 (N_1885,N_1484,In_783);
nand U1886 (N_1886,In_1839,N_1633);
and U1887 (N_1887,In_1120,N_1724);
xor U1888 (N_1888,In_2736,N_1309);
and U1889 (N_1889,N_1694,N_975);
nor U1890 (N_1890,In_2459,N_1558);
nor U1891 (N_1891,In_1049,In_612);
xor U1892 (N_1892,N_1627,N_1419);
xnor U1893 (N_1893,N_526,N_1506);
or U1894 (N_1894,N_1335,N_1460);
nor U1895 (N_1895,N_607,N_1794);
nor U1896 (N_1896,N_1451,In_1378);
or U1897 (N_1897,In_262,N_809);
nor U1898 (N_1898,N_1719,N_1755);
and U1899 (N_1899,N_477,N_1710);
xor U1900 (N_1900,N_1720,In_1062);
xor U1901 (N_1901,N_1583,N_1307);
nor U1902 (N_1902,N_1433,In_303);
or U1903 (N_1903,N_1017,In_2646);
and U1904 (N_1904,N_1054,N_1712);
or U1905 (N_1905,In_2782,In_2890);
nand U1906 (N_1906,N_1279,N_335);
and U1907 (N_1907,In_2044,N_1439);
xor U1908 (N_1908,In_1880,In_898);
nand U1909 (N_1909,N_1726,N_49);
nor U1910 (N_1910,N_1569,N_829);
or U1911 (N_1911,N_1327,N_1150);
or U1912 (N_1912,N_1572,In_2057);
xnor U1913 (N_1913,N_1525,N_245);
nand U1914 (N_1914,N_1418,In_2192);
xor U1915 (N_1915,N_1701,N_1560);
and U1916 (N_1916,N_1638,In_2039);
or U1917 (N_1917,N_504,N_834);
nor U1918 (N_1918,N_1566,N_1416);
xnor U1919 (N_1919,In_208,N_909);
and U1920 (N_1920,N_1148,N_1218);
nand U1921 (N_1921,N_284,N_187);
nand U1922 (N_1922,In_1058,N_1757);
and U1923 (N_1923,In_207,N_640);
nand U1924 (N_1924,In_980,N_19);
or U1925 (N_1925,In_154,In_0);
and U1926 (N_1926,In_1512,In_15);
nand U1927 (N_1927,N_1352,In_2991);
xor U1928 (N_1928,N_448,In_151);
and U1929 (N_1929,In_2274,In_1090);
and U1930 (N_1930,N_499,N_1452);
and U1931 (N_1931,N_1066,N_297);
and U1932 (N_1932,In_2450,N_1609);
nor U1933 (N_1933,N_1302,N_897);
nand U1934 (N_1934,In_2930,In_2955);
xnor U1935 (N_1935,In_2053,N_1131);
nand U1936 (N_1936,N_1596,In_1831);
and U1937 (N_1937,N_1243,In_408);
xnor U1938 (N_1938,N_1308,N_37);
xor U1939 (N_1939,N_1636,N_530);
nand U1940 (N_1940,In_2142,N_1704);
and U1941 (N_1941,In_1848,N_1677);
and U1942 (N_1942,N_482,In_1569);
nor U1943 (N_1943,In_2302,In_88);
or U1944 (N_1944,N_735,In_1981);
or U1945 (N_1945,In_2341,In_527);
and U1946 (N_1946,N_1440,N_833);
nand U1947 (N_1947,N_1354,N_1751);
or U1948 (N_1948,N_1659,N_1386);
nand U1949 (N_1949,In_2076,N_883);
nand U1950 (N_1950,N_1728,N_946);
nor U1951 (N_1951,In_189,In_639);
nand U1952 (N_1952,In_2860,N_736);
nand U1953 (N_1953,N_848,N_1430);
nor U1954 (N_1954,N_625,N_94);
nand U1955 (N_1955,N_1197,N_1731);
xor U1956 (N_1956,In_2402,In_1313);
or U1957 (N_1957,In_2499,N_1582);
or U1958 (N_1958,N_1578,In_2574);
nor U1959 (N_1959,N_1169,In_2270);
nor U1960 (N_1960,In_1574,In_1239);
or U1961 (N_1961,N_1687,N_1595);
xnor U1962 (N_1962,In_752,N_1789);
nor U1963 (N_1963,N_669,N_758);
nand U1964 (N_1964,N_1646,N_1067);
nor U1965 (N_1965,In_1939,N_778);
or U1966 (N_1966,In_2824,In_2177);
nand U1967 (N_1967,In_176,N_1630);
or U1968 (N_1968,N_1543,N_1598);
nand U1969 (N_1969,N_1678,In_1774);
xor U1970 (N_1970,N_1186,N_1342);
nor U1971 (N_1971,N_1576,In_642);
nor U1972 (N_1972,In_1674,N_1328);
and U1973 (N_1973,N_1428,N_1562);
nor U1974 (N_1974,N_1610,N_1524);
nand U1975 (N_1975,In_452,N_364);
nand U1976 (N_1976,N_1425,In_2606);
xor U1977 (N_1977,N_1372,N_1570);
nand U1978 (N_1978,N_1644,N_970);
or U1979 (N_1979,N_1247,In_2466);
xnor U1980 (N_1980,N_1777,N_1231);
or U1981 (N_1981,N_823,N_1708);
nand U1982 (N_1982,N_1396,N_1742);
nand U1983 (N_1983,N_1286,N_1639);
and U1984 (N_1984,N_1698,N_382);
nor U1985 (N_1985,N_1647,In_1231);
and U1986 (N_1986,N_1565,In_2474);
xor U1987 (N_1987,N_744,In_953);
nor U1988 (N_1988,N_141,N_1643);
or U1989 (N_1989,N_1671,In_2096);
nor U1990 (N_1990,N_1454,N_997);
xnor U1991 (N_1991,In_2760,N_1748);
or U1992 (N_1992,N_983,In_2720);
and U1993 (N_1993,N_775,N_1507);
xor U1994 (N_1994,In_1739,N_206);
xnor U1995 (N_1995,N_650,N_1656);
xor U1996 (N_1996,N_1202,N_1371);
nor U1997 (N_1997,N_1224,N_1123);
and U1998 (N_1998,N_1166,In_827);
nand U1999 (N_1999,N_1414,N_1784);
nand U2000 (N_2000,In_431,N_1512);
nor U2001 (N_2001,N_1763,N_616);
or U2002 (N_2002,N_1513,N_1778);
and U2003 (N_2003,N_405,N_788);
nand U2004 (N_2004,N_1094,N_545);
or U2005 (N_2005,N_1511,In_1297);
or U2006 (N_2006,In_71,In_177);
and U2007 (N_2007,N_553,In_2995);
xnor U2008 (N_2008,N_1116,N_1036);
or U2009 (N_2009,N_1471,In_267);
and U2010 (N_2010,In_2029,N_1618);
or U2011 (N_2011,N_1693,N_990);
nand U2012 (N_2012,N_1174,N_876);
and U2013 (N_2013,In_765,N_1155);
and U2014 (N_2014,N_1391,N_1457);
nand U2015 (N_2015,N_1217,N_1736);
or U2016 (N_2016,N_1669,N_1456);
or U2017 (N_2017,N_502,N_548);
xnor U2018 (N_2018,In_1973,In_2613);
xnor U2019 (N_2019,N_1284,N_1650);
xnor U2020 (N_2020,In_1944,N_1684);
and U2021 (N_2021,In_344,N_774);
nor U2022 (N_2022,N_1020,In_1801);
xor U2023 (N_2023,N_1492,N_1614);
nand U2024 (N_2024,N_1537,In_1551);
nor U2025 (N_2025,N_1510,In_1342);
or U2026 (N_2026,N_615,In_916);
xor U2027 (N_2027,N_1564,In_1879);
xor U2028 (N_2028,In_1802,N_769);
nor U2029 (N_2029,In_643,N_1660);
xor U2030 (N_2030,N_1681,N_1690);
nand U2031 (N_2031,N_1466,In_490);
or U2032 (N_2032,In_367,N_1594);
or U2033 (N_2033,N_1503,In_314);
nand U2034 (N_2034,N_1550,N_1181);
xor U2035 (N_2035,N_648,N_456);
and U2036 (N_2036,N_1463,N_808);
and U2037 (N_2037,N_1257,N_1555);
nand U2038 (N_2038,N_1670,In_2769);
and U2039 (N_2039,N_1631,N_1167);
xnor U2040 (N_2040,N_1615,N_1138);
and U2041 (N_2041,In_2014,N_1124);
nand U2042 (N_2042,In_503,In_2899);
or U2043 (N_2043,N_1541,N_915);
or U2044 (N_2044,In_1142,N_1745);
nand U2045 (N_2045,N_932,N_1655);
nand U2046 (N_2046,In_494,N_1367);
nor U2047 (N_2047,N_1520,In_2159);
or U2048 (N_2048,N_354,N_1651);
or U2049 (N_2049,N_1281,N_1674);
or U2050 (N_2050,In_440,N_497);
nand U2051 (N_2051,N_1697,N_1790);
or U2052 (N_2052,N_1600,N_1743);
nand U2053 (N_2053,In_274,N_562);
nand U2054 (N_2054,N_319,In_2563);
and U2055 (N_2055,N_940,In_428);
and U2056 (N_2056,In_2633,N_256);
or U2057 (N_2057,In_486,In_2202);
nand U2058 (N_2058,N_687,N_1339);
or U2059 (N_2059,In_1365,In_83);
nand U2060 (N_2060,In_2922,N_1182);
and U2061 (N_2061,In_926,In_2729);
nor U2062 (N_2062,N_1642,In_2040);
xor U2063 (N_2063,In_173,N_1523);
nand U2064 (N_2064,N_1427,In_400);
nor U2065 (N_2065,N_1409,In_2060);
nor U2066 (N_2066,N_0,N_1384);
nor U2067 (N_2067,In_2797,N_643);
and U2068 (N_2068,In_417,In_326);
nand U2069 (N_2069,N_1658,N_1488);
nand U2070 (N_2070,N_1556,N_966);
or U2071 (N_2071,In_2228,N_1325);
and U2072 (N_2072,N_64,In_358);
or U2073 (N_2073,In_2062,N_1584);
nor U2074 (N_2074,N_1429,N_1529);
xor U2075 (N_2075,N_1019,N_1269);
xor U2076 (N_2076,In_943,In_2628);
or U2077 (N_2077,In_445,N_884);
nor U2078 (N_2078,In_505,N_1675);
nor U2079 (N_2079,N_1563,In_2352);
or U2080 (N_2080,N_1739,N_1191);
nor U2081 (N_2081,N_1621,In_1745);
or U2082 (N_2082,In_457,N_1344);
or U2083 (N_2083,N_457,N_1262);
and U2084 (N_2084,N_1130,N_1261);
xnor U2085 (N_2085,N_1193,N_1740);
nor U2086 (N_2086,N_317,N_1441);
nand U2087 (N_2087,N_1229,N_1341);
or U2088 (N_2088,N_1753,N_1756);
xor U2089 (N_2089,N_1761,N_1759);
nand U2090 (N_2090,N_1518,In_1229);
nand U2091 (N_2091,In_2674,N_1276);
and U2092 (N_2092,N_1086,N_78);
nand U2093 (N_2093,N_232,N_1496);
or U2094 (N_2094,N_604,N_1245);
nor U2095 (N_2095,In_871,N_1539);
xnor U2096 (N_2096,N_1356,In_1055);
or U2097 (N_2097,N_1733,N_1773);
nor U2098 (N_2098,N_1587,N_1725);
or U2099 (N_2099,In_2642,N_1549);
nor U2100 (N_2100,N_2076,N_106);
nand U2101 (N_2101,N_1406,N_2031);
or U2102 (N_2102,N_1163,N_1979);
xnor U2103 (N_2103,In_2965,N_801);
xnor U2104 (N_2104,In_2704,N_1239);
nor U2105 (N_2105,N_1863,N_54);
and U2106 (N_2106,In_634,N_912);
xor U2107 (N_2107,N_2022,N_1476);
xnor U2108 (N_2108,N_2083,N_1068);
nand U2109 (N_2109,N_1867,N_690);
nor U2110 (N_2110,N_1847,N_1453);
nor U2111 (N_2111,N_1001,In_1205);
nand U2112 (N_2112,In_1721,N_1968);
or U2113 (N_2113,In_2269,In_33);
or U2114 (N_2114,N_2012,N_1683);
and U2115 (N_2115,N_1871,N_1468);
or U2116 (N_2116,N_1424,N_2052);
or U2117 (N_2117,N_1912,N_2020);
and U2118 (N_2118,In_1227,In_914);
xor U2119 (N_2119,N_1504,In_2240);
or U2120 (N_2120,N_988,N_1826);
nand U2121 (N_2121,N_2023,In_1082);
nand U2122 (N_2122,N_2080,N_1919);
nand U2123 (N_2123,N_1664,N_1295);
and U2124 (N_2124,In_2854,In_2884);
nor U2125 (N_2125,In_2597,In_2655);
nand U2126 (N_2126,In_1669,N_1938);
nor U2127 (N_2127,In_1133,N_1225);
and U2128 (N_2128,N_1128,N_836);
and U2129 (N_2129,N_1461,N_1988);
xnor U2130 (N_2130,N_686,In_904);
nor U2131 (N_2131,N_1483,N_1521);
nand U2132 (N_2132,N_1103,N_1957);
nand U2133 (N_2133,In_1542,N_995);
or U2134 (N_2134,N_1945,N_1747);
nand U2135 (N_2135,N_1839,N_2038);
xnor U2136 (N_2136,N_1946,N_1921);
or U2137 (N_2137,In_1132,N_1991);
nand U2138 (N_2138,In_2853,N_2099);
nor U2139 (N_2139,N_1929,N_1254);
nand U2140 (N_2140,In_186,N_388);
and U2141 (N_2141,N_1141,N_1953);
nor U2142 (N_2142,N_1821,N_1667);
nand U2143 (N_2143,N_2062,N_1553);
or U2144 (N_2144,N_1490,N_1884);
or U2145 (N_2145,N_2036,N_1364);
nor U2146 (N_2146,N_1986,N_1412);
nand U2147 (N_2147,N_1392,N_1718);
xnor U2148 (N_2148,N_969,N_738);
nand U2149 (N_2149,N_1707,In_2487);
and U2150 (N_2150,N_1509,In_1020);
nor U2151 (N_2151,N_1880,N_692);
or U2152 (N_2152,N_1477,N_1387);
xor U2153 (N_2153,N_439,N_2018);
nor U2154 (N_2154,N_1956,N_1505);
and U2155 (N_2155,N_1161,In_1174);
xor U2156 (N_2156,N_1845,N_244);
and U2157 (N_2157,N_2030,N_1907);
xnor U2158 (N_2158,N_352,In_252);
xnor U2159 (N_2159,N_1085,In_828);
and U2160 (N_2160,N_1270,N_1978);
nand U2161 (N_2161,N_1672,N_2009);
and U2162 (N_2162,N_90,N_1850);
xor U2163 (N_2163,N_1653,N_2071);
and U2164 (N_2164,In_354,N_1916);
nand U2165 (N_2165,N_639,N_2007);
nand U2166 (N_2166,N_1223,N_1925);
xnor U2167 (N_2167,N_1987,In_222);
and U2168 (N_2168,N_2058,N_1823);
nor U2169 (N_2169,N_1854,In_1394);
nor U2170 (N_2170,N_1960,N_950);
nor U2171 (N_2171,N_1469,In_787);
or U2172 (N_2172,N_1554,N_2094);
nor U2173 (N_2173,N_1063,N_191);
or U2174 (N_2174,In_2398,In_2690);
nor U2175 (N_2175,N_1752,In_1804);
and U2176 (N_2176,N_1447,N_1899);
or U2177 (N_2177,N_2079,N_1611);
or U2178 (N_2178,N_1498,N_1283);
nor U2179 (N_2179,N_586,N_1983);
xnor U2180 (N_2180,N_1714,N_1861);
nor U2181 (N_2181,N_1668,N_1932);
and U2182 (N_2182,In_1043,In_541);
or U2183 (N_2183,N_1835,N_879);
xnor U2184 (N_2184,N_1027,In_2677);
and U2185 (N_2185,N_1951,N_2002);
xnor U2186 (N_2186,N_1862,In_2059);
xor U2187 (N_2187,N_1119,N_1890);
and U2188 (N_2188,N_724,N_2078);
nor U2189 (N_2189,N_2053,N_1819);
nor U2190 (N_2190,N_1970,N_880);
and U2191 (N_2191,In_2388,N_2000);
or U2192 (N_2192,N_838,N_1347);
or U2193 (N_2193,N_1475,N_1029);
and U2194 (N_2194,In_1637,N_1923);
nor U2195 (N_2195,In_1643,N_1775);
xor U2196 (N_2196,In_815,N_1947);
xnor U2197 (N_2197,N_1735,In_1746);
and U2198 (N_2198,N_1470,N_1914);
nor U2199 (N_2199,N_1804,N_1039);
xnor U2200 (N_2200,In_1756,N_1832);
nand U2201 (N_2201,N_1767,N_1765);
xnor U2202 (N_2202,N_1272,N_2067);
nand U2203 (N_2203,In_1875,N_1606);
and U2204 (N_2204,N_1338,N_1786);
xnor U2205 (N_2205,N_2075,N_1853);
nor U2206 (N_2206,N_1958,N_1552);
xor U2207 (N_2207,In_1360,N_1769);
nand U2208 (N_2208,N_2034,In_2396);
xnor U2209 (N_2209,In_2241,N_1467);
xor U2210 (N_2210,N_1941,In_1453);
xor U2211 (N_2211,N_1546,N_30);
and U2212 (N_2212,N_1405,N_346);
or U2213 (N_2213,N_1426,N_1210);
and U2214 (N_2214,N_2088,N_1984);
or U2215 (N_2215,In_103,N_1887);
or U2216 (N_2216,N_1028,N_254);
xnor U2217 (N_2217,N_1226,N_1934);
or U2218 (N_2218,N_1087,In_2335);
and U2219 (N_2219,N_374,In_1571);
xor U2220 (N_2220,N_1715,N_1413);
nand U2221 (N_2221,N_1106,N_1237);
nor U2222 (N_2222,N_1389,N_1825);
nand U2223 (N_2223,N_1629,N_1865);
nor U2224 (N_2224,In_1517,N_1795);
and U2225 (N_2225,N_1965,N_1324);
nor U2226 (N_2226,In_1914,N_1220);
nand U2227 (N_2227,In_198,N_1886);
or U2228 (N_2228,N_1227,N_2066);
nand U2229 (N_2229,N_1770,N_1906);
and U2230 (N_2230,N_2017,N_1877);
and U2231 (N_2231,In_1240,N_1021);
and U2232 (N_2232,N_274,In_1325);
or U2233 (N_2233,N_1974,In_1481);
or U2234 (N_2234,In_2021,In_204);
and U2235 (N_2235,N_1900,N_524);
nand U2236 (N_2236,N_1771,N_2039);
nor U2237 (N_2237,In_376,N_1859);
or U2238 (N_2238,N_609,N_715);
or U2239 (N_2239,N_1776,N_1635);
or U2240 (N_2240,N_664,N_1869);
or U2241 (N_2241,N_1840,N_1781);
nand U2242 (N_2242,N_1993,N_1431);
nand U2243 (N_2243,N_1897,In_949);
and U2244 (N_2244,N_913,N_1336);
nand U2245 (N_2245,In_1355,N_1966);
nand U2246 (N_2246,N_1494,N_1073);
xor U2247 (N_2247,In_2186,N_1700);
nor U2248 (N_2248,N_1913,N_1632);
nor U2249 (N_2249,N_1076,N_417);
or U2250 (N_2250,N_1896,N_2050);
and U2251 (N_2251,N_618,N_1822);
nand U2252 (N_2252,N_2097,N_710);
nor U2253 (N_2253,N_1816,N_2005);
xor U2254 (N_2254,N_1891,N_1545);
and U2255 (N_2255,N_937,N_2001);
nor U2256 (N_2256,In_165,N_1031);
nor U2257 (N_2257,N_2045,N_1531);
xnor U2258 (N_2258,N_1612,N_2046);
or U2259 (N_2259,N_1948,In_1710);
nand U2260 (N_2260,N_1303,In_479);
nor U2261 (N_2261,N_1240,N_159);
or U2262 (N_2262,N_1190,N_1881);
nor U2263 (N_2263,N_1806,N_1278);
and U2264 (N_2264,In_905,N_16);
or U2265 (N_2265,N_1723,N_544);
and U2266 (N_2266,N_1375,N_1937);
and U2267 (N_2267,N_1721,In_1575);
xor U2268 (N_2268,In_1248,N_1943);
and U2269 (N_2269,N_1259,N_1959);
nand U2270 (N_2270,N_1811,N_1575);
xor U2271 (N_2271,N_2095,N_36);
or U2272 (N_2272,N_1738,N_1857);
or U2273 (N_2273,In_1039,N_1274);
nor U2274 (N_2274,In_2454,N_1446);
xnor U2275 (N_2275,N_85,N_1055);
nor U2276 (N_2276,N_1812,In_2136);
nand U2277 (N_2277,In_796,N_1904);
and U2278 (N_2278,In_1607,N_1911);
nand U2279 (N_2279,N_959,N_1903);
nor U2280 (N_2280,N_1472,In_402);
and U2281 (N_2281,N_1268,In_1448);
xnor U2282 (N_2282,N_858,In_2840);
nand U2283 (N_2283,N_1820,N_2091);
or U2284 (N_2284,N_1995,N_1580);
and U2285 (N_2285,N_1333,N_1515);
or U2286 (N_2286,N_1942,In_2207);
nor U2287 (N_2287,In_2432,N_2026);
xnor U2288 (N_2288,N_1915,N_1212);
or U2289 (N_2289,N_2028,In_2722);
or U2290 (N_2290,In_1228,N_617);
and U2291 (N_2291,N_1603,In_1683);
xor U2292 (N_2292,In_2033,N_570);
nor U2293 (N_2293,N_1597,N_1954);
xor U2294 (N_2294,In_1742,N_1442);
nand U2295 (N_2295,N_1605,N_1872);
xor U2296 (N_2296,N_1624,N_1814);
or U2297 (N_2297,In_1081,N_2060);
nor U2298 (N_2298,N_1878,In_2280);
or U2299 (N_2299,N_993,N_84);
nand U2300 (N_2300,N_1856,N_1699);
or U2301 (N_2301,N_591,N_2065);
xnor U2302 (N_2302,N_1935,N_1590);
and U2303 (N_2303,N_1933,In_2336);
or U2304 (N_2304,N_513,N_1551);
xnor U2305 (N_2305,N_1011,N_1895);
or U2306 (N_2306,N_1696,In_4);
xnor U2307 (N_2307,In_1945,N_1885);
nand U2308 (N_2308,N_1033,N_1267);
and U2309 (N_2309,N_1990,N_2092);
and U2310 (N_2310,In_2921,N_1964);
nor U2311 (N_2311,In_1877,N_1831);
xnor U2312 (N_2312,N_1855,N_2090);
or U2313 (N_2313,N_904,N_1559);
and U2314 (N_2314,In_298,N_1357);
nand U2315 (N_2315,N_2010,N_1369);
xnor U2316 (N_2316,N_1749,N_2096);
or U2317 (N_2317,In_673,N_1289);
or U2318 (N_2318,N_1713,In_1526);
nor U2319 (N_2319,In_2896,N_1841);
xnor U2320 (N_2320,In_854,N_1532);
xor U2321 (N_2321,N_2074,N_569);
xnor U2322 (N_2322,N_173,In_686);
nand U2323 (N_2323,N_2084,N_1393);
and U2324 (N_2324,N_1961,N_1249);
xnor U2325 (N_2325,N_1385,In_945);
or U2326 (N_2326,In_291,In_1612);
or U2327 (N_2327,In_2498,N_1499);
nor U2328 (N_2328,N_1474,In_491);
or U2329 (N_2329,N_1894,N_2025);
nand U2330 (N_2330,N_1373,N_982);
or U2331 (N_2331,In_218,N_713);
nor U2332 (N_2332,N_826,N_1219);
and U2333 (N_2333,N_1592,N_1994);
and U2334 (N_2334,N_1764,N_409);
and U2335 (N_2335,N_1730,N_1567);
nand U2336 (N_2336,N_1808,N_1917);
and U2337 (N_2337,In_2564,N_2003);
xnor U2338 (N_2338,N_1892,In_1329);
nor U2339 (N_2339,N_1996,N_1800);
nand U2340 (N_2340,N_1061,N_1577);
and U2341 (N_2341,N_1081,N_899);
or U2342 (N_2342,In_1198,N_174);
and U2343 (N_2343,In_194,N_2048);
nor U2344 (N_2344,N_1608,N_1105);
or U2345 (N_2345,N_1172,N_1801);
nor U2346 (N_2346,In_2847,In_1541);
or U2347 (N_2347,N_266,In_1359);
nor U2348 (N_2348,N_1905,N_2011);
or U2349 (N_2349,N_2059,N_363);
or U2350 (N_2350,N_2073,N_2057);
nor U2351 (N_2351,N_2014,N_1702);
nor U2352 (N_2352,N_1949,N_1234);
nand U2353 (N_2353,N_1963,N_2093);
or U2354 (N_2354,N_2077,N_1864);
and U2355 (N_2355,N_1999,N_96);
xnor U2356 (N_2356,N_1838,N_1879);
or U2357 (N_2357,N_2029,N_1902);
or U2358 (N_2358,In_14,In_1353);
or U2359 (N_2359,In_1412,In_2281);
and U2360 (N_2360,N_1717,N_1500);
nand U2361 (N_2361,In_2627,In_1144);
nand U2362 (N_2362,N_2087,N_1682);
xor U2363 (N_2363,N_1709,N_1534);
nor U2364 (N_2364,N_1744,N_2019);
nand U2365 (N_2365,In_2550,N_1830);
nor U2366 (N_2366,N_1910,N_672);
or U2367 (N_2367,In_219,N_1936);
and U2368 (N_2368,N_1798,N_2037);
nand U2369 (N_2369,N_242,N_1976);
or U2370 (N_2370,N_1992,In_436);
xor U2371 (N_2371,N_539,In_2298);
and U2372 (N_2372,In_1384,N_264);
or U2373 (N_2373,N_2044,N_1782);
nor U2374 (N_2374,N_1722,N_1432);
or U2375 (N_2375,N_1588,N_730);
xor U2376 (N_2376,N_1927,N_1661);
xnor U2377 (N_2377,N_1037,N_1918);
xnor U2378 (N_2378,N_1849,N_1686);
and U2379 (N_2379,N_1544,N_1486);
xnor U2380 (N_2380,N_1766,N_1557);
xnor U2381 (N_2381,N_1685,In_2439);
nor U2382 (N_2382,In_2203,In_991);
or U2383 (N_2383,N_1093,N_1591);
nand U2384 (N_2384,In_2362,N_2021);
or U2385 (N_2385,N_1846,N_1619);
xor U2386 (N_2386,N_161,N_491);
xor U2387 (N_2387,N_2056,N_1788);
nand U2388 (N_2388,N_397,N_2015);
and U2389 (N_2389,N_1772,N_1673);
or U2390 (N_2390,N_1177,N_1680);
nand U2391 (N_2391,N_1358,N_355);
nand U2392 (N_2392,N_1101,N_1833);
and U2393 (N_2393,N_2063,N_602);
nand U2394 (N_2394,In_782,N_1950);
xor U2395 (N_2395,N_2004,In_1115);
or U2396 (N_2396,N_1329,In_2963);
nor U2397 (N_2397,In_973,In_706);
and U2398 (N_2398,N_2042,N_1873);
xnor U2399 (N_2399,N_1842,In_1037);
and U2400 (N_2400,N_2142,N_1985);
xor U2401 (N_2401,In_2775,In_2702);
nand U2402 (N_2402,N_1866,N_2197);
nand U2403 (N_2403,N_1977,N_1628);
nor U2404 (N_2404,N_2324,N_1944);
and U2405 (N_2405,N_2301,N_2296);
nand U2406 (N_2406,N_1641,N_1858);
nor U2407 (N_2407,N_2362,In_1931);
xor U2408 (N_2408,N_2204,N_1803);
nand U2409 (N_2409,N_1253,N_379);
and U2410 (N_2410,N_2192,N_2232);
and U2411 (N_2411,N_706,N_2013);
or U2412 (N_2412,N_1370,N_1692);
and U2413 (N_2413,In_1744,N_2363);
or U2414 (N_2414,N_1829,N_385);
nand U2415 (N_2415,N_1802,N_2309);
nand U2416 (N_2416,N_1617,N_2255);
and U2417 (N_2417,N_1634,N_2006);
or U2418 (N_2418,N_2398,N_1981);
and U2419 (N_2419,N_2122,N_2143);
nand U2420 (N_2420,N_934,N_2310);
nand U2421 (N_2421,N_1288,N_2323);
xnor U2422 (N_2422,N_1530,N_2229);
nand U2423 (N_2423,N_923,N_2375);
nor U2424 (N_2424,N_1648,N_1330);
nor U2425 (N_2425,N_2394,N_2106);
nand U2426 (N_2426,N_2384,In_2214);
nand U2427 (N_2427,In_729,N_2275);
nor U2428 (N_2428,N_2115,N_2109);
and U2429 (N_2429,N_2245,N_2315);
or U2430 (N_2430,N_1616,N_2266);
and U2431 (N_2431,In_919,N_2348);
nand U2432 (N_2432,N_1034,N_1924);
nor U2433 (N_2433,N_1209,N_1729);
or U2434 (N_2434,N_2209,N_1889);
nor U2435 (N_2435,In_1992,N_2070);
and U2436 (N_2436,N_2198,N_2200);
nand U2437 (N_2437,N_1207,N_2327);
or U2438 (N_2438,N_2306,N_1455);
xnor U2439 (N_2439,N_2027,N_663);
xnor U2440 (N_2440,In_2409,N_2370);
nor U2441 (N_2441,N_2203,N_1750);
xnor U2442 (N_2442,N_2341,N_2082);
or U2443 (N_2443,N_1360,In_329);
nor U2444 (N_2444,N_2215,N_1975);
nand U2445 (N_2445,N_2043,N_2141);
nand U2446 (N_2446,N_2239,N_1928);
or U2447 (N_2447,N_428,In_843);
and U2448 (N_2448,N_2267,N_2113);
nand U2449 (N_2449,N_2161,N_2118);
nor U2450 (N_2450,N_2168,N_1982);
nand U2451 (N_2451,N_308,N_2347);
xor U2452 (N_2452,N_2146,N_1705);
or U2453 (N_2453,N_2123,N_2366);
nand U2454 (N_2454,N_1263,N_262);
nor U2455 (N_2455,N_2369,N_1282);
nor U2456 (N_2456,N_2243,N_2008);
nor U2457 (N_2457,N_1561,N_1908);
and U2458 (N_2458,N_1868,N_2265);
xor U2459 (N_2459,N_2317,N_2322);
nor U2460 (N_2460,N_2179,N_2041);
nand U2461 (N_2461,N_2228,N_637);
and U2462 (N_2462,In_2365,N_2376);
or U2463 (N_2463,N_2247,N_2374);
nor U2464 (N_2464,N_1415,N_2140);
and U2465 (N_2465,N_1939,N_1997);
nand U2466 (N_2466,N_2292,N_2325);
or U2467 (N_2467,N_2175,N_1016);
nand U2468 (N_2468,N_2253,N_1920);
xnor U2469 (N_2469,N_1791,N_1931);
nand U2470 (N_2470,N_2389,N_1809);
and U2471 (N_2471,N_2205,N_2136);
nand U2472 (N_2472,N_1799,N_1422);
xor U2473 (N_2473,N_2358,In_1172);
nor U2474 (N_2474,In_1960,N_282);
or U2475 (N_2475,N_2206,In_2119);
nand U2476 (N_2476,N_1508,N_1337);
nor U2477 (N_2477,N_1818,N_1882);
xnor U2478 (N_2478,In_2184,N_1383);
nor U2479 (N_2479,N_2246,N_133);
and U2480 (N_2480,N_1844,N_2276);
xor U2481 (N_2481,N_2211,N_2284);
xor U2482 (N_2482,N_905,N_2178);
and U2483 (N_2483,N_361,N_2193);
or U2484 (N_2484,N_2166,N_2258);
or U2485 (N_2485,N_2033,N_2278);
or U2486 (N_2486,N_2240,N_2261);
and U2487 (N_2487,N_2051,N_2280);
or U2488 (N_2488,N_2157,N_2064);
xnor U2489 (N_2489,N_2349,N_1909);
nor U2490 (N_2490,N_2264,In_2735);
or U2491 (N_2491,N_2298,N_143);
nor U2492 (N_2492,N_2170,N_1926);
or U2493 (N_2493,N_2314,N_2125);
or U2494 (N_2494,N_2299,N_2367);
and U2495 (N_2495,N_854,N_2241);
nor U2496 (N_2496,N_1517,N_2069);
nor U2497 (N_2497,N_1813,N_2167);
nand U2498 (N_2498,N_2355,N_2195);
xnor U2499 (N_2499,N_1851,N_2293);
nor U2500 (N_2500,N_2257,N_2368);
nand U2501 (N_2501,N_2225,N_1955);
and U2502 (N_2502,N_2199,N_2254);
xor U2503 (N_2503,In_6,N_1622);
xor U2504 (N_2504,N_1810,N_2102);
nor U2505 (N_2505,N_2328,N_2387);
xnor U2506 (N_2506,N_2286,N_2272);
nand U2507 (N_2507,N_1176,N_2343);
nand U2508 (N_2508,N_2182,N_2357);
and U2509 (N_2509,N_1901,N_2233);
nor U2510 (N_2510,N_1805,N_2016);
and U2511 (N_2511,N_2227,N_2236);
xnor U2512 (N_2512,N_1843,In_2547);
xor U2513 (N_2513,N_2068,N_120);
nor U2514 (N_2514,N_2149,N_1852);
xor U2515 (N_2515,N_2373,N_930);
or U2516 (N_2516,N_2133,N_1679);
nor U2517 (N_2517,N_2270,N_1568);
nor U2518 (N_2518,N_2103,N_2271);
nand U2519 (N_2519,N_1497,N_2399);
nand U2520 (N_2520,N_2072,In_2073);
nor U2521 (N_2521,N_2259,N_2216);
xor U2522 (N_2522,N_1666,N_1390);
xnor U2523 (N_2523,N_2107,N_2235);
nand U2524 (N_2524,N_2263,In_994);
xor U2525 (N_2525,N_2121,N_1438);
xor U2526 (N_2526,N_2165,In_205);
or U2527 (N_2527,In_1254,N_1980);
and U2528 (N_2528,N_2162,N_2285);
nor U2529 (N_2529,N_1785,N_2226);
nand U2530 (N_2530,N_1737,N_1827);
and U2531 (N_2531,N_2219,N_2282);
nand U2532 (N_2532,N_2155,In_558);
nor U2533 (N_2533,N_1883,N_2279);
nor U2534 (N_2534,In_2848,N_2174);
nor U2535 (N_2535,N_1407,N_2196);
xnor U2536 (N_2536,In_1913,N_2184);
nand U2537 (N_2537,N_1940,N_2316);
nand U2538 (N_2538,In_1959,In_1611);
and U2539 (N_2539,N_2352,N_2382);
and U2540 (N_2540,N_2105,N_2152);
xor U2541 (N_2541,N_2134,N_2111);
nand U2542 (N_2542,N_1898,N_578);
nand U2543 (N_2543,N_1420,N_2130);
nor U2544 (N_2544,N_1971,N_537);
nor U2545 (N_2545,In_206,N_2128);
or U2546 (N_2546,N_2365,N_2331);
nand U2547 (N_2547,In_2951,N_2221);
nor U2548 (N_2548,N_2172,N_2371);
nand U2549 (N_2549,N_1536,N_2342);
or U2550 (N_2550,N_2303,In_947);
nand U2551 (N_2551,N_890,N_2386);
nand U2552 (N_2552,N_2378,N_2148);
xnor U2553 (N_2553,N_2248,N_137);
nand U2554 (N_2554,N_2260,N_2144);
and U2555 (N_2555,N_2188,N_2024);
nand U2556 (N_2556,N_2202,N_2220);
or U2557 (N_2557,N_2132,N_2159);
nand U2558 (N_2558,In_1696,N_2190);
nor U2559 (N_2559,N_1888,N_1706);
and U2560 (N_2560,N_1107,N_1637);
nor U2561 (N_2561,In_1884,N_2308);
and U2562 (N_2562,N_1807,N_1538);
xnor U2563 (N_2563,N_2290,N_327);
nand U2564 (N_2564,N_2163,N_2339);
and U2565 (N_2565,N_2390,N_2124);
xnor U2566 (N_2566,N_2112,N_1754);
and U2567 (N_2567,N_1998,N_2249);
or U2568 (N_2568,N_1316,N_2114);
xor U2569 (N_2569,N_2153,N_1298);
nor U2570 (N_2570,N_2185,N_1836);
xor U2571 (N_2571,N_1930,N_2218);
nand U2572 (N_2572,N_2250,N_2150);
nand U2573 (N_2573,In_2380,N_2381);
nand U2574 (N_2574,N_2337,In_2532);
or U2575 (N_2575,In_1990,N_2291);
nand U2576 (N_2576,N_2158,N_2098);
nand U2577 (N_2577,N_1542,N_1205);
nor U2578 (N_2578,In_1752,N_1824);
or U2579 (N_2579,N_2126,N_1657);
or U2580 (N_2580,N_2283,N_2393);
and U2581 (N_2581,N_2164,N_635);
and U2582 (N_2582,N_2201,N_2305);
and U2583 (N_2583,N_2,N_1797);
nor U2584 (N_2584,N_158,In_1245);
nor U2585 (N_2585,N_1973,N_2268);
nand U2586 (N_2586,N_612,N_2212);
nor U2587 (N_2587,N_1817,N_2117);
xor U2588 (N_2588,N_2289,In_1097);
nor U2589 (N_2589,N_2085,N_2234);
nor U2590 (N_2590,N_2345,N_2252);
or U2591 (N_2591,N_964,N_211);
nand U2592 (N_2592,In_1866,N_2120);
nand U2593 (N_2593,N_957,N_1602);
or U2594 (N_2594,N_2313,N_2274);
or U2595 (N_2595,N_2119,N_2224);
xor U2596 (N_2596,N_597,N_1134);
or U2597 (N_2597,N_763,N_2297);
or U2598 (N_2598,N_2156,N_2237);
xor U2599 (N_2599,N_2356,N_802);
and U2600 (N_2600,N_2288,N_2032);
xnor U2601 (N_2601,N_2304,N_2127);
and U2602 (N_2602,N_1828,N_2319);
nor U2603 (N_2603,N_1489,N_2397);
nand U2604 (N_2604,In_1344,N_31);
or U2605 (N_2605,N_2180,N_2210);
or U2606 (N_2606,N_2391,N_2329);
nor U2607 (N_2607,N_306,N_2104);
or U2608 (N_2608,N_1962,N_1762);
nor U2609 (N_2609,In_276,N_2049);
nor U2610 (N_2610,In_2678,N_1780);
and U2611 (N_2611,N_2217,In_694);
and U2612 (N_2612,N_2035,N_2187);
xnor U2613 (N_2613,N_2340,N_1989);
nor U2614 (N_2614,N_1478,N_2230);
or U2615 (N_2615,N_1793,N_2383);
and U2616 (N_2616,N_1734,N_1599);
nor U2617 (N_2617,N_2320,N_2147);
nor U2618 (N_2618,N_2396,N_1535);
nand U2619 (N_2619,N_2047,N_676);
nand U2620 (N_2620,N_2214,N_2273);
or U2621 (N_2621,N_1640,N_654);
xnor U2622 (N_2622,In_2573,N_2131);
nor U2623 (N_2623,N_1860,N_2388);
nor U2624 (N_2624,N_1874,N_2181);
or U2625 (N_2625,N_1242,N_1967);
xor U2626 (N_2626,N_2194,N_2361);
xor U2627 (N_2627,N_2392,N_2330);
nand U2628 (N_2628,N_610,N_2251);
and U2629 (N_2629,N_2262,N_2333);
nand U2630 (N_2630,N_1196,N_321);
and U2631 (N_2631,N_2336,N_1285);
nand U2632 (N_2632,N_2186,N_2081);
nand U2633 (N_2633,N_2287,N_1787);
and U2634 (N_2634,N_2055,N_2372);
or U2635 (N_2635,N_2318,N_691);
nand U2636 (N_2636,N_2346,In_223);
xor U2637 (N_2637,N_1522,N_2183);
xnor U2638 (N_2638,N_2231,N_2177);
or U2639 (N_2639,N_2302,N_1676);
xnor U2640 (N_2640,N_2294,N_2351);
or U2641 (N_2641,N_2207,N_2311);
nor U2642 (N_2642,N_1815,In_1788);
nor U2643 (N_2643,N_339,N_2089);
xnor U2644 (N_2644,N_2222,N_1662);
nor U2645 (N_2645,N_2138,N_1293);
nand U2646 (N_2646,N_2335,N_2334);
and U2647 (N_2647,N_1012,N_1779);
or U2648 (N_2648,In_2753,N_2380);
xor U2649 (N_2649,N_1834,N_1922);
nor U2650 (N_2650,N_1482,N_286);
xor U2651 (N_2651,N_2191,In_1306);
nor U2652 (N_2652,N_1876,N_2360);
nand U2653 (N_2653,N_2269,N_2086);
xnor U2654 (N_2654,N_2385,N_1689);
or U2655 (N_2655,N_2054,N_2326);
or U2656 (N_2656,N_1058,N_2160);
xor U2657 (N_2657,N_2244,N_2379);
nand U2658 (N_2658,N_1875,N_2139);
or U2659 (N_2659,N_1626,In_2171);
xnor U2660 (N_2660,In_1096,N_1969);
or U2661 (N_2661,N_1716,N_2213);
xnor U2662 (N_2662,N_2151,N_1402);
and U2663 (N_2663,N_2223,N_2359);
or U2664 (N_2664,N_2364,N_2377);
xnor U2665 (N_2665,In_1531,N_2040);
and U2666 (N_2666,N_2169,N_1183);
xor U2667 (N_2667,N_2108,N_2176);
or U2668 (N_2668,N_2353,N_2350);
or U2669 (N_2669,N_2145,N_2238);
xor U2670 (N_2670,N_475,In_1872);
nand U2671 (N_2671,N_1613,N_2332);
xor U2672 (N_2672,N_2100,N_2189);
nand U2673 (N_2673,N_2173,N_2101);
or U2674 (N_2674,N_2344,N_1952);
and U2675 (N_2675,N_349,N_2395);
and U2676 (N_2676,N_2135,N_2312);
nor U2677 (N_2677,In_832,N_2295);
nand U2678 (N_2678,N_2354,N_1164);
nand U2679 (N_2679,N_2242,N_2110);
nor U2680 (N_2680,N_901,N_1589);
nand U2681 (N_2681,N_1206,N_2307);
nor U2682 (N_2682,In_2123,N_2208);
nor U2683 (N_2683,In_2804,N_1893);
or U2684 (N_2684,In_1477,N_1848);
xnor U2685 (N_2685,N_2154,N_2300);
xor U2686 (N_2686,In_567,N_1870);
and U2687 (N_2687,N_2338,N_2277);
nand U2688 (N_2688,N_1758,N_2116);
or U2689 (N_2689,N_177,N_1574);
nor U2690 (N_2690,N_1972,N_2321);
nor U2691 (N_2691,N_71,N_1732);
and U2692 (N_2692,N_1145,N_2061);
or U2693 (N_2693,N_2137,N_2171);
or U2694 (N_2694,In_2980,N_1235);
nand U2695 (N_2695,N_2281,N_1528);
nand U2696 (N_2696,N_1837,N_1005);
or U2697 (N_2697,N_1320,N_2129);
nor U2698 (N_2698,N_2256,In_2629);
xor U2699 (N_2699,In_1982,N_1625);
xor U2700 (N_2700,N_2682,N_2619);
nor U2701 (N_2701,N_2519,N_2654);
nand U2702 (N_2702,N_2448,N_2464);
nor U2703 (N_2703,N_2475,N_2628);
nand U2704 (N_2704,N_2529,N_2407);
and U2705 (N_2705,N_2492,N_2653);
or U2706 (N_2706,N_2563,N_2510);
nand U2707 (N_2707,N_2651,N_2517);
and U2708 (N_2708,N_2587,N_2616);
or U2709 (N_2709,N_2440,N_2692);
or U2710 (N_2710,N_2441,N_2545);
and U2711 (N_2711,N_2466,N_2561);
nor U2712 (N_2712,N_2627,N_2662);
nand U2713 (N_2713,N_2611,N_2494);
nor U2714 (N_2714,N_2465,N_2579);
nor U2715 (N_2715,N_2637,N_2690);
nand U2716 (N_2716,N_2659,N_2671);
or U2717 (N_2717,N_2696,N_2412);
or U2718 (N_2718,N_2456,N_2687);
or U2719 (N_2719,N_2567,N_2639);
and U2720 (N_2720,N_2461,N_2427);
nand U2721 (N_2721,N_2485,N_2585);
nor U2722 (N_2722,N_2689,N_2525);
and U2723 (N_2723,N_2406,N_2454);
nand U2724 (N_2724,N_2468,N_2531);
nand U2725 (N_2725,N_2450,N_2413);
or U2726 (N_2726,N_2566,N_2697);
nor U2727 (N_2727,N_2430,N_2562);
xnor U2728 (N_2728,N_2649,N_2449);
and U2729 (N_2729,N_2433,N_2674);
and U2730 (N_2730,N_2679,N_2578);
and U2731 (N_2731,N_2535,N_2400);
nand U2732 (N_2732,N_2688,N_2591);
or U2733 (N_2733,N_2534,N_2685);
or U2734 (N_2734,N_2621,N_2589);
or U2735 (N_2735,N_2558,N_2451);
nor U2736 (N_2736,N_2644,N_2571);
nand U2737 (N_2737,N_2486,N_2640);
nand U2738 (N_2738,N_2452,N_2540);
nor U2739 (N_2739,N_2565,N_2421);
or U2740 (N_2740,N_2559,N_2469);
nor U2741 (N_2741,N_2414,N_2513);
nor U2742 (N_2742,N_2583,N_2691);
nand U2743 (N_2743,N_2522,N_2613);
or U2744 (N_2744,N_2422,N_2553);
or U2745 (N_2745,N_2698,N_2472);
xnor U2746 (N_2746,N_2680,N_2675);
nor U2747 (N_2747,N_2439,N_2425);
nor U2748 (N_2748,N_2624,N_2676);
nand U2749 (N_2749,N_2474,N_2408);
and U2750 (N_2750,N_2462,N_2532);
nor U2751 (N_2751,N_2600,N_2602);
and U2752 (N_2752,N_2577,N_2645);
and U2753 (N_2753,N_2409,N_2515);
xnor U2754 (N_2754,N_2542,N_2614);
and U2755 (N_2755,N_2509,N_2521);
or U2756 (N_2756,N_2656,N_2516);
and U2757 (N_2757,N_2479,N_2547);
xor U2758 (N_2758,N_2543,N_2592);
and U2759 (N_2759,N_2491,N_2481);
nand U2760 (N_2760,N_2463,N_2514);
and U2761 (N_2761,N_2677,N_2528);
or U2762 (N_2762,N_2555,N_2503);
xor U2763 (N_2763,N_2478,N_2695);
nor U2764 (N_2764,N_2620,N_2664);
or U2765 (N_2765,N_2416,N_2554);
and U2766 (N_2766,N_2551,N_2699);
nand U2767 (N_2767,N_2552,N_2437);
and U2768 (N_2768,N_2593,N_2471);
and U2769 (N_2769,N_2467,N_2537);
nand U2770 (N_2770,N_2663,N_2693);
nor U2771 (N_2771,N_2536,N_2527);
nor U2772 (N_2772,N_2588,N_2505);
xnor U2773 (N_2773,N_2499,N_2501);
xnor U2774 (N_2774,N_2569,N_2584);
nand U2775 (N_2775,N_2580,N_2417);
nor U2776 (N_2776,N_2670,N_2657);
nand U2777 (N_2777,N_2520,N_2502);
or U2778 (N_2778,N_2668,N_2405);
nor U2779 (N_2779,N_2590,N_2538);
or U2780 (N_2780,N_2477,N_2420);
and U2781 (N_2781,N_2442,N_2672);
xor U2782 (N_2782,N_2546,N_2606);
nand U2783 (N_2783,N_2630,N_2429);
and U2784 (N_2784,N_2594,N_2678);
nand U2785 (N_2785,N_2550,N_2493);
and U2786 (N_2786,N_2660,N_2576);
or U2787 (N_2787,N_2453,N_2431);
xnor U2788 (N_2788,N_2560,N_2496);
or U2789 (N_2789,N_2597,N_2459);
and U2790 (N_2790,N_2632,N_2615);
and U2791 (N_2791,N_2419,N_2548);
nor U2792 (N_2792,N_2596,N_2638);
nand U2793 (N_2793,N_2432,N_2618);
or U2794 (N_2794,N_2473,N_2426);
or U2795 (N_2795,N_2488,N_2612);
or U2796 (N_2796,N_2610,N_2533);
nand U2797 (N_2797,N_2623,N_2666);
and U2798 (N_2798,N_2633,N_2444);
nand U2799 (N_2799,N_2411,N_2457);
nand U2800 (N_2800,N_2557,N_2530);
nor U2801 (N_2801,N_2617,N_2476);
nand U2802 (N_2802,N_2482,N_2625);
or U2803 (N_2803,N_2603,N_2631);
nand U2804 (N_2804,N_2498,N_2490);
or U2805 (N_2805,N_2646,N_2575);
nor U2806 (N_2806,N_2549,N_2683);
xor U2807 (N_2807,N_2572,N_2489);
xor U2808 (N_2808,N_2665,N_2605);
or U2809 (N_2809,N_2655,N_2641);
nor U2810 (N_2810,N_2402,N_2629);
and U2811 (N_2811,N_2673,N_2595);
nand U2812 (N_2812,N_2667,N_2460);
or U2813 (N_2813,N_2648,N_2573);
or U2814 (N_2814,N_2607,N_2508);
nand U2815 (N_2815,N_2523,N_2404);
or U2816 (N_2816,N_2650,N_2445);
and U2817 (N_2817,N_2446,N_2434);
xnor U2818 (N_2818,N_2541,N_2506);
nor U2819 (N_2819,N_2470,N_2599);
xor U2820 (N_2820,N_2669,N_2511);
nand U2821 (N_2821,N_2626,N_2608);
or U2822 (N_2822,N_2410,N_2694);
and U2823 (N_2823,N_2568,N_2539);
nor U2824 (N_2824,N_2647,N_2681);
nor U2825 (N_2825,N_2643,N_2661);
xnor U2826 (N_2826,N_2497,N_2526);
or U2827 (N_2827,N_2642,N_2423);
and U2828 (N_2828,N_2604,N_2564);
or U2829 (N_2829,N_2458,N_2487);
and U2830 (N_2830,N_2636,N_2447);
and U2831 (N_2831,N_2480,N_2544);
nor U2832 (N_2832,N_2512,N_2652);
and U2833 (N_2833,N_2609,N_2428);
or U2834 (N_2834,N_2518,N_2635);
nand U2835 (N_2835,N_2483,N_2436);
or U2836 (N_2836,N_2401,N_2443);
nor U2837 (N_2837,N_2438,N_2686);
or U2838 (N_2838,N_2582,N_2418);
xor U2839 (N_2839,N_2570,N_2524);
nand U2840 (N_2840,N_2598,N_2581);
nor U2841 (N_2841,N_2424,N_2601);
nand U2842 (N_2842,N_2507,N_2500);
nor U2843 (N_2843,N_2658,N_2495);
xor U2844 (N_2844,N_2415,N_2622);
nand U2845 (N_2845,N_2484,N_2455);
nor U2846 (N_2846,N_2435,N_2684);
xor U2847 (N_2847,N_2556,N_2504);
nor U2848 (N_2848,N_2634,N_2586);
and U2849 (N_2849,N_2403,N_2574);
nor U2850 (N_2850,N_2450,N_2544);
nand U2851 (N_2851,N_2458,N_2472);
or U2852 (N_2852,N_2530,N_2534);
or U2853 (N_2853,N_2642,N_2496);
or U2854 (N_2854,N_2584,N_2623);
or U2855 (N_2855,N_2597,N_2564);
nor U2856 (N_2856,N_2469,N_2633);
nor U2857 (N_2857,N_2638,N_2463);
nand U2858 (N_2858,N_2582,N_2444);
and U2859 (N_2859,N_2403,N_2540);
or U2860 (N_2860,N_2678,N_2570);
xor U2861 (N_2861,N_2626,N_2501);
and U2862 (N_2862,N_2412,N_2453);
nor U2863 (N_2863,N_2578,N_2427);
and U2864 (N_2864,N_2538,N_2474);
and U2865 (N_2865,N_2539,N_2684);
or U2866 (N_2866,N_2400,N_2438);
nand U2867 (N_2867,N_2554,N_2443);
nand U2868 (N_2868,N_2625,N_2606);
nand U2869 (N_2869,N_2697,N_2514);
xnor U2870 (N_2870,N_2419,N_2471);
xnor U2871 (N_2871,N_2470,N_2420);
nand U2872 (N_2872,N_2419,N_2624);
xnor U2873 (N_2873,N_2617,N_2548);
or U2874 (N_2874,N_2672,N_2525);
xor U2875 (N_2875,N_2630,N_2434);
and U2876 (N_2876,N_2503,N_2407);
nand U2877 (N_2877,N_2683,N_2669);
nand U2878 (N_2878,N_2504,N_2419);
xor U2879 (N_2879,N_2443,N_2457);
nor U2880 (N_2880,N_2568,N_2676);
xnor U2881 (N_2881,N_2626,N_2485);
xnor U2882 (N_2882,N_2564,N_2429);
or U2883 (N_2883,N_2658,N_2419);
and U2884 (N_2884,N_2584,N_2421);
nand U2885 (N_2885,N_2447,N_2456);
or U2886 (N_2886,N_2480,N_2645);
nor U2887 (N_2887,N_2666,N_2557);
nand U2888 (N_2888,N_2692,N_2405);
nor U2889 (N_2889,N_2421,N_2661);
xnor U2890 (N_2890,N_2570,N_2654);
nor U2891 (N_2891,N_2698,N_2547);
xor U2892 (N_2892,N_2641,N_2640);
or U2893 (N_2893,N_2667,N_2404);
xor U2894 (N_2894,N_2669,N_2630);
nand U2895 (N_2895,N_2459,N_2519);
xor U2896 (N_2896,N_2624,N_2412);
or U2897 (N_2897,N_2628,N_2584);
and U2898 (N_2898,N_2467,N_2425);
xor U2899 (N_2899,N_2552,N_2635);
nand U2900 (N_2900,N_2628,N_2664);
or U2901 (N_2901,N_2483,N_2503);
or U2902 (N_2902,N_2437,N_2587);
nor U2903 (N_2903,N_2574,N_2652);
xor U2904 (N_2904,N_2585,N_2572);
and U2905 (N_2905,N_2541,N_2574);
or U2906 (N_2906,N_2557,N_2551);
xor U2907 (N_2907,N_2570,N_2539);
and U2908 (N_2908,N_2525,N_2575);
xnor U2909 (N_2909,N_2451,N_2478);
nor U2910 (N_2910,N_2524,N_2568);
nand U2911 (N_2911,N_2442,N_2414);
nor U2912 (N_2912,N_2408,N_2674);
xnor U2913 (N_2913,N_2650,N_2560);
nand U2914 (N_2914,N_2423,N_2668);
nor U2915 (N_2915,N_2492,N_2445);
and U2916 (N_2916,N_2472,N_2688);
nand U2917 (N_2917,N_2525,N_2476);
or U2918 (N_2918,N_2666,N_2411);
nor U2919 (N_2919,N_2508,N_2411);
and U2920 (N_2920,N_2503,N_2432);
nor U2921 (N_2921,N_2598,N_2517);
nand U2922 (N_2922,N_2444,N_2673);
xnor U2923 (N_2923,N_2483,N_2460);
and U2924 (N_2924,N_2563,N_2542);
nor U2925 (N_2925,N_2634,N_2506);
xor U2926 (N_2926,N_2556,N_2588);
nand U2927 (N_2927,N_2682,N_2465);
and U2928 (N_2928,N_2477,N_2415);
nor U2929 (N_2929,N_2500,N_2662);
and U2930 (N_2930,N_2403,N_2473);
or U2931 (N_2931,N_2663,N_2457);
nand U2932 (N_2932,N_2470,N_2593);
and U2933 (N_2933,N_2417,N_2640);
nand U2934 (N_2934,N_2404,N_2493);
nor U2935 (N_2935,N_2598,N_2461);
or U2936 (N_2936,N_2505,N_2439);
nor U2937 (N_2937,N_2698,N_2490);
xnor U2938 (N_2938,N_2535,N_2508);
xnor U2939 (N_2939,N_2436,N_2548);
and U2940 (N_2940,N_2643,N_2652);
nor U2941 (N_2941,N_2502,N_2424);
nor U2942 (N_2942,N_2421,N_2516);
nor U2943 (N_2943,N_2444,N_2609);
and U2944 (N_2944,N_2638,N_2438);
or U2945 (N_2945,N_2632,N_2576);
nand U2946 (N_2946,N_2537,N_2564);
xnor U2947 (N_2947,N_2400,N_2530);
nor U2948 (N_2948,N_2405,N_2457);
nor U2949 (N_2949,N_2474,N_2555);
and U2950 (N_2950,N_2586,N_2633);
and U2951 (N_2951,N_2659,N_2490);
xor U2952 (N_2952,N_2690,N_2604);
and U2953 (N_2953,N_2414,N_2531);
nor U2954 (N_2954,N_2592,N_2552);
or U2955 (N_2955,N_2559,N_2576);
xnor U2956 (N_2956,N_2637,N_2487);
nor U2957 (N_2957,N_2661,N_2537);
or U2958 (N_2958,N_2493,N_2428);
nor U2959 (N_2959,N_2583,N_2501);
nand U2960 (N_2960,N_2479,N_2541);
or U2961 (N_2961,N_2601,N_2667);
nor U2962 (N_2962,N_2503,N_2695);
or U2963 (N_2963,N_2531,N_2603);
nand U2964 (N_2964,N_2563,N_2468);
nand U2965 (N_2965,N_2402,N_2669);
xnor U2966 (N_2966,N_2535,N_2579);
nand U2967 (N_2967,N_2609,N_2433);
or U2968 (N_2968,N_2551,N_2431);
and U2969 (N_2969,N_2495,N_2558);
or U2970 (N_2970,N_2639,N_2525);
nand U2971 (N_2971,N_2462,N_2529);
nand U2972 (N_2972,N_2635,N_2532);
xor U2973 (N_2973,N_2417,N_2491);
and U2974 (N_2974,N_2529,N_2535);
nand U2975 (N_2975,N_2509,N_2615);
nor U2976 (N_2976,N_2469,N_2641);
or U2977 (N_2977,N_2441,N_2429);
or U2978 (N_2978,N_2632,N_2657);
nand U2979 (N_2979,N_2552,N_2675);
and U2980 (N_2980,N_2522,N_2618);
and U2981 (N_2981,N_2488,N_2638);
nand U2982 (N_2982,N_2557,N_2624);
or U2983 (N_2983,N_2665,N_2569);
or U2984 (N_2984,N_2495,N_2667);
xnor U2985 (N_2985,N_2626,N_2599);
xnor U2986 (N_2986,N_2688,N_2578);
and U2987 (N_2987,N_2591,N_2417);
nand U2988 (N_2988,N_2498,N_2519);
nor U2989 (N_2989,N_2681,N_2453);
xnor U2990 (N_2990,N_2413,N_2503);
and U2991 (N_2991,N_2640,N_2610);
nor U2992 (N_2992,N_2549,N_2561);
and U2993 (N_2993,N_2618,N_2470);
nor U2994 (N_2994,N_2552,N_2422);
nor U2995 (N_2995,N_2506,N_2659);
and U2996 (N_2996,N_2417,N_2456);
nor U2997 (N_2997,N_2574,N_2482);
nor U2998 (N_2998,N_2545,N_2468);
xnor U2999 (N_2999,N_2423,N_2431);
and U3000 (N_3000,N_2845,N_2933);
nand U3001 (N_3001,N_2816,N_2736);
nand U3002 (N_3002,N_2829,N_2946);
nand U3003 (N_3003,N_2938,N_2777);
or U3004 (N_3004,N_2744,N_2835);
nand U3005 (N_3005,N_2909,N_2717);
nor U3006 (N_3006,N_2735,N_2770);
xor U3007 (N_3007,N_2935,N_2721);
xnor U3008 (N_3008,N_2997,N_2983);
nor U3009 (N_3009,N_2928,N_2906);
or U3010 (N_3010,N_2807,N_2895);
nor U3011 (N_3011,N_2888,N_2806);
nor U3012 (N_3012,N_2804,N_2950);
nor U3013 (N_3013,N_2746,N_2989);
xor U3014 (N_3014,N_2964,N_2755);
nor U3015 (N_3015,N_2756,N_2759);
nand U3016 (N_3016,N_2903,N_2738);
nand U3017 (N_3017,N_2971,N_2968);
xnor U3018 (N_3018,N_2712,N_2982);
nand U3019 (N_3019,N_2802,N_2977);
xnor U3020 (N_3020,N_2726,N_2711);
nand U3021 (N_3021,N_2958,N_2793);
nor U3022 (N_3022,N_2956,N_2841);
nand U3023 (N_3023,N_2832,N_2762);
xor U3024 (N_3024,N_2716,N_2889);
nor U3025 (N_3025,N_2809,N_2942);
xor U3026 (N_3026,N_2857,N_2827);
nor U3027 (N_3027,N_2723,N_2820);
and U3028 (N_3028,N_2969,N_2800);
nor U3029 (N_3029,N_2730,N_2913);
or U3030 (N_3030,N_2996,N_2731);
xor U3031 (N_3031,N_2954,N_2885);
nor U3032 (N_3032,N_2779,N_2824);
and U3033 (N_3033,N_2704,N_2877);
xor U3034 (N_3034,N_2880,N_2702);
or U3035 (N_3035,N_2973,N_2776);
nand U3036 (N_3036,N_2797,N_2853);
or U3037 (N_3037,N_2878,N_2765);
and U3038 (N_3038,N_2749,N_2761);
and U3039 (N_3039,N_2992,N_2972);
and U3040 (N_3040,N_2985,N_2767);
nor U3041 (N_3041,N_2825,N_2862);
and U3042 (N_3042,N_2796,N_2760);
and U3043 (N_3043,N_2917,N_2894);
and U3044 (N_3044,N_2805,N_2869);
nand U3045 (N_3045,N_2907,N_2720);
xnor U3046 (N_3046,N_2941,N_2739);
nand U3047 (N_3047,N_2791,N_2848);
or U3048 (N_3048,N_2863,N_2833);
nand U3049 (N_3049,N_2814,N_2734);
xor U3050 (N_3050,N_2953,N_2998);
xnor U3051 (N_3051,N_2844,N_2701);
nor U3052 (N_3052,N_2748,N_2811);
nor U3053 (N_3053,N_2999,N_2715);
and U3054 (N_3054,N_2929,N_2801);
and U3055 (N_3055,N_2974,N_2925);
and U3056 (N_3056,N_2708,N_2790);
or U3057 (N_3057,N_2817,N_2775);
nor U3058 (N_3058,N_2963,N_2764);
nor U3059 (N_3059,N_2706,N_2781);
or U3060 (N_3060,N_2849,N_2991);
nor U3061 (N_3061,N_2927,N_2709);
nand U3062 (N_3062,N_2873,N_2766);
nand U3063 (N_3063,N_2831,N_2856);
or U3064 (N_3064,N_2947,N_2826);
and U3065 (N_3065,N_2897,N_2919);
xnor U3066 (N_3066,N_2965,N_2931);
nor U3067 (N_3067,N_2784,N_2923);
nand U3068 (N_3068,N_2966,N_2828);
nand U3069 (N_3069,N_2741,N_2733);
nand U3070 (N_3070,N_2757,N_2910);
xnor U3071 (N_3071,N_2945,N_2851);
xnor U3072 (N_3072,N_2879,N_2768);
nand U3073 (N_3073,N_2700,N_2934);
xnor U3074 (N_3074,N_2978,N_2798);
nor U3075 (N_3075,N_2957,N_2850);
xnor U3076 (N_3076,N_2890,N_2914);
and U3077 (N_3077,N_2728,N_2887);
nor U3078 (N_3078,N_2815,N_2854);
nor U3079 (N_3079,N_2944,N_2955);
or U3080 (N_3080,N_2898,N_2799);
xor U3081 (N_3081,N_2896,N_2745);
nor U3082 (N_3082,N_2703,N_2724);
nand U3083 (N_3083,N_2994,N_2922);
nand U3084 (N_3084,N_2722,N_2782);
nor U3085 (N_3085,N_2740,N_2818);
or U3086 (N_3086,N_2905,N_2795);
xnor U3087 (N_3087,N_2876,N_2714);
xnor U3088 (N_3088,N_2866,N_2838);
nand U3089 (N_3089,N_2836,N_2892);
or U3090 (N_3090,N_2752,N_2840);
or U3091 (N_3091,N_2803,N_2773);
xor U3092 (N_3092,N_2860,N_2732);
nor U3093 (N_3093,N_2900,N_2753);
or U3094 (N_3094,N_2839,N_2940);
xnor U3095 (N_3095,N_2912,N_2769);
nor U3096 (N_3096,N_2859,N_2995);
or U3097 (N_3097,N_2864,N_2976);
xor U3098 (N_3098,N_2975,N_2774);
nand U3099 (N_3099,N_2908,N_2719);
nand U3100 (N_3100,N_2710,N_2743);
and U3101 (N_3101,N_2987,N_2727);
xor U3102 (N_3102,N_2874,N_2785);
and U3103 (N_3103,N_2808,N_2871);
and U3104 (N_3104,N_2902,N_2921);
or U3105 (N_3105,N_2884,N_2962);
nand U3106 (N_3106,N_2812,N_2932);
and U3107 (N_3107,N_2705,N_2920);
nor U3108 (N_3108,N_2868,N_2883);
or U3109 (N_3109,N_2891,N_2783);
or U3110 (N_3110,N_2961,N_2916);
nor U3111 (N_3111,N_2911,N_2821);
or U3112 (N_3112,N_2758,N_2990);
and U3113 (N_3113,N_2926,N_2980);
or U3114 (N_3114,N_2788,N_2875);
and U3115 (N_3115,N_2915,N_2713);
and U3116 (N_3116,N_2904,N_2842);
nor U3117 (N_3117,N_2936,N_2967);
xor U3118 (N_3118,N_2948,N_2852);
and U3119 (N_3119,N_2794,N_2846);
or U3120 (N_3120,N_2867,N_2729);
xnor U3121 (N_3121,N_2789,N_2886);
or U3122 (N_3122,N_2882,N_2893);
and U3123 (N_3123,N_2861,N_2718);
or U3124 (N_3124,N_2855,N_2949);
or U3125 (N_3125,N_2813,N_2858);
nand U3126 (N_3126,N_2899,N_2986);
nor U3127 (N_3127,N_2725,N_2970);
or U3128 (N_3128,N_2747,N_2754);
and U3129 (N_3129,N_2837,N_2865);
nand U3130 (N_3130,N_2772,N_2930);
nor U3131 (N_3131,N_2939,N_2918);
and U3132 (N_3132,N_2843,N_2834);
or U3133 (N_3133,N_2901,N_2771);
nand U3134 (N_3134,N_2822,N_2737);
and U3135 (N_3135,N_2707,N_2881);
or U3136 (N_3136,N_2872,N_2810);
and U3137 (N_3137,N_2786,N_2952);
nand U3138 (N_3138,N_2951,N_2787);
nor U3139 (N_3139,N_2778,N_2847);
or U3140 (N_3140,N_2830,N_2792);
or U3141 (N_3141,N_2984,N_2751);
nor U3142 (N_3142,N_2742,N_2981);
and U3143 (N_3143,N_2993,N_2937);
nand U3144 (N_3144,N_2763,N_2819);
and U3145 (N_3145,N_2750,N_2780);
nor U3146 (N_3146,N_2979,N_2870);
and U3147 (N_3147,N_2988,N_2960);
nand U3148 (N_3148,N_2943,N_2959);
nor U3149 (N_3149,N_2823,N_2924);
nor U3150 (N_3150,N_2982,N_2903);
xnor U3151 (N_3151,N_2820,N_2810);
or U3152 (N_3152,N_2832,N_2789);
or U3153 (N_3153,N_2888,N_2730);
nor U3154 (N_3154,N_2844,N_2711);
and U3155 (N_3155,N_2771,N_2970);
nand U3156 (N_3156,N_2788,N_2893);
or U3157 (N_3157,N_2942,N_2720);
or U3158 (N_3158,N_2720,N_2794);
nor U3159 (N_3159,N_2810,N_2992);
xnor U3160 (N_3160,N_2720,N_2851);
nand U3161 (N_3161,N_2888,N_2793);
and U3162 (N_3162,N_2916,N_2915);
nor U3163 (N_3163,N_2833,N_2834);
xnor U3164 (N_3164,N_2983,N_2970);
xor U3165 (N_3165,N_2967,N_2881);
and U3166 (N_3166,N_2787,N_2883);
and U3167 (N_3167,N_2990,N_2818);
xor U3168 (N_3168,N_2796,N_2710);
and U3169 (N_3169,N_2906,N_2980);
nand U3170 (N_3170,N_2947,N_2788);
and U3171 (N_3171,N_2833,N_2937);
nor U3172 (N_3172,N_2895,N_2931);
xnor U3173 (N_3173,N_2814,N_2995);
and U3174 (N_3174,N_2908,N_2896);
xor U3175 (N_3175,N_2972,N_2880);
xor U3176 (N_3176,N_2730,N_2814);
nor U3177 (N_3177,N_2973,N_2705);
or U3178 (N_3178,N_2911,N_2732);
xnor U3179 (N_3179,N_2743,N_2962);
or U3180 (N_3180,N_2731,N_2730);
xnor U3181 (N_3181,N_2812,N_2979);
and U3182 (N_3182,N_2732,N_2773);
and U3183 (N_3183,N_2703,N_2842);
and U3184 (N_3184,N_2727,N_2909);
xnor U3185 (N_3185,N_2752,N_2800);
xor U3186 (N_3186,N_2748,N_2834);
nor U3187 (N_3187,N_2883,N_2783);
and U3188 (N_3188,N_2950,N_2810);
and U3189 (N_3189,N_2931,N_2850);
nand U3190 (N_3190,N_2899,N_2739);
xor U3191 (N_3191,N_2959,N_2808);
or U3192 (N_3192,N_2958,N_2888);
or U3193 (N_3193,N_2706,N_2755);
xor U3194 (N_3194,N_2999,N_2868);
nor U3195 (N_3195,N_2733,N_2980);
or U3196 (N_3196,N_2907,N_2791);
or U3197 (N_3197,N_2972,N_2709);
nor U3198 (N_3198,N_2728,N_2755);
or U3199 (N_3199,N_2762,N_2725);
or U3200 (N_3200,N_2920,N_2815);
nor U3201 (N_3201,N_2702,N_2962);
xnor U3202 (N_3202,N_2836,N_2891);
nor U3203 (N_3203,N_2950,N_2709);
nor U3204 (N_3204,N_2884,N_2859);
and U3205 (N_3205,N_2873,N_2993);
xnor U3206 (N_3206,N_2954,N_2785);
xor U3207 (N_3207,N_2955,N_2941);
nand U3208 (N_3208,N_2912,N_2956);
and U3209 (N_3209,N_2754,N_2769);
nor U3210 (N_3210,N_2872,N_2958);
and U3211 (N_3211,N_2911,N_2962);
and U3212 (N_3212,N_2989,N_2835);
and U3213 (N_3213,N_2808,N_2887);
or U3214 (N_3214,N_2819,N_2958);
nand U3215 (N_3215,N_2877,N_2718);
nor U3216 (N_3216,N_2846,N_2968);
nand U3217 (N_3217,N_2843,N_2719);
or U3218 (N_3218,N_2958,N_2922);
or U3219 (N_3219,N_2907,N_2854);
or U3220 (N_3220,N_2734,N_2765);
and U3221 (N_3221,N_2764,N_2912);
xnor U3222 (N_3222,N_2759,N_2922);
and U3223 (N_3223,N_2735,N_2736);
or U3224 (N_3224,N_2919,N_2816);
nand U3225 (N_3225,N_2724,N_2727);
nand U3226 (N_3226,N_2967,N_2998);
nor U3227 (N_3227,N_2883,N_2797);
xnor U3228 (N_3228,N_2903,N_2864);
xnor U3229 (N_3229,N_2722,N_2854);
or U3230 (N_3230,N_2804,N_2998);
and U3231 (N_3231,N_2794,N_2874);
and U3232 (N_3232,N_2703,N_2943);
and U3233 (N_3233,N_2980,N_2762);
or U3234 (N_3234,N_2753,N_2721);
and U3235 (N_3235,N_2722,N_2967);
nor U3236 (N_3236,N_2759,N_2817);
nand U3237 (N_3237,N_2767,N_2839);
xor U3238 (N_3238,N_2763,N_2973);
or U3239 (N_3239,N_2908,N_2756);
or U3240 (N_3240,N_2875,N_2842);
or U3241 (N_3241,N_2713,N_2981);
xnor U3242 (N_3242,N_2795,N_2907);
xor U3243 (N_3243,N_2851,N_2743);
and U3244 (N_3244,N_2857,N_2944);
nor U3245 (N_3245,N_2803,N_2883);
xnor U3246 (N_3246,N_2804,N_2748);
xor U3247 (N_3247,N_2897,N_2926);
or U3248 (N_3248,N_2824,N_2741);
xor U3249 (N_3249,N_2718,N_2828);
and U3250 (N_3250,N_2738,N_2796);
nor U3251 (N_3251,N_2812,N_2946);
nor U3252 (N_3252,N_2931,N_2992);
nor U3253 (N_3253,N_2949,N_2911);
and U3254 (N_3254,N_2747,N_2954);
nor U3255 (N_3255,N_2728,N_2710);
nand U3256 (N_3256,N_2972,N_2945);
or U3257 (N_3257,N_2846,N_2895);
nor U3258 (N_3258,N_2797,N_2898);
nor U3259 (N_3259,N_2972,N_2776);
nand U3260 (N_3260,N_2868,N_2885);
nand U3261 (N_3261,N_2747,N_2845);
nand U3262 (N_3262,N_2955,N_2845);
nor U3263 (N_3263,N_2952,N_2744);
xor U3264 (N_3264,N_2942,N_2943);
or U3265 (N_3265,N_2739,N_2808);
nor U3266 (N_3266,N_2764,N_2783);
nand U3267 (N_3267,N_2766,N_2789);
xnor U3268 (N_3268,N_2878,N_2796);
nand U3269 (N_3269,N_2839,N_2842);
nand U3270 (N_3270,N_2872,N_2908);
or U3271 (N_3271,N_2831,N_2980);
and U3272 (N_3272,N_2757,N_2723);
nand U3273 (N_3273,N_2835,N_2917);
xnor U3274 (N_3274,N_2906,N_2875);
and U3275 (N_3275,N_2930,N_2964);
nand U3276 (N_3276,N_2917,N_2985);
or U3277 (N_3277,N_2968,N_2872);
and U3278 (N_3278,N_2955,N_2863);
or U3279 (N_3279,N_2825,N_2982);
nor U3280 (N_3280,N_2892,N_2718);
nand U3281 (N_3281,N_2803,N_2717);
or U3282 (N_3282,N_2985,N_2726);
and U3283 (N_3283,N_2968,N_2825);
nor U3284 (N_3284,N_2793,N_2997);
xnor U3285 (N_3285,N_2920,N_2965);
nor U3286 (N_3286,N_2980,N_2975);
nand U3287 (N_3287,N_2898,N_2858);
nand U3288 (N_3288,N_2838,N_2796);
xnor U3289 (N_3289,N_2754,N_2954);
or U3290 (N_3290,N_2888,N_2988);
nand U3291 (N_3291,N_2980,N_2851);
and U3292 (N_3292,N_2714,N_2986);
and U3293 (N_3293,N_2868,N_2717);
or U3294 (N_3294,N_2955,N_2700);
and U3295 (N_3295,N_2958,N_2844);
nand U3296 (N_3296,N_2901,N_2759);
xor U3297 (N_3297,N_2786,N_2909);
nor U3298 (N_3298,N_2947,N_2951);
nand U3299 (N_3299,N_2726,N_2977);
xor U3300 (N_3300,N_3143,N_3096);
nand U3301 (N_3301,N_3038,N_3190);
or U3302 (N_3302,N_3159,N_3211);
nand U3303 (N_3303,N_3101,N_3138);
and U3304 (N_3304,N_3031,N_3186);
xor U3305 (N_3305,N_3149,N_3081);
nor U3306 (N_3306,N_3039,N_3108);
and U3307 (N_3307,N_3178,N_3153);
nand U3308 (N_3308,N_3253,N_3046);
nor U3309 (N_3309,N_3237,N_3158);
or U3310 (N_3310,N_3268,N_3181);
nor U3311 (N_3311,N_3242,N_3209);
nand U3312 (N_3312,N_3239,N_3142);
nand U3313 (N_3313,N_3174,N_3000);
and U3314 (N_3314,N_3063,N_3210);
nor U3315 (N_3315,N_3292,N_3119);
or U3316 (N_3316,N_3191,N_3020);
or U3317 (N_3317,N_3025,N_3150);
nand U3318 (N_3318,N_3040,N_3255);
nand U3319 (N_3319,N_3018,N_3092);
xor U3320 (N_3320,N_3276,N_3224);
and U3321 (N_3321,N_3064,N_3118);
or U3322 (N_3322,N_3011,N_3198);
or U3323 (N_3323,N_3244,N_3116);
nor U3324 (N_3324,N_3107,N_3157);
nor U3325 (N_3325,N_3279,N_3284);
xor U3326 (N_3326,N_3023,N_3016);
nand U3327 (N_3327,N_3007,N_3259);
xor U3328 (N_3328,N_3221,N_3275);
nand U3329 (N_3329,N_3067,N_3085);
nand U3330 (N_3330,N_3228,N_3294);
and U3331 (N_3331,N_3299,N_3047);
xor U3332 (N_3332,N_3124,N_3089);
xor U3333 (N_3333,N_3044,N_3225);
and U3334 (N_3334,N_3072,N_3162);
or U3335 (N_3335,N_3014,N_3182);
or U3336 (N_3336,N_3263,N_3298);
or U3337 (N_3337,N_3097,N_3117);
or U3338 (N_3338,N_3283,N_3206);
and U3339 (N_3339,N_3111,N_3013);
nor U3340 (N_3340,N_3261,N_3029);
nand U3341 (N_3341,N_3069,N_3288);
nand U3342 (N_3342,N_3098,N_3274);
xor U3343 (N_3343,N_3037,N_3144);
nor U3344 (N_3344,N_3235,N_3132);
nor U3345 (N_3345,N_3219,N_3160);
nand U3346 (N_3346,N_3155,N_3278);
or U3347 (N_3347,N_3262,N_3257);
nor U3348 (N_3348,N_3084,N_3269);
nand U3349 (N_3349,N_3080,N_3141);
or U3350 (N_3350,N_3002,N_3168);
nor U3351 (N_3351,N_3060,N_3215);
or U3352 (N_3352,N_3114,N_3019);
nand U3353 (N_3353,N_3035,N_3282);
nor U3354 (N_3354,N_3083,N_3280);
and U3355 (N_3355,N_3133,N_3171);
or U3356 (N_3356,N_3055,N_3166);
nand U3357 (N_3357,N_3012,N_3199);
nand U3358 (N_3358,N_3200,N_3105);
nand U3359 (N_3359,N_3252,N_3277);
xnor U3360 (N_3360,N_3147,N_3066);
and U3361 (N_3361,N_3214,N_3126);
xor U3362 (N_3362,N_3267,N_3043);
nand U3363 (N_3363,N_3249,N_3074);
or U3364 (N_3364,N_3054,N_3091);
or U3365 (N_3365,N_3183,N_3193);
nand U3366 (N_3366,N_3227,N_3231);
or U3367 (N_3367,N_3078,N_3194);
nor U3368 (N_3368,N_3172,N_3295);
nand U3369 (N_3369,N_3045,N_3256);
xor U3370 (N_3370,N_3030,N_3058);
or U3371 (N_3371,N_3165,N_3205);
nand U3372 (N_3372,N_3061,N_3129);
xor U3373 (N_3373,N_3015,N_3109);
and U3374 (N_3374,N_3192,N_3120);
nand U3375 (N_3375,N_3289,N_3123);
xor U3376 (N_3376,N_3139,N_3076);
xnor U3377 (N_3377,N_3003,N_3163);
nand U3378 (N_3378,N_3115,N_3042);
xnor U3379 (N_3379,N_3273,N_3093);
nor U3380 (N_3380,N_3296,N_3176);
nand U3381 (N_3381,N_3090,N_3232);
or U3382 (N_3382,N_3184,N_3195);
nor U3383 (N_3383,N_3135,N_3201);
xnor U3384 (N_3384,N_3033,N_3001);
nor U3385 (N_3385,N_3017,N_3075);
xor U3386 (N_3386,N_3286,N_3285);
or U3387 (N_3387,N_3112,N_3265);
and U3388 (N_3388,N_3202,N_3204);
nand U3389 (N_3389,N_3208,N_3071);
or U3390 (N_3390,N_3233,N_3036);
xnor U3391 (N_3391,N_3140,N_3099);
nand U3392 (N_3392,N_3173,N_3087);
nor U3393 (N_3393,N_3222,N_3290);
nand U3394 (N_3394,N_3052,N_3131);
nand U3395 (N_3395,N_3266,N_3254);
xor U3396 (N_3396,N_3041,N_3216);
nand U3397 (N_3397,N_3230,N_3152);
nor U3398 (N_3398,N_3170,N_3247);
and U3399 (N_3399,N_3229,N_3006);
and U3400 (N_3400,N_3212,N_3250);
or U3401 (N_3401,N_3125,N_3034);
nor U3402 (N_3402,N_3027,N_3024);
nor U3403 (N_3403,N_3258,N_3100);
and U3404 (N_3404,N_3010,N_3213);
xnor U3405 (N_3405,N_3028,N_3245);
and U3406 (N_3406,N_3136,N_3248);
or U3407 (N_3407,N_3271,N_3134);
nor U3408 (N_3408,N_3243,N_3110);
nor U3409 (N_3409,N_3022,N_3187);
xnor U3410 (N_3410,N_3161,N_3226);
nand U3411 (N_3411,N_3197,N_3217);
nor U3412 (N_3412,N_3137,N_3051);
xnor U3413 (N_3413,N_3106,N_3048);
xor U3414 (N_3414,N_3146,N_3009);
or U3415 (N_3415,N_3095,N_3234);
nor U3416 (N_3416,N_3121,N_3005);
xnor U3417 (N_3417,N_3026,N_3196);
nor U3418 (N_3418,N_3236,N_3082);
xor U3419 (N_3419,N_3287,N_3180);
nand U3420 (N_3420,N_3103,N_3070);
or U3421 (N_3421,N_3297,N_3088);
xor U3422 (N_3422,N_3102,N_3246);
xor U3423 (N_3423,N_3073,N_3050);
nor U3424 (N_3424,N_3175,N_3151);
nor U3425 (N_3425,N_3223,N_3004);
nand U3426 (N_3426,N_3203,N_3128);
or U3427 (N_3427,N_3240,N_3164);
nand U3428 (N_3428,N_3293,N_3104);
nand U3429 (N_3429,N_3086,N_3281);
and U3430 (N_3430,N_3156,N_3053);
nor U3431 (N_3431,N_3188,N_3065);
xnor U3432 (N_3432,N_3113,N_3218);
and U3433 (N_3433,N_3127,N_3154);
xnor U3434 (N_3434,N_3207,N_3179);
and U3435 (N_3435,N_3264,N_3270);
and U3436 (N_3436,N_3177,N_3291);
or U3437 (N_3437,N_3272,N_3068);
and U3438 (N_3438,N_3169,N_3238);
nand U3439 (N_3439,N_3057,N_3049);
nor U3440 (N_3440,N_3032,N_3122);
xnor U3441 (N_3441,N_3241,N_3008);
and U3442 (N_3442,N_3251,N_3077);
or U3443 (N_3443,N_3167,N_3145);
xor U3444 (N_3444,N_3059,N_3056);
and U3445 (N_3445,N_3220,N_3094);
and U3446 (N_3446,N_3130,N_3021);
or U3447 (N_3447,N_3079,N_3185);
xnor U3448 (N_3448,N_3189,N_3260);
or U3449 (N_3449,N_3062,N_3148);
and U3450 (N_3450,N_3039,N_3202);
xor U3451 (N_3451,N_3052,N_3205);
or U3452 (N_3452,N_3095,N_3236);
xor U3453 (N_3453,N_3181,N_3271);
or U3454 (N_3454,N_3239,N_3095);
or U3455 (N_3455,N_3004,N_3161);
xor U3456 (N_3456,N_3183,N_3069);
and U3457 (N_3457,N_3120,N_3091);
and U3458 (N_3458,N_3171,N_3053);
nor U3459 (N_3459,N_3064,N_3050);
xor U3460 (N_3460,N_3250,N_3001);
xnor U3461 (N_3461,N_3152,N_3094);
nand U3462 (N_3462,N_3265,N_3128);
or U3463 (N_3463,N_3061,N_3139);
xnor U3464 (N_3464,N_3217,N_3216);
xor U3465 (N_3465,N_3093,N_3241);
and U3466 (N_3466,N_3106,N_3158);
xor U3467 (N_3467,N_3123,N_3030);
nor U3468 (N_3468,N_3127,N_3073);
or U3469 (N_3469,N_3213,N_3274);
nor U3470 (N_3470,N_3143,N_3273);
xor U3471 (N_3471,N_3161,N_3188);
nor U3472 (N_3472,N_3094,N_3020);
xnor U3473 (N_3473,N_3124,N_3229);
xor U3474 (N_3474,N_3054,N_3043);
nand U3475 (N_3475,N_3159,N_3224);
nor U3476 (N_3476,N_3293,N_3248);
nand U3477 (N_3477,N_3238,N_3246);
xnor U3478 (N_3478,N_3027,N_3244);
xnor U3479 (N_3479,N_3259,N_3114);
nor U3480 (N_3480,N_3225,N_3059);
nor U3481 (N_3481,N_3236,N_3197);
nor U3482 (N_3482,N_3127,N_3121);
and U3483 (N_3483,N_3195,N_3185);
xnor U3484 (N_3484,N_3079,N_3174);
and U3485 (N_3485,N_3184,N_3128);
and U3486 (N_3486,N_3294,N_3191);
and U3487 (N_3487,N_3267,N_3002);
nor U3488 (N_3488,N_3028,N_3225);
nor U3489 (N_3489,N_3297,N_3153);
xnor U3490 (N_3490,N_3280,N_3141);
or U3491 (N_3491,N_3129,N_3054);
and U3492 (N_3492,N_3237,N_3072);
nor U3493 (N_3493,N_3159,N_3252);
xor U3494 (N_3494,N_3204,N_3151);
nor U3495 (N_3495,N_3262,N_3196);
xnor U3496 (N_3496,N_3291,N_3083);
xnor U3497 (N_3497,N_3159,N_3297);
or U3498 (N_3498,N_3128,N_3281);
or U3499 (N_3499,N_3283,N_3031);
xnor U3500 (N_3500,N_3033,N_3089);
and U3501 (N_3501,N_3272,N_3286);
and U3502 (N_3502,N_3298,N_3245);
and U3503 (N_3503,N_3183,N_3006);
nor U3504 (N_3504,N_3039,N_3025);
or U3505 (N_3505,N_3272,N_3082);
and U3506 (N_3506,N_3244,N_3020);
and U3507 (N_3507,N_3103,N_3295);
xor U3508 (N_3508,N_3233,N_3120);
nor U3509 (N_3509,N_3024,N_3183);
or U3510 (N_3510,N_3237,N_3140);
or U3511 (N_3511,N_3251,N_3171);
and U3512 (N_3512,N_3094,N_3024);
nor U3513 (N_3513,N_3169,N_3124);
nor U3514 (N_3514,N_3257,N_3296);
and U3515 (N_3515,N_3043,N_3114);
or U3516 (N_3516,N_3177,N_3257);
and U3517 (N_3517,N_3114,N_3160);
xor U3518 (N_3518,N_3016,N_3168);
nor U3519 (N_3519,N_3258,N_3087);
or U3520 (N_3520,N_3100,N_3030);
or U3521 (N_3521,N_3106,N_3084);
or U3522 (N_3522,N_3261,N_3064);
and U3523 (N_3523,N_3166,N_3077);
nand U3524 (N_3524,N_3252,N_3181);
or U3525 (N_3525,N_3292,N_3183);
and U3526 (N_3526,N_3210,N_3038);
xor U3527 (N_3527,N_3133,N_3299);
and U3528 (N_3528,N_3197,N_3233);
nor U3529 (N_3529,N_3084,N_3237);
nand U3530 (N_3530,N_3249,N_3096);
xnor U3531 (N_3531,N_3277,N_3193);
and U3532 (N_3532,N_3185,N_3282);
or U3533 (N_3533,N_3130,N_3125);
nor U3534 (N_3534,N_3030,N_3176);
and U3535 (N_3535,N_3057,N_3031);
or U3536 (N_3536,N_3280,N_3122);
nand U3537 (N_3537,N_3027,N_3255);
xor U3538 (N_3538,N_3188,N_3149);
nand U3539 (N_3539,N_3109,N_3296);
xor U3540 (N_3540,N_3068,N_3072);
and U3541 (N_3541,N_3274,N_3002);
nand U3542 (N_3542,N_3122,N_3017);
nor U3543 (N_3543,N_3255,N_3228);
nand U3544 (N_3544,N_3121,N_3214);
nand U3545 (N_3545,N_3287,N_3243);
nor U3546 (N_3546,N_3172,N_3125);
nand U3547 (N_3547,N_3140,N_3181);
xor U3548 (N_3548,N_3221,N_3194);
or U3549 (N_3549,N_3221,N_3083);
or U3550 (N_3550,N_3234,N_3272);
and U3551 (N_3551,N_3071,N_3077);
nor U3552 (N_3552,N_3058,N_3146);
or U3553 (N_3553,N_3082,N_3127);
nand U3554 (N_3554,N_3267,N_3225);
or U3555 (N_3555,N_3070,N_3160);
nor U3556 (N_3556,N_3261,N_3297);
and U3557 (N_3557,N_3233,N_3214);
nand U3558 (N_3558,N_3224,N_3025);
nor U3559 (N_3559,N_3160,N_3283);
nor U3560 (N_3560,N_3212,N_3015);
nand U3561 (N_3561,N_3110,N_3008);
nor U3562 (N_3562,N_3240,N_3250);
or U3563 (N_3563,N_3209,N_3230);
nor U3564 (N_3564,N_3081,N_3181);
xnor U3565 (N_3565,N_3150,N_3179);
nor U3566 (N_3566,N_3048,N_3214);
and U3567 (N_3567,N_3188,N_3150);
nand U3568 (N_3568,N_3208,N_3160);
nand U3569 (N_3569,N_3183,N_3214);
or U3570 (N_3570,N_3202,N_3133);
xor U3571 (N_3571,N_3119,N_3173);
or U3572 (N_3572,N_3149,N_3017);
xor U3573 (N_3573,N_3037,N_3031);
or U3574 (N_3574,N_3201,N_3124);
xor U3575 (N_3575,N_3215,N_3182);
nand U3576 (N_3576,N_3006,N_3145);
nor U3577 (N_3577,N_3224,N_3108);
and U3578 (N_3578,N_3026,N_3249);
and U3579 (N_3579,N_3125,N_3064);
xor U3580 (N_3580,N_3138,N_3059);
nor U3581 (N_3581,N_3134,N_3256);
nor U3582 (N_3582,N_3200,N_3077);
or U3583 (N_3583,N_3289,N_3053);
nor U3584 (N_3584,N_3167,N_3107);
xnor U3585 (N_3585,N_3254,N_3101);
or U3586 (N_3586,N_3173,N_3246);
or U3587 (N_3587,N_3152,N_3208);
or U3588 (N_3588,N_3269,N_3290);
and U3589 (N_3589,N_3175,N_3266);
nand U3590 (N_3590,N_3097,N_3162);
xor U3591 (N_3591,N_3217,N_3288);
nor U3592 (N_3592,N_3080,N_3079);
or U3593 (N_3593,N_3022,N_3292);
and U3594 (N_3594,N_3227,N_3159);
nor U3595 (N_3595,N_3241,N_3193);
and U3596 (N_3596,N_3161,N_3173);
xnor U3597 (N_3597,N_3215,N_3281);
xor U3598 (N_3598,N_3153,N_3005);
nand U3599 (N_3599,N_3137,N_3004);
and U3600 (N_3600,N_3348,N_3513);
xnor U3601 (N_3601,N_3432,N_3312);
or U3602 (N_3602,N_3526,N_3542);
xnor U3603 (N_3603,N_3480,N_3551);
xnor U3604 (N_3604,N_3326,N_3468);
nor U3605 (N_3605,N_3450,N_3557);
or U3606 (N_3606,N_3584,N_3406);
nor U3607 (N_3607,N_3453,N_3516);
nor U3608 (N_3608,N_3457,N_3420);
and U3609 (N_3609,N_3474,N_3390);
or U3610 (N_3610,N_3395,N_3338);
nor U3611 (N_3611,N_3591,N_3417);
xnor U3612 (N_3612,N_3583,N_3366);
and U3613 (N_3613,N_3456,N_3573);
or U3614 (N_3614,N_3426,N_3484);
and U3615 (N_3615,N_3303,N_3412);
nand U3616 (N_3616,N_3429,N_3349);
xnor U3617 (N_3617,N_3413,N_3428);
and U3618 (N_3618,N_3581,N_3567);
xnor U3619 (N_3619,N_3396,N_3536);
and U3620 (N_3620,N_3388,N_3594);
or U3621 (N_3621,N_3559,N_3404);
and U3622 (N_3622,N_3397,N_3554);
nor U3623 (N_3623,N_3494,N_3552);
nand U3624 (N_3624,N_3441,N_3452);
and U3625 (N_3625,N_3446,N_3501);
or U3626 (N_3626,N_3389,N_3488);
xor U3627 (N_3627,N_3391,N_3300);
xnor U3628 (N_3628,N_3320,N_3469);
xnor U3629 (N_3629,N_3544,N_3586);
nor U3630 (N_3630,N_3534,N_3330);
xor U3631 (N_3631,N_3470,N_3560);
nand U3632 (N_3632,N_3458,N_3409);
and U3633 (N_3633,N_3569,N_3527);
nand U3634 (N_3634,N_3333,N_3346);
and U3635 (N_3635,N_3462,N_3547);
or U3636 (N_3636,N_3443,N_3497);
nand U3637 (N_3637,N_3347,N_3354);
nor U3638 (N_3638,N_3461,N_3363);
nor U3639 (N_3639,N_3493,N_3332);
or U3640 (N_3640,N_3335,N_3570);
xnor U3641 (N_3641,N_3444,N_3435);
xor U3642 (N_3642,N_3492,N_3310);
or U3643 (N_3643,N_3418,N_3599);
and U3644 (N_3644,N_3362,N_3422);
nand U3645 (N_3645,N_3342,N_3355);
nor U3646 (N_3646,N_3485,N_3402);
xnor U3647 (N_3647,N_3509,N_3318);
or U3648 (N_3648,N_3382,N_3510);
nand U3649 (N_3649,N_3368,N_3357);
xnor U3650 (N_3650,N_3356,N_3419);
and U3651 (N_3651,N_3472,N_3481);
and U3652 (N_3652,N_3373,N_3562);
nor U3653 (N_3653,N_3555,N_3520);
nand U3654 (N_3654,N_3378,N_3371);
and U3655 (N_3655,N_3490,N_3425);
xor U3656 (N_3656,N_3370,N_3329);
xnor U3657 (N_3657,N_3538,N_3561);
nor U3658 (N_3658,N_3524,N_3575);
and U3659 (N_3659,N_3314,N_3424);
nor U3660 (N_3660,N_3597,N_3553);
xor U3661 (N_3661,N_3504,N_3578);
or U3662 (N_3662,N_3340,N_3414);
nand U3663 (N_3663,N_3523,N_3433);
or U3664 (N_3664,N_3519,N_3448);
or U3665 (N_3665,N_3336,N_3372);
nand U3666 (N_3666,N_3595,N_3393);
nor U3667 (N_3667,N_3486,N_3352);
nor U3668 (N_3668,N_3339,N_3307);
xnor U3669 (N_3669,N_3565,N_3437);
or U3670 (N_3670,N_3498,N_3459);
or U3671 (N_3671,N_3427,N_3380);
and U3672 (N_3672,N_3589,N_3549);
nor U3673 (N_3673,N_3506,N_3434);
nor U3674 (N_3674,N_3598,N_3574);
nand U3675 (N_3675,N_3582,N_3539);
xor U3676 (N_3676,N_3491,N_3487);
nor U3677 (N_3677,N_3405,N_3464);
nand U3678 (N_3678,N_3367,N_3325);
nand U3679 (N_3679,N_3479,N_3596);
nand U3680 (N_3680,N_3416,N_3499);
xor U3681 (N_3681,N_3571,N_3358);
and U3682 (N_3682,N_3337,N_3535);
or U3683 (N_3683,N_3563,N_3411);
and U3684 (N_3684,N_3546,N_3541);
xor U3685 (N_3685,N_3530,N_3502);
and U3686 (N_3686,N_3521,N_3556);
nand U3687 (N_3687,N_3386,N_3564);
xnor U3688 (N_3688,N_3537,N_3445);
xnor U3689 (N_3689,N_3496,N_3345);
nor U3690 (N_3690,N_3592,N_3309);
nand U3691 (N_3691,N_3507,N_3588);
nand U3692 (N_3692,N_3447,N_3317);
or U3693 (N_3693,N_3381,N_3467);
or U3694 (N_3694,N_3532,N_3403);
or U3695 (N_3695,N_3315,N_3511);
nand U3696 (N_3696,N_3376,N_3415);
and U3697 (N_3697,N_3387,N_3301);
nor U3698 (N_3698,N_3438,N_3517);
nand U3699 (N_3699,N_3306,N_3465);
and U3700 (N_3700,N_3334,N_3383);
nor U3701 (N_3701,N_3473,N_3369);
or U3702 (N_3702,N_3305,N_3400);
and U3703 (N_3703,N_3328,N_3364);
nor U3704 (N_3704,N_3533,N_3385);
and U3705 (N_3705,N_3550,N_3455);
nand U3706 (N_3706,N_3477,N_3440);
and U3707 (N_3707,N_3577,N_3407);
nor U3708 (N_3708,N_3505,N_3319);
nor U3709 (N_3709,N_3394,N_3558);
xnor U3710 (N_3710,N_3331,N_3344);
and U3711 (N_3711,N_3360,N_3466);
or U3712 (N_3712,N_3460,N_3398);
nor U3713 (N_3713,N_3476,N_3327);
nand U3714 (N_3714,N_3436,N_3500);
nor U3715 (N_3715,N_3442,N_3515);
nor U3716 (N_3716,N_3311,N_3304);
nand U3717 (N_3717,N_3463,N_3316);
and U3718 (N_3718,N_3324,N_3529);
xor U3719 (N_3719,N_3580,N_3430);
or U3720 (N_3720,N_3401,N_3540);
and U3721 (N_3721,N_3384,N_3590);
xnor U3722 (N_3722,N_3478,N_3514);
or U3723 (N_3723,N_3341,N_3375);
and U3724 (N_3724,N_3566,N_3359);
and U3725 (N_3725,N_3374,N_3323);
nor U3726 (N_3726,N_3587,N_3343);
or U3727 (N_3727,N_3392,N_3576);
or U3728 (N_3728,N_3512,N_3379);
nand U3729 (N_3729,N_3483,N_3454);
and U3730 (N_3730,N_3365,N_3350);
xor U3731 (N_3731,N_3545,N_3451);
and U3732 (N_3732,N_3439,N_3399);
or U3733 (N_3733,N_3593,N_3353);
or U3734 (N_3734,N_3489,N_3322);
xnor U3735 (N_3735,N_3531,N_3508);
xor U3736 (N_3736,N_3475,N_3568);
and U3737 (N_3737,N_3377,N_3308);
xnor U3738 (N_3738,N_3361,N_3525);
or U3739 (N_3739,N_3313,N_3410);
and U3740 (N_3740,N_3302,N_3522);
xnor U3741 (N_3741,N_3421,N_3528);
or U3742 (N_3742,N_3431,N_3518);
xor U3743 (N_3743,N_3585,N_3449);
xnor U3744 (N_3744,N_3503,N_3572);
xnor U3745 (N_3745,N_3548,N_3579);
or U3746 (N_3746,N_3351,N_3471);
and U3747 (N_3747,N_3482,N_3321);
nor U3748 (N_3748,N_3543,N_3495);
nor U3749 (N_3749,N_3408,N_3423);
xor U3750 (N_3750,N_3360,N_3425);
and U3751 (N_3751,N_3350,N_3492);
xnor U3752 (N_3752,N_3312,N_3534);
nor U3753 (N_3753,N_3367,N_3448);
xnor U3754 (N_3754,N_3306,N_3535);
or U3755 (N_3755,N_3492,N_3388);
nand U3756 (N_3756,N_3577,N_3511);
nor U3757 (N_3757,N_3466,N_3471);
or U3758 (N_3758,N_3406,N_3363);
nor U3759 (N_3759,N_3569,N_3387);
xor U3760 (N_3760,N_3364,N_3487);
nand U3761 (N_3761,N_3572,N_3334);
and U3762 (N_3762,N_3597,N_3414);
nand U3763 (N_3763,N_3309,N_3557);
or U3764 (N_3764,N_3593,N_3496);
or U3765 (N_3765,N_3506,N_3406);
and U3766 (N_3766,N_3533,N_3396);
or U3767 (N_3767,N_3366,N_3321);
nand U3768 (N_3768,N_3318,N_3536);
xnor U3769 (N_3769,N_3551,N_3581);
and U3770 (N_3770,N_3578,N_3329);
or U3771 (N_3771,N_3409,N_3511);
nand U3772 (N_3772,N_3413,N_3523);
or U3773 (N_3773,N_3456,N_3361);
and U3774 (N_3774,N_3436,N_3517);
and U3775 (N_3775,N_3456,N_3551);
or U3776 (N_3776,N_3362,N_3304);
xnor U3777 (N_3777,N_3505,N_3438);
nor U3778 (N_3778,N_3348,N_3469);
or U3779 (N_3779,N_3394,N_3425);
nand U3780 (N_3780,N_3583,N_3478);
and U3781 (N_3781,N_3470,N_3305);
nand U3782 (N_3782,N_3451,N_3596);
and U3783 (N_3783,N_3546,N_3512);
or U3784 (N_3784,N_3508,N_3498);
and U3785 (N_3785,N_3342,N_3300);
xor U3786 (N_3786,N_3379,N_3346);
nand U3787 (N_3787,N_3599,N_3535);
and U3788 (N_3788,N_3381,N_3435);
and U3789 (N_3789,N_3506,N_3483);
or U3790 (N_3790,N_3316,N_3303);
or U3791 (N_3791,N_3561,N_3364);
nor U3792 (N_3792,N_3355,N_3337);
and U3793 (N_3793,N_3448,N_3535);
nand U3794 (N_3794,N_3324,N_3474);
xnor U3795 (N_3795,N_3434,N_3547);
nor U3796 (N_3796,N_3424,N_3336);
or U3797 (N_3797,N_3332,N_3436);
nor U3798 (N_3798,N_3362,N_3312);
nor U3799 (N_3799,N_3412,N_3589);
and U3800 (N_3800,N_3519,N_3403);
or U3801 (N_3801,N_3545,N_3428);
nor U3802 (N_3802,N_3501,N_3562);
or U3803 (N_3803,N_3347,N_3361);
nand U3804 (N_3804,N_3476,N_3382);
xor U3805 (N_3805,N_3489,N_3379);
nor U3806 (N_3806,N_3426,N_3445);
or U3807 (N_3807,N_3499,N_3481);
nand U3808 (N_3808,N_3342,N_3380);
nand U3809 (N_3809,N_3536,N_3526);
nand U3810 (N_3810,N_3370,N_3339);
and U3811 (N_3811,N_3568,N_3590);
or U3812 (N_3812,N_3429,N_3398);
and U3813 (N_3813,N_3381,N_3408);
xor U3814 (N_3814,N_3586,N_3553);
or U3815 (N_3815,N_3546,N_3410);
nand U3816 (N_3816,N_3595,N_3366);
and U3817 (N_3817,N_3302,N_3555);
or U3818 (N_3818,N_3378,N_3459);
and U3819 (N_3819,N_3418,N_3504);
or U3820 (N_3820,N_3457,N_3384);
and U3821 (N_3821,N_3393,N_3564);
nor U3822 (N_3822,N_3396,N_3576);
nand U3823 (N_3823,N_3321,N_3417);
nand U3824 (N_3824,N_3540,N_3321);
nor U3825 (N_3825,N_3543,N_3317);
and U3826 (N_3826,N_3391,N_3324);
xor U3827 (N_3827,N_3379,N_3372);
nand U3828 (N_3828,N_3392,N_3417);
nand U3829 (N_3829,N_3393,N_3356);
and U3830 (N_3830,N_3445,N_3397);
and U3831 (N_3831,N_3332,N_3489);
nand U3832 (N_3832,N_3412,N_3433);
nand U3833 (N_3833,N_3428,N_3530);
xor U3834 (N_3834,N_3483,N_3381);
and U3835 (N_3835,N_3371,N_3427);
nor U3836 (N_3836,N_3516,N_3564);
nor U3837 (N_3837,N_3397,N_3436);
nor U3838 (N_3838,N_3513,N_3576);
nor U3839 (N_3839,N_3485,N_3300);
nand U3840 (N_3840,N_3484,N_3456);
nand U3841 (N_3841,N_3306,N_3444);
or U3842 (N_3842,N_3301,N_3425);
and U3843 (N_3843,N_3346,N_3308);
xnor U3844 (N_3844,N_3341,N_3533);
or U3845 (N_3845,N_3439,N_3588);
nor U3846 (N_3846,N_3307,N_3341);
or U3847 (N_3847,N_3560,N_3400);
nor U3848 (N_3848,N_3496,N_3327);
and U3849 (N_3849,N_3520,N_3560);
and U3850 (N_3850,N_3543,N_3517);
and U3851 (N_3851,N_3330,N_3418);
and U3852 (N_3852,N_3497,N_3598);
xnor U3853 (N_3853,N_3586,N_3580);
nand U3854 (N_3854,N_3540,N_3579);
nand U3855 (N_3855,N_3358,N_3543);
nor U3856 (N_3856,N_3511,N_3379);
nor U3857 (N_3857,N_3328,N_3365);
or U3858 (N_3858,N_3355,N_3550);
or U3859 (N_3859,N_3334,N_3491);
nand U3860 (N_3860,N_3392,N_3473);
nor U3861 (N_3861,N_3420,N_3482);
nand U3862 (N_3862,N_3544,N_3519);
and U3863 (N_3863,N_3320,N_3523);
and U3864 (N_3864,N_3341,N_3528);
xnor U3865 (N_3865,N_3357,N_3367);
xor U3866 (N_3866,N_3580,N_3332);
nor U3867 (N_3867,N_3554,N_3358);
or U3868 (N_3868,N_3592,N_3507);
nor U3869 (N_3869,N_3487,N_3328);
and U3870 (N_3870,N_3554,N_3475);
or U3871 (N_3871,N_3447,N_3507);
or U3872 (N_3872,N_3474,N_3343);
nor U3873 (N_3873,N_3355,N_3349);
xnor U3874 (N_3874,N_3359,N_3482);
nor U3875 (N_3875,N_3468,N_3418);
nor U3876 (N_3876,N_3404,N_3487);
or U3877 (N_3877,N_3469,N_3495);
xor U3878 (N_3878,N_3300,N_3558);
nand U3879 (N_3879,N_3348,N_3420);
xnor U3880 (N_3880,N_3532,N_3322);
xnor U3881 (N_3881,N_3359,N_3497);
or U3882 (N_3882,N_3533,N_3380);
nor U3883 (N_3883,N_3365,N_3370);
nor U3884 (N_3884,N_3434,N_3376);
nand U3885 (N_3885,N_3349,N_3379);
or U3886 (N_3886,N_3432,N_3499);
xor U3887 (N_3887,N_3315,N_3543);
xor U3888 (N_3888,N_3426,N_3541);
or U3889 (N_3889,N_3425,N_3474);
and U3890 (N_3890,N_3318,N_3516);
and U3891 (N_3891,N_3599,N_3404);
nor U3892 (N_3892,N_3536,N_3326);
and U3893 (N_3893,N_3518,N_3389);
or U3894 (N_3894,N_3437,N_3456);
or U3895 (N_3895,N_3468,N_3580);
nor U3896 (N_3896,N_3548,N_3417);
or U3897 (N_3897,N_3534,N_3439);
nand U3898 (N_3898,N_3375,N_3333);
nor U3899 (N_3899,N_3340,N_3334);
or U3900 (N_3900,N_3868,N_3842);
or U3901 (N_3901,N_3692,N_3671);
or U3902 (N_3902,N_3602,N_3849);
xor U3903 (N_3903,N_3624,N_3614);
nand U3904 (N_3904,N_3850,N_3699);
and U3905 (N_3905,N_3672,N_3688);
and U3906 (N_3906,N_3799,N_3822);
nor U3907 (N_3907,N_3656,N_3690);
nand U3908 (N_3908,N_3859,N_3724);
and U3909 (N_3909,N_3616,N_3860);
xor U3910 (N_3910,N_3797,N_3780);
xnor U3911 (N_3911,N_3705,N_3856);
and U3912 (N_3912,N_3711,N_3834);
xor U3913 (N_3913,N_3631,N_3652);
nor U3914 (N_3914,N_3871,N_3740);
xnor U3915 (N_3915,N_3792,N_3710);
and U3916 (N_3916,N_3835,N_3865);
or U3917 (N_3917,N_3864,N_3702);
and U3918 (N_3918,N_3653,N_3726);
and U3919 (N_3919,N_3613,N_3720);
nor U3920 (N_3920,N_3679,N_3661);
nand U3921 (N_3921,N_3722,N_3638);
or U3922 (N_3922,N_3814,N_3879);
or U3923 (N_3923,N_3843,N_3839);
and U3924 (N_3924,N_3853,N_3830);
nand U3925 (N_3925,N_3791,N_3649);
or U3926 (N_3926,N_3645,N_3881);
or U3927 (N_3927,N_3776,N_3886);
and U3928 (N_3928,N_3811,N_3634);
nor U3929 (N_3929,N_3793,N_3732);
nor U3930 (N_3930,N_3681,N_3659);
xor U3931 (N_3931,N_3801,N_3765);
xnor U3932 (N_3932,N_3889,N_3749);
xor U3933 (N_3933,N_3821,N_3862);
xnor U3934 (N_3934,N_3618,N_3639);
and U3935 (N_3935,N_3844,N_3771);
nor U3936 (N_3936,N_3826,N_3683);
nor U3937 (N_3937,N_3769,N_3617);
xor U3938 (N_3938,N_3640,N_3609);
or U3939 (N_3939,N_3697,N_3633);
xnor U3940 (N_3940,N_3636,N_3685);
or U3941 (N_3941,N_3810,N_3861);
xnor U3942 (N_3942,N_3838,N_3777);
nand U3943 (N_3943,N_3745,N_3763);
and U3944 (N_3944,N_3682,N_3759);
and U3945 (N_3945,N_3727,N_3802);
nor U3946 (N_3946,N_3737,N_3878);
nor U3947 (N_3947,N_3698,N_3798);
or U3948 (N_3948,N_3746,N_3619);
nand U3949 (N_3949,N_3731,N_3678);
nor U3950 (N_3950,N_3627,N_3800);
and U3951 (N_3951,N_3758,N_3611);
nor U3952 (N_3952,N_3806,N_3808);
nand U3953 (N_3953,N_3620,N_3686);
or U3954 (N_3954,N_3774,N_3600);
xor U3955 (N_3955,N_3676,N_3657);
and U3956 (N_3956,N_3701,N_3827);
or U3957 (N_3957,N_3654,N_3812);
nand U3958 (N_3958,N_3695,N_3641);
and U3959 (N_3959,N_3768,N_3742);
nor U3960 (N_3960,N_3615,N_3887);
nand U3961 (N_3961,N_3757,N_3779);
or U3962 (N_3962,N_3610,N_3706);
and U3963 (N_3963,N_3719,N_3845);
nor U3964 (N_3964,N_3635,N_3770);
nand U3965 (N_3965,N_3736,N_3663);
and U3966 (N_3966,N_3718,N_3787);
nand U3967 (N_3967,N_3693,N_3760);
or U3968 (N_3968,N_3781,N_3899);
or U3969 (N_3969,N_3622,N_3747);
xnor U3970 (N_3970,N_3788,N_3607);
and U3971 (N_3971,N_3825,N_3873);
nor U3972 (N_3972,N_3863,N_3643);
nand U3973 (N_3973,N_3738,N_3890);
or U3974 (N_3974,N_3896,N_3809);
or U3975 (N_3975,N_3744,N_3729);
nor U3976 (N_3976,N_3828,N_3601);
nor U3977 (N_3977,N_3813,N_3847);
and U3978 (N_3978,N_3832,N_3794);
nor U3979 (N_3979,N_3755,N_3716);
or U3980 (N_3980,N_3816,N_3664);
nor U3981 (N_3981,N_3851,N_3725);
nand U3982 (N_3982,N_3767,N_3668);
nor U3983 (N_3983,N_3642,N_3867);
xor U3984 (N_3984,N_3628,N_3795);
nand U3985 (N_3985,N_3677,N_3876);
and U3986 (N_3986,N_3888,N_3665);
nand U3987 (N_3987,N_3714,N_3773);
xnor U3988 (N_3988,N_3625,N_3629);
and U3989 (N_3989,N_3778,N_3761);
and U3990 (N_3990,N_3687,N_3623);
nor U3991 (N_3991,N_3723,N_3784);
or U3992 (N_3992,N_3658,N_3833);
or U3993 (N_3993,N_3632,N_3892);
xor U3994 (N_3994,N_3750,N_3855);
nand U3995 (N_3995,N_3852,N_3637);
and U3996 (N_3996,N_3841,N_3789);
nor U3997 (N_3997,N_3782,N_3748);
and U3998 (N_3998,N_3675,N_3805);
or U3999 (N_3999,N_3829,N_3817);
and U4000 (N_4000,N_3605,N_3612);
nand U4001 (N_4001,N_3877,N_3894);
and U4002 (N_4002,N_3669,N_3846);
xnor U4003 (N_4003,N_3824,N_3647);
nand U4004 (N_4004,N_3870,N_3854);
xor U4005 (N_4005,N_3733,N_3786);
nor U4006 (N_4006,N_3836,N_3662);
xnor U4007 (N_4007,N_3709,N_3772);
xnor U4008 (N_4008,N_3882,N_3753);
xnor U4009 (N_4009,N_3898,N_3650);
and U4010 (N_4010,N_3707,N_3885);
or U4011 (N_4011,N_3604,N_3869);
nor U4012 (N_4012,N_3673,N_3752);
nand U4013 (N_4013,N_3803,N_3655);
nand U4014 (N_4014,N_3762,N_3626);
nand U4015 (N_4015,N_3840,N_3880);
and U4016 (N_4016,N_3646,N_3667);
or U4017 (N_4017,N_3735,N_3754);
nor U4018 (N_4018,N_3857,N_3666);
nor U4019 (N_4019,N_3730,N_3712);
nand U4020 (N_4020,N_3734,N_3608);
and U4021 (N_4021,N_3815,N_3775);
xnor U4022 (N_4022,N_3874,N_3895);
or U4023 (N_4023,N_3603,N_3721);
or U4024 (N_4024,N_3848,N_3713);
xor U4025 (N_4025,N_3872,N_3891);
or U4026 (N_4026,N_3837,N_3621);
and U4027 (N_4027,N_3796,N_3700);
nand U4028 (N_4028,N_3807,N_3790);
nand U4029 (N_4029,N_3875,N_3648);
xnor U4030 (N_4030,N_3893,N_3743);
and U4031 (N_4031,N_3751,N_3897);
and U4032 (N_4032,N_3820,N_3674);
and U4033 (N_4033,N_3858,N_3670);
and U4034 (N_4034,N_3818,N_3883);
nor U4035 (N_4035,N_3819,N_3630);
or U4036 (N_4036,N_3606,N_3660);
nor U4037 (N_4037,N_3785,N_3703);
and U4038 (N_4038,N_3741,N_3766);
nor U4039 (N_4039,N_3696,N_3756);
nor U4040 (N_4040,N_3764,N_3684);
xor U4041 (N_4041,N_3831,N_3717);
nand U4042 (N_4042,N_3715,N_3804);
nor U4043 (N_4043,N_3728,N_3691);
nor U4044 (N_4044,N_3644,N_3739);
and U4045 (N_4045,N_3708,N_3884);
nor U4046 (N_4046,N_3651,N_3689);
or U4047 (N_4047,N_3866,N_3783);
nor U4048 (N_4048,N_3704,N_3680);
and U4049 (N_4049,N_3694,N_3823);
or U4050 (N_4050,N_3743,N_3878);
or U4051 (N_4051,N_3855,N_3663);
nand U4052 (N_4052,N_3879,N_3638);
nand U4053 (N_4053,N_3841,N_3727);
nor U4054 (N_4054,N_3734,N_3644);
or U4055 (N_4055,N_3723,N_3836);
or U4056 (N_4056,N_3816,N_3724);
xor U4057 (N_4057,N_3644,N_3874);
nand U4058 (N_4058,N_3753,N_3744);
nor U4059 (N_4059,N_3882,N_3788);
xnor U4060 (N_4060,N_3891,N_3879);
and U4061 (N_4061,N_3856,N_3776);
nor U4062 (N_4062,N_3756,N_3881);
xor U4063 (N_4063,N_3600,N_3768);
or U4064 (N_4064,N_3857,N_3687);
nand U4065 (N_4065,N_3681,N_3800);
nand U4066 (N_4066,N_3778,N_3730);
and U4067 (N_4067,N_3830,N_3832);
xor U4068 (N_4068,N_3840,N_3609);
nand U4069 (N_4069,N_3706,N_3877);
nand U4070 (N_4070,N_3760,N_3711);
xor U4071 (N_4071,N_3693,N_3861);
nor U4072 (N_4072,N_3651,N_3852);
and U4073 (N_4073,N_3736,N_3831);
and U4074 (N_4074,N_3643,N_3635);
or U4075 (N_4075,N_3826,N_3616);
nand U4076 (N_4076,N_3835,N_3651);
or U4077 (N_4077,N_3642,N_3707);
xnor U4078 (N_4078,N_3820,N_3631);
nand U4079 (N_4079,N_3614,N_3866);
nand U4080 (N_4080,N_3863,N_3740);
or U4081 (N_4081,N_3642,N_3664);
or U4082 (N_4082,N_3736,N_3725);
nor U4083 (N_4083,N_3830,N_3601);
and U4084 (N_4084,N_3829,N_3893);
nor U4085 (N_4085,N_3663,N_3786);
and U4086 (N_4086,N_3700,N_3838);
nor U4087 (N_4087,N_3847,N_3668);
nand U4088 (N_4088,N_3876,N_3644);
and U4089 (N_4089,N_3763,N_3653);
nor U4090 (N_4090,N_3662,N_3877);
or U4091 (N_4091,N_3648,N_3887);
nand U4092 (N_4092,N_3627,N_3805);
xor U4093 (N_4093,N_3897,N_3763);
nand U4094 (N_4094,N_3853,N_3603);
xor U4095 (N_4095,N_3629,N_3806);
or U4096 (N_4096,N_3763,N_3605);
nand U4097 (N_4097,N_3623,N_3821);
nand U4098 (N_4098,N_3774,N_3623);
xnor U4099 (N_4099,N_3649,N_3608);
nor U4100 (N_4100,N_3601,N_3845);
xor U4101 (N_4101,N_3845,N_3604);
or U4102 (N_4102,N_3772,N_3615);
nor U4103 (N_4103,N_3725,N_3621);
or U4104 (N_4104,N_3824,N_3646);
xnor U4105 (N_4105,N_3826,N_3781);
nand U4106 (N_4106,N_3865,N_3665);
and U4107 (N_4107,N_3620,N_3800);
nand U4108 (N_4108,N_3653,N_3715);
nand U4109 (N_4109,N_3687,N_3660);
nand U4110 (N_4110,N_3863,N_3864);
or U4111 (N_4111,N_3894,N_3742);
nor U4112 (N_4112,N_3657,N_3739);
nand U4113 (N_4113,N_3851,N_3793);
xnor U4114 (N_4114,N_3620,N_3718);
nand U4115 (N_4115,N_3667,N_3601);
xor U4116 (N_4116,N_3899,N_3651);
nor U4117 (N_4117,N_3792,N_3791);
and U4118 (N_4118,N_3670,N_3743);
or U4119 (N_4119,N_3649,N_3800);
and U4120 (N_4120,N_3851,N_3741);
nor U4121 (N_4121,N_3847,N_3671);
nor U4122 (N_4122,N_3709,N_3634);
or U4123 (N_4123,N_3864,N_3743);
xor U4124 (N_4124,N_3865,N_3622);
or U4125 (N_4125,N_3743,N_3728);
xnor U4126 (N_4126,N_3789,N_3838);
nand U4127 (N_4127,N_3806,N_3628);
or U4128 (N_4128,N_3708,N_3628);
nor U4129 (N_4129,N_3608,N_3775);
or U4130 (N_4130,N_3685,N_3868);
and U4131 (N_4131,N_3613,N_3891);
nor U4132 (N_4132,N_3824,N_3808);
nand U4133 (N_4133,N_3848,N_3899);
nor U4134 (N_4134,N_3839,N_3713);
nor U4135 (N_4135,N_3734,N_3609);
and U4136 (N_4136,N_3613,N_3699);
and U4137 (N_4137,N_3628,N_3650);
and U4138 (N_4138,N_3756,N_3629);
nand U4139 (N_4139,N_3760,N_3817);
nand U4140 (N_4140,N_3742,N_3761);
and U4141 (N_4141,N_3673,N_3625);
nor U4142 (N_4142,N_3668,N_3830);
xnor U4143 (N_4143,N_3803,N_3715);
nor U4144 (N_4144,N_3623,N_3750);
and U4145 (N_4145,N_3631,N_3601);
or U4146 (N_4146,N_3854,N_3711);
and U4147 (N_4147,N_3796,N_3696);
and U4148 (N_4148,N_3796,N_3806);
xnor U4149 (N_4149,N_3716,N_3659);
and U4150 (N_4150,N_3796,N_3642);
nand U4151 (N_4151,N_3840,N_3628);
nand U4152 (N_4152,N_3784,N_3718);
nand U4153 (N_4153,N_3796,N_3729);
nand U4154 (N_4154,N_3613,N_3853);
or U4155 (N_4155,N_3863,N_3812);
xor U4156 (N_4156,N_3754,N_3732);
or U4157 (N_4157,N_3698,N_3761);
nor U4158 (N_4158,N_3687,N_3776);
nand U4159 (N_4159,N_3641,N_3629);
and U4160 (N_4160,N_3843,N_3600);
nand U4161 (N_4161,N_3839,N_3674);
or U4162 (N_4162,N_3725,N_3756);
and U4163 (N_4163,N_3890,N_3837);
nor U4164 (N_4164,N_3767,N_3632);
or U4165 (N_4165,N_3833,N_3698);
xnor U4166 (N_4166,N_3878,N_3769);
nand U4167 (N_4167,N_3715,N_3670);
nor U4168 (N_4168,N_3847,N_3610);
nand U4169 (N_4169,N_3882,N_3874);
and U4170 (N_4170,N_3705,N_3762);
xor U4171 (N_4171,N_3619,N_3675);
xnor U4172 (N_4172,N_3888,N_3628);
and U4173 (N_4173,N_3793,N_3854);
nand U4174 (N_4174,N_3660,N_3727);
xor U4175 (N_4175,N_3646,N_3715);
nand U4176 (N_4176,N_3705,N_3788);
nand U4177 (N_4177,N_3885,N_3847);
nand U4178 (N_4178,N_3870,N_3864);
and U4179 (N_4179,N_3604,N_3723);
and U4180 (N_4180,N_3809,N_3801);
and U4181 (N_4181,N_3780,N_3796);
xor U4182 (N_4182,N_3681,N_3656);
or U4183 (N_4183,N_3667,N_3754);
and U4184 (N_4184,N_3688,N_3637);
xnor U4185 (N_4185,N_3601,N_3651);
xnor U4186 (N_4186,N_3786,N_3824);
nor U4187 (N_4187,N_3793,N_3739);
nor U4188 (N_4188,N_3843,N_3624);
or U4189 (N_4189,N_3606,N_3719);
and U4190 (N_4190,N_3677,N_3815);
or U4191 (N_4191,N_3641,N_3643);
and U4192 (N_4192,N_3827,N_3841);
and U4193 (N_4193,N_3892,N_3857);
nand U4194 (N_4194,N_3615,N_3844);
xnor U4195 (N_4195,N_3609,N_3732);
and U4196 (N_4196,N_3625,N_3805);
xnor U4197 (N_4197,N_3743,N_3799);
or U4198 (N_4198,N_3719,N_3757);
and U4199 (N_4199,N_3780,N_3807);
or U4200 (N_4200,N_4123,N_4158);
nand U4201 (N_4201,N_4180,N_4010);
and U4202 (N_4202,N_4048,N_3940);
or U4203 (N_4203,N_4138,N_4162);
xnor U4204 (N_4204,N_3944,N_3929);
xor U4205 (N_4205,N_4141,N_3996);
xor U4206 (N_4206,N_4095,N_4065);
and U4207 (N_4207,N_4110,N_4003);
and U4208 (N_4208,N_4001,N_3921);
or U4209 (N_4209,N_4017,N_4081);
nor U4210 (N_4210,N_4056,N_3915);
nor U4211 (N_4211,N_4076,N_4103);
nor U4212 (N_4212,N_4027,N_3965);
xor U4213 (N_4213,N_4169,N_4052);
xnor U4214 (N_4214,N_4070,N_4038);
or U4215 (N_4215,N_3906,N_3982);
and U4216 (N_4216,N_3989,N_4140);
and U4217 (N_4217,N_4080,N_4178);
and U4218 (N_4218,N_4090,N_4062);
or U4219 (N_4219,N_4088,N_4036);
or U4220 (N_4220,N_4008,N_4196);
and U4221 (N_4221,N_4152,N_3936);
nor U4222 (N_4222,N_4054,N_4114);
or U4223 (N_4223,N_3995,N_4113);
xor U4224 (N_4224,N_4142,N_4105);
nor U4225 (N_4225,N_3903,N_4031);
and U4226 (N_4226,N_4032,N_4084);
nor U4227 (N_4227,N_3961,N_4013);
or U4228 (N_4228,N_4074,N_3960);
nand U4229 (N_4229,N_4148,N_4073);
nor U4230 (N_4230,N_4184,N_3981);
nor U4231 (N_4231,N_3992,N_3938);
xor U4232 (N_4232,N_4028,N_3931);
nor U4233 (N_4233,N_4185,N_4000);
nor U4234 (N_4234,N_4072,N_3914);
or U4235 (N_4235,N_4015,N_4101);
nand U4236 (N_4236,N_3972,N_4099);
and U4237 (N_4237,N_4174,N_3946);
nand U4238 (N_4238,N_4045,N_4087);
and U4239 (N_4239,N_4006,N_4033);
xor U4240 (N_4240,N_4191,N_4153);
nand U4241 (N_4241,N_3980,N_4047);
xnor U4242 (N_4242,N_3937,N_4069);
nand U4243 (N_4243,N_4107,N_3985);
xor U4244 (N_4244,N_4195,N_3966);
nor U4245 (N_4245,N_3999,N_3924);
and U4246 (N_4246,N_4130,N_4179);
or U4247 (N_4247,N_3911,N_4112);
or U4248 (N_4248,N_4023,N_4135);
or U4249 (N_4249,N_3964,N_4150);
xor U4250 (N_4250,N_3956,N_4083);
or U4251 (N_4251,N_4139,N_3950);
and U4252 (N_4252,N_4005,N_3920);
xor U4253 (N_4253,N_3913,N_3998);
nand U4254 (N_4254,N_3919,N_4146);
nor U4255 (N_4255,N_3932,N_4068);
or U4256 (N_4256,N_4137,N_4024);
or U4257 (N_4257,N_3917,N_4098);
nor U4258 (N_4258,N_4154,N_4044);
and U4259 (N_4259,N_4159,N_3904);
xnor U4260 (N_4260,N_4160,N_4041);
nor U4261 (N_4261,N_4089,N_3976);
nand U4262 (N_4262,N_4051,N_3947);
and U4263 (N_4263,N_4168,N_3916);
nand U4264 (N_4264,N_4119,N_4022);
or U4265 (N_4265,N_4149,N_4131);
nand U4266 (N_4266,N_3987,N_3900);
and U4267 (N_4267,N_4172,N_4190);
or U4268 (N_4268,N_3948,N_4144);
or U4269 (N_4269,N_4034,N_4011);
and U4270 (N_4270,N_3934,N_3952);
xnor U4271 (N_4271,N_4166,N_4170);
xor U4272 (N_4272,N_4189,N_4025);
and U4273 (N_4273,N_4116,N_3984);
or U4274 (N_4274,N_3926,N_4177);
or U4275 (N_4275,N_4155,N_3977);
nor U4276 (N_4276,N_4053,N_4058);
nor U4277 (N_4277,N_4121,N_4128);
nor U4278 (N_4278,N_4111,N_4082);
xnor U4279 (N_4279,N_4043,N_4094);
xnor U4280 (N_4280,N_4157,N_4163);
nand U4281 (N_4281,N_4040,N_3907);
and U4282 (N_4282,N_3993,N_4050);
and U4283 (N_4283,N_3951,N_4039);
and U4284 (N_4284,N_4061,N_3986);
or U4285 (N_4285,N_4183,N_4042);
and U4286 (N_4286,N_4018,N_3971);
or U4287 (N_4287,N_4020,N_4132);
xnor U4288 (N_4288,N_4085,N_3963);
nor U4289 (N_4289,N_4091,N_4182);
nand U4290 (N_4290,N_4037,N_3909);
and U4291 (N_4291,N_4127,N_4125);
or U4292 (N_4292,N_3988,N_4117);
nor U4293 (N_4293,N_4064,N_3910);
and U4294 (N_4294,N_4165,N_3930);
or U4295 (N_4295,N_4021,N_3959);
xnor U4296 (N_4296,N_4104,N_4106);
and U4297 (N_4297,N_4057,N_4115);
xnor U4298 (N_4298,N_4029,N_4133);
and U4299 (N_4299,N_3974,N_4046);
and U4300 (N_4300,N_3983,N_4067);
xnor U4301 (N_4301,N_4109,N_4147);
nand U4302 (N_4302,N_4030,N_4071);
or U4303 (N_4303,N_3949,N_3905);
and U4304 (N_4304,N_4171,N_4019);
or U4305 (N_4305,N_3954,N_4016);
and U4306 (N_4306,N_3945,N_4134);
nor U4307 (N_4307,N_4164,N_4145);
nand U4308 (N_4308,N_3962,N_4012);
or U4309 (N_4309,N_4055,N_4060);
nand U4310 (N_4310,N_4188,N_4059);
xor U4311 (N_4311,N_4187,N_4175);
nand U4312 (N_4312,N_4193,N_4118);
or U4313 (N_4313,N_3969,N_4122);
nand U4314 (N_4314,N_4100,N_4136);
or U4315 (N_4315,N_4096,N_4126);
xnor U4316 (N_4316,N_3997,N_3955);
or U4317 (N_4317,N_4092,N_4066);
and U4318 (N_4318,N_4192,N_3943);
and U4319 (N_4319,N_3975,N_3991);
and U4320 (N_4320,N_4097,N_3933);
or U4321 (N_4321,N_3953,N_4026);
and U4322 (N_4322,N_3958,N_3902);
and U4323 (N_4323,N_4161,N_4198);
and U4324 (N_4324,N_3941,N_4077);
nor U4325 (N_4325,N_3925,N_4129);
or U4326 (N_4326,N_4194,N_4014);
nand U4327 (N_4327,N_3942,N_3901);
nor U4328 (N_4328,N_4186,N_4004);
or U4329 (N_4329,N_3908,N_4007);
nor U4330 (N_4330,N_3923,N_4124);
nand U4331 (N_4331,N_4151,N_3935);
nand U4332 (N_4332,N_3922,N_3967);
nand U4333 (N_4333,N_3918,N_4078);
and U4334 (N_4334,N_4197,N_4143);
nand U4335 (N_4335,N_3928,N_4173);
and U4336 (N_4336,N_4108,N_4063);
nand U4337 (N_4337,N_3968,N_4102);
xnor U4338 (N_4338,N_3970,N_3973);
xor U4339 (N_4339,N_4093,N_4167);
xor U4340 (N_4340,N_3912,N_3978);
and U4341 (N_4341,N_4156,N_4176);
and U4342 (N_4342,N_3939,N_4009);
nor U4343 (N_4343,N_3927,N_3957);
and U4344 (N_4344,N_3990,N_4120);
or U4345 (N_4345,N_4079,N_3994);
nand U4346 (N_4346,N_4049,N_4181);
xnor U4347 (N_4347,N_4075,N_4199);
xor U4348 (N_4348,N_3979,N_4086);
and U4349 (N_4349,N_4035,N_4002);
nor U4350 (N_4350,N_3945,N_4034);
nand U4351 (N_4351,N_4109,N_4185);
and U4352 (N_4352,N_3916,N_3955);
nor U4353 (N_4353,N_4185,N_4148);
and U4354 (N_4354,N_3955,N_4142);
nor U4355 (N_4355,N_4018,N_3936);
nand U4356 (N_4356,N_4140,N_3961);
nor U4357 (N_4357,N_4167,N_4052);
or U4358 (N_4358,N_4052,N_4152);
or U4359 (N_4359,N_4000,N_3903);
nor U4360 (N_4360,N_4053,N_4147);
nand U4361 (N_4361,N_4186,N_4164);
xnor U4362 (N_4362,N_4028,N_4111);
nand U4363 (N_4363,N_3987,N_3947);
and U4364 (N_4364,N_4117,N_4095);
or U4365 (N_4365,N_3938,N_4106);
or U4366 (N_4366,N_4162,N_4003);
nand U4367 (N_4367,N_3936,N_3980);
and U4368 (N_4368,N_3971,N_4082);
nor U4369 (N_4369,N_4115,N_4082);
or U4370 (N_4370,N_4035,N_4187);
nor U4371 (N_4371,N_4129,N_4151);
nand U4372 (N_4372,N_4022,N_3948);
nand U4373 (N_4373,N_4113,N_4175);
xor U4374 (N_4374,N_3924,N_4012);
nand U4375 (N_4375,N_4056,N_4185);
nor U4376 (N_4376,N_4077,N_3959);
and U4377 (N_4377,N_4060,N_4152);
xnor U4378 (N_4378,N_4125,N_4184);
nor U4379 (N_4379,N_4053,N_4127);
nand U4380 (N_4380,N_4140,N_4149);
nand U4381 (N_4381,N_4092,N_4001);
or U4382 (N_4382,N_4158,N_4166);
or U4383 (N_4383,N_4022,N_4094);
and U4384 (N_4384,N_4098,N_4113);
and U4385 (N_4385,N_4009,N_3941);
xor U4386 (N_4386,N_3946,N_4103);
xor U4387 (N_4387,N_4003,N_4130);
or U4388 (N_4388,N_3990,N_4108);
nand U4389 (N_4389,N_4065,N_3907);
nor U4390 (N_4390,N_3972,N_4060);
and U4391 (N_4391,N_4008,N_4086);
and U4392 (N_4392,N_4197,N_4157);
and U4393 (N_4393,N_4185,N_4180);
xor U4394 (N_4394,N_3991,N_4016);
nor U4395 (N_4395,N_3981,N_4040);
xnor U4396 (N_4396,N_4142,N_4136);
xnor U4397 (N_4397,N_3945,N_3992);
nor U4398 (N_4398,N_3980,N_4024);
xnor U4399 (N_4399,N_4194,N_4033);
and U4400 (N_4400,N_4192,N_4165);
nand U4401 (N_4401,N_4128,N_3960);
nand U4402 (N_4402,N_4188,N_4105);
or U4403 (N_4403,N_3955,N_3920);
or U4404 (N_4404,N_4169,N_3953);
nand U4405 (N_4405,N_4142,N_4171);
and U4406 (N_4406,N_4032,N_4136);
nand U4407 (N_4407,N_3949,N_4003);
xor U4408 (N_4408,N_3932,N_4139);
xnor U4409 (N_4409,N_4196,N_3908);
and U4410 (N_4410,N_4145,N_3907);
xor U4411 (N_4411,N_4018,N_4193);
nor U4412 (N_4412,N_4131,N_4165);
xnor U4413 (N_4413,N_4015,N_4128);
and U4414 (N_4414,N_3905,N_4034);
nand U4415 (N_4415,N_4113,N_3972);
xor U4416 (N_4416,N_3991,N_3985);
xor U4417 (N_4417,N_4173,N_3955);
nor U4418 (N_4418,N_3960,N_3908);
nor U4419 (N_4419,N_4094,N_4069);
xor U4420 (N_4420,N_4067,N_4185);
or U4421 (N_4421,N_4017,N_4175);
xnor U4422 (N_4422,N_4013,N_4016);
and U4423 (N_4423,N_3987,N_3939);
nand U4424 (N_4424,N_4039,N_4027);
or U4425 (N_4425,N_3906,N_4119);
and U4426 (N_4426,N_3955,N_4041);
or U4427 (N_4427,N_4089,N_4169);
or U4428 (N_4428,N_4158,N_3986);
and U4429 (N_4429,N_4087,N_4081);
nor U4430 (N_4430,N_3925,N_4183);
nor U4431 (N_4431,N_4046,N_4166);
and U4432 (N_4432,N_3996,N_3956);
xor U4433 (N_4433,N_4137,N_4050);
nand U4434 (N_4434,N_3977,N_3909);
nand U4435 (N_4435,N_3990,N_3978);
nand U4436 (N_4436,N_3907,N_4071);
and U4437 (N_4437,N_4098,N_3931);
and U4438 (N_4438,N_4009,N_4126);
nand U4439 (N_4439,N_3952,N_4094);
nor U4440 (N_4440,N_4120,N_4195);
and U4441 (N_4441,N_3997,N_4001);
nand U4442 (N_4442,N_4087,N_3997);
nor U4443 (N_4443,N_4093,N_3923);
and U4444 (N_4444,N_4059,N_4180);
nor U4445 (N_4445,N_4132,N_4155);
nand U4446 (N_4446,N_4002,N_4069);
or U4447 (N_4447,N_4066,N_4139);
and U4448 (N_4448,N_4083,N_4159);
xor U4449 (N_4449,N_4128,N_4139);
or U4450 (N_4450,N_4039,N_4156);
and U4451 (N_4451,N_4089,N_3926);
nor U4452 (N_4452,N_4187,N_3914);
nand U4453 (N_4453,N_3961,N_4056);
and U4454 (N_4454,N_3938,N_3962);
and U4455 (N_4455,N_3935,N_3953);
and U4456 (N_4456,N_4003,N_3999);
or U4457 (N_4457,N_3906,N_3961);
or U4458 (N_4458,N_4014,N_4148);
and U4459 (N_4459,N_3962,N_4186);
nand U4460 (N_4460,N_4070,N_3910);
nor U4461 (N_4461,N_3974,N_3931);
or U4462 (N_4462,N_3987,N_4091);
xnor U4463 (N_4463,N_4007,N_4000);
or U4464 (N_4464,N_4130,N_3946);
or U4465 (N_4465,N_4047,N_4143);
xnor U4466 (N_4466,N_3969,N_4179);
nor U4467 (N_4467,N_3928,N_4047);
and U4468 (N_4468,N_4077,N_3958);
and U4469 (N_4469,N_4105,N_4042);
xor U4470 (N_4470,N_3906,N_4000);
and U4471 (N_4471,N_4152,N_3958);
nor U4472 (N_4472,N_3992,N_4045);
xnor U4473 (N_4473,N_4007,N_3997);
or U4474 (N_4474,N_3940,N_4113);
xor U4475 (N_4475,N_4051,N_3912);
or U4476 (N_4476,N_4163,N_4189);
nand U4477 (N_4477,N_4180,N_3941);
or U4478 (N_4478,N_4049,N_4030);
and U4479 (N_4479,N_3912,N_4066);
xor U4480 (N_4480,N_4155,N_3990);
nor U4481 (N_4481,N_4027,N_4157);
nor U4482 (N_4482,N_4031,N_4156);
nand U4483 (N_4483,N_4118,N_4108);
xor U4484 (N_4484,N_3924,N_4121);
nor U4485 (N_4485,N_4117,N_4150);
nand U4486 (N_4486,N_3949,N_4187);
and U4487 (N_4487,N_3985,N_4124);
nor U4488 (N_4488,N_4144,N_4145);
and U4489 (N_4489,N_4131,N_4167);
xor U4490 (N_4490,N_3960,N_4030);
and U4491 (N_4491,N_4112,N_4076);
xnor U4492 (N_4492,N_3963,N_4181);
nand U4493 (N_4493,N_4134,N_4198);
and U4494 (N_4494,N_3970,N_4044);
xor U4495 (N_4495,N_3931,N_4089);
nor U4496 (N_4496,N_4007,N_3938);
and U4497 (N_4497,N_3991,N_4051);
xor U4498 (N_4498,N_4124,N_4129);
or U4499 (N_4499,N_4067,N_4163);
nor U4500 (N_4500,N_4475,N_4441);
xnor U4501 (N_4501,N_4378,N_4479);
nand U4502 (N_4502,N_4205,N_4332);
and U4503 (N_4503,N_4458,N_4482);
xor U4504 (N_4504,N_4296,N_4243);
nor U4505 (N_4505,N_4328,N_4455);
nand U4506 (N_4506,N_4464,N_4496);
nor U4507 (N_4507,N_4476,N_4355);
xnor U4508 (N_4508,N_4420,N_4215);
xnor U4509 (N_4509,N_4467,N_4321);
and U4510 (N_4510,N_4335,N_4316);
or U4511 (N_4511,N_4260,N_4214);
or U4512 (N_4512,N_4303,N_4320);
nor U4513 (N_4513,N_4370,N_4450);
and U4514 (N_4514,N_4213,N_4392);
or U4515 (N_4515,N_4406,N_4411);
and U4516 (N_4516,N_4346,N_4493);
nand U4517 (N_4517,N_4326,N_4389);
nand U4518 (N_4518,N_4301,N_4404);
xor U4519 (N_4519,N_4307,N_4202);
xor U4520 (N_4520,N_4402,N_4401);
nor U4521 (N_4521,N_4363,N_4414);
nand U4522 (N_4522,N_4403,N_4366);
and U4523 (N_4523,N_4294,N_4227);
nand U4524 (N_4524,N_4255,N_4290);
nand U4525 (N_4525,N_4257,N_4345);
or U4526 (N_4526,N_4422,N_4423);
xor U4527 (N_4527,N_4436,N_4372);
nand U4528 (N_4528,N_4437,N_4418);
and U4529 (N_4529,N_4409,N_4208);
and U4530 (N_4530,N_4367,N_4369);
xor U4531 (N_4531,N_4211,N_4480);
nor U4532 (N_4532,N_4415,N_4288);
xnor U4533 (N_4533,N_4276,N_4271);
nor U4534 (N_4534,N_4265,N_4241);
nor U4535 (N_4535,N_4413,N_4314);
nand U4536 (N_4536,N_4306,N_4274);
or U4537 (N_4537,N_4275,N_4286);
or U4538 (N_4538,N_4311,N_4249);
nand U4539 (N_4539,N_4349,N_4305);
nor U4540 (N_4540,N_4492,N_4262);
nand U4541 (N_4541,N_4439,N_4235);
or U4542 (N_4542,N_4353,N_4253);
or U4543 (N_4543,N_4416,N_4282);
and U4544 (N_4544,N_4310,N_4499);
and U4545 (N_4545,N_4484,N_4309);
and U4546 (N_4546,N_4435,N_4239);
nor U4547 (N_4547,N_4487,N_4340);
or U4548 (N_4548,N_4228,N_4261);
or U4549 (N_4549,N_4299,N_4448);
and U4550 (N_4550,N_4379,N_4352);
xnor U4551 (N_4551,N_4250,N_4421);
and U4552 (N_4552,N_4277,N_4319);
and U4553 (N_4553,N_4291,N_4390);
xnor U4554 (N_4554,N_4270,N_4331);
nor U4555 (N_4555,N_4407,N_4452);
or U4556 (N_4556,N_4217,N_4242);
nand U4557 (N_4557,N_4295,N_4221);
nand U4558 (N_4558,N_4490,N_4333);
xor U4559 (N_4559,N_4495,N_4298);
nand U4560 (N_4560,N_4327,N_4342);
nor U4561 (N_4561,N_4469,N_4445);
nand U4562 (N_4562,N_4489,N_4336);
nor U4563 (N_4563,N_4456,N_4280);
nand U4564 (N_4564,N_4417,N_4426);
xnor U4565 (N_4565,N_4494,N_4498);
xor U4566 (N_4566,N_4337,N_4451);
xor U4567 (N_4567,N_4364,N_4386);
or U4568 (N_4568,N_4473,N_4430);
nand U4569 (N_4569,N_4383,N_4240);
xnor U4570 (N_4570,N_4488,N_4396);
nand U4571 (N_4571,N_4442,N_4247);
xnor U4572 (N_4572,N_4334,N_4219);
and U4573 (N_4573,N_4491,N_4233);
nand U4574 (N_4574,N_4238,N_4210);
nand U4575 (N_4575,N_4360,N_4244);
nand U4576 (N_4576,N_4359,N_4324);
or U4577 (N_4577,N_4264,N_4229);
and U4578 (N_4578,N_4478,N_4382);
and U4579 (N_4579,N_4472,N_4431);
and U4580 (N_4580,N_4344,N_4209);
and U4581 (N_4581,N_4350,N_4222);
or U4582 (N_4582,N_4251,N_4485);
or U4583 (N_4583,N_4308,N_4373);
nand U4584 (N_4584,N_4293,N_4325);
nand U4585 (N_4585,N_4252,N_4384);
nand U4586 (N_4586,N_4405,N_4374);
nor U4587 (N_4587,N_4440,N_4388);
and U4588 (N_4588,N_4203,N_4393);
nor U4589 (N_4589,N_4394,N_4234);
nor U4590 (N_4590,N_4361,N_4377);
nor U4591 (N_4591,N_4471,N_4323);
or U4592 (N_4592,N_4269,N_4232);
and U4593 (N_4593,N_4343,N_4444);
nand U4594 (N_4594,N_4330,N_4297);
xor U4595 (N_4595,N_4284,N_4272);
xnor U4596 (N_4596,N_4236,N_4231);
nand U4597 (N_4597,N_4339,N_4216);
xnor U4598 (N_4598,N_4387,N_4462);
nand U4599 (N_4599,N_4438,N_4258);
xor U4600 (N_4600,N_4283,N_4453);
nand U4601 (N_4601,N_4317,N_4226);
and U4602 (N_4602,N_4245,N_4463);
or U4603 (N_4603,N_4425,N_4225);
and U4604 (N_4604,N_4347,N_4486);
or U4605 (N_4605,N_4220,N_4292);
or U4606 (N_4606,N_4304,N_4279);
nand U4607 (N_4607,N_4399,N_4204);
nand U4608 (N_4608,N_4454,N_4380);
nor U4609 (N_4609,N_4230,N_4300);
or U4610 (N_4610,N_4200,N_4313);
and U4611 (N_4611,N_4398,N_4443);
nor U4612 (N_4612,N_4424,N_4474);
or U4613 (N_4613,N_4268,N_4248);
nand U4614 (N_4614,N_4285,N_4302);
nor U4615 (N_4615,N_4206,N_4312);
xor U4616 (N_4616,N_4446,N_4212);
nand U4617 (N_4617,N_4254,N_4348);
nor U4618 (N_4618,N_4412,N_4362);
xor U4619 (N_4619,N_4322,N_4427);
nand U4620 (N_4620,N_4391,N_4429);
nor U4621 (N_4621,N_4281,N_4358);
nand U4622 (N_4622,N_4483,N_4477);
nor U4623 (N_4623,N_4461,N_4357);
nor U4624 (N_4624,N_4237,N_4267);
xnor U4625 (N_4625,N_4201,N_4428);
nor U4626 (N_4626,N_4341,N_4218);
and U4627 (N_4627,N_4223,N_4449);
and U4628 (N_4628,N_4224,N_4256);
and U4629 (N_4629,N_4259,N_4263);
and U4630 (N_4630,N_4419,N_4338);
or U4631 (N_4631,N_4356,N_4273);
or U4632 (N_4632,N_4376,N_4447);
and U4633 (N_4633,N_4395,N_4466);
or U4634 (N_4634,N_4365,N_4408);
nor U4635 (N_4635,N_4278,N_4481);
nor U4636 (N_4636,N_4468,N_4287);
and U4637 (N_4637,N_4459,N_4266);
or U4638 (N_4638,N_4351,N_4371);
and U4639 (N_4639,N_4432,N_4433);
nor U4640 (N_4640,N_4470,N_4207);
xnor U4641 (N_4641,N_4457,N_4497);
or U4642 (N_4642,N_4385,N_4246);
xor U4643 (N_4643,N_4329,N_4460);
xor U4644 (N_4644,N_4400,N_4397);
nor U4645 (N_4645,N_4318,N_4434);
nand U4646 (N_4646,N_4368,N_4410);
nor U4647 (N_4647,N_4465,N_4289);
nand U4648 (N_4648,N_4354,N_4375);
nor U4649 (N_4649,N_4315,N_4381);
xnor U4650 (N_4650,N_4399,N_4324);
nand U4651 (N_4651,N_4488,N_4292);
xor U4652 (N_4652,N_4483,N_4431);
or U4653 (N_4653,N_4326,N_4333);
or U4654 (N_4654,N_4411,N_4369);
nand U4655 (N_4655,N_4394,N_4229);
nor U4656 (N_4656,N_4362,N_4317);
and U4657 (N_4657,N_4298,N_4442);
and U4658 (N_4658,N_4227,N_4321);
and U4659 (N_4659,N_4210,N_4381);
xor U4660 (N_4660,N_4334,N_4314);
nor U4661 (N_4661,N_4222,N_4404);
xnor U4662 (N_4662,N_4212,N_4210);
nand U4663 (N_4663,N_4428,N_4423);
xor U4664 (N_4664,N_4409,N_4324);
nand U4665 (N_4665,N_4321,N_4435);
or U4666 (N_4666,N_4442,N_4372);
and U4667 (N_4667,N_4231,N_4443);
nand U4668 (N_4668,N_4455,N_4374);
nand U4669 (N_4669,N_4490,N_4323);
and U4670 (N_4670,N_4395,N_4427);
xor U4671 (N_4671,N_4482,N_4253);
or U4672 (N_4672,N_4499,N_4234);
nor U4673 (N_4673,N_4284,N_4261);
or U4674 (N_4674,N_4346,N_4473);
nor U4675 (N_4675,N_4384,N_4311);
nand U4676 (N_4676,N_4489,N_4390);
or U4677 (N_4677,N_4416,N_4421);
and U4678 (N_4678,N_4481,N_4288);
or U4679 (N_4679,N_4476,N_4450);
or U4680 (N_4680,N_4314,N_4268);
or U4681 (N_4681,N_4328,N_4380);
nor U4682 (N_4682,N_4313,N_4467);
xor U4683 (N_4683,N_4297,N_4481);
and U4684 (N_4684,N_4248,N_4223);
or U4685 (N_4685,N_4354,N_4469);
xnor U4686 (N_4686,N_4274,N_4428);
or U4687 (N_4687,N_4367,N_4443);
nor U4688 (N_4688,N_4300,N_4231);
and U4689 (N_4689,N_4290,N_4320);
nand U4690 (N_4690,N_4268,N_4430);
nor U4691 (N_4691,N_4494,N_4203);
xnor U4692 (N_4692,N_4287,N_4217);
nand U4693 (N_4693,N_4327,N_4398);
nor U4694 (N_4694,N_4218,N_4219);
and U4695 (N_4695,N_4231,N_4226);
nand U4696 (N_4696,N_4233,N_4483);
nor U4697 (N_4697,N_4238,N_4440);
or U4698 (N_4698,N_4265,N_4347);
or U4699 (N_4699,N_4456,N_4481);
nor U4700 (N_4700,N_4460,N_4452);
nor U4701 (N_4701,N_4459,N_4216);
nor U4702 (N_4702,N_4369,N_4451);
xnor U4703 (N_4703,N_4476,N_4210);
or U4704 (N_4704,N_4288,N_4450);
nand U4705 (N_4705,N_4294,N_4214);
nand U4706 (N_4706,N_4391,N_4395);
nand U4707 (N_4707,N_4346,N_4423);
nor U4708 (N_4708,N_4381,N_4249);
nand U4709 (N_4709,N_4464,N_4379);
and U4710 (N_4710,N_4298,N_4337);
nor U4711 (N_4711,N_4486,N_4485);
or U4712 (N_4712,N_4227,N_4382);
and U4713 (N_4713,N_4444,N_4263);
or U4714 (N_4714,N_4376,N_4430);
or U4715 (N_4715,N_4210,N_4365);
or U4716 (N_4716,N_4402,N_4251);
or U4717 (N_4717,N_4453,N_4240);
xor U4718 (N_4718,N_4337,N_4330);
and U4719 (N_4719,N_4286,N_4356);
xor U4720 (N_4720,N_4270,N_4272);
nand U4721 (N_4721,N_4436,N_4250);
xnor U4722 (N_4722,N_4371,N_4343);
xnor U4723 (N_4723,N_4342,N_4406);
and U4724 (N_4724,N_4330,N_4201);
and U4725 (N_4725,N_4268,N_4338);
nand U4726 (N_4726,N_4220,N_4343);
nand U4727 (N_4727,N_4476,N_4453);
xnor U4728 (N_4728,N_4416,N_4407);
nor U4729 (N_4729,N_4295,N_4297);
nand U4730 (N_4730,N_4434,N_4425);
or U4731 (N_4731,N_4206,N_4247);
nor U4732 (N_4732,N_4275,N_4456);
or U4733 (N_4733,N_4276,N_4435);
xnor U4734 (N_4734,N_4341,N_4346);
xor U4735 (N_4735,N_4275,N_4287);
and U4736 (N_4736,N_4329,N_4240);
nor U4737 (N_4737,N_4430,N_4479);
nor U4738 (N_4738,N_4224,N_4357);
nor U4739 (N_4739,N_4298,N_4214);
nor U4740 (N_4740,N_4429,N_4373);
xor U4741 (N_4741,N_4437,N_4310);
and U4742 (N_4742,N_4228,N_4202);
nand U4743 (N_4743,N_4448,N_4226);
xor U4744 (N_4744,N_4331,N_4252);
xnor U4745 (N_4745,N_4322,N_4313);
xor U4746 (N_4746,N_4367,N_4323);
nor U4747 (N_4747,N_4367,N_4349);
nand U4748 (N_4748,N_4209,N_4355);
or U4749 (N_4749,N_4251,N_4394);
and U4750 (N_4750,N_4203,N_4272);
nand U4751 (N_4751,N_4430,N_4250);
nor U4752 (N_4752,N_4331,N_4295);
or U4753 (N_4753,N_4450,N_4283);
and U4754 (N_4754,N_4461,N_4302);
nand U4755 (N_4755,N_4301,N_4375);
and U4756 (N_4756,N_4467,N_4407);
or U4757 (N_4757,N_4422,N_4233);
or U4758 (N_4758,N_4215,N_4336);
and U4759 (N_4759,N_4413,N_4363);
and U4760 (N_4760,N_4362,N_4212);
nor U4761 (N_4761,N_4449,N_4377);
or U4762 (N_4762,N_4277,N_4430);
and U4763 (N_4763,N_4483,N_4344);
xnor U4764 (N_4764,N_4457,N_4399);
and U4765 (N_4765,N_4432,N_4465);
nand U4766 (N_4766,N_4304,N_4420);
xor U4767 (N_4767,N_4263,N_4279);
nand U4768 (N_4768,N_4227,N_4410);
nand U4769 (N_4769,N_4489,N_4303);
nor U4770 (N_4770,N_4493,N_4453);
nor U4771 (N_4771,N_4303,N_4334);
xor U4772 (N_4772,N_4282,N_4255);
xnor U4773 (N_4773,N_4465,N_4288);
nor U4774 (N_4774,N_4203,N_4240);
or U4775 (N_4775,N_4380,N_4434);
or U4776 (N_4776,N_4331,N_4431);
nand U4777 (N_4777,N_4367,N_4432);
and U4778 (N_4778,N_4301,N_4439);
and U4779 (N_4779,N_4460,N_4486);
nor U4780 (N_4780,N_4236,N_4323);
and U4781 (N_4781,N_4273,N_4334);
xnor U4782 (N_4782,N_4413,N_4205);
nor U4783 (N_4783,N_4318,N_4268);
and U4784 (N_4784,N_4374,N_4251);
nor U4785 (N_4785,N_4472,N_4498);
xnor U4786 (N_4786,N_4415,N_4240);
nand U4787 (N_4787,N_4405,N_4494);
nor U4788 (N_4788,N_4455,N_4439);
nand U4789 (N_4789,N_4241,N_4379);
or U4790 (N_4790,N_4437,N_4315);
or U4791 (N_4791,N_4280,N_4399);
nor U4792 (N_4792,N_4425,N_4491);
or U4793 (N_4793,N_4357,N_4441);
or U4794 (N_4794,N_4482,N_4443);
nand U4795 (N_4795,N_4310,N_4220);
or U4796 (N_4796,N_4368,N_4408);
and U4797 (N_4797,N_4282,N_4384);
nand U4798 (N_4798,N_4352,N_4259);
or U4799 (N_4799,N_4365,N_4325);
or U4800 (N_4800,N_4547,N_4646);
xnor U4801 (N_4801,N_4531,N_4794);
xor U4802 (N_4802,N_4691,N_4769);
or U4803 (N_4803,N_4654,N_4557);
or U4804 (N_4804,N_4696,N_4663);
nand U4805 (N_4805,N_4608,N_4510);
nor U4806 (N_4806,N_4614,N_4522);
nor U4807 (N_4807,N_4552,N_4788);
xnor U4808 (N_4808,N_4661,N_4752);
or U4809 (N_4809,N_4618,N_4509);
and U4810 (N_4810,N_4605,N_4591);
and U4811 (N_4811,N_4527,N_4520);
nand U4812 (N_4812,N_4683,N_4727);
nor U4813 (N_4813,N_4664,N_4759);
nor U4814 (N_4814,N_4740,N_4659);
nor U4815 (N_4815,N_4561,N_4785);
or U4816 (N_4816,N_4538,N_4628);
nor U4817 (N_4817,N_4519,N_4559);
and U4818 (N_4818,N_4710,N_4736);
or U4819 (N_4819,N_4501,N_4513);
nor U4820 (N_4820,N_4641,N_4745);
and U4821 (N_4821,N_4570,N_4731);
xor U4822 (N_4822,N_4762,N_4582);
and U4823 (N_4823,N_4596,N_4542);
xnor U4824 (N_4824,N_4624,N_4611);
nand U4825 (N_4825,N_4755,N_4653);
or U4826 (N_4826,N_4524,N_4715);
and U4827 (N_4827,N_4790,N_4535);
or U4828 (N_4828,N_4729,N_4717);
nand U4829 (N_4829,N_4604,N_4616);
or U4830 (N_4830,N_4636,N_4598);
and U4831 (N_4831,N_4627,N_4673);
or U4832 (N_4832,N_4669,N_4503);
and U4833 (N_4833,N_4766,N_4656);
nor U4834 (N_4834,N_4723,N_4711);
and U4835 (N_4835,N_4692,N_4568);
nor U4836 (N_4836,N_4774,N_4776);
xor U4837 (N_4837,N_4595,N_4645);
nor U4838 (N_4838,N_4599,N_4639);
nor U4839 (N_4839,N_4697,N_4625);
or U4840 (N_4840,N_4682,N_4584);
and U4841 (N_4841,N_4630,N_4648);
or U4842 (N_4842,N_4667,N_4617);
and U4843 (N_4843,N_4665,N_4734);
nor U4844 (N_4844,N_4721,N_4743);
and U4845 (N_4845,N_4702,N_4797);
and U4846 (N_4846,N_4754,N_4571);
nand U4847 (N_4847,N_4508,N_4767);
nor U4848 (N_4848,N_4747,N_4716);
and U4849 (N_4849,N_4576,N_4647);
xor U4850 (N_4850,N_4791,N_4670);
xor U4851 (N_4851,N_4578,N_4744);
nand U4852 (N_4852,N_4675,N_4523);
nand U4853 (N_4853,N_4572,N_4703);
or U4854 (N_4854,N_4735,N_4511);
nor U4855 (N_4855,N_4560,N_4534);
or U4856 (N_4856,N_4550,N_4640);
and U4857 (N_4857,N_4622,N_4589);
xnor U4858 (N_4858,N_4719,N_4540);
nand U4859 (N_4859,N_4699,N_4554);
nor U4860 (N_4860,N_4693,N_4521);
or U4861 (N_4861,N_4565,N_4756);
and U4862 (N_4862,N_4563,N_4603);
nor U4863 (N_4863,N_4761,N_4671);
xnor U4864 (N_4864,N_4757,N_4526);
and U4865 (N_4865,N_4587,N_4546);
or U4866 (N_4866,N_4753,N_4748);
nor U4867 (N_4867,N_4606,N_4610);
nand U4868 (N_4868,N_4738,N_4585);
and U4869 (N_4869,N_4631,N_4718);
nor U4870 (N_4870,N_4662,N_4643);
and U4871 (N_4871,N_4732,N_4629);
nand U4872 (N_4872,N_4679,N_4515);
nand U4873 (N_4873,N_4537,N_4666);
or U4874 (N_4874,N_4658,N_4607);
nand U4875 (N_4875,N_4741,N_4613);
nand U4876 (N_4876,N_4650,N_4612);
xnor U4877 (N_4877,N_4601,N_4507);
or U4878 (N_4878,N_4566,N_4698);
nor U4879 (N_4879,N_4765,N_4768);
xor U4880 (N_4880,N_4724,N_4713);
xor U4881 (N_4881,N_4660,N_4701);
nor U4882 (N_4882,N_4553,N_4620);
nor U4883 (N_4883,N_4548,N_4581);
xor U4884 (N_4884,N_4615,N_4635);
nor U4885 (N_4885,N_4798,N_4712);
nand U4886 (N_4886,N_4577,N_4760);
xnor U4887 (N_4887,N_4708,N_4651);
or U4888 (N_4888,N_4782,N_4784);
nor U4889 (N_4889,N_4539,N_4558);
and U4890 (N_4890,N_4792,N_4525);
or U4891 (N_4891,N_4771,N_4586);
and U4892 (N_4892,N_4500,N_4725);
nand U4893 (N_4893,N_4544,N_4677);
xor U4894 (N_4894,N_4714,N_4530);
nand U4895 (N_4895,N_4730,N_4728);
nor U4896 (N_4896,N_4583,N_4686);
or U4897 (N_4897,N_4632,N_4580);
xor U4898 (N_4898,N_4750,N_4770);
xor U4899 (N_4899,N_4758,N_4781);
nand U4900 (N_4900,N_4700,N_4705);
xnor U4901 (N_4901,N_4786,N_4795);
nand U4902 (N_4902,N_4609,N_4575);
nand U4903 (N_4903,N_4574,N_4742);
and U4904 (N_4904,N_4678,N_4739);
nand U4905 (N_4905,N_4545,N_4655);
or U4906 (N_4906,N_4516,N_4668);
nand U4907 (N_4907,N_4555,N_4778);
nor U4908 (N_4908,N_4514,N_4690);
nand U4909 (N_4909,N_4592,N_4796);
or U4910 (N_4910,N_4681,N_4504);
nor U4911 (N_4911,N_4532,N_4619);
or U4912 (N_4912,N_4597,N_4689);
xnor U4913 (N_4913,N_4564,N_4777);
and U4914 (N_4914,N_4556,N_4623);
nor U4915 (N_4915,N_4704,N_4793);
xnor U4916 (N_4916,N_4528,N_4707);
nor U4917 (N_4917,N_4685,N_4764);
nor U4918 (N_4918,N_4680,N_4674);
or U4919 (N_4919,N_4621,N_4789);
nor U4920 (N_4920,N_4652,N_4644);
xor U4921 (N_4921,N_4517,N_4657);
xor U4922 (N_4922,N_4783,N_4694);
nand U4923 (N_4923,N_4590,N_4518);
xnor U4924 (N_4924,N_4506,N_4749);
or U4925 (N_4925,N_4773,N_4746);
xor U4926 (N_4926,N_4751,N_4649);
and U4927 (N_4927,N_4638,N_4763);
nand U4928 (N_4928,N_4688,N_4672);
nand U4929 (N_4929,N_4512,N_4775);
nor U4930 (N_4930,N_4551,N_4573);
xnor U4931 (N_4931,N_4549,N_4541);
nor U4932 (N_4932,N_4634,N_4709);
nand U4933 (N_4933,N_4733,N_4772);
nor U4934 (N_4934,N_4600,N_4799);
or U4935 (N_4935,N_4676,N_4593);
nand U4936 (N_4936,N_4684,N_4787);
nor U4937 (N_4937,N_4726,N_4569);
nand U4938 (N_4938,N_4637,N_4780);
nand U4939 (N_4939,N_4687,N_4633);
nand U4940 (N_4940,N_4642,N_4588);
nand U4941 (N_4941,N_4562,N_4533);
and U4942 (N_4942,N_4720,N_4722);
or U4943 (N_4943,N_4737,N_4695);
nor U4944 (N_4944,N_4505,N_4706);
nand U4945 (N_4945,N_4602,N_4536);
xnor U4946 (N_4946,N_4529,N_4594);
nand U4947 (N_4947,N_4543,N_4502);
nor U4948 (N_4948,N_4626,N_4567);
nor U4949 (N_4949,N_4779,N_4579);
nor U4950 (N_4950,N_4649,N_4589);
and U4951 (N_4951,N_4749,N_4709);
or U4952 (N_4952,N_4516,N_4721);
nand U4953 (N_4953,N_4781,N_4530);
nand U4954 (N_4954,N_4783,N_4546);
or U4955 (N_4955,N_4720,N_4781);
nand U4956 (N_4956,N_4583,N_4683);
xor U4957 (N_4957,N_4631,N_4588);
or U4958 (N_4958,N_4778,N_4559);
or U4959 (N_4959,N_4542,N_4582);
nand U4960 (N_4960,N_4772,N_4648);
nor U4961 (N_4961,N_4562,N_4737);
nand U4962 (N_4962,N_4621,N_4622);
or U4963 (N_4963,N_4659,N_4772);
xor U4964 (N_4964,N_4762,N_4785);
nand U4965 (N_4965,N_4523,N_4603);
or U4966 (N_4966,N_4766,N_4660);
and U4967 (N_4967,N_4601,N_4712);
xnor U4968 (N_4968,N_4749,N_4531);
nand U4969 (N_4969,N_4735,N_4683);
and U4970 (N_4970,N_4784,N_4517);
nand U4971 (N_4971,N_4703,N_4539);
nor U4972 (N_4972,N_4588,N_4548);
xor U4973 (N_4973,N_4530,N_4690);
xnor U4974 (N_4974,N_4728,N_4539);
and U4975 (N_4975,N_4692,N_4758);
or U4976 (N_4976,N_4614,N_4770);
nand U4977 (N_4977,N_4581,N_4655);
nor U4978 (N_4978,N_4527,N_4777);
nor U4979 (N_4979,N_4759,N_4576);
nor U4980 (N_4980,N_4666,N_4791);
nor U4981 (N_4981,N_4548,N_4619);
nand U4982 (N_4982,N_4518,N_4724);
nand U4983 (N_4983,N_4631,N_4501);
nor U4984 (N_4984,N_4750,N_4715);
xor U4985 (N_4985,N_4571,N_4703);
or U4986 (N_4986,N_4561,N_4707);
nor U4987 (N_4987,N_4595,N_4664);
xor U4988 (N_4988,N_4602,N_4555);
and U4989 (N_4989,N_4615,N_4755);
nand U4990 (N_4990,N_4585,N_4678);
nand U4991 (N_4991,N_4534,N_4705);
and U4992 (N_4992,N_4619,N_4757);
nor U4993 (N_4993,N_4526,N_4793);
and U4994 (N_4994,N_4675,N_4588);
and U4995 (N_4995,N_4625,N_4556);
and U4996 (N_4996,N_4504,N_4654);
and U4997 (N_4997,N_4713,N_4542);
and U4998 (N_4998,N_4584,N_4706);
nor U4999 (N_4999,N_4694,N_4628);
and U5000 (N_5000,N_4657,N_4688);
or U5001 (N_5001,N_4739,N_4530);
or U5002 (N_5002,N_4517,N_4744);
nand U5003 (N_5003,N_4660,N_4683);
nor U5004 (N_5004,N_4652,N_4593);
xor U5005 (N_5005,N_4790,N_4646);
nand U5006 (N_5006,N_4773,N_4754);
nor U5007 (N_5007,N_4666,N_4617);
nor U5008 (N_5008,N_4501,N_4607);
xnor U5009 (N_5009,N_4660,N_4591);
or U5010 (N_5010,N_4518,N_4755);
nor U5011 (N_5011,N_4541,N_4707);
xnor U5012 (N_5012,N_4771,N_4729);
nand U5013 (N_5013,N_4706,N_4647);
nand U5014 (N_5014,N_4712,N_4527);
nand U5015 (N_5015,N_4790,N_4684);
xor U5016 (N_5016,N_4540,N_4546);
nand U5017 (N_5017,N_4661,N_4624);
and U5018 (N_5018,N_4764,N_4780);
xor U5019 (N_5019,N_4612,N_4587);
and U5020 (N_5020,N_4693,N_4606);
xnor U5021 (N_5021,N_4600,N_4538);
and U5022 (N_5022,N_4598,N_4524);
nand U5023 (N_5023,N_4663,N_4695);
nor U5024 (N_5024,N_4703,N_4760);
nor U5025 (N_5025,N_4608,N_4671);
nor U5026 (N_5026,N_4515,N_4799);
nand U5027 (N_5027,N_4660,N_4549);
nand U5028 (N_5028,N_4672,N_4633);
or U5029 (N_5029,N_4705,N_4604);
nor U5030 (N_5030,N_4650,N_4754);
and U5031 (N_5031,N_4685,N_4586);
or U5032 (N_5032,N_4504,N_4501);
nor U5033 (N_5033,N_4624,N_4758);
or U5034 (N_5034,N_4573,N_4786);
and U5035 (N_5035,N_4718,N_4754);
and U5036 (N_5036,N_4682,N_4516);
nor U5037 (N_5037,N_4514,N_4783);
xnor U5038 (N_5038,N_4671,N_4711);
and U5039 (N_5039,N_4714,N_4688);
nand U5040 (N_5040,N_4704,N_4631);
nand U5041 (N_5041,N_4546,N_4534);
and U5042 (N_5042,N_4517,N_4678);
xnor U5043 (N_5043,N_4537,N_4755);
nand U5044 (N_5044,N_4796,N_4564);
xor U5045 (N_5045,N_4731,N_4687);
nand U5046 (N_5046,N_4535,N_4765);
and U5047 (N_5047,N_4540,N_4570);
nor U5048 (N_5048,N_4603,N_4578);
nand U5049 (N_5049,N_4708,N_4662);
or U5050 (N_5050,N_4632,N_4721);
nor U5051 (N_5051,N_4714,N_4766);
nand U5052 (N_5052,N_4613,N_4665);
xnor U5053 (N_5053,N_4703,N_4687);
xnor U5054 (N_5054,N_4686,N_4660);
and U5055 (N_5055,N_4763,N_4539);
and U5056 (N_5056,N_4675,N_4716);
xor U5057 (N_5057,N_4637,N_4668);
nor U5058 (N_5058,N_4664,N_4659);
nand U5059 (N_5059,N_4632,N_4548);
nand U5060 (N_5060,N_4716,N_4627);
or U5061 (N_5061,N_4764,N_4787);
and U5062 (N_5062,N_4735,N_4770);
nand U5063 (N_5063,N_4606,N_4540);
nand U5064 (N_5064,N_4761,N_4730);
nand U5065 (N_5065,N_4636,N_4783);
nand U5066 (N_5066,N_4694,N_4645);
and U5067 (N_5067,N_4775,N_4649);
and U5068 (N_5068,N_4581,N_4664);
xor U5069 (N_5069,N_4777,N_4551);
nand U5070 (N_5070,N_4761,N_4676);
nor U5071 (N_5071,N_4767,N_4742);
xor U5072 (N_5072,N_4612,N_4744);
nand U5073 (N_5073,N_4607,N_4505);
or U5074 (N_5074,N_4500,N_4637);
xnor U5075 (N_5075,N_4633,N_4778);
and U5076 (N_5076,N_4613,N_4628);
xor U5077 (N_5077,N_4736,N_4612);
or U5078 (N_5078,N_4540,N_4738);
nand U5079 (N_5079,N_4659,N_4681);
and U5080 (N_5080,N_4660,N_4691);
nor U5081 (N_5081,N_4527,N_4737);
nand U5082 (N_5082,N_4775,N_4589);
and U5083 (N_5083,N_4703,N_4511);
and U5084 (N_5084,N_4769,N_4581);
nand U5085 (N_5085,N_4661,N_4548);
nor U5086 (N_5086,N_4665,N_4554);
nor U5087 (N_5087,N_4698,N_4791);
nor U5088 (N_5088,N_4699,N_4639);
xnor U5089 (N_5089,N_4612,N_4737);
xor U5090 (N_5090,N_4740,N_4503);
nand U5091 (N_5091,N_4610,N_4750);
and U5092 (N_5092,N_4777,N_4623);
or U5093 (N_5093,N_4546,N_4635);
nor U5094 (N_5094,N_4544,N_4757);
nand U5095 (N_5095,N_4739,N_4789);
xnor U5096 (N_5096,N_4552,N_4610);
xor U5097 (N_5097,N_4693,N_4790);
or U5098 (N_5098,N_4500,N_4641);
xor U5099 (N_5099,N_4753,N_4559);
xnor U5100 (N_5100,N_5064,N_4876);
nor U5101 (N_5101,N_4883,N_5059);
and U5102 (N_5102,N_4811,N_4822);
or U5103 (N_5103,N_5016,N_5046);
nor U5104 (N_5104,N_4870,N_4878);
nand U5105 (N_5105,N_4961,N_4980);
or U5106 (N_5106,N_5006,N_4999);
nor U5107 (N_5107,N_4918,N_5002);
xnor U5108 (N_5108,N_5092,N_4902);
xnor U5109 (N_5109,N_4917,N_4867);
or U5110 (N_5110,N_4879,N_4926);
xor U5111 (N_5111,N_4916,N_4937);
and U5112 (N_5112,N_4979,N_4829);
xnor U5113 (N_5113,N_4852,N_4825);
nand U5114 (N_5114,N_4969,N_5095);
xor U5115 (N_5115,N_4975,N_4983);
or U5116 (N_5116,N_5099,N_4903);
xor U5117 (N_5117,N_4855,N_5063);
nor U5118 (N_5118,N_4977,N_5083);
xor U5119 (N_5119,N_4843,N_4858);
nand U5120 (N_5120,N_5061,N_4828);
and U5121 (N_5121,N_4890,N_4891);
nand U5122 (N_5122,N_4957,N_4945);
or U5123 (N_5123,N_5060,N_5055);
nor U5124 (N_5124,N_4846,N_4987);
xor U5125 (N_5125,N_5057,N_4837);
and U5126 (N_5126,N_4992,N_4869);
nor U5127 (N_5127,N_5039,N_4936);
nor U5128 (N_5128,N_4899,N_4838);
nand U5129 (N_5129,N_4857,N_5081);
nand U5130 (N_5130,N_5037,N_5028);
xor U5131 (N_5131,N_5021,N_4823);
xor U5132 (N_5132,N_4818,N_4928);
and U5133 (N_5133,N_4904,N_4845);
nor U5134 (N_5134,N_5050,N_4915);
and U5135 (N_5135,N_4802,N_5068);
or U5136 (N_5136,N_4976,N_5071);
and U5137 (N_5137,N_4955,N_4910);
or U5138 (N_5138,N_4873,N_4972);
nand U5139 (N_5139,N_4908,N_4820);
or U5140 (N_5140,N_4839,N_4944);
or U5141 (N_5141,N_4804,N_4931);
xnor U5142 (N_5142,N_5056,N_4875);
and U5143 (N_5143,N_5031,N_5051);
xnor U5144 (N_5144,N_4991,N_5003);
or U5145 (N_5145,N_4889,N_4964);
and U5146 (N_5146,N_4914,N_5089);
nor U5147 (N_5147,N_5069,N_4895);
xor U5148 (N_5148,N_4860,N_5075);
nand U5149 (N_5149,N_4927,N_4968);
or U5150 (N_5150,N_5004,N_5033);
or U5151 (N_5151,N_5088,N_5080);
or U5152 (N_5152,N_5024,N_5085);
nor U5153 (N_5153,N_4901,N_4805);
and U5154 (N_5154,N_4863,N_4933);
and U5155 (N_5155,N_4947,N_5045);
nand U5156 (N_5156,N_4880,N_4884);
nor U5157 (N_5157,N_4866,N_4803);
and U5158 (N_5158,N_5008,N_4827);
nor U5159 (N_5159,N_4960,N_4978);
xor U5160 (N_5160,N_4924,N_5066);
and U5161 (N_5161,N_4922,N_5078);
or U5162 (N_5162,N_5035,N_4907);
nor U5163 (N_5163,N_5011,N_4913);
or U5164 (N_5164,N_4848,N_4942);
nand U5165 (N_5165,N_5026,N_5093);
or U5166 (N_5166,N_4851,N_5043);
and U5167 (N_5167,N_5030,N_5079);
xnor U5168 (N_5168,N_5023,N_4836);
nor U5169 (N_5169,N_5067,N_4919);
nor U5170 (N_5170,N_4994,N_4952);
and U5171 (N_5171,N_4993,N_5047);
nand U5172 (N_5172,N_4959,N_4988);
nand U5173 (N_5173,N_5005,N_4941);
nand U5174 (N_5174,N_4830,N_4864);
nand U5175 (N_5175,N_5074,N_4953);
and U5176 (N_5176,N_5013,N_5082);
or U5177 (N_5177,N_5084,N_5049);
nor U5178 (N_5178,N_5042,N_5040);
xnor U5179 (N_5179,N_4989,N_4990);
or U5180 (N_5180,N_4974,N_5032);
xor U5181 (N_5181,N_4859,N_4842);
or U5182 (N_5182,N_5025,N_4935);
nand U5183 (N_5183,N_4810,N_4970);
nor U5184 (N_5184,N_4963,N_4939);
or U5185 (N_5185,N_4886,N_4923);
and U5186 (N_5186,N_4949,N_4824);
or U5187 (N_5187,N_4985,N_4865);
nand U5188 (N_5188,N_4814,N_5077);
and U5189 (N_5189,N_4800,N_4853);
and U5190 (N_5190,N_4819,N_4854);
and U5191 (N_5191,N_5072,N_4995);
nor U5192 (N_5192,N_5010,N_4841);
nand U5193 (N_5193,N_4956,N_4940);
nor U5194 (N_5194,N_4905,N_4815);
nor U5195 (N_5195,N_4967,N_4888);
nand U5196 (N_5196,N_5034,N_5041);
nor U5197 (N_5197,N_5058,N_5022);
xor U5198 (N_5198,N_4998,N_4898);
nand U5199 (N_5199,N_4920,N_4816);
or U5200 (N_5200,N_5027,N_4821);
and U5201 (N_5201,N_4809,N_5019);
and U5202 (N_5202,N_4951,N_4881);
xor U5203 (N_5203,N_4877,N_5044);
and U5204 (N_5204,N_4965,N_4911);
and U5205 (N_5205,N_4892,N_4906);
and U5206 (N_5206,N_5017,N_5014);
or U5207 (N_5207,N_4982,N_5029);
or U5208 (N_5208,N_4826,N_5009);
xnor U5209 (N_5209,N_5054,N_4887);
xnor U5210 (N_5210,N_4997,N_4954);
xor U5211 (N_5211,N_4948,N_4958);
nor U5212 (N_5212,N_4835,N_4834);
xnor U5213 (N_5213,N_4847,N_4943);
xor U5214 (N_5214,N_4946,N_4882);
or U5215 (N_5215,N_4850,N_5062);
nor U5216 (N_5216,N_4801,N_4981);
or U5217 (N_5217,N_5073,N_4996);
nor U5218 (N_5218,N_5087,N_4909);
and U5219 (N_5219,N_5070,N_5097);
nand U5220 (N_5220,N_4806,N_4984);
nand U5221 (N_5221,N_4900,N_4874);
xor U5222 (N_5222,N_4813,N_5007);
nand U5223 (N_5223,N_5065,N_5052);
nand U5224 (N_5224,N_5098,N_4950);
xor U5225 (N_5225,N_4925,N_4832);
and U5226 (N_5226,N_5096,N_4840);
xor U5227 (N_5227,N_4833,N_4812);
nand U5228 (N_5228,N_5053,N_5038);
xor U5229 (N_5229,N_4849,N_4885);
or U5230 (N_5230,N_5076,N_5048);
nor U5231 (N_5231,N_4966,N_4844);
or U5232 (N_5232,N_4808,N_4896);
nor U5233 (N_5233,N_5090,N_4986);
or U5234 (N_5234,N_4897,N_4932);
xnor U5235 (N_5235,N_5094,N_4971);
nor U5236 (N_5236,N_4856,N_5012);
nor U5237 (N_5237,N_4930,N_5036);
or U5238 (N_5238,N_5001,N_4817);
and U5239 (N_5239,N_4893,N_4962);
nor U5240 (N_5240,N_5086,N_4862);
xnor U5241 (N_5241,N_4831,N_4938);
nand U5242 (N_5242,N_5091,N_5000);
nor U5243 (N_5243,N_4868,N_5018);
xor U5244 (N_5244,N_4894,N_4934);
or U5245 (N_5245,N_4929,N_5020);
xor U5246 (N_5246,N_4912,N_4872);
nand U5247 (N_5247,N_4807,N_4861);
nand U5248 (N_5248,N_4871,N_5015);
nor U5249 (N_5249,N_4973,N_4921);
nor U5250 (N_5250,N_5035,N_4968);
nand U5251 (N_5251,N_5026,N_5014);
nor U5252 (N_5252,N_4812,N_4851);
and U5253 (N_5253,N_4872,N_4995);
nor U5254 (N_5254,N_5065,N_5016);
nor U5255 (N_5255,N_5082,N_4925);
xor U5256 (N_5256,N_5087,N_4885);
or U5257 (N_5257,N_4926,N_4995);
xor U5258 (N_5258,N_4912,N_5072);
nand U5259 (N_5259,N_4922,N_5014);
xor U5260 (N_5260,N_4832,N_4989);
nor U5261 (N_5261,N_5087,N_5054);
nor U5262 (N_5262,N_4991,N_4962);
nor U5263 (N_5263,N_4925,N_4978);
and U5264 (N_5264,N_4873,N_5005);
nand U5265 (N_5265,N_4827,N_4962);
xor U5266 (N_5266,N_4836,N_4883);
nor U5267 (N_5267,N_4977,N_4947);
or U5268 (N_5268,N_4849,N_4834);
or U5269 (N_5269,N_4911,N_4981);
nand U5270 (N_5270,N_4900,N_5087);
nand U5271 (N_5271,N_4893,N_5027);
or U5272 (N_5272,N_5001,N_4890);
and U5273 (N_5273,N_4938,N_5013);
and U5274 (N_5274,N_4988,N_4904);
and U5275 (N_5275,N_4936,N_4827);
xor U5276 (N_5276,N_5055,N_4962);
nand U5277 (N_5277,N_4800,N_4842);
nor U5278 (N_5278,N_5054,N_4807);
nor U5279 (N_5279,N_4938,N_5035);
and U5280 (N_5280,N_5065,N_4827);
xor U5281 (N_5281,N_5033,N_4998);
xor U5282 (N_5282,N_5063,N_4919);
nor U5283 (N_5283,N_4965,N_4902);
xnor U5284 (N_5284,N_5005,N_4800);
nor U5285 (N_5285,N_4869,N_5045);
or U5286 (N_5286,N_4843,N_4919);
nor U5287 (N_5287,N_4895,N_4819);
xnor U5288 (N_5288,N_4899,N_4927);
nand U5289 (N_5289,N_4809,N_5053);
nand U5290 (N_5290,N_4838,N_5012);
nand U5291 (N_5291,N_4905,N_4987);
nand U5292 (N_5292,N_4904,N_4947);
and U5293 (N_5293,N_4857,N_4819);
xnor U5294 (N_5294,N_4897,N_4933);
nor U5295 (N_5295,N_5059,N_4848);
nand U5296 (N_5296,N_5067,N_4838);
xor U5297 (N_5297,N_4925,N_5012);
nor U5298 (N_5298,N_4821,N_4822);
xor U5299 (N_5299,N_4931,N_4883);
xnor U5300 (N_5300,N_4846,N_4951);
xnor U5301 (N_5301,N_4862,N_4978);
or U5302 (N_5302,N_4898,N_4861);
nand U5303 (N_5303,N_5009,N_4843);
or U5304 (N_5304,N_5057,N_4946);
nand U5305 (N_5305,N_4844,N_4818);
and U5306 (N_5306,N_4995,N_5060);
and U5307 (N_5307,N_4840,N_4876);
and U5308 (N_5308,N_4983,N_4887);
xor U5309 (N_5309,N_4964,N_4897);
xor U5310 (N_5310,N_5006,N_4937);
xnor U5311 (N_5311,N_5001,N_5008);
and U5312 (N_5312,N_4825,N_4943);
xor U5313 (N_5313,N_5060,N_5005);
nor U5314 (N_5314,N_4873,N_5079);
xnor U5315 (N_5315,N_4841,N_5052);
nand U5316 (N_5316,N_4893,N_5075);
and U5317 (N_5317,N_5069,N_5038);
xnor U5318 (N_5318,N_4816,N_4919);
and U5319 (N_5319,N_4821,N_4888);
or U5320 (N_5320,N_4904,N_5067);
xnor U5321 (N_5321,N_4969,N_4942);
and U5322 (N_5322,N_5077,N_5076);
nor U5323 (N_5323,N_5099,N_5036);
nor U5324 (N_5324,N_4800,N_4919);
nand U5325 (N_5325,N_4973,N_5042);
and U5326 (N_5326,N_5083,N_4936);
or U5327 (N_5327,N_4913,N_4815);
nor U5328 (N_5328,N_4970,N_4993);
xor U5329 (N_5329,N_4851,N_4829);
and U5330 (N_5330,N_4852,N_5017);
nand U5331 (N_5331,N_4888,N_4996);
and U5332 (N_5332,N_4814,N_4854);
nor U5333 (N_5333,N_4934,N_4979);
xor U5334 (N_5334,N_4817,N_5006);
and U5335 (N_5335,N_4860,N_4847);
nand U5336 (N_5336,N_5013,N_4935);
and U5337 (N_5337,N_4981,N_4962);
and U5338 (N_5338,N_4897,N_4994);
or U5339 (N_5339,N_4847,N_5053);
nor U5340 (N_5340,N_5061,N_4900);
and U5341 (N_5341,N_4927,N_4998);
nand U5342 (N_5342,N_4933,N_4983);
or U5343 (N_5343,N_5094,N_5046);
and U5344 (N_5344,N_4828,N_4824);
or U5345 (N_5345,N_4843,N_5064);
nand U5346 (N_5346,N_4827,N_5046);
and U5347 (N_5347,N_4875,N_4987);
nand U5348 (N_5348,N_5097,N_4892);
nor U5349 (N_5349,N_4810,N_4978);
nand U5350 (N_5350,N_5050,N_5091);
or U5351 (N_5351,N_4986,N_4959);
xnor U5352 (N_5352,N_5089,N_4983);
nand U5353 (N_5353,N_5020,N_4998);
xor U5354 (N_5354,N_5006,N_4896);
and U5355 (N_5355,N_4970,N_4988);
nor U5356 (N_5356,N_5039,N_4993);
nor U5357 (N_5357,N_5030,N_4960);
and U5358 (N_5358,N_4839,N_4932);
nor U5359 (N_5359,N_5097,N_5050);
nand U5360 (N_5360,N_5051,N_5065);
xnor U5361 (N_5361,N_5060,N_4861);
and U5362 (N_5362,N_4987,N_4979);
nor U5363 (N_5363,N_4940,N_4803);
xnor U5364 (N_5364,N_4948,N_5064);
or U5365 (N_5365,N_5098,N_4998);
nor U5366 (N_5366,N_4832,N_5049);
and U5367 (N_5367,N_4920,N_4830);
or U5368 (N_5368,N_4975,N_4932);
and U5369 (N_5369,N_4960,N_4878);
or U5370 (N_5370,N_4883,N_4913);
nor U5371 (N_5371,N_4906,N_4930);
and U5372 (N_5372,N_4959,N_4990);
nor U5373 (N_5373,N_4918,N_4888);
nor U5374 (N_5374,N_4861,N_5002);
nand U5375 (N_5375,N_5075,N_4903);
and U5376 (N_5376,N_4969,N_4817);
nand U5377 (N_5377,N_4940,N_4847);
and U5378 (N_5378,N_4928,N_4826);
or U5379 (N_5379,N_4857,N_5062);
nor U5380 (N_5380,N_4940,N_4880);
and U5381 (N_5381,N_4885,N_4934);
xor U5382 (N_5382,N_4886,N_5090);
xor U5383 (N_5383,N_4839,N_5082);
and U5384 (N_5384,N_4805,N_4895);
or U5385 (N_5385,N_4970,N_4974);
nand U5386 (N_5386,N_4900,N_4970);
xor U5387 (N_5387,N_5002,N_4939);
nor U5388 (N_5388,N_4911,N_5008);
xor U5389 (N_5389,N_4930,N_4840);
nand U5390 (N_5390,N_5000,N_4855);
nor U5391 (N_5391,N_5017,N_4828);
xnor U5392 (N_5392,N_4996,N_4891);
nand U5393 (N_5393,N_5087,N_4880);
xor U5394 (N_5394,N_4847,N_4914);
xnor U5395 (N_5395,N_4997,N_4956);
or U5396 (N_5396,N_4825,N_5052);
and U5397 (N_5397,N_4827,N_5075);
nor U5398 (N_5398,N_4963,N_4945);
and U5399 (N_5399,N_4835,N_4841);
or U5400 (N_5400,N_5175,N_5218);
or U5401 (N_5401,N_5185,N_5387);
xnor U5402 (N_5402,N_5174,N_5372);
and U5403 (N_5403,N_5297,N_5266);
or U5404 (N_5404,N_5350,N_5319);
nand U5405 (N_5405,N_5109,N_5231);
nor U5406 (N_5406,N_5283,N_5219);
nand U5407 (N_5407,N_5395,N_5230);
xnor U5408 (N_5408,N_5203,N_5178);
nor U5409 (N_5409,N_5285,N_5383);
nand U5410 (N_5410,N_5288,N_5399);
nor U5411 (N_5411,N_5132,N_5149);
or U5412 (N_5412,N_5275,N_5200);
xnor U5413 (N_5413,N_5199,N_5188);
nor U5414 (N_5414,N_5211,N_5336);
xnor U5415 (N_5415,N_5258,N_5168);
nor U5416 (N_5416,N_5257,N_5296);
or U5417 (N_5417,N_5201,N_5118);
and U5418 (N_5418,N_5346,N_5310);
or U5419 (N_5419,N_5381,N_5291);
or U5420 (N_5420,N_5194,N_5281);
or U5421 (N_5421,N_5298,N_5277);
nand U5422 (N_5422,N_5358,N_5364);
xnor U5423 (N_5423,N_5113,N_5311);
xnor U5424 (N_5424,N_5315,N_5376);
xnor U5425 (N_5425,N_5228,N_5159);
nand U5426 (N_5426,N_5127,N_5324);
and U5427 (N_5427,N_5136,N_5389);
xor U5428 (N_5428,N_5312,N_5348);
or U5429 (N_5429,N_5322,N_5371);
or U5430 (N_5430,N_5171,N_5359);
nand U5431 (N_5431,N_5183,N_5397);
xor U5432 (N_5432,N_5344,N_5162);
and U5433 (N_5433,N_5261,N_5256);
nand U5434 (N_5434,N_5313,N_5209);
xor U5435 (N_5435,N_5363,N_5130);
or U5436 (N_5436,N_5318,N_5192);
xor U5437 (N_5437,N_5213,N_5239);
nand U5438 (N_5438,N_5120,N_5169);
nand U5439 (N_5439,N_5144,N_5244);
and U5440 (N_5440,N_5375,N_5332);
xnor U5441 (N_5441,N_5260,N_5167);
or U5442 (N_5442,N_5137,N_5181);
nor U5443 (N_5443,N_5102,N_5386);
xnor U5444 (N_5444,N_5339,N_5274);
xor U5445 (N_5445,N_5151,N_5259);
xor U5446 (N_5446,N_5366,N_5202);
nand U5447 (N_5447,N_5370,N_5365);
xor U5448 (N_5448,N_5196,N_5294);
and U5449 (N_5449,N_5122,N_5119);
nor U5450 (N_5450,N_5352,N_5210);
nor U5451 (N_5451,N_5378,N_5155);
xor U5452 (N_5452,N_5327,N_5272);
xnor U5453 (N_5453,N_5304,N_5262);
or U5454 (N_5454,N_5112,N_5191);
nand U5455 (N_5455,N_5148,N_5360);
nor U5456 (N_5456,N_5245,N_5237);
nor U5457 (N_5457,N_5126,N_5341);
xor U5458 (N_5458,N_5131,N_5117);
or U5459 (N_5459,N_5320,N_5111);
nand U5460 (N_5460,N_5116,N_5100);
xnor U5461 (N_5461,N_5104,N_5152);
or U5462 (N_5462,N_5212,N_5345);
nand U5463 (N_5463,N_5314,N_5355);
and U5464 (N_5464,N_5163,N_5101);
and U5465 (N_5465,N_5161,N_5225);
nor U5466 (N_5466,N_5187,N_5128);
or U5467 (N_5467,N_5248,N_5247);
or U5468 (N_5468,N_5138,N_5103);
and U5469 (N_5469,N_5226,N_5221);
or U5470 (N_5470,N_5114,N_5160);
or U5471 (N_5471,N_5385,N_5156);
and U5472 (N_5472,N_5170,N_5217);
or U5473 (N_5473,N_5166,N_5353);
xnor U5474 (N_5474,N_5216,N_5369);
nand U5475 (N_5475,N_5110,N_5254);
and U5476 (N_5476,N_5134,N_5368);
or U5477 (N_5477,N_5306,N_5265);
or U5478 (N_5478,N_5198,N_5220);
or U5479 (N_5479,N_5269,N_5309);
and U5480 (N_5480,N_5321,N_5173);
or U5481 (N_5481,N_5164,N_5242);
or U5482 (N_5482,N_5235,N_5308);
and U5483 (N_5483,N_5271,N_5293);
nand U5484 (N_5484,N_5325,N_5382);
or U5485 (N_5485,N_5384,N_5253);
xor U5486 (N_5486,N_5316,N_5273);
xnor U5487 (N_5487,N_5195,N_5330);
and U5488 (N_5488,N_5121,N_5133);
nor U5489 (N_5489,N_5186,N_5394);
xor U5490 (N_5490,N_5232,N_5143);
xnor U5491 (N_5491,N_5165,N_5179);
nand U5492 (N_5492,N_5295,N_5205);
xor U5493 (N_5493,N_5264,N_5147);
and U5494 (N_5494,N_5227,N_5289);
nor U5495 (N_5495,N_5249,N_5391);
xor U5496 (N_5496,N_5267,N_5343);
nor U5497 (N_5497,N_5124,N_5367);
and U5498 (N_5498,N_5300,N_5252);
nor U5499 (N_5499,N_5307,N_5377);
nor U5500 (N_5500,N_5299,N_5215);
nor U5501 (N_5501,N_5190,N_5214);
and U5502 (N_5502,N_5177,N_5140);
or U5503 (N_5503,N_5331,N_5398);
xnor U5504 (N_5504,N_5234,N_5393);
nor U5505 (N_5505,N_5125,N_5270);
nand U5506 (N_5506,N_5292,N_5197);
and U5507 (N_5507,N_5263,N_5284);
nand U5508 (N_5508,N_5189,N_5207);
nor U5509 (N_5509,N_5396,N_5157);
or U5510 (N_5510,N_5141,N_5323);
xor U5511 (N_5511,N_5280,N_5184);
nor U5512 (N_5512,N_5337,N_5278);
nor U5513 (N_5513,N_5224,N_5317);
nor U5514 (N_5514,N_5240,N_5105);
or U5515 (N_5515,N_5276,N_5392);
and U5516 (N_5516,N_5373,N_5123);
nor U5517 (N_5517,N_5340,N_5333);
and U5518 (N_5518,N_5357,N_5279);
nand U5519 (N_5519,N_5390,N_5338);
and U5520 (N_5520,N_5305,N_5286);
or U5521 (N_5521,N_5241,N_5326);
or U5522 (N_5522,N_5356,N_5255);
nand U5523 (N_5523,N_5229,N_5329);
nand U5524 (N_5524,N_5223,N_5362);
xnor U5525 (N_5525,N_5290,N_5158);
or U5526 (N_5526,N_5142,N_5115);
or U5527 (N_5527,N_5342,N_5335);
nor U5528 (N_5528,N_5154,N_5246);
xnor U5529 (N_5529,N_5238,N_5374);
nor U5530 (N_5530,N_5347,N_5233);
nor U5531 (N_5531,N_5107,N_5243);
or U5532 (N_5532,N_5106,N_5222);
and U5533 (N_5533,N_5251,N_5354);
or U5534 (N_5534,N_5236,N_5129);
nand U5535 (N_5535,N_5182,N_5388);
nand U5536 (N_5536,N_5379,N_5380);
and U5537 (N_5537,N_5303,N_5334);
nand U5538 (N_5538,N_5172,N_5206);
xnor U5539 (N_5539,N_5302,N_5153);
or U5540 (N_5540,N_5193,N_5287);
nor U5541 (N_5541,N_5361,N_5180);
xnor U5542 (N_5542,N_5282,N_5135);
and U5543 (N_5543,N_5351,N_5349);
and U5544 (N_5544,N_5139,N_5301);
nand U5545 (N_5545,N_5268,N_5150);
or U5546 (N_5546,N_5108,N_5208);
nor U5547 (N_5547,N_5176,N_5328);
or U5548 (N_5548,N_5250,N_5146);
or U5549 (N_5549,N_5204,N_5145);
xnor U5550 (N_5550,N_5324,N_5185);
or U5551 (N_5551,N_5119,N_5126);
nand U5552 (N_5552,N_5124,N_5214);
xor U5553 (N_5553,N_5126,N_5369);
or U5554 (N_5554,N_5260,N_5262);
or U5555 (N_5555,N_5208,N_5306);
xor U5556 (N_5556,N_5366,N_5325);
and U5557 (N_5557,N_5148,N_5155);
or U5558 (N_5558,N_5177,N_5242);
or U5559 (N_5559,N_5385,N_5290);
and U5560 (N_5560,N_5229,N_5344);
and U5561 (N_5561,N_5339,N_5191);
and U5562 (N_5562,N_5319,N_5199);
nor U5563 (N_5563,N_5279,N_5359);
nor U5564 (N_5564,N_5216,N_5133);
or U5565 (N_5565,N_5236,N_5202);
nor U5566 (N_5566,N_5295,N_5226);
or U5567 (N_5567,N_5388,N_5305);
and U5568 (N_5568,N_5175,N_5103);
xnor U5569 (N_5569,N_5114,N_5187);
xor U5570 (N_5570,N_5206,N_5364);
xor U5571 (N_5571,N_5229,N_5306);
or U5572 (N_5572,N_5198,N_5271);
or U5573 (N_5573,N_5355,N_5261);
nor U5574 (N_5574,N_5109,N_5222);
xor U5575 (N_5575,N_5376,N_5205);
and U5576 (N_5576,N_5374,N_5132);
and U5577 (N_5577,N_5335,N_5368);
nand U5578 (N_5578,N_5101,N_5229);
nor U5579 (N_5579,N_5248,N_5298);
or U5580 (N_5580,N_5391,N_5201);
or U5581 (N_5581,N_5190,N_5161);
and U5582 (N_5582,N_5215,N_5122);
nor U5583 (N_5583,N_5260,N_5177);
nand U5584 (N_5584,N_5259,N_5237);
xor U5585 (N_5585,N_5183,N_5135);
and U5586 (N_5586,N_5203,N_5220);
nor U5587 (N_5587,N_5354,N_5273);
and U5588 (N_5588,N_5349,N_5286);
and U5589 (N_5589,N_5354,N_5175);
nand U5590 (N_5590,N_5359,N_5323);
or U5591 (N_5591,N_5230,N_5114);
nor U5592 (N_5592,N_5305,N_5279);
nand U5593 (N_5593,N_5398,N_5265);
nand U5594 (N_5594,N_5330,N_5220);
and U5595 (N_5595,N_5243,N_5384);
nor U5596 (N_5596,N_5366,N_5188);
nand U5597 (N_5597,N_5102,N_5256);
nand U5598 (N_5598,N_5240,N_5183);
xor U5599 (N_5599,N_5351,N_5184);
xnor U5600 (N_5600,N_5325,N_5118);
or U5601 (N_5601,N_5298,N_5236);
nor U5602 (N_5602,N_5359,N_5161);
or U5603 (N_5603,N_5375,N_5281);
nor U5604 (N_5604,N_5174,N_5267);
nor U5605 (N_5605,N_5175,N_5292);
or U5606 (N_5606,N_5226,N_5237);
and U5607 (N_5607,N_5244,N_5245);
nand U5608 (N_5608,N_5163,N_5368);
xor U5609 (N_5609,N_5379,N_5135);
xor U5610 (N_5610,N_5125,N_5151);
or U5611 (N_5611,N_5164,N_5147);
or U5612 (N_5612,N_5249,N_5193);
and U5613 (N_5613,N_5283,N_5151);
nor U5614 (N_5614,N_5111,N_5308);
or U5615 (N_5615,N_5144,N_5120);
or U5616 (N_5616,N_5161,N_5237);
xor U5617 (N_5617,N_5251,N_5141);
nand U5618 (N_5618,N_5124,N_5171);
nor U5619 (N_5619,N_5174,N_5204);
nor U5620 (N_5620,N_5385,N_5159);
and U5621 (N_5621,N_5391,N_5206);
xor U5622 (N_5622,N_5151,N_5257);
and U5623 (N_5623,N_5178,N_5185);
nor U5624 (N_5624,N_5132,N_5171);
nand U5625 (N_5625,N_5376,N_5374);
nor U5626 (N_5626,N_5368,N_5243);
nand U5627 (N_5627,N_5153,N_5147);
and U5628 (N_5628,N_5163,N_5167);
or U5629 (N_5629,N_5250,N_5139);
nor U5630 (N_5630,N_5256,N_5116);
or U5631 (N_5631,N_5213,N_5397);
or U5632 (N_5632,N_5243,N_5283);
or U5633 (N_5633,N_5190,N_5102);
nand U5634 (N_5634,N_5267,N_5245);
nand U5635 (N_5635,N_5397,N_5279);
or U5636 (N_5636,N_5309,N_5270);
xor U5637 (N_5637,N_5394,N_5226);
xnor U5638 (N_5638,N_5248,N_5194);
and U5639 (N_5639,N_5269,N_5113);
or U5640 (N_5640,N_5282,N_5163);
nand U5641 (N_5641,N_5233,N_5109);
or U5642 (N_5642,N_5233,N_5393);
nand U5643 (N_5643,N_5117,N_5184);
nand U5644 (N_5644,N_5295,N_5174);
nand U5645 (N_5645,N_5215,N_5295);
or U5646 (N_5646,N_5138,N_5121);
and U5647 (N_5647,N_5179,N_5304);
nand U5648 (N_5648,N_5213,N_5207);
or U5649 (N_5649,N_5170,N_5288);
xnor U5650 (N_5650,N_5283,N_5200);
xor U5651 (N_5651,N_5224,N_5276);
nand U5652 (N_5652,N_5378,N_5165);
or U5653 (N_5653,N_5100,N_5135);
nor U5654 (N_5654,N_5208,N_5194);
xnor U5655 (N_5655,N_5138,N_5111);
and U5656 (N_5656,N_5252,N_5240);
or U5657 (N_5657,N_5377,N_5287);
or U5658 (N_5658,N_5344,N_5212);
or U5659 (N_5659,N_5260,N_5315);
nor U5660 (N_5660,N_5163,N_5353);
nor U5661 (N_5661,N_5315,N_5160);
nand U5662 (N_5662,N_5382,N_5177);
nand U5663 (N_5663,N_5354,N_5350);
and U5664 (N_5664,N_5152,N_5258);
or U5665 (N_5665,N_5282,N_5182);
nor U5666 (N_5666,N_5356,N_5218);
xor U5667 (N_5667,N_5306,N_5193);
xor U5668 (N_5668,N_5364,N_5239);
and U5669 (N_5669,N_5189,N_5109);
and U5670 (N_5670,N_5255,N_5230);
xor U5671 (N_5671,N_5130,N_5382);
and U5672 (N_5672,N_5241,N_5387);
nor U5673 (N_5673,N_5374,N_5214);
or U5674 (N_5674,N_5165,N_5130);
or U5675 (N_5675,N_5150,N_5267);
xor U5676 (N_5676,N_5229,N_5322);
or U5677 (N_5677,N_5153,N_5144);
or U5678 (N_5678,N_5150,N_5310);
nand U5679 (N_5679,N_5386,N_5255);
and U5680 (N_5680,N_5247,N_5172);
and U5681 (N_5681,N_5246,N_5103);
xnor U5682 (N_5682,N_5385,N_5283);
xnor U5683 (N_5683,N_5322,N_5117);
nor U5684 (N_5684,N_5394,N_5161);
nor U5685 (N_5685,N_5110,N_5210);
or U5686 (N_5686,N_5273,N_5103);
or U5687 (N_5687,N_5113,N_5302);
and U5688 (N_5688,N_5329,N_5231);
nand U5689 (N_5689,N_5376,N_5287);
nand U5690 (N_5690,N_5288,N_5144);
or U5691 (N_5691,N_5356,N_5191);
or U5692 (N_5692,N_5330,N_5361);
and U5693 (N_5693,N_5372,N_5228);
and U5694 (N_5694,N_5261,N_5184);
nand U5695 (N_5695,N_5145,N_5316);
nand U5696 (N_5696,N_5210,N_5159);
nor U5697 (N_5697,N_5234,N_5341);
and U5698 (N_5698,N_5337,N_5211);
nor U5699 (N_5699,N_5282,N_5393);
nor U5700 (N_5700,N_5492,N_5563);
or U5701 (N_5701,N_5516,N_5684);
nand U5702 (N_5702,N_5494,N_5535);
nor U5703 (N_5703,N_5624,N_5598);
nor U5704 (N_5704,N_5580,N_5465);
nor U5705 (N_5705,N_5456,N_5448);
and U5706 (N_5706,N_5466,N_5446);
xnor U5707 (N_5707,N_5468,N_5649);
nor U5708 (N_5708,N_5634,N_5420);
xnor U5709 (N_5709,N_5609,N_5678);
nor U5710 (N_5710,N_5515,N_5425);
xor U5711 (N_5711,N_5571,N_5587);
nand U5712 (N_5712,N_5542,N_5472);
nor U5713 (N_5713,N_5558,N_5655);
nor U5714 (N_5714,N_5493,N_5540);
or U5715 (N_5715,N_5543,N_5569);
nand U5716 (N_5716,N_5443,N_5513);
nor U5717 (N_5717,N_5610,N_5663);
xor U5718 (N_5718,N_5536,N_5618);
xnor U5719 (N_5719,N_5581,N_5602);
and U5720 (N_5720,N_5686,N_5522);
or U5721 (N_5721,N_5442,N_5670);
or U5722 (N_5722,N_5632,N_5413);
xnor U5723 (N_5723,N_5652,N_5500);
nand U5724 (N_5724,N_5570,N_5672);
nor U5725 (N_5725,N_5483,N_5628);
nor U5726 (N_5726,N_5556,N_5668);
xor U5727 (N_5727,N_5635,N_5695);
nor U5728 (N_5728,N_5653,N_5585);
xnor U5729 (N_5729,N_5476,N_5694);
and U5730 (N_5730,N_5449,N_5667);
nor U5731 (N_5731,N_5407,N_5596);
or U5732 (N_5732,N_5552,N_5669);
nand U5733 (N_5733,N_5533,N_5677);
nand U5734 (N_5734,N_5429,N_5421);
xnor U5735 (N_5735,N_5441,N_5671);
nand U5736 (N_5736,N_5640,N_5625);
xnor U5737 (N_5737,N_5647,N_5477);
and U5738 (N_5738,N_5660,N_5605);
and U5739 (N_5739,N_5544,N_5498);
xnor U5740 (N_5740,N_5665,N_5532);
nor U5741 (N_5741,N_5599,N_5428);
and U5742 (N_5742,N_5683,N_5415);
or U5743 (N_5743,N_5620,N_5664);
and U5744 (N_5744,N_5588,N_5511);
nor U5745 (N_5745,N_5505,N_5507);
nand U5746 (N_5746,N_5597,N_5519);
xor U5747 (N_5747,N_5478,N_5530);
and U5748 (N_5748,N_5661,N_5528);
or U5749 (N_5749,N_5490,N_5659);
xor U5750 (N_5750,N_5502,N_5481);
xnor U5751 (N_5751,N_5523,N_5401);
nor U5752 (N_5752,N_5619,N_5525);
or U5753 (N_5753,N_5693,N_5560);
or U5754 (N_5754,N_5537,N_5583);
nand U5755 (N_5755,N_5538,N_5613);
xnor U5756 (N_5756,N_5403,N_5648);
and U5757 (N_5757,N_5408,N_5461);
xnor U5758 (N_5758,N_5574,N_5557);
and U5759 (N_5759,N_5546,N_5676);
nand U5760 (N_5760,N_5512,N_5457);
xor U5761 (N_5761,N_5549,N_5555);
xnor U5762 (N_5762,N_5612,N_5462);
xor U5763 (N_5763,N_5447,N_5651);
nand U5764 (N_5764,N_5489,N_5627);
xnor U5765 (N_5765,N_5504,N_5690);
nand U5766 (N_5766,N_5467,N_5517);
and U5767 (N_5767,N_5586,N_5554);
xor U5768 (N_5768,N_5471,N_5450);
xnor U5769 (N_5769,N_5590,N_5444);
nor U5770 (N_5770,N_5501,N_5514);
nand U5771 (N_5771,N_5642,N_5527);
xor U5772 (N_5772,N_5582,N_5688);
nand U5773 (N_5773,N_5682,N_5487);
nand U5774 (N_5774,N_5687,N_5545);
nand U5775 (N_5775,N_5521,N_5475);
xnor U5776 (N_5776,N_5548,N_5623);
nor U5777 (N_5777,N_5400,N_5680);
xnor U5778 (N_5778,N_5404,N_5430);
nor U5779 (N_5779,N_5604,N_5626);
nand U5780 (N_5780,N_5479,N_5697);
xor U5781 (N_5781,N_5611,N_5518);
and U5782 (N_5782,N_5464,N_5650);
nor U5783 (N_5783,N_5474,N_5416);
or U5784 (N_5784,N_5573,N_5509);
xor U5785 (N_5785,N_5534,N_5641);
nor U5786 (N_5786,N_5578,N_5458);
nor U5787 (N_5787,N_5454,N_5636);
nand U5788 (N_5788,N_5455,N_5491);
nand U5789 (N_5789,N_5427,N_5691);
and U5790 (N_5790,N_5414,N_5526);
nor U5791 (N_5791,N_5488,N_5572);
or U5792 (N_5792,N_5601,N_5435);
nand U5793 (N_5793,N_5411,N_5418);
xnor U5794 (N_5794,N_5459,N_5484);
and U5795 (N_5795,N_5410,N_5595);
and U5796 (N_5796,N_5562,N_5575);
nor U5797 (N_5797,N_5423,N_5480);
and U5798 (N_5798,N_5426,N_5412);
nand U5799 (N_5799,N_5674,N_5644);
or U5800 (N_5800,N_5692,N_5439);
or U5801 (N_5801,N_5654,N_5675);
nor U5802 (N_5802,N_5629,N_5436);
nor U5803 (N_5803,N_5657,N_5470);
nand U5804 (N_5804,N_5422,N_5630);
or U5805 (N_5805,N_5589,N_5594);
nand U5806 (N_5806,N_5424,N_5608);
nor U5807 (N_5807,N_5638,N_5565);
nand U5808 (N_5808,N_5531,N_5579);
nand U5809 (N_5809,N_5576,N_5432);
nor U5810 (N_5810,N_5445,N_5419);
nand U5811 (N_5811,N_5417,N_5524);
xnor U5812 (N_5812,N_5643,N_5431);
nor U5813 (N_5813,N_5409,N_5506);
or U5814 (N_5814,N_5405,N_5606);
and U5815 (N_5815,N_5406,N_5633);
nor U5816 (N_5816,N_5437,N_5566);
or U5817 (N_5817,N_5696,N_5499);
xor U5818 (N_5818,N_5681,N_5645);
xnor U5819 (N_5819,N_5550,N_5553);
nand U5820 (N_5820,N_5434,N_5658);
nand U5821 (N_5821,N_5616,N_5591);
nand U5822 (N_5822,N_5473,N_5469);
nor U5823 (N_5823,N_5577,N_5551);
nor U5824 (N_5824,N_5402,N_5520);
xor U5825 (N_5825,N_5541,N_5495);
or U5826 (N_5826,N_5460,N_5503);
nand U5827 (N_5827,N_5453,N_5637);
nor U5828 (N_5828,N_5600,N_5685);
and U5829 (N_5829,N_5539,N_5440);
nor U5830 (N_5830,N_5568,N_5485);
or U5831 (N_5831,N_5559,N_5451);
nor U5832 (N_5832,N_5621,N_5631);
xor U5833 (N_5833,N_5438,N_5567);
nor U5834 (N_5834,N_5639,N_5614);
nand U5835 (N_5835,N_5662,N_5615);
nand U5836 (N_5836,N_5584,N_5656);
xnor U5837 (N_5837,N_5646,N_5497);
xor U5838 (N_5838,N_5496,N_5433);
nand U5839 (N_5839,N_5508,N_5486);
xor U5840 (N_5840,N_5673,N_5698);
nor U5841 (N_5841,N_5463,N_5561);
and U5842 (N_5842,N_5529,N_5510);
or U5843 (N_5843,N_5592,N_5622);
xor U5844 (N_5844,N_5452,N_5593);
nor U5845 (N_5845,N_5617,N_5603);
nor U5846 (N_5846,N_5564,N_5699);
and U5847 (N_5847,N_5679,N_5482);
nor U5848 (N_5848,N_5689,N_5607);
xnor U5849 (N_5849,N_5666,N_5547);
nand U5850 (N_5850,N_5526,N_5428);
and U5851 (N_5851,N_5673,N_5503);
or U5852 (N_5852,N_5659,N_5589);
nand U5853 (N_5853,N_5545,N_5438);
xnor U5854 (N_5854,N_5564,N_5529);
nor U5855 (N_5855,N_5491,N_5661);
nand U5856 (N_5856,N_5463,N_5504);
xor U5857 (N_5857,N_5660,N_5600);
xor U5858 (N_5858,N_5514,N_5625);
xor U5859 (N_5859,N_5490,N_5498);
and U5860 (N_5860,N_5662,N_5488);
nor U5861 (N_5861,N_5686,N_5564);
xor U5862 (N_5862,N_5544,N_5444);
nor U5863 (N_5863,N_5616,N_5673);
xor U5864 (N_5864,N_5576,N_5498);
xnor U5865 (N_5865,N_5644,N_5578);
nand U5866 (N_5866,N_5400,N_5577);
or U5867 (N_5867,N_5576,N_5458);
or U5868 (N_5868,N_5671,N_5691);
nand U5869 (N_5869,N_5443,N_5686);
or U5870 (N_5870,N_5424,N_5476);
xor U5871 (N_5871,N_5626,N_5600);
or U5872 (N_5872,N_5476,N_5415);
nand U5873 (N_5873,N_5442,N_5644);
or U5874 (N_5874,N_5636,N_5556);
and U5875 (N_5875,N_5466,N_5587);
or U5876 (N_5876,N_5557,N_5636);
nor U5877 (N_5877,N_5635,N_5407);
nor U5878 (N_5878,N_5479,N_5663);
nand U5879 (N_5879,N_5458,N_5640);
nand U5880 (N_5880,N_5465,N_5477);
nand U5881 (N_5881,N_5571,N_5514);
nor U5882 (N_5882,N_5664,N_5433);
and U5883 (N_5883,N_5424,N_5489);
xor U5884 (N_5884,N_5470,N_5524);
nand U5885 (N_5885,N_5422,N_5605);
and U5886 (N_5886,N_5566,N_5620);
or U5887 (N_5887,N_5503,N_5485);
xor U5888 (N_5888,N_5685,N_5583);
xnor U5889 (N_5889,N_5406,N_5607);
nand U5890 (N_5890,N_5513,N_5630);
nor U5891 (N_5891,N_5507,N_5699);
nor U5892 (N_5892,N_5612,N_5444);
nor U5893 (N_5893,N_5461,N_5412);
nor U5894 (N_5894,N_5555,N_5670);
nor U5895 (N_5895,N_5583,N_5415);
and U5896 (N_5896,N_5606,N_5576);
and U5897 (N_5897,N_5512,N_5690);
xor U5898 (N_5898,N_5554,N_5647);
and U5899 (N_5899,N_5423,N_5682);
nand U5900 (N_5900,N_5620,N_5569);
and U5901 (N_5901,N_5405,N_5649);
and U5902 (N_5902,N_5551,N_5498);
or U5903 (N_5903,N_5421,N_5579);
or U5904 (N_5904,N_5513,N_5462);
and U5905 (N_5905,N_5489,N_5599);
xor U5906 (N_5906,N_5481,N_5618);
xnor U5907 (N_5907,N_5476,N_5405);
xor U5908 (N_5908,N_5468,N_5682);
and U5909 (N_5909,N_5631,N_5543);
nor U5910 (N_5910,N_5663,N_5587);
nand U5911 (N_5911,N_5606,N_5617);
nand U5912 (N_5912,N_5423,N_5541);
xor U5913 (N_5913,N_5554,N_5466);
nand U5914 (N_5914,N_5485,N_5445);
nor U5915 (N_5915,N_5697,N_5673);
nand U5916 (N_5916,N_5405,N_5471);
and U5917 (N_5917,N_5449,N_5585);
or U5918 (N_5918,N_5534,N_5559);
or U5919 (N_5919,N_5486,N_5415);
nand U5920 (N_5920,N_5592,N_5591);
and U5921 (N_5921,N_5542,N_5509);
xnor U5922 (N_5922,N_5613,N_5450);
and U5923 (N_5923,N_5474,N_5469);
or U5924 (N_5924,N_5473,N_5443);
or U5925 (N_5925,N_5614,N_5550);
nand U5926 (N_5926,N_5486,N_5470);
xnor U5927 (N_5927,N_5415,N_5536);
or U5928 (N_5928,N_5427,N_5554);
or U5929 (N_5929,N_5655,N_5691);
and U5930 (N_5930,N_5674,N_5432);
or U5931 (N_5931,N_5581,N_5653);
nor U5932 (N_5932,N_5529,N_5598);
nor U5933 (N_5933,N_5651,N_5499);
nor U5934 (N_5934,N_5522,N_5531);
nor U5935 (N_5935,N_5438,N_5646);
nand U5936 (N_5936,N_5519,N_5419);
and U5937 (N_5937,N_5525,N_5665);
nand U5938 (N_5938,N_5606,N_5509);
nand U5939 (N_5939,N_5516,N_5406);
nand U5940 (N_5940,N_5440,N_5519);
nand U5941 (N_5941,N_5553,N_5565);
and U5942 (N_5942,N_5695,N_5667);
or U5943 (N_5943,N_5656,N_5604);
xor U5944 (N_5944,N_5593,N_5602);
xnor U5945 (N_5945,N_5557,N_5400);
xor U5946 (N_5946,N_5695,N_5603);
xnor U5947 (N_5947,N_5537,N_5567);
nor U5948 (N_5948,N_5401,N_5624);
nor U5949 (N_5949,N_5516,N_5620);
nor U5950 (N_5950,N_5641,N_5513);
xnor U5951 (N_5951,N_5569,N_5519);
xor U5952 (N_5952,N_5472,N_5475);
or U5953 (N_5953,N_5515,N_5612);
nand U5954 (N_5954,N_5502,N_5425);
nand U5955 (N_5955,N_5582,N_5594);
or U5956 (N_5956,N_5639,N_5560);
nor U5957 (N_5957,N_5440,N_5441);
and U5958 (N_5958,N_5598,N_5493);
nand U5959 (N_5959,N_5580,N_5477);
nor U5960 (N_5960,N_5525,N_5604);
nor U5961 (N_5961,N_5542,N_5461);
or U5962 (N_5962,N_5579,N_5682);
nor U5963 (N_5963,N_5413,N_5566);
nand U5964 (N_5964,N_5549,N_5685);
or U5965 (N_5965,N_5641,N_5427);
xnor U5966 (N_5966,N_5434,N_5634);
nand U5967 (N_5967,N_5488,N_5615);
nand U5968 (N_5968,N_5439,N_5634);
and U5969 (N_5969,N_5609,N_5610);
nand U5970 (N_5970,N_5489,N_5566);
xor U5971 (N_5971,N_5564,N_5569);
nand U5972 (N_5972,N_5671,N_5672);
nand U5973 (N_5973,N_5491,N_5632);
or U5974 (N_5974,N_5420,N_5529);
nor U5975 (N_5975,N_5489,N_5681);
nor U5976 (N_5976,N_5546,N_5666);
xnor U5977 (N_5977,N_5468,N_5627);
nand U5978 (N_5978,N_5578,N_5530);
xnor U5979 (N_5979,N_5584,N_5423);
nand U5980 (N_5980,N_5565,N_5427);
nor U5981 (N_5981,N_5577,N_5401);
nor U5982 (N_5982,N_5504,N_5433);
or U5983 (N_5983,N_5668,N_5638);
xor U5984 (N_5984,N_5640,N_5517);
nor U5985 (N_5985,N_5544,N_5609);
or U5986 (N_5986,N_5440,N_5671);
nor U5987 (N_5987,N_5455,N_5675);
nor U5988 (N_5988,N_5504,N_5417);
xnor U5989 (N_5989,N_5458,N_5441);
and U5990 (N_5990,N_5456,N_5586);
nand U5991 (N_5991,N_5538,N_5642);
or U5992 (N_5992,N_5540,N_5674);
or U5993 (N_5993,N_5531,N_5639);
and U5994 (N_5994,N_5506,N_5614);
nand U5995 (N_5995,N_5511,N_5494);
xor U5996 (N_5996,N_5656,N_5484);
or U5997 (N_5997,N_5412,N_5498);
nor U5998 (N_5998,N_5557,N_5520);
nand U5999 (N_5999,N_5629,N_5555);
nand U6000 (N_6000,N_5786,N_5726);
or U6001 (N_6001,N_5912,N_5969);
or U6002 (N_6002,N_5754,N_5970);
xnor U6003 (N_6003,N_5837,N_5723);
nand U6004 (N_6004,N_5987,N_5760);
xnor U6005 (N_6005,N_5914,N_5994);
nand U6006 (N_6006,N_5979,N_5765);
or U6007 (N_6007,N_5834,N_5784);
and U6008 (N_6008,N_5818,N_5909);
nor U6009 (N_6009,N_5761,N_5932);
or U6010 (N_6010,N_5880,N_5976);
nor U6011 (N_6011,N_5958,N_5783);
or U6012 (N_6012,N_5770,N_5702);
and U6013 (N_6013,N_5758,N_5798);
xnor U6014 (N_6014,N_5944,N_5893);
nor U6015 (N_6015,N_5737,N_5771);
nor U6016 (N_6016,N_5945,N_5779);
nand U6017 (N_6017,N_5789,N_5925);
xor U6018 (N_6018,N_5719,N_5928);
or U6019 (N_6019,N_5857,N_5806);
and U6020 (N_6020,N_5750,N_5825);
or U6021 (N_6021,N_5860,N_5830);
nand U6022 (N_6022,N_5731,N_5707);
and U6023 (N_6023,N_5990,N_5950);
nand U6024 (N_6024,N_5882,N_5924);
and U6025 (N_6025,N_5910,N_5862);
xnor U6026 (N_6026,N_5817,N_5748);
nand U6027 (N_6027,N_5892,N_5858);
xor U6028 (N_6028,N_5900,N_5949);
nor U6029 (N_6029,N_5951,N_5870);
and U6030 (N_6030,N_5968,N_5859);
nor U6031 (N_6031,N_5923,N_5971);
xnor U6032 (N_6032,N_5795,N_5742);
nor U6033 (N_6033,N_5764,N_5952);
xnor U6034 (N_6034,N_5794,N_5919);
xor U6035 (N_6035,N_5883,N_5777);
nand U6036 (N_6036,N_5939,N_5986);
xor U6037 (N_6037,N_5703,N_5845);
nor U6038 (N_6038,N_5943,N_5811);
nand U6039 (N_6039,N_5984,N_5772);
nand U6040 (N_6040,N_5955,N_5962);
and U6041 (N_6041,N_5889,N_5948);
nand U6042 (N_6042,N_5769,N_5807);
nand U6043 (N_6043,N_5728,N_5868);
and U6044 (N_6044,N_5897,N_5753);
or U6045 (N_6045,N_5774,N_5793);
xnor U6046 (N_6046,N_5936,N_5978);
and U6047 (N_6047,N_5908,N_5822);
nand U6048 (N_6048,N_5716,N_5850);
nand U6049 (N_6049,N_5814,N_5813);
nand U6050 (N_6050,N_5757,N_5823);
or U6051 (N_6051,N_5735,N_5838);
xor U6052 (N_6052,N_5810,N_5864);
nor U6053 (N_6053,N_5841,N_5714);
or U6054 (N_6054,N_5740,N_5998);
nand U6055 (N_6055,N_5824,N_5993);
and U6056 (N_6056,N_5808,N_5964);
nor U6057 (N_6057,N_5729,N_5856);
nor U6058 (N_6058,N_5773,N_5886);
nor U6059 (N_6059,N_5981,N_5861);
or U6060 (N_6060,N_5790,N_5941);
nand U6061 (N_6061,N_5996,N_5960);
nand U6062 (N_6062,N_5805,N_5744);
and U6063 (N_6063,N_5835,N_5930);
nor U6064 (N_6064,N_5927,N_5706);
nor U6065 (N_6065,N_5878,N_5871);
nand U6066 (N_6066,N_5855,N_5710);
xor U6067 (N_6067,N_5872,N_5839);
nand U6068 (N_6068,N_5741,N_5942);
xor U6069 (N_6069,N_5711,N_5852);
and U6070 (N_6070,N_5926,N_5887);
xnor U6071 (N_6071,N_5791,N_5977);
or U6072 (N_6072,N_5898,N_5847);
or U6073 (N_6073,N_5727,N_5766);
and U6074 (N_6074,N_5809,N_5920);
xnor U6075 (N_6075,N_5730,N_5891);
xor U6076 (N_6076,N_5752,N_5812);
and U6077 (N_6077,N_5775,N_5989);
nand U6078 (N_6078,N_5866,N_5840);
and U6079 (N_6079,N_5995,N_5785);
nor U6080 (N_6080,N_5906,N_5999);
xnor U6081 (N_6081,N_5846,N_5946);
nand U6082 (N_6082,N_5738,N_5934);
or U6083 (N_6083,N_5875,N_5827);
xnor U6084 (N_6084,N_5983,N_5724);
xnor U6085 (N_6085,N_5718,N_5828);
or U6086 (N_6086,N_5991,N_5853);
nor U6087 (N_6087,N_5782,N_5863);
xnor U6088 (N_6088,N_5954,N_5833);
nand U6089 (N_6089,N_5778,N_5781);
nor U6090 (N_6090,N_5736,N_5751);
nor U6091 (N_6091,N_5756,N_5953);
or U6092 (N_6092,N_5988,N_5762);
xnor U6093 (N_6093,N_5816,N_5929);
nor U6094 (N_6094,N_5966,N_5869);
nor U6095 (N_6095,N_5937,N_5963);
nor U6096 (N_6096,N_5913,N_5959);
nand U6097 (N_6097,N_5961,N_5876);
or U6098 (N_6098,N_5907,N_5787);
or U6099 (N_6099,N_5901,N_5938);
nor U6100 (N_6100,N_5747,N_5836);
xor U6101 (N_6101,N_5973,N_5917);
xor U6102 (N_6102,N_5902,N_5739);
nor U6103 (N_6103,N_5715,N_5733);
and U6104 (N_6104,N_5734,N_5801);
xor U6105 (N_6105,N_5849,N_5704);
nand U6106 (N_6106,N_5896,N_5842);
xor U6107 (N_6107,N_5899,N_5722);
and U6108 (N_6108,N_5877,N_5780);
nand U6109 (N_6109,N_5884,N_5820);
or U6110 (N_6110,N_5985,N_5815);
and U6111 (N_6111,N_5796,N_5918);
and U6112 (N_6112,N_5831,N_5745);
and U6113 (N_6113,N_5865,N_5746);
and U6114 (N_6114,N_5804,N_5915);
nand U6115 (N_6115,N_5709,N_5732);
nand U6116 (N_6116,N_5705,N_5854);
or U6117 (N_6117,N_5931,N_5749);
xnor U6118 (N_6118,N_5922,N_5851);
and U6119 (N_6119,N_5997,N_5717);
nand U6120 (N_6120,N_5921,N_5972);
nand U6121 (N_6121,N_5916,N_5792);
nor U6122 (N_6122,N_5800,N_5956);
or U6123 (N_6123,N_5873,N_5874);
nand U6124 (N_6124,N_5843,N_5957);
nand U6125 (N_6125,N_5879,N_5895);
and U6126 (N_6126,N_5867,N_5992);
xor U6127 (N_6127,N_5982,N_5763);
and U6128 (N_6128,N_5725,N_5975);
xnor U6129 (N_6129,N_5799,N_5935);
xnor U6130 (N_6130,N_5890,N_5803);
and U6131 (N_6131,N_5903,N_5940);
or U6132 (N_6132,N_5802,N_5888);
and U6133 (N_6133,N_5947,N_5911);
and U6134 (N_6134,N_5788,N_5776);
nand U6135 (N_6135,N_5980,N_5768);
and U6136 (N_6136,N_5821,N_5708);
nor U6137 (N_6137,N_5881,N_5819);
xnor U6138 (N_6138,N_5720,N_5767);
xnor U6139 (N_6139,N_5829,N_5832);
or U6140 (N_6140,N_5712,N_5974);
nor U6141 (N_6141,N_5967,N_5885);
nor U6142 (N_6142,N_5713,N_5700);
or U6143 (N_6143,N_5904,N_5721);
or U6144 (N_6144,N_5759,N_5826);
nor U6145 (N_6145,N_5701,N_5743);
xnor U6146 (N_6146,N_5894,N_5844);
nand U6147 (N_6147,N_5965,N_5905);
and U6148 (N_6148,N_5755,N_5933);
and U6149 (N_6149,N_5848,N_5797);
nand U6150 (N_6150,N_5803,N_5989);
nor U6151 (N_6151,N_5792,N_5863);
nor U6152 (N_6152,N_5742,N_5950);
nand U6153 (N_6153,N_5770,N_5834);
and U6154 (N_6154,N_5938,N_5846);
xor U6155 (N_6155,N_5816,N_5886);
nor U6156 (N_6156,N_5970,N_5927);
xnor U6157 (N_6157,N_5927,N_5791);
xor U6158 (N_6158,N_5712,N_5981);
xnor U6159 (N_6159,N_5865,N_5905);
and U6160 (N_6160,N_5708,N_5834);
or U6161 (N_6161,N_5767,N_5925);
and U6162 (N_6162,N_5780,N_5747);
nand U6163 (N_6163,N_5891,N_5745);
nand U6164 (N_6164,N_5748,N_5727);
or U6165 (N_6165,N_5884,N_5843);
or U6166 (N_6166,N_5794,N_5962);
nor U6167 (N_6167,N_5942,N_5969);
and U6168 (N_6168,N_5769,N_5758);
xnor U6169 (N_6169,N_5763,N_5739);
nor U6170 (N_6170,N_5974,N_5853);
or U6171 (N_6171,N_5835,N_5961);
or U6172 (N_6172,N_5769,N_5768);
nor U6173 (N_6173,N_5721,N_5884);
nor U6174 (N_6174,N_5877,N_5843);
nor U6175 (N_6175,N_5970,N_5725);
and U6176 (N_6176,N_5965,N_5731);
nand U6177 (N_6177,N_5930,N_5805);
xnor U6178 (N_6178,N_5713,N_5847);
xnor U6179 (N_6179,N_5893,N_5772);
and U6180 (N_6180,N_5857,N_5741);
nand U6181 (N_6181,N_5799,N_5825);
and U6182 (N_6182,N_5754,N_5932);
nand U6183 (N_6183,N_5793,N_5873);
nor U6184 (N_6184,N_5920,N_5905);
nor U6185 (N_6185,N_5863,N_5845);
xnor U6186 (N_6186,N_5755,N_5946);
and U6187 (N_6187,N_5989,N_5964);
nor U6188 (N_6188,N_5957,N_5797);
or U6189 (N_6189,N_5935,N_5837);
or U6190 (N_6190,N_5835,N_5886);
or U6191 (N_6191,N_5861,N_5829);
or U6192 (N_6192,N_5730,N_5962);
and U6193 (N_6193,N_5991,N_5712);
and U6194 (N_6194,N_5836,N_5781);
or U6195 (N_6195,N_5754,N_5767);
xor U6196 (N_6196,N_5840,N_5891);
xnor U6197 (N_6197,N_5809,N_5927);
and U6198 (N_6198,N_5834,N_5828);
xnor U6199 (N_6199,N_5728,N_5741);
nor U6200 (N_6200,N_5843,N_5973);
nand U6201 (N_6201,N_5993,N_5777);
nor U6202 (N_6202,N_5749,N_5994);
nand U6203 (N_6203,N_5871,N_5725);
nand U6204 (N_6204,N_5797,N_5983);
and U6205 (N_6205,N_5960,N_5934);
nor U6206 (N_6206,N_5729,N_5882);
nor U6207 (N_6207,N_5713,N_5844);
or U6208 (N_6208,N_5994,N_5855);
nor U6209 (N_6209,N_5955,N_5739);
nor U6210 (N_6210,N_5944,N_5728);
nand U6211 (N_6211,N_5916,N_5743);
nor U6212 (N_6212,N_5900,N_5761);
nand U6213 (N_6213,N_5985,N_5973);
nand U6214 (N_6214,N_5928,N_5892);
xnor U6215 (N_6215,N_5906,N_5712);
and U6216 (N_6216,N_5859,N_5944);
xnor U6217 (N_6217,N_5945,N_5836);
xnor U6218 (N_6218,N_5877,N_5864);
and U6219 (N_6219,N_5921,N_5751);
nand U6220 (N_6220,N_5830,N_5955);
or U6221 (N_6221,N_5801,N_5970);
nand U6222 (N_6222,N_5796,N_5739);
and U6223 (N_6223,N_5884,N_5962);
nand U6224 (N_6224,N_5868,N_5901);
and U6225 (N_6225,N_5948,N_5824);
and U6226 (N_6226,N_5855,N_5912);
or U6227 (N_6227,N_5843,N_5961);
nor U6228 (N_6228,N_5824,N_5792);
nand U6229 (N_6229,N_5725,N_5752);
or U6230 (N_6230,N_5770,N_5944);
or U6231 (N_6231,N_5899,N_5825);
and U6232 (N_6232,N_5769,N_5863);
nor U6233 (N_6233,N_5817,N_5763);
nor U6234 (N_6234,N_5769,N_5992);
nor U6235 (N_6235,N_5819,N_5893);
nor U6236 (N_6236,N_5771,N_5762);
or U6237 (N_6237,N_5768,N_5898);
and U6238 (N_6238,N_5914,N_5982);
or U6239 (N_6239,N_5709,N_5979);
nor U6240 (N_6240,N_5708,N_5746);
nor U6241 (N_6241,N_5893,N_5804);
nand U6242 (N_6242,N_5713,N_5826);
and U6243 (N_6243,N_5786,N_5732);
nand U6244 (N_6244,N_5826,N_5953);
nand U6245 (N_6245,N_5830,N_5927);
nor U6246 (N_6246,N_5905,N_5967);
nand U6247 (N_6247,N_5805,N_5977);
nor U6248 (N_6248,N_5821,N_5714);
xnor U6249 (N_6249,N_5787,N_5791);
xnor U6250 (N_6250,N_5758,N_5773);
or U6251 (N_6251,N_5967,N_5746);
nor U6252 (N_6252,N_5878,N_5724);
or U6253 (N_6253,N_5808,N_5885);
nor U6254 (N_6254,N_5766,N_5821);
nand U6255 (N_6255,N_5751,N_5719);
xnor U6256 (N_6256,N_5860,N_5812);
or U6257 (N_6257,N_5711,N_5855);
nand U6258 (N_6258,N_5958,N_5835);
nand U6259 (N_6259,N_5759,N_5815);
and U6260 (N_6260,N_5905,N_5884);
or U6261 (N_6261,N_5710,N_5716);
or U6262 (N_6262,N_5958,N_5876);
and U6263 (N_6263,N_5735,N_5944);
xor U6264 (N_6264,N_5926,N_5976);
nor U6265 (N_6265,N_5742,N_5962);
nand U6266 (N_6266,N_5739,N_5980);
nor U6267 (N_6267,N_5821,N_5710);
nor U6268 (N_6268,N_5720,N_5895);
and U6269 (N_6269,N_5934,N_5915);
or U6270 (N_6270,N_5710,N_5817);
nand U6271 (N_6271,N_5760,N_5764);
nand U6272 (N_6272,N_5968,N_5728);
nor U6273 (N_6273,N_5914,N_5901);
nand U6274 (N_6274,N_5917,N_5961);
nand U6275 (N_6275,N_5796,N_5843);
nor U6276 (N_6276,N_5958,N_5744);
or U6277 (N_6277,N_5762,N_5748);
or U6278 (N_6278,N_5897,N_5941);
nor U6279 (N_6279,N_5745,N_5857);
or U6280 (N_6280,N_5771,N_5901);
and U6281 (N_6281,N_5704,N_5782);
nand U6282 (N_6282,N_5975,N_5853);
or U6283 (N_6283,N_5931,N_5746);
nand U6284 (N_6284,N_5920,N_5722);
or U6285 (N_6285,N_5700,N_5976);
or U6286 (N_6286,N_5993,N_5876);
or U6287 (N_6287,N_5831,N_5915);
or U6288 (N_6288,N_5701,N_5861);
nand U6289 (N_6289,N_5729,N_5998);
nand U6290 (N_6290,N_5766,N_5700);
or U6291 (N_6291,N_5897,N_5814);
and U6292 (N_6292,N_5840,N_5753);
or U6293 (N_6293,N_5707,N_5968);
and U6294 (N_6294,N_5852,N_5721);
or U6295 (N_6295,N_5830,N_5966);
xnor U6296 (N_6296,N_5985,N_5803);
xor U6297 (N_6297,N_5709,N_5936);
xnor U6298 (N_6298,N_5782,N_5956);
and U6299 (N_6299,N_5742,N_5714);
and U6300 (N_6300,N_6159,N_6074);
xnor U6301 (N_6301,N_6066,N_6138);
nor U6302 (N_6302,N_6147,N_6030);
nor U6303 (N_6303,N_6108,N_6180);
nand U6304 (N_6304,N_6255,N_6179);
or U6305 (N_6305,N_6188,N_6068);
and U6306 (N_6306,N_6232,N_6099);
xor U6307 (N_6307,N_6128,N_6004);
nor U6308 (N_6308,N_6149,N_6216);
xnor U6309 (N_6309,N_6191,N_6069);
xnor U6310 (N_6310,N_6297,N_6195);
and U6311 (N_6311,N_6111,N_6194);
xor U6312 (N_6312,N_6220,N_6127);
or U6313 (N_6313,N_6018,N_6198);
nor U6314 (N_6314,N_6235,N_6257);
nor U6315 (N_6315,N_6061,N_6243);
xor U6316 (N_6316,N_6221,N_6283);
nor U6317 (N_6317,N_6040,N_6222);
and U6318 (N_6318,N_6279,N_6148);
nor U6319 (N_6319,N_6087,N_6082);
or U6320 (N_6320,N_6201,N_6086);
xnor U6321 (N_6321,N_6136,N_6067);
xnor U6322 (N_6322,N_6072,N_6126);
nor U6323 (N_6323,N_6178,N_6223);
nor U6324 (N_6324,N_6181,N_6175);
xnor U6325 (N_6325,N_6185,N_6121);
xor U6326 (N_6326,N_6055,N_6015);
and U6327 (N_6327,N_6239,N_6139);
nor U6328 (N_6328,N_6215,N_6197);
and U6329 (N_6329,N_6098,N_6059);
nor U6330 (N_6330,N_6267,N_6282);
or U6331 (N_6331,N_6037,N_6058);
nor U6332 (N_6332,N_6025,N_6045);
or U6333 (N_6333,N_6230,N_6287);
or U6334 (N_6334,N_6106,N_6020);
and U6335 (N_6335,N_6065,N_6112);
xnor U6336 (N_6336,N_6034,N_6047);
and U6337 (N_6337,N_6078,N_6118);
nand U6338 (N_6338,N_6039,N_6295);
nor U6339 (N_6339,N_6123,N_6203);
and U6340 (N_6340,N_6049,N_6102);
or U6341 (N_6341,N_6023,N_6116);
nor U6342 (N_6342,N_6135,N_6044);
or U6343 (N_6343,N_6006,N_6028);
and U6344 (N_6344,N_6009,N_6146);
nor U6345 (N_6345,N_6027,N_6211);
or U6346 (N_6346,N_6226,N_6085);
xnor U6347 (N_6347,N_6160,N_6164);
xnor U6348 (N_6348,N_6225,N_6036);
nand U6349 (N_6349,N_6228,N_6005);
or U6350 (N_6350,N_6129,N_6212);
nor U6351 (N_6351,N_6210,N_6280);
xor U6352 (N_6352,N_6268,N_6131);
and U6353 (N_6353,N_6094,N_6275);
or U6354 (N_6354,N_6251,N_6016);
and U6355 (N_6355,N_6029,N_6177);
xnor U6356 (N_6356,N_6270,N_6064);
xor U6357 (N_6357,N_6184,N_6240);
nand U6358 (N_6358,N_6233,N_6293);
and U6359 (N_6359,N_6110,N_6153);
nand U6360 (N_6360,N_6114,N_6217);
xor U6361 (N_6361,N_6076,N_6026);
nor U6362 (N_6362,N_6238,N_6001);
and U6363 (N_6363,N_6079,N_6218);
nand U6364 (N_6364,N_6017,N_6043);
nor U6365 (N_6365,N_6057,N_6134);
nor U6366 (N_6366,N_6115,N_6281);
xnor U6367 (N_6367,N_6003,N_6167);
or U6368 (N_6368,N_6219,N_6075);
xor U6369 (N_6369,N_6091,N_6196);
and U6370 (N_6370,N_6161,N_6289);
nor U6371 (N_6371,N_6286,N_6248);
xor U6372 (N_6372,N_6207,N_6093);
nor U6373 (N_6373,N_6254,N_6182);
xnor U6374 (N_6374,N_6236,N_6272);
nand U6375 (N_6375,N_6252,N_6002);
or U6376 (N_6376,N_6033,N_6193);
or U6377 (N_6377,N_6176,N_6224);
xnor U6378 (N_6378,N_6296,N_6032);
xor U6379 (N_6379,N_6204,N_6097);
xnor U6380 (N_6380,N_6105,N_6260);
or U6381 (N_6381,N_6284,N_6051);
xnor U6382 (N_6382,N_6213,N_6038);
nor U6383 (N_6383,N_6261,N_6088);
nand U6384 (N_6384,N_6187,N_6155);
nand U6385 (N_6385,N_6151,N_6273);
and U6386 (N_6386,N_6062,N_6071);
and U6387 (N_6387,N_6258,N_6011);
nor U6388 (N_6388,N_6200,N_6092);
nand U6389 (N_6389,N_6141,N_6237);
xnor U6390 (N_6390,N_6299,N_6171);
or U6391 (N_6391,N_6170,N_6206);
nor U6392 (N_6392,N_6168,N_6124);
or U6393 (N_6393,N_6205,N_6137);
xnor U6394 (N_6394,N_6262,N_6000);
nor U6395 (N_6395,N_6104,N_6089);
and U6396 (N_6396,N_6107,N_6172);
nor U6397 (N_6397,N_6035,N_6142);
or U6398 (N_6398,N_6140,N_6242);
and U6399 (N_6399,N_6183,N_6090);
nand U6400 (N_6400,N_6103,N_6259);
and U6401 (N_6401,N_6249,N_6250);
or U6402 (N_6402,N_6241,N_6169);
or U6403 (N_6403,N_6073,N_6133);
xnor U6404 (N_6404,N_6010,N_6143);
nand U6405 (N_6405,N_6285,N_6042);
and U6406 (N_6406,N_6291,N_6165);
nand U6407 (N_6407,N_6292,N_6070);
nand U6408 (N_6408,N_6276,N_6048);
xnor U6409 (N_6409,N_6095,N_6046);
and U6410 (N_6410,N_6202,N_6278);
or U6411 (N_6411,N_6150,N_6122);
and U6412 (N_6412,N_6246,N_6125);
nor U6413 (N_6413,N_6190,N_6060);
nor U6414 (N_6414,N_6231,N_6083);
xor U6415 (N_6415,N_6157,N_6156);
and U6416 (N_6416,N_6052,N_6084);
or U6417 (N_6417,N_6008,N_6096);
xor U6418 (N_6418,N_6264,N_6119);
nor U6419 (N_6419,N_6063,N_6120);
and U6420 (N_6420,N_6199,N_6288);
nand U6421 (N_6421,N_6132,N_6152);
xnor U6422 (N_6422,N_6166,N_6209);
xnor U6423 (N_6423,N_6244,N_6274);
and U6424 (N_6424,N_6080,N_6247);
or U6425 (N_6425,N_6214,N_6245);
and U6426 (N_6426,N_6298,N_6294);
or U6427 (N_6427,N_6266,N_6173);
or U6428 (N_6428,N_6109,N_6144);
or U6429 (N_6429,N_6208,N_6192);
xor U6430 (N_6430,N_6229,N_6054);
and U6431 (N_6431,N_6101,N_6277);
xor U6432 (N_6432,N_6163,N_6265);
nand U6433 (N_6433,N_6117,N_6263);
or U6434 (N_6434,N_6050,N_6234);
and U6435 (N_6435,N_6162,N_6012);
nand U6436 (N_6436,N_6019,N_6041);
nor U6437 (N_6437,N_6158,N_6014);
and U6438 (N_6438,N_6186,N_6100);
or U6439 (N_6439,N_6013,N_6113);
xnor U6440 (N_6440,N_6271,N_6253);
nand U6441 (N_6441,N_6022,N_6130);
xnor U6442 (N_6442,N_6021,N_6053);
xor U6443 (N_6443,N_6024,N_6290);
or U6444 (N_6444,N_6056,N_6145);
nor U6445 (N_6445,N_6189,N_6256);
and U6446 (N_6446,N_6077,N_6227);
and U6447 (N_6447,N_6081,N_6269);
or U6448 (N_6448,N_6031,N_6174);
and U6449 (N_6449,N_6007,N_6154);
nand U6450 (N_6450,N_6210,N_6208);
nor U6451 (N_6451,N_6119,N_6043);
nor U6452 (N_6452,N_6258,N_6114);
nand U6453 (N_6453,N_6067,N_6016);
nor U6454 (N_6454,N_6208,N_6202);
and U6455 (N_6455,N_6106,N_6226);
and U6456 (N_6456,N_6032,N_6287);
xor U6457 (N_6457,N_6106,N_6165);
and U6458 (N_6458,N_6045,N_6243);
nor U6459 (N_6459,N_6144,N_6176);
xor U6460 (N_6460,N_6144,N_6286);
or U6461 (N_6461,N_6008,N_6124);
or U6462 (N_6462,N_6128,N_6235);
or U6463 (N_6463,N_6286,N_6278);
nand U6464 (N_6464,N_6209,N_6021);
or U6465 (N_6465,N_6151,N_6296);
or U6466 (N_6466,N_6264,N_6034);
nand U6467 (N_6467,N_6286,N_6111);
and U6468 (N_6468,N_6285,N_6053);
and U6469 (N_6469,N_6199,N_6040);
nor U6470 (N_6470,N_6124,N_6014);
or U6471 (N_6471,N_6170,N_6080);
xnor U6472 (N_6472,N_6170,N_6065);
nand U6473 (N_6473,N_6090,N_6052);
nor U6474 (N_6474,N_6131,N_6046);
or U6475 (N_6475,N_6231,N_6136);
or U6476 (N_6476,N_6119,N_6222);
or U6477 (N_6477,N_6013,N_6143);
nor U6478 (N_6478,N_6014,N_6021);
nor U6479 (N_6479,N_6110,N_6126);
nand U6480 (N_6480,N_6155,N_6103);
and U6481 (N_6481,N_6117,N_6122);
and U6482 (N_6482,N_6198,N_6012);
xnor U6483 (N_6483,N_6292,N_6055);
and U6484 (N_6484,N_6290,N_6014);
nand U6485 (N_6485,N_6041,N_6017);
or U6486 (N_6486,N_6159,N_6233);
xor U6487 (N_6487,N_6171,N_6148);
xnor U6488 (N_6488,N_6244,N_6131);
and U6489 (N_6489,N_6104,N_6218);
or U6490 (N_6490,N_6287,N_6278);
xnor U6491 (N_6491,N_6060,N_6188);
and U6492 (N_6492,N_6016,N_6026);
and U6493 (N_6493,N_6258,N_6229);
nand U6494 (N_6494,N_6207,N_6147);
nand U6495 (N_6495,N_6175,N_6232);
xor U6496 (N_6496,N_6060,N_6264);
nor U6497 (N_6497,N_6190,N_6199);
nand U6498 (N_6498,N_6095,N_6281);
nor U6499 (N_6499,N_6066,N_6115);
or U6500 (N_6500,N_6007,N_6168);
nor U6501 (N_6501,N_6262,N_6192);
nand U6502 (N_6502,N_6016,N_6278);
or U6503 (N_6503,N_6296,N_6171);
nor U6504 (N_6504,N_6050,N_6260);
xor U6505 (N_6505,N_6022,N_6137);
nor U6506 (N_6506,N_6142,N_6045);
nor U6507 (N_6507,N_6232,N_6036);
nor U6508 (N_6508,N_6012,N_6182);
xnor U6509 (N_6509,N_6027,N_6206);
and U6510 (N_6510,N_6152,N_6104);
and U6511 (N_6511,N_6009,N_6132);
xor U6512 (N_6512,N_6203,N_6009);
xnor U6513 (N_6513,N_6169,N_6174);
nor U6514 (N_6514,N_6222,N_6046);
xnor U6515 (N_6515,N_6299,N_6120);
xor U6516 (N_6516,N_6046,N_6029);
nand U6517 (N_6517,N_6140,N_6157);
nor U6518 (N_6518,N_6155,N_6072);
or U6519 (N_6519,N_6011,N_6248);
nor U6520 (N_6520,N_6012,N_6126);
xor U6521 (N_6521,N_6264,N_6232);
or U6522 (N_6522,N_6292,N_6215);
nand U6523 (N_6523,N_6005,N_6056);
nand U6524 (N_6524,N_6091,N_6176);
or U6525 (N_6525,N_6264,N_6001);
or U6526 (N_6526,N_6272,N_6284);
xnor U6527 (N_6527,N_6035,N_6294);
xor U6528 (N_6528,N_6055,N_6052);
nand U6529 (N_6529,N_6194,N_6167);
and U6530 (N_6530,N_6290,N_6216);
nor U6531 (N_6531,N_6056,N_6121);
nand U6532 (N_6532,N_6059,N_6149);
and U6533 (N_6533,N_6115,N_6079);
or U6534 (N_6534,N_6274,N_6025);
and U6535 (N_6535,N_6201,N_6008);
nor U6536 (N_6536,N_6036,N_6242);
or U6537 (N_6537,N_6166,N_6071);
and U6538 (N_6538,N_6131,N_6202);
xnor U6539 (N_6539,N_6126,N_6238);
nand U6540 (N_6540,N_6273,N_6226);
xnor U6541 (N_6541,N_6039,N_6126);
xnor U6542 (N_6542,N_6022,N_6021);
nor U6543 (N_6543,N_6053,N_6078);
xnor U6544 (N_6544,N_6185,N_6122);
nand U6545 (N_6545,N_6061,N_6028);
and U6546 (N_6546,N_6011,N_6217);
xnor U6547 (N_6547,N_6194,N_6088);
nand U6548 (N_6548,N_6142,N_6067);
nor U6549 (N_6549,N_6185,N_6267);
nand U6550 (N_6550,N_6205,N_6149);
xnor U6551 (N_6551,N_6087,N_6013);
xnor U6552 (N_6552,N_6224,N_6191);
xnor U6553 (N_6553,N_6236,N_6129);
and U6554 (N_6554,N_6177,N_6125);
nor U6555 (N_6555,N_6036,N_6299);
and U6556 (N_6556,N_6037,N_6043);
and U6557 (N_6557,N_6235,N_6093);
xnor U6558 (N_6558,N_6223,N_6289);
nor U6559 (N_6559,N_6134,N_6229);
xnor U6560 (N_6560,N_6286,N_6032);
nand U6561 (N_6561,N_6226,N_6294);
and U6562 (N_6562,N_6037,N_6119);
nor U6563 (N_6563,N_6242,N_6136);
nand U6564 (N_6564,N_6158,N_6219);
nand U6565 (N_6565,N_6131,N_6297);
xnor U6566 (N_6566,N_6097,N_6119);
xnor U6567 (N_6567,N_6150,N_6212);
and U6568 (N_6568,N_6165,N_6222);
nor U6569 (N_6569,N_6166,N_6019);
xnor U6570 (N_6570,N_6032,N_6133);
xnor U6571 (N_6571,N_6269,N_6112);
nor U6572 (N_6572,N_6076,N_6165);
nor U6573 (N_6573,N_6143,N_6086);
nor U6574 (N_6574,N_6280,N_6058);
xor U6575 (N_6575,N_6128,N_6043);
xnor U6576 (N_6576,N_6239,N_6130);
nand U6577 (N_6577,N_6067,N_6137);
and U6578 (N_6578,N_6260,N_6121);
xor U6579 (N_6579,N_6197,N_6053);
or U6580 (N_6580,N_6088,N_6126);
xor U6581 (N_6581,N_6199,N_6148);
and U6582 (N_6582,N_6190,N_6071);
xor U6583 (N_6583,N_6031,N_6249);
nor U6584 (N_6584,N_6286,N_6011);
or U6585 (N_6585,N_6098,N_6202);
nor U6586 (N_6586,N_6288,N_6188);
or U6587 (N_6587,N_6098,N_6209);
nor U6588 (N_6588,N_6255,N_6212);
nand U6589 (N_6589,N_6213,N_6046);
nor U6590 (N_6590,N_6090,N_6059);
nor U6591 (N_6591,N_6294,N_6206);
or U6592 (N_6592,N_6173,N_6271);
xnor U6593 (N_6593,N_6195,N_6166);
nand U6594 (N_6594,N_6237,N_6103);
xor U6595 (N_6595,N_6098,N_6254);
or U6596 (N_6596,N_6221,N_6216);
nand U6597 (N_6597,N_6266,N_6262);
nand U6598 (N_6598,N_6289,N_6207);
nand U6599 (N_6599,N_6152,N_6143);
and U6600 (N_6600,N_6492,N_6408);
nor U6601 (N_6601,N_6437,N_6511);
xnor U6602 (N_6602,N_6585,N_6525);
and U6603 (N_6603,N_6570,N_6329);
nand U6604 (N_6604,N_6400,N_6555);
nand U6605 (N_6605,N_6598,N_6327);
nand U6606 (N_6606,N_6491,N_6481);
xor U6607 (N_6607,N_6342,N_6427);
nand U6608 (N_6608,N_6444,N_6463);
and U6609 (N_6609,N_6411,N_6338);
nand U6610 (N_6610,N_6488,N_6592);
xnor U6611 (N_6611,N_6460,N_6371);
nor U6612 (N_6612,N_6431,N_6343);
nor U6613 (N_6613,N_6542,N_6521);
or U6614 (N_6614,N_6453,N_6550);
and U6615 (N_6615,N_6347,N_6302);
xnor U6616 (N_6616,N_6530,N_6455);
xnor U6617 (N_6617,N_6500,N_6505);
nand U6618 (N_6618,N_6375,N_6573);
nor U6619 (N_6619,N_6425,N_6357);
or U6620 (N_6620,N_6580,N_6504);
or U6621 (N_6621,N_6370,N_6313);
nor U6622 (N_6622,N_6379,N_6372);
nand U6623 (N_6623,N_6499,N_6507);
and U6624 (N_6624,N_6556,N_6386);
nor U6625 (N_6625,N_6354,N_6330);
nor U6626 (N_6626,N_6441,N_6325);
nor U6627 (N_6627,N_6515,N_6367);
xnor U6628 (N_6628,N_6454,N_6422);
and U6629 (N_6629,N_6595,N_6418);
and U6630 (N_6630,N_6552,N_6377);
and U6631 (N_6631,N_6383,N_6502);
and U6632 (N_6632,N_6308,N_6331);
nor U6633 (N_6633,N_6486,N_6541);
xor U6634 (N_6634,N_6423,N_6495);
nor U6635 (N_6635,N_6412,N_6467);
or U6636 (N_6636,N_6519,N_6376);
and U6637 (N_6637,N_6527,N_6513);
xor U6638 (N_6638,N_6588,N_6385);
nor U6639 (N_6639,N_6353,N_6483);
nor U6640 (N_6640,N_6341,N_6350);
and U6641 (N_6641,N_6438,N_6593);
xor U6642 (N_6642,N_6493,N_6594);
or U6643 (N_6643,N_6496,N_6449);
nor U6644 (N_6644,N_6458,N_6416);
and U6645 (N_6645,N_6567,N_6373);
xnor U6646 (N_6646,N_6554,N_6576);
nand U6647 (N_6647,N_6413,N_6464);
and U6648 (N_6648,N_6477,N_6524);
nor U6649 (N_6649,N_6361,N_6497);
nand U6650 (N_6650,N_6402,N_6434);
and U6651 (N_6651,N_6316,N_6475);
nand U6652 (N_6652,N_6459,N_6345);
nor U6653 (N_6653,N_6597,N_6539);
and U6654 (N_6654,N_6443,N_6358);
and U6655 (N_6655,N_6532,N_6424);
xnor U6656 (N_6656,N_6322,N_6533);
and U6657 (N_6657,N_6473,N_6366);
or U6658 (N_6658,N_6520,N_6328);
xnor U6659 (N_6659,N_6575,N_6392);
and U6660 (N_6660,N_6336,N_6476);
and U6661 (N_6661,N_6510,N_6572);
nand U6662 (N_6662,N_6586,N_6339);
and U6663 (N_6663,N_6384,N_6494);
xor U6664 (N_6664,N_6560,N_6440);
and U6665 (N_6665,N_6472,N_6360);
xnor U6666 (N_6666,N_6596,N_6523);
and U6667 (N_6667,N_6536,N_6528);
or U6668 (N_6668,N_6406,N_6566);
xnor U6669 (N_6669,N_6479,N_6590);
xor U6670 (N_6670,N_6421,N_6403);
or U6671 (N_6671,N_6387,N_6432);
xnor U6672 (N_6672,N_6482,N_6485);
xor U6673 (N_6673,N_6388,N_6396);
or U6674 (N_6674,N_6417,N_6317);
nor U6675 (N_6675,N_6518,N_6462);
xor U6676 (N_6676,N_6314,N_6538);
xnor U6677 (N_6677,N_6506,N_6436);
and U6678 (N_6678,N_6551,N_6516);
or U6679 (N_6679,N_6522,N_6351);
xnor U6680 (N_6680,N_6583,N_6321);
or U6681 (N_6681,N_6509,N_6445);
or U6682 (N_6682,N_6582,N_6562);
or U6683 (N_6683,N_6490,N_6334);
nor U6684 (N_6684,N_6461,N_6569);
or U6685 (N_6685,N_6531,N_6340);
or U6686 (N_6686,N_6355,N_6581);
xor U6687 (N_6687,N_6352,N_6315);
nand U6688 (N_6688,N_6407,N_6577);
nor U6689 (N_6689,N_6429,N_6318);
xor U6690 (N_6690,N_6584,N_6587);
nand U6691 (N_6691,N_6571,N_6549);
and U6692 (N_6692,N_6470,N_6565);
nor U6693 (N_6693,N_6397,N_6404);
xnor U6694 (N_6694,N_6394,N_6450);
nand U6695 (N_6695,N_6545,N_6517);
xor U6696 (N_6696,N_6333,N_6324);
and U6697 (N_6697,N_6484,N_6419);
and U6698 (N_6698,N_6480,N_6568);
or U6699 (N_6699,N_6382,N_6303);
nor U6700 (N_6700,N_6362,N_6442);
and U6701 (N_6701,N_6364,N_6415);
and U6702 (N_6702,N_6557,N_6301);
nor U6703 (N_6703,N_6380,N_6471);
and U6704 (N_6704,N_6448,N_6381);
and U6705 (N_6705,N_6563,N_6420);
nor U6706 (N_6706,N_6300,N_6501);
nand U6707 (N_6707,N_6564,N_6306);
and U6708 (N_6708,N_6365,N_6398);
or U6709 (N_6709,N_6319,N_6537);
nor U6710 (N_6710,N_6466,N_6410);
xnor U6711 (N_6711,N_6326,N_6428);
or U6712 (N_6712,N_6558,N_6369);
xnor U6713 (N_6713,N_6498,N_6469);
nor U6714 (N_6714,N_6363,N_6399);
and U6715 (N_6715,N_6544,N_6426);
or U6716 (N_6716,N_6478,N_6447);
nand U6717 (N_6717,N_6401,N_6307);
or U6718 (N_6718,N_6547,N_6435);
nor U6719 (N_6719,N_6579,N_6457);
and U6720 (N_6720,N_6474,N_6344);
nand U6721 (N_6721,N_6512,N_6323);
nand U6722 (N_6722,N_6335,N_6368);
nand U6723 (N_6723,N_6589,N_6439);
xnor U6724 (N_6724,N_6348,N_6446);
nor U6725 (N_6725,N_6312,N_6346);
xnor U6726 (N_6726,N_6395,N_6389);
nor U6727 (N_6727,N_6526,N_6559);
nor U6728 (N_6728,N_6390,N_6574);
nor U6729 (N_6729,N_6468,N_6487);
nor U6730 (N_6730,N_6320,N_6543);
nor U6731 (N_6731,N_6374,N_6503);
and U6732 (N_6732,N_6489,N_6465);
nand U6733 (N_6733,N_6405,N_6356);
or U6734 (N_6734,N_6535,N_6378);
and U6735 (N_6735,N_6304,N_6591);
xnor U6736 (N_6736,N_6534,N_6529);
nand U6737 (N_6737,N_6546,N_6451);
nor U6738 (N_6738,N_6311,N_6508);
or U6739 (N_6739,N_6349,N_6452);
nand U6740 (N_6740,N_6553,N_6599);
nand U6741 (N_6741,N_6332,N_6337);
nand U6742 (N_6742,N_6409,N_6540);
xor U6743 (N_6743,N_6393,N_6456);
xnor U6744 (N_6744,N_6548,N_6578);
and U6745 (N_6745,N_6310,N_6359);
nor U6746 (N_6746,N_6391,N_6305);
xor U6747 (N_6747,N_6514,N_6430);
or U6748 (N_6748,N_6433,N_6309);
nand U6749 (N_6749,N_6561,N_6414);
or U6750 (N_6750,N_6335,N_6483);
and U6751 (N_6751,N_6468,N_6438);
nand U6752 (N_6752,N_6563,N_6484);
or U6753 (N_6753,N_6335,N_6470);
and U6754 (N_6754,N_6581,N_6563);
nor U6755 (N_6755,N_6438,N_6528);
nand U6756 (N_6756,N_6398,N_6596);
nand U6757 (N_6757,N_6396,N_6597);
or U6758 (N_6758,N_6391,N_6357);
xnor U6759 (N_6759,N_6327,N_6445);
or U6760 (N_6760,N_6485,N_6384);
nand U6761 (N_6761,N_6367,N_6490);
or U6762 (N_6762,N_6312,N_6303);
and U6763 (N_6763,N_6340,N_6543);
nand U6764 (N_6764,N_6565,N_6482);
or U6765 (N_6765,N_6532,N_6547);
and U6766 (N_6766,N_6562,N_6322);
nand U6767 (N_6767,N_6400,N_6537);
nand U6768 (N_6768,N_6581,N_6313);
xnor U6769 (N_6769,N_6359,N_6331);
nor U6770 (N_6770,N_6542,N_6549);
or U6771 (N_6771,N_6555,N_6517);
xor U6772 (N_6772,N_6459,N_6462);
xnor U6773 (N_6773,N_6434,N_6582);
nand U6774 (N_6774,N_6492,N_6439);
or U6775 (N_6775,N_6415,N_6508);
nand U6776 (N_6776,N_6391,N_6566);
xor U6777 (N_6777,N_6355,N_6393);
xnor U6778 (N_6778,N_6319,N_6484);
or U6779 (N_6779,N_6360,N_6375);
or U6780 (N_6780,N_6507,N_6486);
or U6781 (N_6781,N_6581,N_6584);
nor U6782 (N_6782,N_6437,N_6494);
and U6783 (N_6783,N_6463,N_6490);
and U6784 (N_6784,N_6300,N_6576);
nor U6785 (N_6785,N_6338,N_6330);
xnor U6786 (N_6786,N_6431,N_6593);
nor U6787 (N_6787,N_6473,N_6330);
or U6788 (N_6788,N_6326,N_6361);
xnor U6789 (N_6789,N_6550,N_6327);
or U6790 (N_6790,N_6330,N_6550);
nand U6791 (N_6791,N_6376,N_6383);
xnor U6792 (N_6792,N_6501,N_6398);
and U6793 (N_6793,N_6386,N_6442);
nand U6794 (N_6794,N_6559,N_6408);
xor U6795 (N_6795,N_6333,N_6396);
or U6796 (N_6796,N_6529,N_6316);
nor U6797 (N_6797,N_6593,N_6500);
and U6798 (N_6798,N_6587,N_6520);
or U6799 (N_6799,N_6548,N_6580);
nor U6800 (N_6800,N_6541,N_6356);
and U6801 (N_6801,N_6436,N_6452);
nor U6802 (N_6802,N_6377,N_6505);
or U6803 (N_6803,N_6361,N_6560);
and U6804 (N_6804,N_6418,N_6495);
nor U6805 (N_6805,N_6591,N_6328);
xor U6806 (N_6806,N_6511,N_6433);
xnor U6807 (N_6807,N_6586,N_6305);
nand U6808 (N_6808,N_6475,N_6496);
xnor U6809 (N_6809,N_6418,N_6320);
nand U6810 (N_6810,N_6373,N_6515);
or U6811 (N_6811,N_6354,N_6470);
and U6812 (N_6812,N_6439,N_6367);
and U6813 (N_6813,N_6349,N_6556);
or U6814 (N_6814,N_6342,N_6571);
nand U6815 (N_6815,N_6411,N_6500);
and U6816 (N_6816,N_6536,N_6356);
or U6817 (N_6817,N_6494,N_6568);
xor U6818 (N_6818,N_6523,N_6433);
nand U6819 (N_6819,N_6438,N_6589);
nor U6820 (N_6820,N_6486,N_6591);
and U6821 (N_6821,N_6307,N_6530);
or U6822 (N_6822,N_6571,N_6564);
and U6823 (N_6823,N_6534,N_6448);
or U6824 (N_6824,N_6462,N_6407);
and U6825 (N_6825,N_6463,N_6358);
or U6826 (N_6826,N_6457,N_6516);
xor U6827 (N_6827,N_6519,N_6577);
and U6828 (N_6828,N_6309,N_6407);
xnor U6829 (N_6829,N_6592,N_6562);
nor U6830 (N_6830,N_6359,N_6332);
xor U6831 (N_6831,N_6390,N_6474);
xnor U6832 (N_6832,N_6339,N_6446);
and U6833 (N_6833,N_6549,N_6421);
or U6834 (N_6834,N_6482,N_6314);
and U6835 (N_6835,N_6344,N_6591);
or U6836 (N_6836,N_6563,N_6320);
nand U6837 (N_6837,N_6376,N_6523);
nand U6838 (N_6838,N_6474,N_6371);
nand U6839 (N_6839,N_6469,N_6434);
xnor U6840 (N_6840,N_6411,N_6476);
nand U6841 (N_6841,N_6490,N_6526);
or U6842 (N_6842,N_6442,N_6487);
nor U6843 (N_6843,N_6408,N_6503);
and U6844 (N_6844,N_6322,N_6559);
nand U6845 (N_6845,N_6406,N_6578);
or U6846 (N_6846,N_6449,N_6551);
xor U6847 (N_6847,N_6445,N_6407);
xnor U6848 (N_6848,N_6535,N_6423);
and U6849 (N_6849,N_6434,N_6488);
xor U6850 (N_6850,N_6572,N_6314);
nand U6851 (N_6851,N_6535,N_6583);
or U6852 (N_6852,N_6552,N_6407);
and U6853 (N_6853,N_6565,N_6506);
xor U6854 (N_6854,N_6316,N_6512);
nor U6855 (N_6855,N_6508,N_6359);
nand U6856 (N_6856,N_6417,N_6362);
and U6857 (N_6857,N_6416,N_6424);
nor U6858 (N_6858,N_6427,N_6382);
or U6859 (N_6859,N_6536,N_6474);
nor U6860 (N_6860,N_6388,N_6465);
or U6861 (N_6861,N_6374,N_6593);
and U6862 (N_6862,N_6510,N_6375);
and U6863 (N_6863,N_6495,N_6578);
and U6864 (N_6864,N_6597,N_6579);
nor U6865 (N_6865,N_6554,N_6537);
nor U6866 (N_6866,N_6585,N_6416);
and U6867 (N_6867,N_6376,N_6506);
nand U6868 (N_6868,N_6304,N_6590);
nand U6869 (N_6869,N_6424,N_6521);
nand U6870 (N_6870,N_6467,N_6368);
or U6871 (N_6871,N_6560,N_6594);
or U6872 (N_6872,N_6523,N_6435);
xor U6873 (N_6873,N_6351,N_6559);
nand U6874 (N_6874,N_6477,N_6476);
and U6875 (N_6875,N_6330,N_6405);
xor U6876 (N_6876,N_6532,N_6389);
xor U6877 (N_6877,N_6352,N_6562);
xnor U6878 (N_6878,N_6501,N_6399);
and U6879 (N_6879,N_6552,N_6595);
xnor U6880 (N_6880,N_6329,N_6524);
xor U6881 (N_6881,N_6423,N_6582);
nor U6882 (N_6882,N_6542,N_6369);
or U6883 (N_6883,N_6417,N_6586);
and U6884 (N_6884,N_6320,N_6374);
nand U6885 (N_6885,N_6353,N_6512);
xor U6886 (N_6886,N_6580,N_6471);
and U6887 (N_6887,N_6476,N_6472);
nor U6888 (N_6888,N_6430,N_6526);
and U6889 (N_6889,N_6359,N_6348);
or U6890 (N_6890,N_6594,N_6327);
and U6891 (N_6891,N_6506,N_6304);
nand U6892 (N_6892,N_6445,N_6558);
and U6893 (N_6893,N_6562,N_6316);
and U6894 (N_6894,N_6544,N_6354);
or U6895 (N_6895,N_6373,N_6405);
nand U6896 (N_6896,N_6545,N_6463);
nand U6897 (N_6897,N_6585,N_6399);
and U6898 (N_6898,N_6387,N_6505);
nand U6899 (N_6899,N_6460,N_6561);
and U6900 (N_6900,N_6664,N_6772);
xnor U6901 (N_6901,N_6693,N_6787);
xnor U6902 (N_6902,N_6609,N_6706);
nand U6903 (N_6903,N_6886,N_6845);
and U6904 (N_6904,N_6663,N_6839);
xor U6905 (N_6905,N_6615,N_6805);
xnor U6906 (N_6906,N_6876,N_6620);
and U6907 (N_6907,N_6846,N_6653);
or U6908 (N_6908,N_6822,N_6753);
or U6909 (N_6909,N_6742,N_6874);
nor U6910 (N_6910,N_6825,N_6868);
nor U6911 (N_6911,N_6789,N_6847);
or U6912 (N_6912,N_6679,N_6644);
nor U6913 (N_6913,N_6752,N_6866);
nand U6914 (N_6914,N_6818,N_6783);
or U6915 (N_6915,N_6600,N_6697);
xnor U6916 (N_6916,N_6833,N_6654);
or U6917 (N_6917,N_6638,N_6767);
xor U6918 (N_6918,N_6850,N_6680);
or U6919 (N_6919,N_6823,N_6899);
nor U6920 (N_6920,N_6834,N_6743);
nor U6921 (N_6921,N_6735,N_6729);
and U6922 (N_6922,N_6812,N_6619);
and U6923 (N_6923,N_6701,N_6746);
nor U6924 (N_6924,N_6696,N_6657);
nor U6925 (N_6925,N_6853,N_6763);
or U6926 (N_6926,N_6712,N_6618);
or U6927 (N_6927,N_6758,N_6625);
xnor U6928 (N_6928,N_6750,N_6608);
or U6929 (N_6929,N_6670,N_6708);
nand U6930 (N_6930,N_6762,N_6754);
nor U6931 (N_6931,N_6613,N_6793);
nand U6932 (N_6932,N_6830,N_6826);
nor U6933 (N_6933,N_6804,N_6809);
and U6934 (N_6934,N_6810,N_6678);
and U6935 (N_6935,N_6786,N_6666);
nand U6936 (N_6936,N_6884,N_6871);
and U6937 (N_6937,N_6689,N_6688);
and U6938 (N_6938,N_6860,N_6837);
nand U6939 (N_6939,N_6673,N_6864);
and U6940 (N_6940,N_6842,N_6617);
or U6941 (N_6941,N_6740,N_6623);
and U6942 (N_6942,N_6851,N_6637);
nor U6943 (N_6943,N_6709,N_6797);
or U6944 (N_6944,N_6677,N_6603);
and U6945 (N_6945,N_6785,N_6814);
and U6946 (N_6946,N_6643,N_6704);
nor U6947 (N_6947,N_6737,N_6776);
and U6948 (N_6948,N_6836,N_6628);
nand U6949 (N_6949,N_6824,N_6878);
xor U6950 (N_6950,N_6683,N_6872);
nor U6951 (N_6951,N_6734,N_6770);
and U6952 (N_6952,N_6832,N_6640);
nand U6953 (N_6953,N_6650,N_6621);
nand U6954 (N_6954,N_6759,N_6720);
nor U6955 (N_6955,N_6831,N_6893);
nor U6956 (N_6956,N_6710,N_6700);
xnor U6957 (N_6957,N_6724,N_6631);
nor U6958 (N_6958,N_6888,N_6791);
xnor U6959 (N_6959,N_6835,N_6633);
nor U6960 (N_6960,N_6726,N_6792);
nand U6961 (N_6961,N_6764,N_6869);
xnor U6962 (N_6962,N_6674,N_6801);
nor U6963 (N_6963,N_6802,N_6691);
or U6964 (N_6964,N_6757,N_6690);
nand U6965 (N_6965,N_6894,N_6799);
xor U6966 (N_6966,N_6605,N_6857);
xnor U6967 (N_6967,N_6741,N_6719);
and U6968 (N_6968,N_6703,N_6671);
or U6969 (N_6969,N_6736,N_6858);
and U6970 (N_6970,N_6747,N_6639);
nand U6971 (N_6971,N_6642,N_6612);
nand U6972 (N_6972,N_6755,N_6796);
xor U6973 (N_6973,N_6766,N_6879);
or U6974 (N_6974,N_6892,N_6775);
xnor U6975 (N_6975,N_6707,N_6685);
nand U6976 (N_6976,N_6744,N_6828);
nor U6977 (N_6977,N_6760,N_6658);
xnor U6978 (N_6978,N_6774,N_6800);
xnor U6979 (N_6979,N_6780,N_6607);
xor U6980 (N_6980,N_6610,N_6773);
nand U6981 (N_6981,N_6629,N_6897);
and U6982 (N_6982,N_6777,N_6635);
or U6983 (N_6983,N_6821,N_6636);
and U6984 (N_6984,N_6718,N_6651);
xor U6985 (N_6985,N_6855,N_6881);
nor U6986 (N_6986,N_6655,N_6732);
xor U6987 (N_6987,N_6728,N_6676);
xnor U6988 (N_6988,N_6725,N_6727);
xnor U6989 (N_6989,N_6748,N_6778);
nor U6990 (N_6990,N_6803,N_6795);
or U6991 (N_6991,N_6721,N_6813);
or U6992 (N_6992,N_6816,N_6820);
and U6993 (N_6993,N_6626,N_6875);
nand U6994 (N_6994,N_6854,N_6692);
and U6995 (N_6995,N_6715,N_6733);
xnor U6996 (N_6996,N_6705,N_6817);
xnor U6997 (N_6997,N_6684,N_6632);
xor U6998 (N_6998,N_6889,N_6861);
xor U6999 (N_6999,N_6849,N_6641);
xnor U7000 (N_7000,N_6867,N_6765);
or U7001 (N_7001,N_6856,N_6667);
xor U7002 (N_7002,N_6761,N_6604);
and U7003 (N_7003,N_6790,N_6843);
nor U7004 (N_7004,N_6859,N_6788);
nand U7005 (N_7005,N_6738,N_6771);
nor U7006 (N_7006,N_6716,N_6711);
nor U7007 (N_7007,N_6624,N_6882);
nor U7008 (N_7008,N_6756,N_6887);
xnor U7009 (N_7009,N_6781,N_6768);
or U7010 (N_7010,N_6769,N_6611);
nand U7011 (N_7011,N_6659,N_6616);
or U7012 (N_7012,N_6848,N_6687);
or U7013 (N_7013,N_6745,N_6806);
nand U7014 (N_7014,N_6895,N_6630);
or U7015 (N_7015,N_6896,N_6601);
and U7016 (N_7016,N_6827,N_6695);
nor U7017 (N_7017,N_6602,N_6713);
nand U7018 (N_7018,N_6751,N_6698);
and U7019 (N_7019,N_6782,N_6699);
and U7020 (N_7020,N_6808,N_6665);
or U7021 (N_7021,N_6870,N_6798);
nor U7022 (N_7022,N_6811,N_6686);
or U7023 (N_7023,N_6661,N_6898);
nor U7024 (N_7024,N_6873,N_6749);
nand U7025 (N_7025,N_6841,N_6645);
or U7026 (N_7026,N_6863,N_6669);
and U7027 (N_7027,N_6731,N_6862);
nor U7028 (N_7028,N_6794,N_6662);
xor U7029 (N_7029,N_6890,N_6722);
and U7030 (N_7030,N_6652,N_6660);
and U7031 (N_7031,N_6852,N_6681);
nor U7032 (N_7032,N_6675,N_6702);
or U7033 (N_7033,N_6891,N_6880);
nand U7034 (N_7034,N_6714,N_6829);
xnor U7035 (N_7035,N_6883,N_6648);
nand U7036 (N_7036,N_6885,N_6865);
or U7037 (N_7037,N_6656,N_6606);
nand U7038 (N_7038,N_6723,N_6649);
xor U7039 (N_7039,N_6739,N_6784);
or U7040 (N_7040,N_6672,N_6614);
nand U7041 (N_7041,N_6627,N_6682);
nand U7042 (N_7042,N_6717,N_6622);
nand U7043 (N_7043,N_6647,N_6877);
xor U7044 (N_7044,N_6807,N_6634);
and U7045 (N_7045,N_6694,N_6838);
and U7046 (N_7046,N_6819,N_6646);
nor U7047 (N_7047,N_6730,N_6779);
nand U7048 (N_7048,N_6844,N_6840);
nand U7049 (N_7049,N_6668,N_6815);
and U7050 (N_7050,N_6848,N_6617);
nor U7051 (N_7051,N_6761,N_6666);
and U7052 (N_7052,N_6634,N_6865);
or U7053 (N_7053,N_6775,N_6634);
and U7054 (N_7054,N_6625,N_6635);
nor U7055 (N_7055,N_6887,N_6729);
and U7056 (N_7056,N_6746,N_6690);
nor U7057 (N_7057,N_6717,N_6809);
nor U7058 (N_7058,N_6755,N_6724);
nor U7059 (N_7059,N_6649,N_6836);
or U7060 (N_7060,N_6690,N_6731);
nor U7061 (N_7061,N_6679,N_6784);
nor U7062 (N_7062,N_6788,N_6657);
or U7063 (N_7063,N_6866,N_6690);
nand U7064 (N_7064,N_6691,N_6603);
and U7065 (N_7065,N_6806,N_6853);
nor U7066 (N_7066,N_6865,N_6737);
nand U7067 (N_7067,N_6742,N_6659);
nor U7068 (N_7068,N_6888,N_6665);
and U7069 (N_7069,N_6664,N_6745);
nand U7070 (N_7070,N_6672,N_6624);
nand U7071 (N_7071,N_6640,N_6602);
nand U7072 (N_7072,N_6649,N_6780);
or U7073 (N_7073,N_6899,N_6781);
or U7074 (N_7074,N_6794,N_6717);
or U7075 (N_7075,N_6748,N_6765);
or U7076 (N_7076,N_6663,N_6833);
or U7077 (N_7077,N_6781,N_6712);
nand U7078 (N_7078,N_6801,N_6662);
nor U7079 (N_7079,N_6740,N_6895);
or U7080 (N_7080,N_6692,N_6832);
and U7081 (N_7081,N_6891,N_6687);
nand U7082 (N_7082,N_6728,N_6805);
and U7083 (N_7083,N_6637,N_6788);
nor U7084 (N_7084,N_6707,N_6636);
xnor U7085 (N_7085,N_6689,N_6763);
and U7086 (N_7086,N_6795,N_6750);
and U7087 (N_7087,N_6724,N_6702);
and U7088 (N_7088,N_6675,N_6643);
and U7089 (N_7089,N_6714,N_6675);
nand U7090 (N_7090,N_6842,N_6866);
nand U7091 (N_7091,N_6723,N_6635);
xor U7092 (N_7092,N_6816,N_6692);
or U7093 (N_7093,N_6896,N_6646);
and U7094 (N_7094,N_6845,N_6785);
nor U7095 (N_7095,N_6682,N_6634);
nand U7096 (N_7096,N_6600,N_6632);
nand U7097 (N_7097,N_6624,N_6868);
or U7098 (N_7098,N_6601,N_6698);
and U7099 (N_7099,N_6895,N_6858);
xnor U7100 (N_7100,N_6668,N_6679);
nand U7101 (N_7101,N_6617,N_6705);
nor U7102 (N_7102,N_6749,N_6816);
nor U7103 (N_7103,N_6612,N_6809);
nand U7104 (N_7104,N_6658,N_6683);
xor U7105 (N_7105,N_6896,N_6824);
or U7106 (N_7106,N_6646,N_6735);
nand U7107 (N_7107,N_6640,N_6632);
nand U7108 (N_7108,N_6829,N_6717);
or U7109 (N_7109,N_6734,N_6733);
xor U7110 (N_7110,N_6770,N_6670);
nand U7111 (N_7111,N_6801,N_6628);
nor U7112 (N_7112,N_6759,N_6631);
and U7113 (N_7113,N_6877,N_6762);
xor U7114 (N_7114,N_6670,N_6758);
nand U7115 (N_7115,N_6841,N_6858);
and U7116 (N_7116,N_6870,N_6681);
xor U7117 (N_7117,N_6824,N_6643);
and U7118 (N_7118,N_6857,N_6838);
nor U7119 (N_7119,N_6751,N_6703);
nand U7120 (N_7120,N_6658,N_6786);
and U7121 (N_7121,N_6745,N_6694);
or U7122 (N_7122,N_6644,N_6650);
and U7123 (N_7123,N_6687,N_6628);
xnor U7124 (N_7124,N_6855,N_6742);
and U7125 (N_7125,N_6868,N_6636);
or U7126 (N_7126,N_6894,N_6695);
and U7127 (N_7127,N_6726,N_6644);
nand U7128 (N_7128,N_6600,N_6628);
xnor U7129 (N_7129,N_6643,N_6758);
or U7130 (N_7130,N_6685,N_6810);
nand U7131 (N_7131,N_6761,N_6855);
nor U7132 (N_7132,N_6626,N_6782);
nor U7133 (N_7133,N_6680,N_6684);
and U7134 (N_7134,N_6823,N_6841);
and U7135 (N_7135,N_6733,N_6679);
nor U7136 (N_7136,N_6669,N_6872);
nand U7137 (N_7137,N_6813,N_6868);
xnor U7138 (N_7138,N_6810,N_6651);
nand U7139 (N_7139,N_6682,N_6857);
and U7140 (N_7140,N_6723,N_6693);
xor U7141 (N_7141,N_6660,N_6621);
nand U7142 (N_7142,N_6683,N_6824);
nand U7143 (N_7143,N_6761,N_6701);
nand U7144 (N_7144,N_6805,N_6842);
nor U7145 (N_7145,N_6822,N_6614);
nor U7146 (N_7146,N_6772,N_6890);
or U7147 (N_7147,N_6888,N_6771);
or U7148 (N_7148,N_6775,N_6860);
nor U7149 (N_7149,N_6831,N_6640);
or U7150 (N_7150,N_6658,N_6712);
xnor U7151 (N_7151,N_6779,N_6855);
nor U7152 (N_7152,N_6642,N_6772);
nor U7153 (N_7153,N_6704,N_6660);
and U7154 (N_7154,N_6707,N_6776);
or U7155 (N_7155,N_6672,N_6674);
or U7156 (N_7156,N_6674,N_6766);
xor U7157 (N_7157,N_6820,N_6649);
nor U7158 (N_7158,N_6732,N_6689);
and U7159 (N_7159,N_6655,N_6738);
and U7160 (N_7160,N_6669,N_6751);
nand U7161 (N_7161,N_6847,N_6753);
or U7162 (N_7162,N_6739,N_6664);
and U7163 (N_7163,N_6669,N_6776);
and U7164 (N_7164,N_6794,N_6673);
nor U7165 (N_7165,N_6770,N_6815);
nor U7166 (N_7166,N_6773,N_6659);
nor U7167 (N_7167,N_6699,N_6837);
xnor U7168 (N_7168,N_6731,N_6664);
nor U7169 (N_7169,N_6886,N_6743);
or U7170 (N_7170,N_6658,N_6704);
nor U7171 (N_7171,N_6810,N_6853);
or U7172 (N_7172,N_6780,N_6697);
nor U7173 (N_7173,N_6789,N_6636);
nand U7174 (N_7174,N_6688,N_6827);
nand U7175 (N_7175,N_6718,N_6662);
and U7176 (N_7176,N_6849,N_6699);
and U7177 (N_7177,N_6776,N_6722);
or U7178 (N_7178,N_6687,N_6751);
nor U7179 (N_7179,N_6760,N_6819);
xor U7180 (N_7180,N_6700,N_6632);
xor U7181 (N_7181,N_6875,N_6674);
or U7182 (N_7182,N_6864,N_6755);
nand U7183 (N_7183,N_6642,N_6614);
or U7184 (N_7184,N_6631,N_6718);
xnor U7185 (N_7185,N_6793,N_6871);
and U7186 (N_7186,N_6783,N_6774);
or U7187 (N_7187,N_6818,N_6813);
nor U7188 (N_7188,N_6844,N_6839);
nor U7189 (N_7189,N_6666,N_6815);
xor U7190 (N_7190,N_6786,N_6686);
nand U7191 (N_7191,N_6731,N_6889);
nand U7192 (N_7192,N_6781,N_6821);
or U7193 (N_7193,N_6810,N_6829);
nor U7194 (N_7194,N_6741,N_6756);
and U7195 (N_7195,N_6738,N_6797);
nor U7196 (N_7196,N_6825,N_6831);
xnor U7197 (N_7197,N_6882,N_6828);
xor U7198 (N_7198,N_6680,N_6757);
and U7199 (N_7199,N_6610,N_6734);
nor U7200 (N_7200,N_6946,N_7114);
or U7201 (N_7201,N_7093,N_7113);
nand U7202 (N_7202,N_7111,N_7035);
or U7203 (N_7203,N_6921,N_7049);
and U7204 (N_7204,N_6962,N_7105);
or U7205 (N_7205,N_7032,N_7086);
nor U7206 (N_7206,N_7197,N_7062);
nor U7207 (N_7207,N_6908,N_7104);
xor U7208 (N_7208,N_7112,N_6958);
nand U7209 (N_7209,N_7120,N_6941);
nand U7210 (N_7210,N_7024,N_7136);
nand U7211 (N_7211,N_6910,N_7056);
or U7212 (N_7212,N_6943,N_7174);
nor U7213 (N_7213,N_7155,N_7045);
nor U7214 (N_7214,N_7154,N_7029);
nor U7215 (N_7215,N_7166,N_7100);
or U7216 (N_7216,N_6956,N_6952);
nor U7217 (N_7217,N_7143,N_6965);
nand U7218 (N_7218,N_6901,N_6909);
nand U7219 (N_7219,N_6976,N_6996);
nand U7220 (N_7220,N_7025,N_7134);
nand U7221 (N_7221,N_7193,N_7194);
nor U7222 (N_7222,N_7168,N_7021);
and U7223 (N_7223,N_7043,N_7140);
and U7224 (N_7224,N_7198,N_6940);
and U7225 (N_7225,N_7087,N_7098);
xnor U7226 (N_7226,N_7047,N_7102);
and U7227 (N_7227,N_7195,N_7191);
nor U7228 (N_7228,N_6988,N_6973);
or U7229 (N_7229,N_7141,N_7122);
or U7230 (N_7230,N_7097,N_7108);
and U7231 (N_7231,N_7146,N_7132);
nand U7232 (N_7232,N_6948,N_6925);
nor U7233 (N_7233,N_7152,N_6954);
or U7234 (N_7234,N_7026,N_7013);
and U7235 (N_7235,N_6918,N_7088);
or U7236 (N_7236,N_7075,N_7060);
or U7237 (N_7237,N_6907,N_7116);
nand U7238 (N_7238,N_7038,N_7145);
nor U7239 (N_7239,N_7007,N_7138);
xor U7240 (N_7240,N_7040,N_7095);
nand U7241 (N_7241,N_7149,N_6972);
nand U7242 (N_7242,N_7142,N_7018);
and U7243 (N_7243,N_6969,N_7171);
nor U7244 (N_7244,N_7080,N_6916);
nand U7245 (N_7245,N_7002,N_7096);
nor U7246 (N_7246,N_6905,N_7044);
nor U7247 (N_7247,N_6906,N_6938);
and U7248 (N_7248,N_7169,N_7031);
and U7249 (N_7249,N_7127,N_7067);
nand U7250 (N_7250,N_7058,N_7020);
nand U7251 (N_7251,N_7010,N_7066);
nor U7252 (N_7252,N_7054,N_6902);
nor U7253 (N_7253,N_6937,N_6917);
xnor U7254 (N_7254,N_7070,N_7071);
nand U7255 (N_7255,N_7009,N_6977);
or U7256 (N_7256,N_7180,N_6992);
and U7257 (N_7257,N_7139,N_7089);
or U7258 (N_7258,N_7034,N_6953);
or U7259 (N_7259,N_7176,N_7137);
nand U7260 (N_7260,N_6914,N_6928);
and U7261 (N_7261,N_7012,N_7161);
and U7262 (N_7262,N_6951,N_6944);
and U7263 (N_7263,N_6990,N_6987);
nor U7264 (N_7264,N_6945,N_7053);
nand U7265 (N_7265,N_7153,N_6927);
and U7266 (N_7266,N_7182,N_7084);
nand U7267 (N_7267,N_7051,N_7017);
nand U7268 (N_7268,N_7189,N_6959);
or U7269 (N_7269,N_7039,N_7046);
nor U7270 (N_7270,N_7186,N_6998);
nand U7271 (N_7271,N_7094,N_7006);
nor U7272 (N_7272,N_7076,N_6995);
nand U7273 (N_7273,N_7181,N_7109);
xor U7274 (N_7274,N_7055,N_6904);
or U7275 (N_7275,N_7023,N_6971);
nand U7276 (N_7276,N_7150,N_7099);
nor U7277 (N_7277,N_6915,N_6966);
nor U7278 (N_7278,N_7052,N_6933);
nand U7279 (N_7279,N_6967,N_6935);
and U7280 (N_7280,N_6981,N_7185);
or U7281 (N_7281,N_7011,N_7057);
nor U7282 (N_7282,N_6930,N_7144);
or U7283 (N_7283,N_7178,N_7077);
nor U7284 (N_7284,N_6903,N_6994);
xnor U7285 (N_7285,N_7172,N_7179);
xor U7286 (N_7286,N_7110,N_6932);
nor U7287 (N_7287,N_6957,N_7048);
and U7288 (N_7288,N_6961,N_7175);
xor U7289 (N_7289,N_7027,N_7064);
nor U7290 (N_7290,N_7003,N_7158);
nand U7291 (N_7291,N_6968,N_7117);
and U7292 (N_7292,N_7118,N_7000);
nand U7293 (N_7293,N_7129,N_7033);
xor U7294 (N_7294,N_7173,N_7082);
and U7295 (N_7295,N_7123,N_7078);
nor U7296 (N_7296,N_6931,N_7106);
or U7297 (N_7297,N_7041,N_6984);
nor U7298 (N_7298,N_6991,N_6964);
xnor U7299 (N_7299,N_7091,N_7159);
nand U7300 (N_7300,N_6942,N_6983);
xor U7301 (N_7301,N_6974,N_7036);
nor U7302 (N_7302,N_7190,N_7119);
xnor U7303 (N_7303,N_7059,N_7103);
xor U7304 (N_7304,N_7028,N_7184);
or U7305 (N_7305,N_6980,N_6950);
and U7306 (N_7306,N_6947,N_7073);
nor U7307 (N_7307,N_7163,N_6929);
or U7308 (N_7308,N_6923,N_6985);
nand U7309 (N_7309,N_7125,N_6936);
or U7310 (N_7310,N_6949,N_7037);
nor U7311 (N_7311,N_6986,N_7107);
and U7312 (N_7312,N_7085,N_7121);
and U7313 (N_7313,N_7074,N_7005);
xor U7314 (N_7314,N_6920,N_6911);
nand U7315 (N_7315,N_7126,N_6926);
xnor U7316 (N_7316,N_7157,N_6989);
nor U7317 (N_7317,N_6978,N_7050);
nand U7318 (N_7318,N_7188,N_7196);
xor U7319 (N_7319,N_7156,N_6975);
nand U7320 (N_7320,N_7081,N_6900);
nor U7321 (N_7321,N_6960,N_7199);
nand U7322 (N_7322,N_7115,N_7160);
xnor U7323 (N_7323,N_6963,N_7042);
and U7324 (N_7324,N_6922,N_6919);
or U7325 (N_7325,N_6982,N_7004);
xor U7326 (N_7326,N_7162,N_6912);
xor U7327 (N_7327,N_7015,N_7092);
nand U7328 (N_7328,N_7177,N_7090);
and U7329 (N_7329,N_7065,N_7030);
or U7330 (N_7330,N_7133,N_6924);
or U7331 (N_7331,N_7147,N_7187);
nor U7332 (N_7332,N_7130,N_7061);
xnor U7333 (N_7333,N_7183,N_7069);
or U7334 (N_7334,N_7101,N_7164);
or U7335 (N_7335,N_7063,N_7124);
or U7336 (N_7336,N_7008,N_6970);
nor U7337 (N_7337,N_7131,N_7192);
and U7338 (N_7338,N_6939,N_6993);
nand U7339 (N_7339,N_7001,N_6999);
nor U7340 (N_7340,N_7068,N_7072);
and U7341 (N_7341,N_7022,N_6913);
xor U7342 (N_7342,N_6934,N_6979);
nor U7343 (N_7343,N_7165,N_6997);
xnor U7344 (N_7344,N_7148,N_7079);
nand U7345 (N_7345,N_7083,N_6955);
nor U7346 (N_7346,N_7167,N_7019);
and U7347 (N_7347,N_7135,N_7170);
or U7348 (N_7348,N_7128,N_7151);
and U7349 (N_7349,N_7014,N_7016);
xnor U7350 (N_7350,N_6917,N_7171);
xnor U7351 (N_7351,N_7017,N_6915);
nor U7352 (N_7352,N_7086,N_6998);
and U7353 (N_7353,N_6960,N_7197);
nor U7354 (N_7354,N_6902,N_6961);
xor U7355 (N_7355,N_6999,N_6915);
or U7356 (N_7356,N_7165,N_7185);
and U7357 (N_7357,N_7115,N_7012);
nor U7358 (N_7358,N_7167,N_7024);
nand U7359 (N_7359,N_7188,N_6953);
and U7360 (N_7360,N_7027,N_7070);
or U7361 (N_7361,N_7043,N_7034);
xnor U7362 (N_7362,N_7025,N_7179);
xor U7363 (N_7363,N_7198,N_7076);
nor U7364 (N_7364,N_7060,N_7107);
nand U7365 (N_7365,N_7069,N_6903);
or U7366 (N_7366,N_6964,N_6987);
and U7367 (N_7367,N_7155,N_7085);
xnor U7368 (N_7368,N_7131,N_7121);
or U7369 (N_7369,N_7167,N_7072);
nand U7370 (N_7370,N_7186,N_7083);
and U7371 (N_7371,N_7127,N_7191);
nand U7372 (N_7372,N_7044,N_7077);
nand U7373 (N_7373,N_7130,N_7044);
or U7374 (N_7374,N_7141,N_7035);
nand U7375 (N_7375,N_7170,N_7143);
nand U7376 (N_7376,N_7118,N_7071);
nand U7377 (N_7377,N_7196,N_7171);
and U7378 (N_7378,N_7103,N_6969);
or U7379 (N_7379,N_6937,N_6936);
xnor U7380 (N_7380,N_7156,N_7176);
nand U7381 (N_7381,N_7124,N_7131);
nand U7382 (N_7382,N_7002,N_7072);
or U7383 (N_7383,N_7024,N_6985);
xor U7384 (N_7384,N_7154,N_6970);
or U7385 (N_7385,N_7104,N_6913);
nor U7386 (N_7386,N_6976,N_7136);
or U7387 (N_7387,N_7079,N_6970);
and U7388 (N_7388,N_6962,N_7026);
and U7389 (N_7389,N_6926,N_7104);
nor U7390 (N_7390,N_7030,N_6998);
xnor U7391 (N_7391,N_7091,N_7092);
or U7392 (N_7392,N_7060,N_7135);
and U7393 (N_7393,N_7108,N_6908);
nor U7394 (N_7394,N_6980,N_6947);
nand U7395 (N_7395,N_7129,N_7141);
or U7396 (N_7396,N_6931,N_6947);
nand U7397 (N_7397,N_7052,N_7166);
or U7398 (N_7398,N_6909,N_7138);
and U7399 (N_7399,N_7122,N_7029);
nor U7400 (N_7400,N_6932,N_7035);
nor U7401 (N_7401,N_7190,N_7121);
and U7402 (N_7402,N_7162,N_7131);
nand U7403 (N_7403,N_6910,N_7119);
xnor U7404 (N_7404,N_7065,N_7097);
or U7405 (N_7405,N_6914,N_6913);
xor U7406 (N_7406,N_6935,N_7103);
and U7407 (N_7407,N_6946,N_6933);
xnor U7408 (N_7408,N_6967,N_7055);
nor U7409 (N_7409,N_7115,N_7164);
nand U7410 (N_7410,N_7196,N_6998);
and U7411 (N_7411,N_6995,N_6965);
and U7412 (N_7412,N_7079,N_7027);
xnor U7413 (N_7413,N_6919,N_6928);
and U7414 (N_7414,N_7000,N_7036);
nand U7415 (N_7415,N_6960,N_7055);
nor U7416 (N_7416,N_6974,N_7181);
nor U7417 (N_7417,N_7147,N_7076);
or U7418 (N_7418,N_7137,N_7002);
and U7419 (N_7419,N_6935,N_6972);
nand U7420 (N_7420,N_7194,N_6925);
nor U7421 (N_7421,N_7122,N_7175);
nor U7422 (N_7422,N_7103,N_6964);
xor U7423 (N_7423,N_7075,N_7034);
xor U7424 (N_7424,N_7065,N_7053);
nor U7425 (N_7425,N_7157,N_7022);
and U7426 (N_7426,N_7109,N_7035);
nor U7427 (N_7427,N_7159,N_6972);
nand U7428 (N_7428,N_6955,N_6975);
nand U7429 (N_7429,N_7155,N_7044);
or U7430 (N_7430,N_7043,N_7036);
or U7431 (N_7431,N_6903,N_6941);
or U7432 (N_7432,N_7049,N_6933);
or U7433 (N_7433,N_7072,N_7149);
or U7434 (N_7434,N_7155,N_7114);
nand U7435 (N_7435,N_7009,N_6945);
or U7436 (N_7436,N_7018,N_6968);
and U7437 (N_7437,N_6998,N_6928);
xnor U7438 (N_7438,N_6953,N_7176);
and U7439 (N_7439,N_7169,N_7111);
xnor U7440 (N_7440,N_7025,N_6972);
or U7441 (N_7441,N_7093,N_7183);
nand U7442 (N_7442,N_6979,N_6965);
and U7443 (N_7443,N_6985,N_6922);
nand U7444 (N_7444,N_6939,N_7059);
xnor U7445 (N_7445,N_7165,N_7073);
or U7446 (N_7446,N_7030,N_6985);
or U7447 (N_7447,N_7103,N_7053);
xnor U7448 (N_7448,N_7187,N_6909);
nor U7449 (N_7449,N_7012,N_6959);
nand U7450 (N_7450,N_7131,N_7073);
xor U7451 (N_7451,N_7008,N_7034);
or U7452 (N_7452,N_7169,N_6914);
or U7453 (N_7453,N_6929,N_7087);
and U7454 (N_7454,N_6988,N_6901);
nand U7455 (N_7455,N_6995,N_7034);
nand U7456 (N_7456,N_7061,N_7133);
nand U7457 (N_7457,N_6914,N_7173);
nor U7458 (N_7458,N_7071,N_7150);
nor U7459 (N_7459,N_7143,N_7135);
nand U7460 (N_7460,N_7073,N_7036);
nand U7461 (N_7461,N_7121,N_6985);
nand U7462 (N_7462,N_7185,N_7177);
nand U7463 (N_7463,N_7173,N_7045);
nand U7464 (N_7464,N_6937,N_6945);
nand U7465 (N_7465,N_6989,N_7099);
nor U7466 (N_7466,N_7021,N_7029);
nand U7467 (N_7467,N_6927,N_7109);
xor U7468 (N_7468,N_7008,N_7074);
xor U7469 (N_7469,N_7011,N_7178);
and U7470 (N_7470,N_7173,N_7063);
or U7471 (N_7471,N_6935,N_6928);
nand U7472 (N_7472,N_6911,N_7031);
or U7473 (N_7473,N_6907,N_7195);
or U7474 (N_7474,N_6953,N_6920);
and U7475 (N_7475,N_7087,N_7082);
nor U7476 (N_7476,N_7008,N_6951);
nand U7477 (N_7477,N_7042,N_7039);
and U7478 (N_7478,N_6953,N_7103);
or U7479 (N_7479,N_7160,N_7063);
or U7480 (N_7480,N_6997,N_6929);
and U7481 (N_7481,N_7004,N_7036);
or U7482 (N_7482,N_6910,N_7092);
xnor U7483 (N_7483,N_7099,N_7061);
and U7484 (N_7484,N_7017,N_7070);
xnor U7485 (N_7485,N_7025,N_7171);
nor U7486 (N_7486,N_6924,N_7000);
nand U7487 (N_7487,N_7109,N_6929);
and U7488 (N_7488,N_7065,N_7034);
nand U7489 (N_7489,N_7121,N_7084);
nor U7490 (N_7490,N_7009,N_6916);
and U7491 (N_7491,N_7112,N_6912);
xnor U7492 (N_7492,N_6989,N_6967);
xnor U7493 (N_7493,N_7068,N_7111);
and U7494 (N_7494,N_7171,N_7163);
nand U7495 (N_7495,N_7122,N_7181);
and U7496 (N_7496,N_7047,N_6900);
nand U7497 (N_7497,N_7134,N_6907);
nor U7498 (N_7498,N_6947,N_7083);
nor U7499 (N_7499,N_6969,N_7155);
and U7500 (N_7500,N_7279,N_7433);
nand U7501 (N_7501,N_7221,N_7378);
and U7502 (N_7502,N_7216,N_7390);
xor U7503 (N_7503,N_7213,N_7244);
nand U7504 (N_7504,N_7264,N_7370);
xor U7505 (N_7505,N_7401,N_7234);
nand U7506 (N_7506,N_7203,N_7439);
and U7507 (N_7507,N_7325,N_7349);
and U7508 (N_7508,N_7223,N_7200);
and U7509 (N_7509,N_7313,N_7407);
or U7510 (N_7510,N_7317,N_7487);
and U7511 (N_7511,N_7278,N_7478);
xor U7512 (N_7512,N_7410,N_7385);
or U7513 (N_7513,N_7287,N_7379);
xor U7514 (N_7514,N_7217,N_7432);
and U7515 (N_7515,N_7483,N_7323);
nor U7516 (N_7516,N_7292,N_7434);
nand U7517 (N_7517,N_7399,N_7276);
and U7518 (N_7518,N_7305,N_7335);
xnor U7519 (N_7519,N_7319,N_7242);
and U7520 (N_7520,N_7492,N_7255);
nor U7521 (N_7521,N_7253,N_7333);
or U7522 (N_7522,N_7398,N_7228);
nand U7523 (N_7523,N_7306,N_7374);
nor U7524 (N_7524,N_7286,N_7201);
or U7525 (N_7525,N_7329,N_7465);
nand U7526 (N_7526,N_7263,N_7428);
nor U7527 (N_7527,N_7405,N_7402);
or U7528 (N_7528,N_7260,N_7283);
or U7529 (N_7529,N_7373,N_7249);
nand U7530 (N_7530,N_7484,N_7215);
or U7531 (N_7531,N_7489,N_7365);
nand U7532 (N_7532,N_7209,N_7359);
nor U7533 (N_7533,N_7426,N_7411);
nor U7534 (N_7534,N_7392,N_7207);
nor U7535 (N_7535,N_7372,N_7477);
nand U7536 (N_7536,N_7262,N_7346);
or U7537 (N_7537,N_7290,N_7357);
and U7538 (N_7538,N_7413,N_7336);
nor U7539 (N_7539,N_7225,N_7499);
xnor U7540 (N_7540,N_7285,N_7224);
nand U7541 (N_7541,N_7204,N_7471);
xnor U7542 (N_7542,N_7376,N_7414);
and U7543 (N_7543,N_7348,N_7269);
and U7544 (N_7544,N_7397,N_7481);
or U7545 (N_7545,N_7396,N_7364);
or U7546 (N_7546,N_7496,N_7356);
xnor U7547 (N_7547,N_7441,N_7450);
and U7548 (N_7548,N_7476,N_7408);
and U7549 (N_7549,N_7246,N_7380);
xnor U7550 (N_7550,N_7424,N_7486);
nand U7551 (N_7551,N_7247,N_7237);
nor U7552 (N_7552,N_7475,N_7321);
nand U7553 (N_7553,N_7420,N_7241);
and U7554 (N_7554,N_7493,N_7377);
and U7555 (N_7555,N_7256,N_7482);
xor U7556 (N_7556,N_7238,N_7363);
nor U7557 (N_7557,N_7274,N_7498);
nor U7558 (N_7558,N_7316,N_7229);
nand U7559 (N_7559,N_7231,N_7354);
nand U7560 (N_7560,N_7448,N_7344);
xnor U7561 (N_7561,N_7400,N_7425);
nand U7562 (N_7562,N_7341,N_7446);
and U7563 (N_7563,N_7350,N_7409);
xnor U7564 (N_7564,N_7435,N_7273);
and U7565 (N_7565,N_7314,N_7371);
or U7566 (N_7566,N_7230,N_7308);
nand U7567 (N_7567,N_7296,N_7497);
xor U7568 (N_7568,N_7267,N_7208);
xor U7569 (N_7569,N_7464,N_7239);
and U7570 (N_7570,N_7459,N_7445);
nand U7571 (N_7571,N_7252,N_7270);
or U7572 (N_7572,N_7266,N_7220);
nand U7573 (N_7573,N_7418,N_7383);
and U7574 (N_7574,N_7210,N_7447);
or U7575 (N_7575,N_7494,N_7381);
or U7576 (N_7576,N_7312,N_7258);
xnor U7577 (N_7577,N_7389,N_7265);
nor U7578 (N_7578,N_7332,N_7452);
and U7579 (N_7579,N_7340,N_7275);
or U7580 (N_7580,N_7235,N_7394);
xor U7581 (N_7581,N_7470,N_7416);
nand U7582 (N_7582,N_7358,N_7236);
nor U7583 (N_7583,N_7437,N_7485);
nor U7584 (N_7584,N_7472,N_7315);
xor U7585 (N_7585,N_7423,N_7490);
or U7586 (N_7586,N_7431,N_7355);
nand U7587 (N_7587,N_7303,N_7387);
nand U7588 (N_7588,N_7466,N_7386);
and U7589 (N_7589,N_7328,N_7330);
or U7590 (N_7590,N_7284,N_7421);
or U7591 (N_7591,N_7429,N_7298);
nand U7592 (N_7592,N_7320,N_7360);
or U7593 (N_7593,N_7302,N_7388);
nor U7594 (N_7594,N_7419,N_7310);
or U7595 (N_7595,N_7226,N_7214);
and U7596 (N_7596,N_7261,N_7361);
xor U7597 (N_7597,N_7322,N_7455);
nor U7598 (N_7598,N_7288,N_7307);
or U7599 (N_7599,N_7282,N_7259);
nor U7600 (N_7600,N_7347,N_7289);
or U7601 (N_7601,N_7440,N_7339);
and U7602 (N_7602,N_7248,N_7473);
nand U7603 (N_7603,N_7222,N_7211);
xor U7604 (N_7604,N_7458,N_7393);
xnor U7605 (N_7605,N_7301,N_7353);
and U7606 (N_7606,N_7495,N_7311);
nand U7607 (N_7607,N_7362,N_7254);
xor U7608 (N_7608,N_7243,N_7338);
nor U7609 (N_7609,N_7300,N_7369);
or U7610 (N_7610,N_7295,N_7436);
nor U7611 (N_7611,N_7460,N_7251);
or U7612 (N_7612,N_7212,N_7304);
xnor U7613 (N_7613,N_7384,N_7294);
and U7614 (N_7614,N_7309,N_7271);
nor U7615 (N_7615,N_7293,N_7202);
xor U7616 (N_7616,N_7240,N_7206);
nor U7617 (N_7617,N_7272,N_7351);
and U7618 (N_7618,N_7451,N_7327);
xor U7619 (N_7619,N_7250,N_7467);
xnor U7620 (N_7620,N_7427,N_7219);
or U7621 (N_7621,N_7479,N_7257);
nor U7622 (N_7622,N_7366,N_7461);
xnor U7623 (N_7623,N_7233,N_7412);
nand U7624 (N_7624,N_7342,N_7218);
nand U7625 (N_7625,N_7277,N_7324);
and U7626 (N_7626,N_7417,N_7331);
nand U7627 (N_7627,N_7291,N_7375);
nor U7628 (N_7628,N_7343,N_7456);
and U7629 (N_7629,N_7345,N_7444);
or U7630 (N_7630,N_7453,N_7454);
xnor U7631 (N_7631,N_7403,N_7391);
nor U7632 (N_7632,N_7299,N_7367);
or U7633 (N_7633,N_7268,N_7480);
nand U7634 (N_7634,N_7457,N_7469);
nand U7635 (N_7635,N_7438,N_7449);
nand U7636 (N_7636,N_7281,N_7462);
nor U7637 (N_7637,N_7245,N_7488);
or U7638 (N_7638,N_7368,N_7415);
nor U7639 (N_7639,N_7280,N_7442);
nor U7640 (N_7640,N_7227,N_7463);
xnor U7641 (N_7641,N_7382,N_7334);
and U7642 (N_7642,N_7443,N_7352);
nand U7643 (N_7643,N_7337,N_7205);
xnor U7644 (N_7644,N_7430,N_7395);
or U7645 (N_7645,N_7318,N_7422);
or U7646 (N_7646,N_7232,N_7404);
xor U7647 (N_7647,N_7474,N_7491);
nand U7648 (N_7648,N_7406,N_7326);
nand U7649 (N_7649,N_7468,N_7297);
or U7650 (N_7650,N_7436,N_7357);
nand U7651 (N_7651,N_7391,N_7331);
or U7652 (N_7652,N_7342,N_7458);
and U7653 (N_7653,N_7381,N_7308);
or U7654 (N_7654,N_7217,N_7336);
or U7655 (N_7655,N_7422,N_7273);
xnor U7656 (N_7656,N_7208,N_7313);
nor U7657 (N_7657,N_7496,N_7455);
nor U7658 (N_7658,N_7366,N_7207);
nor U7659 (N_7659,N_7299,N_7431);
nand U7660 (N_7660,N_7249,N_7284);
nor U7661 (N_7661,N_7214,N_7358);
xnor U7662 (N_7662,N_7208,N_7210);
or U7663 (N_7663,N_7229,N_7459);
and U7664 (N_7664,N_7377,N_7335);
nor U7665 (N_7665,N_7482,N_7249);
xor U7666 (N_7666,N_7458,N_7322);
and U7667 (N_7667,N_7210,N_7299);
nand U7668 (N_7668,N_7295,N_7415);
or U7669 (N_7669,N_7292,N_7498);
or U7670 (N_7670,N_7333,N_7360);
nor U7671 (N_7671,N_7277,N_7487);
nand U7672 (N_7672,N_7340,N_7242);
and U7673 (N_7673,N_7423,N_7412);
and U7674 (N_7674,N_7362,N_7404);
or U7675 (N_7675,N_7494,N_7206);
xor U7676 (N_7676,N_7498,N_7373);
and U7677 (N_7677,N_7209,N_7409);
or U7678 (N_7678,N_7412,N_7495);
nor U7679 (N_7679,N_7486,N_7321);
nor U7680 (N_7680,N_7318,N_7241);
nand U7681 (N_7681,N_7285,N_7274);
xnor U7682 (N_7682,N_7329,N_7354);
or U7683 (N_7683,N_7289,N_7209);
and U7684 (N_7684,N_7370,N_7205);
nor U7685 (N_7685,N_7269,N_7374);
and U7686 (N_7686,N_7468,N_7465);
or U7687 (N_7687,N_7395,N_7345);
xor U7688 (N_7688,N_7330,N_7290);
xnor U7689 (N_7689,N_7491,N_7310);
nor U7690 (N_7690,N_7210,N_7342);
xnor U7691 (N_7691,N_7372,N_7336);
xor U7692 (N_7692,N_7455,N_7253);
xor U7693 (N_7693,N_7225,N_7303);
nor U7694 (N_7694,N_7456,N_7367);
nand U7695 (N_7695,N_7494,N_7256);
and U7696 (N_7696,N_7482,N_7440);
and U7697 (N_7697,N_7405,N_7365);
or U7698 (N_7698,N_7403,N_7277);
nand U7699 (N_7699,N_7268,N_7309);
and U7700 (N_7700,N_7437,N_7458);
xnor U7701 (N_7701,N_7498,N_7468);
xor U7702 (N_7702,N_7436,N_7394);
nand U7703 (N_7703,N_7406,N_7394);
or U7704 (N_7704,N_7349,N_7215);
nor U7705 (N_7705,N_7224,N_7376);
nor U7706 (N_7706,N_7215,N_7231);
xnor U7707 (N_7707,N_7221,N_7244);
nand U7708 (N_7708,N_7499,N_7240);
nand U7709 (N_7709,N_7471,N_7282);
nand U7710 (N_7710,N_7406,N_7369);
xnor U7711 (N_7711,N_7394,N_7390);
xor U7712 (N_7712,N_7221,N_7414);
nor U7713 (N_7713,N_7226,N_7418);
nor U7714 (N_7714,N_7215,N_7305);
nand U7715 (N_7715,N_7364,N_7295);
or U7716 (N_7716,N_7347,N_7491);
or U7717 (N_7717,N_7410,N_7423);
or U7718 (N_7718,N_7277,N_7427);
or U7719 (N_7719,N_7211,N_7372);
or U7720 (N_7720,N_7279,N_7417);
or U7721 (N_7721,N_7252,N_7313);
and U7722 (N_7722,N_7406,N_7347);
and U7723 (N_7723,N_7329,N_7421);
nand U7724 (N_7724,N_7346,N_7354);
nor U7725 (N_7725,N_7326,N_7338);
and U7726 (N_7726,N_7475,N_7431);
and U7727 (N_7727,N_7254,N_7418);
or U7728 (N_7728,N_7384,N_7299);
nor U7729 (N_7729,N_7356,N_7297);
xor U7730 (N_7730,N_7284,N_7346);
and U7731 (N_7731,N_7368,N_7409);
or U7732 (N_7732,N_7296,N_7454);
nand U7733 (N_7733,N_7399,N_7394);
and U7734 (N_7734,N_7421,N_7377);
nand U7735 (N_7735,N_7257,N_7407);
nand U7736 (N_7736,N_7217,N_7409);
xor U7737 (N_7737,N_7234,N_7392);
or U7738 (N_7738,N_7290,N_7430);
xnor U7739 (N_7739,N_7368,N_7259);
and U7740 (N_7740,N_7267,N_7236);
xor U7741 (N_7741,N_7355,N_7423);
xnor U7742 (N_7742,N_7445,N_7289);
nand U7743 (N_7743,N_7284,N_7318);
nand U7744 (N_7744,N_7372,N_7297);
xnor U7745 (N_7745,N_7283,N_7289);
and U7746 (N_7746,N_7399,N_7420);
nand U7747 (N_7747,N_7238,N_7446);
and U7748 (N_7748,N_7404,N_7408);
xnor U7749 (N_7749,N_7391,N_7317);
and U7750 (N_7750,N_7261,N_7389);
nor U7751 (N_7751,N_7428,N_7446);
nand U7752 (N_7752,N_7288,N_7272);
or U7753 (N_7753,N_7205,N_7332);
xor U7754 (N_7754,N_7482,N_7235);
and U7755 (N_7755,N_7440,N_7296);
xor U7756 (N_7756,N_7367,N_7494);
nand U7757 (N_7757,N_7440,N_7479);
and U7758 (N_7758,N_7230,N_7410);
xnor U7759 (N_7759,N_7429,N_7297);
and U7760 (N_7760,N_7262,N_7439);
and U7761 (N_7761,N_7258,N_7231);
nand U7762 (N_7762,N_7278,N_7485);
and U7763 (N_7763,N_7493,N_7396);
nor U7764 (N_7764,N_7335,N_7381);
xnor U7765 (N_7765,N_7496,N_7221);
xor U7766 (N_7766,N_7308,N_7370);
nor U7767 (N_7767,N_7429,N_7432);
xor U7768 (N_7768,N_7330,N_7474);
nand U7769 (N_7769,N_7208,N_7379);
nor U7770 (N_7770,N_7470,N_7468);
xor U7771 (N_7771,N_7299,N_7425);
and U7772 (N_7772,N_7412,N_7254);
xor U7773 (N_7773,N_7375,N_7488);
xnor U7774 (N_7774,N_7204,N_7364);
or U7775 (N_7775,N_7242,N_7499);
and U7776 (N_7776,N_7490,N_7465);
or U7777 (N_7777,N_7234,N_7444);
or U7778 (N_7778,N_7311,N_7226);
nand U7779 (N_7779,N_7361,N_7426);
or U7780 (N_7780,N_7227,N_7374);
xnor U7781 (N_7781,N_7284,N_7237);
xnor U7782 (N_7782,N_7498,N_7417);
xor U7783 (N_7783,N_7334,N_7437);
xnor U7784 (N_7784,N_7247,N_7203);
and U7785 (N_7785,N_7388,N_7295);
or U7786 (N_7786,N_7375,N_7349);
xnor U7787 (N_7787,N_7378,N_7230);
or U7788 (N_7788,N_7415,N_7251);
xor U7789 (N_7789,N_7339,N_7487);
or U7790 (N_7790,N_7442,N_7348);
or U7791 (N_7791,N_7432,N_7420);
nor U7792 (N_7792,N_7296,N_7321);
or U7793 (N_7793,N_7316,N_7361);
or U7794 (N_7794,N_7252,N_7297);
nand U7795 (N_7795,N_7489,N_7372);
and U7796 (N_7796,N_7275,N_7390);
or U7797 (N_7797,N_7405,N_7269);
and U7798 (N_7798,N_7459,N_7461);
nor U7799 (N_7799,N_7288,N_7267);
or U7800 (N_7800,N_7766,N_7524);
or U7801 (N_7801,N_7688,N_7754);
or U7802 (N_7802,N_7619,N_7641);
and U7803 (N_7803,N_7677,N_7547);
and U7804 (N_7804,N_7546,N_7665);
nor U7805 (N_7805,N_7747,N_7722);
nor U7806 (N_7806,N_7519,N_7762);
nor U7807 (N_7807,N_7668,N_7724);
nor U7808 (N_7808,N_7718,N_7663);
nand U7809 (N_7809,N_7588,N_7582);
and U7810 (N_7810,N_7571,N_7504);
or U7811 (N_7811,N_7732,N_7567);
nand U7812 (N_7812,N_7760,N_7702);
and U7813 (N_7813,N_7520,N_7683);
nand U7814 (N_7814,N_7552,N_7703);
and U7815 (N_7815,N_7518,N_7787);
nand U7816 (N_7816,N_7507,N_7666);
and U7817 (N_7817,N_7799,N_7587);
xor U7818 (N_7818,N_7629,N_7778);
or U7819 (N_7819,N_7513,N_7605);
xnor U7820 (N_7820,N_7728,N_7651);
xor U7821 (N_7821,N_7646,N_7572);
nor U7822 (N_7822,N_7661,N_7624);
or U7823 (N_7823,N_7639,N_7773);
and U7824 (N_7824,N_7511,N_7537);
and U7825 (N_7825,N_7767,N_7670);
xor U7826 (N_7826,N_7725,N_7573);
xor U7827 (N_7827,N_7505,N_7752);
and U7828 (N_7828,N_7740,N_7649);
xor U7829 (N_7829,N_7554,N_7727);
or U7830 (N_7830,N_7786,N_7764);
and U7831 (N_7831,N_7769,N_7638);
nand U7832 (N_7832,N_7550,N_7656);
nor U7833 (N_7833,N_7788,N_7525);
nand U7834 (N_7834,N_7654,N_7535);
nand U7835 (N_7835,N_7763,N_7659);
nor U7836 (N_7836,N_7607,N_7575);
nand U7837 (N_7837,N_7642,N_7771);
xnor U7838 (N_7838,N_7791,N_7585);
nor U7839 (N_7839,N_7539,N_7509);
nor U7840 (N_7840,N_7751,N_7647);
nor U7841 (N_7841,N_7730,N_7700);
nand U7842 (N_7842,N_7528,N_7757);
or U7843 (N_7843,N_7570,N_7652);
nor U7844 (N_7844,N_7601,N_7704);
nor U7845 (N_7845,N_7542,N_7620);
or U7846 (N_7846,N_7614,N_7741);
and U7847 (N_7847,N_7779,N_7578);
nor U7848 (N_7848,N_7776,N_7560);
nand U7849 (N_7849,N_7521,N_7508);
or U7850 (N_7850,N_7758,N_7556);
or U7851 (N_7851,N_7631,N_7785);
nand U7852 (N_7852,N_7600,N_7723);
and U7853 (N_7853,N_7739,N_7711);
nor U7854 (N_7854,N_7783,N_7617);
xnor U7855 (N_7855,N_7549,N_7708);
xor U7856 (N_7856,N_7565,N_7709);
xnor U7857 (N_7857,N_7640,N_7583);
or U7858 (N_7858,N_7609,N_7584);
and U7859 (N_7859,N_7589,N_7742);
or U7860 (N_7860,N_7678,N_7695);
nor U7861 (N_7861,N_7653,N_7676);
nand U7862 (N_7862,N_7612,N_7595);
or U7863 (N_7863,N_7794,N_7645);
nand U7864 (N_7864,N_7627,N_7798);
and U7865 (N_7865,N_7777,N_7564);
and U7866 (N_7866,N_7768,N_7598);
or U7867 (N_7867,N_7710,N_7715);
and U7868 (N_7868,N_7544,N_7626);
xnor U7869 (N_7869,N_7574,N_7780);
nor U7870 (N_7870,N_7613,N_7749);
xor U7871 (N_7871,N_7632,N_7603);
and U7872 (N_7872,N_7596,N_7591);
and U7873 (N_7873,N_7781,N_7697);
xor U7874 (N_7874,N_7685,N_7658);
nand U7875 (N_7875,N_7608,N_7536);
or U7876 (N_7876,N_7716,N_7753);
xor U7877 (N_7877,N_7541,N_7784);
or U7878 (N_7878,N_7736,N_7743);
nor U7879 (N_7879,N_7623,N_7569);
and U7880 (N_7880,N_7579,N_7599);
nor U7881 (N_7881,N_7557,N_7737);
nand U7882 (N_7882,N_7755,N_7712);
xnor U7883 (N_7883,N_7705,N_7533);
and U7884 (N_7884,N_7506,N_7733);
and U7885 (N_7885,N_7706,N_7553);
nand U7886 (N_7886,N_7750,N_7782);
xor U7887 (N_7887,N_7684,N_7500);
nand U7888 (N_7888,N_7650,N_7673);
and U7889 (N_7889,N_7698,N_7622);
or U7890 (N_7890,N_7610,N_7693);
nor U7891 (N_7891,N_7746,N_7713);
nor U7892 (N_7892,N_7770,N_7721);
nand U7893 (N_7893,N_7534,N_7615);
xor U7894 (N_7894,N_7618,N_7674);
nor U7895 (N_7895,N_7526,N_7795);
nand U7896 (N_7896,N_7679,N_7566);
nor U7897 (N_7897,N_7562,N_7580);
nor U7898 (N_7898,N_7633,N_7761);
nor U7899 (N_7899,N_7682,N_7745);
nand U7900 (N_7900,N_7735,N_7555);
xnor U7901 (N_7901,N_7687,N_7616);
and U7902 (N_7902,N_7529,N_7694);
nand U7903 (N_7903,N_7717,N_7531);
and U7904 (N_7904,N_7561,N_7548);
nor U7905 (N_7905,N_7738,N_7581);
or U7906 (N_7906,N_7503,N_7686);
xor U7907 (N_7907,N_7611,N_7635);
nor U7908 (N_7908,N_7734,N_7680);
xnor U7909 (N_7909,N_7636,N_7563);
nand U7910 (N_7910,N_7793,N_7593);
and U7911 (N_7911,N_7558,N_7514);
nor U7912 (N_7912,N_7576,N_7691);
and U7913 (N_7913,N_7726,N_7775);
or U7914 (N_7914,N_7699,N_7523);
nand U7915 (N_7915,N_7594,N_7664);
xor U7916 (N_7916,N_7714,N_7696);
and U7917 (N_7917,N_7527,N_7621);
or U7918 (N_7918,N_7660,N_7644);
nor U7919 (N_7919,N_7648,N_7720);
xor U7920 (N_7920,N_7515,N_7796);
and U7921 (N_7921,N_7729,N_7592);
and U7922 (N_7922,N_7628,N_7671);
and U7923 (N_7923,N_7538,N_7790);
xnor U7924 (N_7924,N_7669,N_7744);
or U7925 (N_7925,N_7675,N_7667);
nand U7926 (N_7926,N_7637,N_7568);
nor U7927 (N_7927,N_7772,N_7543);
xor U7928 (N_7928,N_7662,N_7597);
xnor U7929 (N_7929,N_7797,N_7759);
nand U7930 (N_7930,N_7765,N_7690);
or U7931 (N_7931,N_7630,N_7551);
nor U7932 (N_7932,N_7792,N_7586);
nor U7933 (N_7933,N_7577,N_7545);
or U7934 (N_7934,N_7657,N_7774);
and U7935 (N_7935,N_7692,N_7501);
nor U7936 (N_7936,N_7789,N_7655);
nand U7937 (N_7937,N_7634,N_7512);
or U7938 (N_7938,N_7530,N_7719);
nand U7939 (N_7939,N_7701,N_7559);
nor U7940 (N_7940,N_7748,N_7502);
xor U7941 (N_7941,N_7540,N_7590);
nand U7942 (N_7942,N_7756,N_7672);
nor U7943 (N_7943,N_7625,N_7707);
or U7944 (N_7944,N_7532,N_7689);
or U7945 (N_7945,N_7604,N_7510);
and U7946 (N_7946,N_7681,N_7517);
nor U7947 (N_7947,N_7731,N_7643);
xnor U7948 (N_7948,N_7516,N_7602);
and U7949 (N_7949,N_7606,N_7522);
xor U7950 (N_7950,N_7699,N_7757);
nor U7951 (N_7951,N_7735,N_7720);
nand U7952 (N_7952,N_7709,N_7637);
xnor U7953 (N_7953,N_7711,N_7651);
nor U7954 (N_7954,N_7536,N_7753);
or U7955 (N_7955,N_7605,N_7590);
nand U7956 (N_7956,N_7724,N_7549);
or U7957 (N_7957,N_7611,N_7739);
xor U7958 (N_7958,N_7626,N_7631);
or U7959 (N_7959,N_7789,N_7769);
nand U7960 (N_7960,N_7547,N_7580);
xnor U7961 (N_7961,N_7646,N_7640);
or U7962 (N_7962,N_7730,N_7742);
nor U7963 (N_7963,N_7537,N_7548);
and U7964 (N_7964,N_7733,N_7771);
xnor U7965 (N_7965,N_7691,N_7546);
nand U7966 (N_7966,N_7716,N_7637);
or U7967 (N_7967,N_7639,N_7707);
nor U7968 (N_7968,N_7693,N_7788);
or U7969 (N_7969,N_7783,N_7658);
nand U7970 (N_7970,N_7670,N_7731);
or U7971 (N_7971,N_7786,N_7736);
nor U7972 (N_7972,N_7699,N_7513);
nor U7973 (N_7973,N_7582,N_7729);
and U7974 (N_7974,N_7758,N_7636);
xor U7975 (N_7975,N_7647,N_7760);
or U7976 (N_7976,N_7643,N_7514);
xnor U7977 (N_7977,N_7770,N_7564);
xor U7978 (N_7978,N_7763,N_7623);
nand U7979 (N_7979,N_7646,N_7663);
nand U7980 (N_7980,N_7636,N_7633);
xnor U7981 (N_7981,N_7635,N_7555);
nor U7982 (N_7982,N_7589,N_7641);
nor U7983 (N_7983,N_7524,N_7744);
nand U7984 (N_7984,N_7566,N_7711);
nor U7985 (N_7985,N_7695,N_7590);
or U7986 (N_7986,N_7771,N_7693);
or U7987 (N_7987,N_7651,N_7776);
xnor U7988 (N_7988,N_7544,N_7768);
and U7989 (N_7989,N_7699,N_7741);
xor U7990 (N_7990,N_7784,N_7520);
or U7991 (N_7991,N_7624,N_7784);
nor U7992 (N_7992,N_7607,N_7529);
or U7993 (N_7993,N_7578,N_7544);
xor U7994 (N_7994,N_7518,N_7676);
and U7995 (N_7995,N_7671,N_7762);
and U7996 (N_7996,N_7502,N_7567);
or U7997 (N_7997,N_7610,N_7718);
or U7998 (N_7998,N_7631,N_7642);
xnor U7999 (N_7999,N_7790,N_7537);
or U8000 (N_8000,N_7717,N_7773);
and U8001 (N_8001,N_7740,N_7570);
or U8002 (N_8002,N_7762,N_7635);
nand U8003 (N_8003,N_7675,N_7658);
nand U8004 (N_8004,N_7794,N_7704);
nor U8005 (N_8005,N_7519,N_7788);
nand U8006 (N_8006,N_7734,N_7525);
nor U8007 (N_8007,N_7638,N_7600);
or U8008 (N_8008,N_7678,N_7511);
and U8009 (N_8009,N_7783,N_7791);
and U8010 (N_8010,N_7506,N_7668);
nor U8011 (N_8011,N_7506,N_7541);
and U8012 (N_8012,N_7726,N_7591);
or U8013 (N_8013,N_7684,N_7610);
or U8014 (N_8014,N_7547,N_7608);
nor U8015 (N_8015,N_7676,N_7562);
nand U8016 (N_8016,N_7586,N_7654);
xnor U8017 (N_8017,N_7522,N_7695);
xnor U8018 (N_8018,N_7605,N_7781);
xor U8019 (N_8019,N_7744,N_7703);
or U8020 (N_8020,N_7668,N_7707);
xnor U8021 (N_8021,N_7667,N_7640);
nor U8022 (N_8022,N_7528,N_7709);
nor U8023 (N_8023,N_7734,N_7618);
xor U8024 (N_8024,N_7686,N_7603);
and U8025 (N_8025,N_7631,N_7619);
and U8026 (N_8026,N_7622,N_7564);
or U8027 (N_8027,N_7558,N_7615);
or U8028 (N_8028,N_7742,N_7578);
nand U8029 (N_8029,N_7582,N_7553);
and U8030 (N_8030,N_7607,N_7617);
or U8031 (N_8031,N_7516,N_7569);
or U8032 (N_8032,N_7532,N_7676);
nand U8033 (N_8033,N_7511,N_7568);
xnor U8034 (N_8034,N_7706,N_7578);
or U8035 (N_8035,N_7643,N_7610);
or U8036 (N_8036,N_7714,N_7752);
and U8037 (N_8037,N_7518,N_7607);
or U8038 (N_8038,N_7622,N_7550);
or U8039 (N_8039,N_7730,N_7529);
nand U8040 (N_8040,N_7762,N_7739);
nor U8041 (N_8041,N_7692,N_7662);
nand U8042 (N_8042,N_7548,N_7794);
nor U8043 (N_8043,N_7573,N_7532);
xor U8044 (N_8044,N_7725,N_7749);
xor U8045 (N_8045,N_7635,N_7773);
nor U8046 (N_8046,N_7733,N_7670);
xnor U8047 (N_8047,N_7538,N_7791);
nand U8048 (N_8048,N_7698,N_7549);
nand U8049 (N_8049,N_7766,N_7513);
and U8050 (N_8050,N_7534,N_7537);
xor U8051 (N_8051,N_7655,N_7543);
or U8052 (N_8052,N_7764,N_7699);
or U8053 (N_8053,N_7666,N_7664);
nor U8054 (N_8054,N_7633,N_7676);
xor U8055 (N_8055,N_7725,N_7597);
or U8056 (N_8056,N_7659,N_7587);
nand U8057 (N_8057,N_7751,N_7621);
nand U8058 (N_8058,N_7684,N_7611);
or U8059 (N_8059,N_7785,N_7569);
or U8060 (N_8060,N_7693,N_7576);
and U8061 (N_8061,N_7745,N_7771);
nor U8062 (N_8062,N_7516,N_7703);
or U8063 (N_8063,N_7783,N_7597);
and U8064 (N_8064,N_7543,N_7785);
nor U8065 (N_8065,N_7549,N_7796);
nand U8066 (N_8066,N_7603,N_7706);
nor U8067 (N_8067,N_7786,N_7696);
xor U8068 (N_8068,N_7550,N_7751);
xor U8069 (N_8069,N_7754,N_7549);
xor U8070 (N_8070,N_7582,N_7621);
and U8071 (N_8071,N_7506,N_7731);
xor U8072 (N_8072,N_7540,N_7746);
nor U8073 (N_8073,N_7682,N_7642);
nand U8074 (N_8074,N_7755,N_7543);
or U8075 (N_8075,N_7547,N_7724);
xnor U8076 (N_8076,N_7627,N_7514);
or U8077 (N_8077,N_7678,N_7629);
nand U8078 (N_8078,N_7760,N_7616);
and U8079 (N_8079,N_7550,N_7624);
xor U8080 (N_8080,N_7574,N_7692);
and U8081 (N_8081,N_7732,N_7608);
and U8082 (N_8082,N_7584,N_7677);
and U8083 (N_8083,N_7656,N_7788);
or U8084 (N_8084,N_7560,N_7677);
xor U8085 (N_8085,N_7627,N_7555);
nand U8086 (N_8086,N_7666,N_7608);
nor U8087 (N_8087,N_7674,N_7592);
nor U8088 (N_8088,N_7785,N_7767);
xor U8089 (N_8089,N_7504,N_7626);
xor U8090 (N_8090,N_7555,N_7656);
nand U8091 (N_8091,N_7561,N_7628);
and U8092 (N_8092,N_7531,N_7619);
and U8093 (N_8093,N_7670,N_7621);
or U8094 (N_8094,N_7512,N_7736);
xor U8095 (N_8095,N_7728,N_7515);
nand U8096 (N_8096,N_7724,N_7590);
nor U8097 (N_8097,N_7633,N_7774);
nand U8098 (N_8098,N_7737,N_7542);
xor U8099 (N_8099,N_7599,N_7731);
nor U8100 (N_8100,N_7872,N_7957);
nand U8101 (N_8101,N_7908,N_7956);
or U8102 (N_8102,N_7968,N_7869);
xor U8103 (N_8103,N_7945,N_7987);
and U8104 (N_8104,N_8095,N_8001);
or U8105 (N_8105,N_8087,N_7954);
or U8106 (N_8106,N_8050,N_8024);
nand U8107 (N_8107,N_7824,N_7856);
nor U8108 (N_8108,N_7922,N_7996);
nand U8109 (N_8109,N_7835,N_7823);
nand U8110 (N_8110,N_8068,N_7928);
nand U8111 (N_8111,N_7983,N_7925);
xor U8112 (N_8112,N_8042,N_8000);
nor U8113 (N_8113,N_7969,N_7955);
nor U8114 (N_8114,N_7938,N_7897);
nor U8115 (N_8115,N_7967,N_8061);
nor U8116 (N_8116,N_7865,N_8079);
and U8117 (N_8117,N_7936,N_8058);
xor U8118 (N_8118,N_8051,N_8028);
xor U8119 (N_8119,N_7933,N_8093);
or U8120 (N_8120,N_8082,N_7907);
nand U8121 (N_8121,N_7826,N_7975);
nand U8122 (N_8122,N_7802,N_7923);
nand U8123 (N_8123,N_7934,N_7986);
and U8124 (N_8124,N_7931,N_7951);
and U8125 (N_8125,N_7855,N_7803);
or U8126 (N_8126,N_7812,N_7810);
or U8127 (N_8127,N_7952,N_7866);
nand U8128 (N_8128,N_7960,N_7962);
nor U8129 (N_8129,N_7927,N_7919);
or U8130 (N_8130,N_7997,N_7913);
xnor U8131 (N_8131,N_8086,N_7868);
and U8132 (N_8132,N_7876,N_8053);
nor U8133 (N_8133,N_8033,N_7830);
and U8134 (N_8134,N_7822,N_7905);
nand U8135 (N_8135,N_7992,N_7970);
and U8136 (N_8136,N_7892,N_7867);
nor U8137 (N_8137,N_8013,N_7980);
nor U8138 (N_8138,N_8098,N_7929);
and U8139 (N_8139,N_7881,N_7893);
nand U8140 (N_8140,N_8083,N_7946);
or U8141 (N_8141,N_7948,N_7806);
nor U8142 (N_8142,N_8046,N_7832);
or U8143 (N_8143,N_7808,N_8032);
or U8144 (N_8144,N_8091,N_8005);
and U8145 (N_8145,N_8072,N_8022);
and U8146 (N_8146,N_8077,N_7889);
and U8147 (N_8147,N_7801,N_7860);
and U8148 (N_8148,N_7845,N_7819);
nor U8149 (N_8149,N_7836,N_7877);
and U8150 (N_8150,N_7906,N_8043);
nand U8151 (N_8151,N_7871,N_7984);
xor U8152 (N_8152,N_8034,N_7800);
or U8153 (N_8153,N_7921,N_7879);
nand U8154 (N_8154,N_7890,N_7976);
nand U8155 (N_8155,N_8047,N_7891);
nand U8156 (N_8156,N_7900,N_8003);
or U8157 (N_8157,N_7973,N_8085);
and U8158 (N_8158,N_7941,N_7809);
xnor U8159 (N_8159,N_7961,N_7989);
or U8160 (N_8160,N_8063,N_7886);
xor U8161 (N_8161,N_8020,N_7972);
or U8162 (N_8162,N_8048,N_8088);
nand U8163 (N_8163,N_8015,N_8065);
or U8164 (N_8164,N_7994,N_7862);
xnor U8165 (N_8165,N_7846,N_7943);
or U8166 (N_8166,N_8014,N_7998);
nor U8167 (N_8167,N_7979,N_8070);
and U8168 (N_8168,N_8074,N_7971);
and U8169 (N_8169,N_8002,N_8059);
xor U8170 (N_8170,N_7834,N_7880);
and U8171 (N_8171,N_7844,N_7829);
nand U8172 (N_8172,N_8052,N_8094);
and U8173 (N_8173,N_7870,N_7939);
nand U8174 (N_8174,N_7804,N_7974);
xor U8175 (N_8175,N_7878,N_8078);
nand U8176 (N_8176,N_8011,N_7841);
and U8177 (N_8177,N_8096,N_7859);
or U8178 (N_8178,N_8060,N_8017);
and U8179 (N_8179,N_7937,N_7902);
and U8180 (N_8180,N_7833,N_7942);
nand U8181 (N_8181,N_7932,N_7904);
xnor U8182 (N_8182,N_7837,N_8069);
nor U8183 (N_8183,N_8090,N_7926);
or U8184 (N_8184,N_8009,N_8075);
nand U8185 (N_8185,N_7842,N_7895);
or U8186 (N_8186,N_7818,N_7982);
nor U8187 (N_8187,N_7914,N_8027);
and U8188 (N_8188,N_7817,N_8073);
nand U8189 (N_8189,N_7944,N_7838);
nor U8190 (N_8190,N_7857,N_7827);
xnor U8191 (N_8191,N_8039,N_7848);
xnor U8192 (N_8192,N_8025,N_7816);
or U8193 (N_8193,N_7920,N_7851);
nor U8194 (N_8194,N_7940,N_7917);
nand U8195 (N_8195,N_7847,N_7874);
xor U8196 (N_8196,N_7911,N_8023);
and U8197 (N_8197,N_7959,N_8036);
xor U8198 (N_8198,N_8057,N_7915);
nand U8199 (N_8199,N_7977,N_7805);
nor U8200 (N_8200,N_8016,N_7853);
xnor U8201 (N_8201,N_8071,N_8097);
nor U8202 (N_8202,N_8038,N_7811);
xnor U8203 (N_8203,N_8054,N_7815);
and U8204 (N_8204,N_7843,N_7888);
xnor U8205 (N_8205,N_7873,N_7883);
nand U8206 (N_8206,N_8008,N_7950);
and U8207 (N_8207,N_7985,N_8018);
nand U8208 (N_8208,N_7947,N_7899);
nand U8209 (N_8209,N_8076,N_7953);
nand U8210 (N_8210,N_7918,N_8030);
xor U8211 (N_8211,N_7882,N_7978);
nand U8212 (N_8212,N_8006,N_7850);
nor U8213 (N_8213,N_8007,N_7864);
or U8214 (N_8214,N_7820,N_7993);
xnor U8215 (N_8215,N_8026,N_7903);
nor U8216 (N_8216,N_8044,N_7958);
nand U8217 (N_8217,N_8056,N_8031);
and U8218 (N_8218,N_7924,N_7909);
nand U8219 (N_8219,N_7840,N_7964);
nand U8220 (N_8220,N_7949,N_8062);
or U8221 (N_8221,N_8092,N_8067);
or U8222 (N_8222,N_7963,N_7828);
or U8223 (N_8223,N_7898,N_7916);
xnor U8224 (N_8224,N_8019,N_7930);
xor U8225 (N_8225,N_7910,N_8012);
or U8226 (N_8226,N_7912,N_8037);
nand U8227 (N_8227,N_7813,N_7814);
or U8228 (N_8228,N_7901,N_8064);
and U8229 (N_8229,N_8004,N_7807);
nor U8230 (N_8230,N_8066,N_8029);
nand U8231 (N_8231,N_8041,N_7884);
xnor U8232 (N_8232,N_7863,N_7935);
nand U8233 (N_8233,N_7852,N_7849);
or U8234 (N_8234,N_7990,N_7999);
nand U8235 (N_8235,N_7858,N_7991);
nand U8236 (N_8236,N_8089,N_7821);
xor U8237 (N_8237,N_7896,N_8045);
xnor U8238 (N_8238,N_7966,N_7885);
or U8239 (N_8239,N_7887,N_8080);
or U8240 (N_8240,N_8099,N_7981);
nor U8241 (N_8241,N_7825,N_7965);
and U8242 (N_8242,N_7831,N_8049);
xnor U8243 (N_8243,N_8035,N_8084);
or U8244 (N_8244,N_7854,N_7839);
nand U8245 (N_8245,N_8010,N_7861);
nand U8246 (N_8246,N_8021,N_7894);
or U8247 (N_8247,N_7875,N_8040);
and U8248 (N_8248,N_8055,N_7988);
xnor U8249 (N_8249,N_8081,N_7995);
or U8250 (N_8250,N_7915,N_7940);
nand U8251 (N_8251,N_7846,N_7896);
nor U8252 (N_8252,N_7843,N_7877);
and U8253 (N_8253,N_7917,N_7832);
or U8254 (N_8254,N_7821,N_7971);
or U8255 (N_8255,N_7954,N_8013);
xor U8256 (N_8256,N_8037,N_7949);
xor U8257 (N_8257,N_7882,N_7879);
and U8258 (N_8258,N_8064,N_7806);
nand U8259 (N_8259,N_8021,N_8062);
nand U8260 (N_8260,N_8091,N_8012);
xnor U8261 (N_8261,N_7899,N_7908);
nor U8262 (N_8262,N_7948,N_7816);
nor U8263 (N_8263,N_7821,N_7913);
or U8264 (N_8264,N_8048,N_7958);
xnor U8265 (N_8265,N_7974,N_7809);
and U8266 (N_8266,N_7859,N_8030);
nor U8267 (N_8267,N_7913,N_8088);
or U8268 (N_8268,N_7805,N_7819);
nor U8269 (N_8269,N_7917,N_7977);
and U8270 (N_8270,N_7875,N_7920);
or U8271 (N_8271,N_8037,N_7938);
xnor U8272 (N_8272,N_7975,N_7810);
nand U8273 (N_8273,N_7969,N_7981);
nor U8274 (N_8274,N_7964,N_7958);
or U8275 (N_8275,N_7806,N_7933);
nor U8276 (N_8276,N_7966,N_7893);
or U8277 (N_8277,N_7901,N_8003);
nand U8278 (N_8278,N_7829,N_7822);
and U8279 (N_8279,N_8011,N_7944);
and U8280 (N_8280,N_8005,N_8072);
nor U8281 (N_8281,N_7801,N_7904);
and U8282 (N_8282,N_7950,N_7834);
xor U8283 (N_8283,N_8008,N_8021);
or U8284 (N_8284,N_8003,N_7961);
nor U8285 (N_8285,N_7921,N_8060);
nor U8286 (N_8286,N_7893,N_8041);
or U8287 (N_8287,N_7927,N_7928);
and U8288 (N_8288,N_7946,N_7827);
xor U8289 (N_8289,N_7904,N_7825);
nand U8290 (N_8290,N_7947,N_7985);
nand U8291 (N_8291,N_8075,N_7999);
nand U8292 (N_8292,N_7900,N_8068);
xnor U8293 (N_8293,N_7818,N_8099);
nand U8294 (N_8294,N_7802,N_7934);
or U8295 (N_8295,N_7894,N_7917);
nand U8296 (N_8296,N_7832,N_7810);
nand U8297 (N_8297,N_8048,N_7984);
xor U8298 (N_8298,N_7851,N_7921);
nand U8299 (N_8299,N_7883,N_8014);
or U8300 (N_8300,N_7961,N_8045);
nand U8301 (N_8301,N_7876,N_7972);
nor U8302 (N_8302,N_7821,N_7980);
and U8303 (N_8303,N_8096,N_8053);
nor U8304 (N_8304,N_7902,N_7826);
or U8305 (N_8305,N_8058,N_7876);
nand U8306 (N_8306,N_7835,N_7892);
or U8307 (N_8307,N_8072,N_8034);
nand U8308 (N_8308,N_7898,N_7927);
nor U8309 (N_8309,N_7900,N_7814);
nand U8310 (N_8310,N_7986,N_7807);
nand U8311 (N_8311,N_7969,N_8014);
nand U8312 (N_8312,N_8060,N_7886);
nor U8313 (N_8313,N_8035,N_8099);
or U8314 (N_8314,N_7905,N_7849);
nand U8315 (N_8315,N_8084,N_7857);
xor U8316 (N_8316,N_7866,N_7955);
xnor U8317 (N_8317,N_7807,N_8096);
and U8318 (N_8318,N_7883,N_8036);
nand U8319 (N_8319,N_7832,N_8023);
and U8320 (N_8320,N_7936,N_8060);
xnor U8321 (N_8321,N_7974,N_7950);
and U8322 (N_8322,N_8092,N_7892);
nor U8323 (N_8323,N_7948,N_7857);
nand U8324 (N_8324,N_8046,N_7957);
nand U8325 (N_8325,N_7989,N_7969);
or U8326 (N_8326,N_7871,N_7829);
nand U8327 (N_8327,N_7901,N_7913);
nand U8328 (N_8328,N_7929,N_7913);
nand U8329 (N_8329,N_7818,N_7966);
xor U8330 (N_8330,N_8036,N_7988);
nand U8331 (N_8331,N_7953,N_7836);
xnor U8332 (N_8332,N_7817,N_7906);
nor U8333 (N_8333,N_7988,N_7894);
nor U8334 (N_8334,N_7833,N_8085);
or U8335 (N_8335,N_8034,N_7905);
nand U8336 (N_8336,N_7943,N_7981);
nand U8337 (N_8337,N_7801,N_7999);
and U8338 (N_8338,N_7891,N_7997);
or U8339 (N_8339,N_8023,N_7918);
xnor U8340 (N_8340,N_7877,N_7927);
nor U8341 (N_8341,N_7970,N_8062);
nand U8342 (N_8342,N_7964,N_7845);
and U8343 (N_8343,N_8019,N_7831);
xor U8344 (N_8344,N_7975,N_7850);
nor U8345 (N_8345,N_8096,N_7879);
or U8346 (N_8346,N_8025,N_7818);
nand U8347 (N_8347,N_8083,N_7881);
nor U8348 (N_8348,N_7889,N_7974);
or U8349 (N_8349,N_7812,N_7830);
nand U8350 (N_8350,N_7936,N_7823);
nand U8351 (N_8351,N_7840,N_7977);
and U8352 (N_8352,N_7825,N_8022);
nor U8353 (N_8353,N_7884,N_7832);
and U8354 (N_8354,N_7943,N_7918);
nand U8355 (N_8355,N_8014,N_8091);
or U8356 (N_8356,N_8073,N_7884);
and U8357 (N_8357,N_7862,N_7873);
or U8358 (N_8358,N_7973,N_8005);
or U8359 (N_8359,N_8083,N_8017);
and U8360 (N_8360,N_7967,N_7963);
and U8361 (N_8361,N_8036,N_8050);
and U8362 (N_8362,N_7821,N_8030);
and U8363 (N_8363,N_8030,N_7853);
nand U8364 (N_8364,N_8022,N_7919);
or U8365 (N_8365,N_7923,N_7934);
and U8366 (N_8366,N_8000,N_8059);
nor U8367 (N_8367,N_7804,N_8006);
xnor U8368 (N_8368,N_8068,N_7873);
nor U8369 (N_8369,N_7999,N_7910);
and U8370 (N_8370,N_7951,N_7954);
nor U8371 (N_8371,N_7986,N_7846);
xnor U8372 (N_8372,N_7898,N_8003);
nand U8373 (N_8373,N_7970,N_7997);
nand U8374 (N_8374,N_8007,N_8084);
nand U8375 (N_8375,N_8027,N_7945);
and U8376 (N_8376,N_8006,N_8062);
and U8377 (N_8377,N_7824,N_7835);
nand U8378 (N_8378,N_7970,N_7883);
xnor U8379 (N_8379,N_7906,N_7865);
or U8380 (N_8380,N_7964,N_8009);
xor U8381 (N_8381,N_7987,N_8089);
or U8382 (N_8382,N_7804,N_7966);
or U8383 (N_8383,N_8027,N_7968);
or U8384 (N_8384,N_8099,N_7980);
and U8385 (N_8385,N_8067,N_8095);
xor U8386 (N_8386,N_7920,N_7824);
and U8387 (N_8387,N_7967,N_8045);
and U8388 (N_8388,N_7888,N_7977);
xnor U8389 (N_8389,N_7851,N_8009);
nand U8390 (N_8390,N_7953,N_7925);
nor U8391 (N_8391,N_8070,N_8097);
and U8392 (N_8392,N_7934,N_7956);
nor U8393 (N_8393,N_7894,N_7805);
nand U8394 (N_8394,N_7895,N_8028);
nand U8395 (N_8395,N_7988,N_8000);
nand U8396 (N_8396,N_7962,N_8084);
and U8397 (N_8397,N_8020,N_7874);
and U8398 (N_8398,N_7837,N_8084);
nand U8399 (N_8399,N_7828,N_8036);
or U8400 (N_8400,N_8372,N_8229);
or U8401 (N_8401,N_8174,N_8121);
nand U8402 (N_8402,N_8267,N_8338);
nand U8403 (N_8403,N_8398,N_8220);
or U8404 (N_8404,N_8193,N_8232);
or U8405 (N_8405,N_8138,N_8110);
and U8406 (N_8406,N_8360,N_8391);
nand U8407 (N_8407,N_8176,N_8265);
nand U8408 (N_8408,N_8393,N_8242);
and U8409 (N_8409,N_8339,N_8368);
nor U8410 (N_8410,N_8126,N_8266);
xnor U8411 (N_8411,N_8227,N_8216);
nor U8412 (N_8412,N_8109,N_8334);
and U8413 (N_8413,N_8268,N_8178);
or U8414 (N_8414,N_8112,N_8206);
xnor U8415 (N_8415,N_8326,N_8210);
and U8416 (N_8416,N_8134,N_8374);
or U8417 (N_8417,N_8256,N_8188);
xor U8418 (N_8418,N_8284,N_8328);
and U8419 (N_8419,N_8342,N_8155);
nand U8420 (N_8420,N_8355,N_8335);
or U8421 (N_8421,N_8396,N_8141);
xor U8422 (N_8422,N_8129,N_8181);
nand U8423 (N_8423,N_8128,N_8204);
or U8424 (N_8424,N_8389,N_8226);
xor U8425 (N_8425,N_8249,N_8202);
and U8426 (N_8426,N_8333,N_8386);
or U8427 (N_8427,N_8297,N_8315);
nand U8428 (N_8428,N_8157,N_8296);
xnor U8429 (N_8429,N_8382,N_8292);
xor U8430 (N_8430,N_8131,N_8158);
nor U8431 (N_8431,N_8303,N_8218);
xor U8432 (N_8432,N_8246,N_8160);
nor U8433 (N_8433,N_8214,N_8252);
xor U8434 (N_8434,N_8180,N_8179);
or U8435 (N_8435,N_8195,N_8230);
or U8436 (N_8436,N_8197,N_8279);
nor U8437 (N_8437,N_8211,N_8212);
nand U8438 (N_8438,N_8100,N_8271);
nor U8439 (N_8439,N_8111,N_8270);
and U8440 (N_8440,N_8171,N_8104);
or U8441 (N_8441,N_8184,N_8235);
nand U8442 (N_8442,N_8283,N_8194);
or U8443 (N_8443,N_8170,N_8311);
xnor U8444 (N_8444,N_8125,N_8263);
nand U8445 (N_8445,N_8352,N_8224);
nor U8446 (N_8446,N_8161,N_8213);
xnor U8447 (N_8447,N_8369,N_8375);
nand U8448 (N_8448,N_8124,N_8319);
nand U8449 (N_8449,N_8321,N_8277);
nor U8450 (N_8450,N_8346,N_8127);
and U8451 (N_8451,N_8231,N_8240);
and U8452 (N_8452,N_8164,N_8349);
xor U8453 (N_8453,N_8278,N_8365);
and U8454 (N_8454,N_8172,N_8169);
and U8455 (N_8455,N_8247,N_8376);
nor U8456 (N_8456,N_8120,N_8244);
or U8457 (N_8457,N_8237,N_8183);
xor U8458 (N_8458,N_8384,N_8275);
xnor U8459 (N_8459,N_8136,N_8307);
xor U8460 (N_8460,N_8113,N_8239);
nor U8461 (N_8461,N_8133,N_8222);
xnor U8462 (N_8462,N_8156,N_8289);
and U8463 (N_8463,N_8258,N_8312);
or U8464 (N_8464,N_8103,N_8234);
and U8465 (N_8465,N_8253,N_8395);
xnor U8466 (N_8466,N_8152,N_8225);
nor U8467 (N_8467,N_8381,N_8264);
or U8468 (N_8468,N_8219,N_8101);
and U8469 (N_8469,N_8228,N_8288);
and U8470 (N_8470,N_8354,N_8119);
and U8471 (N_8471,N_8371,N_8168);
nor U8472 (N_8472,N_8347,N_8191);
nand U8473 (N_8473,N_8313,N_8196);
xor U8474 (N_8474,N_8116,N_8105);
nand U8475 (N_8475,N_8345,N_8397);
and U8476 (N_8476,N_8135,N_8337);
nor U8477 (N_8477,N_8325,N_8379);
and U8478 (N_8478,N_8273,N_8286);
nand U8479 (N_8479,N_8150,N_8274);
xor U8480 (N_8480,N_8107,N_8329);
nand U8481 (N_8481,N_8336,N_8380);
nand U8482 (N_8482,N_8254,N_8309);
xor U8483 (N_8483,N_8317,N_8294);
nand U8484 (N_8484,N_8366,N_8177);
nand U8485 (N_8485,N_8159,N_8318);
nand U8486 (N_8486,N_8358,N_8241);
and U8487 (N_8487,N_8377,N_8282);
xor U8488 (N_8488,N_8373,N_8167);
nor U8489 (N_8489,N_8359,N_8139);
or U8490 (N_8490,N_8122,N_8298);
xor U8491 (N_8491,N_8162,N_8387);
nor U8492 (N_8492,N_8272,N_8343);
or U8493 (N_8493,N_8291,N_8245);
xnor U8494 (N_8494,N_8378,N_8327);
or U8495 (N_8495,N_8189,N_8163);
nand U8496 (N_8496,N_8285,N_8305);
nand U8497 (N_8497,N_8123,N_8302);
xor U8498 (N_8498,N_8262,N_8146);
or U8499 (N_8499,N_8293,N_8306);
and U8500 (N_8500,N_8165,N_8259);
and U8501 (N_8501,N_8173,N_8115);
xor U8502 (N_8502,N_8310,N_8323);
nand U8503 (N_8503,N_8370,N_8186);
or U8504 (N_8504,N_8332,N_8207);
and U8505 (N_8505,N_8132,N_8215);
and U8506 (N_8506,N_8390,N_8320);
nor U8507 (N_8507,N_8185,N_8209);
and U8508 (N_8508,N_8314,N_8153);
and U8509 (N_8509,N_8200,N_8394);
xor U8510 (N_8510,N_8149,N_8399);
or U8511 (N_8511,N_8348,N_8144);
xnor U8512 (N_8512,N_8203,N_8248);
and U8513 (N_8513,N_8148,N_8290);
xnor U8514 (N_8514,N_8357,N_8299);
or U8515 (N_8515,N_8205,N_8117);
nor U8516 (N_8516,N_8356,N_8316);
xor U8517 (N_8517,N_8145,N_8322);
and U8518 (N_8518,N_8243,N_8341);
nor U8519 (N_8519,N_8208,N_8182);
nand U8520 (N_8520,N_8269,N_8287);
xnor U8521 (N_8521,N_8154,N_8143);
xnor U8522 (N_8522,N_8166,N_8392);
xor U8523 (N_8523,N_8192,N_8137);
nor U8524 (N_8524,N_8175,N_8276);
xnor U8525 (N_8525,N_8304,N_8367);
nand U8526 (N_8526,N_8114,N_8142);
xor U8527 (N_8527,N_8187,N_8217);
nand U8528 (N_8528,N_8364,N_8118);
or U8529 (N_8529,N_8190,N_8223);
and U8530 (N_8530,N_8324,N_8221);
or U8531 (N_8531,N_8300,N_8238);
and U8532 (N_8532,N_8151,N_8363);
and U8533 (N_8533,N_8130,N_8261);
nor U8534 (N_8534,N_8388,N_8280);
xnor U8535 (N_8535,N_8353,N_8383);
nand U8536 (N_8536,N_8255,N_8260);
or U8537 (N_8537,N_8330,N_8362);
xor U8538 (N_8538,N_8295,N_8331);
and U8539 (N_8539,N_8340,N_8102);
or U8540 (N_8540,N_8281,N_8385);
nand U8541 (N_8541,N_8140,N_8361);
nand U8542 (N_8542,N_8147,N_8108);
nand U8543 (N_8543,N_8251,N_8301);
nand U8544 (N_8544,N_8106,N_8250);
or U8545 (N_8545,N_8236,N_8233);
and U8546 (N_8546,N_8308,N_8199);
nor U8547 (N_8547,N_8350,N_8351);
nor U8548 (N_8548,N_8257,N_8198);
nor U8549 (N_8549,N_8344,N_8201);
nand U8550 (N_8550,N_8387,N_8117);
or U8551 (N_8551,N_8170,N_8167);
or U8552 (N_8552,N_8186,N_8188);
and U8553 (N_8553,N_8183,N_8352);
xnor U8554 (N_8554,N_8361,N_8271);
nor U8555 (N_8555,N_8128,N_8379);
nand U8556 (N_8556,N_8132,N_8363);
or U8557 (N_8557,N_8122,N_8355);
nor U8558 (N_8558,N_8251,N_8164);
or U8559 (N_8559,N_8285,N_8217);
and U8560 (N_8560,N_8218,N_8118);
and U8561 (N_8561,N_8162,N_8388);
nor U8562 (N_8562,N_8301,N_8393);
nor U8563 (N_8563,N_8141,N_8308);
or U8564 (N_8564,N_8228,N_8305);
nor U8565 (N_8565,N_8113,N_8230);
nand U8566 (N_8566,N_8231,N_8193);
xnor U8567 (N_8567,N_8215,N_8319);
xnor U8568 (N_8568,N_8307,N_8221);
nor U8569 (N_8569,N_8155,N_8379);
and U8570 (N_8570,N_8111,N_8295);
and U8571 (N_8571,N_8349,N_8353);
or U8572 (N_8572,N_8210,N_8284);
nor U8573 (N_8573,N_8249,N_8376);
or U8574 (N_8574,N_8104,N_8339);
and U8575 (N_8575,N_8168,N_8126);
and U8576 (N_8576,N_8174,N_8382);
and U8577 (N_8577,N_8345,N_8169);
and U8578 (N_8578,N_8243,N_8322);
nand U8579 (N_8579,N_8209,N_8103);
nand U8580 (N_8580,N_8181,N_8126);
xor U8581 (N_8581,N_8370,N_8181);
nor U8582 (N_8582,N_8370,N_8379);
nand U8583 (N_8583,N_8174,N_8113);
and U8584 (N_8584,N_8243,N_8202);
or U8585 (N_8585,N_8271,N_8328);
nand U8586 (N_8586,N_8158,N_8208);
nor U8587 (N_8587,N_8129,N_8255);
and U8588 (N_8588,N_8340,N_8115);
nand U8589 (N_8589,N_8201,N_8320);
or U8590 (N_8590,N_8339,N_8214);
xnor U8591 (N_8591,N_8226,N_8138);
nor U8592 (N_8592,N_8305,N_8226);
nand U8593 (N_8593,N_8329,N_8376);
or U8594 (N_8594,N_8211,N_8106);
nand U8595 (N_8595,N_8327,N_8113);
or U8596 (N_8596,N_8224,N_8216);
nand U8597 (N_8597,N_8214,N_8165);
or U8598 (N_8598,N_8155,N_8246);
xor U8599 (N_8599,N_8295,N_8250);
xnor U8600 (N_8600,N_8121,N_8386);
nand U8601 (N_8601,N_8246,N_8217);
nand U8602 (N_8602,N_8347,N_8217);
xnor U8603 (N_8603,N_8213,N_8137);
nand U8604 (N_8604,N_8120,N_8254);
and U8605 (N_8605,N_8382,N_8154);
xnor U8606 (N_8606,N_8103,N_8228);
or U8607 (N_8607,N_8125,N_8231);
nand U8608 (N_8608,N_8195,N_8243);
xor U8609 (N_8609,N_8148,N_8384);
nor U8610 (N_8610,N_8282,N_8294);
and U8611 (N_8611,N_8368,N_8270);
or U8612 (N_8612,N_8365,N_8169);
xor U8613 (N_8613,N_8131,N_8107);
nor U8614 (N_8614,N_8360,N_8242);
nor U8615 (N_8615,N_8307,N_8210);
or U8616 (N_8616,N_8359,N_8244);
xnor U8617 (N_8617,N_8247,N_8312);
and U8618 (N_8618,N_8222,N_8121);
or U8619 (N_8619,N_8145,N_8397);
xor U8620 (N_8620,N_8166,N_8267);
nor U8621 (N_8621,N_8346,N_8241);
or U8622 (N_8622,N_8390,N_8349);
xor U8623 (N_8623,N_8186,N_8140);
and U8624 (N_8624,N_8263,N_8382);
xnor U8625 (N_8625,N_8301,N_8148);
nor U8626 (N_8626,N_8186,N_8143);
nor U8627 (N_8627,N_8172,N_8112);
and U8628 (N_8628,N_8114,N_8289);
or U8629 (N_8629,N_8218,N_8338);
nand U8630 (N_8630,N_8383,N_8242);
nand U8631 (N_8631,N_8118,N_8232);
and U8632 (N_8632,N_8102,N_8232);
xnor U8633 (N_8633,N_8341,N_8149);
xor U8634 (N_8634,N_8246,N_8151);
or U8635 (N_8635,N_8230,N_8348);
or U8636 (N_8636,N_8382,N_8225);
and U8637 (N_8637,N_8178,N_8351);
and U8638 (N_8638,N_8189,N_8340);
and U8639 (N_8639,N_8150,N_8382);
and U8640 (N_8640,N_8142,N_8229);
and U8641 (N_8641,N_8206,N_8236);
nand U8642 (N_8642,N_8393,N_8215);
xor U8643 (N_8643,N_8249,N_8207);
xnor U8644 (N_8644,N_8319,N_8200);
nor U8645 (N_8645,N_8209,N_8214);
or U8646 (N_8646,N_8155,N_8237);
nand U8647 (N_8647,N_8301,N_8367);
nand U8648 (N_8648,N_8132,N_8118);
or U8649 (N_8649,N_8112,N_8240);
nor U8650 (N_8650,N_8105,N_8244);
xnor U8651 (N_8651,N_8189,N_8169);
xnor U8652 (N_8652,N_8291,N_8382);
or U8653 (N_8653,N_8336,N_8105);
nor U8654 (N_8654,N_8309,N_8186);
nand U8655 (N_8655,N_8154,N_8376);
nor U8656 (N_8656,N_8139,N_8196);
nand U8657 (N_8657,N_8106,N_8272);
xnor U8658 (N_8658,N_8146,N_8143);
xnor U8659 (N_8659,N_8232,N_8274);
xor U8660 (N_8660,N_8289,N_8325);
nand U8661 (N_8661,N_8101,N_8221);
and U8662 (N_8662,N_8199,N_8399);
and U8663 (N_8663,N_8399,N_8342);
or U8664 (N_8664,N_8104,N_8251);
xnor U8665 (N_8665,N_8187,N_8383);
xor U8666 (N_8666,N_8134,N_8218);
xor U8667 (N_8667,N_8160,N_8266);
or U8668 (N_8668,N_8265,N_8356);
xor U8669 (N_8669,N_8343,N_8256);
nor U8670 (N_8670,N_8178,N_8153);
or U8671 (N_8671,N_8144,N_8303);
nor U8672 (N_8672,N_8312,N_8131);
nor U8673 (N_8673,N_8180,N_8165);
xnor U8674 (N_8674,N_8261,N_8195);
xnor U8675 (N_8675,N_8267,N_8236);
nor U8676 (N_8676,N_8245,N_8363);
and U8677 (N_8677,N_8329,N_8212);
nor U8678 (N_8678,N_8160,N_8197);
xor U8679 (N_8679,N_8256,N_8332);
and U8680 (N_8680,N_8355,N_8210);
nor U8681 (N_8681,N_8303,N_8161);
and U8682 (N_8682,N_8153,N_8327);
nor U8683 (N_8683,N_8184,N_8206);
xor U8684 (N_8684,N_8329,N_8233);
xor U8685 (N_8685,N_8338,N_8253);
xor U8686 (N_8686,N_8371,N_8175);
xnor U8687 (N_8687,N_8388,N_8317);
or U8688 (N_8688,N_8167,N_8361);
or U8689 (N_8689,N_8213,N_8333);
nand U8690 (N_8690,N_8174,N_8235);
nor U8691 (N_8691,N_8353,N_8389);
nand U8692 (N_8692,N_8315,N_8139);
or U8693 (N_8693,N_8203,N_8307);
and U8694 (N_8694,N_8396,N_8369);
and U8695 (N_8695,N_8207,N_8323);
nand U8696 (N_8696,N_8281,N_8299);
and U8697 (N_8697,N_8135,N_8254);
nor U8698 (N_8698,N_8246,N_8148);
nor U8699 (N_8699,N_8104,N_8141);
or U8700 (N_8700,N_8416,N_8583);
nor U8701 (N_8701,N_8697,N_8579);
xor U8702 (N_8702,N_8445,N_8414);
xor U8703 (N_8703,N_8454,N_8550);
nand U8704 (N_8704,N_8568,N_8566);
or U8705 (N_8705,N_8594,N_8654);
and U8706 (N_8706,N_8402,N_8430);
xnor U8707 (N_8707,N_8538,N_8493);
or U8708 (N_8708,N_8422,N_8496);
nor U8709 (N_8709,N_8500,N_8601);
xnor U8710 (N_8710,N_8606,N_8668);
and U8711 (N_8711,N_8597,N_8415);
and U8712 (N_8712,N_8464,N_8541);
xor U8713 (N_8713,N_8684,N_8623);
nor U8714 (N_8714,N_8656,N_8551);
and U8715 (N_8715,N_8643,N_8636);
and U8716 (N_8716,N_8535,N_8463);
or U8717 (N_8717,N_8460,N_8452);
nor U8718 (N_8718,N_8404,N_8588);
nand U8719 (N_8719,N_8652,N_8562);
and U8720 (N_8720,N_8521,N_8455);
or U8721 (N_8721,N_8598,N_8631);
nand U8722 (N_8722,N_8479,N_8457);
nand U8723 (N_8723,N_8696,N_8456);
xnor U8724 (N_8724,N_8518,N_8548);
nor U8725 (N_8725,N_8688,N_8593);
or U8726 (N_8726,N_8474,N_8401);
nor U8727 (N_8727,N_8462,N_8638);
or U8728 (N_8728,N_8685,N_8622);
xor U8729 (N_8729,N_8425,N_8611);
and U8730 (N_8730,N_8530,N_8438);
or U8731 (N_8731,N_8630,N_8660);
nand U8732 (N_8732,N_8676,N_8419);
and U8733 (N_8733,N_8617,N_8512);
nor U8734 (N_8734,N_8525,N_8644);
and U8735 (N_8735,N_8675,N_8527);
nor U8736 (N_8736,N_8413,N_8648);
xor U8737 (N_8737,N_8540,N_8699);
nor U8738 (N_8738,N_8466,N_8449);
nor U8739 (N_8739,N_8624,N_8567);
or U8740 (N_8740,N_8475,N_8483);
nand U8741 (N_8741,N_8524,N_8687);
and U8742 (N_8742,N_8665,N_8646);
and U8743 (N_8743,N_8637,N_8534);
nand U8744 (N_8744,N_8561,N_8504);
nor U8745 (N_8745,N_8477,N_8600);
nand U8746 (N_8746,N_8532,N_8658);
xnor U8747 (N_8747,N_8545,N_8647);
or U8748 (N_8748,N_8608,N_8424);
or U8749 (N_8749,N_8664,N_8412);
or U8750 (N_8750,N_8410,N_8471);
xnor U8751 (N_8751,N_8436,N_8511);
and U8752 (N_8752,N_8501,N_8632);
nor U8753 (N_8753,N_8437,N_8552);
nor U8754 (N_8754,N_8543,N_8519);
nor U8755 (N_8755,N_8633,N_8686);
nor U8756 (N_8756,N_8693,N_8408);
and U8757 (N_8757,N_8592,N_8558);
and U8758 (N_8758,N_8431,N_8400);
and U8759 (N_8759,N_8440,N_8546);
nand U8760 (N_8760,N_8528,N_8553);
and U8761 (N_8761,N_8453,N_8426);
or U8762 (N_8762,N_8667,N_8577);
nor U8763 (N_8763,N_8490,N_8607);
nand U8764 (N_8764,N_8672,N_8616);
nand U8765 (N_8765,N_8522,N_8458);
and U8766 (N_8766,N_8520,N_8581);
nand U8767 (N_8767,N_8576,N_8486);
nor U8768 (N_8768,N_8694,N_8671);
or U8769 (N_8769,N_8678,N_8661);
and U8770 (N_8770,N_8418,N_8582);
nand U8771 (N_8771,N_8507,N_8485);
nand U8772 (N_8772,N_8692,N_8602);
or U8773 (N_8773,N_8621,N_8645);
nor U8774 (N_8774,N_8523,N_8429);
or U8775 (N_8775,N_8639,N_8407);
nand U8776 (N_8776,N_8683,N_8587);
nand U8777 (N_8777,N_8509,N_8533);
nor U8778 (N_8778,N_8650,N_8603);
nand U8779 (N_8779,N_8498,N_8599);
xor U8780 (N_8780,N_8409,N_8565);
nor U8781 (N_8781,N_8495,N_8690);
or U8782 (N_8782,N_8605,N_8497);
nand U8783 (N_8783,N_8516,N_8669);
and U8784 (N_8784,N_8591,N_8572);
and U8785 (N_8785,N_8443,N_8641);
or U8786 (N_8786,N_8657,N_8482);
or U8787 (N_8787,N_8555,N_8469);
xor U8788 (N_8788,N_8478,N_8689);
xnor U8789 (N_8789,N_8674,N_8405);
or U8790 (N_8790,N_8585,N_8557);
xor U8791 (N_8791,N_8406,N_8526);
nor U8792 (N_8792,N_8434,N_8554);
and U8793 (N_8793,N_8492,N_8514);
or U8794 (N_8794,N_8439,N_8515);
xnor U8795 (N_8795,N_8433,N_8564);
nor U8796 (N_8796,N_8489,N_8612);
nor U8797 (N_8797,N_8560,N_8503);
nor U8798 (N_8798,N_8470,N_8580);
and U8799 (N_8799,N_8573,N_8595);
nand U8800 (N_8800,N_8590,N_8691);
nor U8801 (N_8801,N_8448,N_8620);
xor U8802 (N_8802,N_8544,N_8467);
nand U8803 (N_8803,N_8662,N_8575);
xor U8804 (N_8804,N_8472,N_8626);
nor U8805 (N_8805,N_8653,N_8635);
xor U8806 (N_8806,N_8539,N_8420);
and U8807 (N_8807,N_8670,N_8627);
nor U8808 (N_8808,N_8484,N_8640);
nor U8809 (N_8809,N_8513,N_8655);
nor U8810 (N_8810,N_8571,N_8559);
nand U8811 (N_8811,N_8629,N_8542);
and U8812 (N_8812,N_8491,N_8451);
or U8813 (N_8813,N_8649,N_8417);
nand U8814 (N_8814,N_8428,N_8610);
nor U8815 (N_8815,N_8677,N_8673);
and U8816 (N_8816,N_8574,N_8547);
nor U8817 (N_8817,N_8666,N_8446);
and U8818 (N_8818,N_8614,N_8570);
or U8819 (N_8819,N_8403,N_8589);
nand U8820 (N_8820,N_8663,N_8698);
xor U8821 (N_8821,N_8569,N_8411);
nor U8822 (N_8822,N_8619,N_8615);
nor U8823 (N_8823,N_8427,N_8695);
or U8824 (N_8824,N_8441,N_8473);
and U8825 (N_8825,N_8421,N_8679);
or U8826 (N_8826,N_8505,N_8468);
nor U8827 (N_8827,N_8465,N_8681);
xor U8828 (N_8828,N_8461,N_8517);
or U8829 (N_8829,N_8423,N_8502);
nand U8830 (N_8830,N_8578,N_8529);
nand U8831 (N_8831,N_8680,N_8556);
nand U8832 (N_8832,N_8596,N_8432);
xor U8833 (N_8833,N_8609,N_8613);
or U8834 (N_8834,N_8586,N_8536);
nor U8835 (N_8835,N_8604,N_8499);
nor U8836 (N_8836,N_8625,N_8494);
nor U8837 (N_8837,N_8549,N_8651);
nand U8838 (N_8838,N_8682,N_8628);
and U8839 (N_8839,N_8634,N_8508);
and U8840 (N_8840,N_8510,N_8659);
nand U8841 (N_8841,N_8618,N_8444);
and U8842 (N_8842,N_8480,N_8447);
xnor U8843 (N_8843,N_8487,N_8584);
and U8844 (N_8844,N_8435,N_8642);
nor U8845 (N_8845,N_8488,N_8476);
nand U8846 (N_8846,N_8450,N_8531);
nand U8847 (N_8847,N_8481,N_8506);
or U8848 (N_8848,N_8563,N_8442);
nor U8849 (N_8849,N_8459,N_8537);
and U8850 (N_8850,N_8560,N_8573);
nor U8851 (N_8851,N_8618,N_8565);
nor U8852 (N_8852,N_8431,N_8478);
nand U8853 (N_8853,N_8690,N_8691);
and U8854 (N_8854,N_8630,N_8646);
xnor U8855 (N_8855,N_8404,N_8481);
and U8856 (N_8856,N_8581,N_8689);
nand U8857 (N_8857,N_8465,N_8691);
xor U8858 (N_8858,N_8696,N_8470);
nand U8859 (N_8859,N_8408,N_8688);
nor U8860 (N_8860,N_8517,N_8567);
nand U8861 (N_8861,N_8536,N_8631);
xnor U8862 (N_8862,N_8437,N_8576);
and U8863 (N_8863,N_8432,N_8551);
xor U8864 (N_8864,N_8413,N_8437);
and U8865 (N_8865,N_8585,N_8589);
nand U8866 (N_8866,N_8542,N_8490);
xnor U8867 (N_8867,N_8411,N_8689);
nand U8868 (N_8868,N_8432,N_8506);
and U8869 (N_8869,N_8607,N_8552);
xor U8870 (N_8870,N_8575,N_8471);
nor U8871 (N_8871,N_8611,N_8409);
and U8872 (N_8872,N_8404,N_8571);
nand U8873 (N_8873,N_8566,N_8633);
nand U8874 (N_8874,N_8607,N_8685);
nand U8875 (N_8875,N_8681,N_8618);
or U8876 (N_8876,N_8680,N_8544);
xnor U8877 (N_8877,N_8400,N_8496);
and U8878 (N_8878,N_8442,N_8514);
or U8879 (N_8879,N_8616,N_8687);
nand U8880 (N_8880,N_8625,N_8437);
nor U8881 (N_8881,N_8448,N_8654);
or U8882 (N_8882,N_8685,N_8584);
or U8883 (N_8883,N_8469,N_8501);
or U8884 (N_8884,N_8629,N_8679);
and U8885 (N_8885,N_8419,N_8569);
xnor U8886 (N_8886,N_8530,N_8644);
or U8887 (N_8887,N_8524,N_8471);
nand U8888 (N_8888,N_8637,N_8618);
xnor U8889 (N_8889,N_8652,N_8673);
nand U8890 (N_8890,N_8661,N_8641);
nor U8891 (N_8891,N_8504,N_8538);
or U8892 (N_8892,N_8613,N_8501);
nand U8893 (N_8893,N_8523,N_8479);
nand U8894 (N_8894,N_8422,N_8454);
xor U8895 (N_8895,N_8697,N_8413);
xnor U8896 (N_8896,N_8415,N_8527);
xnor U8897 (N_8897,N_8516,N_8465);
nor U8898 (N_8898,N_8443,N_8629);
and U8899 (N_8899,N_8444,N_8560);
nand U8900 (N_8900,N_8460,N_8418);
and U8901 (N_8901,N_8482,N_8452);
nand U8902 (N_8902,N_8684,N_8449);
nor U8903 (N_8903,N_8603,N_8653);
nor U8904 (N_8904,N_8472,N_8685);
nand U8905 (N_8905,N_8443,N_8442);
or U8906 (N_8906,N_8699,N_8507);
nand U8907 (N_8907,N_8532,N_8493);
xor U8908 (N_8908,N_8411,N_8476);
nor U8909 (N_8909,N_8511,N_8664);
and U8910 (N_8910,N_8648,N_8697);
nand U8911 (N_8911,N_8571,N_8445);
or U8912 (N_8912,N_8520,N_8640);
nand U8913 (N_8913,N_8575,N_8495);
or U8914 (N_8914,N_8638,N_8628);
nor U8915 (N_8915,N_8603,N_8549);
nor U8916 (N_8916,N_8495,N_8661);
and U8917 (N_8917,N_8692,N_8546);
and U8918 (N_8918,N_8404,N_8567);
or U8919 (N_8919,N_8494,N_8602);
or U8920 (N_8920,N_8595,N_8564);
xnor U8921 (N_8921,N_8469,N_8616);
or U8922 (N_8922,N_8566,N_8574);
and U8923 (N_8923,N_8548,N_8671);
nand U8924 (N_8924,N_8525,N_8517);
and U8925 (N_8925,N_8575,N_8597);
xor U8926 (N_8926,N_8647,N_8510);
and U8927 (N_8927,N_8554,N_8506);
nand U8928 (N_8928,N_8468,N_8694);
nor U8929 (N_8929,N_8537,N_8597);
nor U8930 (N_8930,N_8632,N_8509);
nand U8931 (N_8931,N_8604,N_8459);
xnor U8932 (N_8932,N_8600,N_8651);
nand U8933 (N_8933,N_8608,N_8442);
or U8934 (N_8934,N_8499,N_8699);
xor U8935 (N_8935,N_8610,N_8586);
nand U8936 (N_8936,N_8408,N_8557);
or U8937 (N_8937,N_8685,N_8545);
nand U8938 (N_8938,N_8589,N_8462);
and U8939 (N_8939,N_8527,N_8420);
xor U8940 (N_8940,N_8469,N_8690);
nand U8941 (N_8941,N_8698,N_8453);
xor U8942 (N_8942,N_8520,N_8565);
nor U8943 (N_8943,N_8696,N_8648);
nor U8944 (N_8944,N_8526,N_8472);
xor U8945 (N_8945,N_8647,N_8590);
and U8946 (N_8946,N_8613,N_8509);
nor U8947 (N_8947,N_8444,N_8676);
nand U8948 (N_8948,N_8694,N_8467);
nor U8949 (N_8949,N_8544,N_8671);
nand U8950 (N_8950,N_8587,N_8500);
nor U8951 (N_8951,N_8426,N_8636);
xnor U8952 (N_8952,N_8431,N_8463);
nor U8953 (N_8953,N_8404,N_8625);
nor U8954 (N_8954,N_8507,N_8519);
or U8955 (N_8955,N_8476,N_8445);
xor U8956 (N_8956,N_8545,N_8462);
nor U8957 (N_8957,N_8447,N_8494);
and U8958 (N_8958,N_8586,N_8607);
nand U8959 (N_8959,N_8518,N_8549);
or U8960 (N_8960,N_8676,N_8460);
or U8961 (N_8961,N_8688,N_8475);
and U8962 (N_8962,N_8576,N_8485);
nand U8963 (N_8963,N_8522,N_8641);
nor U8964 (N_8964,N_8634,N_8477);
and U8965 (N_8965,N_8646,N_8514);
nand U8966 (N_8966,N_8671,N_8665);
nor U8967 (N_8967,N_8606,N_8636);
and U8968 (N_8968,N_8578,N_8479);
xor U8969 (N_8969,N_8555,N_8556);
xor U8970 (N_8970,N_8602,N_8605);
xnor U8971 (N_8971,N_8631,N_8683);
xor U8972 (N_8972,N_8482,N_8662);
and U8973 (N_8973,N_8652,N_8638);
or U8974 (N_8974,N_8667,N_8529);
or U8975 (N_8975,N_8495,N_8478);
or U8976 (N_8976,N_8504,N_8531);
and U8977 (N_8977,N_8640,N_8495);
and U8978 (N_8978,N_8583,N_8636);
or U8979 (N_8979,N_8554,N_8555);
nor U8980 (N_8980,N_8559,N_8618);
nand U8981 (N_8981,N_8524,N_8691);
and U8982 (N_8982,N_8480,N_8400);
and U8983 (N_8983,N_8592,N_8619);
xnor U8984 (N_8984,N_8535,N_8629);
and U8985 (N_8985,N_8535,N_8677);
nor U8986 (N_8986,N_8548,N_8424);
and U8987 (N_8987,N_8601,N_8614);
xnor U8988 (N_8988,N_8631,N_8437);
and U8989 (N_8989,N_8417,N_8636);
or U8990 (N_8990,N_8674,N_8546);
nand U8991 (N_8991,N_8635,N_8497);
or U8992 (N_8992,N_8413,N_8581);
nor U8993 (N_8993,N_8531,N_8697);
nor U8994 (N_8994,N_8477,N_8604);
nand U8995 (N_8995,N_8410,N_8461);
nand U8996 (N_8996,N_8517,N_8677);
xor U8997 (N_8997,N_8676,N_8699);
xor U8998 (N_8998,N_8596,N_8684);
nor U8999 (N_8999,N_8661,N_8623);
xnor U9000 (N_9000,N_8986,N_8775);
nor U9001 (N_9001,N_8872,N_8883);
nor U9002 (N_9002,N_8847,N_8874);
nor U9003 (N_9003,N_8972,N_8752);
xor U9004 (N_9004,N_8702,N_8746);
and U9005 (N_9005,N_8837,N_8731);
xor U9006 (N_9006,N_8811,N_8794);
xor U9007 (N_9007,N_8768,N_8866);
nor U9008 (N_9008,N_8992,N_8817);
or U9009 (N_9009,N_8849,N_8922);
nand U9010 (N_9010,N_8877,N_8935);
xor U9011 (N_9011,N_8806,N_8818);
and U9012 (N_9012,N_8723,N_8982);
and U9013 (N_9013,N_8733,N_8782);
or U9014 (N_9014,N_8961,N_8748);
nor U9015 (N_9015,N_8893,N_8720);
nor U9016 (N_9016,N_8975,N_8984);
xor U9017 (N_9017,N_8985,N_8950);
nor U9018 (N_9018,N_8844,N_8708);
and U9019 (N_9019,N_8734,N_8842);
and U9020 (N_9020,N_8916,N_8846);
nand U9021 (N_9021,N_8960,N_8839);
xor U9022 (N_9022,N_8964,N_8716);
or U9023 (N_9023,N_8735,N_8741);
nand U9024 (N_9024,N_8882,N_8971);
and U9025 (N_9025,N_8946,N_8804);
nand U9026 (N_9026,N_8903,N_8925);
and U9027 (N_9027,N_8914,N_8881);
nand U9028 (N_9028,N_8906,N_8722);
nand U9029 (N_9029,N_8712,N_8875);
nor U9030 (N_9030,N_8841,N_8788);
or U9031 (N_9031,N_8711,N_8947);
nand U9032 (N_9032,N_8949,N_8802);
xnor U9033 (N_9033,N_8710,N_8776);
or U9034 (N_9034,N_8886,N_8803);
nand U9035 (N_9035,N_8999,N_8898);
or U9036 (N_9036,N_8828,N_8718);
nor U9037 (N_9037,N_8894,N_8765);
nand U9038 (N_9038,N_8927,N_8757);
or U9039 (N_9039,N_8742,N_8967);
xnor U9040 (N_9040,N_8853,N_8915);
nor U9041 (N_9041,N_8871,N_8879);
xnor U9042 (N_9042,N_8957,N_8890);
nor U9043 (N_9043,N_8850,N_8859);
or U9044 (N_9044,N_8709,N_8948);
nand U9045 (N_9045,N_8969,N_8807);
xnor U9046 (N_9046,N_8980,N_8873);
and U9047 (N_9047,N_8834,N_8705);
xnor U9048 (N_9048,N_8838,N_8825);
nor U9049 (N_9049,N_8848,N_8706);
nand U9050 (N_9050,N_8805,N_8988);
nor U9051 (N_9051,N_8885,N_8786);
nor U9052 (N_9052,N_8899,N_8700);
xor U9053 (N_9053,N_8815,N_8730);
nor U9054 (N_9054,N_8989,N_8816);
nand U9055 (N_9055,N_8767,N_8738);
or U9056 (N_9056,N_8981,N_8953);
or U9057 (N_9057,N_8789,N_8895);
nor U9058 (N_9058,N_8760,N_8926);
nor U9059 (N_9059,N_8778,N_8913);
and U9060 (N_9060,N_8819,N_8995);
nand U9061 (N_9061,N_8861,N_8756);
and U9062 (N_9062,N_8755,N_8833);
and U9063 (N_9063,N_8715,N_8860);
and U9064 (N_9064,N_8744,N_8973);
xnor U9065 (N_9065,N_8942,N_8729);
or U9066 (N_9066,N_8766,N_8704);
nor U9067 (N_9067,N_8707,N_8745);
xnor U9068 (N_9068,N_8905,N_8809);
or U9069 (N_9069,N_8996,N_8761);
nor U9070 (N_9070,N_8764,N_8884);
and U9071 (N_9071,N_8908,N_8897);
nand U9072 (N_9072,N_8824,N_8962);
or U9073 (N_9073,N_8901,N_8864);
xor U9074 (N_9074,N_8868,N_8772);
and U9075 (N_9075,N_8754,N_8959);
xor U9076 (N_9076,N_8714,N_8832);
and U9077 (N_9077,N_8936,N_8727);
nand U9078 (N_9078,N_8831,N_8880);
nor U9079 (N_9079,N_8790,N_8791);
nand U9080 (N_9080,N_8826,N_8867);
or U9081 (N_9081,N_8787,N_8813);
nand U9082 (N_9082,N_8854,N_8923);
nor U9083 (N_9083,N_8909,N_8750);
and U9084 (N_9084,N_8793,N_8934);
nor U9085 (N_9085,N_8919,N_8955);
xnor U9086 (N_9086,N_8954,N_8938);
xnor U9087 (N_9087,N_8974,N_8783);
nor U9088 (N_9088,N_8777,N_8940);
xnor U9089 (N_9089,N_8878,N_8944);
and U9090 (N_9090,N_8970,N_8845);
xnor U9091 (N_9091,N_8785,N_8751);
and U9092 (N_9092,N_8958,N_8758);
nand U9093 (N_9093,N_8943,N_8812);
nand U9094 (N_9094,N_8843,N_8869);
xnor U9095 (N_9095,N_8827,N_8997);
nand U9096 (N_9096,N_8798,N_8774);
xor U9097 (N_9097,N_8719,N_8945);
nor U9098 (N_9098,N_8726,N_8740);
or U9099 (N_9099,N_8852,N_8703);
nor U9100 (N_9100,N_8917,N_8814);
xor U9101 (N_9101,N_8952,N_8956);
xnor U9102 (N_9102,N_8921,N_8769);
xor U9103 (N_9103,N_8951,N_8737);
and U9104 (N_9104,N_8998,N_8931);
nor U9105 (N_9105,N_8763,N_8991);
and U9106 (N_9106,N_8924,N_8968);
and U9107 (N_9107,N_8732,N_8933);
and U9108 (N_9108,N_8990,N_8887);
nor U9109 (N_9109,N_8808,N_8979);
xnor U9110 (N_9110,N_8910,N_8835);
nor U9111 (N_9111,N_8963,N_8701);
or U9112 (N_9112,N_8784,N_8937);
or U9113 (N_9113,N_8918,N_8865);
or U9114 (N_9114,N_8771,N_8976);
xor U9115 (N_9115,N_8939,N_8840);
nor U9116 (N_9116,N_8994,N_8821);
nand U9117 (N_9117,N_8747,N_8965);
xnor U9118 (N_9118,N_8779,N_8888);
xor U9119 (N_9119,N_8823,N_8721);
nand U9120 (N_9120,N_8891,N_8770);
nand U9121 (N_9121,N_8912,N_8749);
nor U9122 (N_9122,N_8851,N_8858);
or U9123 (N_9123,N_8907,N_8930);
and U9124 (N_9124,N_8728,N_8941);
or U9125 (N_9125,N_8863,N_8724);
xnor U9126 (N_9126,N_8822,N_8773);
xnor U9127 (N_9127,N_8796,N_8792);
nor U9128 (N_9128,N_8799,N_8862);
nor U9129 (N_9129,N_8932,N_8736);
nor U9130 (N_9130,N_8800,N_8904);
and U9131 (N_9131,N_8753,N_8928);
nor U9132 (N_9132,N_8987,N_8830);
and U9133 (N_9133,N_8762,N_8713);
nor U9134 (N_9134,N_8900,N_8820);
nor U9135 (N_9135,N_8829,N_8836);
nor U9136 (N_9136,N_8725,N_8920);
and U9137 (N_9137,N_8966,N_8977);
and U9138 (N_9138,N_8857,N_8892);
and U9139 (N_9139,N_8993,N_8929);
or U9140 (N_9140,N_8810,N_8743);
nor U9141 (N_9141,N_8902,N_8876);
and U9142 (N_9142,N_8795,N_8717);
nor U9143 (N_9143,N_8781,N_8978);
nor U9144 (N_9144,N_8983,N_8889);
nor U9145 (N_9145,N_8780,N_8855);
nand U9146 (N_9146,N_8797,N_8856);
nand U9147 (N_9147,N_8870,N_8896);
and U9148 (N_9148,N_8759,N_8801);
nand U9149 (N_9149,N_8739,N_8911);
and U9150 (N_9150,N_8726,N_8948);
nor U9151 (N_9151,N_8773,N_8856);
nand U9152 (N_9152,N_8827,N_8927);
nor U9153 (N_9153,N_8860,N_8750);
xnor U9154 (N_9154,N_8731,N_8891);
and U9155 (N_9155,N_8921,N_8895);
or U9156 (N_9156,N_8864,N_8905);
nand U9157 (N_9157,N_8829,N_8825);
nand U9158 (N_9158,N_8986,N_8825);
nand U9159 (N_9159,N_8706,N_8704);
xnor U9160 (N_9160,N_8986,N_8895);
or U9161 (N_9161,N_8970,N_8828);
nand U9162 (N_9162,N_8869,N_8949);
or U9163 (N_9163,N_8788,N_8734);
and U9164 (N_9164,N_8887,N_8933);
or U9165 (N_9165,N_8912,N_8919);
or U9166 (N_9166,N_8772,N_8832);
and U9167 (N_9167,N_8820,N_8902);
or U9168 (N_9168,N_8896,N_8795);
and U9169 (N_9169,N_8933,N_8706);
or U9170 (N_9170,N_8777,N_8889);
nand U9171 (N_9171,N_8763,N_8813);
nand U9172 (N_9172,N_8711,N_8750);
nor U9173 (N_9173,N_8904,N_8995);
nand U9174 (N_9174,N_8752,N_8979);
xnor U9175 (N_9175,N_8762,N_8765);
or U9176 (N_9176,N_8868,N_8973);
nor U9177 (N_9177,N_8728,N_8708);
or U9178 (N_9178,N_8892,N_8837);
nand U9179 (N_9179,N_8957,N_8760);
nor U9180 (N_9180,N_8916,N_8872);
or U9181 (N_9181,N_8742,N_8948);
and U9182 (N_9182,N_8761,N_8729);
xor U9183 (N_9183,N_8929,N_8920);
nor U9184 (N_9184,N_8914,N_8823);
or U9185 (N_9185,N_8914,N_8933);
or U9186 (N_9186,N_8870,N_8710);
nor U9187 (N_9187,N_8732,N_8966);
or U9188 (N_9188,N_8916,N_8767);
or U9189 (N_9189,N_8970,N_8967);
or U9190 (N_9190,N_8855,N_8943);
xor U9191 (N_9191,N_8945,N_8777);
and U9192 (N_9192,N_8797,N_8929);
nand U9193 (N_9193,N_8993,N_8840);
or U9194 (N_9194,N_8886,N_8859);
nand U9195 (N_9195,N_8701,N_8983);
nor U9196 (N_9196,N_8927,N_8734);
xnor U9197 (N_9197,N_8713,N_8868);
or U9198 (N_9198,N_8719,N_8854);
and U9199 (N_9199,N_8836,N_8946);
and U9200 (N_9200,N_8969,N_8843);
xor U9201 (N_9201,N_8842,N_8973);
or U9202 (N_9202,N_8811,N_8916);
nor U9203 (N_9203,N_8984,N_8879);
or U9204 (N_9204,N_8907,N_8834);
or U9205 (N_9205,N_8946,N_8783);
nor U9206 (N_9206,N_8782,N_8750);
nand U9207 (N_9207,N_8760,N_8997);
xnor U9208 (N_9208,N_8794,N_8700);
xnor U9209 (N_9209,N_8816,N_8804);
and U9210 (N_9210,N_8908,N_8819);
and U9211 (N_9211,N_8703,N_8850);
xor U9212 (N_9212,N_8889,N_8968);
nor U9213 (N_9213,N_8880,N_8739);
nand U9214 (N_9214,N_8722,N_8749);
nor U9215 (N_9215,N_8733,N_8808);
nand U9216 (N_9216,N_8876,N_8888);
xnor U9217 (N_9217,N_8945,N_8828);
or U9218 (N_9218,N_8709,N_8733);
nor U9219 (N_9219,N_8721,N_8770);
and U9220 (N_9220,N_8761,N_8714);
xnor U9221 (N_9221,N_8996,N_8937);
nor U9222 (N_9222,N_8972,N_8769);
xnor U9223 (N_9223,N_8880,N_8898);
nor U9224 (N_9224,N_8703,N_8998);
or U9225 (N_9225,N_8783,N_8944);
xor U9226 (N_9226,N_8883,N_8756);
and U9227 (N_9227,N_8948,N_8918);
xor U9228 (N_9228,N_8766,N_8893);
nand U9229 (N_9229,N_8722,N_8761);
xnor U9230 (N_9230,N_8890,N_8807);
nand U9231 (N_9231,N_8754,N_8781);
nor U9232 (N_9232,N_8916,N_8714);
nor U9233 (N_9233,N_8790,N_8793);
nand U9234 (N_9234,N_8983,N_8772);
nand U9235 (N_9235,N_8783,N_8847);
xor U9236 (N_9236,N_8990,N_8917);
or U9237 (N_9237,N_8849,N_8962);
nand U9238 (N_9238,N_8793,N_8808);
and U9239 (N_9239,N_8954,N_8779);
or U9240 (N_9240,N_8919,N_8922);
or U9241 (N_9241,N_8952,N_8794);
or U9242 (N_9242,N_8955,N_8773);
xnor U9243 (N_9243,N_8880,N_8794);
xnor U9244 (N_9244,N_8814,N_8898);
nand U9245 (N_9245,N_8835,N_8853);
nand U9246 (N_9246,N_8917,N_8785);
and U9247 (N_9247,N_8986,N_8814);
nor U9248 (N_9248,N_8860,N_8841);
or U9249 (N_9249,N_8914,N_8757);
and U9250 (N_9250,N_8706,N_8796);
nor U9251 (N_9251,N_8893,N_8933);
nand U9252 (N_9252,N_8702,N_8709);
or U9253 (N_9253,N_8887,N_8924);
and U9254 (N_9254,N_8898,N_8893);
xnor U9255 (N_9255,N_8967,N_8722);
xnor U9256 (N_9256,N_8905,N_8726);
xnor U9257 (N_9257,N_8756,N_8753);
or U9258 (N_9258,N_8948,N_8999);
or U9259 (N_9259,N_8716,N_8824);
and U9260 (N_9260,N_8722,N_8754);
and U9261 (N_9261,N_8755,N_8895);
or U9262 (N_9262,N_8776,N_8733);
nor U9263 (N_9263,N_8759,N_8943);
and U9264 (N_9264,N_8904,N_8894);
xnor U9265 (N_9265,N_8937,N_8777);
or U9266 (N_9266,N_8880,N_8928);
nor U9267 (N_9267,N_8897,N_8775);
and U9268 (N_9268,N_8955,N_8716);
and U9269 (N_9269,N_8790,N_8838);
xnor U9270 (N_9270,N_8810,N_8952);
nor U9271 (N_9271,N_8920,N_8712);
xnor U9272 (N_9272,N_8853,N_8973);
or U9273 (N_9273,N_8922,N_8987);
and U9274 (N_9274,N_8977,N_8980);
or U9275 (N_9275,N_8916,N_8883);
or U9276 (N_9276,N_8812,N_8865);
and U9277 (N_9277,N_8804,N_8726);
or U9278 (N_9278,N_8911,N_8824);
xor U9279 (N_9279,N_8777,N_8793);
nor U9280 (N_9280,N_8881,N_8852);
and U9281 (N_9281,N_8829,N_8884);
or U9282 (N_9282,N_8922,N_8991);
or U9283 (N_9283,N_8871,N_8819);
nor U9284 (N_9284,N_8926,N_8836);
nand U9285 (N_9285,N_8925,N_8732);
nand U9286 (N_9286,N_8941,N_8706);
xor U9287 (N_9287,N_8704,N_8906);
and U9288 (N_9288,N_8853,N_8954);
or U9289 (N_9289,N_8961,N_8962);
nor U9290 (N_9290,N_8912,N_8799);
or U9291 (N_9291,N_8708,N_8778);
nor U9292 (N_9292,N_8920,N_8906);
or U9293 (N_9293,N_8823,N_8830);
nor U9294 (N_9294,N_8728,N_8715);
and U9295 (N_9295,N_8801,N_8890);
nand U9296 (N_9296,N_8981,N_8715);
nand U9297 (N_9297,N_8745,N_8878);
nor U9298 (N_9298,N_8717,N_8879);
or U9299 (N_9299,N_8960,N_8959);
or U9300 (N_9300,N_9129,N_9198);
nand U9301 (N_9301,N_9138,N_9202);
and U9302 (N_9302,N_9076,N_9005);
and U9303 (N_9303,N_9155,N_9180);
nand U9304 (N_9304,N_9050,N_9064);
nand U9305 (N_9305,N_9237,N_9099);
nor U9306 (N_9306,N_9094,N_9043);
nand U9307 (N_9307,N_9222,N_9269);
nand U9308 (N_9308,N_9022,N_9151);
xor U9309 (N_9309,N_9248,N_9046);
and U9310 (N_9310,N_9037,N_9068);
nand U9311 (N_9311,N_9108,N_9193);
or U9312 (N_9312,N_9058,N_9278);
or U9313 (N_9313,N_9103,N_9139);
and U9314 (N_9314,N_9072,N_9289);
nand U9315 (N_9315,N_9171,N_9090);
and U9316 (N_9316,N_9262,N_9261);
nor U9317 (N_9317,N_9002,N_9247);
xor U9318 (N_9318,N_9223,N_9128);
nor U9319 (N_9319,N_9297,N_9283);
xnor U9320 (N_9320,N_9086,N_9188);
or U9321 (N_9321,N_9294,N_9109);
nor U9322 (N_9322,N_9290,N_9275);
xnor U9323 (N_9323,N_9147,N_9277);
nor U9324 (N_9324,N_9291,N_9066);
and U9325 (N_9325,N_9210,N_9061);
xor U9326 (N_9326,N_9008,N_9161);
nor U9327 (N_9327,N_9246,N_9021);
nand U9328 (N_9328,N_9113,N_9007);
or U9329 (N_9329,N_9144,N_9150);
xor U9330 (N_9330,N_9203,N_9221);
and U9331 (N_9331,N_9231,N_9137);
xor U9332 (N_9332,N_9217,N_9204);
or U9333 (N_9333,N_9160,N_9131);
nand U9334 (N_9334,N_9084,N_9241);
nand U9335 (N_9335,N_9265,N_9228);
xor U9336 (N_9336,N_9256,N_9199);
nor U9337 (N_9337,N_9284,N_9266);
nand U9338 (N_9338,N_9238,N_9279);
or U9339 (N_9339,N_9006,N_9179);
or U9340 (N_9340,N_9140,N_9181);
nor U9341 (N_9341,N_9242,N_9148);
and U9342 (N_9342,N_9095,N_9239);
and U9343 (N_9343,N_9010,N_9166);
xnor U9344 (N_9344,N_9141,N_9184);
nor U9345 (N_9345,N_9127,N_9057);
nor U9346 (N_9346,N_9081,N_9101);
nor U9347 (N_9347,N_9153,N_9136);
and U9348 (N_9348,N_9017,N_9038);
nor U9349 (N_9349,N_9011,N_9115);
nor U9350 (N_9350,N_9102,N_9107);
nor U9351 (N_9351,N_9226,N_9078);
xor U9352 (N_9352,N_9192,N_9097);
and U9353 (N_9353,N_9167,N_9031);
xnor U9354 (N_9354,N_9287,N_9177);
or U9355 (N_9355,N_9253,N_9267);
or U9356 (N_9356,N_9168,N_9268);
xor U9357 (N_9357,N_9183,N_9232);
nand U9358 (N_9358,N_9118,N_9252);
or U9359 (N_9359,N_9030,N_9035);
nand U9360 (N_9360,N_9286,N_9083);
nand U9361 (N_9361,N_9062,N_9285);
nand U9362 (N_9362,N_9216,N_9276);
and U9363 (N_9363,N_9074,N_9132);
xnor U9364 (N_9364,N_9200,N_9004);
or U9365 (N_9365,N_9280,N_9234);
xor U9366 (N_9366,N_9055,N_9093);
or U9367 (N_9367,N_9213,N_9070);
or U9368 (N_9368,N_9048,N_9013);
nor U9369 (N_9369,N_9026,N_9196);
nand U9370 (N_9370,N_9163,N_9025);
xor U9371 (N_9371,N_9045,N_9032);
nor U9372 (N_9372,N_9236,N_9034);
or U9373 (N_9373,N_9014,N_9251);
xor U9374 (N_9374,N_9172,N_9225);
xnor U9375 (N_9375,N_9077,N_9119);
xnor U9376 (N_9376,N_9096,N_9130);
xnor U9377 (N_9377,N_9124,N_9000);
and U9378 (N_9378,N_9069,N_9281);
xnor U9379 (N_9379,N_9075,N_9067);
or U9380 (N_9380,N_9159,N_9092);
xnor U9381 (N_9381,N_9040,N_9257);
xor U9382 (N_9382,N_9133,N_9015);
nand U9383 (N_9383,N_9080,N_9047);
nand U9384 (N_9384,N_9125,N_9149);
nor U9385 (N_9385,N_9001,N_9170);
nor U9386 (N_9386,N_9063,N_9110);
or U9387 (N_9387,N_9121,N_9174);
or U9388 (N_9388,N_9263,N_9016);
nor U9389 (N_9389,N_9089,N_9197);
xor U9390 (N_9390,N_9208,N_9056);
xnor U9391 (N_9391,N_9027,N_9003);
or U9392 (N_9392,N_9191,N_9162);
xor U9393 (N_9393,N_9215,N_9165);
and U9394 (N_9394,N_9088,N_9255);
and U9395 (N_9395,N_9189,N_9049);
and U9396 (N_9396,N_9019,N_9041);
nor U9397 (N_9397,N_9206,N_9085);
and U9398 (N_9398,N_9274,N_9134);
xnor U9399 (N_9399,N_9036,N_9227);
xnor U9400 (N_9400,N_9024,N_9187);
nand U9401 (N_9401,N_9194,N_9106);
xnor U9402 (N_9402,N_9243,N_9218);
nor U9403 (N_9403,N_9271,N_9100);
and U9404 (N_9404,N_9028,N_9135);
nand U9405 (N_9405,N_9259,N_9122);
nand U9406 (N_9406,N_9186,N_9173);
or U9407 (N_9407,N_9065,N_9178);
and U9408 (N_9408,N_9020,N_9249);
nand U9409 (N_9409,N_9288,N_9211);
xnor U9410 (N_9410,N_9156,N_9052);
nand U9411 (N_9411,N_9229,N_9120);
and U9412 (N_9412,N_9207,N_9042);
and U9413 (N_9413,N_9182,N_9176);
or U9414 (N_9414,N_9082,N_9114);
xnor U9415 (N_9415,N_9250,N_9087);
nand U9416 (N_9416,N_9091,N_9212);
xor U9417 (N_9417,N_9264,N_9012);
xnor U9418 (N_9418,N_9111,N_9146);
and U9419 (N_9419,N_9220,N_9235);
and U9420 (N_9420,N_9143,N_9071);
and U9421 (N_9421,N_9023,N_9009);
and U9422 (N_9422,N_9272,N_9190);
nand U9423 (N_9423,N_9299,N_9039);
and U9424 (N_9424,N_9105,N_9018);
xor U9425 (N_9425,N_9126,N_9154);
and U9426 (N_9426,N_9054,N_9164);
nand U9427 (N_9427,N_9185,N_9104);
nor U9428 (N_9428,N_9033,N_9152);
and U9429 (N_9429,N_9158,N_9175);
or U9430 (N_9430,N_9292,N_9296);
xnor U9431 (N_9431,N_9293,N_9245);
nand U9432 (N_9432,N_9209,N_9273);
xnor U9433 (N_9433,N_9098,N_9240);
or U9434 (N_9434,N_9254,N_9282);
nand U9435 (N_9435,N_9295,N_9051);
or U9436 (N_9436,N_9157,N_9053);
or U9437 (N_9437,N_9079,N_9270);
and U9438 (N_9438,N_9044,N_9230);
nor U9439 (N_9439,N_9258,N_9201);
and U9440 (N_9440,N_9195,N_9219);
or U9441 (N_9441,N_9214,N_9205);
xnor U9442 (N_9442,N_9117,N_9123);
nor U9443 (N_9443,N_9059,N_9224);
nor U9444 (N_9444,N_9233,N_9073);
or U9445 (N_9445,N_9260,N_9029);
and U9446 (N_9446,N_9112,N_9169);
nor U9447 (N_9447,N_9145,N_9060);
xor U9448 (N_9448,N_9116,N_9244);
or U9449 (N_9449,N_9142,N_9298);
xor U9450 (N_9450,N_9291,N_9288);
or U9451 (N_9451,N_9167,N_9143);
nand U9452 (N_9452,N_9252,N_9131);
nor U9453 (N_9453,N_9069,N_9265);
nand U9454 (N_9454,N_9182,N_9017);
nor U9455 (N_9455,N_9128,N_9282);
or U9456 (N_9456,N_9086,N_9255);
nand U9457 (N_9457,N_9027,N_9186);
and U9458 (N_9458,N_9047,N_9183);
or U9459 (N_9459,N_9154,N_9004);
nand U9460 (N_9460,N_9141,N_9242);
and U9461 (N_9461,N_9145,N_9058);
nand U9462 (N_9462,N_9191,N_9112);
xnor U9463 (N_9463,N_9101,N_9255);
xnor U9464 (N_9464,N_9203,N_9234);
nor U9465 (N_9465,N_9053,N_9162);
nand U9466 (N_9466,N_9117,N_9170);
or U9467 (N_9467,N_9009,N_9177);
xnor U9468 (N_9468,N_9094,N_9218);
nor U9469 (N_9469,N_9231,N_9091);
or U9470 (N_9470,N_9180,N_9061);
and U9471 (N_9471,N_9075,N_9124);
nand U9472 (N_9472,N_9082,N_9013);
or U9473 (N_9473,N_9048,N_9297);
nor U9474 (N_9474,N_9103,N_9149);
and U9475 (N_9475,N_9089,N_9212);
xnor U9476 (N_9476,N_9160,N_9197);
nor U9477 (N_9477,N_9177,N_9214);
or U9478 (N_9478,N_9058,N_9134);
xnor U9479 (N_9479,N_9022,N_9156);
xor U9480 (N_9480,N_9032,N_9200);
and U9481 (N_9481,N_9261,N_9232);
and U9482 (N_9482,N_9047,N_9209);
or U9483 (N_9483,N_9063,N_9031);
xnor U9484 (N_9484,N_9277,N_9136);
nand U9485 (N_9485,N_9070,N_9030);
nor U9486 (N_9486,N_9249,N_9054);
nor U9487 (N_9487,N_9044,N_9110);
or U9488 (N_9488,N_9031,N_9224);
xnor U9489 (N_9489,N_9167,N_9136);
or U9490 (N_9490,N_9206,N_9004);
xnor U9491 (N_9491,N_9195,N_9189);
nor U9492 (N_9492,N_9251,N_9272);
xor U9493 (N_9493,N_9194,N_9271);
and U9494 (N_9494,N_9277,N_9101);
nor U9495 (N_9495,N_9033,N_9190);
and U9496 (N_9496,N_9224,N_9070);
and U9497 (N_9497,N_9065,N_9250);
nor U9498 (N_9498,N_9060,N_9152);
nand U9499 (N_9499,N_9230,N_9226);
and U9500 (N_9500,N_9221,N_9156);
nor U9501 (N_9501,N_9091,N_9253);
and U9502 (N_9502,N_9074,N_9212);
or U9503 (N_9503,N_9275,N_9113);
or U9504 (N_9504,N_9122,N_9216);
and U9505 (N_9505,N_9042,N_9094);
nand U9506 (N_9506,N_9060,N_9013);
and U9507 (N_9507,N_9073,N_9154);
and U9508 (N_9508,N_9058,N_9289);
xor U9509 (N_9509,N_9200,N_9193);
nor U9510 (N_9510,N_9033,N_9057);
nor U9511 (N_9511,N_9241,N_9140);
nor U9512 (N_9512,N_9253,N_9062);
nor U9513 (N_9513,N_9142,N_9197);
nand U9514 (N_9514,N_9164,N_9249);
or U9515 (N_9515,N_9198,N_9117);
xnor U9516 (N_9516,N_9107,N_9053);
and U9517 (N_9517,N_9072,N_9063);
xnor U9518 (N_9518,N_9257,N_9205);
and U9519 (N_9519,N_9124,N_9014);
and U9520 (N_9520,N_9199,N_9242);
nor U9521 (N_9521,N_9260,N_9086);
nand U9522 (N_9522,N_9146,N_9272);
xnor U9523 (N_9523,N_9278,N_9203);
nand U9524 (N_9524,N_9028,N_9043);
or U9525 (N_9525,N_9104,N_9285);
nor U9526 (N_9526,N_9037,N_9171);
nor U9527 (N_9527,N_9117,N_9137);
nand U9528 (N_9528,N_9028,N_9060);
xnor U9529 (N_9529,N_9262,N_9165);
xor U9530 (N_9530,N_9194,N_9262);
nand U9531 (N_9531,N_9245,N_9266);
nand U9532 (N_9532,N_9068,N_9159);
or U9533 (N_9533,N_9045,N_9206);
nor U9534 (N_9534,N_9260,N_9143);
xnor U9535 (N_9535,N_9240,N_9116);
or U9536 (N_9536,N_9234,N_9161);
or U9537 (N_9537,N_9297,N_9287);
nor U9538 (N_9538,N_9060,N_9226);
and U9539 (N_9539,N_9049,N_9124);
or U9540 (N_9540,N_9137,N_9203);
or U9541 (N_9541,N_9183,N_9136);
and U9542 (N_9542,N_9005,N_9208);
nor U9543 (N_9543,N_9012,N_9186);
xor U9544 (N_9544,N_9151,N_9224);
xnor U9545 (N_9545,N_9019,N_9252);
and U9546 (N_9546,N_9021,N_9118);
xor U9547 (N_9547,N_9221,N_9261);
nand U9548 (N_9548,N_9123,N_9023);
nor U9549 (N_9549,N_9151,N_9128);
nor U9550 (N_9550,N_9081,N_9270);
and U9551 (N_9551,N_9186,N_9200);
xor U9552 (N_9552,N_9298,N_9007);
nor U9553 (N_9553,N_9168,N_9233);
or U9554 (N_9554,N_9116,N_9142);
or U9555 (N_9555,N_9074,N_9170);
nand U9556 (N_9556,N_9123,N_9108);
or U9557 (N_9557,N_9097,N_9282);
nand U9558 (N_9558,N_9160,N_9220);
nor U9559 (N_9559,N_9180,N_9065);
xor U9560 (N_9560,N_9278,N_9207);
nand U9561 (N_9561,N_9113,N_9273);
xor U9562 (N_9562,N_9154,N_9138);
nor U9563 (N_9563,N_9095,N_9106);
nand U9564 (N_9564,N_9172,N_9186);
and U9565 (N_9565,N_9127,N_9036);
or U9566 (N_9566,N_9170,N_9284);
nor U9567 (N_9567,N_9245,N_9097);
nor U9568 (N_9568,N_9140,N_9029);
nor U9569 (N_9569,N_9287,N_9135);
or U9570 (N_9570,N_9067,N_9173);
xor U9571 (N_9571,N_9178,N_9052);
nor U9572 (N_9572,N_9298,N_9180);
and U9573 (N_9573,N_9249,N_9282);
and U9574 (N_9574,N_9046,N_9066);
nand U9575 (N_9575,N_9138,N_9134);
and U9576 (N_9576,N_9106,N_9282);
nor U9577 (N_9577,N_9066,N_9083);
xnor U9578 (N_9578,N_9139,N_9094);
nand U9579 (N_9579,N_9065,N_9215);
nand U9580 (N_9580,N_9004,N_9032);
nand U9581 (N_9581,N_9085,N_9139);
or U9582 (N_9582,N_9265,N_9037);
and U9583 (N_9583,N_9181,N_9139);
nand U9584 (N_9584,N_9064,N_9282);
xor U9585 (N_9585,N_9049,N_9042);
nor U9586 (N_9586,N_9293,N_9135);
and U9587 (N_9587,N_9135,N_9151);
xnor U9588 (N_9588,N_9191,N_9116);
and U9589 (N_9589,N_9219,N_9247);
nor U9590 (N_9590,N_9172,N_9217);
nand U9591 (N_9591,N_9213,N_9104);
or U9592 (N_9592,N_9023,N_9150);
and U9593 (N_9593,N_9046,N_9152);
and U9594 (N_9594,N_9094,N_9148);
nand U9595 (N_9595,N_9089,N_9003);
or U9596 (N_9596,N_9157,N_9073);
xor U9597 (N_9597,N_9287,N_9153);
nand U9598 (N_9598,N_9205,N_9050);
and U9599 (N_9599,N_9267,N_9034);
or U9600 (N_9600,N_9481,N_9360);
and U9601 (N_9601,N_9316,N_9414);
nand U9602 (N_9602,N_9405,N_9433);
or U9603 (N_9603,N_9324,N_9581);
or U9604 (N_9604,N_9341,N_9458);
nor U9605 (N_9605,N_9514,N_9484);
nor U9606 (N_9606,N_9544,N_9353);
and U9607 (N_9607,N_9529,N_9462);
and U9608 (N_9608,N_9432,N_9317);
nand U9609 (N_9609,N_9323,N_9322);
and U9610 (N_9610,N_9493,N_9496);
or U9611 (N_9611,N_9564,N_9314);
and U9612 (N_9612,N_9446,N_9315);
nand U9613 (N_9613,N_9318,N_9460);
nand U9614 (N_9614,N_9569,N_9371);
nand U9615 (N_9615,N_9457,N_9557);
xnor U9616 (N_9616,N_9369,N_9494);
or U9617 (N_9617,N_9308,N_9395);
or U9618 (N_9618,N_9391,N_9503);
xnor U9619 (N_9619,N_9389,N_9358);
nor U9620 (N_9620,N_9438,N_9357);
and U9621 (N_9621,N_9429,N_9513);
nor U9622 (N_9622,N_9576,N_9392);
nor U9623 (N_9623,N_9593,N_9393);
xor U9624 (N_9624,N_9472,N_9586);
and U9625 (N_9625,N_9394,N_9597);
or U9626 (N_9626,N_9455,N_9338);
and U9627 (N_9627,N_9594,N_9456);
xnor U9628 (N_9628,N_9304,N_9373);
and U9629 (N_9629,N_9319,N_9473);
and U9630 (N_9630,N_9443,N_9554);
or U9631 (N_9631,N_9583,N_9363);
xor U9632 (N_9632,N_9515,N_9431);
xnor U9633 (N_9633,N_9582,N_9374);
nand U9634 (N_9634,N_9417,N_9459);
nor U9635 (N_9635,N_9483,N_9384);
or U9636 (N_9636,N_9416,N_9528);
xnor U9637 (N_9637,N_9587,N_9420);
xnor U9638 (N_9638,N_9495,N_9300);
or U9639 (N_9639,N_9551,N_9359);
xnor U9640 (N_9640,N_9599,N_9535);
nor U9641 (N_9641,N_9592,N_9453);
xor U9642 (N_9642,N_9388,N_9510);
or U9643 (N_9643,N_9509,N_9415);
and U9644 (N_9644,N_9356,N_9502);
or U9645 (N_9645,N_9465,N_9355);
or U9646 (N_9646,N_9546,N_9596);
nand U9647 (N_9647,N_9404,N_9320);
and U9648 (N_9648,N_9452,N_9331);
nand U9649 (N_9649,N_9342,N_9590);
and U9650 (N_9650,N_9476,N_9306);
nor U9651 (N_9651,N_9527,N_9497);
or U9652 (N_9652,N_9367,N_9343);
nor U9653 (N_9653,N_9467,N_9567);
nor U9654 (N_9654,N_9463,N_9517);
xnor U9655 (N_9655,N_9553,N_9425);
xnor U9656 (N_9656,N_9507,N_9534);
nand U9657 (N_9657,N_9475,N_9408);
and U9658 (N_9658,N_9538,N_9570);
nor U9659 (N_9659,N_9488,N_9519);
xnor U9660 (N_9660,N_9589,N_9485);
xor U9661 (N_9661,N_9327,N_9337);
xnor U9662 (N_9662,N_9444,N_9464);
or U9663 (N_9663,N_9500,N_9411);
nand U9664 (N_9664,N_9413,N_9498);
xor U9665 (N_9665,N_9402,N_9346);
nand U9666 (N_9666,N_9365,N_9491);
xnor U9667 (N_9667,N_9435,N_9563);
nor U9668 (N_9668,N_9577,N_9386);
xor U9669 (N_9669,N_9480,N_9526);
nor U9670 (N_9670,N_9471,N_9328);
nor U9671 (N_9671,N_9440,N_9591);
nand U9672 (N_9672,N_9424,N_9301);
xor U9673 (N_9673,N_9504,N_9451);
xor U9674 (N_9674,N_9518,N_9347);
xor U9675 (N_9675,N_9409,N_9558);
or U9676 (N_9676,N_9313,N_9489);
nand U9677 (N_9677,N_9520,N_9348);
and U9678 (N_9678,N_9545,N_9580);
xor U9679 (N_9679,N_9536,N_9382);
xor U9680 (N_9680,N_9366,N_9506);
xor U9681 (N_9681,N_9321,N_9378);
or U9682 (N_9682,N_9543,N_9352);
or U9683 (N_9683,N_9430,N_9379);
and U9684 (N_9684,N_9312,N_9548);
or U9685 (N_9685,N_9501,N_9588);
or U9686 (N_9686,N_9595,N_9561);
xnor U9687 (N_9687,N_9533,N_9585);
nand U9688 (N_9688,N_9449,N_9335);
or U9689 (N_9689,N_9511,N_9550);
nand U9690 (N_9690,N_9372,N_9436);
nor U9691 (N_9691,N_9336,N_9499);
or U9692 (N_9692,N_9547,N_9364);
nand U9693 (N_9693,N_9428,N_9477);
and U9694 (N_9694,N_9571,N_9445);
or U9695 (N_9695,N_9385,N_9562);
xor U9696 (N_9696,N_9530,N_9383);
and U9697 (N_9697,N_9361,N_9325);
xor U9698 (N_9698,N_9339,N_9486);
xnor U9699 (N_9699,N_9351,N_9332);
or U9700 (N_9700,N_9397,N_9419);
or U9701 (N_9701,N_9540,N_9447);
xor U9702 (N_9702,N_9302,N_9375);
or U9703 (N_9703,N_9354,N_9478);
and U9704 (N_9704,N_9390,N_9349);
xnor U9705 (N_9705,N_9406,N_9307);
or U9706 (N_9706,N_9555,N_9454);
xnor U9707 (N_9707,N_9303,N_9552);
nand U9708 (N_9708,N_9334,N_9512);
nand U9709 (N_9709,N_9423,N_9568);
xor U9710 (N_9710,N_9565,N_9575);
or U9711 (N_9711,N_9524,N_9434);
nand U9712 (N_9712,N_9466,N_9377);
xor U9713 (N_9713,N_9468,N_9407);
nor U9714 (N_9714,N_9398,N_9400);
and U9715 (N_9715,N_9560,N_9345);
nor U9716 (N_9716,N_9556,N_9559);
nor U9717 (N_9717,N_9329,N_9549);
or U9718 (N_9718,N_9450,N_9508);
or U9719 (N_9719,N_9523,N_9525);
and U9720 (N_9720,N_9412,N_9309);
xnor U9721 (N_9721,N_9441,N_9469);
nor U9722 (N_9722,N_9310,N_9492);
nand U9723 (N_9723,N_9396,N_9461);
nor U9724 (N_9724,N_9573,N_9479);
xor U9725 (N_9725,N_9566,N_9410);
or U9726 (N_9726,N_9344,N_9532);
nand U9727 (N_9727,N_9537,N_9574);
nand U9728 (N_9728,N_9387,N_9539);
nand U9729 (N_9729,N_9401,N_9305);
nand U9730 (N_9730,N_9376,N_9437);
nand U9731 (N_9731,N_9418,N_9362);
and U9732 (N_9732,N_9370,N_9579);
and U9733 (N_9733,N_9521,N_9522);
xnor U9734 (N_9734,N_9541,N_9427);
or U9735 (N_9735,N_9482,N_9531);
nor U9736 (N_9736,N_9403,N_9380);
xor U9737 (N_9737,N_9330,N_9474);
nor U9738 (N_9738,N_9368,N_9542);
or U9739 (N_9739,N_9487,N_9442);
nor U9740 (N_9740,N_9311,N_9490);
and U9741 (N_9741,N_9439,N_9381);
nor U9742 (N_9742,N_9399,N_9516);
xnor U9743 (N_9743,N_9333,N_9505);
nand U9744 (N_9744,N_9326,N_9598);
and U9745 (N_9745,N_9572,N_9470);
nand U9746 (N_9746,N_9422,N_9578);
or U9747 (N_9747,N_9421,N_9426);
nor U9748 (N_9748,N_9584,N_9350);
nand U9749 (N_9749,N_9340,N_9448);
nor U9750 (N_9750,N_9304,N_9402);
xor U9751 (N_9751,N_9569,N_9415);
xor U9752 (N_9752,N_9495,N_9337);
nor U9753 (N_9753,N_9483,N_9594);
nor U9754 (N_9754,N_9432,N_9446);
xnor U9755 (N_9755,N_9492,N_9363);
nand U9756 (N_9756,N_9591,N_9358);
and U9757 (N_9757,N_9558,N_9555);
xor U9758 (N_9758,N_9409,N_9425);
nand U9759 (N_9759,N_9545,N_9494);
and U9760 (N_9760,N_9568,N_9305);
xor U9761 (N_9761,N_9512,N_9411);
xnor U9762 (N_9762,N_9524,N_9469);
or U9763 (N_9763,N_9582,N_9580);
and U9764 (N_9764,N_9578,N_9582);
or U9765 (N_9765,N_9523,N_9564);
nand U9766 (N_9766,N_9393,N_9492);
xor U9767 (N_9767,N_9425,N_9350);
xnor U9768 (N_9768,N_9418,N_9501);
and U9769 (N_9769,N_9432,N_9441);
nand U9770 (N_9770,N_9515,N_9379);
or U9771 (N_9771,N_9536,N_9325);
and U9772 (N_9772,N_9545,N_9365);
nand U9773 (N_9773,N_9545,N_9515);
and U9774 (N_9774,N_9533,N_9352);
and U9775 (N_9775,N_9315,N_9598);
xor U9776 (N_9776,N_9306,N_9598);
or U9777 (N_9777,N_9458,N_9472);
or U9778 (N_9778,N_9463,N_9343);
nand U9779 (N_9779,N_9438,N_9463);
nand U9780 (N_9780,N_9370,N_9563);
xor U9781 (N_9781,N_9411,N_9441);
xnor U9782 (N_9782,N_9306,N_9554);
and U9783 (N_9783,N_9313,N_9533);
nor U9784 (N_9784,N_9535,N_9320);
nor U9785 (N_9785,N_9518,N_9407);
xor U9786 (N_9786,N_9589,N_9384);
nor U9787 (N_9787,N_9472,N_9317);
and U9788 (N_9788,N_9585,N_9364);
and U9789 (N_9789,N_9393,N_9474);
and U9790 (N_9790,N_9312,N_9441);
and U9791 (N_9791,N_9330,N_9401);
or U9792 (N_9792,N_9556,N_9431);
or U9793 (N_9793,N_9322,N_9305);
and U9794 (N_9794,N_9502,N_9318);
and U9795 (N_9795,N_9485,N_9372);
nand U9796 (N_9796,N_9577,N_9558);
or U9797 (N_9797,N_9516,N_9452);
or U9798 (N_9798,N_9305,N_9339);
nor U9799 (N_9799,N_9438,N_9589);
or U9800 (N_9800,N_9318,N_9466);
xnor U9801 (N_9801,N_9348,N_9307);
and U9802 (N_9802,N_9385,N_9541);
and U9803 (N_9803,N_9406,N_9399);
xor U9804 (N_9804,N_9404,N_9462);
nor U9805 (N_9805,N_9486,N_9452);
xnor U9806 (N_9806,N_9522,N_9476);
and U9807 (N_9807,N_9431,N_9533);
nor U9808 (N_9808,N_9306,N_9470);
or U9809 (N_9809,N_9395,N_9317);
nand U9810 (N_9810,N_9505,N_9362);
or U9811 (N_9811,N_9428,N_9480);
or U9812 (N_9812,N_9386,N_9540);
and U9813 (N_9813,N_9327,N_9531);
nand U9814 (N_9814,N_9386,N_9517);
or U9815 (N_9815,N_9318,N_9446);
or U9816 (N_9816,N_9302,N_9548);
xnor U9817 (N_9817,N_9445,N_9493);
or U9818 (N_9818,N_9440,N_9584);
or U9819 (N_9819,N_9452,N_9598);
xnor U9820 (N_9820,N_9506,N_9420);
or U9821 (N_9821,N_9528,N_9432);
or U9822 (N_9822,N_9585,N_9405);
nor U9823 (N_9823,N_9421,N_9326);
nand U9824 (N_9824,N_9335,N_9315);
or U9825 (N_9825,N_9428,N_9435);
nor U9826 (N_9826,N_9479,N_9477);
and U9827 (N_9827,N_9396,N_9311);
xnor U9828 (N_9828,N_9344,N_9329);
and U9829 (N_9829,N_9580,N_9502);
xnor U9830 (N_9830,N_9413,N_9404);
nor U9831 (N_9831,N_9509,N_9409);
nor U9832 (N_9832,N_9464,N_9442);
nor U9833 (N_9833,N_9526,N_9497);
and U9834 (N_9834,N_9356,N_9340);
nor U9835 (N_9835,N_9514,N_9535);
nor U9836 (N_9836,N_9343,N_9455);
or U9837 (N_9837,N_9441,N_9345);
and U9838 (N_9838,N_9571,N_9529);
or U9839 (N_9839,N_9457,N_9373);
and U9840 (N_9840,N_9351,N_9457);
xor U9841 (N_9841,N_9470,N_9567);
nor U9842 (N_9842,N_9533,N_9329);
and U9843 (N_9843,N_9453,N_9588);
xnor U9844 (N_9844,N_9439,N_9584);
xnor U9845 (N_9845,N_9402,N_9535);
and U9846 (N_9846,N_9410,N_9567);
nor U9847 (N_9847,N_9518,N_9596);
nand U9848 (N_9848,N_9565,N_9320);
or U9849 (N_9849,N_9446,N_9476);
nand U9850 (N_9850,N_9385,N_9461);
nand U9851 (N_9851,N_9400,N_9415);
nor U9852 (N_9852,N_9368,N_9515);
and U9853 (N_9853,N_9330,N_9348);
and U9854 (N_9854,N_9402,N_9532);
xnor U9855 (N_9855,N_9347,N_9346);
nand U9856 (N_9856,N_9563,N_9559);
or U9857 (N_9857,N_9495,N_9539);
or U9858 (N_9858,N_9455,N_9440);
nor U9859 (N_9859,N_9508,N_9552);
nor U9860 (N_9860,N_9405,N_9314);
nor U9861 (N_9861,N_9468,N_9539);
nor U9862 (N_9862,N_9433,N_9503);
or U9863 (N_9863,N_9481,N_9398);
nor U9864 (N_9864,N_9388,N_9374);
nor U9865 (N_9865,N_9520,N_9432);
nor U9866 (N_9866,N_9592,N_9552);
and U9867 (N_9867,N_9457,N_9422);
nor U9868 (N_9868,N_9569,N_9473);
nand U9869 (N_9869,N_9303,N_9483);
or U9870 (N_9870,N_9398,N_9414);
xnor U9871 (N_9871,N_9472,N_9502);
and U9872 (N_9872,N_9347,N_9302);
nor U9873 (N_9873,N_9463,N_9361);
or U9874 (N_9874,N_9356,N_9324);
nand U9875 (N_9875,N_9325,N_9335);
and U9876 (N_9876,N_9433,N_9345);
and U9877 (N_9877,N_9302,N_9447);
nor U9878 (N_9878,N_9302,N_9499);
nand U9879 (N_9879,N_9510,N_9381);
xor U9880 (N_9880,N_9323,N_9311);
nand U9881 (N_9881,N_9521,N_9398);
nand U9882 (N_9882,N_9586,N_9464);
and U9883 (N_9883,N_9596,N_9566);
nand U9884 (N_9884,N_9516,N_9545);
nor U9885 (N_9885,N_9336,N_9592);
nor U9886 (N_9886,N_9574,N_9568);
xnor U9887 (N_9887,N_9305,N_9383);
or U9888 (N_9888,N_9440,N_9599);
nor U9889 (N_9889,N_9481,N_9483);
or U9890 (N_9890,N_9573,N_9579);
nand U9891 (N_9891,N_9521,N_9460);
nand U9892 (N_9892,N_9413,N_9500);
xnor U9893 (N_9893,N_9573,N_9490);
nand U9894 (N_9894,N_9535,N_9325);
or U9895 (N_9895,N_9573,N_9494);
or U9896 (N_9896,N_9562,N_9357);
nand U9897 (N_9897,N_9508,N_9415);
nor U9898 (N_9898,N_9462,N_9328);
nand U9899 (N_9899,N_9415,N_9574);
or U9900 (N_9900,N_9855,N_9680);
nor U9901 (N_9901,N_9856,N_9668);
and U9902 (N_9902,N_9811,N_9741);
xnor U9903 (N_9903,N_9871,N_9842);
and U9904 (N_9904,N_9647,N_9733);
xnor U9905 (N_9905,N_9762,N_9663);
nand U9906 (N_9906,N_9694,N_9667);
xnor U9907 (N_9907,N_9878,N_9675);
xnor U9908 (N_9908,N_9773,N_9823);
and U9909 (N_9909,N_9784,N_9777);
nand U9910 (N_9910,N_9779,N_9879);
nand U9911 (N_9911,N_9833,N_9843);
xnor U9912 (N_9912,N_9854,N_9845);
nor U9913 (N_9913,N_9883,N_9793);
nor U9914 (N_9914,N_9660,N_9665);
nor U9915 (N_9915,N_9635,N_9723);
xor U9916 (N_9916,N_9863,N_9600);
nand U9917 (N_9917,N_9791,N_9801);
nand U9918 (N_9918,N_9829,N_9656);
nand U9919 (N_9919,N_9673,N_9857);
xnor U9920 (N_9920,N_9753,N_9848);
or U9921 (N_9921,N_9804,N_9818);
xnor U9922 (N_9922,N_9807,N_9729);
xor U9923 (N_9923,N_9870,N_9638);
nand U9924 (N_9924,N_9698,N_9825);
or U9925 (N_9925,N_9645,N_9880);
and U9926 (N_9926,N_9712,N_9744);
or U9927 (N_9927,N_9882,N_9742);
or U9928 (N_9928,N_9687,N_9633);
or U9929 (N_9929,N_9643,N_9612);
or U9930 (N_9930,N_9689,N_9814);
nand U9931 (N_9931,N_9866,N_9819);
xnor U9932 (N_9932,N_9674,N_9619);
nand U9933 (N_9933,N_9704,N_9624);
nand U9934 (N_9934,N_9695,N_9731);
or U9935 (N_9935,N_9640,N_9810);
and U9936 (N_9936,N_9722,N_9726);
nor U9937 (N_9937,N_9679,N_9724);
xor U9938 (N_9938,N_9636,N_9891);
xor U9939 (N_9939,N_9678,N_9708);
or U9940 (N_9940,N_9683,N_9877);
xnor U9941 (N_9941,N_9743,N_9828);
and U9942 (N_9942,N_9691,N_9763);
xnor U9943 (N_9943,N_9839,N_9651);
xnor U9944 (N_9944,N_9795,N_9699);
or U9945 (N_9945,N_9890,N_9644);
or U9946 (N_9946,N_9853,N_9888);
xnor U9947 (N_9947,N_9613,N_9727);
and U9948 (N_9948,N_9693,N_9802);
and U9949 (N_9949,N_9766,N_9813);
nor U9950 (N_9950,N_9885,N_9849);
xor U9951 (N_9951,N_9785,N_9838);
nor U9952 (N_9952,N_9628,N_9800);
nand U9953 (N_9953,N_9815,N_9641);
nor U9954 (N_9954,N_9701,N_9610);
xnor U9955 (N_9955,N_9601,N_9739);
xnor U9956 (N_9956,N_9720,N_9756);
nand U9957 (N_9957,N_9661,N_9821);
nor U9958 (N_9958,N_9782,N_9835);
and U9959 (N_9959,N_9899,N_9809);
xor U9960 (N_9960,N_9799,N_9875);
nor U9961 (N_9961,N_9616,N_9719);
or U9962 (N_9962,N_9755,N_9778);
or U9963 (N_9963,N_9803,N_9609);
nor U9964 (N_9964,N_9666,N_9735);
nand U9965 (N_9965,N_9844,N_9794);
xor U9966 (N_9966,N_9715,N_9884);
xor U9967 (N_9967,N_9757,N_9713);
nand U9968 (N_9968,N_9869,N_9780);
or U9969 (N_9969,N_9770,N_9622);
and U9970 (N_9970,N_9632,N_9604);
nor U9971 (N_9971,N_9669,N_9837);
nor U9972 (N_9972,N_9623,N_9740);
or U9973 (N_9973,N_9841,N_9617);
xnor U9974 (N_9974,N_9629,N_9816);
and U9975 (N_9975,N_9758,N_9750);
nand U9976 (N_9976,N_9772,N_9897);
xor U9977 (N_9977,N_9650,N_9730);
xor U9978 (N_9978,N_9658,N_9659);
and U9979 (N_9979,N_9747,N_9867);
and U9980 (N_9980,N_9876,N_9664);
or U9981 (N_9981,N_9787,N_9671);
or U9982 (N_9982,N_9752,N_9625);
nand U9983 (N_9983,N_9826,N_9868);
and U9984 (N_9984,N_9860,N_9771);
xor U9985 (N_9985,N_9874,N_9776);
nand U9986 (N_9986,N_9627,N_9685);
nor U9987 (N_9987,N_9754,N_9892);
and U9988 (N_9988,N_9677,N_9748);
nand U9989 (N_9989,N_9728,N_9702);
nand U9990 (N_9990,N_9655,N_9711);
and U9991 (N_9991,N_9709,N_9717);
nand U9992 (N_9992,N_9707,N_9654);
nor U9993 (N_9993,N_9895,N_9865);
xnor U9994 (N_9994,N_9615,N_9789);
xnor U9995 (N_9995,N_9710,N_9642);
or U9996 (N_9996,N_9852,N_9670);
nor U9997 (N_9997,N_9796,N_9652);
nor U9998 (N_9998,N_9706,N_9792);
or U9999 (N_9999,N_9686,N_9716);
or U10000 (N_10000,N_9832,N_9672);
and U10001 (N_10001,N_9760,N_9649);
xor U10002 (N_10002,N_9618,N_9751);
nor U10003 (N_10003,N_9775,N_9630);
xor U10004 (N_10004,N_9893,N_9692);
and U10005 (N_10005,N_9761,N_9737);
or U10006 (N_10006,N_9631,N_9690);
or U10007 (N_10007,N_9746,N_9851);
nand U10008 (N_10008,N_9831,N_9768);
or U10009 (N_10009,N_9834,N_9657);
nor U10010 (N_10010,N_9798,N_9620);
or U10011 (N_10011,N_9824,N_9611);
or U10012 (N_10012,N_9840,N_9606);
nand U10013 (N_10013,N_9898,N_9774);
xor U10014 (N_10014,N_9725,N_9682);
xor U10015 (N_10015,N_9738,N_9602);
nand U10016 (N_10016,N_9697,N_9603);
or U10017 (N_10017,N_9684,N_9859);
xor U10018 (N_10018,N_9648,N_9830);
nor U10019 (N_10019,N_9872,N_9688);
or U10020 (N_10020,N_9783,N_9806);
or U10021 (N_10021,N_9820,N_9608);
xor U10022 (N_10022,N_9788,N_9808);
and U10023 (N_10023,N_9850,N_9881);
and U10024 (N_10024,N_9614,N_9607);
nor U10025 (N_10025,N_9646,N_9676);
nor U10026 (N_10026,N_9805,N_9894);
nor U10027 (N_10027,N_9862,N_9653);
nand U10028 (N_10028,N_9714,N_9873);
xnor U10029 (N_10029,N_9846,N_9817);
and U10030 (N_10030,N_9749,N_9732);
and U10031 (N_10031,N_9764,N_9889);
xnor U10032 (N_10032,N_9887,N_9734);
nor U10033 (N_10033,N_9639,N_9705);
and U10034 (N_10034,N_9721,N_9786);
nor U10035 (N_10035,N_9896,N_9696);
and U10036 (N_10036,N_9797,N_9861);
nand U10037 (N_10037,N_9886,N_9790);
and U10038 (N_10038,N_9662,N_9858);
xor U10039 (N_10039,N_9745,N_9700);
or U10040 (N_10040,N_9781,N_9812);
or U10041 (N_10041,N_9637,N_9847);
xor U10042 (N_10042,N_9681,N_9605);
nor U10043 (N_10043,N_9621,N_9765);
nand U10044 (N_10044,N_9864,N_9718);
xor U10045 (N_10045,N_9634,N_9767);
xnor U10046 (N_10046,N_9836,N_9626);
and U10047 (N_10047,N_9736,N_9827);
nand U10048 (N_10048,N_9703,N_9769);
or U10049 (N_10049,N_9759,N_9822);
nor U10050 (N_10050,N_9760,N_9886);
or U10051 (N_10051,N_9734,N_9767);
nand U10052 (N_10052,N_9867,N_9720);
or U10053 (N_10053,N_9898,N_9884);
or U10054 (N_10054,N_9793,N_9737);
xnor U10055 (N_10055,N_9861,N_9681);
nor U10056 (N_10056,N_9743,N_9633);
and U10057 (N_10057,N_9672,N_9650);
xnor U10058 (N_10058,N_9824,N_9674);
or U10059 (N_10059,N_9816,N_9668);
xor U10060 (N_10060,N_9807,N_9694);
nor U10061 (N_10061,N_9801,N_9824);
and U10062 (N_10062,N_9862,N_9800);
nor U10063 (N_10063,N_9756,N_9626);
nand U10064 (N_10064,N_9875,N_9667);
or U10065 (N_10065,N_9834,N_9669);
nor U10066 (N_10066,N_9614,N_9880);
nand U10067 (N_10067,N_9646,N_9758);
nand U10068 (N_10068,N_9813,N_9698);
and U10069 (N_10069,N_9859,N_9621);
nor U10070 (N_10070,N_9727,N_9861);
nand U10071 (N_10071,N_9824,N_9678);
or U10072 (N_10072,N_9839,N_9790);
and U10073 (N_10073,N_9798,N_9654);
xor U10074 (N_10074,N_9609,N_9797);
and U10075 (N_10075,N_9615,N_9723);
or U10076 (N_10076,N_9868,N_9721);
xnor U10077 (N_10077,N_9685,N_9819);
xnor U10078 (N_10078,N_9813,N_9710);
nand U10079 (N_10079,N_9825,N_9640);
xnor U10080 (N_10080,N_9779,N_9833);
and U10081 (N_10081,N_9662,N_9842);
nand U10082 (N_10082,N_9820,N_9869);
nand U10083 (N_10083,N_9806,N_9856);
or U10084 (N_10084,N_9786,N_9656);
nand U10085 (N_10085,N_9628,N_9651);
and U10086 (N_10086,N_9854,N_9833);
nand U10087 (N_10087,N_9789,N_9663);
nor U10088 (N_10088,N_9734,N_9732);
nor U10089 (N_10089,N_9796,N_9897);
nor U10090 (N_10090,N_9657,N_9776);
nor U10091 (N_10091,N_9638,N_9688);
or U10092 (N_10092,N_9782,N_9831);
nand U10093 (N_10093,N_9681,N_9817);
xor U10094 (N_10094,N_9719,N_9689);
nand U10095 (N_10095,N_9836,N_9677);
nand U10096 (N_10096,N_9813,N_9862);
nand U10097 (N_10097,N_9761,N_9856);
and U10098 (N_10098,N_9877,N_9774);
and U10099 (N_10099,N_9651,N_9846);
nor U10100 (N_10100,N_9767,N_9603);
and U10101 (N_10101,N_9849,N_9718);
nor U10102 (N_10102,N_9755,N_9621);
or U10103 (N_10103,N_9865,N_9788);
nand U10104 (N_10104,N_9898,N_9725);
nor U10105 (N_10105,N_9649,N_9706);
nand U10106 (N_10106,N_9753,N_9603);
xor U10107 (N_10107,N_9846,N_9895);
nand U10108 (N_10108,N_9897,N_9886);
nor U10109 (N_10109,N_9761,N_9615);
nor U10110 (N_10110,N_9770,N_9682);
or U10111 (N_10111,N_9633,N_9648);
and U10112 (N_10112,N_9679,N_9641);
nor U10113 (N_10113,N_9843,N_9835);
and U10114 (N_10114,N_9824,N_9705);
nor U10115 (N_10115,N_9666,N_9749);
or U10116 (N_10116,N_9736,N_9713);
and U10117 (N_10117,N_9658,N_9863);
and U10118 (N_10118,N_9752,N_9772);
nand U10119 (N_10119,N_9645,N_9846);
nor U10120 (N_10120,N_9844,N_9603);
and U10121 (N_10121,N_9640,N_9612);
or U10122 (N_10122,N_9688,N_9601);
or U10123 (N_10123,N_9656,N_9686);
nor U10124 (N_10124,N_9866,N_9737);
nand U10125 (N_10125,N_9746,N_9613);
and U10126 (N_10126,N_9702,N_9805);
and U10127 (N_10127,N_9674,N_9781);
nor U10128 (N_10128,N_9630,N_9856);
nand U10129 (N_10129,N_9826,N_9734);
and U10130 (N_10130,N_9862,N_9661);
and U10131 (N_10131,N_9670,N_9636);
and U10132 (N_10132,N_9841,N_9663);
or U10133 (N_10133,N_9819,N_9710);
or U10134 (N_10134,N_9693,N_9613);
and U10135 (N_10135,N_9730,N_9635);
and U10136 (N_10136,N_9810,N_9633);
and U10137 (N_10137,N_9708,N_9859);
xnor U10138 (N_10138,N_9805,N_9671);
xnor U10139 (N_10139,N_9897,N_9696);
nor U10140 (N_10140,N_9856,N_9752);
and U10141 (N_10141,N_9608,N_9797);
xor U10142 (N_10142,N_9874,N_9698);
xnor U10143 (N_10143,N_9891,N_9621);
and U10144 (N_10144,N_9604,N_9682);
or U10145 (N_10145,N_9837,N_9608);
nand U10146 (N_10146,N_9857,N_9871);
or U10147 (N_10147,N_9788,N_9784);
xnor U10148 (N_10148,N_9638,N_9785);
nor U10149 (N_10149,N_9740,N_9696);
nor U10150 (N_10150,N_9750,N_9640);
and U10151 (N_10151,N_9864,N_9709);
xor U10152 (N_10152,N_9818,N_9787);
nand U10153 (N_10153,N_9850,N_9715);
and U10154 (N_10154,N_9726,N_9873);
or U10155 (N_10155,N_9632,N_9701);
or U10156 (N_10156,N_9705,N_9654);
or U10157 (N_10157,N_9657,N_9771);
nor U10158 (N_10158,N_9652,N_9615);
nor U10159 (N_10159,N_9692,N_9750);
or U10160 (N_10160,N_9827,N_9600);
nor U10161 (N_10161,N_9767,N_9821);
nand U10162 (N_10162,N_9814,N_9729);
xnor U10163 (N_10163,N_9769,N_9750);
and U10164 (N_10164,N_9650,N_9752);
and U10165 (N_10165,N_9795,N_9756);
nand U10166 (N_10166,N_9691,N_9689);
xnor U10167 (N_10167,N_9649,N_9715);
nand U10168 (N_10168,N_9647,N_9608);
nand U10169 (N_10169,N_9653,N_9657);
and U10170 (N_10170,N_9696,N_9892);
nand U10171 (N_10171,N_9742,N_9801);
nor U10172 (N_10172,N_9899,N_9729);
nand U10173 (N_10173,N_9629,N_9688);
and U10174 (N_10174,N_9669,N_9739);
xor U10175 (N_10175,N_9727,N_9796);
and U10176 (N_10176,N_9812,N_9884);
nand U10177 (N_10177,N_9648,N_9707);
xor U10178 (N_10178,N_9682,N_9697);
xnor U10179 (N_10179,N_9674,N_9758);
or U10180 (N_10180,N_9764,N_9683);
and U10181 (N_10181,N_9740,N_9639);
or U10182 (N_10182,N_9648,N_9862);
nor U10183 (N_10183,N_9646,N_9806);
nand U10184 (N_10184,N_9879,N_9800);
or U10185 (N_10185,N_9763,N_9864);
xnor U10186 (N_10186,N_9780,N_9772);
xnor U10187 (N_10187,N_9673,N_9843);
xnor U10188 (N_10188,N_9733,N_9706);
xor U10189 (N_10189,N_9749,N_9777);
or U10190 (N_10190,N_9686,N_9722);
nor U10191 (N_10191,N_9833,N_9639);
xor U10192 (N_10192,N_9855,N_9724);
nor U10193 (N_10193,N_9889,N_9791);
nor U10194 (N_10194,N_9742,N_9681);
nor U10195 (N_10195,N_9868,N_9655);
or U10196 (N_10196,N_9859,N_9834);
nor U10197 (N_10197,N_9883,N_9696);
and U10198 (N_10198,N_9632,N_9877);
and U10199 (N_10199,N_9715,N_9888);
or U10200 (N_10200,N_10067,N_10013);
nor U10201 (N_10201,N_9917,N_10003);
and U10202 (N_10202,N_10001,N_10096);
and U10203 (N_10203,N_9976,N_10161);
xnor U10204 (N_10204,N_10023,N_10092);
nor U10205 (N_10205,N_9914,N_10146);
or U10206 (N_10206,N_9967,N_9935);
nor U10207 (N_10207,N_10139,N_9962);
xnor U10208 (N_10208,N_9980,N_10058);
nand U10209 (N_10209,N_10109,N_10048);
or U10210 (N_10210,N_10129,N_10120);
and U10211 (N_10211,N_9906,N_10021);
or U10212 (N_10212,N_10007,N_10119);
or U10213 (N_10213,N_9989,N_9918);
nand U10214 (N_10214,N_10081,N_9938);
nand U10215 (N_10215,N_10110,N_10085);
or U10216 (N_10216,N_9975,N_10101);
nand U10217 (N_10217,N_10070,N_9940);
and U10218 (N_10218,N_9908,N_10187);
nor U10219 (N_10219,N_9921,N_10106);
nor U10220 (N_10220,N_10133,N_10183);
nand U10221 (N_10221,N_10193,N_10071);
and U10222 (N_10222,N_10136,N_10167);
xnor U10223 (N_10223,N_10004,N_10164);
nor U10224 (N_10224,N_10195,N_9911);
xnor U10225 (N_10225,N_9916,N_10037);
and U10226 (N_10226,N_10141,N_10180);
nand U10227 (N_10227,N_9970,N_9953);
or U10228 (N_10228,N_9946,N_9944);
nor U10229 (N_10229,N_10075,N_10163);
or U10230 (N_10230,N_10131,N_10114);
or U10231 (N_10231,N_10017,N_9960);
xor U10232 (N_10232,N_9900,N_10145);
xor U10233 (N_10233,N_10198,N_9901);
nand U10234 (N_10234,N_9905,N_10154);
and U10235 (N_10235,N_10186,N_9963);
or U10236 (N_10236,N_10086,N_10020);
nor U10237 (N_10237,N_10172,N_9930);
nand U10238 (N_10238,N_9922,N_9902);
nand U10239 (N_10239,N_9997,N_9987);
nand U10240 (N_10240,N_10157,N_10147);
nand U10241 (N_10241,N_9928,N_10043);
and U10242 (N_10242,N_10057,N_10107);
and U10243 (N_10243,N_10000,N_10192);
and U10244 (N_10244,N_10012,N_9981);
xnor U10245 (N_10245,N_10138,N_10051);
nand U10246 (N_10246,N_10045,N_10185);
nand U10247 (N_10247,N_9923,N_9986);
nand U10248 (N_10248,N_9985,N_10103);
xnor U10249 (N_10249,N_9998,N_9925);
nand U10250 (N_10250,N_10165,N_9996);
xnor U10251 (N_10251,N_10079,N_10135);
nor U10252 (N_10252,N_10010,N_10199);
and U10253 (N_10253,N_9974,N_10076);
or U10254 (N_10254,N_10171,N_10052);
xor U10255 (N_10255,N_9973,N_10005);
nor U10256 (N_10256,N_10031,N_10046);
or U10257 (N_10257,N_10044,N_10065);
nand U10258 (N_10258,N_10082,N_9999);
xor U10259 (N_10259,N_10130,N_9927);
nor U10260 (N_10260,N_10009,N_10056);
xnor U10261 (N_10261,N_9942,N_10144);
and U10262 (N_10262,N_10011,N_9959);
and U10263 (N_10263,N_9994,N_9984);
nand U10264 (N_10264,N_10089,N_10176);
and U10265 (N_10265,N_10094,N_10034);
or U10266 (N_10266,N_10059,N_10064);
and U10267 (N_10267,N_10140,N_10162);
nand U10268 (N_10268,N_9948,N_10068);
or U10269 (N_10269,N_9992,N_10159);
and U10270 (N_10270,N_10033,N_10049);
nor U10271 (N_10271,N_10078,N_10022);
and U10272 (N_10272,N_10170,N_9934);
nand U10273 (N_10273,N_9982,N_9958);
xor U10274 (N_10274,N_10190,N_10143);
xor U10275 (N_10275,N_10090,N_10196);
nand U10276 (N_10276,N_9990,N_10156);
and U10277 (N_10277,N_10122,N_9955);
and U10278 (N_10278,N_10024,N_10053);
xor U10279 (N_10279,N_9945,N_9966);
and U10280 (N_10280,N_10108,N_10066);
nor U10281 (N_10281,N_10050,N_9924);
nand U10282 (N_10282,N_9991,N_9941);
xor U10283 (N_10283,N_10168,N_10069);
or U10284 (N_10284,N_9936,N_9913);
xor U10285 (N_10285,N_10173,N_10124);
nor U10286 (N_10286,N_10063,N_10178);
nand U10287 (N_10287,N_10153,N_10137);
nand U10288 (N_10288,N_10041,N_10166);
and U10289 (N_10289,N_9904,N_10029);
and U10290 (N_10290,N_9972,N_9937);
or U10291 (N_10291,N_10019,N_9909);
nor U10292 (N_10292,N_10128,N_10098);
or U10293 (N_10293,N_10188,N_10189);
nand U10294 (N_10294,N_9949,N_9993);
or U10295 (N_10295,N_9933,N_10061);
xor U10296 (N_10296,N_10184,N_9952);
xor U10297 (N_10297,N_10030,N_10142);
or U10298 (N_10298,N_10008,N_9968);
nor U10299 (N_10299,N_10072,N_10006);
and U10300 (N_10300,N_10093,N_10113);
xnor U10301 (N_10301,N_10036,N_10102);
xnor U10302 (N_10302,N_10018,N_10152);
or U10303 (N_10303,N_10027,N_10039);
nor U10304 (N_10304,N_10084,N_10121);
or U10305 (N_10305,N_10123,N_9983);
nor U10306 (N_10306,N_10077,N_10177);
or U10307 (N_10307,N_10194,N_9979);
nor U10308 (N_10308,N_10126,N_10015);
nand U10309 (N_10309,N_9954,N_9964);
nand U10310 (N_10310,N_9920,N_10118);
and U10311 (N_10311,N_9961,N_10055);
nand U10312 (N_10312,N_9965,N_10179);
nor U10313 (N_10313,N_10026,N_10155);
nand U10314 (N_10314,N_9950,N_9956);
and U10315 (N_10315,N_10016,N_10062);
nor U10316 (N_10316,N_9915,N_9903);
or U10317 (N_10317,N_10150,N_10095);
xor U10318 (N_10318,N_10158,N_10083);
nor U10319 (N_10319,N_9969,N_10047);
xor U10320 (N_10320,N_10035,N_9939);
and U10321 (N_10321,N_10073,N_9931);
xor U10322 (N_10322,N_10028,N_10148);
xor U10323 (N_10323,N_10038,N_10032);
xnor U10324 (N_10324,N_9978,N_10025);
nand U10325 (N_10325,N_10100,N_10197);
nand U10326 (N_10326,N_10060,N_10097);
and U10327 (N_10327,N_9951,N_10169);
nor U10328 (N_10328,N_10117,N_9947);
or U10329 (N_10329,N_10002,N_9932);
nor U10330 (N_10330,N_9907,N_10132);
xnor U10331 (N_10331,N_10099,N_9995);
xnor U10332 (N_10332,N_10191,N_10080);
nor U10333 (N_10333,N_10160,N_10111);
nor U10334 (N_10334,N_10042,N_10040);
and U10335 (N_10335,N_10054,N_10014);
and U10336 (N_10336,N_10091,N_10175);
nand U10337 (N_10337,N_10134,N_10125);
or U10338 (N_10338,N_10174,N_9977);
nand U10339 (N_10339,N_9912,N_10181);
nand U10340 (N_10340,N_9929,N_10149);
and U10341 (N_10341,N_9971,N_10087);
and U10342 (N_10342,N_9919,N_10116);
nor U10343 (N_10343,N_10112,N_9943);
xnor U10344 (N_10344,N_10104,N_10088);
nor U10345 (N_10345,N_10151,N_10182);
xnor U10346 (N_10346,N_9957,N_10127);
and U10347 (N_10347,N_10115,N_9988);
or U10348 (N_10348,N_9910,N_10105);
xnor U10349 (N_10349,N_10074,N_9926);
xor U10350 (N_10350,N_10099,N_10187);
nand U10351 (N_10351,N_9925,N_10037);
nand U10352 (N_10352,N_10029,N_10179);
nand U10353 (N_10353,N_9922,N_10155);
and U10354 (N_10354,N_10009,N_9993);
and U10355 (N_10355,N_10025,N_10091);
nand U10356 (N_10356,N_9946,N_10115);
nor U10357 (N_10357,N_9996,N_9933);
nand U10358 (N_10358,N_10024,N_10171);
xnor U10359 (N_10359,N_9990,N_10127);
xnor U10360 (N_10360,N_9906,N_9931);
or U10361 (N_10361,N_10192,N_10177);
and U10362 (N_10362,N_10054,N_10112);
or U10363 (N_10363,N_9947,N_10028);
nand U10364 (N_10364,N_10007,N_10103);
and U10365 (N_10365,N_10146,N_10103);
nor U10366 (N_10366,N_9968,N_10184);
or U10367 (N_10367,N_10191,N_9975);
and U10368 (N_10368,N_10196,N_9942);
or U10369 (N_10369,N_9936,N_9967);
xnor U10370 (N_10370,N_10075,N_9966);
or U10371 (N_10371,N_9936,N_9907);
nor U10372 (N_10372,N_10049,N_10068);
nand U10373 (N_10373,N_10066,N_9965);
nor U10374 (N_10374,N_10150,N_10031);
xnor U10375 (N_10375,N_9960,N_9979);
nor U10376 (N_10376,N_10005,N_10138);
and U10377 (N_10377,N_10100,N_9977);
nor U10378 (N_10378,N_10039,N_10160);
or U10379 (N_10379,N_9958,N_10169);
xnor U10380 (N_10380,N_10014,N_9996);
or U10381 (N_10381,N_9928,N_9909);
xor U10382 (N_10382,N_9940,N_9953);
nor U10383 (N_10383,N_9912,N_10130);
nand U10384 (N_10384,N_10081,N_9901);
xnor U10385 (N_10385,N_9983,N_9900);
xnor U10386 (N_10386,N_10161,N_9964);
nand U10387 (N_10387,N_9911,N_10188);
and U10388 (N_10388,N_9950,N_9992);
xnor U10389 (N_10389,N_9950,N_10050);
or U10390 (N_10390,N_10183,N_10082);
and U10391 (N_10391,N_10182,N_10082);
nand U10392 (N_10392,N_10062,N_9970);
nand U10393 (N_10393,N_10122,N_9908);
nor U10394 (N_10394,N_10082,N_10123);
xor U10395 (N_10395,N_10100,N_10045);
or U10396 (N_10396,N_10023,N_10059);
nand U10397 (N_10397,N_10092,N_10136);
or U10398 (N_10398,N_9968,N_9930);
nand U10399 (N_10399,N_10083,N_10190);
nand U10400 (N_10400,N_10194,N_9920);
and U10401 (N_10401,N_9958,N_10147);
and U10402 (N_10402,N_10085,N_9922);
nand U10403 (N_10403,N_10000,N_10193);
nor U10404 (N_10404,N_9978,N_10199);
nand U10405 (N_10405,N_9929,N_10031);
and U10406 (N_10406,N_10077,N_10091);
nor U10407 (N_10407,N_9993,N_10117);
xnor U10408 (N_10408,N_10177,N_10072);
nor U10409 (N_10409,N_10078,N_9902);
and U10410 (N_10410,N_10064,N_10107);
xor U10411 (N_10411,N_9973,N_10176);
or U10412 (N_10412,N_10116,N_10045);
and U10413 (N_10413,N_10080,N_10078);
or U10414 (N_10414,N_10108,N_9902);
xnor U10415 (N_10415,N_10108,N_10044);
or U10416 (N_10416,N_10012,N_9920);
nand U10417 (N_10417,N_10146,N_10149);
or U10418 (N_10418,N_9907,N_10130);
or U10419 (N_10419,N_10109,N_9913);
or U10420 (N_10420,N_10063,N_10060);
xnor U10421 (N_10421,N_10031,N_10054);
nor U10422 (N_10422,N_10106,N_9923);
or U10423 (N_10423,N_9901,N_9900);
xnor U10424 (N_10424,N_10193,N_10079);
xnor U10425 (N_10425,N_9944,N_10187);
or U10426 (N_10426,N_10115,N_10055);
and U10427 (N_10427,N_10141,N_10027);
and U10428 (N_10428,N_10064,N_9965);
or U10429 (N_10429,N_10027,N_10091);
and U10430 (N_10430,N_10113,N_10031);
and U10431 (N_10431,N_10038,N_10048);
and U10432 (N_10432,N_9930,N_10052);
and U10433 (N_10433,N_9911,N_10168);
and U10434 (N_10434,N_9999,N_9948);
nand U10435 (N_10435,N_9955,N_10096);
xor U10436 (N_10436,N_10111,N_10014);
or U10437 (N_10437,N_10171,N_10180);
nor U10438 (N_10438,N_9955,N_10138);
and U10439 (N_10439,N_10153,N_10182);
xnor U10440 (N_10440,N_9996,N_10052);
nand U10441 (N_10441,N_9921,N_10061);
or U10442 (N_10442,N_9965,N_10069);
xnor U10443 (N_10443,N_10144,N_10095);
nor U10444 (N_10444,N_9908,N_9947);
nand U10445 (N_10445,N_10154,N_10058);
or U10446 (N_10446,N_10085,N_10120);
nand U10447 (N_10447,N_9916,N_9938);
and U10448 (N_10448,N_10165,N_10099);
nor U10449 (N_10449,N_10187,N_10148);
nand U10450 (N_10450,N_9902,N_10080);
or U10451 (N_10451,N_9972,N_10143);
or U10452 (N_10452,N_9950,N_9934);
nor U10453 (N_10453,N_9905,N_10018);
nor U10454 (N_10454,N_10165,N_10039);
nor U10455 (N_10455,N_10041,N_10091);
or U10456 (N_10456,N_10124,N_10073);
nand U10457 (N_10457,N_10058,N_10152);
and U10458 (N_10458,N_9977,N_9913);
nand U10459 (N_10459,N_9903,N_10030);
xor U10460 (N_10460,N_9945,N_10005);
nor U10461 (N_10461,N_9936,N_10025);
and U10462 (N_10462,N_9907,N_10049);
xnor U10463 (N_10463,N_9999,N_9933);
nor U10464 (N_10464,N_9948,N_9990);
or U10465 (N_10465,N_9933,N_9927);
and U10466 (N_10466,N_10125,N_10181);
and U10467 (N_10467,N_10061,N_10026);
nand U10468 (N_10468,N_10181,N_9979);
nor U10469 (N_10469,N_10195,N_10016);
nand U10470 (N_10470,N_10167,N_10050);
xor U10471 (N_10471,N_10132,N_9994);
nor U10472 (N_10472,N_10173,N_10050);
nand U10473 (N_10473,N_10185,N_9983);
nor U10474 (N_10474,N_9986,N_10074);
and U10475 (N_10475,N_10108,N_9981);
or U10476 (N_10476,N_9975,N_10027);
nor U10477 (N_10477,N_9928,N_9952);
or U10478 (N_10478,N_9934,N_10046);
nand U10479 (N_10479,N_9999,N_10088);
nand U10480 (N_10480,N_10023,N_9964);
nor U10481 (N_10481,N_9970,N_10067);
nor U10482 (N_10482,N_10034,N_10138);
and U10483 (N_10483,N_10109,N_10049);
xor U10484 (N_10484,N_10061,N_10088);
and U10485 (N_10485,N_10195,N_9932);
nor U10486 (N_10486,N_10071,N_9935);
nand U10487 (N_10487,N_10194,N_10011);
xnor U10488 (N_10488,N_9924,N_10173);
and U10489 (N_10489,N_10188,N_10030);
and U10490 (N_10490,N_10032,N_9934);
xnor U10491 (N_10491,N_9910,N_10103);
nand U10492 (N_10492,N_9970,N_9990);
and U10493 (N_10493,N_10031,N_10067);
nor U10494 (N_10494,N_10027,N_10083);
and U10495 (N_10495,N_10066,N_10199);
nor U10496 (N_10496,N_10073,N_10050);
and U10497 (N_10497,N_9993,N_10010);
nand U10498 (N_10498,N_10199,N_10079);
or U10499 (N_10499,N_9958,N_10074);
or U10500 (N_10500,N_10248,N_10449);
nand U10501 (N_10501,N_10492,N_10387);
or U10502 (N_10502,N_10208,N_10299);
and U10503 (N_10503,N_10431,N_10301);
xor U10504 (N_10504,N_10309,N_10348);
and U10505 (N_10505,N_10412,N_10496);
xor U10506 (N_10506,N_10298,N_10358);
or U10507 (N_10507,N_10370,N_10371);
nand U10508 (N_10508,N_10398,N_10267);
nor U10509 (N_10509,N_10380,N_10364);
or U10510 (N_10510,N_10469,N_10273);
and U10511 (N_10511,N_10354,N_10243);
or U10512 (N_10512,N_10264,N_10302);
or U10513 (N_10513,N_10305,N_10310);
or U10514 (N_10514,N_10234,N_10219);
nand U10515 (N_10515,N_10488,N_10369);
xor U10516 (N_10516,N_10448,N_10377);
xor U10517 (N_10517,N_10265,N_10434);
nand U10518 (N_10518,N_10419,N_10421);
xnor U10519 (N_10519,N_10294,N_10226);
and U10520 (N_10520,N_10455,N_10222);
xor U10521 (N_10521,N_10470,N_10390);
nand U10522 (N_10522,N_10446,N_10317);
or U10523 (N_10523,N_10463,N_10220);
nor U10524 (N_10524,N_10318,N_10315);
or U10525 (N_10525,N_10335,N_10406);
nand U10526 (N_10526,N_10375,N_10461);
or U10527 (N_10527,N_10439,N_10232);
nor U10528 (N_10528,N_10306,N_10435);
or U10529 (N_10529,N_10295,N_10352);
and U10530 (N_10530,N_10414,N_10473);
xnor U10531 (N_10531,N_10246,N_10253);
and U10532 (N_10532,N_10351,N_10437);
nor U10533 (N_10533,N_10451,N_10224);
or U10534 (N_10534,N_10415,N_10280);
nor U10535 (N_10535,N_10237,N_10472);
nand U10536 (N_10536,N_10320,N_10256);
nor U10537 (N_10537,N_10250,N_10429);
xor U10538 (N_10538,N_10485,N_10445);
and U10539 (N_10539,N_10402,N_10326);
xnor U10540 (N_10540,N_10204,N_10282);
nand U10541 (N_10541,N_10303,N_10279);
xor U10542 (N_10542,N_10423,N_10262);
nor U10543 (N_10543,N_10454,N_10339);
xor U10544 (N_10544,N_10424,N_10286);
nor U10545 (N_10545,N_10458,N_10484);
nand U10546 (N_10546,N_10374,N_10291);
and U10547 (N_10547,N_10331,N_10213);
nor U10548 (N_10548,N_10378,N_10479);
or U10549 (N_10549,N_10201,N_10347);
and U10550 (N_10550,N_10440,N_10361);
nor U10551 (N_10551,N_10413,N_10323);
xnor U10552 (N_10552,N_10225,N_10408);
xnor U10553 (N_10553,N_10202,N_10355);
and U10554 (N_10554,N_10399,N_10211);
or U10555 (N_10555,N_10365,N_10235);
or U10556 (N_10556,N_10283,N_10272);
nor U10557 (N_10557,N_10288,N_10290);
nand U10558 (N_10558,N_10209,N_10251);
and U10559 (N_10559,N_10245,N_10316);
nand U10560 (N_10560,N_10456,N_10478);
xor U10561 (N_10561,N_10254,N_10376);
nor U10562 (N_10562,N_10382,N_10383);
or U10563 (N_10563,N_10452,N_10255);
or U10564 (N_10564,N_10244,N_10236);
nor U10565 (N_10565,N_10268,N_10312);
or U10566 (N_10566,N_10210,N_10327);
xnor U10567 (N_10567,N_10203,N_10436);
nor U10568 (N_10568,N_10462,N_10494);
xor U10569 (N_10569,N_10239,N_10276);
xor U10570 (N_10570,N_10486,N_10442);
nor U10571 (N_10571,N_10223,N_10341);
xnor U10572 (N_10572,N_10395,N_10285);
and U10573 (N_10573,N_10308,N_10403);
nand U10574 (N_10574,N_10433,N_10468);
or U10575 (N_10575,N_10360,N_10405);
and U10576 (N_10576,N_10444,N_10200);
nand U10577 (N_10577,N_10464,N_10495);
nand U10578 (N_10578,N_10293,N_10418);
or U10579 (N_10579,N_10396,N_10259);
nand U10580 (N_10580,N_10384,N_10465);
and U10581 (N_10581,N_10490,N_10428);
or U10582 (N_10582,N_10214,N_10404);
xnor U10583 (N_10583,N_10252,N_10350);
and U10584 (N_10584,N_10389,N_10471);
nor U10585 (N_10585,N_10416,N_10297);
xnor U10586 (N_10586,N_10432,N_10411);
nor U10587 (N_10587,N_10231,N_10319);
nand U10588 (N_10588,N_10271,N_10460);
xnor U10589 (N_10589,N_10438,N_10443);
nand U10590 (N_10590,N_10487,N_10330);
nor U10591 (N_10591,N_10270,N_10205);
xor U10592 (N_10592,N_10221,N_10373);
or U10593 (N_10593,N_10427,N_10356);
xor U10594 (N_10594,N_10275,N_10313);
or U10595 (N_10595,N_10475,N_10314);
or U10596 (N_10596,N_10333,N_10385);
xnor U10597 (N_10597,N_10277,N_10409);
or U10598 (N_10598,N_10338,N_10359);
nand U10599 (N_10599,N_10420,N_10366);
xnor U10600 (N_10600,N_10450,N_10241);
or U10601 (N_10601,N_10362,N_10332);
nand U10602 (N_10602,N_10489,N_10324);
nor U10603 (N_10603,N_10466,N_10346);
nand U10604 (N_10604,N_10284,N_10422);
nand U10605 (N_10605,N_10353,N_10242);
nand U10606 (N_10606,N_10497,N_10388);
nor U10607 (N_10607,N_10228,N_10328);
nand U10608 (N_10608,N_10477,N_10349);
nand U10609 (N_10609,N_10215,N_10278);
nand U10610 (N_10610,N_10474,N_10400);
nor U10611 (N_10611,N_10397,N_10311);
xnor U10612 (N_10612,N_10340,N_10329);
and U10613 (N_10613,N_10266,N_10257);
or U10614 (N_10614,N_10322,N_10357);
or U10615 (N_10615,N_10334,N_10274);
or U10616 (N_10616,N_10263,N_10410);
nand U10617 (N_10617,N_10337,N_10227);
nor U10618 (N_10618,N_10426,N_10281);
xor U10619 (N_10619,N_10481,N_10394);
or U10620 (N_10620,N_10392,N_10206);
nand U10621 (N_10621,N_10480,N_10476);
nor U10622 (N_10622,N_10381,N_10417);
or U10623 (N_10623,N_10482,N_10391);
xnor U10624 (N_10624,N_10336,N_10207);
nor U10625 (N_10625,N_10249,N_10344);
and U10626 (N_10626,N_10240,N_10296);
xnor U10627 (N_10627,N_10321,N_10363);
and U10628 (N_10628,N_10300,N_10407);
and U10629 (N_10629,N_10499,N_10238);
nand U10630 (N_10630,N_10260,N_10325);
nor U10631 (N_10631,N_10393,N_10217);
or U10632 (N_10632,N_10230,N_10483);
nor U10633 (N_10633,N_10368,N_10441);
nor U10634 (N_10634,N_10498,N_10491);
or U10635 (N_10635,N_10216,N_10304);
xnor U10636 (N_10636,N_10379,N_10342);
and U10637 (N_10637,N_10493,N_10425);
nor U10638 (N_10638,N_10258,N_10233);
or U10639 (N_10639,N_10457,N_10261);
nand U10640 (N_10640,N_10247,N_10307);
nor U10641 (N_10641,N_10289,N_10386);
xor U10642 (N_10642,N_10229,N_10372);
and U10643 (N_10643,N_10401,N_10287);
nand U10644 (N_10644,N_10345,N_10218);
and U10645 (N_10645,N_10343,N_10269);
nand U10646 (N_10646,N_10453,N_10367);
nand U10647 (N_10647,N_10467,N_10459);
or U10648 (N_10648,N_10430,N_10292);
nor U10649 (N_10649,N_10447,N_10212);
nand U10650 (N_10650,N_10292,N_10385);
nand U10651 (N_10651,N_10396,N_10392);
or U10652 (N_10652,N_10412,N_10324);
and U10653 (N_10653,N_10321,N_10268);
or U10654 (N_10654,N_10268,N_10208);
nand U10655 (N_10655,N_10379,N_10317);
xor U10656 (N_10656,N_10235,N_10264);
nor U10657 (N_10657,N_10388,N_10429);
nand U10658 (N_10658,N_10223,N_10411);
xnor U10659 (N_10659,N_10336,N_10333);
and U10660 (N_10660,N_10330,N_10477);
or U10661 (N_10661,N_10262,N_10268);
xor U10662 (N_10662,N_10245,N_10265);
nor U10663 (N_10663,N_10331,N_10216);
xnor U10664 (N_10664,N_10363,N_10334);
and U10665 (N_10665,N_10232,N_10474);
xnor U10666 (N_10666,N_10375,N_10414);
nor U10667 (N_10667,N_10410,N_10288);
or U10668 (N_10668,N_10399,N_10421);
nand U10669 (N_10669,N_10369,N_10226);
nand U10670 (N_10670,N_10302,N_10495);
nor U10671 (N_10671,N_10447,N_10268);
xor U10672 (N_10672,N_10263,N_10445);
or U10673 (N_10673,N_10353,N_10264);
or U10674 (N_10674,N_10239,N_10318);
nor U10675 (N_10675,N_10358,N_10339);
and U10676 (N_10676,N_10450,N_10245);
nor U10677 (N_10677,N_10465,N_10247);
or U10678 (N_10678,N_10233,N_10272);
nand U10679 (N_10679,N_10272,N_10243);
nand U10680 (N_10680,N_10469,N_10292);
or U10681 (N_10681,N_10296,N_10416);
or U10682 (N_10682,N_10245,N_10393);
or U10683 (N_10683,N_10409,N_10250);
and U10684 (N_10684,N_10246,N_10291);
nor U10685 (N_10685,N_10335,N_10217);
nor U10686 (N_10686,N_10214,N_10458);
xnor U10687 (N_10687,N_10200,N_10263);
and U10688 (N_10688,N_10362,N_10285);
nand U10689 (N_10689,N_10377,N_10460);
nand U10690 (N_10690,N_10396,N_10443);
or U10691 (N_10691,N_10314,N_10447);
nor U10692 (N_10692,N_10418,N_10272);
xnor U10693 (N_10693,N_10223,N_10380);
nand U10694 (N_10694,N_10200,N_10468);
or U10695 (N_10695,N_10349,N_10297);
nand U10696 (N_10696,N_10432,N_10265);
or U10697 (N_10697,N_10432,N_10434);
or U10698 (N_10698,N_10392,N_10446);
nor U10699 (N_10699,N_10380,N_10409);
and U10700 (N_10700,N_10214,N_10363);
nor U10701 (N_10701,N_10351,N_10209);
nor U10702 (N_10702,N_10296,N_10242);
and U10703 (N_10703,N_10415,N_10393);
or U10704 (N_10704,N_10289,N_10419);
or U10705 (N_10705,N_10309,N_10355);
or U10706 (N_10706,N_10366,N_10253);
nor U10707 (N_10707,N_10382,N_10267);
xnor U10708 (N_10708,N_10336,N_10308);
nor U10709 (N_10709,N_10217,N_10397);
nor U10710 (N_10710,N_10448,N_10402);
nand U10711 (N_10711,N_10215,N_10258);
or U10712 (N_10712,N_10487,N_10320);
xnor U10713 (N_10713,N_10239,N_10278);
nor U10714 (N_10714,N_10316,N_10348);
nand U10715 (N_10715,N_10274,N_10446);
and U10716 (N_10716,N_10381,N_10238);
nor U10717 (N_10717,N_10210,N_10399);
or U10718 (N_10718,N_10259,N_10377);
xnor U10719 (N_10719,N_10459,N_10266);
and U10720 (N_10720,N_10412,N_10241);
xor U10721 (N_10721,N_10361,N_10461);
and U10722 (N_10722,N_10463,N_10208);
and U10723 (N_10723,N_10412,N_10342);
nand U10724 (N_10724,N_10471,N_10255);
xor U10725 (N_10725,N_10341,N_10421);
xnor U10726 (N_10726,N_10312,N_10481);
or U10727 (N_10727,N_10348,N_10499);
or U10728 (N_10728,N_10408,N_10484);
nor U10729 (N_10729,N_10297,N_10282);
xor U10730 (N_10730,N_10376,N_10241);
or U10731 (N_10731,N_10254,N_10240);
or U10732 (N_10732,N_10351,N_10349);
and U10733 (N_10733,N_10200,N_10312);
nor U10734 (N_10734,N_10452,N_10203);
or U10735 (N_10735,N_10473,N_10337);
nor U10736 (N_10736,N_10484,N_10219);
xnor U10737 (N_10737,N_10490,N_10451);
nand U10738 (N_10738,N_10440,N_10370);
xnor U10739 (N_10739,N_10209,N_10457);
and U10740 (N_10740,N_10321,N_10368);
or U10741 (N_10741,N_10390,N_10346);
and U10742 (N_10742,N_10223,N_10267);
and U10743 (N_10743,N_10302,N_10221);
nand U10744 (N_10744,N_10425,N_10395);
or U10745 (N_10745,N_10364,N_10373);
nand U10746 (N_10746,N_10362,N_10284);
and U10747 (N_10747,N_10285,N_10260);
nor U10748 (N_10748,N_10238,N_10235);
nand U10749 (N_10749,N_10213,N_10359);
nand U10750 (N_10750,N_10493,N_10214);
and U10751 (N_10751,N_10384,N_10457);
or U10752 (N_10752,N_10475,N_10212);
and U10753 (N_10753,N_10491,N_10463);
nor U10754 (N_10754,N_10278,N_10380);
nand U10755 (N_10755,N_10361,N_10381);
nand U10756 (N_10756,N_10494,N_10471);
and U10757 (N_10757,N_10243,N_10336);
nand U10758 (N_10758,N_10318,N_10249);
nand U10759 (N_10759,N_10498,N_10461);
and U10760 (N_10760,N_10419,N_10284);
nand U10761 (N_10761,N_10440,N_10241);
nand U10762 (N_10762,N_10304,N_10360);
nand U10763 (N_10763,N_10230,N_10441);
xnor U10764 (N_10764,N_10384,N_10293);
or U10765 (N_10765,N_10232,N_10286);
or U10766 (N_10766,N_10326,N_10285);
and U10767 (N_10767,N_10214,N_10338);
nor U10768 (N_10768,N_10446,N_10305);
and U10769 (N_10769,N_10362,N_10369);
nand U10770 (N_10770,N_10482,N_10348);
xnor U10771 (N_10771,N_10245,N_10209);
and U10772 (N_10772,N_10379,N_10212);
and U10773 (N_10773,N_10404,N_10243);
nor U10774 (N_10774,N_10416,N_10362);
nor U10775 (N_10775,N_10257,N_10472);
nor U10776 (N_10776,N_10318,N_10263);
nor U10777 (N_10777,N_10480,N_10310);
nand U10778 (N_10778,N_10213,N_10391);
or U10779 (N_10779,N_10311,N_10367);
xor U10780 (N_10780,N_10341,N_10275);
xnor U10781 (N_10781,N_10488,N_10498);
xnor U10782 (N_10782,N_10216,N_10448);
nor U10783 (N_10783,N_10209,N_10224);
or U10784 (N_10784,N_10215,N_10201);
or U10785 (N_10785,N_10290,N_10255);
or U10786 (N_10786,N_10421,N_10488);
nor U10787 (N_10787,N_10462,N_10377);
and U10788 (N_10788,N_10257,N_10278);
and U10789 (N_10789,N_10295,N_10414);
xor U10790 (N_10790,N_10317,N_10295);
or U10791 (N_10791,N_10444,N_10255);
nand U10792 (N_10792,N_10228,N_10324);
and U10793 (N_10793,N_10416,N_10338);
nor U10794 (N_10794,N_10343,N_10348);
nand U10795 (N_10795,N_10271,N_10265);
nor U10796 (N_10796,N_10409,N_10473);
nor U10797 (N_10797,N_10332,N_10424);
nor U10798 (N_10798,N_10339,N_10479);
xor U10799 (N_10799,N_10395,N_10259);
nor U10800 (N_10800,N_10694,N_10519);
nor U10801 (N_10801,N_10726,N_10633);
xor U10802 (N_10802,N_10763,N_10594);
or U10803 (N_10803,N_10799,N_10780);
or U10804 (N_10804,N_10585,N_10567);
and U10805 (N_10805,N_10697,N_10739);
xnor U10806 (N_10806,N_10584,N_10632);
nand U10807 (N_10807,N_10647,N_10678);
xor U10808 (N_10808,N_10604,N_10655);
nand U10809 (N_10809,N_10574,N_10589);
xor U10810 (N_10810,N_10675,N_10717);
or U10811 (N_10811,N_10532,N_10564);
nor U10812 (N_10812,N_10586,N_10699);
and U10813 (N_10813,N_10738,N_10745);
or U10814 (N_10814,N_10679,N_10515);
nor U10815 (N_10815,N_10746,N_10751);
or U10816 (N_10816,N_10591,N_10536);
nor U10817 (N_10817,N_10514,N_10702);
or U10818 (N_10818,N_10797,N_10686);
or U10819 (N_10819,N_10565,N_10507);
or U10820 (N_10820,N_10557,N_10768);
xnor U10821 (N_10821,N_10669,N_10545);
nand U10822 (N_10822,N_10628,N_10561);
nor U10823 (N_10823,N_10527,N_10641);
xnor U10824 (N_10824,N_10575,N_10710);
nand U10825 (N_10825,N_10605,N_10523);
nand U10826 (N_10826,N_10755,N_10779);
or U10827 (N_10827,N_10613,N_10725);
and U10828 (N_10828,N_10793,N_10533);
nor U10829 (N_10829,N_10511,N_10764);
or U10830 (N_10830,N_10539,N_10620);
or U10831 (N_10831,N_10707,N_10769);
nand U10832 (N_10832,N_10791,N_10549);
xnor U10833 (N_10833,N_10609,N_10625);
nor U10834 (N_10834,N_10602,N_10503);
nor U10835 (N_10835,N_10508,N_10681);
nand U10836 (N_10836,N_10538,N_10618);
and U10837 (N_10837,N_10524,N_10553);
or U10838 (N_10838,N_10798,N_10658);
nand U10839 (N_10839,N_10588,N_10719);
and U10840 (N_10840,N_10770,N_10667);
and U10841 (N_10841,N_10704,N_10502);
nor U10842 (N_10842,N_10795,N_10547);
or U10843 (N_10843,N_10747,N_10651);
and U10844 (N_10844,N_10551,N_10715);
and U10845 (N_10845,N_10504,N_10711);
nor U10846 (N_10846,N_10505,N_10501);
or U10847 (N_10847,N_10695,N_10785);
or U10848 (N_10848,N_10560,N_10762);
and U10849 (N_10849,N_10736,N_10767);
nor U10850 (N_10850,N_10629,N_10534);
and U10851 (N_10851,N_10643,N_10624);
nand U10852 (N_10852,N_10544,N_10740);
or U10853 (N_10853,N_10787,N_10786);
nand U10854 (N_10854,N_10776,N_10592);
nand U10855 (N_10855,N_10580,N_10646);
or U10856 (N_10856,N_10705,N_10639);
xnor U10857 (N_10857,N_10645,N_10743);
and U10858 (N_10858,N_10610,N_10753);
xor U10859 (N_10859,N_10509,N_10656);
nand U10860 (N_10860,N_10759,N_10765);
or U10861 (N_10861,N_10771,N_10525);
or U10862 (N_10862,N_10714,N_10615);
or U10863 (N_10863,N_10558,N_10706);
nor U10864 (N_10864,N_10723,N_10576);
and U10865 (N_10865,N_10742,N_10626);
xnor U10866 (N_10866,N_10690,N_10607);
and U10867 (N_10867,N_10598,N_10622);
and U10868 (N_10868,N_10573,N_10783);
or U10869 (N_10869,N_10563,N_10623);
or U10870 (N_10870,N_10520,N_10683);
or U10871 (N_10871,N_10708,N_10569);
nand U10872 (N_10872,N_10582,N_10603);
nand U10873 (N_10873,N_10550,N_10506);
or U10874 (N_10874,N_10546,N_10730);
nor U10875 (N_10875,N_10530,N_10516);
xnor U10876 (N_10876,N_10552,N_10542);
or U10877 (N_10877,N_10619,N_10654);
or U10878 (N_10878,N_10721,N_10577);
nand U10879 (N_10879,N_10631,N_10790);
or U10880 (N_10880,N_10616,N_10757);
nor U10881 (N_10881,N_10663,N_10748);
and U10882 (N_10882,N_10665,N_10548);
or U10883 (N_10883,N_10522,N_10664);
xor U10884 (N_10884,N_10526,N_10579);
xor U10885 (N_10885,N_10781,N_10652);
nor U10886 (N_10886,N_10718,N_10649);
and U10887 (N_10887,N_10578,N_10627);
nor U10888 (N_10888,N_10559,N_10720);
nand U10889 (N_10889,N_10572,N_10513);
xnor U10890 (N_10890,N_10693,N_10642);
and U10891 (N_10891,N_10662,N_10630);
nand U10892 (N_10892,N_10556,N_10635);
or U10893 (N_10893,N_10518,N_10703);
and U10894 (N_10894,N_10744,N_10614);
and U10895 (N_10895,N_10670,N_10731);
or U10896 (N_10896,N_10608,N_10775);
nor U10897 (N_10897,N_10660,N_10650);
xor U10898 (N_10898,N_10570,N_10682);
nor U10899 (N_10899,N_10777,N_10644);
xnor U10900 (N_10900,N_10766,N_10612);
nand U10901 (N_10901,N_10684,N_10732);
nand U10902 (N_10902,N_10760,N_10788);
nor U10903 (N_10903,N_10713,N_10648);
nor U10904 (N_10904,N_10774,N_10680);
nor U10905 (N_10905,N_10691,N_10535);
or U10906 (N_10906,N_10555,N_10789);
and U10907 (N_10907,N_10701,N_10674);
nor U10908 (N_10908,N_10709,N_10537);
nor U10909 (N_10909,N_10566,N_10601);
nand U10910 (N_10910,N_10792,N_10571);
xnor U10911 (N_10911,N_10541,N_10758);
or U10912 (N_10912,N_10599,N_10593);
nor U10913 (N_10913,N_10727,N_10510);
nand U10914 (N_10914,N_10722,N_10782);
nor U10915 (N_10915,N_10672,N_10794);
nor U10916 (N_10916,N_10756,N_10712);
and U10917 (N_10917,N_10761,N_10636);
and U10918 (N_10918,N_10671,N_10638);
xnor U10919 (N_10919,N_10597,N_10617);
or U10920 (N_10920,N_10696,N_10688);
nor U10921 (N_10921,N_10554,N_10676);
nand U10922 (N_10922,N_10772,N_10666);
nor U10923 (N_10923,N_10752,N_10583);
nand U10924 (N_10924,N_10621,N_10728);
nor U10925 (N_10925,N_10596,N_10521);
xor U10926 (N_10926,N_10737,N_10653);
and U10927 (N_10927,N_10687,N_10606);
or U10928 (N_10928,N_10528,N_10540);
xor U10929 (N_10929,N_10529,N_10661);
nand U10930 (N_10930,N_10784,N_10600);
and U10931 (N_10931,N_10668,N_10716);
nor U10932 (N_10932,N_10698,N_10724);
nor U10933 (N_10933,N_10673,N_10685);
nor U10934 (N_10934,N_10735,N_10637);
or U10935 (N_10935,N_10640,N_10657);
or U10936 (N_10936,N_10729,N_10517);
xor U10937 (N_10937,N_10500,N_10733);
and U10938 (N_10938,N_10749,N_10754);
nor U10939 (N_10939,N_10692,N_10796);
and U10940 (N_10940,N_10581,N_10562);
nor U10941 (N_10941,N_10659,N_10568);
nor U10942 (N_10942,N_10531,N_10700);
or U10943 (N_10943,N_10634,N_10689);
nand U10944 (N_10944,N_10543,N_10590);
xnor U10945 (N_10945,N_10741,N_10512);
or U10946 (N_10946,N_10773,N_10587);
nand U10947 (N_10947,N_10677,N_10778);
and U10948 (N_10948,N_10595,N_10750);
or U10949 (N_10949,N_10734,N_10611);
nor U10950 (N_10950,N_10510,N_10581);
and U10951 (N_10951,N_10600,N_10766);
and U10952 (N_10952,N_10524,N_10616);
xor U10953 (N_10953,N_10636,N_10677);
nand U10954 (N_10954,N_10758,N_10508);
nand U10955 (N_10955,N_10734,N_10594);
nand U10956 (N_10956,N_10539,N_10635);
and U10957 (N_10957,N_10608,N_10509);
xnor U10958 (N_10958,N_10726,N_10602);
nor U10959 (N_10959,N_10775,N_10719);
xnor U10960 (N_10960,N_10574,N_10500);
or U10961 (N_10961,N_10613,N_10690);
xor U10962 (N_10962,N_10609,N_10525);
nor U10963 (N_10963,N_10739,N_10637);
xor U10964 (N_10964,N_10779,N_10578);
nor U10965 (N_10965,N_10532,N_10596);
xor U10966 (N_10966,N_10572,N_10630);
or U10967 (N_10967,N_10730,N_10647);
or U10968 (N_10968,N_10755,N_10703);
xor U10969 (N_10969,N_10723,N_10529);
nor U10970 (N_10970,N_10551,N_10758);
and U10971 (N_10971,N_10536,N_10566);
xnor U10972 (N_10972,N_10603,N_10722);
xor U10973 (N_10973,N_10516,N_10788);
nand U10974 (N_10974,N_10602,N_10569);
or U10975 (N_10975,N_10536,N_10742);
nand U10976 (N_10976,N_10506,N_10685);
xnor U10977 (N_10977,N_10790,N_10549);
or U10978 (N_10978,N_10672,N_10605);
and U10979 (N_10979,N_10642,N_10729);
nand U10980 (N_10980,N_10757,N_10597);
xor U10981 (N_10981,N_10576,N_10739);
xnor U10982 (N_10982,N_10672,N_10508);
nand U10983 (N_10983,N_10747,N_10734);
nand U10984 (N_10984,N_10674,N_10627);
or U10985 (N_10985,N_10770,N_10590);
nand U10986 (N_10986,N_10618,N_10566);
and U10987 (N_10987,N_10685,N_10703);
nand U10988 (N_10988,N_10529,N_10537);
nor U10989 (N_10989,N_10687,N_10655);
and U10990 (N_10990,N_10589,N_10632);
nand U10991 (N_10991,N_10751,N_10799);
or U10992 (N_10992,N_10653,N_10629);
nand U10993 (N_10993,N_10695,N_10618);
or U10994 (N_10994,N_10534,N_10526);
nand U10995 (N_10995,N_10576,N_10710);
or U10996 (N_10996,N_10608,N_10585);
or U10997 (N_10997,N_10726,N_10667);
or U10998 (N_10998,N_10552,N_10686);
and U10999 (N_10999,N_10615,N_10734);
or U11000 (N_11000,N_10744,N_10787);
nor U11001 (N_11001,N_10688,N_10719);
nand U11002 (N_11002,N_10750,N_10722);
xor U11003 (N_11003,N_10704,N_10695);
and U11004 (N_11004,N_10581,N_10620);
nor U11005 (N_11005,N_10653,N_10695);
or U11006 (N_11006,N_10629,N_10591);
xnor U11007 (N_11007,N_10531,N_10705);
nand U11008 (N_11008,N_10517,N_10671);
nand U11009 (N_11009,N_10687,N_10683);
nor U11010 (N_11010,N_10753,N_10689);
xor U11011 (N_11011,N_10511,N_10660);
and U11012 (N_11012,N_10797,N_10616);
nor U11013 (N_11013,N_10724,N_10599);
nor U11014 (N_11014,N_10607,N_10766);
or U11015 (N_11015,N_10573,N_10530);
nor U11016 (N_11016,N_10637,N_10586);
nor U11017 (N_11017,N_10635,N_10759);
nor U11018 (N_11018,N_10759,N_10723);
xor U11019 (N_11019,N_10683,N_10674);
nor U11020 (N_11020,N_10545,N_10653);
and U11021 (N_11021,N_10570,N_10741);
or U11022 (N_11022,N_10615,N_10569);
nand U11023 (N_11023,N_10543,N_10669);
or U11024 (N_11024,N_10605,N_10622);
and U11025 (N_11025,N_10704,N_10687);
or U11026 (N_11026,N_10546,N_10768);
and U11027 (N_11027,N_10723,N_10510);
or U11028 (N_11028,N_10596,N_10500);
and U11029 (N_11029,N_10537,N_10615);
nor U11030 (N_11030,N_10522,N_10623);
nand U11031 (N_11031,N_10672,N_10676);
or U11032 (N_11032,N_10649,N_10767);
or U11033 (N_11033,N_10698,N_10520);
or U11034 (N_11034,N_10628,N_10668);
xnor U11035 (N_11035,N_10735,N_10726);
and U11036 (N_11036,N_10736,N_10730);
xnor U11037 (N_11037,N_10709,N_10710);
nand U11038 (N_11038,N_10758,N_10546);
nor U11039 (N_11039,N_10611,N_10511);
nand U11040 (N_11040,N_10677,N_10614);
and U11041 (N_11041,N_10649,N_10669);
nand U11042 (N_11042,N_10751,N_10719);
xnor U11043 (N_11043,N_10684,N_10532);
and U11044 (N_11044,N_10519,N_10746);
and U11045 (N_11045,N_10549,N_10616);
xor U11046 (N_11046,N_10736,N_10632);
nor U11047 (N_11047,N_10710,N_10520);
or U11048 (N_11048,N_10769,N_10569);
nand U11049 (N_11049,N_10791,N_10522);
and U11050 (N_11050,N_10628,N_10797);
nor U11051 (N_11051,N_10791,N_10781);
and U11052 (N_11052,N_10554,N_10601);
xnor U11053 (N_11053,N_10519,N_10555);
and U11054 (N_11054,N_10713,N_10628);
nand U11055 (N_11055,N_10583,N_10650);
xnor U11056 (N_11056,N_10614,N_10699);
or U11057 (N_11057,N_10723,N_10592);
nor U11058 (N_11058,N_10740,N_10535);
or U11059 (N_11059,N_10723,N_10689);
and U11060 (N_11060,N_10760,N_10670);
or U11061 (N_11061,N_10770,N_10721);
nor U11062 (N_11062,N_10786,N_10669);
or U11063 (N_11063,N_10733,N_10717);
nor U11064 (N_11064,N_10578,N_10764);
xor U11065 (N_11065,N_10514,N_10789);
nand U11066 (N_11066,N_10765,N_10751);
xnor U11067 (N_11067,N_10765,N_10640);
nand U11068 (N_11068,N_10580,N_10774);
nor U11069 (N_11069,N_10592,N_10598);
xnor U11070 (N_11070,N_10613,N_10534);
or U11071 (N_11071,N_10687,N_10721);
or U11072 (N_11072,N_10504,N_10620);
or U11073 (N_11073,N_10511,N_10567);
xnor U11074 (N_11074,N_10624,N_10693);
xor U11075 (N_11075,N_10690,N_10550);
and U11076 (N_11076,N_10504,N_10761);
nand U11077 (N_11077,N_10783,N_10622);
xnor U11078 (N_11078,N_10511,N_10780);
xor U11079 (N_11079,N_10510,N_10798);
nand U11080 (N_11080,N_10534,N_10543);
nor U11081 (N_11081,N_10654,N_10746);
and U11082 (N_11082,N_10580,N_10695);
nor U11083 (N_11083,N_10685,N_10662);
nand U11084 (N_11084,N_10651,N_10779);
xor U11085 (N_11085,N_10631,N_10637);
xnor U11086 (N_11086,N_10561,N_10622);
and U11087 (N_11087,N_10542,N_10546);
xnor U11088 (N_11088,N_10628,N_10760);
and U11089 (N_11089,N_10556,N_10700);
xnor U11090 (N_11090,N_10575,N_10553);
or U11091 (N_11091,N_10664,N_10688);
nor U11092 (N_11092,N_10686,N_10606);
nand U11093 (N_11093,N_10514,N_10600);
or U11094 (N_11094,N_10505,N_10508);
nor U11095 (N_11095,N_10528,N_10768);
xnor U11096 (N_11096,N_10673,N_10679);
nor U11097 (N_11097,N_10628,N_10655);
xnor U11098 (N_11098,N_10760,N_10752);
nand U11099 (N_11099,N_10504,N_10554);
xnor U11100 (N_11100,N_10950,N_11026);
nand U11101 (N_11101,N_10856,N_10886);
or U11102 (N_11102,N_10922,N_10910);
or U11103 (N_11103,N_10938,N_11039);
xor U11104 (N_11104,N_11006,N_11022);
or U11105 (N_11105,N_11048,N_11001);
or U11106 (N_11106,N_11052,N_10906);
nand U11107 (N_11107,N_11099,N_10872);
or U11108 (N_11108,N_10951,N_11075);
xor U11109 (N_11109,N_11080,N_10835);
nand U11110 (N_11110,N_11072,N_10963);
or U11111 (N_11111,N_10860,N_10810);
and U11112 (N_11112,N_10878,N_11030);
nor U11113 (N_11113,N_10898,N_11057);
xor U11114 (N_11114,N_10865,N_11093);
nor U11115 (N_11115,N_11069,N_10889);
and U11116 (N_11116,N_10894,N_10828);
nand U11117 (N_11117,N_10901,N_11017);
nor U11118 (N_11118,N_11047,N_10831);
nor U11119 (N_11119,N_10907,N_10843);
xnor U11120 (N_11120,N_11061,N_11004);
nor U11121 (N_11121,N_10937,N_10999);
and U11122 (N_11122,N_10837,N_10885);
xor U11123 (N_11123,N_10909,N_11095);
nor U11124 (N_11124,N_11078,N_10957);
nor U11125 (N_11125,N_11009,N_10903);
nor U11126 (N_11126,N_10829,N_11012);
or U11127 (N_11127,N_10945,N_10952);
or U11128 (N_11128,N_10968,N_10832);
and U11129 (N_11129,N_10859,N_11088);
nor U11130 (N_11130,N_10953,N_11033);
and U11131 (N_11131,N_10942,N_10918);
and U11132 (N_11132,N_10845,N_10955);
xor U11133 (N_11133,N_10858,N_11065);
and U11134 (N_11134,N_10993,N_11070);
nand U11135 (N_11135,N_10992,N_11096);
or U11136 (N_11136,N_10987,N_10958);
xnor U11137 (N_11137,N_11021,N_11032);
nor U11138 (N_11138,N_10959,N_11015);
nor U11139 (N_11139,N_10905,N_11034);
nor U11140 (N_11140,N_11092,N_10913);
nand U11141 (N_11141,N_10869,N_10979);
nor U11142 (N_11142,N_10805,N_10853);
nand U11143 (N_11143,N_10931,N_10917);
or U11144 (N_11144,N_11036,N_10804);
xnor U11145 (N_11145,N_10874,N_10912);
or U11146 (N_11146,N_10916,N_10949);
and U11147 (N_11147,N_10815,N_10868);
xnor U11148 (N_11148,N_10940,N_11037);
and U11149 (N_11149,N_11086,N_11005);
or U11150 (N_11150,N_11077,N_10873);
or U11151 (N_11151,N_11087,N_10974);
nor U11152 (N_11152,N_10944,N_11044);
nand U11153 (N_11153,N_10911,N_10883);
or U11154 (N_11154,N_10930,N_11008);
xor U11155 (N_11155,N_11066,N_11079);
and U11156 (N_11156,N_11059,N_11050);
xnor U11157 (N_11157,N_11067,N_11029);
xnor U11158 (N_11158,N_10855,N_10947);
or U11159 (N_11159,N_10862,N_10818);
or U11160 (N_11160,N_10991,N_11028);
xor U11161 (N_11161,N_10854,N_10943);
nor U11162 (N_11162,N_11054,N_10978);
nand U11163 (N_11163,N_10802,N_10971);
nor U11164 (N_11164,N_10961,N_10866);
nand U11165 (N_11165,N_10984,N_10891);
and U11166 (N_11166,N_10813,N_10820);
nand U11167 (N_11167,N_10990,N_11056);
nand U11168 (N_11168,N_10836,N_10882);
and U11169 (N_11169,N_10844,N_10988);
or U11170 (N_11170,N_10871,N_10933);
xor U11171 (N_11171,N_10842,N_10876);
nor U11172 (N_11172,N_10819,N_10877);
xor U11173 (N_11173,N_11000,N_10975);
or U11174 (N_11174,N_10850,N_10928);
or U11175 (N_11175,N_10956,N_11098);
xnor U11176 (N_11176,N_10879,N_10807);
or U11177 (N_11177,N_10921,N_10900);
nor U11178 (N_11178,N_11083,N_10960);
xor U11179 (N_11179,N_11035,N_10896);
nor U11180 (N_11180,N_10801,N_10884);
nand U11181 (N_11181,N_10816,N_10981);
nor U11182 (N_11182,N_10852,N_11081);
and U11183 (N_11183,N_11082,N_10895);
xor U11184 (N_11184,N_10887,N_10899);
nor U11185 (N_11185,N_11042,N_10936);
or U11186 (N_11186,N_11068,N_10998);
nand U11187 (N_11187,N_11063,N_10821);
nor U11188 (N_11188,N_10825,N_11031);
nand U11189 (N_11189,N_10934,N_11002);
nand U11190 (N_11190,N_11014,N_10980);
nor U11191 (N_11191,N_10851,N_10808);
xor U11192 (N_11192,N_11094,N_10983);
or U11193 (N_11193,N_10946,N_10939);
or U11194 (N_11194,N_11010,N_10966);
xor U11195 (N_11195,N_11018,N_10897);
or U11196 (N_11196,N_10809,N_10817);
and U11197 (N_11197,N_11074,N_10997);
xor U11198 (N_11198,N_11053,N_11097);
and U11199 (N_11199,N_11013,N_10830);
nor U11200 (N_11200,N_10919,N_11046);
nor U11201 (N_11201,N_11071,N_10904);
nand U11202 (N_11202,N_10824,N_11016);
or U11203 (N_11203,N_10822,N_10989);
and U11204 (N_11204,N_10941,N_10827);
or U11205 (N_11205,N_10811,N_11089);
nand U11206 (N_11206,N_10970,N_11058);
or U11207 (N_11207,N_11038,N_11040);
nand U11208 (N_11208,N_10929,N_10881);
and U11209 (N_11209,N_11060,N_10995);
nor U11210 (N_11210,N_10838,N_10863);
or U11211 (N_11211,N_10846,N_10977);
xor U11212 (N_11212,N_11003,N_10996);
or U11213 (N_11213,N_11020,N_10926);
nand U11214 (N_11214,N_10880,N_10849);
or U11215 (N_11215,N_11011,N_10840);
or U11216 (N_11216,N_10932,N_10800);
or U11217 (N_11217,N_10834,N_10925);
nor U11218 (N_11218,N_10915,N_11064);
nand U11219 (N_11219,N_10848,N_11024);
and U11220 (N_11220,N_10976,N_10841);
nor U11221 (N_11221,N_10973,N_10833);
and U11222 (N_11222,N_10861,N_10972);
or U11223 (N_11223,N_10964,N_11073);
and U11224 (N_11224,N_10924,N_10920);
nor U11225 (N_11225,N_10948,N_11051);
xor U11226 (N_11226,N_10847,N_10857);
nand U11227 (N_11227,N_10965,N_10982);
nor U11228 (N_11228,N_11023,N_10875);
xor U11229 (N_11229,N_10806,N_11019);
nand U11230 (N_11230,N_10893,N_11041);
or U11231 (N_11231,N_11062,N_10864);
nand U11232 (N_11232,N_10870,N_10986);
nor U11233 (N_11233,N_11043,N_10985);
and U11234 (N_11234,N_10935,N_11084);
and U11235 (N_11235,N_10954,N_10908);
nand U11236 (N_11236,N_10902,N_10888);
and U11237 (N_11237,N_11007,N_11045);
nand U11238 (N_11238,N_10969,N_10814);
xor U11239 (N_11239,N_10867,N_11049);
nor U11240 (N_11240,N_10914,N_10923);
nor U11241 (N_11241,N_10803,N_10839);
xor U11242 (N_11242,N_10994,N_10962);
and U11243 (N_11243,N_10927,N_11076);
or U11244 (N_11244,N_10892,N_11025);
or U11245 (N_11245,N_10890,N_11091);
xnor U11246 (N_11246,N_10826,N_10812);
nor U11247 (N_11247,N_11055,N_11090);
or U11248 (N_11248,N_11085,N_10823);
and U11249 (N_11249,N_11027,N_10967);
or U11250 (N_11250,N_10852,N_10994);
nor U11251 (N_11251,N_10937,N_10942);
xnor U11252 (N_11252,N_10919,N_10992);
xnor U11253 (N_11253,N_10870,N_10913);
nor U11254 (N_11254,N_11019,N_11070);
xor U11255 (N_11255,N_10962,N_11041);
nor U11256 (N_11256,N_10862,N_10999);
xnor U11257 (N_11257,N_11033,N_10931);
xor U11258 (N_11258,N_11037,N_11025);
xnor U11259 (N_11259,N_11016,N_10940);
and U11260 (N_11260,N_11067,N_10964);
or U11261 (N_11261,N_10948,N_10954);
nand U11262 (N_11262,N_10990,N_11062);
xnor U11263 (N_11263,N_10916,N_10971);
nand U11264 (N_11264,N_10856,N_10860);
or U11265 (N_11265,N_11078,N_11059);
xnor U11266 (N_11266,N_11045,N_10973);
and U11267 (N_11267,N_11018,N_10831);
or U11268 (N_11268,N_11091,N_11065);
and U11269 (N_11269,N_11015,N_10800);
nor U11270 (N_11270,N_10848,N_11081);
and U11271 (N_11271,N_11076,N_10900);
nand U11272 (N_11272,N_11092,N_10987);
nand U11273 (N_11273,N_10895,N_11075);
nand U11274 (N_11274,N_10836,N_10941);
xnor U11275 (N_11275,N_10923,N_10839);
and U11276 (N_11276,N_10946,N_11023);
nand U11277 (N_11277,N_11062,N_10950);
or U11278 (N_11278,N_11021,N_11091);
xor U11279 (N_11279,N_10900,N_11032);
and U11280 (N_11280,N_10801,N_10992);
xnor U11281 (N_11281,N_11032,N_11071);
and U11282 (N_11282,N_10893,N_11019);
xnor U11283 (N_11283,N_10982,N_10810);
nand U11284 (N_11284,N_11043,N_11040);
and U11285 (N_11285,N_10940,N_11028);
and U11286 (N_11286,N_11019,N_10857);
or U11287 (N_11287,N_11087,N_10813);
xnor U11288 (N_11288,N_10807,N_11004);
and U11289 (N_11289,N_10859,N_10997);
nand U11290 (N_11290,N_11033,N_10869);
and U11291 (N_11291,N_10800,N_10897);
nand U11292 (N_11292,N_10948,N_11054);
xnor U11293 (N_11293,N_10983,N_10814);
or U11294 (N_11294,N_11042,N_11081);
nand U11295 (N_11295,N_10988,N_11058);
xor U11296 (N_11296,N_10979,N_10829);
nor U11297 (N_11297,N_10922,N_10802);
nor U11298 (N_11298,N_10995,N_10932);
or U11299 (N_11299,N_11025,N_11071);
nand U11300 (N_11300,N_10800,N_10902);
nand U11301 (N_11301,N_10924,N_11082);
and U11302 (N_11302,N_10880,N_11050);
xnor U11303 (N_11303,N_10826,N_10931);
xor U11304 (N_11304,N_10822,N_11085);
or U11305 (N_11305,N_11022,N_11076);
nor U11306 (N_11306,N_10854,N_10993);
nand U11307 (N_11307,N_11065,N_11033);
and U11308 (N_11308,N_11093,N_11073);
and U11309 (N_11309,N_10843,N_11074);
xor U11310 (N_11310,N_11048,N_11029);
and U11311 (N_11311,N_10991,N_11099);
nand U11312 (N_11312,N_10916,N_10965);
nor U11313 (N_11313,N_10854,N_10863);
xnor U11314 (N_11314,N_10974,N_10801);
nand U11315 (N_11315,N_10890,N_11080);
or U11316 (N_11316,N_10836,N_10872);
xnor U11317 (N_11317,N_10856,N_11089);
and U11318 (N_11318,N_11006,N_11093);
and U11319 (N_11319,N_11023,N_10825);
nand U11320 (N_11320,N_10921,N_11032);
xor U11321 (N_11321,N_11012,N_10958);
and U11322 (N_11322,N_10832,N_10866);
and U11323 (N_11323,N_10899,N_11090);
or U11324 (N_11324,N_10802,N_11066);
nor U11325 (N_11325,N_10855,N_10972);
nand U11326 (N_11326,N_10992,N_10817);
or U11327 (N_11327,N_10966,N_11093);
xnor U11328 (N_11328,N_10984,N_10972);
xnor U11329 (N_11329,N_10896,N_10880);
xnor U11330 (N_11330,N_10997,N_10943);
or U11331 (N_11331,N_11086,N_10907);
nand U11332 (N_11332,N_10831,N_10836);
nor U11333 (N_11333,N_10879,N_10835);
nor U11334 (N_11334,N_11014,N_11062);
xnor U11335 (N_11335,N_10891,N_10874);
and U11336 (N_11336,N_11065,N_10966);
nor U11337 (N_11337,N_10806,N_11054);
nand U11338 (N_11338,N_10838,N_11036);
or U11339 (N_11339,N_11068,N_10972);
and U11340 (N_11340,N_10948,N_11000);
or U11341 (N_11341,N_10818,N_10955);
or U11342 (N_11342,N_11046,N_10934);
nand U11343 (N_11343,N_10878,N_10837);
xor U11344 (N_11344,N_10906,N_11005);
or U11345 (N_11345,N_10902,N_11091);
or U11346 (N_11346,N_10878,N_10824);
or U11347 (N_11347,N_11063,N_10842);
nand U11348 (N_11348,N_11044,N_10912);
and U11349 (N_11349,N_11096,N_11049);
or U11350 (N_11350,N_11066,N_11067);
xor U11351 (N_11351,N_10907,N_11037);
nor U11352 (N_11352,N_10989,N_10970);
nor U11353 (N_11353,N_11049,N_10983);
xnor U11354 (N_11354,N_10979,N_11071);
and U11355 (N_11355,N_10893,N_10885);
nor U11356 (N_11356,N_10898,N_11011);
xor U11357 (N_11357,N_10832,N_10954);
nand U11358 (N_11358,N_10939,N_11059);
nor U11359 (N_11359,N_10860,N_11050);
xor U11360 (N_11360,N_10851,N_10887);
and U11361 (N_11361,N_11031,N_10901);
xnor U11362 (N_11362,N_10943,N_11016);
and U11363 (N_11363,N_10921,N_10982);
and U11364 (N_11364,N_10990,N_10834);
xnor U11365 (N_11365,N_10984,N_10918);
xor U11366 (N_11366,N_10868,N_10922);
nand U11367 (N_11367,N_10999,N_10939);
xor U11368 (N_11368,N_11095,N_10916);
or U11369 (N_11369,N_10840,N_10859);
xnor U11370 (N_11370,N_10940,N_11000);
nor U11371 (N_11371,N_10952,N_10922);
and U11372 (N_11372,N_10953,N_11052);
nor U11373 (N_11373,N_10977,N_11043);
and U11374 (N_11374,N_10992,N_10822);
and U11375 (N_11375,N_11015,N_11003);
nor U11376 (N_11376,N_10815,N_11018);
xnor U11377 (N_11377,N_11076,N_11001);
and U11378 (N_11378,N_10829,N_10901);
or U11379 (N_11379,N_11004,N_10886);
nand U11380 (N_11380,N_11084,N_11088);
nor U11381 (N_11381,N_11014,N_11061);
and U11382 (N_11382,N_11081,N_10988);
xnor U11383 (N_11383,N_11012,N_11029);
and U11384 (N_11384,N_11067,N_11092);
or U11385 (N_11385,N_10990,N_10905);
xor U11386 (N_11386,N_11010,N_10909);
and U11387 (N_11387,N_10896,N_10851);
or U11388 (N_11388,N_10932,N_10883);
nor U11389 (N_11389,N_10969,N_10910);
nor U11390 (N_11390,N_11036,N_11017);
or U11391 (N_11391,N_10958,N_10810);
xnor U11392 (N_11392,N_10864,N_10848);
xnor U11393 (N_11393,N_10941,N_10962);
and U11394 (N_11394,N_10905,N_10969);
nor U11395 (N_11395,N_10855,N_10951);
nor U11396 (N_11396,N_11009,N_10945);
or U11397 (N_11397,N_11024,N_10869);
xor U11398 (N_11398,N_11081,N_10822);
nor U11399 (N_11399,N_11017,N_10907);
or U11400 (N_11400,N_11370,N_11273);
nand U11401 (N_11401,N_11238,N_11354);
xnor U11402 (N_11402,N_11169,N_11216);
and U11403 (N_11403,N_11358,N_11153);
or U11404 (N_11404,N_11395,N_11367);
nand U11405 (N_11405,N_11309,N_11340);
and U11406 (N_11406,N_11294,N_11124);
and U11407 (N_11407,N_11311,N_11160);
nand U11408 (N_11408,N_11297,N_11194);
and U11409 (N_11409,N_11338,N_11165);
or U11410 (N_11410,N_11138,N_11135);
and U11411 (N_11411,N_11260,N_11356);
and U11412 (N_11412,N_11334,N_11236);
nand U11413 (N_11413,N_11264,N_11119);
nand U11414 (N_11414,N_11226,N_11346);
or U11415 (N_11415,N_11310,N_11318);
xor U11416 (N_11416,N_11156,N_11145);
and U11417 (N_11417,N_11139,N_11140);
or U11418 (N_11418,N_11333,N_11376);
nor U11419 (N_11419,N_11265,N_11148);
xnor U11420 (N_11420,N_11234,N_11117);
and U11421 (N_11421,N_11157,N_11206);
and U11422 (N_11422,N_11191,N_11313);
and U11423 (N_11423,N_11230,N_11278);
and U11424 (N_11424,N_11232,N_11254);
nor U11425 (N_11425,N_11162,N_11106);
and U11426 (N_11426,N_11239,N_11126);
xor U11427 (N_11427,N_11251,N_11364);
and U11428 (N_11428,N_11352,N_11231);
xor U11429 (N_11429,N_11286,N_11320);
or U11430 (N_11430,N_11287,N_11322);
nand U11431 (N_11431,N_11315,N_11387);
nor U11432 (N_11432,N_11362,N_11131);
and U11433 (N_11433,N_11125,N_11211);
or U11434 (N_11434,N_11281,N_11142);
nand U11435 (N_11435,N_11130,N_11328);
or U11436 (N_11436,N_11290,N_11351);
xor U11437 (N_11437,N_11336,N_11147);
nand U11438 (N_11438,N_11209,N_11144);
and U11439 (N_11439,N_11382,N_11296);
and U11440 (N_11440,N_11366,N_11357);
nor U11441 (N_11441,N_11212,N_11198);
nand U11442 (N_11442,N_11104,N_11196);
nand U11443 (N_11443,N_11255,N_11378);
and U11444 (N_11444,N_11176,N_11240);
xor U11445 (N_11445,N_11244,N_11298);
nor U11446 (N_11446,N_11258,N_11171);
nor U11447 (N_11447,N_11303,N_11306);
nand U11448 (N_11448,N_11183,N_11159);
xor U11449 (N_11449,N_11103,N_11282);
nand U11450 (N_11450,N_11284,N_11396);
or U11451 (N_11451,N_11149,N_11246);
xor U11452 (N_11452,N_11179,N_11245);
nor U11453 (N_11453,N_11204,N_11291);
and U11454 (N_11454,N_11200,N_11243);
xnor U11455 (N_11455,N_11319,N_11329);
and U11456 (N_11456,N_11173,N_11108);
nand U11457 (N_11457,N_11266,N_11220);
or U11458 (N_11458,N_11188,N_11189);
or U11459 (N_11459,N_11347,N_11172);
nor U11460 (N_11460,N_11210,N_11307);
nand U11461 (N_11461,N_11288,N_11348);
nand U11462 (N_11462,N_11305,N_11304);
xnor U11463 (N_11463,N_11228,N_11229);
nand U11464 (N_11464,N_11374,N_11143);
nor U11465 (N_11465,N_11224,N_11375);
nand U11466 (N_11466,N_11280,N_11112);
nand U11467 (N_11467,N_11178,N_11202);
xnor U11468 (N_11468,N_11267,N_11208);
xnor U11469 (N_11469,N_11301,N_11277);
or U11470 (N_11470,N_11353,N_11134);
and U11471 (N_11471,N_11213,N_11377);
xnor U11472 (N_11472,N_11215,N_11343);
or U11473 (N_11473,N_11289,N_11359);
or U11474 (N_11474,N_11295,N_11312);
or U11475 (N_11475,N_11270,N_11355);
xnor U11476 (N_11476,N_11127,N_11170);
xor U11477 (N_11477,N_11337,N_11368);
xor U11478 (N_11478,N_11203,N_11326);
or U11479 (N_11479,N_11107,N_11293);
xor U11480 (N_11480,N_11242,N_11350);
nand U11481 (N_11481,N_11201,N_11256);
and U11482 (N_11482,N_11190,N_11394);
and U11483 (N_11483,N_11187,N_11398);
nand U11484 (N_11484,N_11389,N_11360);
and U11485 (N_11485,N_11122,N_11133);
nor U11486 (N_11486,N_11399,N_11252);
or U11487 (N_11487,N_11365,N_11372);
nand U11488 (N_11488,N_11369,N_11261);
and U11489 (N_11489,N_11101,N_11123);
or U11490 (N_11490,N_11308,N_11175);
xor U11491 (N_11491,N_11113,N_11314);
xor U11492 (N_11492,N_11193,N_11186);
xor U11493 (N_11493,N_11120,N_11109);
xor U11494 (N_11494,N_11332,N_11218);
nor U11495 (N_11495,N_11214,N_11383);
nor U11496 (N_11496,N_11327,N_11259);
nand U11497 (N_11497,N_11146,N_11249);
and U11498 (N_11498,N_11152,N_11136);
nor U11499 (N_11499,N_11250,N_11192);
nor U11500 (N_11500,N_11154,N_11222);
xor U11501 (N_11501,N_11257,N_11339);
nor U11502 (N_11502,N_11317,N_11237);
or U11503 (N_11503,N_11115,N_11241);
or U11504 (N_11504,N_11151,N_11393);
or U11505 (N_11505,N_11342,N_11180);
or U11506 (N_11506,N_11129,N_11235);
xor U11507 (N_11507,N_11274,N_11150);
or U11508 (N_11508,N_11379,N_11279);
nand U11509 (N_11509,N_11302,N_11330);
xor U11510 (N_11510,N_11102,N_11184);
nor U11511 (N_11511,N_11269,N_11205);
and U11512 (N_11512,N_11321,N_11181);
nand U11513 (N_11513,N_11141,N_11248);
and U11514 (N_11514,N_11373,N_11324);
nor U11515 (N_11515,N_11361,N_11137);
or U11516 (N_11516,N_11391,N_11118);
or U11517 (N_11517,N_11253,N_11199);
xnor U11518 (N_11518,N_11397,N_11167);
or U11519 (N_11519,N_11110,N_11363);
or U11520 (N_11520,N_11223,N_11177);
nor U11521 (N_11521,N_11388,N_11331);
nand U11522 (N_11522,N_11105,N_11285);
or U11523 (N_11523,N_11132,N_11316);
xor U11524 (N_11524,N_11128,N_11349);
and U11525 (N_11525,N_11219,N_11275);
nor U11526 (N_11526,N_11168,N_11161);
and U11527 (N_11527,N_11185,N_11174);
nor U11528 (N_11528,N_11335,N_11381);
nand U11529 (N_11529,N_11392,N_11233);
nand U11530 (N_11530,N_11325,N_11371);
or U11531 (N_11531,N_11345,N_11268);
or U11532 (N_11532,N_11221,N_11386);
or U11533 (N_11533,N_11380,N_11344);
xnor U11534 (N_11534,N_11163,N_11271);
nor U11535 (N_11535,N_11195,N_11111);
xnor U11536 (N_11536,N_11217,N_11158);
xnor U11537 (N_11537,N_11225,N_11155);
nor U11538 (N_11538,N_11164,N_11227);
and U11539 (N_11539,N_11247,N_11207);
nor U11540 (N_11540,N_11182,N_11116);
nand U11541 (N_11541,N_11292,N_11197);
and U11542 (N_11542,N_11385,N_11384);
nand U11543 (N_11543,N_11300,N_11114);
or U11544 (N_11544,N_11323,N_11263);
and U11545 (N_11545,N_11100,N_11262);
or U11546 (N_11546,N_11299,N_11272);
nor U11547 (N_11547,N_11121,N_11166);
xnor U11548 (N_11548,N_11276,N_11283);
xnor U11549 (N_11549,N_11341,N_11390);
nor U11550 (N_11550,N_11254,N_11306);
or U11551 (N_11551,N_11337,N_11371);
nand U11552 (N_11552,N_11109,N_11122);
nor U11553 (N_11553,N_11188,N_11387);
nand U11554 (N_11554,N_11381,N_11366);
and U11555 (N_11555,N_11368,N_11143);
xnor U11556 (N_11556,N_11241,N_11315);
or U11557 (N_11557,N_11128,N_11204);
or U11558 (N_11558,N_11332,N_11394);
xor U11559 (N_11559,N_11126,N_11330);
and U11560 (N_11560,N_11297,N_11373);
nor U11561 (N_11561,N_11326,N_11256);
xnor U11562 (N_11562,N_11235,N_11393);
or U11563 (N_11563,N_11144,N_11355);
nor U11564 (N_11564,N_11371,N_11230);
and U11565 (N_11565,N_11100,N_11298);
or U11566 (N_11566,N_11304,N_11321);
xnor U11567 (N_11567,N_11382,N_11234);
xnor U11568 (N_11568,N_11270,N_11202);
and U11569 (N_11569,N_11180,N_11204);
xor U11570 (N_11570,N_11121,N_11388);
xnor U11571 (N_11571,N_11250,N_11198);
or U11572 (N_11572,N_11100,N_11101);
nand U11573 (N_11573,N_11327,N_11190);
or U11574 (N_11574,N_11108,N_11152);
nor U11575 (N_11575,N_11110,N_11204);
and U11576 (N_11576,N_11330,N_11296);
and U11577 (N_11577,N_11284,N_11115);
or U11578 (N_11578,N_11253,N_11135);
or U11579 (N_11579,N_11220,N_11200);
or U11580 (N_11580,N_11257,N_11199);
and U11581 (N_11581,N_11161,N_11239);
xor U11582 (N_11582,N_11352,N_11203);
or U11583 (N_11583,N_11102,N_11328);
or U11584 (N_11584,N_11305,N_11242);
xnor U11585 (N_11585,N_11221,N_11399);
xor U11586 (N_11586,N_11311,N_11363);
nand U11587 (N_11587,N_11334,N_11231);
or U11588 (N_11588,N_11333,N_11291);
or U11589 (N_11589,N_11147,N_11219);
and U11590 (N_11590,N_11228,N_11353);
and U11591 (N_11591,N_11259,N_11203);
nor U11592 (N_11592,N_11357,N_11337);
xnor U11593 (N_11593,N_11335,N_11236);
xnor U11594 (N_11594,N_11119,N_11248);
or U11595 (N_11595,N_11368,N_11113);
nor U11596 (N_11596,N_11250,N_11178);
xnor U11597 (N_11597,N_11118,N_11121);
or U11598 (N_11598,N_11377,N_11130);
or U11599 (N_11599,N_11389,N_11190);
xnor U11600 (N_11600,N_11108,N_11343);
and U11601 (N_11601,N_11221,N_11179);
or U11602 (N_11602,N_11286,N_11265);
nor U11603 (N_11603,N_11284,N_11229);
xor U11604 (N_11604,N_11200,N_11269);
nor U11605 (N_11605,N_11335,N_11162);
and U11606 (N_11606,N_11387,N_11141);
nand U11607 (N_11607,N_11197,N_11181);
xnor U11608 (N_11608,N_11350,N_11315);
nor U11609 (N_11609,N_11297,N_11121);
and U11610 (N_11610,N_11242,N_11325);
or U11611 (N_11611,N_11251,N_11222);
nor U11612 (N_11612,N_11311,N_11102);
or U11613 (N_11613,N_11374,N_11286);
or U11614 (N_11614,N_11272,N_11263);
and U11615 (N_11615,N_11227,N_11372);
and U11616 (N_11616,N_11278,N_11363);
xor U11617 (N_11617,N_11368,N_11173);
nor U11618 (N_11618,N_11126,N_11289);
nand U11619 (N_11619,N_11292,N_11142);
nand U11620 (N_11620,N_11287,N_11204);
or U11621 (N_11621,N_11270,N_11229);
xor U11622 (N_11622,N_11112,N_11293);
or U11623 (N_11623,N_11254,N_11312);
xor U11624 (N_11624,N_11376,N_11211);
nand U11625 (N_11625,N_11355,N_11302);
nor U11626 (N_11626,N_11246,N_11218);
or U11627 (N_11627,N_11348,N_11253);
or U11628 (N_11628,N_11148,N_11392);
nor U11629 (N_11629,N_11162,N_11122);
and U11630 (N_11630,N_11362,N_11267);
and U11631 (N_11631,N_11287,N_11142);
xor U11632 (N_11632,N_11342,N_11328);
xnor U11633 (N_11633,N_11198,N_11306);
xnor U11634 (N_11634,N_11321,N_11160);
and U11635 (N_11635,N_11245,N_11206);
xnor U11636 (N_11636,N_11300,N_11161);
xor U11637 (N_11637,N_11210,N_11245);
nand U11638 (N_11638,N_11354,N_11291);
nor U11639 (N_11639,N_11305,N_11349);
nand U11640 (N_11640,N_11165,N_11190);
and U11641 (N_11641,N_11181,N_11223);
and U11642 (N_11642,N_11105,N_11164);
and U11643 (N_11643,N_11281,N_11129);
nor U11644 (N_11644,N_11327,N_11197);
and U11645 (N_11645,N_11261,N_11383);
xor U11646 (N_11646,N_11174,N_11221);
xnor U11647 (N_11647,N_11289,N_11387);
nand U11648 (N_11648,N_11339,N_11172);
and U11649 (N_11649,N_11349,N_11172);
and U11650 (N_11650,N_11128,N_11187);
or U11651 (N_11651,N_11139,N_11284);
xnor U11652 (N_11652,N_11338,N_11125);
and U11653 (N_11653,N_11134,N_11171);
and U11654 (N_11654,N_11245,N_11273);
xnor U11655 (N_11655,N_11379,N_11370);
nand U11656 (N_11656,N_11168,N_11276);
nand U11657 (N_11657,N_11175,N_11138);
and U11658 (N_11658,N_11215,N_11322);
nand U11659 (N_11659,N_11347,N_11379);
nor U11660 (N_11660,N_11151,N_11252);
or U11661 (N_11661,N_11373,N_11166);
nand U11662 (N_11662,N_11226,N_11191);
nor U11663 (N_11663,N_11372,N_11349);
nor U11664 (N_11664,N_11282,N_11391);
xnor U11665 (N_11665,N_11337,N_11249);
xor U11666 (N_11666,N_11111,N_11334);
nand U11667 (N_11667,N_11103,N_11126);
nand U11668 (N_11668,N_11346,N_11156);
or U11669 (N_11669,N_11307,N_11300);
and U11670 (N_11670,N_11259,N_11381);
xnor U11671 (N_11671,N_11388,N_11294);
nor U11672 (N_11672,N_11163,N_11329);
nand U11673 (N_11673,N_11338,N_11367);
and U11674 (N_11674,N_11266,N_11294);
and U11675 (N_11675,N_11327,N_11230);
xnor U11676 (N_11676,N_11290,N_11122);
nand U11677 (N_11677,N_11247,N_11137);
or U11678 (N_11678,N_11109,N_11373);
nand U11679 (N_11679,N_11232,N_11184);
nand U11680 (N_11680,N_11399,N_11384);
nor U11681 (N_11681,N_11220,N_11379);
and U11682 (N_11682,N_11172,N_11289);
or U11683 (N_11683,N_11155,N_11141);
nand U11684 (N_11684,N_11340,N_11314);
nor U11685 (N_11685,N_11341,N_11225);
nand U11686 (N_11686,N_11317,N_11113);
nor U11687 (N_11687,N_11385,N_11193);
and U11688 (N_11688,N_11384,N_11243);
and U11689 (N_11689,N_11141,N_11319);
xnor U11690 (N_11690,N_11135,N_11203);
or U11691 (N_11691,N_11224,N_11344);
nand U11692 (N_11692,N_11276,N_11317);
xnor U11693 (N_11693,N_11121,N_11190);
or U11694 (N_11694,N_11389,N_11383);
xnor U11695 (N_11695,N_11249,N_11140);
or U11696 (N_11696,N_11135,N_11181);
nand U11697 (N_11697,N_11369,N_11131);
nand U11698 (N_11698,N_11205,N_11159);
xor U11699 (N_11699,N_11386,N_11158);
or U11700 (N_11700,N_11606,N_11504);
nor U11701 (N_11701,N_11605,N_11632);
and U11702 (N_11702,N_11691,N_11547);
and U11703 (N_11703,N_11469,N_11499);
xor U11704 (N_11704,N_11566,N_11636);
nand U11705 (N_11705,N_11588,N_11450);
xor U11706 (N_11706,N_11608,N_11492);
nand U11707 (N_11707,N_11640,N_11459);
or U11708 (N_11708,N_11674,N_11622);
or U11709 (N_11709,N_11637,N_11573);
nor U11710 (N_11710,N_11522,N_11653);
xnor U11711 (N_11711,N_11457,N_11501);
nor U11712 (N_11712,N_11631,N_11663);
and U11713 (N_11713,N_11496,N_11462);
or U11714 (N_11714,N_11687,N_11667);
and U11715 (N_11715,N_11480,N_11426);
and U11716 (N_11716,N_11555,N_11515);
xnor U11717 (N_11717,N_11562,N_11530);
nor U11718 (N_11718,N_11455,N_11671);
and U11719 (N_11719,N_11623,N_11537);
nor U11720 (N_11720,N_11543,N_11624);
and U11721 (N_11721,N_11656,N_11603);
xnor U11722 (N_11722,N_11581,N_11604);
or U11723 (N_11723,N_11595,N_11629);
and U11724 (N_11724,N_11690,N_11675);
nor U11725 (N_11725,N_11415,N_11633);
nor U11726 (N_11726,N_11490,N_11488);
nand U11727 (N_11727,N_11615,N_11402);
or U11728 (N_11728,N_11585,N_11645);
nor U11729 (N_11729,N_11693,N_11472);
or U11730 (N_11730,N_11429,N_11500);
and U11731 (N_11731,N_11525,N_11463);
nor U11732 (N_11732,N_11494,N_11614);
nand U11733 (N_11733,N_11422,N_11590);
nor U11734 (N_11734,N_11541,N_11613);
and U11735 (N_11735,N_11669,N_11695);
xor U11736 (N_11736,N_11424,N_11616);
and U11737 (N_11737,N_11578,N_11418);
or U11738 (N_11738,N_11523,N_11567);
xor U11739 (N_11739,N_11602,N_11458);
and U11740 (N_11740,N_11516,N_11617);
xnor U11741 (N_11741,N_11404,N_11688);
and U11742 (N_11742,N_11546,N_11431);
nand U11743 (N_11743,N_11611,N_11412);
nand U11744 (N_11744,N_11460,N_11527);
or U11745 (N_11745,N_11420,N_11502);
and U11746 (N_11746,N_11630,N_11526);
nand U11747 (N_11747,N_11445,N_11430);
and U11748 (N_11748,N_11452,N_11580);
and U11749 (N_11749,N_11503,N_11564);
or U11750 (N_11750,N_11427,N_11493);
and U11751 (N_11751,N_11621,N_11444);
and U11752 (N_11752,N_11536,N_11448);
or U11753 (N_11753,N_11405,N_11654);
nor U11754 (N_11754,N_11435,N_11419);
nand U11755 (N_11755,N_11644,N_11540);
nor U11756 (N_11756,N_11681,N_11533);
nand U11757 (N_11757,N_11416,N_11495);
and U11758 (N_11758,N_11483,N_11627);
or U11759 (N_11759,N_11507,N_11454);
or U11760 (N_11760,N_11571,N_11679);
nand U11761 (N_11761,N_11570,N_11549);
nand U11762 (N_11762,N_11465,N_11620);
and U11763 (N_11763,N_11414,N_11572);
nor U11764 (N_11764,N_11409,N_11598);
xnor U11765 (N_11765,N_11521,N_11650);
nand U11766 (N_11766,N_11639,N_11408);
or U11767 (N_11767,N_11531,N_11596);
nand U11768 (N_11768,N_11664,N_11489);
or U11769 (N_11769,N_11649,N_11635);
nor U11770 (N_11770,N_11586,N_11642);
nand U11771 (N_11771,N_11619,N_11625);
xor U11772 (N_11772,N_11478,N_11474);
xor U11773 (N_11773,N_11591,N_11468);
or U11774 (N_11774,N_11432,N_11610);
xnor U11775 (N_11775,N_11689,N_11439);
or U11776 (N_11776,N_11456,N_11648);
nand U11777 (N_11777,N_11647,N_11660);
nand U11778 (N_11778,N_11423,N_11400);
nand U11779 (N_11779,N_11498,N_11612);
nand U11780 (N_11780,N_11421,N_11593);
or U11781 (N_11781,N_11662,N_11582);
and U11782 (N_11782,N_11532,N_11659);
nor U11783 (N_11783,N_11479,N_11668);
nand U11784 (N_11784,N_11511,N_11512);
and U11785 (N_11785,N_11554,N_11491);
and U11786 (N_11786,N_11584,N_11477);
or U11787 (N_11787,N_11678,N_11634);
or U11788 (N_11788,N_11411,N_11673);
and U11789 (N_11789,N_11410,N_11481);
xor U11790 (N_11790,N_11524,N_11626);
xor U11791 (N_11791,N_11529,N_11406);
nand U11792 (N_11792,N_11535,N_11594);
or U11793 (N_11793,N_11552,N_11550);
xor U11794 (N_11794,N_11484,N_11470);
xor U11795 (N_11795,N_11651,N_11449);
xnor U11796 (N_11796,N_11561,N_11607);
or U11797 (N_11797,N_11519,N_11518);
nor U11798 (N_11798,N_11506,N_11609);
or U11799 (N_11799,N_11425,N_11497);
xnor U11800 (N_11800,N_11438,N_11646);
nand U11801 (N_11801,N_11677,N_11553);
nor U11802 (N_11802,N_11583,N_11509);
nor U11803 (N_11803,N_11413,N_11436);
or U11804 (N_11804,N_11514,N_11403);
and U11805 (N_11805,N_11539,N_11579);
and U11806 (N_11806,N_11447,N_11538);
or U11807 (N_11807,N_11434,N_11428);
xnor U11808 (N_11808,N_11560,N_11505);
or U11809 (N_11809,N_11587,N_11464);
xnor U11810 (N_11810,N_11685,N_11682);
nand U11811 (N_11811,N_11569,N_11551);
nand U11812 (N_11812,N_11655,N_11442);
nor U11813 (N_11813,N_11513,N_11577);
nand U11814 (N_11814,N_11597,N_11565);
xor U11815 (N_11815,N_11510,N_11600);
nand U11816 (N_11816,N_11574,N_11433);
or U11817 (N_11817,N_11544,N_11443);
xor U11818 (N_11818,N_11699,N_11661);
and U11819 (N_11819,N_11558,N_11446);
nor U11820 (N_11820,N_11638,N_11601);
or U11821 (N_11821,N_11401,N_11618);
nor U11822 (N_11822,N_11476,N_11697);
xnor U11823 (N_11823,N_11520,N_11592);
nor U11824 (N_11824,N_11696,N_11508);
nor U11825 (N_11825,N_11684,N_11517);
xnor U11826 (N_11826,N_11575,N_11576);
nand U11827 (N_11827,N_11665,N_11440);
and U11828 (N_11828,N_11482,N_11643);
or U11829 (N_11829,N_11467,N_11485);
or U11830 (N_11830,N_11487,N_11694);
nand U11831 (N_11831,N_11473,N_11676);
or U11832 (N_11832,N_11563,N_11568);
and U11833 (N_11833,N_11658,N_11486);
and U11834 (N_11834,N_11641,N_11441);
nor U11835 (N_11835,N_11692,N_11672);
nor U11836 (N_11836,N_11417,N_11534);
and U11837 (N_11837,N_11698,N_11407);
nor U11838 (N_11838,N_11451,N_11686);
nor U11839 (N_11839,N_11548,N_11542);
nor U11840 (N_11840,N_11475,N_11466);
xnor U11841 (N_11841,N_11599,N_11559);
or U11842 (N_11842,N_11670,N_11556);
and U11843 (N_11843,N_11557,N_11652);
nor U11844 (N_11844,N_11589,N_11471);
and U11845 (N_11845,N_11683,N_11453);
xor U11846 (N_11846,N_11680,N_11628);
nand U11847 (N_11847,N_11437,N_11657);
nand U11848 (N_11848,N_11528,N_11461);
and U11849 (N_11849,N_11545,N_11666);
nand U11850 (N_11850,N_11662,N_11606);
xnor U11851 (N_11851,N_11601,N_11470);
and U11852 (N_11852,N_11545,N_11489);
nor U11853 (N_11853,N_11457,N_11579);
nand U11854 (N_11854,N_11467,N_11443);
nand U11855 (N_11855,N_11490,N_11435);
nor U11856 (N_11856,N_11560,N_11646);
or U11857 (N_11857,N_11474,N_11573);
and U11858 (N_11858,N_11667,N_11592);
or U11859 (N_11859,N_11693,N_11654);
and U11860 (N_11860,N_11446,N_11419);
xnor U11861 (N_11861,N_11414,N_11654);
or U11862 (N_11862,N_11651,N_11558);
or U11863 (N_11863,N_11629,N_11414);
xnor U11864 (N_11864,N_11559,N_11523);
nor U11865 (N_11865,N_11633,N_11491);
and U11866 (N_11866,N_11632,N_11535);
nor U11867 (N_11867,N_11563,N_11668);
xnor U11868 (N_11868,N_11587,N_11582);
or U11869 (N_11869,N_11616,N_11578);
nor U11870 (N_11870,N_11470,N_11486);
and U11871 (N_11871,N_11512,N_11667);
nor U11872 (N_11872,N_11431,N_11575);
nand U11873 (N_11873,N_11541,N_11699);
and U11874 (N_11874,N_11608,N_11511);
and U11875 (N_11875,N_11534,N_11408);
xnor U11876 (N_11876,N_11656,N_11663);
xnor U11877 (N_11877,N_11503,N_11675);
xnor U11878 (N_11878,N_11475,N_11512);
xor U11879 (N_11879,N_11621,N_11527);
nand U11880 (N_11880,N_11506,N_11457);
and U11881 (N_11881,N_11690,N_11660);
or U11882 (N_11882,N_11676,N_11457);
nor U11883 (N_11883,N_11690,N_11438);
nand U11884 (N_11884,N_11671,N_11524);
nand U11885 (N_11885,N_11696,N_11556);
or U11886 (N_11886,N_11615,N_11595);
nand U11887 (N_11887,N_11631,N_11433);
xnor U11888 (N_11888,N_11633,N_11596);
xnor U11889 (N_11889,N_11655,N_11696);
or U11890 (N_11890,N_11461,N_11531);
or U11891 (N_11891,N_11412,N_11683);
or U11892 (N_11892,N_11423,N_11476);
nor U11893 (N_11893,N_11574,N_11558);
or U11894 (N_11894,N_11500,N_11640);
or U11895 (N_11895,N_11549,N_11686);
or U11896 (N_11896,N_11486,N_11497);
xnor U11897 (N_11897,N_11603,N_11619);
nor U11898 (N_11898,N_11594,N_11489);
nand U11899 (N_11899,N_11418,N_11638);
and U11900 (N_11900,N_11406,N_11621);
and U11901 (N_11901,N_11573,N_11601);
or U11902 (N_11902,N_11594,N_11674);
and U11903 (N_11903,N_11485,N_11620);
and U11904 (N_11904,N_11414,N_11689);
nand U11905 (N_11905,N_11543,N_11550);
xnor U11906 (N_11906,N_11434,N_11657);
or U11907 (N_11907,N_11602,N_11684);
and U11908 (N_11908,N_11640,N_11414);
nor U11909 (N_11909,N_11623,N_11472);
nand U11910 (N_11910,N_11512,N_11605);
xor U11911 (N_11911,N_11481,N_11446);
or U11912 (N_11912,N_11683,N_11602);
nand U11913 (N_11913,N_11443,N_11608);
and U11914 (N_11914,N_11538,N_11416);
or U11915 (N_11915,N_11610,N_11590);
and U11916 (N_11916,N_11507,N_11668);
xor U11917 (N_11917,N_11697,N_11699);
nor U11918 (N_11918,N_11443,N_11691);
nor U11919 (N_11919,N_11422,N_11439);
nor U11920 (N_11920,N_11471,N_11461);
xor U11921 (N_11921,N_11448,N_11580);
nor U11922 (N_11922,N_11576,N_11418);
nor U11923 (N_11923,N_11672,N_11600);
or U11924 (N_11924,N_11659,N_11488);
xnor U11925 (N_11925,N_11585,N_11559);
nor U11926 (N_11926,N_11431,N_11665);
and U11927 (N_11927,N_11536,N_11575);
and U11928 (N_11928,N_11689,N_11549);
nor U11929 (N_11929,N_11489,N_11618);
or U11930 (N_11930,N_11418,N_11407);
nand U11931 (N_11931,N_11679,N_11463);
and U11932 (N_11932,N_11584,N_11551);
nor U11933 (N_11933,N_11642,N_11501);
and U11934 (N_11934,N_11573,N_11627);
xor U11935 (N_11935,N_11591,N_11697);
or U11936 (N_11936,N_11510,N_11466);
nand U11937 (N_11937,N_11603,N_11582);
and U11938 (N_11938,N_11482,N_11488);
xnor U11939 (N_11939,N_11638,N_11560);
nor U11940 (N_11940,N_11459,N_11601);
and U11941 (N_11941,N_11477,N_11452);
or U11942 (N_11942,N_11662,N_11505);
and U11943 (N_11943,N_11627,N_11509);
nor U11944 (N_11944,N_11627,N_11557);
xor U11945 (N_11945,N_11609,N_11479);
and U11946 (N_11946,N_11556,N_11562);
xor U11947 (N_11947,N_11542,N_11653);
xnor U11948 (N_11948,N_11601,N_11541);
and U11949 (N_11949,N_11685,N_11649);
and U11950 (N_11950,N_11581,N_11626);
nor U11951 (N_11951,N_11514,N_11593);
or U11952 (N_11952,N_11670,N_11437);
nor U11953 (N_11953,N_11590,N_11476);
and U11954 (N_11954,N_11423,N_11553);
and U11955 (N_11955,N_11636,N_11632);
and U11956 (N_11956,N_11410,N_11672);
nand U11957 (N_11957,N_11536,N_11522);
nand U11958 (N_11958,N_11622,N_11599);
nand U11959 (N_11959,N_11584,N_11571);
or U11960 (N_11960,N_11623,N_11670);
xor U11961 (N_11961,N_11409,N_11676);
nor U11962 (N_11962,N_11449,N_11699);
nand U11963 (N_11963,N_11623,N_11615);
or U11964 (N_11964,N_11558,N_11504);
or U11965 (N_11965,N_11414,N_11420);
xnor U11966 (N_11966,N_11630,N_11416);
or U11967 (N_11967,N_11663,N_11678);
nand U11968 (N_11968,N_11570,N_11400);
or U11969 (N_11969,N_11693,N_11442);
xnor U11970 (N_11970,N_11469,N_11653);
nor U11971 (N_11971,N_11573,N_11429);
xnor U11972 (N_11972,N_11409,N_11689);
nor U11973 (N_11973,N_11439,N_11486);
nand U11974 (N_11974,N_11638,N_11575);
or U11975 (N_11975,N_11549,N_11598);
xor U11976 (N_11976,N_11565,N_11616);
and U11977 (N_11977,N_11407,N_11652);
nor U11978 (N_11978,N_11605,N_11637);
xor U11979 (N_11979,N_11584,N_11520);
and U11980 (N_11980,N_11515,N_11610);
or U11981 (N_11981,N_11651,N_11567);
nor U11982 (N_11982,N_11418,N_11412);
nand U11983 (N_11983,N_11442,N_11609);
xor U11984 (N_11984,N_11513,N_11410);
nor U11985 (N_11985,N_11667,N_11676);
nand U11986 (N_11986,N_11667,N_11619);
or U11987 (N_11987,N_11646,N_11572);
nor U11988 (N_11988,N_11496,N_11409);
xnor U11989 (N_11989,N_11618,N_11692);
xor U11990 (N_11990,N_11550,N_11631);
nor U11991 (N_11991,N_11634,N_11426);
nand U11992 (N_11992,N_11451,N_11615);
xor U11993 (N_11993,N_11446,N_11658);
xnor U11994 (N_11994,N_11542,N_11458);
xnor U11995 (N_11995,N_11651,N_11432);
and U11996 (N_11996,N_11448,N_11484);
or U11997 (N_11997,N_11605,N_11650);
nor U11998 (N_11998,N_11603,N_11443);
or U11999 (N_11999,N_11485,N_11566);
nand U12000 (N_12000,N_11988,N_11865);
nor U12001 (N_12001,N_11962,N_11918);
nand U12002 (N_12002,N_11750,N_11718);
or U12003 (N_12003,N_11761,N_11730);
or U12004 (N_12004,N_11782,N_11808);
and U12005 (N_12005,N_11846,N_11900);
and U12006 (N_12006,N_11897,N_11763);
nand U12007 (N_12007,N_11714,N_11876);
and U12008 (N_12008,N_11705,N_11956);
nor U12009 (N_12009,N_11810,N_11935);
nand U12010 (N_12010,N_11845,N_11886);
nand U12011 (N_12011,N_11723,N_11993);
xor U12012 (N_12012,N_11771,N_11825);
and U12013 (N_12013,N_11751,N_11816);
nand U12014 (N_12014,N_11767,N_11707);
nor U12015 (N_12015,N_11955,N_11754);
or U12016 (N_12016,N_11938,N_11933);
or U12017 (N_12017,N_11848,N_11983);
xnor U12018 (N_12018,N_11952,N_11857);
or U12019 (N_12019,N_11824,N_11871);
or U12020 (N_12020,N_11787,N_11743);
or U12021 (N_12021,N_11881,N_11940);
xnor U12022 (N_12022,N_11758,N_11789);
or U12023 (N_12023,N_11880,N_11817);
nand U12024 (N_12024,N_11986,N_11995);
xnor U12025 (N_12025,N_11796,N_11928);
xnor U12026 (N_12026,N_11741,N_11890);
and U12027 (N_12027,N_11854,N_11856);
or U12028 (N_12028,N_11981,N_11711);
nor U12029 (N_12029,N_11913,N_11728);
nand U12030 (N_12030,N_11852,N_11954);
nor U12031 (N_12031,N_11894,N_11906);
or U12032 (N_12032,N_11899,N_11802);
nand U12033 (N_12033,N_11943,N_11922);
and U12034 (N_12034,N_11972,N_11964);
and U12035 (N_12035,N_11729,N_11720);
nand U12036 (N_12036,N_11722,N_11831);
and U12037 (N_12037,N_11827,N_11828);
nand U12038 (N_12038,N_11923,N_11987);
and U12039 (N_12039,N_11721,N_11779);
xnor U12040 (N_12040,N_11991,N_11748);
and U12041 (N_12041,N_11959,N_11901);
nor U12042 (N_12042,N_11836,N_11781);
or U12043 (N_12043,N_11821,N_11826);
xnor U12044 (N_12044,N_11910,N_11708);
and U12045 (N_12045,N_11919,N_11784);
nor U12046 (N_12046,N_11920,N_11701);
and U12047 (N_12047,N_11765,N_11949);
nor U12048 (N_12048,N_11961,N_11934);
nor U12049 (N_12049,N_11855,N_11841);
and U12050 (N_12050,N_11804,N_11835);
nand U12051 (N_12051,N_11889,N_11719);
or U12052 (N_12052,N_11715,N_11950);
nor U12053 (N_12053,N_11752,N_11747);
or U12054 (N_12054,N_11878,N_11870);
nor U12055 (N_12055,N_11905,N_11927);
nor U12056 (N_12056,N_11944,N_11974);
or U12057 (N_12057,N_11992,N_11851);
nand U12058 (N_12058,N_11980,N_11749);
xnor U12059 (N_12059,N_11775,N_11853);
and U12060 (N_12060,N_11939,N_11932);
xnor U12061 (N_12061,N_11960,N_11700);
and U12062 (N_12062,N_11760,N_11908);
nand U12063 (N_12063,N_11736,N_11764);
nand U12064 (N_12064,N_11953,N_11734);
nand U12065 (N_12065,N_11970,N_11975);
or U12066 (N_12066,N_11702,N_11822);
nor U12067 (N_12067,N_11921,N_11724);
and U12068 (N_12068,N_11850,N_11811);
nor U12069 (N_12069,N_11777,N_11772);
nand U12070 (N_12070,N_11805,N_11731);
or U12071 (N_12071,N_11757,N_11874);
or U12072 (N_12072,N_11903,N_11829);
and U12073 (N_12073,N_11832,N_11909);
nand U12074 (N_12074,N_11792,N_11717);
or U12075 (N_12075,N_11769,N_11797);
or U12076 (N_12076,N_11873,N_11931);
xor U12077 (N_12077,N_11907,N_11898);
or U12078 (N_12078,N_11716,N_11713);
or U12079 (N_12079,N_11895,N_11925);
or U12080 (N_12080,N_11996,N_11785);
and U12081 (N_12081,N_11997,N_11887);
xor U12082 (N_12082,N_11869,N_11776);
nor U12083 (N_12083,N_11867,N_11888);
nand U12084 (N_12084,N_11778,N_11742);
nand U12085 (N_12085,N_11893,N_11967);
nand U12086 (N_12086,N_11877,N_11947);
and U12087 (N_12087,N_11774,N_11725);
or U12088 (N_12088,N_11969,N_11866);
nor U12089 (N_12089,N_11814,N_11799);
xnor U12090 (N_12090,N_11842,N_11755);
nor U12091 (N_12091,N_11840,N_11712);
xor U12092 (N_12092,N_11976,N_11803);
nor U12093 (N_12093,N_11809,N_11963);
or U12094 (N_12094,N_11818,N_11946);
and U12095 (N_12095,N_11930,N_11830);
nor U12096 (N_12096,N_11733,N_11912);
or U12097 (N_12097,N_11773,N_11861);
nand U12098 (N_12098,N_11982,N_11783);
nand U12099 (N_12099,N_11892,N_11756);
and U12100 (N_12100,N_11801,N_11790);
nand U12101 (N_12101,N_11911,N_11948);
and U12102 (N_12102,N_11989,N_11859);
and U12103 (N_12103,N_11977,N_11902);
nor U12104 (N_12104,N_11999,N_11727);
and U12105 (N_12105,N_11968,N_11709);
xor U12106 (N_12106,N_11914,N_11978);
xor U12107 (N_12107,N_11896,N_11745);
and U12108 (N_12108,N_11726,N_11844);
and U12109 (N_12109,N_11915,N_11847);
nor U12110 (N_12110,N_11863,N_11823);
and U12111 (N_12111,N_11762,N_11891);
or U12112 (N_12112,N_11990,N_11917);
or U12113 (N_12113,N_11735,N_11740);
nand U12114 (N_12114,N_11703,N_11885);
nor U12115 (N_12115,N_11807,N_11957);
nand U12116 (N_12116,N_11704,N_11786);
nand U12117 (N_12117,N_11746,N_11812);
nor U12118 (N_12118,N_11936,N_11780);
nand U12119 (N_12119,N_11904,N_11916);
and U12120 (N_12120,N_11973,N_11806);
or U12121 (N_12121,N_11833,N_11737);
or U12122 (N_12122,N_11860,N_11958);
xnor U12123 (N_12123,N_11872,N_11965);
and U12124 (N_12124,N_11744,N_11985);
or U12125 (N_12125,N_11998,N_11862);
and U12126 (N_12126,N_11794,N_11984);
xor U12127 (N_12127,N_11710,N_11979);
nor U12128 (N_12128,N_11929,N_11971);
and U12129 (N_12129,N_11770,N_11788);
and U12130 (N_12130,N_11868,N_11768);
nor U12131 (N_12131,N_11738,N_11795);
xor U12132 (N_12132,N_11800,N_11883);
or U12133 (N_12133,N_11834,N_11813);
nor U12134 (N_12134,N_11879,N_11864);
and U12135 (N_12135,N_11759,N_11839);
xor U12136 (N_12136,N_11926,N_11994);
and U12137 (N_12137,N_11884,N_11766);
xor U12138 (N_12138,N_11843,N_11706);
and U12139 (N_12139,N_11837,N_11793);
nor U12140 (N_12140,N_11945,N_11941);
xor U12141 (N_12141,N_11966,N_11937);
or U12142 (N_12142,N_11924,N_11875);
xnor U12143 (N_12143,N_11951,N_11798);
and U12144 (N_12144,N_11732,N_11858);
nor U12145 (N_12145,N_11820,N_11942);
xnor U12146 (N_12146,N_11882,N_11838);
and U12147 (N_12147,N_11791,N_11849);
or U12148 (N_12148,N_11739,N_11815);
nand U12149 (N_12149,N_11819,N_11753);
and U12150 (N_12150,N_11707,N_11882);
nand U12151 (N_12151,N_11788,N_11939);
and U12152 (N_12152,N_11856,N_11872);
and U12153 (N_12153,N_11952,N_11939);
xnor U12154 (N_12154,N_11865,N_11714);
nand U12155 (N_12155,N_11707,N_11921);
xnor U12156 (N_12156,N_11986,N_11909);
nor U12157 (N_12157,N_11827,N_11917);
xor U12158 (N_12158,N_11750,N_11769);
nand U12159 (N_12159,N_11708,N_11970);
nor U12160 (N_12160,N_11942,N_11993);
xnor U12161 (N_12161,N_11824,N_11832);
nor U12162 (N_12162,N_11927,N_11882);
nor U12163 (N_12163,N_11900,N_11915);
and U12164 (N_12164,N_11961,N_11887);
and U12165 (N_12165,N_11983,N_11771);
nand U12166 (N_12166,N_11913,N_11796);
nand U12167 (N_12167,N_11941,N_11708);
nor U12168 (N_12168,N_11909,N_11972);
and U12169 (N_12169,N_11912,N_11943);
xor U12170 (N_12170,N_11885,N_11701);
or U12171 (N_12171,N_11973,N_11783);
nand U12172 (N_12172,N_11781,N_11972);
xnor U12173 (N_12173,N_11939,N_11924);
nand U12174 (N_12174,N_11863,N_11957);
xor U12175 (N_12175,N_11938,N_11866);
nand U12176 (N_12176,N_11705,N_11903);
nand U12177 (N_12177,N_11708,N_11907);
and U12178 (N_12178,N_11899,N_11925);
nand U12179 (N_12179,N_11945,N_11706);
xnor U12180 (N_12180,N_11996,N_11758);
or U12181 (N_12181,N_11956,N_11997);
nor U12182 (N_12182,N_11710,N_11836);
and U12183 (N_12183,N_11903,N_11793);
nor U12184 (N_12184,N_11794,N_11983);
or U12185 (N_12185,N_11787,N_11768);
and U12186 (N_12186,N_11998,N_11853);
and U12187 (N_12187,N_11980,N_11883);
nand U12188 (N_12188,N_11914,N_11761);
or U12189 (N_12189,N_11753,N_11841);
nand U12190 (N_12190,N_11831,N_11758);
and U12191 (N_12191,N_11991,N_11872);
nand U12192 (N_12192,N_11842,N_11883);
nand U12193 (N_12193,N_11997,N_11988);
nand U12194 (N_12194,N_11832,N_11971);
and U12195 (N_12195,N_11808,N_11875);
and U12196 (N_12196,N_11982,N_11765);
xor U12197 (N_12197,N_11873,N_11755);
and U12198 (N_12198,N_11824,N_11760);
nand U12199 (N_12199,N_11738,N_11845);
nand U12200 (N_12200,N_11853,N_11762);
and U12201 (N_12201,N_11712,N_11969);
nor U12202 (N_12202,N_11809,N_11928);
xnor U12203 (N_12203,N_11755,N_11780);
nor U12204 (N_12204,N_11761,N_11800);
and U12205 (N_12205,N_11873,N_11803);
nand U12206 (N_12206,N_11846,N_11974);
xnor U12207 (N_12207,N_11857,N_11887);
nand U12208 (N_12208,N_11951,N_11765);
nor U12209 (N_12209,N_11790,N_11798);
xor U12210 (N_12210,N_11700,N_11968);
and U12211 (N_12211,N_11919,N_11968);
and U12212 (N_12212,N_11911,N_11986);
or U12213 (N_12213,N_11796,N_11921);
nand U12214 (N_12214,N_11847,N_11977);
nor U12215 (N_12215,N_11933,N_11790);
and U12216 (N_12216,N_11732,N_11829);
or U12217 (N_12217,N_11869,N_11905);
xor U12218 (N_12218,N_11957,N_11842);
and U12219 (N_12219,N_11841,N_11800);
nor U12220 (N_12220,N_11775,N_11862);
xor U12221 (N_12221,N_11773,N_11740);
or U12222 (N_12222,N_11793,N_11945);
xnor U12223 (N_12223,N_11828,N_11898);
and U12224 (N_12224,N_11760,N_11961);
nand U12225 (N_12225,N_11724,N_11729);
or U12226 (N_12226,N_11784,N_11861);
nand U12227 (N_12227,N_11916,N_11959);
nand U12228 (N_12228,N_11946,N_11985);
or U12229 (N_12229,N_11784,N_11977);
xor U12230 (N_12230,N_11916,N_11781);
or U12231 (N_12231,N_11946,N_11952);
and U12232 (N_12232,N_11964,N_11767);
or U12233 (N_12233,N_11826,N_11976);
or U12234 (N_12234,N_11989,N_11746);
or U12235 (N_12235,N_11860,N_11868);
nand U12236 (N_12236,N_11924,N_11823);
nand U12237 (N_12237,N_11949,N_11720);
nor U12238 (N_12238,N_11873,N_11968);
xnor U12239 (N_12239,N_11929,N_11728);
nand U12240 (N_12240,N_11883,N_11705);
and U12241 (N_12241,N_11993,N_11795);
xnor U12242 (N_12242,N_11764,N_11844);
and U12243 (N_12243,N_11701,N_11732);
and U12244 (N_12244,N_11985,N_11938);
and U12245 (N_12245,N_11718,N_11938);
nand U12246 (N_12246,N_11713,N_11995);
nand U12247 (N_12247,N_11817,N_11967);
nand U12248 (N_12248,N_11941,N_11808);
nand U12249 (N_12249,N_11970,N_11906);
and U12250 (N_12250,N_11916,N_11974);
nand U12251 (N_12251,N_11981,N_11917);
or U12252 (N_12252,N_11785,N_11958);
xnor U12253 (N_12253,N_11923,N_11902);
or U12254 (N_12254,N_11837,N_11815);
xor U12255 (N_12255,N_11861,N_11958);
nand U12256 (N_12256,N_11875,N_11750);
or U12257 (N_12257,N_11748,N_11756);
or U12258 (N_12258,N_11780,N_11964);
xnor U12259 (N_12259,N_11979,N_11904);
nand U12260 (N_12260,N_11829,N_11868);
nor U12261 (N_12261,N_11945,N_11831);
and U12262 (N_12262,N_11836,N_11817);
xnor U12263 (N_12263,N_11996,N_11977);
xor U12264 (N_12264,N_11932,N_11975);
xnor U12265 (N_12265,N_11718,N_11706);
or U12266 (N_12266,N_11798,N_11747);
nand U12267 (N_12267,N_11800,N_11864);
nor U12268 (N_12268,N_11862,N_11711);
xnor U12269 (N_12269,N_11840,N_11921);
and U12270 (N_12270,N_11759,N_11912);
and U12271 (N_12271,N_11957,N_11768);
nor U12272 (N_12272,N_11815,N_11970);
nand U12273 (N_12273,N_11943,N_11910);
nand U12274 (N_12274,N_11789,N_11838);
and U12275 (N_12275,N_11984,N_11848);
nand U12276 (N_12276,N_11737,N_11963);
xnor U12277 (N_12277,N_11980,N_11812);
nor U12278 (N_12278,N_11939,N_11748);
nor U12279 (N_12279,N_11760,N_11874);
nand U12280 (N_12280,N_11776,N_11821);
and U12281 (N_12281,N_11842,N_11781);
nand U12282 (N_12282,N_11739,N_11706);
and U12283 (N_12283,N_11926,N_11806);
nor U12284 (N_12284,N_11791,N_11761);
nand U12285 (N_12285,N_11923,N_11928);
nor U12286 (N_12286,N_11706,N_11791);
xnor U12287 (N_12287,N_11994,N_11846);
xor U12288 (N_12288,N_11777,N_11980);
xnor U12289 (N_12289,N_11918,N_11932);
or U12290 (N_12290,N_11818,N_11923);
xnor U12291 (N_12291,N_11954,N_11913);
or U12292 (N_12292,N_11835,N_11969);
xor U12293 (N_12293,N_11809,N_11750);
or U12294 (N_12294,N_11911,N_11897);
and U12295 (N_12295,N_11994,N_11819);
nor U12296 (N_12296,N_11795,N_11897);
or U12297 (N_12297,N_11855,N_11972);
nand U12298 (N_12298,N_11774,N_11786);
and U12299 (N_12299,N_11900,N_11765);
xor U12300 (N_12300,N_12197,N_12281);
xnor U12301 (N_12301,N_12073,N_12104);
and U12302 (N_12302,N_12019,N_12156);
nor U12303 (N_12303,N_12222,N_12256);
nand U12304 (N_12304,N_12078,N_12214);
nor U12305 (N_12305,N_12145,N_12259);
and U12306 (N_12306,N_12223,N_12040);
and U12307 (N_12307,N_12075,N_12097);
xor U12308 (N_12308,N_12129,N_12157);
xnor U12309 (N_12309,N_12143,N_12125);
xor U12310 (N_12310,N_12174,N_12043);
and U12311 (N_12311,N_12207,N_12182);
nor U12312 (N_12312,N_12224,N_12120);
and U12313 (N_12313,N_12263,N_12124);
nor U12314 (N_12314,N_12116,N_12258);
nand U12315 (N_12315,N_12006,N_12204);
xor U12316 (N_12316,N_12053,N_12277);
nand U12317 (N_12317,N_12250,N_12049);
and U12318 (N_12318,N_12242,N_12159);
nor U12319 (N_12319,N_12035,N_12177);
and U12320 (N_12320,N_12131,N_12192);
and U12321 (N_12321,N_12213,N_12126);
or U12322 (N_12322,N_12220,N_12121);
nand U12323 (N_12323,N_12058,N_12024);
or U12324 (N_12324,N_12070,N_12202);
nor U12325 (N_12325,N_12168,N_12099);
nor U12326 (N_12326,N_12090,N_12028);
nor U12327 (N_12327,N_12151,N_12030);
nor U12328 (N_12328,N_12173,N_12096);
nand U12329 (N_12329,N_12294,N_12023);
nor U12330 (N_12330,N_12094,N_12178);
xor U12331 (N_12331,N_12188,N_12257);
nor U12332 (N_12332,N_12288,N_12239);
and U12333 (N_12333,N_12016,N_12240);
nand U12334 (N_12334,N_12119,N_12015);
xnor U12335 (N_12335,N_12252,N_12087);
nand U12336 (N_12336,N_12198,N_12051);
nand U12337 (N_12337,N_12191,N_12065);
xor U12338 (N_12338,N_12228,N_12147);
nor U12339 (N_12339,N_12152,N_12260);
xor U12340 (N_12340,N_12068,N_12295);
xor U12341 (N_12341,N_12190,N_12158);
nand U12342 (N_12342,N_12175,N_12215);
and U12343 (N_12343,N_12055,N_12000);
xnor U12344 (N_12344,N_12025,N_12086);
nor U12345 (N_12345,N_12088,N_12118);
or U12346 (N_12346,N_12271,N_12013);
or U12347 (N_12347,N_12117,N_12128);
nand U12348 (N_12348,N_12272,N_12189);
xnor U12349 (N_12349,N_12140,N_12203);
nor U12350 (N_12350,N_12251,N_12005);
nand U12351 (N_12351,N_12185,N_12243);
and U12352 (N_12352,N_12254,N_12122);
and U12353 (N_12353,N_12267,N_12238);
or U12354 (N_12354,N_12180,N_12225);
or U12355 (N_12355,N_12210,N_12160);
and U12356 (N_12356,N_12027,N_12166);
and U12357 (N_12357,N_12150,N_12226);
nor U12358 (N_12358,N_12093,N_12001);
nor U12359 (N_12359,N_12020,N_12249);
nor U12360 (N_12360,N_12276,N_12183);
or U12361 (N_12361,N_12036,N_12021);
and U12362 (N_12362,N_12261,N_12084);
nor U12363 (N_12363,N_12039,N_12031);
xor U12364 (N_12364,N_12292,N_12149);
xor U12365 (N_12365,N_12007,N_12161);
nor U12366 (N_12366,N_12022,N_12184);
or U12367 (N_12367,N_12237,N_12244);
xor U12368 (N_12368,N_12136,N_12110);
and U12369 (N_12369,N_12103,N_12217);
or U12370 (N_12370,N_12176,N_12056);
nand U12371 (N_12371,N_12010,N_12105);
and U12372 (N_12372,N_12195,N_12127);
nand U12373 (N_12373,N_12080,N_12113);
xnor U12374 (N_12374,N_12245,N_12106);
xnor U12375 (N_12375,N_12285,N_12011);
or U12376 (N_12376,N_12045,N_12123);
xnor U12377 (N_12377,N_12264,N_12199);
xnor U12378 (N_12378,N_12268,N_12229);
xnor U12379 (N_12379,N_12227,N_12208);
nand U12380 (N_12380,N_12026,N_12231);
nand U12381 (N_12381,N_12291,N_12059);
nor U12382 (N_12382,N_12091,N_12050);
or U12383 (N_12383,N_12092,N_12296);
xnor U12384 (N_12384,N_12179,N_12003);
nor U12385 (N_12385,N_12109,N_12139);
xor U12386 (N_12386,N_12141,N_12172);
nor U12387 (N_12387,N_12289,N_12034);
nor U12388 (N_12388,N_12241,N_12200);
nand U12389 (N_12389,N_12062,N_12299);
nor U12390 (N_12390,N_12235,N_12262);
nand U12391 (N_12391,N_12008,N_12218);
nor U12392 (N_12392,N_12234,N_12163);
nand U12393 (N_12393,N_12298,N_12077);
xor U12394 (N_12394,N_12282,N_12221);
or U12395 (N_12395,N_12293,N_12212);
and U12396 (N_12396,N_12046,N_12201);
nor U12397 (N_12397,N_12082,N_12108);
and U12398 (N_12398,N_12095,N_12002);
nand U12399 (N_12399,N_12209,N_12057);
xor U12400 (N_12400,N_12287,N_12278);
and U12401 (N_12401,N_12134,N_12089);
or U12402 (N_12402,N_12297,N_12211);
and U12403 (N_12403,N_12255,N_12048);
or U12404 (N_12404,N_12194,N_12133);
nor U12405 (N_12405,N_12266,N_12098);
nor U12406 (N_12406,N_12083,N_12216);
xnor U12407 (N_12407,N_12066,N_12004);
xor U12408 (N_12408,N_12279,N_12232);
xnor U12409 (N_12409,N_12033,N_12085);
or U12410 (N_12410,N_12269,N_12193);
nand U12411 (N_12411,N_12196,N_12018);
xnor U12412 (N_12412,N_12069,N_12165);
nor U12413 (N_12413,N_12072,N_12067);
or U12414 (N_12414,N_12270,N_12012);
nand U12415 (N_12415,N_12038,N_12187);
nand U12416 (N_12416,N_12162,N_12060);
or U12417 (N_12417,N_12061,N_12169);
nand U12418 (N_12418,N_12181,N_12219);
and U12419 (N_12419,N_12107,N_12284);
or U12420 (N_12420,N_12236,N_12064);
or U12421 (N_12421,N_12047,N_12273);
xor U12422 (N_12422,N_12167,N_12074);
nand U12423 (N_12423,N_12206,N_12014);
xnor U12424 (N_12424,N_12171,N_12044);
nor U12425 (N_12425,N_12114,N_12265);
nand U12426 (N_12426,N_12029,N_12164);
nor U12427 (N_12427,N_12286,N_12246);
xnor U12428 (N_12428,N_12233,N_12230);
and U12429 (N_12429,N_12155,N_12081);
and U12430 (N_12430,N_12100,N_12115);
nor U12431 (N_12431,N_12132,N_12076);
or U12432 (N_12432,N_12041,N_12135);
xor U12433 (N_12433,N_12042,N_12130);
xor U12434 (N_12434,N_12148,N_12253);
nand U12435 (N_12435,N_12146,N_12138);
nand U12436 (N_12436,N_12079,N_12102);
nand U12437 (N_12437,N_12186,N_12111);
and U12438 (N_12438,N_12032,N_12280);
or U12439 (N_12439,N_12063,N_12137);
and U12440 (N_12440,N_12142,N_12054);
or U12441 (N_12441,N_12283,N_12037);
nand U12442 (N_12442,N_12290,N_12017);
nor U12443 (N_12443,N_12248,N_12071);
or U12444 (N_12444,N_12247,N_12144);
nor U12445 (N_12445,N_12153,N_12274);
nand U12446 (N_12446,N_12052,N_12170);
nand U12447 (N_12447,N_12205,N_12154);
nor U12448 (N_12448,N_12275,N_12101);
and U12449 (N_12449,N_12112,N_12009);
and U12450 (N_12450,N_12100,N_12237);
nand U12451 (N_12451,N_12287,N_12006);
and U12452 (N_12452,N_12106,N_12023);
and U12453 (N_12453,N_12136,N_12170);
xor U12454 (N_12454,N_12068,N_12117);
xor U12455 (N_12455,N_12125,N_12169);
and U12456 (N_12456,N_12290,N_12129);
and U12457 (N_12457,N_12018,N_12044);
and U12458 (N_12458,N_12071,N_12186);
nor U12459 (N_12459,N_12169,N_12111);
and U12460 (N_12460,N_12085,N_12159);
or U12461 (N_12461,N_12215,N_12177);
or U12462 (N_12462,N_12204,N_12187);
or U12463 (N_12463,N_12201,N_12247);
nor U12464 (N_12464,N_12284,N_12066);
nand U12465 (N_12465,N_12223,N_12139);
or U12466 (N_12466,N_12096,N_12126);
nand U12467 (N_12467,N_12231,N_12162);
or U12468 (N_12468,N_12282,N_12169);
nor U12469 (N_12469,N_12209,N_12151);
xnor U12470 (N_12470,N_12157,N_12131);
nor U12471 (N_12471,N_12272,N_12099);
or U12472 (N_12472,N_12161,N_12098);
and U12473 (N_12473,N_12131,N_12051);
nand U12474 (N_12474,N_12111,N_12139);
and U12475 (N_12475,N_12040,N_12042);
and U12476 (N_12476,N_12015,N_12128);
nor U12477 (N_12477,N_12192,N_12278);
xnor U12478 (N_12478,N_12292,N_12257);
nand U12479 (N_12479,N_12197,N_12206);
or U12480 (N_12480,N_12122,N_12296);
xnor U12481 (N_12481,N_12017,N_12175);
and U12482 (N_12482,N_12254,N_12256);
nand U12483 (N_12483,N_12238,N_12199);
nand U12484 (N_12484,N_12136,N_12298);
nor U12485 (N_12485,N_12249,N_12251);
xnor U12486 (N_12486,N_12298,N_12254);
nor U12487 (N_12487,N_12284,N_12115);
xor U12488 (N_12488,N_12107,N_12137);
nand U12489 (N_12489,N_12158,N_12096);
and U12490 (N_12490,N_12005,N_12101);
and U12491 (N_12491,N_12252,N_12223);
nand U12492 (N_12492,N_12272,N_12081);
xor U12493 (N_12493,N_12029,N_12094);
xnor U12494 (N_12494,N_12052,N_12261);
and U12495 (N_12495,N_12243,N_12118);
or U12496 (N_12496,N_12162,N_12033);
xnor U12497 (N_12497,N_12188,N_12047);
nor U12498 (N_12498,N_12239,N_12059);
nand U12499 (N_12499,N_12204,N_12284);
xnor U12500 (N_12500,N_12089,N_12265);
xor U12501 (N_12501,N_12064,N_12267);
nor U12502 (N_12502,N_12075,N_12199);
nand U12503 (N_12503,N_12197,N_12019);
and U12504 (N_12504,N_12264,N_12194);
and U12505 (N_12505,N_12044,N_12169);
nand U12506 (N_12506,N_12063,N_12062);
or U12507 (N_12507,N_12014,N_12236);
or U12508 (N_12508,N_12121,N_12113);
nor U12509 (N_12509,N_12006,N_12154);
nand U12510 (N_12510,N_12024,N_12083);
nor U12511 (N_12511,N_12248,N_12047);
nor U12512 (N_12512,N_12045,N_12199);
and U12513 (N_12513,N_12299,N_12144);
nor U12514 (N_12514,N_12224,N_12106);
nor U12515 (N_12515,N_12280,N_12034);
nand U12516 (N_12516,N_12207,N_12293);
nor U12517 (N_12517,N_12149,N_12169);
nand U12518 (N_12518,N_12185,N_12147);
or U12519 (N_12519,N_12082,N_12166);
and U12520 (N_12520,N_12183,N_12130);
nand U12521 (N_12521,N_12194,N_12285);
nand U12522 (N_12522,N_12188,N_12076);
or U12523 (N_12523,N_12079,N_12004);
nor U12524 (N_12524,N_12245,N_12287);
nor U12525 (N_12525,N_12110,N_12062);
and U12526 (N_12526,N_12019,N_12089);
xor U12527 (N_12527,N_12274,N_12288);
or U12528 (N_12528,N_12298,N_12162);
nor U12529 (N_12529,N_12238,N_12090);
and U12530 (N_12530,N_12219,N_12030);
or U12531 (N_12531,N_12276,N_12207);
nor U12532 (N_12532,N_12250,N_12041);
nand U12533 (N_12533,N_12097,N_12112);
nor U12534 (N_12534,N_12247,N_12269);
xnor U12535 (N_12535,N_12148,N_12124);
xor U12536 (N_12536,N_12202,N_12156);
nand U12537 (N_12537,N_12157,N_12244);
and U12538 (N_12538,N_12267,N_12233);
xor U12539 (N_12539,N_12228,N_12194);
and U12540 (N_12540,N_12126,N_12085);
nand U12541 (N_12541,N_12013,N_12156);
or U12542 (N_12542,N_12215,N_12146);
and U12543 (N_12543,N_12053,N_12046);
or U12544 (N_12544,N_12007,N_12273);
xnor U12545 (N_12545,N_12028,N_12197);
nand U12546 (N_12546,N_12149,N_12259);
or U12547 (N_12547,N_12045,N_12155);
and U12548 (N_12548,N_12032,N_12019);
xnor U12549 (N_12549,N_12277,N_12117);
or U12550 (N_12550,N_12108,N_12165);
or U12551 (N_12551,N_12275,N_12090);
nand U12552 (N_12552,N_12034,N_12288);
nor U12553 (N_12553,N_12206,N_12130);
nor U12554 (N_12554,N_12273,N_12160);
or U12555 (N_12555,N_12266,N_12097);
nand U12556 (N_12556,N_12238,N_12214);
nor U12557 (N_12557,N_12033,N_12029);
nand U12558 (N_12558,N_12032,N_12067);
or U12559 (N_12559,N_12205,N_12078);
and U12560 (N_12560,N_12124,N_12186);
and U12561 (N_12561,N_12124,N_12072);
and U12562 (N_12562,N_12182,N_12049);
or U12563 (N_12563,N_12010,N_12144);
and U12564 (N_12564,N_12256,N_12161);
xnor U12565 (N_12565,N_12211,N_12137);
xor U12566 (N_12566,N_12032,N_12178);
nor U12567 (N_12567,N_12275,N_12178);
nor U12568 (N_12568,N_12185,N_12180);
and U12569 (N_12569,N_12080,N_12284);
and U12570 (N_12570,N_12008,N_12269);
and U12571 (N_12571,N_12115,N_12288);
nor U12572 (N_12572,N_12255,N_12036);
or U12573 (N_12573,N_12226,N_12274);
and U12574 (N_12574,N_12129,N_12219);
xor U12575 (N_12575,N_12282,N_12010);
xnor U12576 (N_12576,N_12040,N_12147);
and U12577 (N_12577,N_12092,N_12114);
nand U12578 (N_12578,N_12090,N_12248);
nor U12579 (N_12579,N_12018,N_12263);
nand U12580 (N_12580,N_12113,N_12256);
nor U12581 (N_12581,N_12204,N_12064);
and U12582 (N_12582,N_12290,N_12014);
or U12583 (N_12583,N_12128,N_12140);
nor U12584 (N_12584,N_12217,N_12040);
nor U12585 (N_12585,N_12194,N_12041);
nor U12586 (N_12586,N_12199,N_12122);
xnor U12587 (N_12587,N_12224,N_12040);
or U12588 (N_12588,N_12098,N_12240);
nor U12589 (N_12589,N_12242,N_12295);
nand U12590 (N_12590,N_12083,N_12093);
nand U12591 (N_12591,N_12232,N_12130);
and U12592 (N_12592,N_12271,N_12079);
nor U12593 (N_12593,N_12231,N_12224);
or U12594 (N_12594,N_12118,N_12179);
and U12595 (N_12595,N_12135,N_12042);
nand U12596 (N_12596,N_12164,N_12106);
nor U12597 (N_12597,N_12017,N_12083);
xnor U12598 (N_12598,N_12251,N_12000);
and U12599 (N_12599,N_12063,N_12068);
nand U12600 (N_12600,N_12568,N_12400);
xnor U12601 (N_12601,N_12499,N_12432);
nand U12602 (N_12602,N_12488,N_12367);
and U12603 (N_12603,N_12575,N_12375);
or U12604 (N_12604,N_12403,N_12550);
nand U12605 (N_12605,N_12387,N_12438);
nand U12606 (N_12606,N_12360,N_12402);
xor U12607 (N_12607,N_12474,N_12406);
xor U12608 (N_12608,N_12490,N_12439);
and U12609 (N_12609,N_12519,N_12437);
xor U12610 (N_12610,N_12413,N_12527);
nand U12611 (N_12611,N_12487,N_12492);
xor U12612 (N_12612,N_12334,N_12396);
nand U12613 (N_12613,N_12530,N_12392);
nor U12614 (N_12614,N_12513,N_12498);
nor U12615 (N_12615,N_12484,N_12370);
nand U12616 (N_12616,N_12470,N_12328);
or U12617 (N_12617,N_12539,N_12430);
or U12618 (N_12618,N_12457,N_12566);
and U12619 (N_12619,N_12503,N_12314);
nor U12620 (N_12620,N_12338,N_12471);
nand U12621 (N_12621,N_12572,N_12570);
nand U12622 (N_12622,N_12386,N_12401);
xor U12623 (N_12623,N_12565,N_12586);
xnor U12624 (N_12624,N_12440,N_12311);
and U12625 (N_12625,N_12379,N_12455);
xor U12626 (N_12626,N_12497,N_12461);
nor U12627 (N_12627,N_12306,N_12472);
or U12628 (N_12628,N_12502,N_12380);
and U12629 (N_12629,N_12300,N_12535);
and U12630 (N_12630,N_12336,N_12398);
or U12631 (N_12631,N_12344,N_12468);
nand U12632 (N_12632,N_12592,N_12473);
nor U12633 (N_12633,N_12394,N_12359);
and U12634 (N_12634,N_12365,N_12424);
nand U12635 (N_12635,N_12304,N_12485);
or U12636 (N_12636,N_12463,N_12573);
nand U12637 (N_12637,N_12378,N_12558);
nor U12638 (N_12638,N_12361,N_12441);
or U12639 (N_12639,N_12552,N_12525);
nor U12640 (N_12640,N_12511,N_12557);
or U12641 (N_12641,N_12559,N_12467);
and U12642 (N_12642,N_12416,N_12547);
xnor U12643 (N_12643,N_12358,N_12397);
nand U12644 (N_12644,N_12518,N_12579);
and U12645 (N_12645,N_12594,N_12551);
nand U12646 (N_12646,N_12301,N_12506);
nand U12647 (N_12647,N_12451,N_12454);
or U12648 (N_12648,N_12352,N_12313);
and U12649 (N_12649,N_12521,N_12390);
nor U12650 (N_12650,N_12408,N_12417);
nand U12651 (N_12651,N_12371,N_12409);
or U12652 (N_12652,N_12383,N_12372);
xnor U12653 (N_12653,N_12320,N_12373);
xnor U12654 (N_12654,N_12464,N_12353);
nor U12655 (N_12655,N_12590,N_12593);
and U12656 (N_12656,N_12449,N_12549);
or U12657 (N_12657,N_12486,N_12308);
nor U12658 (N_12658,N_12591,N_12391);
or U12659 (N_12659,N_12429,N_12374);
nand U12660 (N_12660,N_12421,N_12447);
and U12661 (N_12661,N_12460,N_12480);
nor U12662 (N_12662,N_12567,N_12536);
or U12663 (N_12663,N_12330,N_12562);
and U12664 (N_12664,N_12310,N_12415);
nand U12665 (N_12665,N_12369,N_12302);
nor U12666 (N_12666,N_12450,N_12425);
or U12667 (N_12667,N_12532,N_12571);
or U12668 (N_12668,N_12305,N_12587);
nand U12669 (N_12669,N_12393,N_12541);
or U12670 (N_12670,N_12595,N_12599);
nor U12671 (N_12671,N_12533,N_12509);
or U12672 (N_12672,N_12520,N_12433);
or U12673 (N_12673,N_12462,N_12517);
and U12674 (N_12674,N_12459,N_12428);
and U12675 (N_12675,N_12577,N_12576);
and U12676 (N_12676,N_12582,N_12312);
nor U12677 (N_12677,N_12381,N_12508);
or U12678 (N_12678,N_12355,N_12544);
nor U12679 (N_12679,N_12411,N_12340);
or U12680 (N_12680,N_12585,N_12448);
nor U12681 (N_12681,N_12588,N_12366);
nor U12682 (N_12682,N_12356,N_12423);
nand U12683 (N_12683,N_12345,N_12598);
and U12684 (N_12684,N_12542,N_12404);
nand U12685 (N_12685,N_12466,N_12507);
nor U12686 (N_12686,N_12325,N_12548);
nor U12687 (N_12687,N_12555,N_12427);
xor U12688 (N_12688,N_12405,N_12434);
and U12689 (N_12689,N_12368,N_12540);
and U12690 (N_12690,N_12331,N_12563);
nor U12691 (N_12691,N_12420,N_12335);
nand U12692 (N_12692,N_12316,N_12389);
nor U12693 (N_12693,N_12435,N_12496);
nor U12694 (N_12694,N_12426,N_12343);
or U12695 (N_12695,N_12333,N_12538);
and U12696 (N_12696,N_12436,N_12456);
nor U12697 (N_12697,N_12317,N_12537);
xor U12698 (N_12698,N_12357,N_12418);
or U12699 (N_12699,N_12349,N_12385);
or U12700 (N_12700,N_12578,N_12307);
nor U12701 (N_12701,N_12554,N_12510);
xor U12702 (N_12702,N_12443,N_12553);
and U12703 (N_12703,N_12322,N_12442);
nor U12704 (N_12704,N_12494,N_12363);
and U12705 (N_12705,N_12476,N_12339);
or U12706 (N_12706,N_12465,N_12501);
or U12707 (N_12707,N_12453,N_12581);
nor U12708 (N_12708,N_12388,N_12522);
nand U12709 (N_12709,N_12399,N_12446);
and U12710 (N_12710,N_12444,N_12412);
xor U12711 (N_12711,N_12584,N_12445);
nor U12712 (N_12712,N_12376,N_12545);
nand U12713 (N_12713,N_12303,N_12597);
and U12714 (N_12714,N_12348,N_12337);
nand U12715 (N_12715,N_12534,N_12431);
nand U12716 (N_12716,N_12351,N_12469);
and U12717 (N_12717,N_12481,N_12362);
nor U12718 (N_12718,N_12482,N_12524);
nand U12719 (N_12719,N_12419,N_12309);
or U12720 (N_12720,N_12318,N_12346);
xnor U12721 (N_12721,N_12543,N_12364);
and U12722 (N_12722,N_12479,N_12329);
xnor U12723 (N_12723,N_12504,N_12512);
nand U12724 (N_12724,N_12347,N_12327);
xor U12725 (N_12725,N_12560,N_12546);
nor U12726 (N_12726,N_12382,N_12324);
and U12727 (N_12727,N_12514,N_12458);
and U12728 (N_12728,N_12589,N_12452);
nor U12729 (N_12729,N_12332,N_12564);
or U12730 (N_12730,N_12477,N_12516);
or U12731 (N_12731,N_12515,N_12414);
nor U12732 (N_12732,N_12377,N_12596);
nand U12733 (N_12733,N_12354,N_12495);
and U12734 (N_12734,N_12528,N_12489);
nand U12735 (N_12735,N_12326,N_12531);
xnor U12736 (N_12736,N_12583,N_12321);
xnor U12737 (N_12737,N_12523,N_12556);
xnor U12738 (N_12738,N_12491,N_12384);
nor U12739 (N_12739,N_12315,N_12422);
xnor U12740 (N_12740,N_12319,N_12407);
xor U12741 (N_12741,N_12478,N_12574);
nand U12742 (N_12742,N_12341,N_12529);
nand U12743 (N_12743,N_12410,N_12350);
and U12744 (N_12744,N_12561,N_12580);
or U12745 (N_12745,N_12323,N_12526);
or U12746 (N_12746,N_12505,N_12493);
or U12747 (N_12747,N_12475,N_12483);
or U12748 (N_12748,N_12500,N_12342);
xnor U12749 (N_12749,N_12569,N_12395);
or U12750 (N_12750,N_12582,N_12482);
nand U12751 (N_12751,N_12472,N_12573);
nand U12752 (N_12752,N_12445,N_12499);
xor U12753 (N_12753,N_12561,N_12454);
or U12754 (N_12754,N_12342,N_12309);
or U12755 (N_12755,N_12571,N_12415);
and U12756 (N_12756,N_12429,N_12396);
or U12757 (N_12757,N_12311,N_12319);
and U12758 (N_12758,N_12389,N_12335);
or U12759 (N_12759,N_12341,N_12362);
nand U12760 (N_12760,N_12492,N_12348);
nand U12761 (N_12761,N_12450,N_12542);
nor U12762 (N_12762,N_12395,N_12439);
nor U12763 (N_12763,N_12385,N_12386);
and U12764 (N_12764,N_12350,N_12523);
and U12765 (N_12765,N_12486,N_12585);
xor U12766 (N_12766,N_12516,N_12416);
or U12767 (N_12767,N_12395,N_12418);
nand U12768 (N_12768,N_12405,N_12303);
or U12769 (N_12769,N_12355,N_12562);
or U12770 (N_12770,N_12588,N_12473);
xnor U12771 (N_12771,N_12305,N_12468);
and U12772 (N_12772,N_12523,N_12398);
or U12773 (N_12773,N_12306,N_12404);
nand U12774 (N_12774,N_12337,N_12419);
xnor U12775 (N_12775,N_12508,N_12396);
xnor U12776 (N_12776,N_12379,N_12573);
or U12777 (N_12777,N_12471,N_12475);
xor U12778 (N_12778,N_12395,N_12448);
or U12779 (N_12779,N_12438,N_12497);
or U12780 (N_12780,N_12314,N_12523);
and U12781 (N_12781,N_12390,N_12519);
and U12782 (N_12782,N_12305,N_12504);
or U12783 (N_12783,N_12304,N_12443);
or U12784 (N_12784,N_12446,N_12586);
xnor U12785 (N_12785,N_12496,N_12423);
xnor U12786 (N_12786,N_12363,N_12411);
nand U12787 (N_12787,N_12359,N_12474);
or U12788 (N_12788,N_12449,N_12452);
xor U12789 (N_12789,N_12330,N_12533);
and U12790 (N_12790,N_12418,N_12572);
and U12791 (N_12791,N_12338,N_12543);
nor U12792 (N_12792,N_12464,N_12574);
nor U12793 (N_12793,N_12306,N_12588);
or U12794 (N_12794,N_12575,N_12494);
and U12795 (N_12795,N_12436,N_12485);
and U12796 (N_12796,N_12460,N_12434);
and U12797 (N_12797,N_12380,N_12599);
and U12798 (N_12798,N_12504,N_12458);
nor U12799 (N_12799,N_12436,N_12473);
or U12800 (N_12800,N_12525,N_12599);
nand U12801 (N_12801,N_12496,N_12320);
nor U12802 (N_12802,N_12599,N_12324);
nor U12803 (N_12803,N_12526,N_12447);
xor U12804 (N_12804,N_12337,N_12382);
xor U12805 (N_12805,N_12309,N_12493);
nand U12806 (N_12806,N_12383,N_12411);
nor U12807 (N_12807,N_12347,N_12436);
xor U12808 (N_12808,N_12450,N_12309);
or U12809 (N_12809,N_12343,N_12407);
or U12810 (N_12810,N_12521,N_12454);
nand U12811 (N_12811,N_12594,N_12472);
xor U12812 (N_12812,N_12482,N_12350);
xor U12813 (N_12813,N_12358,N_12483);
nor U12814 (N_12814,N_12462,N_12465);
or U12815 (N_12815,N_12524,N_12326);
nor U12816 (N_12816,N_12555,N_12465);
and U12817 (N_12817,N_12326,N_12500);
nor U12818 (N_12818,N_12369,N_12474);
nor U12819 (N_12819,N_12472,N_12490);
xor U12820 (N_12820,N_12566,N_12305);
nand U12821 (N_12821,N_12462,N_12410);
and U12822 (N_12822,N_12574,N_12437);
nor U12823 (N_12823,N_12369,N_12389);
xor U12824 (N_12824,N_12316,N_12592);
nand U12825 (N_12825,N_12342,N_12323);
nor U12826 (N_12826,N_12450,N_12338);
nand U12827 (N_12827,N_12501,N_12587);
nor U12828 (N_12828,N_12493,N_12301);
nor U12829 (N_12829,N_12388,N_12311);
and U12830 (N_12830,N_12586,N_12579);
or U12831 (N_12831,N_12367,N_12475);
and U12832 (N_12832,N_12326,N_12428);
xor U12833 (N_12833,N_12418,N_12522);
nor U12834 (N_12834,N_12593,N_12350);
and U12835 (N_12835,N_12361,N_12322);
xor U12836 (N_12836,N_12423,N_12537);
xnor U12837 (N_12837,N_12595,N_12542);
or U12838 (N_12838,N_12397,N_12518);
and U12839 (N_12839,N_12592,N_12455);
and U12840 (N_12840,N_12581,N_12479);
nand U12841 (N_12841,N_12374,N_12584);
nor U12842 (N_12842,N_12568,N_12316);
and U12843 (N_12843,N_12488,N_12325);
xor U12844 (N_12844,N_12516,N_12573);
xnor U12845 (N_12845,N_12526,N_12303);
nand U12846 (N_12846,N_12563,N_12414);
and U12847 (N_12847,N_12343,N_12583);
or U12848 (N_12848,N_12348,N_12429);
nor U12849 (N_12849,N_12328,N_12316);
xnor U12850 (N_12850,N_12490,N_12401);
and U12851 (N_12851,N_12328,N_12523);
nand U12852 (N_12852,N_12417,N_12521);
nand U12853 (N_12853,N_12575,N_12429);
and U12854 (N_12854,N_12459,N_12433);
or U12855 (N_12855,N_12561,N_12379);
and U12856 (N_12856,N_12338,N_12386);
or U12857 (N_12857,N_12336,N_12327);
or U12858 (N_12858,N_12409,N_12509);
or U12859 (N_12859,N_12401,N_12410);
or U12860 (N_12860,N_12591,N_12587);
nand U12861 (N_12861,N_12346,N_12486);
and U12862 (N_12862,N_12498,N_12439);
nor U12863 (N_12863,N_12473,N_12472);
nand U12864 (N_12864,N_12436,N_12528);
and U12865 (N_12865,N_12532,N_12418);
nand U12866 (N_12866,N_12495,N_12589);
or U12867 (N_12867,N_12545,N_12535);
nor U12868 (N_12868,N_12542,N_12326);
xnor U12869 (N_12869,N_12558,N_12464);
and U12870 (N_12870,N_12500,N_12438);
or U12871 (N_12871,N_12355,N_12599);
or U12872 (N_12872,N_12397,N_12333);
or U12873 (N_12873,N_12466,N_12583);
and U12874 (N_12874,N_12561,N_12587);
nor U12875 (N_12875,N_12418,N_12368);
xor U12876 (N_12876,N_12328,N_12386);
nand U12877 (N_12877,N_12392,N_12303);
nor U12878 (N_12878,N_12321,N_12464);
or U12879 (N_12879,N_12448,N_12576);
nor U12880 (N_12880,N_12385,N_12371);
and U12881 (N_12881,N_12568,N_12545);
nand U12882 (N_12882,N_12397,N_12345);
nand U12883 (N_12883,N_12502,N_12519);
or U12884 (N_12884,N_12306,N_12561);
or U12885 (N_12885,N_12447,N_12511);
nor U12886 (N_12886,N_12410,N_12390);
nand U12887 (N_12887,N_12382,N_12374);
or U12888 (N_12888,N_12414,N_12305);
and U12889 (N_12889,N_12375,N_12544);
or U12890 (N_12890,N_12486,N_12404);
xnor U12891 (N_12891,N_12451,N_12588);
nor U12892 (N_12892,N_12526,N_12398);
xnor U12893 (N_12893,N_12399,N_12332);
nand U12894 (N_12894,N_12449,N_12314);
nand U12895 (N_12895,N_12526,N_12549);
nand U12896 (N_12896,N_12311,N_12513);
nand U12897 (N_12897,N_12389,N_12515);
xor U12898 (N_12898,N_12399,N_12559);
nand U12899 (N_12899,N_12350,N_12566);
xnor U12900 (N_12900,N_12814,N_12897);
and U12901 (N_12901,N_12763,N_12896);
and U12902 (N_12902,N_12734,N_12833);
and U12903 (N_12903,N_12676,N_12788);
xnor U12904 (N_12904,N_12824,N_12672);
nand U12905 (N_12905,N_12632,N_12805);
and U12906 (N_12906,N_12783,N_12646);
or U12907 (N_12907,N_12859,N_12652);
and U12908 (N_12908,N_12670,N_12819);
xnor U12909 (N_12909,N_12848,N_12780);
xor U12910 (N_12910,N_12879,N_12841);
nor U12911 (N_12911,N_12888,N_12750);
or U12912 (N_12912,N_12784,N_12803);
and U12913 (N_12913,N_12615,N_12874);
nor U12914 (N_12914,N_12630,N_12643);
or U12915 (N_12915,N_12785,N_12741);
and U12916 (N_12916,N_12600,N_12886);
nor U12917 (N_12917,N_12872,N_12611);
and U12918 (N_12918,N_12602,N_12873);
and U12919 (N_12919,N_12705,N_12636);
nor U12920 (N_12920,N_12802,N_12877);
and U12921 (N_12921,N_12810,N_12661);
or U12922 (N_12922,N_12826,N_12771);
or U12923 (N_12923,N_12700,N_12601);
or U12924 (N_12924,N_12622,N_12773);
nor U12925 (N_12925,N_12692,N_12857);
nand U12926 (N_12926,N_12608,N_12604);
nor U12927 (N_12927,N_12659,N_12609);
nor U12928 (N_12928,N_12786,N_12796);
or U12929 (N_12929,N_12658,N_12684);
or U12930 (N_12930,N_12791,N_12745);
and U12931 (N_12931,N_12650,N_12603);
nor U12932 (N_12932,N_12770,N_12868);
nor U12933 (N_12933,N_12721,N_12663);
nand U12934 (N_12934,N_12827,N_12756);
xor U12935 (N_12935,N_12719,N_12683);
nor U12936 (N_12936,N_12722,N_12673);
or U12937 (N_12937,N_12669,N_12751);
nor U12938 (N_12938,N_12645,N_12704);
nor U12939 (N_12939,N_12666,N_12739);
nand U12940 (N_12940,N_12727,N_12651);
or U12941 (N_12941,N_12633,N_12730);
nand U12942 (N_12942,N_12618,N_12605);
nand U12943 (N_12943,N_12628,N_12816);
and U12944 (N_12944,N_12708,N_12828);
nand U12945 (N_12945,N_12885,N_12610);
and U12946 (N_12946,N_12712,N_12714);
nor U12947 (N_12947,N_12681,N_12846);
xor U12948 (N_12948,N_12776,N_12717);
or U12949 (N_12949,N_12878,N_12619);
nor U12950 (N_12950,N_12626,N_12893);
or U12951 (N_12951,N_12698,N_12640);
nand U12952 (N_12952,N_12840,N_12800);
xnor U12953 (N_12953,N_12735,N_12845);
nand U12954 (N_12954,N_12862,N_12726);
or U12955 (N_12955,N_12895,N_12778);
and U12956 (N_12956,N_12758,N_12880);
nand U12957 (N_12957,N_12799,N_12691);
nand U12958 (N_12958,N_12664,N_12687);
xnor U12959 (N_12959,N_12774,N_12812);
or U12960 (N_12960,N_12869,N_12641);
and U12961 (N_12961,N_12820,N_12855);
nand U12962 (N_12962,N_12762,N_12858);
or U12963 (N_12963,N_12890,N_12823);
nand U12964 (N_12964,N_12793,N_12635);
nand U12965 (N_12965,N_12861,N_12818);
nand U12966 (N_12966,N_12612,N_12740);
nand U12967 (N_12967,N_12821,N_12744);
nand U12968 (N_12968,N_12679,N_12806);
and U12969 (N_12969,N_12864,N_12715);
and U12970 (N_12970,N_12701,N_12777);
nand U12971 (N_12971,N_12634,N_12836);
and U12972 (N_12972,N_12831,N_12662);
or U12973 (N_12973,N_12648,N_12882);
and U12974 (N_12974,N_12667,N_12738);
xor U12975 (N_12975,N_12627,N_12693);
and U12976 (N_12976,N_12709,N_12716);
or U12977 (N_12977,N_12811,N_12607);
xor U12978 (N_12978,N_12775,N_12844);
or U12979 (N_12979,N_12621,N_12875);
nand U12980 (N_12980,N_12674,N_12733);
xnor U12981 (N_12981,N_12736,N_12637);
nand U12982 (N_12982,N_12737,N_12849);
or U12983 (N_12983,N_12631,N_12718);
nand U12984 (N_12984,N_12729,N_12644);
and U12985 (N_12985,N_12647,N_12746);
nand U12986 (N_12986,N_12665,N_12761);
nand U12987 (N_12987,N_12753,N_12884);
nor U12988 (N_12988,N_12657,N_12798);
and U12989 (N_12989,N_12616,N_12760);
nand U12990 (N_12990,N_12731,N_12696);
and U12991 (N_12991,N_12772,N_12668);
nor U12992 (N_12992,N_12764,N_12689);
and U12993 (N_12993,N_12867,N_12747);
or U12994 (N_12994,N_12702,N_12881);
xnor U12995 (N_12995,N_12829,N_12863);
nor U12996 (N_12996,N_12787,N_12725);
or U12997 (N_12997,N_12624,N_12653);
and U12998 (N_12998,N_12865,N_12732);
xnor U12999 (N_12999,N_12707,N_12695);
nand U13000 (N_13000,N_12832,N_12685);
xor U13001 (N_13001,N_12854,N_12757);
or U13002 (N_13002,N_12682,N_12856);
and U13003 (N_13003,N_12842,N_12795);
xnor U13004 (N_13004,N_12851,N_12629);
or U13005 (N_13005,N_12817,N_12754);
nor U13006 (N_13006,N_12809,N_12688);
and U13007 (N_13007,N_12724,N_12660);
nor U13008 (N_13008,N_12656,N_12639);
nand U13009 (N_13009,N_12769,N_12623);
or U13010 (N_13010,N_12887,N_12871);
and U13011 (N_13011,N_12853,N_12617);
nor U13012 (N_13012,N_12843,N_12749);
xor U13013 (N_13013,N_12852,N_12697);
and U13014 (N_13014,N_12723,N_12625);
xnor U13015 (N_13015,N_12675,N_12898);
and U13016 (N_13016,N_12779,N_12742);
nor U13017 (N_13017,N_12835,N_12678);
or U13018 (N_13018,N_12834,N_12706);
or U13019 (N_13019,N_12613,N_12703);
and U13020 (N_13020,N_12720,N_12752);
nand U13021 (N_13021,N_12755,N_12743);
nand U13022 (N_13022,N_12680,N_12789);
xor U13023 (N_13023,N_12838,N_12765);
nor U13024 (N_13024,N_12759,N_12766);
or U13025 (N_13025,N_12797,N_12699);
xor U13026 (N_13026,N_12850,N_12807);
or U13027 (N_13027,N_12677,N_12614);
and U13028 (N_13028,N_12870,N_12655);
xor U13029 (N_13029,N_12801,N_12649);
nor U13030 (N_13030,N_12839,N_12638);
xor U13031 (N_13031,N_12804,N_12790);
or U13032 (N_13032,N_12710,N_12728);
and U13033 (N_13033,N_12825,N_12686);
nor U13034 (N_13034,N_12894,N_12813);
nor U13035 (N_13035,N_12748,N_12891);
xnor U13036 (N_13036,N_12889,N_12892);
xnor U13037 (N_13037,N_12808,N_12620);
xor U13038 (N_13038,N_12690,N_12847);
nand U13039 (N_13039,N_12866,N_12781);
or U13040 (N_13040,N_12694,N_12830);
or U13041 (N_13041,N_12713,N_12642);
nand U13042 (N_13042,N_12837,N_12822);
or U13043 (N_13043,N_12899,N_12883);
xnor U13044 (N_13044,N_12860,N_12792);
nor U13045 (N_13045,N_12711,N_12768);
nand U13046 (N_13046,N_12815,N_12606);
xnor U13047 (N_13047,N_12671,N_12794);
nand U13048 (N_13048,N_12876,N_12654);
nor U13049 (N_13049,N_12782,N_12767);
and U13050 (N_13050,N_12733,N_12861);
nor U13051 (N_13051,N_12687,N_12794);
nor U13052 (N_13052,N_12793,N_12663);
xor U13053 (N_13053,N_12616,N_12882);
or U13054 (N_13054,N_12858,N_12630);
nand U13055 (N_13055,N_12766,N_12714);
nor U13056 (N_13056,N_12871,N_12830);
nor U13057 (N_13057,N_12815,N_12874);
nand U13058 (N_13058,N_12703,N_12774);
xnor U13059 (N_13059,N_12851,N_12713);
and U13060 (N_13060,N_12704,N_12865);
and U13061 (N_13061,N_12794,N_12696);
and U13062 (N_13062,N_12766,N_12797);
or U13063 (N_13063,N_12714,N_12655);
nor U13064 (N_13064,N_12691,N_12668);
nor U13065 (N_13065,N_12823,N_12730);
xor U13066 (N_13066,N_12648,N_12743);
and U13067 (N_13067,N_12893,N_12616);
and U13068 (N_13068,N_12884,N_12803);
nor U13069 (N_13069,N_12741,N_12678);
or U13070 (N_13070,N_12658,N_12601);
or U13071 (N_13071,N_12759,N_12665);
or U13072 (N_13072,N_12773,N_12761);
or U13073 (N_13073,N_12839,N_12832);
nor U13074 (N_13074,N_12819,N_12895);
nor U13075 (N_13075,N_12694,N_12671);
xor U13076 (N_13076,N_12717,N_12873);
xnor U13077 (N_13077,N_12783,N_12643);
xnor U13078 (N_13078,N_12826,N_12642);
and U13079 (N_13079,N_12625,N_12659);
nor U13080 (N_13080,N_12690,N_12794);
nor U13081 (N_13081,N_12809,N_12700);
or U13082 (N_13082,N_12735,N_12726);
and U13083 (N_13083,N_12893,N_12608);
and U13084 (N_13084,N_12677,N_12694);
or U13085 (N_13085,N_12848,N_12821);
nor U13086 (N_13086,N_12777,N_12739);
nor U13087 (N_13087,N_12880,N_12645);
and U13088 (N_13088,N_12819,N_12850);
and U13089 (N_13089,N_12688,N_12703);
xnor U13090 (N_13090,N_12855,N_12818);
and U13091 (N_13091,N_12801,N_12847);
and U13092 (N_13092,N_12805,N_12667);
nor U13093 (N_13093,N_12605,N_12892);
or U13094 (N_13094,N_12857,N_12701);
xnor U13095 (N_13095,N_12658,N_12608);
nor U13096 (N_13096,N_12628,N_12878);
nor U13097 (N_13097,N_12743,N_12671);
and U13098 (N_13098,N_12862,N_12843);
nand U13099 (N_13099,N_12751,N_12666);
or U13100 (N_13100,N_12720,N_12810);
and U13101 (N_13101,N_12823,N_12831);
or U13102 (N_13102,N_12813,N_12733);
xnor U13103 (N_13103,N_12748,N_12839);
and U13104 (N_13104,N_12667,N_12633);
nor U13105 (N_13105,N_12710,N_12862);
nand U13106 (N_13106,N_12869,N_12603);
nand U13107 (N_13107,N_12844,N_12625);
nor U13108 (N_13108,N_12642,N_12699);
or U13109 (N_13109,N_12808,N_12790);
xnor U13110 (N_13110,N_12771,N_12887);
or U13111 (N_13111,N_12605,N_12784);
nand U13112 (N_13112,N_12742,N_12672);
and U13113 (N_13113,N_12618,N_12636);
and U13114 (N_13114,N_12694,N_12643);
or U13115 (N_13115,N_12635,N_12759);
nand U13116 (N_13116,N_12651,N_12808);
and U13117 (N_13117,N_12651,N_12844);
nand U13118 (N_13118,N_12666,N_12759);
xor U13119 (N_13119,N_12764,N_12618);
nand U13120 (N_13120,N_12748,N_12865);
nand U13121 (N_13121,N_12604,N_12639);
xnor U13122 (N_13122,N_12749,N_12764);
xor U13123 (N_13123,N_12835,N_12638);
nor U13124 (N_13124,N_12855,N_12758);
xor U13125 (N_13125,N_12796,N_12888);
nand U13126 (N_13126,N_12856,N_12758);
or U13127 (N_13127,N_12883,N_12881);
nand U13128 (N_13128,N_12756,N_12733);
nor U13129 (N_13129,N_12622,N_12706);
nand U13130 (N_13130,N_12796,N_12619);
xnor U13131 (N_13131,N_12858,N_12712);
nand U13132 (N_13132,N_12609,N_12751);
nand U13133 (N_13133,N_12899,N_12631);
and U13134 (N_13134,N_12766,N_12828);
nand U13135 (N_13135,N_12738,N_12886);
xor U13136 (N_13136,N_12649,N_12740);
nand U13137 (N_13137,N_12790,N_12854);
nand U13138 (N_13138,N_12629,N_12702);
nand U13139 (N_13139,N_12877,N_12839);
nor U13140 (N_13140,N_12653,N_12646);
and U13141 (N_13141,N_12672,N_12673);
and U13142 (N_13142,N_12814,N_12720);
and U13143 (N_13143,N_12699,N_12623);
xor U13144 (N_13144,N_12667,N_12869);
or U13145 (N_13145,N_12743,N_12626);
nor U13146 (N_13146,N_12619,N_12654);
xor U13147 (N_13147,N_12691,N_12612);
or U13148 (N_13148,N_12826,N_12800);
nand U13149 (N_13149,N_12898,N_12700);
and U13150 (N_13150,N_12859,N_12684);
or U13151 (N_13151,N_12839,N_12643);
xnor U13152 (N_13152,N_12727,N_12612);
or U13153 (N_13153,N_12707,N_12754);
or U13154 (N_13154,N_12836,N_12614);
or U13155 (N_13155,N_12860,N_12752);
nand U13156 (N_13156,N_12779,N_12886);
and U13157 (N_13157,N_12713,N_12779);
and U13158 (N_13158,N_12733,N_12677);
nand U13159 (N_13159,N_12705,N_12738);
or U13160 (N_13160,N_12784,N_12730);
nor U13161 (N_13161,N_12883,N_12687);
nand U13162 (N_13162,N_12823,N_12760);
xnor U13163 (N_13163,N_12642,N_12811);
and U13164 (N_13164,N_12641,N_12776);
and U13165 (N_13165,N_12733,N_12759);
xor U13166 (N_13166,N_12863,N_12850);
and U13167 (N_13167,N_12763,N_12741);
xor U13168 (N_13168,N_12657,N_12638);
or U13169 (N_13169,N_12678,N_12608);
nand U13170 (N_13170,N_12665,N_12816);
nand U13171 (N_13171,N_12822,N_12864);
and U13172 (N_13172,N_12629,N_12704);
nor U13173 (N_13173,N_12897,N_12827);
nor U13174 (N_13174,N_12678,N_12899);
or U13175 (N_13175,N_12782,N_12617);
nor U13176 (N_13176,N_12832,N_12890);
xnor U13177 (N_13177,N_12762,N_12655);
nor U13178 (N_13178,N_12866,N_12775);
or U13179 (N_13179,N_12884,N_12821);
nand U13180 (N_13180,N_12782,N_12674);
nand U13181 (N_13181,N_12803,N_12719);
xnor U13182 (N_13182,N_12896,N_12640);
nand U13183 (N_13183,N_12698,N_12631);
nor U13184 (N_13184,N_12719,N_12743);
nand U13185 (N_13185,N_12776,N_12682);
or U13186 (N_13186,N_12795,N_12733);
or U13187 (N_13187,N_12660,N_12889);
and U13188 (N_13188,N_12777,N_12643);
and U13189 (N_13189,N_12702,N_12774);
or U13190 (N_13190,N_12604,N_12724);
or U13191 (N_13191,N_12771,N_12770);
or U13192 (N_13192,N_12804,N_12772);
or U13193 (N_13193,N_12897,N_12766);
and U13194 (N_13194,N_12838,N_12704);
or U13195 (N_13195,N_12780,N_12822);
nand U13196 (N_13196,N_12897,N_12676);
xnor U13197 (N_13197,N_12729,N_12742);
or U13198 (N_13198,N_12660,N_12866);
nand U13199 (N_13199,N_12859,N_12771);
nor U13200 (N_13200,N_13101,N_13151);
nor U13201 (N_13201,N_13108,N_13188);
nand U13202 (N_13202,N_13058,N_12916);
or U13203 (N_13203,N_12958,N_13075);
or U13204 (N_13204,N_13081,N_13087);
nand U13205 (N_13205,N_12967,N_13054);
xnor U13206 (N_13206,N_12939,N_13193);
and U13207 (N_13207,N_13180,N_13120);
nand U13208 (N_13208,N_13156,N_13140);
and U13209 (N_13209,N_13114,N_13071);
nand U13210 (N_13210,N_12953,N_13137);
or U13211 (N_13211,N_13177,N_12941);
and U13212 (N_13212,N_12972,N_13062);
nand U13213 (N_13213,N_13155,N_13021);
or U13214 (N_13214,N_13149,N_13168);
xnor U13215 (N_13215,N_12935,N_13129);
nor U13216 (N_13216,N_13042,N_13162);
nor U13217 (N_13217,N_13097,N_12968);
nand U13218 (N_13218,N_13109,N_13009);
nor U13219 (N_13219,N_13111,N_13152);
xor U13220 (N_13220,N_12982,N_12984);
and U13221 (N_13221,N_13080,N_12976);
xor U13222 (N_13222,N_12998,N_13088);
nand U13223 (N_13223,N_13037,N_13070);
and U13224 (N_13224,N_12912,N_13000);
xor U13225 (N_13225,N_13063,N_13043);
xor U13226 (N_13226,N_13125,N_13192);
nand U13227 (N_13227,N_13079,N_13161);
or U13228 (N_13228,N_13126,N_13026);
xnor U13229 (N_13229,N_13053,N_13154);
nand U13230 (N_13230,N_13064,N_12943);
xor U13231 (N_13231,N_12944,N_13145);
and U13232 (N_13232,N_13046,N_13121);
or U13233 (N_13233,N_12987,N_12963);
nand U13234 (N_13234,N_12901,N_13024);
and U13235 (N_13235,N_13039,N_13056);
nand U13236 (N_13236,N_13065,N_12914);
nor U13237 (N_13237,N_13007,N_12964);
nor U13238 (N_13238,N_13098,N_12911);
and U13239 (N_13239,N_12980,N_13134);
and U13240 (N_13240,N_12937,N_13113);
xnor U13241 (N_13241,N_12918,N_13057);
and U13242 (N_13242,N_12917,N_12971);
nand U13243 (N_13243,N_13086,N_12924);
and U13244 (N_13244,N_13061,N_13072);
nand U13245 (N_13245,N_12981,N_12951);
xnor U13246 (N_13246,N_12952,N_13095);
nand U13247 (N_13247,N_13052,N_13182);
nor U13248 (N_13248,N_12904,N_13181);
nand U13249 (N_13249,N_13132,N_12996);
xnor U13250 (N_13250,N_13138,N_12946);
nor U13251 (N_13251,N_12902,N_13139);
nor U13252 (N_13252,N_13055,N_12932);
nor U13253 (N_13253,N_12908,N_13084);
and U13254 (N_13254,N_12915,N_13127);
and U13255 (N_13255,N_12929,N_13012);
xnor U13256 (N_13256,N_13128,N_13001);
xor U13257 (N_13257,N_12993,N_13136);
nor U13258 (N_13258,N_13195,N_13141);
and U13259 (N_13259,N_12988,N_13189);
nand U13260 (N_13260,N_13069,N_13076);
or U13261 (N_13261,N_13014,N_13144);
and U13262 (N_13262,N_13169,N_12931);
and U13263 (N_13263,N_12942,N_13003);
or U13264 (N_13264,N_13016,N_13199);
nand U13265 (N_13265,N_13194,N_12919);
nor U13266 (N_13266,N_13027,N_13091);
nor U13267 (N_13267,N_12954,N_13019);
xnor U13268 (N_13268,N_13033,N_13025);
nor U13269 (N_13269,N_13167,N_13175);
nor U13270 (N_13270,N_12913,N_12966);
xor U13271 (N_13271,N_13186,N_12957);
xnor U13272 (N_13272,N_12975,N_13160);
and U13273 (N_13273,N_12956,N_12920);
xnor U13274 (N_13274,N_13112,N_13170);
nand U13275 (N_13275,N_13099,N_12970);
xnor U13276 (N_13276,N_12925,N_12969);
xnor U13277 (N_13277,N_13047,N_13038);
and U13278 (N_13278,N_13190,N_12903);
and U13279 (N_13279,N_13198,N_13032);
xnor U13280 (N_13280,N_13174,N_13171);
nor U13281 (N_13281,N_12992,N_12921);
or U13282 (N_13282,N_13028,N_13068);
nor U13283 (N_13283,N_12962,N_13020);
nand U13284 (N_13284,N_13148,N_13173);
or U13285 (N_13285,N_13102,N_13157);
and U13286 (N_13286,N_13050,N_12978);
nand U13287 (N_13287,N_12959,N_12950);
nand U13288 (N_13288,N_12927,N_12905);
nand U13289 (N_13289,N_13124,N_13179);
or U13290 (N_13290,N_12945,N_13094);
and U13291 (N_13291,N_12965,N_13040);
or U13292 (N_13292,N_13092,N_12991);
xnor U13293 (N_13293,N_13130,N_13165);
or U13294 (N_13294,N_13036,N_12989);
xnor U13295 (N_13295,N_12934,N_13060);
and U13296 (N_13296,N_13030,N_13163);
nor U13297 (N_13297,N_13089,N_12985);
nor U13298 (N_13298,N_12990,N_13066);
nand U13299 (N_13299,N_13122,N_13106);
and U13300 (N_13300,N_13133,N_12986);
nor U13301 (N_13301,N_13191,N_12910);
xnor U13302 (N_13302,N_13184,N_12983);
and U13303 (N_13303,N_13143,N_13017);
nor U13304 (N_13304,N_13018,N_13048);
nand U13305 (N_13305,N_12960,N_13006);
nand U13306 (N_13306,N_13115,N_13083);
or U13307 (N_13307,N_12997,N_13185);
nor U13308 (N_13308,N_12955,N_12933);
nand U13309 (N_13309,N_12999,N_12995);
nor U13310 (N_13310,N_13172,N_13078);
and U13311 (N_13311,N_12907,N_12961);
or U13312 (N_13312,N_12922,N_13034);
xor U13313 (N_13313,N_13011,N_13067);
and U13314 (N_13314,N_13022,N_13059);
nand U13315 (N_13315,N_13142,N_13093);
nor U13316 (N_13316,N_13187,N_13176);
xnor U13317 (N_13317,N_13178,N_13082);
xnor U13318 (N_13318,N_13159,N_13041);
nand U13319 (N_13319,N_13104,N_12994);
nor U13320 (N_13320,N_13023,N_13166);
nor U13321 (N_13321,N_13004,N_13131);
and U13322 (N_13322,N_13008,N_13153);
and U13323 (N_13323,N_13045,N_13158);
and U13324 (N_13324,N_13090,N_13015);
xnor U13325 (N_13325,N_12940,N_13005);
nor U13326 (N_13326,N_12906,N_13044);
nor U13327 (N_13327,N_13035,N_13100);
xnor U13328 (N_13328,N_13051,N_13117);
nor U13329 (N_13329,N_13164,N_12923);
and U13330 (N_13330,N_12977,N_13029);
nand U13331 (N_13331,N_13150,N_12949);
or U13332 (N_13332,N_13013,N_13183);
nor U13333 (N_13333,N_13073,N_12928);
and U13334 (N_13334,N_12948,N_12973);
xnor U13335 (N_13335,N_12926,N_13196);
or U13336 (N_13336,N_13118,N_13105);
xor U13337 (N_13337,N_13103,N_13123);
or U13338 (N_13338,N_13146,N_12936);
nand U13339 (N_13339,N_13096,N_12938);
and U13340 (N_13340,N_13135,N_13031);
or U13341 (N_13341,N_13110,N_13197);
nor U13342 (N_13342,N_12979,N_12930);
nor U13343 (N_13343,N_13116,N_13049);
or U13344 (N_13344,N_12900,N_13119);
xor U13345 (N_13345,N_13147,N_13010);
nor U13346 (N_13346,N_13085,N_13002);
and U13347 (N_13347,N_12974,N_13107);
nor U13348 (N_13348,N_13074,N_12947);
xor U13349 (N_13349,N_12909,N_13077);
nand U13350 (N_13350,N_13189,N_13158);
nor U13351 (N_13351,N_13178,N_12956);
and U13352 (N_13352,N_12929,N_13132);
and U13353 (N_13353,N_12964,N_12992);
xor U13354 (N_13354,N_12973,N_12993);
or U13355 (N_13355,N_13011,N_12976);
nor U13356 (N_13356,N_13001,N_12929);
nand U13357 (N_13357,N_13181,N_13146);
xor U13358 (N_13358,N_13010,N_13099);
and U13359 (N_13359,N_12967,N_13165);
xnor U13360 (N_13360,N_12987,N_13196);
nand U13361 (N_13361,N_13162,N_13174);
nand U13362 (N_13362,N_13196,N_13082);
and U13363 (N_13363,N_12975,N_13043);
xnor U13364 (N_13364,N_13094,N_13100);
or U13365 (N_13365,N_13057,N_13020);
or U13366 (N_13366,N_13148,N_12969);
xor U13367 (N_13367,N_12981,N_12984);
or U13368 (N_13368,N_12928,N_12948);
nand U13369 (N_13369,N_13010,N_12997);
and U13370 (N_13370,N_13174,N_13113);
or U13371 (N_13371,N_13038,N_12950);
or U13372 (N_13372,N_13034,N_12960);
xor U13373 (N_13373,N_12974,N_13069);
and U13374 (N_13374,N_13012,N_12926);
xor U13375 (N_13375,N_13162,N_13100);
xor U13376 (N_13376,N_12998,N_13071);
nor U13377 (N_13377,N_12908,N_13026);
xnor U13378 (N_13378,N_13172,N_13012);
nand U13379 (N_13379,N_13193,N_12997);
or U13380 (N_13380,N_13129,N_12951);
and U13381 (N_13381,N_13015,N_13102);
or U13382 (N_13382,N_12947,N_13195);
nand U13383 (N_13383,N_13085,N_12929);
nor U13384 (N_13384,N_13168,N_12954);
nor U13385 (N_13385,N_13098,N_13173);
nor U13386 (N_13386,N_12940,N_12936);
or U13387 (N_13387,N_12928,N_12953);
nand U13388 (N_13388,N_13088,N_12910);
and U13389 (N_13389,N_13040,N_13060);
or U13390 (N_13390,N_13114,N_12999);
nor U13391 (N_13391,N_12958,N_13087);
nand U13392 (N_13392,N_12972,N_12954);
and U13393 (N_13393,N_13091,N_13097);
nor U13394 (N_13394,N_13133,N_12940);
or U13395 (N_13395,N_12941,N_13179);
nor U13396 (N_13396,N_12932,N_12980);
and U13397 (N_13397,N_12900,N_13083);
or U13398 (N_13398,N_12908,N_13059);
and U13399 (N_13399,N_12969,N_13000);
xnor U13400 (N_13400,N_13023,N_12918);
nor U13401 (N_13401,N_12969,N_12983);
nand U13402 (N_13402,N_13162,N_13023);
and U13403 (N_13403,N_12979,N_13028);
or U13404 (N_13404,N_13091,N_12946);
and U13405 (N_13405,N_12953,N_13089);
nand U13406 (N_13406,N_12910,N_12988);
nand U13407 (N_13407,N_12945,N_12966);
or U13408 (N_13408,N_13076,N_13193);
and U13409 (N_13409,N_13089,N_12937);
xor U13410 (N_13410,N_13111,N_12972);
nand U13411 (N_13411,N_12916,N_13030);
nor U13412 (N_13412,N_12912,N_12931);
nand U13413 (N_13413,N_12955,N_13056);
xnor U13414 (N_13414,N_12937,N_13116);
or U13415 (N_13415,N_12984,N_12932);
nor U13416 (N_13416,N_13137,N_13183);
nor U13417 (N_13417,N_12912,N_12929);
nand U13418 (N_13418,N_13057,N_12936);
or U13419 (N_13419,N_13052,N_13069);
nand U13420 (N_13420,N_13199,N_12926);
and U13421 (N_13421,N_13019,N_12974);
nand U13422 (N_13422,N_13174,N_12920);
nor U13423 (N_13423,N_13163,N_13175);
xnor U13424 (N_13424,N_13043,N_12913);
or U13425 (N_13425,N_12900,N_12913);
and U13426 (N_13426,N_13043,N_13168);
and U13427 (N_13427,N_13186,N_13166);
or U13428 (N_13428,N_12996,N_13172);
and U13429 (N_13429,N_12915,N_13076);
xnor U13430 (N_13430,N_13122,N_13012);
nand U13431 (N_13431,N_12938,N_13172);
nor U13432 (N_13432,N_13059,N_12936);
and U13433 (N_13433,N_13166,N_13005);
nor U13434 (N_13434,N_12960,N_12967);
and U13435 (N_13435,N_13190,N_13193);
xnor U13436 (N_13436,N_13196,N_12930);
or U13437 (N_13437,N_12976,N_13070);
nand U13438 (N_13438,N_13077,N_13189);
xnor U13439 (N_13439,N_13040,N_13161);
and U13440 (N_13440,N_13066,N_12980);
xnor U13441 (N_13441,N_13007,N_13123);
nand U13442 (N_13442,N_13104,N_13192);
nor U13443 (N_13443,N_13076,N_13191);
nand U13444 (N_13444,N_13131,N_12945);
nor U13445 (N_13445,N_13088,N_13187);
xor U13446 (N_13446,N_13049,N_13191);
nor U13447 (N_13447,N_12916,N_13088);
xnor U13448 (N_13448,N_13041,N_12992);
or U13449 (N_13449,N_12983,N_13014);
and U13450 (N_13450,N_13177,N_13054);
xor U13451 (N_13451,N_13015,N_13160);
or U13452 (N_13452,N_13159,N_13063);
nor U13453 (N_13453,N_13012,N_12909);
or U13454 (N_13454,N_12970,N_12950);
and U13455 (N_13455,N_13013,N_12968);
and U13456 (N_13456,N_13037,N_12944);
nand U13457 (N_13457,N_12957,N_12960);
xnor U13458 (N_13458,N_13139,N_13187);
xnor U13459 (N_13459,N_13040,N_13150);
and U13460 (N_13460,N_13139,N_12981);
nor U13461 (N_13461,N_13006,N_13008);
and U13462 (N_13462,N_12960,N_13126);
nand U13463 (N_13463,N_13088,N_13120);
nand U13464 (N_13464,N_13197,N_13191);
nand U13465 (N_13465,N_12928,N_13011);
and U13466 (N_13466,N_13129,N_13069);
nor U13467 (N_13467,N_13065,N_13024);
nor U13468 (N_13468,N_13030,N_13072);
and U13469 (N_13469,N_13126,N_13087);
or U13470 (N_13470,N_13081,N_13039);
xnor U13471 (N_13471,N_13111,N_13092);
and U13472 (N_13472,N_13054,N_12937);
or U13473 (N_13473,N_13084,N_13153);
xnor U13474 (N_13474,N_13176,N_12955);
nor U13475 (N_13475,N_13044,N_13035);
nor U13476 (N_13476,N_13137,N_13120);
and U13477 (N_13477,N_13142,N_13165);
and U13478 (N_13478,N_12936,N_13051);
nand U13479 (N_13479,N_13141,N_13094);
and U13480 (N_13480,N_13153,N_13131);
nand U13481 (N_13481,N_13092,N_13110);
and U13482 (N_13482,N_13173,N_13101);
nand U13483 (N_13483,N_12923,N_12958);
nand U13484 (N_13484,N_13183,N_13023);
nor U13485 (N_13485,N_13095,N_13056);
xnor U13486 (N_13486,N_13162,N_13028);
nor U13487 (N_13487,N_13123,N_13140);
nand U13488 (N_13488,N_12970,N_13056);
nor U13489 (N_13489,N_13071,N_12938);
nor U13490 (N_13490,N_13172,N_13183);
or U13491 (N_13491,N_12900,N_13126);
or U13492 (N_13492,N_13184,N_12998);
xor U13493 (N_13493,N_12943,N_13136);
or U13494 (N_13494,N_13184,N_13053);
nor U13495 (N_13495,N_12964,N_13076);
and U13496 (N_13496,N_12981,N_13064);
nand U13497 (N_13497,N_13187,N_13168);
and U13498 (N_13498,N_13198,N_12980);
and U13499 (N_13499,N_13104,N_12948);
nor U13500 (N_13500,N_13203,N_13208);
nand U13501 (N_13501,N_13479,N_13426);
or U13502 (N_13502,N_13465,N_13259);
and U13503 (N_13503,N_13497,N_13382);
nand U13504 (N_13504,N_13467,N_13248);
nor U13505 (N_13505,N_13430,N_13268);
and U13506 (N_13506,N_13357,N_13267);
nand U13507 (N_13507,N_13481,N_13308);
or U13508 (N_13508,N_13253,N_13491);
and U13509 (N_13509,N_13238,N_13391);
nor U13510 (N_13510,N_13461,N_13339);
and U13511 (N_13511,N_13223,N_13243);
nor U13512 (N_13512,N_13250,N_13459);
xnor U13513 (N_13513,N_13252,N_13387);
xnor U13514 (N_13514,N_13201,N_13494);
nor U13515 (N_13515,N_13424,N_13485);
xor U13516 (N_13516,N_13451,N_13273);
nor U13517 (N_13517,N_13334,N_13269);
and U13518 (N_13518,N_13327,N_13393);
xor U13519 (N_13519,N_13346,N_13431);
or U13520 (N_13520,N_13255,N_13421);
nand U13521 (N_13521,N_13363,N_13296);
nor U13522 (N_13522,N_13263,N_13496);
and U13523 (N_13523,N_13349,N_13412);
or U13524 (N_13524,N_13394,N_13256);
nand U13525 (N_13525,N_13290,N_13202);
or U13526 (N_13526,N_13457,N_13348);
and U13527 (N_13527,N_13381,N_13482);
nor U13528 (N_13528,N_13345,N_13462);
nor U13529 (N_13529,N_13383,N_13280);
nand U13530 (N_13530,N_13315,N_13251);
xnor U13531 (N_13531,N_13298,N_13266);
nor U13532 (N_13532,N_13427,N_13309);
or U13533 (N_13533,N_13450,N_13226);
nor U13534 (N_13534,N_13447,N_13405);
or U13535 (N_13535,N_13257,N_13399);
and U13536 (N_13536,N_13472,N_13215);
or U13537 (N_13537,N_13370,N_13411);
nand U13538 (N_13538,N_13406,N_13305);
nor U13539 (N_13539,N_13204,N_13262);
nand U13540 (N_13540,N_13486,N_13460);
nand U13541 (N_13541,N_13232,N_13355);
nand U13542 (N_13542,N_13474,N_13483);
xor U13543 (N_13543,N_13241,N_13404);
xor U13544 (N_13544,N_13294,N_13407);
or U13545 (N_13545,N_13249,N_13436);
and U13546 (N_13546,N_13480,N_13373);
or U13547 (N_13547,N_13410,N_13335);
or U13548 (N_13548,N_13378,N_13418);
nand U13549 (N_13549,N_13493,N_13217);
nor U13550 (N_13550,N_13282,N_13338);
nor U13551 (N_13551,N_13293,N_13275);
nor U13552 (N_13552,N_13288,N_13299);
or U13553 (N_13553,N_13400,N_13376);
nand U13554 (N_13554,N_13236,N_13358);
xnor U13555 (N_13555,N_13209,N_13316);
or U13556 (N_13556,N_13352,N_13274);
nor U13557 (N_13557,N_13289,N_13435);
xor U13558 (N_13558,N_13401,N_13452);
nor U13559 (N_13559,N_13396,N_13216);
xnor U13560 (N_13560,N_13318,N_13415);
xnor U13561 (N_13561,N_13303,N_13395);
nand U13562 (N_13562,N_13377,N_13281);
nor U13563 (N_13563,N_13423,N_13375);
and U13564 (N_13564,N_13212,N_13227);
and U13565 (N_13565,N_13337,N_13242);
xnor U13566 (N_13566,N_13384,N_13302);
and U13567 (N_13567,N_13287,N_13247);
xor U13568 (N_13568,N_13361,N_13330);
and U13569 (N_13569,N_13283,N_13463);
nand U13570 (N_13570,N_13278,N_13475);
nor U13571 (N_13571,N_13385,N_13398);
or U13572 (N_13572,N_13229,N_13230);
or U13573 (N_13573,N_13487,N_13350);
nor U13574 (N_13574,N_13228,N_13225);
and U13575 (N_13575,N_13333,N_13219);
nor U13576 (N_13576,N_13409,N_13368);
nand U13577 (N_13577,N_13379,N_13408);
xnor U13578 (N_13578,N_13231,N_13336);
nor U13579 (N_13579,N_13419,N_13369);
or U13580 (N_13580,N_13328,N_13469);
and U13581 (N_13581,N_13366,N_13271);
nor U13582 (N_13582,N_13359,N_13218);
xor U13583 (N_13583,N_13222,N_13240);
and U13584 (N_13584,N_13246,N_13417);
nor U13585 (N_13585,N_13207,N_13331);
nor U13586 (N_13586,N_13295,N_13468);
or U13587 (N_13587,N_13392,N_13453);
nand U13588 (N_13588,N_13413,N_13470);
xnor U13589 (N_13589,N_13433,N_13341);
or U13590 (N_13590,N_13322,N_13258);
nor U13591 (N_13591,N_13478,N_13428);
nand U13592 (N_13592,N_13239,N_13319);
or U13593 (N_13593,N_13477,N_13220);
nand U13594 (N_13594,N_13464,N_13362);
nor U13595 (N_13595,N_13441,N_13351);
or U13596 (N_13596,N_13440,N_13321);
nor U13597 (N_13597,N_13402,N_13371);
or U13598 (N_13598,N_13313,N_13432);
and U13599 (N_13599,N_13458,N_13429);
and U13600 (N_13600,N_13320,N_13342);
or U13601 (N_13601,N_13297,N_13476);
nand U13602 (N_13602,N_13221,N_13306);
xor U13603 (N_13603,N_13437,N_13442);
nor U13604 (N_13604,N_13224,N_13364);
nor U13605 (N_13605,N_13438,N_13210);
or U13606 (N_13606,N_13492,N_13353);
nor U13607 (N_13607,N_13264,N_13200);
nor U13608 (N_13608,N_13340,N_13332);
and U13609 (N_13609,N_13272,N_13260);
xnor U13610 (N_13610,N_13284,N_13397);
nand U13611 (N_13611,N_13360,N_13205);
or U13612 (N_13612,N_13254,N_13498);
nand U13613 (N_13613,N_13445,N_13214);
nand U13614 (N_13614,N_13310,N_13244);
nand U13615 (N_13615,N_13265,N_13444);
and U13616 (N_13616,N_13455,N_13312);
nand U13617 (N_13617,N_13311,N_13390);
and U13618 (N_13618,N_13211,N_13206);
nor U13619 (N_13619,N_13279,N_13443);
xnor U13620 (N_13620,N_13324,N_13372);
nand U13621 (N_13621,N_13454,N_13490);
nand U13622 (N_13622,N_13285,N_13488);
or U13623 (N_13623,N_13344,N_13300);
nor U13624 (N_13624,N_13425,N_13473);
nand U13625 (N_13625,N_13489,N_13434);
and U13626 (N_13626,N_13386,N_13403);
nand U13627 (N_13627,N_13276,N_13374);
and U13628 (N_13628,N_13261,N_13292);
or U13629 (N_13629,N_13446,N_13495);
or U13630 (N_13630,N_13439,N_13354);
nor U13631 (N_13631,N_13323,N_13286);
xnor U13632 (N_13632,N_13301,N_13456);
nor U13633 (N_13633,N_13314,N_13389);
or U13634 (N_13634,N_13471,N_13420);
nand U13635 (N_13635,N_13235,N_13270);
or U13636 (N_13636,N_13277,N_13449);
nor U13637 (N_13637,N_13448,N_13245);
nor U13638 (N_13638,N_13347,N_13237);
and U13639 (N_13639,N_13380,N_13291);
and U13640 (N_13640,N_13213,N_13416);
nor U13641 (N_13641,N_13365,N_13484);
nor U13642 (N_13642,N_13307,N_13414);
xor U13643 (N_13643,N_13422,N_13388);
nor U13644 (N_13644,N_13367,N_13466);
nand U13645 (N_13645,N_13499,N_13304);
nand U13646 (N_13646,N_13356,N_13317);
nand U13647 (N_13647,N_13343,N_13329);
nand U13648 (N_13648,N_13234,N_13233);
or U13649 (N_13649,N_13326,N_13325);
or U13650 (N_13650,N_13277,N_13382);
xor U13651 (N_13651,N_13444,N_13432);
and U13652 (N_13652,N_13453,N_13439);
xnor U13653 (N_13653,N_13250,N_13315);
xor U13654 (N_13654,N_13458,N_13393);
xnor U13655 (N_13655,N_13303,N_13225);
nor U13656 (N_13656,N_13286,N_13454);
or U13657 (N_13657,N_13469,N_13339);
nand U13658 (N_13658,N_13441,N_13206);
or U13659 (N_13659,N_13389,N_13370);
nand U13660 (N_13660,N_13276,N_13388);
nand U13661 (N_13661,N_13330,N_13251);
nor U13662 (N_13662,N_13223,N_13230);
or U13663 (N_13663,N_13410,N_13255);
nor U13664 (N_13664,N_13488,N_13399);
xnor U13665 (N_13665,N_13312,N_13266);
or U13666 (N_13666,N_13260,N_13429);
xor U13667 (N_13667,N_13438,N_13333);
xnor U13668 (N_13668,N_13280,N_13412);
nand U13669 (N_13669,N_13289,N_13434);
or U13670 (N_13670,N_13427,N_13462);
and U13671 (N_13671,N_13355,N_13215);
nand U13672 (N_13672,N_13373,N_13315);
nor U13673 (N_13673,N_13323,N_13265);
xnor U13674 (N_13674,N_13425,N_13354);
nor U13675 (N_13675,N_13422,N_13259);
nand U13676 (N_13676,N_13443,N_13232);
xor U13677 (N_13677,N_13482,N_13298);
nand U13678 (N_13678,N_13291,N_13384);
xnor U13679 (N_13679,N_13223,N_13368);
nor U13680 (N_13680,N_13453,N_13231);
and U13681 (N_13681,N_13315,N_13403);
nor U13682 (N_13682,N_13205,N_13459);
nand U13683 (N_13683,N_13493,N_13342);
and U13684 (N_13684,N_13421,N_13248);
or U13685 (N_13685,N_13417,N_13229);
and U13686 (N_13686,N_13487,N_13333);
and U13687 (N_13687,N_13394,N_13359);
and U13688 (N_13688,N_13262,N_13382);
nor U13689 (N_13689,N_13358,N_13256);
nand U13690 (N_13690,N_13479,N_13464);
or U13691 (N_13691,N_13315,N_13419);
and U13692 (N_13692,N_13471,N_13418);
and U13693 (N_13693,N_13492,N_13343);
or U13694 (N_13694,N_13410,N_13302);
or U13695 (N_13695,N_13401,N_13206);
or U13696 (N_13696,N_13277,N_13388);
or U13697 (N_13697,N_13385,N_13380);
and U13698 (N_13698,N_13233,N_13385);
xnor U13699 (N_13699,N_13218,N_13341);
or U13700 (N_13700,N_13310,N_13355);
xor U13701 (N_13701,N_13232,N_13398);
or U13702 (N_13702,N_13405,N_13310);
nor U13703 (N_13703,N_13321,N_13450);
xnor U13704 (N_13704,N_13396,N_13289);
and U13705 (N_13705,N_13451,N_13239);
or U13706 (N_13706,N_13309,N_13362);
xor U13707 (N_13707,N_13494,N_13303);
nor U13708 (N_13708,N_13200,N_13327);
nor U13709 (N_13709,N_13256,N_13474);
nor U13710 (N_13710,N_13398,N_13476);
xnor U13711 (N_13711,N_13290,N_13409);
or U13712 (N_13712,N_13403,N_13357);
or U13713 (N_13713,N_13357,N_13313);
xor U13714 (N_13714,N_13495,N_13308);
or U13715 (N_13715,N_13445,N_13460);
nand U13716 (N_13716,N_13363,N_13306);
nand U13717 (N_13717,N_13414,N_13332);
or U13718 (N_13718,N_13451,N_13241);
nand U13719 (N_13719,N_13427,N_13340);
nor U13720 (N_13720,N_13364,N_13350);
and U13721 (N_13721,N_13362,N_13487);
nand U13722 (N_13722,N_13248,N_13269);
xnor U13723 (N_13723,N_13300,N_13436);
or U13724 (N_13724,N_13281,N_13317);
and U13725 (N_13725,N_13356,N_13446);
or U13726 (N_13726,N_13497,N_13329);
xor U13727 (N_13727,N_13349,N_13497);
xor U13728 (N_13728,N_13409,N_13474);
and U13729 (N_13729,N_13301,N_13352);
xnor U13730 (N_13730,N_13461,N_13311);
and U13731 (N_13731,N_13346,N_13232);
xnor U13732 (N_13732,N_13477,N_13261);
nand U13733 (N_13733,N_13452,N_13474);
nand U13734 (N_13734,N_13217,N_13366);
nand U13735 (N_13735,N_13227,N_13248);
nor U13736 (N_13736,N_13499,N_13443);
xnor U13737 (N_13737,N_13224,N_13480);
nand U13738 (N_13738,N_13437,N_13292);
nor U13739 (N_13739,N_13389,N_13458);
nand U13740 (N_13740,N_13239,N_13473);
nand U13741 (N_13741,N_13208,N_13492);
nor U13742 (N_13742,N_13433,N_13211);
or U13743 (N_13743,N_13289,N_13319);
nor U13744 (N_13744,N_13397,N_13466);
and U13745 (N_13745,N_13201,N_13473);
xnor U13746 (N_13746,N_13279,N_13326);
xor U13747 (N_13747,N_13447,N_13311);
and U13748 (N_13748,N_13276,N_13433);
and U13749 (N_13749,N_13424,N_13397);
or U13750 (N_13750,N_13259,N_13444);
xnor U13751 (N_13751,N_13298,N_13317);
nor U13752 (N_13752,N_13459,N_13273);
or U13753 (N_13753,N_13472,N_13265);
and U13754 (N_13754,N_13238,N_13343);
or U13755 (N_13755,N_13436,N_13220);
nand U13756 (N_13756,N_13409,N_13308);
nand U13757 (N_13757,N_13260,N_13385);
and U13758 (N_13758,N_13413,N_13311);
or U13759 (N_13759,N_13228,N_13310);
or U13760 (N_13760,N_13346,N_13220);
nor U13761 (N_13761,N_13342,N_13354);
nand U13762 (N_13762,N_13371,N_13293);
and U13763 (N_13763,N_13454,N_13483);
or U13764 (N_13764,N_13277,N_13377);
nand U13765 (N_13765,N_13323,N_13426);
nand U13766 (N_13766,N_13270,N_13339);
and U13767 (N_13767,N_13205,N_13294);
or U13768 (N_13768,N_13222,N_13425);
xor U13769 (N_13769,N_13301,N_13306);
nor U13770 (N_13770,N_13309,N_13286);
nand U13771 (N_13771,N_13365,N_13322);
nand U13772 (N_13772,N_13387,N_13326);
and U13773 (N_13773,N_13498,N_13385);
xnor U13774 (N_13774,N_13252,N_13207);
nand U13775 (N_13775,N_13374,N_13247);
or U13776 (N_13776,N_13433,N_13238);
and U13777 (N_13777,N_13376,N_13451);
nor U13778 (N_13778,N_13247,N_13219);
nand U13779 (N_13779,N_13360,N_13444);
or U13780 (N_13780,N_13367,N_13291);
or U13781 (N_13781,N_13311,N_13385);
nand U13782 (N_13782,N_13312,N_13264);
nand U13783 (N_13783,N_13244,N_13333);
and U13784 (N_13784,N_13336,N_13252);
nor U13785 (N_13785,N_13481,N_13375);
nand U13786 (N_13786,N_13460,N_13305);
nor U13787 (N_13787,N_13266,N_13378);
nand U13788 (N_13788,N_13428,N_13331);
or U13789 (N_13789,N_13280,N_13369);
nor U13790 (N_13790,N_13364,N_13218);
and U13791 (N_13791,N_13421,N_13308);
and U13792 (N_13792,N_13451,N_13482);
and U13793 (N_13793,N_13232,N_13370);
and U13794 (N_13794,N_13391,N_13233);
or U13795 (N_13795,N_13439,N_13425);
nand U13796 (N_13796,N_13439,N_13352);
and U13797 (N_13797,N_13217,N_13439);
and U13798 (N_13798,N_13295,N_13331);
and U13799 (N_13799,N_13311,N_13307);
and U13800 (N_13800,N_13642,N_13780);
nor U13801 (N_13801,N_13613,N_13718);
and U13802 (N_13802,N_13592,N_13625);
and U13803 (N_13803,N_13571,N_13644);
nand U13804 (N_13804,N_13566,N_13527);
nand U13805 (N_13805,N_13702,N_13688);
or U13806 (N_13806,N_13725,N_13523);
or U13807 (N_13807,N_13616,N_13786);
or U13808 (N_13808,N_13620,N_13710);
and U13809 (N_13809,N_13678,N_13656);
nor U13810 (N_13810,N_13788,N_13514);
xor U13811 (N_13811,N_13617,N_13673);
or U13812 (N_13812,N_13659,N_13636);
or U13813 (N_13813,N_13793,N_13658);
xor U13814 (N_13814,N_13648,N_13693);
or U13815 (N_13815,N_13502,N_13776);
and U13816 (N_13816,N_13696,N_13739);
xnor U13817 (N_13817,N_13735,N_13761);
nand U13818 (N_13818,N_13500,N_13698);
and U13819 (N_13819,N_13524,N_13533);
nand U13820 (N_13820,N_13717,N_13639);
xnor U13821 (N_13821,N_13614,N_13537);
xor U13822 (N_13822,N_13757,N_13713);
xor U13823 (N_13823,N_13703,N_13584);
and U13824 (N_13824,N_13743,N_13591);
xnor U13825 (N_13825,N_13756,N_13640);
nor U13826 (N_13826,N_13564,N_13545);
or U13827 (N_13827,N_13677,N_13586);
nand U13828 (N_13828,N_13770,N_13531);
or U13829 (N_13829,N_13661,N_13641);
or U13830 (N_13830,N_13745,N_13554);
and U13831 (N_13831,N_13727,N_13645);
nor U13832 (N_13832,N_13730,N_13529);
nand U13833 (N_13833,N_13519,N_13646);
and U13834 (N_13834,N_13582,N_13777);
nor U13835 (N_13835,N_13653,N_13647);
nand U13836 (N_13836,N_13790,N_13627);
or U13837 (N_13837,N_13667,N_13716);
xor U13838 (N_13838,N_13722,N_13797);
nand U13839 (N_13839,N_13555,N_13635);
or U13840 (N_13840,N_13581,N_13556);
and U13841 (N_13841,N_13601,N_13608);
and U13842 (N_13842,N_13738,N_13746);
or U13843 (N_13843,N_13798,N_13781);
and U13844 (N_13844,N_13740,N_13633);
xnor U13845 (N_13845,N_13573,N_13593);
xor U13846 (N_13846,N_13785,N_13512);
and U13847 (N_13847,N_13694,N_13546);
and U13848 (N_13848,N_13682,N_13750);
nor U13849 (N_13849,N_13669,N_13691);
xnor U13850 (N_13850,N_13692,N_13587);
nor U13851 (N_13851,N_13557,N_13513);
nor U13852 (N_13852,N_13578,N_13734);
nand U13853 (N_13853,N_13528,N_13675);
nor U13854 (N_13854,N_13526,N_13530);
nand U13855 (N_13855,N_13649,N_13615);
nor U13856 (N_13856,N_13731,N_13629);
xnor U13857 (N_13857,N_13577,N_13637);
and U13858 (N_13858,N_13631,N_13762);
nand U13859 (N_13859,N_13552,N_13704);
nand U13860 (N_13860,N_13729,N_13736);
and U13861 (N_13861,N_13670,N_13672);
nand U13862 (N_13862,N_13569,N_13604);
and U13863 (N_13863,N_13789,N_13664);
nor U13864 (N_13864,N_13742,N_13791);
or U13865 (N_13865,N_13792,N_13699);
and U13866 (N_13866,N_13598,N_13737);
nor U13867 (N_13867,N_13549,N_13697);
and U13868 (N_13868,N_13663,N_13630);
nor U13869 (N_13869,N_13723,N_13575);
nand U13870 (N_13870,N_13726,N_13687);
and U13871 (N_13871,N_13732,N_13706);
and U13872 (N_13872,N_13755,N_13719);
and U13873 (N_13873,N_13607,N_13685);
and U13874 (N_13874,N_13612,N_13525);
xor U13875 (N_13875,N_13503,N_13515);
or U13876 (N_13876,N_13572,N_13510);
or U13877 (N_13877,N_13563,N_13749);
or U13878 (N_13878,N_13516,N_13606);
nor U13879 (N_13879,N_13695,N_13517);
nand U13880 (N_13880,N_13632,N_13748);
nand U13881 (N_13881,N_13643,N_13654);
and U13882 (N_13882,N_13650,N_13754);
and U13883 (N_13883,N_13522,N_13574);
and U13884 (N_13884,N_13568,N_13520);
xnor U13885 (N_13885,N_13767,N_13634);
xnor U13886 (N_13886,N_13760,N_13714);
nand U13887 (N_13887,N_13747,N_13709);
and U13888 (N_13888,N_13580,N_13759);
xnor U13889 (N_13889,N_13599,N_13768);
nand U13890 (N_13890,N_13787,N_13624);
or U13891 (N_13891,N_13518,N_13751);
or U13892 (N_13892,N_13565,N_13765);
xor U13893 (N_13893,N_13603,N_13595);
and U13894 (N_13894,N_13596,N_13600);
and U13895 (N_13895,N_13626,N_13521);
nor U13896 (N_13896,N_13506,N_13609);
xor U13897 (N_13897,N_13623,N_13576);
and U13898 (N_13898,N_13553,N_13652);
nor U13899 (N_13899,N_13701,N_13544);
nor U13900 (N_13900,N_13618,N_13651);
or U13901 (N_13901,N_13619,N_13542);
or U13902 (N_13902,N_13504,N_13779);
xor U13903 (N_13903,N_13753,N_13708);
nor U13904 (N_13904,N_13684,N_13715);
nand U13905 (N_13905,N_13610,N_13508);
and U13906 (N_13906,N_13501,N_13579);
and U13907 (N_13907,N_13782,N_13605);
xor U13908 (N_13908,N_13666,N_13772);
and U13909 (N_13909,N_13611,N_13562);
xnor U13910 (N_13910,N_13712,N_13536);
or U13911 (N_13911,N_13662,N_13622);
nand U13912 (N_13912,N_13590,N_13671);
nand U13913 (N_13913,N_13548,N_13741);
nand U13914 (N_13914,N_13680,N_13763);
xnor U13915 (N_13915,N_13588,N_13766);
or U13916 (N_13916,N_13660,N_13541);
xor U13917 (N_13917,N_13561,N_13668);
or U13918 (N_13918,N_13543,N_13665);
or U13919 (N_13919,N_13674,N_13724);
nor U13920 (N_13920,N_13681,N_13796);
xor U13921 (N_13921,N_13764,N_13778);
and U13922 (N_13922,N_13507,N_13540);
nor U13923 (N_13923,N_13558,N_13784);
nand U13924 (N_13924,N_13733,N_13655);
or U13925 (N_13925,N_13721,N_13567);
nand U13926 (N_13926,N_13621,N_13657);
and U13927 (N_13927,N_13511,N_13795);
xor U13928 (N_13928,N_13769,N_13690);
and U13929 (N_13929,N_13705,N_13585);
and U13930 (N_13930,N_13771,N_13683);
nand U13931 (N_13931,N_13676,N_13686);
or U13932 (N_13932,N_13551,N_13535);
xnor U13933 (N_13933,N_13794,N_13744);
and U13934 (N_13934,N_13597,N_13638);
or U13935 (N_13935,N_13758,N_13752);
xor U13936 (N_13936,N_13720,N_13711);
xnor U13937 (N_13937,N_13570,N_13547);
or U13938 (N_13938,N_13728,N_13594);
nor U13939 (N_13939,N_13509,N_13628);
nand U13940 (N_13940,N_13538,N_13532);
or U13941 (N_13941,N_13775,N_13774);
or U13942 (N_13942,N_13679,N_13773);
nor U13943 (N_13943,N_13689,N_13602);
nand U13944 (N_13944,N_13505,N_13707);
nor U13945 (N_13945,N_13534,N_13700);
or U13946 (N_13946,N_13799,N_13550);
nand U13947 (N_13947,N_13539,N_13583);
xnor U13948 (N_13948,N_13560,N_13589);
nand U13949 (N_13949,N_13783,N_13559);
xor U13950 (N_13950,N_13604,N_13539);
nor U13951 (N_13951,N_13760,N_13609);
xor U13952 (N_13952,N_13771,N_13555);
or U13953 (N_13953,N_13698,N_13503);
nand U13954 (N_13954,N_13506,N_13719);
or U13955 (N_13955,N_13505,N_13701);
or U13956 (N_13956,N_13680,N_13691);
nand U13957 (N_13957,N_13621,N_13675);
nor U13958 (N_13958,N_13601,N_13747);
and U13959 (N_13959,N_13681,N_13534);
and U13960 (N_13960,N_13567,N_13577);
xnor U13961 (N_13961,N_13664,N_13756);
and U13962 (N_13962,N_13592,N_13508);
or U13963 (N_13963,N_13796,N_13634);
and U13964 (N_13964,N_13760,N_13615);
or U13965 (N_13965,N_13699,N_13621);
or U13966 (N_13966,N_13672,N_13604);
nor U13967 (N_13967,N_13778,N_13741);
nand U13968 (N_13968,N_13749,N_13776);
and U13969 (N_13969,N_13734,N_13768);
nand U13970 (N_13970,N_13559,N_13681);
nor U13971 (N_13971,N_13614,N_13755);
xor U13972 (N_13972,N_13620,N_13657);
nor U13973 (N_13973,N_13661,N_13757);
or U13974 (N_13974,N_13525,N_13750);
and U13975 (N_13975,N_13717,N_13749);
nand U13976 (N_13976,N_13547,N_13744);
xnor U13977 (N_13977,N_13677,N_13595);
or U13978 (N_13978,N_13678,N_13747);
nor U13979 (N_13979,N_13575,N_13664);
and U13980 (N_13980,N_13519,N_13627);
nor U13981 (N_13981,N_13729,N_13711);
and U13982 (N_13982,N_13793,N_13539);
and U13983 (N_13983,N_13732,N_13720);
nor U13984 (N_13984,N_13751,N_13575);
and U13985 (N_13985,N_13566,N_13632);
xor U13986 (N_13986,N_13654,N_13757);
nor U13987 (N_13987,N_13797,N_13680);
nand U13988 (N_13988,N_13708,N_13653);
nand U13989 (N_13989,N_13625,N_13666);
xnor U13990 (N_13990,N_13537,N_13609);
and U13991 (N_13991,N_13542,N_13724);
or U13992 (N_13992,N_13501,N_13778);
xnor U13993 (N_13993,N_13500,N_13594);
or U13994 (N_13994,N_13542,N_13762);
nor U13995 (N_13995,N_13794,N_13688);
xnor U13996 (N_13996,N_13708,N_13764);
nand U13997 (N_13997,N_13741,N_13629);
nand U13998 (N_13998,N_13770,N_13580);
nor U13999 (N_13999,N_13605,N_13671);
xor U14000 (N_14000,N_13684,N_13594);
xor U14001 (N_14001,N_13657,N_13616);
and U14002 (N_14002,N_13572,N_13525);
or U14003 (N_14003,N_13652,N_13736);
nor U14004 (N_14004,N_13704,N_13600);
and U14005 (N_14005,N_13733,N_13670);
and U14006 (N_14006,N_13685,N_13742);
nand U14007 (N_14007,N_13731,N_13659);
and U14008 (N_14008,N_13675,N_13738);
and U14009 (N_14009,N_13772,N_13623);
nor U14010 (N_14010,N_13634,N_13641);
xnor U14011 (N_14011,N_13621,N_13553);
or U14012 (N_14012,N_13657,N_13646);
nor U14013 (N_14013,N_13517,N_13611);
nor U14014 (N_14014,N_13732,N_13627);
nor U14015 (N_14015,N_13771,N_13608);
nor U14016 (N_14016,N_13592,N_13776);
nor U14017 (N_14017,N_13568,N_13696);
xnor U14018 (N_14018,N_13556,N_13774);
nor U14019 (N_14019,N_13677,N_13551);
and U14020 (N_14020,N_13657,N_13772);
nand U14021 (N_14021,N_13642,N_13779);
and U14022 (N_14022,N_13770,N_13769);
nand U14023 (N_14023,N_13762,N_13709);
or U14024 (N_14024,N_13599,N_13659);
or U14025 (N_14025,N_13536,N_13709);
or U14026 (N_14026,N_13689,N_13630);
nor U14027 (N_14027,N_13680,N_13774);
or U14028 (N_14028,N_13660,N_13630);
nor U14029 (N_14029,N_13736,N_13698);
and U14030 (N_14030,N_13528,N_13570);
xor U14031 (N_14031,N_13687,N_13549);
xnor U14032 (N_14032,N_13547,N_13613);
nor U14033 (N_14033,N_13793,N_13657);
nor U14034 (N_14034,N_13758,N_13670);
nand U14035 (N_14035,N_13695,N_13786);
nor U14036 (N_14036,N_13769,N_13679);
nor U14037 (N_14037,N_13588,N_13665);
and U14038 (N_14038,N_13628,N_13771);
and U14039 (N_14039,N_13516,N_13602);
or U14040 (N_14040,N_13659,N_13503);
and U14041 (N_14041,N_13678,N_13549);
nand U14042 (N_14042,N_13505,N_13638);
and U14043 (N_14043,N_13552,N_13629);
or U14044 (N_14044,N_13581,N_13744);
or U14045 (N_14045,N_13749,N_13772);
and U14046 (N_14046,N_13506,N_13710);
and U14047 (N_14047,N_13725,N_13712);
xnor U14048 (N_14048,N_13685,N_13710);
and U14049 (N_14049,N_13533,N_13614);
nand U14050 (N_14050,N_13783,N_13534);
nor U14051 (N_14051,N_13749,N_13694);
or U14052 (N_14052,N_13680,N_13732);
and U14053 (N_14053,N_13544,N_13548);
nand U14054 (N_14054,N_13564,N_13559);
and U14055 (N_14055,N_13506,N_13740);
or U14056 (N_14056,N_13748,N_13623);
or U14057 (N_14057,N_13674,N_13723);
nor U14058 (N_14058,N_13519,N_13580);
and U14059 (N_14059,N_13769,N_13660);
nand U14060 (N_14060,N_13760,N_13679);
or U14061 (N_14061,N_13775,N_13628);
nor U14062 (N_14062,N_13577,N_13580);
and U14063 (N_14063,N_13586,N_13767);
or U14064 (N_14064,N_13597,N_13516);
xor U14065 (N_14065,N_13649,N_13566);
or U14066 (N_14066,N_13637,N_13783);
nor U14067 (N_14067,N_13765,N_13786);
and U14068 (N_14068,N_13774,N_13513);
nand U14069 (N_14069,N_13507,N_13506);
or U14070 (N_14070,N_13785,N_13717);
and U14071 (N_14071,N_13792,N_13662);
nor U14072 (N_14072,N_13535,N_13713);
xnor U14073 (N_14073,N_13731,N_13747);
xnor U14074 (N_14074,N_13782,N_13673);
nor U14075 (N_14075,N_13513,N_13620);
xor U14076 (N_14076,N_13739,N_13543);
nand U14077 (N_14077,N_13643,N_13519);
xor U14078 (N_14078,N_13621,N_13776);
and U14079 (N_14079,N_13622,N_13776);
or U14080 (N_14080,N_13730,N_13761);
and U14081 (N_14081,N_13570,N_13776);
or U14082 (N_14082,N_13583,N_13785);
nand U14083 (N_14083,N_13625,N_13554);
or U14084 (N_14084,N_13793,N_13790);
nor U14085 (N_14085,N_13549,N_13632);
or U14086 (N_14086,N_13782,N_13753);
nand U14087 (N_14087,N_13787,N_13611);
and U14088 (N_14088,N_13727,N_13612);
nand U14089 (N_14089,N_13738,N_13781);
or U14090 (N_14090,N_13631,N_13641);
nor U14091 (N_14091,N_13741,N_13695);
nor U14092 (N_14092,N_13566,N_13612);
xor U14093 (N_14093,N_13695,N_13732);
and U14094 (N_14094,N_13720,N_13532);
nand U14095 (N_14095,N_13602,N_13514);
nor U14096 (N_14096,N_13576,N_13511);
or U14097 (N_14097,N_13513,N_13621);
and U14098 (N_14098,N_13605,N_13711);
or U14099 (N_14099,N_13613,N_13724);
nor U14100 (N_14100,N_13963,N_13855);
and U14101 (N_14101,N_13941,N_14011);
nor U14102 (N_14102,N_13845,N_13812);
nor U14103 (N_14103,N_14051,N_13873);
and U14104 (N_14104,N_13849,N_14058);
xnor U14105 (N_14105,N_13885,N_13924);
or U14106 (N_14106,N_13879,N_13906);
nand U14107 (N_14107,N_14028,N_13828);
nand U14108 (N_14108,N_14088,N_13903);
nand U14109 (N_14109,N_13836,N_14027);
and U14110 (N_14110,N_13881,N_14057);
nor U14111 (N_14111,N_13945,N_14046);
or U14112 (N_14112,N_13908,N_13982);
nor U14113 (N_14113,N_14033,N_14096);
or U14114 (N_14114,N_13859,N_13907);
or U14115 (N_14115,N_13850,N_13992);
nor U14116 (N_14116,N_13886,N_13842);
and U14117 (N_14117,N_14037,N_13882);
nand U14118 (N_14118,N_14066,N_13822);
or U14119 (N_14119,N_13834,N_13977);
and U14120 (N_14120,N_13919,N_14083);
nand U14121 (N_14121,N_14024,N_13966);
and U14122 (N_14122,N_14075,N_13918);
and U14123 (N_14123,N_13837,N_13932);
or U14124 (N_14124,N_14052,N_14004);
nor U14125 (N_14125,N_13937,N_14045);
xnor U14126 (N_14126,N_13833,N_13848);
and U14127 (N_14127,N_14056,N_13930);
xor U14128 (N_14128,N_13984,N_13957);
xor U14129 (N_14129,N_13952,N_14026);
nor U14130 (N_14130,N_13943,N_14076);
nand U14131 (N_14131,N_14097,N_13933);
or U14132 (N_14132,N_13892,N_14007);
nor U14133 (N_14133,N_13814,N_13898);
nand U14134 (N_14134,N_13806,N_14012);
or U14135 (N_14135,N_14038,N_14087);
or U14136 (N_14136,N_13928,N_14069);
nor U14137 (N_14137,N_13994,N_13962);
nor U14138 (N_14138,N_13864,N_14010);
xor U14139 (N_14139,N_13858,N_14073);
and U14140 (N_14140,N_14039,N_14062);
nor U14141 (N_14141,N_13947,N_13980);
xor U14142 (N_14142,N_13832,N_13923);
xor U14143 (N_14143,N_13803,N_13935);
nand U14144 (N_14144,N_14025,N_13893);
and U14145 (N_14145,N_13944,N_13938);
xor U14146 (N_14146,N_14005,N_14018);
and U14147 (N_14147,N_14034,N_13860);
or U14148 (N_14148,N_13874,N_13824);
and U14149 (N_14149,N_13972,N_14080);
or U14150 (N_14150,N_13857,N_13900);
nor U14151 (N_14151,N_14085,N_13851);
xor U14152 (N_14152,N_13807,N_13915);
or U14153 (N_14153,N_13989,N_14016);
xnor U14154 (N_14154,N_14041,N_13926);
and U14155 (N_14155,N_14022,N_13816);
or U14156 (N_14156,N_13958,N_13996);
nor U14157 (N_14157,N_13934,N_13916);
xnor U14158 (N_14158,N_14086,N_13896);
nor U14159 (N_14159,N_13804,N_13959);
nor U14160 (N_14160,N_13987,N_13888);
or U14161 (N_14161,N_13912,N_13844);
nor U14162 (N_14162,N_13846,N_13981);
and U14163 (N_14163,N_13993,N_14002);
nor U14164 (N_14164,N_13838,N_13920);
nand U14165 (N_14165,N_13854,N_14014);
xnor U14166 (N_14166,N_13956,N_14090);
xnor U14167 (N_14167,N_13840,N_13946);
and U14168 (N_14168,N_13868,N_14078);
nand U14169 (N_14169,N_14048,N_13999);
nand U14170 (N_14170,N_14019,N_14023);
nor U14171 (N_14171,N_13931,N_14054);
nand U14172 (N_14172,N_13922,N_14053);
nand U14173 (N_14173,N_13884,N_14036);
and U14174 (N_14174,N_13948,N_13964);
xor U14175 (N_14175,N_13867,N_13883);
nand U14176 (N_14176,N_14095,N_13852);
and U14177 (N_14177,N_13936,N_14092);
nor U14178 (N_14178,N_14091,N_13819);
nor U14179 (N_14179,N_13843,N_13835);
xor U14180 (N_14180,N_13856,N_13974);
or U14181 (N_14181,N_13942,N_13865);
nand U14182 (N_14182,N_14035,N_13950);
nand U14183 (N_14183,N_13809,N_13979);
nand U14184 (N_14184,N_14068,N_13940);
xor U14185 (N_14185,N_13818,N_13927);
xor U14186 (N_14186,N_13967,N_13925);
nand U14187 (N_14187,N_13990,N_13861);
xnor U14188 (N_14188,N_14013,N_14020);
xor U14189 (N_14189,N_13813,N_14001);
xor U14190 (N_14190,N_13902,N_13899);
or U14191 (N_14191,N_14082,N_14077);
nor U14192 (N_14192,N_14044,N_14079);
nand U14193 (N_14193,N_13889,N_13969);
nor U14194 (N_14194,N_14093,N_14060);
and U14195 (N_14195,N_13826,N_13805);
xnor U14196 (N_14196,N_14063,N_13917);
or U14197 (N_14197,N_14055,N_13965);
or U14198 (N_14198,N_14072,N_13904);
and U14199 (N_14199,N_13901,N_13817);
and U14200 (N_14200,N_14029,N_14049);
nor U14201 (N_14201,N_13929,N_13951);
nor U14202 (N_14202,N_13995,N_13880);
nand U14203 (N_14203,N_13876,N_13991);
and U14204 (N_14204,N_14030,N_13983);
nor U14205 (N_14205,N_13862,N_13968);
nand U14206 (N_14206,N_13827,N_14003);
or U14207 (N_14207,N_13953,N_14017);
nor U14208 (N_14208,N_14098,N_13853);
xor U14209 (N_14209,N_13988,N_13985);
or U14210 (N_14210,N_13895,N_13800);
and U14211 (N_14211,N_14047,N_14067);
and U14212 (N_14212,N_14070,N_13975);
nand U14213 (N_14213,N_14074,N_13821);
nor U14214 (N_14214,N_13913,N_13914);
nor U14215 (N_14215,N_13830,N_14081);
and U14216 (N_14216,N_14059,N_14032);
and U14217 (N_14217,N_13970,N_13829);
nand U14218 (N_14218,N_14031,N_13939);
and U14219 (N_14219,N_13954,N_13887);
or U14220 (N_14220,N_13820,N_13811);
or U14221 (N_14221,N_14043,N_13877);
or U14222 (N_14222,N_13808,N_13872);
nand U14223 (N_14223,N_13870,N_13823);
nand U14224 (N_14224,N_13910,N_14006);
nand U14225 (N_14225,N_13955,N_14064);
and U14226 (N_14226,N_13831,N_13894);
xor U14227 (N_14227,N_13905,N_13878);
xor U14228 (N_14228,N_13815,N_13841);
and U14229 (N_14229,N_13949,N_14000);
xnor U14230 (N_14230,N_13960,N_14094);
nand U14231 (N_14231,N_13976,N_13890);
nor U14232 (N_14232,N_13863,N_14021);
and U14233 (N_14233,N_14042,N_13802);
nand U14234 (N_14234,N_13997,N_13891);
xor U14235 (N_14235,N_13978,N_13911);
or U14236 (N_14236,N_14015,N_14050);
nor U14237 (N_14237,N_13971,N_13897);
nand U14238 (N_14238,N_14099,N_14040);
nor U14239 (N_14239,N_13866,N_14009);
xor U14240 (N_14240,N_14084,N_13839);
xnor U14241 (N_14241,N_13801,N_13869);
nand U14242 (N_14242,N_13810,N_13909);
and U14243 (N_14243,N_13961,N_13825);
xor U14244 (N_14244,N_13875,N_13998);
nor U14245 (N_14245,N_13847,N_14061);
nor U14246 (N_14246,N_14008,N_13986);
or U14247 (N_14247,N_13921,N_14065);
or U14248 (N_14248,N_13871,N_13973);
or U14249 (N_14249,N_14071,N_14089);
nor U14250 (N_14250,N_14058,N_13885);
xnor U14251 (N_14251,N_13910,N_14058);
nor U14252 (N_14252,N_13959,N_14049);
nand U14253 (N_14253,N_13910,N_13804);
xor U14254 (N_14254,N_14054,N_13888);
xor U14255 (N_14255,N_13806,N_14043);
or U14256 (N_14256,N_13899,N_13842);
nor U14257 (N_14257,N_13829,N_13825);
or U14258 (N_14258,N_14096,N_14066);
xnor U14259 (N_14259,N_14089,N_13983);
and U14260 (N_14260,N_14020,N_13873);
nand U14261 (N_14261,N_13968,N_13978);
or U14262 (N_14262,N_13920,N_14010);
nor U14263 (N_14263,N_14094,N_13901);
or U14264 (N_14264,N_14007,N_14079);
nand U14265 (N_14265,N_14019,N_13950);
or U14266 (N_14266,N_13899,N_13830);
nand U14267 (N_14267,N_13825,N_13835);
nor U14268 (N_14268,N_14086,N_13917);
or U14269 (N_14269,N_13810,N_13804);
nor U14270 (N_14270,N_13934,N_13920);
xnor U14271 (N_14271,N_13923,N_14030);
nor U14272 (N_14272,N_13856,N_13899);
or U14273 (N_14273,N_14084,N_13807);
and U14274 (N_14274,N_13913,N_14033);
xor U14275 (N_14275,N_14022,N_13977);
or U14276 (N_14276,N_13846,N_13821);
xnor U14277 (N_14277,N_13804,N_14002);
xnor U14278 (N_14278,N_13859,N_13903);
or U14279 (N_14279,N_13815,N_13930);
or U14280 (N_14280,N_13940,N_13886);
or U14281 (N_14281,N_13924,N_14055);
xnor U14282 (N_14282,N_14036,N_14034);
xnor U14283 (N_14283,N_13990,N_13963);
and U14284 (N_14284,N_14002,N_14031);
nand U14285 (N_14285,N_13974,N_13809);
nor U14286 (N_14286,N_13891,N_13976);
and U14287 (N_14287,N_13992,N_14061);
xnor U14288 (N_14288,N_14046,N_13903);
and U14289 (N_14289,N_13954,N_13992);
nor U14290 (N_14290,N_14072,N_13880);
or U14291 (N_14291,N_13892,N_13950);
nor U14292 (N_14292,N_13974,N_14081);
or U14293 (N_14293,N_13920,N_13822);
xnor U14294 (N_14294,N_13961,N_13965);
or U14295 (N_14295,N_14035,N_14087);
nand U14296 (N_14296,N_14026,N_13868);
nand U14297 (N_14297,N_13803,N_13954);
nor U14298 (N_14298,N_13876,N_13842);
nand U14299 (N_14299,N_13912,N_13811);
or U14300 (N_14300,N_13864,N_13809);
and U14301 (N_14301,N_13835,N_14052);
and U14302 (N_14302,N_13883,N_13858);
nand U14303 (N_14303,N_13934,N_14040);
or U14304 (N_14304,N_13949,N_13877);
nand U14305 (N_14305,N_13868,N_14065);
and U14306 (N_14306,N_13880,N_13977);
nor U14307 (N_14307,N_14068,N_13819);
and U14308 (N_14308,N_14027,N_14095);
or U14309 (N_14309,N_13828,N_13873);
and U14310 (N_14310,N_13862,N_13932);
nor U14311 (N_14311,N_13825,N_13941);
and U14312 (N_14312,N_13837,N_13934);
xor U14313 (N_14313,N_13878,N_13970);
xor U14314 (N_14314,N_14056,N_13914);
or U14315 (N_14315,N_13909,N_14019);
and U14316 (N_14316,N_13933,N_14018);
xnor U14317 (N_14317,N_13870,N_13953);
nor U14318 (N_14318,N_13941,N_14074);
nand U14319 (N_14319,N_13913,N_13972);
nand U14320 (N_14320,N_13826,N_13867);
or U14321 (N_14321,N_13918,N_14091);
nor U14322 (N_14322,N_13826,N_13871);
xnor U14323 (N_14323,N_14058,N_13903);
nor U14324 (N_14324,N_14006,N_13947);
nand U14325 (N_14325,N_13884,N_13817);
xor U14326 (N_14326,N_13997,N_13844);
or U14327 (N_14327,N_14022,N_13970);
and U14328 (N_14328,N_14041,N_13952);
nor U14329 (N_14329,N_14039,N_13998);
and U14330 (N_14330,N_13879,N_13963);
xnor U14331 (N_14331,N_13825,N_13995);
or U14332 (N_14332,N_14030,N_13942);
xnor U14333 (N_14333,N_13999,N_13858);
nor U14334 (N_14334,N_13956,N_13855);
or U14335 (N_14335,N_13890,N_13824);
and U14336 (N_14336,N_13880,N_14079);
nor U14337 (N_14337,N_13802,N_14008);
nand U14338 (N_14338,N_13899,N_13877);
xor U14339 (N_14339,N_14085,N_13900);
nor U14340 (N_14340,N_13856,N_13874);
and U14341 (N_14341,N_13946,N_13870);
nor U14342 (N_14342,N_13979,N_13875);
or U14343 (N_14343,N_13960,N_13992);
nand U14344 (N_14344,N_13890,N_13889);
nor U14345 (N_14345,N_13918,N_13818);
xor U14346 (N_14346,N_14007,N_13914);
and U14347 (N_14347,N_13908,N_14072);
and U14348 (N_14348,N_14022,N_14058);
and U14349 (N_14349,N_14073,N_13919);
or U14350 (N_14350,N_13902,N_14093);
nor U14351 (N_14351,N_13947,N_14074);
xor U14352 (N_14352,N_13842,N_13901);
nor U14353 (N_14353,N_13937,N_13979);
and U14354 (N_14354,N_14071,N_14099);
and U14355 (N_14355,N_13835,N_14044);
nand U14356 (N_14356,N_13859,N_13869);
or U14357 (N_14357,N_14057,N_13823);
or U14358 (N_14358,N_14057,N_13815);
nor U14359 (N_14359,N_14076,N_14023);
and U14360 (N_14360,N_13987,N_13901);
nand U14361 (N_14361,N_13831,N_14073);
and U14362 (N_14362,N_13894,N_14077);
nor U14363 (N_14363,N_13905,N_14071);
or U14364 (N_14364,N_13806,N_13876);
nand U14365 (N_14365,N_13935,N_13828);
or U14366 (N_14366,N_13947,N_13892);
and U14367 (N_14367,N_13888,N_14076);
or U14368 (N_14368,N_14040,N_13970);
nor U14369 (N_14369,N_13815,N_13802);
nand U14370 (N_14370,N_13867,N_14073);
xor U14371 (N_14371,N_14047,N_14013);
or U14372 (N_14372,N_13912,N_13966);
nor U14373 (N_14373,N_13824,N_14089);
xnor U14374 (N_14374,N_13868,N_14063);
xor U14375 (N_14375,N_14085,N_14048);
nand U14376 (N_14376,N_14083,N_13943);
or U14377 (N_14377,N_14031,N_14013);
nand U14378 (N_14378,N_13966,N_13876);
xnor U14379 (N_14379,N_13982,N_13996);
nor U14380 (N_14380,N_13892,N_14065);
xnor U14381 (N_14381,N_13922,N_13815);
or U14382 (N_14382,N_14039,N_13899);
nand U14383 (N_14383,N_13821,N_13884);
nand U14384 (N_14384,N_13973,N_13923);
or U14385 (N_14385,N_13864,N_13947);
nand U14386 (N_14386,N_14004,N_14070);
and U14387 (N_14387,N_14001,N_13935);
nand U14388 (N_14388,N_13886,N_13976);
and U14389 (N_14389,N_13891,N_13918);
nand U14390 (N_14390,N_13951,N_13820);
nor U14391 (N_14391,N_14091,N_13951);
nand U14392 (N_14392,N_13819,N_13938);
and U14393 (N_14393,N_14042,N_13903);
and U14394 (N_14394,N_13867,N_13877);
xnor U14395 (N_14395,N_13888,N_14033);
nor U14396 (N_14396,N_13841,N_13965);
nand U14397 (N_14397,N_13853,N_14000);
and U14398 (N_14398,N_13865,N_13876);
nand U14399 (N_14399,N_13982,N_13999);
xnor U14400 (N_14400,N_14303,N_14326);
nor U14401 (N_14401,N_14127,N_14133);
or U14402 (N_14402,N_14392,N_14113);
and U14403 (N_14403,N_14355,N_14226);
nor U14404 (N_14404,N_14117,N_14324);
nor U14405 (N_14405,N_14105,N_14233);
nor U14406 (N_14406,N_14321,N_14311);
or U14407 (N_14407,N_14190,N_14281);
xnor U14408 (N_14408,N_14203,N_14309);
or U14409 (N_14409,N_14371,N_14327);
or U14410 (N_14410,N_14254,N_14108);
xnor U14411 (N_14411,N_14214,N_14363);
xnor U14412 (N_14412,N_14194,N_14393);
xnor U14413 (N_14413,N_14147,N_14273);
and U14414 (N_14414,N_14338,N_14128);
xor U14415 (N_14415,N_14339,N_14302);
xnor U14416 (N_14416,N_14395,N_14143);
nor U14417 (N_14417,N_14232,N_14141);
nor U14418 (N_14418,N_14204,N_14390);
or U14419 (N_14419,N_14140,N_14184);
nor U14420 (N_14420,N_14343,N_14139);
or U14421 (N_14421,N_14360,N_14152);
xnor U14422 (N_14422,N_14283,N_14200);
nand U14423 (N_14423,N_14174,N_14157);
xor U14424 (N_14424,N_14307,N_14196);
or U14425 (N_14425,N_14323,N_14169);
nor U14426 (N_14426,N_14195,N_14336);
and U14427 (N_14427,N_14259,N_14124);
nand U14428 (N_14428,N_14359,N_14236);
nand U14429 (N_14429,N_14367,N_14189);
nand U14430 (N_14430,N_14384,N_14153);
or U14431 (N_14431,N_14347,N_14242);
and U14432 (N_14432,N_14224,N_14261);
and U14433 (N_14433,N_14301,N_14193);
nand U14434 (N_14434,N_14375,N_14315);
and U14435 (N_14435,N_14356,N_14357);
and U14436 (N_14436,N_14154,N_14310);
nor U14437 (N_14437,N_14344,N_14148);
nand U14438 (N_14438,N_14144,N_14378);
or U14439 (N_14439,N_14126,N_14138);
and U14440 (N_14440,N_14364,N_14318);
xor U14441 (N_14441,N_14239,N_14175);
nand U14442 (N_14442,N_14276,N_14192);
xor U14443 (N_14443,N_14216,N_14369);
nand U14444 (N_14444,N_14280,N_14350);
nor U14445 (N_14445,N_14334,N_14372);
and U14446 (N_14446,N_14181,N_14387);
or U14447 (N_14447,N_14304,N_14100);
and U14448 (N_14448,N_14337,N_14349);
nor U14449 (N_14449,N_14180,N_14293);
xnor U14450 (N_14450,N_14149,N_14215);
or U14451 (N_14451,N_14296,N_14109);
and U14452 (N_14452,N_14238,N_14253);
or U14453 (N_14453,N_14201,N_14322);
nor U14454 (N_14454,N_14156,N_14110);
or U14455 (N_14455,N_14185,N_14208);
xor U14456 (N_14456,N_14379,N_14223);
and U14457 (N_14457,N_14289,N_14222);
nand U14458 (N_14458,N_14212,N_14246);
or U14459 (N_14459,N_14329,N_14155);
nand U14460 (N_14460,N_14365,N_14134);
nand U14461 (N_14461,N_14277,N_14166);
and U14462 (N_14462,N_14107,N_14179);
nand U14463 (N_14463,N_14217,N_14111);
nand U14464 (N_14464,N_14167,N_14263);
and U14465 (N_14465,N_14206,N_14219);
nand U14466 (N_14466,N_14243,N_14374);
xor U14467 (N_14467,N_14396,N_14244);
and U14468 (N_14468,N_14299,N_14142);
xnor U14469 (N_14469,N_14399,N_14398);
nor U14470 (N_14470,N_14207,N_14171);
xnor U14471 (N_14471,N_14165,N_14116);
nor U14472 (N_14472,N_14294,N_14397);
xnor U14473 (N_14473,N_14231,N_14377);
and U14474 (N_14474,N_14366,N_14319);
and U14475 (N_14475,N_14255,N_14183);
xor U14476 (N_14476,N_14267,N_14136);
nand U14477 (N_14477,N_14101,N_14227);
nand U14478 (N_14478,N_14146,N_14228);
nor U14479 (N_14479,N_14122,N_14210);
or U14480 (N_14480,N_14320,N_14187);
nor U14481 (N_14481,N_14285,N_14331);
xnor U14482 (N_14482,N_14229,N_14197);
and U14483 (N_14483,N_14330,N_14265);
and U14484 (N_14484,N_14172,N_14115);
and U14485 (N_14485,N_14119,N_14394);
xor U14486 (N_14486,N_14383,N_14264);
nor U14487 (N_14487,N_14177,N_14368);
xnor U14488 (N_14488,N_14158,N_14252);
or U14489 (N_14489,N_14235,N_14328);
xnor U14490 (N_14490,N_14258,N_14354);
or U14491 (N_14491,N_14316,N_14121);
nor U14492 (N_14492,N_14314,N_14389);
nand U14493 (N_14493,N_14295,N_14361);
xor U14494 (N_14494,N_14298,N_14102);
nand U14495 (N_14495,N_14352,N_14256);
and U14496 (N_14496,N_14287,N_14297);
nand U14497 (N_14497,N_14106,N_14345);
nor U14498 (N_14498,N_14151,N_14300);
xor U14499 (N_14499,N_14291,N_14234);
xnor U14500 (N_14500,N_14135,N_14286);
or U14501 (N_14501,N_14353,N_14186);
nand U14502 (N_14502,N_14278,N_14305);
nor U14503 (N_14503,N_14332,N_14198);
nand U14504 (N_14504,N_14351,N_14130);
xor U14505 (N_14505,N_14325,N_14292);
or U14506 (N_14506,N_14274,N_14209);
xnor U14507 (N_14507,N_14218,N_14112);
xor U14508 (N_14508,N_14120,N_14268);
nor U14509 (N_14509,N_14346,N_14103);
xor U14510 (N_14510,N_14241,N_14386);
nor U14511 (N_14511,N_14178,N_14362);
nor U14512 (N_14512,N_14163,N_14131);
and U14513 (N_14513,N_14245,N_14125);
and U14514 (N_14514,N_14247,N_14104);
or U14515 (N_14515,N_14290,N_14176);
xnor U14516 (N_14516,N_14358,N_14317);
nand U14517 (N_14517,N_14257,N_14341);
nand U14518 (N_14518,N_14118,N_14279);
or U14519 (N_14519,N_14342,N_14182);
xor U14520 (N_14520,N_14308,N_14266);
nor U14521 (N_14521,N_14282,N_14260);
and U14522 (N_14522,N_14391,N_14145);
xnor U14523 (N_14523,N_14199,N_14284);
nor U14524 (N_14524,N_14240,N_14312);
and U14525 (N_14525,N_14271,N_14313);
or U14526 (N_14526,N_14225,N_14251);
xor U14527 (N_14527,N_14221,N_14248);
nand U14528 (N_14528,N_14160,N_14205);
and U14529 (N_14529,N_14388,N_14188);
nor U14530 (N_14530,N_14275,N_14173);
and U14531 (N_14531,N_14370,N_14164);
nor U14532 (N_14532,N_14150,N_14340);
nor U14533 (N_14533,N_14262,N_14270);
nand U14534 (N_14534,N_14168,N_14382);
nand U14535 (N_14535,N_14230,N_14161);
nor U14536 (N_14536,N_14385,N_14123);
and U14537 (N_14537,N_14272,N_14202);
nand U14538 (N_14538,N_14333,N_14373);
nand U14539 (N_14539,N_14237,N_14306);
nand U14540 (N_14540,N_14380,N_14269);
nand U14541 (N_14541,N_14132,N_14213);
and U14542 (N_14542,N_14335,N_14220);
xnor U14543 (N_14543,N_14249,N_14129);
or U14544 (N_14544,N_14288,N_14211);
or U14545 (N_14545,N_14191,N_14114);
and U14546 (N_14546,N_14170,N_14381);
nor U14547 (N_14547,N_14137,N_14348);
and U14548 (N_14548,N_14376,N_14162);
nand U14549 (N_14549,N_14250,N_14159);
nand U14550 (N_14550,N_14198,N_14295);
or U14551 (N_14551,N_14196,N_14277);
nand U14552 (N_14552,N_14344,N_14341);
nor U14553 (N_14553,N_14393,N_14374);
and U14554 (N_14554,N_14312,N_14175);
xnor U14555 (N_14555,N_14169,N_14297);
or U14556 (N_14556,N_14156,N_14259);
xor U14557 (N_14557,N_14165,N_14260);
xor U14558 (N_14558,N_14377,N_14270);
and U14559 (N_14559,N_14298,N_14130);
xor U14560 (N_14560,N_14370,N_14272);
and U14561 (N_14561,N_14234,N_14245);
and U14562 (N_14562,N_14187,N_14314);
nor U14563 (N_14563,N_14348,N_14196);
nor U14564 (N_14564,N_14174,N_14101);
nor U14565 (N_14565,N_14283,N_14116);
xnor U14566 (N_14566,N_14266,N_14315);
or U14567 (N_14567,N_14226,N_14314);
nor U14568 (N_14568,N_14153,N_14331);
nor U14569 (N_14569,N_14358,N_14395);
and U14570 (N_14570,N_14323,N_14211);
xor U14571 (N_14571,N_14301,N_14132);
or U14572 (N_14572,N_14246,N_14354);
and U14573 (N_14573,N_14101,N_14294);
xor U14574 (N_14574,N_14177,N_14343);
xor U14575 (N_14575,N_14245,N_14101);
nand U14576 (N_14576,N_14303,N_14308);
or U14577 (N_14577,N_14117,N_14317);
or U14578 (N_14578,N_14160,N_14329);
xor U14579 (N_14579,N_14113,N_14391);
xnor U14580 (N_14580,N_14135,N_14282);
xor U14581 (N_14581,N_14242,N_14112);
and U14582 (N_14582,N_14393,N_14157);
nand U14583 (N_14583,N_14390,N_14155);
xnor U14584 (N_14584,N_14255,N_14382);
nand U14585 (N_14585,N_14368,N_14167);
and U14586 (N_14586,N_14218,N_14282);
and U14587 (N_14587,N_14240,N_14187);
and U14588 (N_14588,N_14315,N_14302);
nand U14589 (N_14589,N_14343,N_14218);
and U14590 (N_14590,N_14312,N_14237);
nor U14591 (N_14591,N_14105,N_14191);
xor U14592 (N_14592,N_14280,N_14329);
xor U14593 (N_14593,N_14386,N_14317);
or U14594 (N_14594,N_14102,N_14121);
or U14595 (N_14595,N_14159,N_14223);
xor U14596 (N_14596,N_14286,N_14331);
or U14597 (N_14597,N_14341,N_14113);
or U14598 (N_14598,N_14106,N_14145);
or U14599 (N_14599,N_14186,N_14143);
or U14600 (N_14600,N_14233,N_14282);
and U14601 (N_14601,N_14398,N_14208);
nand U14602 (N_14602,N_14255,N_14160);
and U14603 (N_14603,N_14267,N_14398);
nand U14604 (N_14604,N_14140,N_14249);
xor U14605 (N_14605,N_14332,N_14179);
nor U14606 (N_14606,N_14379,N_14325);
xor U14607 (N_14607,N_14295,N_14220);
and U14608 (N_14608,N_14180,N_14277);
or U14609 (N_14609,N_14366,N_14231);
xnor U14610 (N_14610,N_14176,N_14251);
xor U14611 (N_14611,N_14230,N_14353);
xor U14612 (N_14612,N_14172,N_14152);
xor U14613 (N_14613,N_14214,N_14287);
nor U14614 (N_14614,N_14308,N_14173);
nand U14615 (N_14615,N_14332,N_14387);
xor U14616 (N_14616,N_14106,N_14360);
xnor U14617 (N_14617,N_14322,N_14242);
nor U14618 (N_14618,N_14177,N_14142);
or U14619 (N_14619,N_14127,N_14193);
xnor U14620 (N_14620,N_14297,N_14191);
or U14621 (N_14621,N_14203,N_14379);
or U14622 (N_14622,N_14393,N_14117);
and U14623 (N_14623,N_14323,N_14124);
or U14624 (N_14624,N_14114,N_14383);
and U14625 (N_14625,N_14252,N_14117);
and U14626 (N_14626,N_14147,N_14163);
nand U14627 (N_14627,N_14174,N_14133);
nand U14628 (N_14628,N_14110,N_14280);
xor U14629 (N_14629,N_14386,N_14139);
nor U14630 (N_14630,N_14353,N_14229);
nand U14631 (N_14631,N_14139,N_14159);
nor U14632 (N_14632,N_14312,N_14399);
nor U14633 (N_14633,N_14220,N_14384);
nand U14634 (N_14634,N_14147,N_14370);
nand U14635 (N_14635,N_14276,N_14269);
xnor U14636 (N_14636,N_14267,N_14274);
and U14637 (N_14637,N_14164,N_14394);
nor U14638 (N_14638,N_14196,N_14227);
and U14639 (N_14639,N_14153,N_14111);
or U14640 (N_14640,N_14228,N_14148);
nand U14641 (N_14641,N_14364,N_14345);
or U14642 (N_14642,N_14316,N_14391);
nor U14643 (N_14643,N_14156,N_14245);
nand U14644 (N_14644,N_14297,N_14199);
or U14645 (N_14645,N_14344,N_14364);
xnor U14646 (N_14646,N_14252,N_14264);
nand U14647 (N_14647,N_14177,N_14190);
xnor U14648 (N_14648,N_14138,N_14342);
nor U14649 (N_14649,N_14236,N_14139);
and U14650 (N_14650,N_14272,N_14247);
or U14651 (N_14651,N_14318,N_14143);
or U14652 (N_14652,N_14189,N_14100);
and U14653 (N_14653,N_14156,N_14302);
nand U14654 (N_14654,N_14364,N_14214);
nand U14655 (N_14655,N_14383,N_14336);
xnor U14656 (N_14656,N_14196,N_14180);
nor U14657 (N_14657,N_14268,N_14304);
xnor U14658 (N_14658,N_14189,N_14261);
nand U14659 (N_14659,N_14188,N_14157);
xnor U14660 (N_14660,N_14206,N_14348);
nor U14661 (N_14661,N_14398,N_14285);
nand U14662 (N_14662,N_14323,N_14271);
xor U14663 (N_14663,N_14373,N_14396);
nor U14664 (N_14664,N_14260,N_14353);
nand U14665 (N_14665,N_14234,N_14114);
nor U14666 (N_14666,N_14100,N_14367);
nor U14667 (N_14667,N_14143,N_14194);
nor U14668 (N_14668,N_14388,N_14317);
nand U14669 (N_14669,N_14162,N_14230);
nor U14670 (N_14670,N_14362,N_14184);
and U14671 (N_14671,N_14189,N_14319);
or U14672 (N_14672,N_14338,N_14319);
nand U14673 (N_14673,N_14225,N_14207);
or U14674 (N_14674,N_14319,N_14267);
and U14675 (N_14675,N_14246,N_14232);
and U14676 (N_14676,N_14242,N_14227);
nor U14677 (N_14677,N_14251,N_14191);
nand U14678 (N_14678,N_14291,N_14371);
xor U14679 (N_14679,N_14331,N_14248);
and U14680 (N_14680,N_14139,N_14247);
or U14681 (N_14681,N_14228,N_14304);
or U14682 (N_14682,N_14288,N_14327);
and U14683 (N_14683,N_14232,N_14151);
nor U14684 (N_14684,N_14157,N_14201);
xor U14685 (N_14685,N_14274,N_14352);
nand U14686 (N_14686,N_14108,N_14288);
nor U14687 (N_14687,N_14338,N_14344);
xnor U14688 (N_14688,N_14167,N_14156);
or U14689 (N_14689,N_14239,N_14186);
or U14690 (N_14690,N_14389,N_14341);
nor U14691 (N_14691,N_14141,N_14199);
xor U14692 (N_14692,N_14249,N_14350);
nor U14693 (N_14693,N_14120,N_14202);
and U14694 (N_14694,N_14119,N_14178);
xnor U14695 (N_14695,N_14393,N_14241);
nor U14696 (N_14696,N_14397,N_14285);
and U14697 (N_14697,N_14213,N_14246);
and U14698 (N_14698,N_14302,N_14216);
xnor U14699 (N_14699,N_14265,N_14379);
nand U14700 (N_14700,N_14685,N_14691);
and U14701 (N_14701,N_14672,N_14525);
xor U14702 (N_14702,N_14689,N_14619);
and U14703 (N_14703,N_14499,N_14526);
and U14704 (N_14704,N_14435,N_14573);
nand U14705 (N_14705,N_14652,N_14637);
nor U14706 (N_14706,N_14469,N_14520);
or U14707 (N_14707,N_14468,N_14661);
xnor U14708 (N_14708,N_14480,N_14698);
xor U14709 (N_14709,N_14549,N_14500);
xnor U14710 (N_14710,N_14627,N_14544);
xor U14711 (N_14711,N_14572,N_14502);
or U14712 (N_14712,N_14460,N_14571);
nor U14713 (N_14713,N_14603,N_14472);
nor U14714 (N_14714,N_14495,N_14583);
or U14715 (N_14715,N_14453,N_14416);
and U14716 (N_14716,N_14431,N_14424);
xor U14717 (N_14717,N_14481,N_14446);
nor U14718 (N_14718,N_14629,N_14442);
xor U14719 (N_14719,N_14479,N_14498);
and U14720 (N_14720,N_14462,N_14546);
nor U14721 (N_14721,N_14615,N_14632);
nand U14722 (N_14722,N_14675,N_14678);
and U14723 (N_14723,N_14686,N_14595);
and U14724 (N_14724,N_14599,N_14579);
nand U14725 (N_14725,N_14411,N_14445);
xor U14726 (N_14726,N_14427,N_14584);
nor U14727 (N_14727,N_14621,N_14659);
nor U14728 (N_14728,N_14646,N_14604);
xnor U14729 (N_14729,N_14475,N_14524);
or U14730 (N_14730,N_14417,N_14485);
or U14731 (N_14731,N_14438,N_14553);
nor U14732 (N_14732,N_14669,N_14602);
nor U14733 (N_14733,N_14641,N_14484);
nand U14734 (N_14734,N_14654,N_14692);
nor U14735 (N_14735,N_14593,N_14666);
nor U14736 (N_14736,N_14492,N_14664);
nor U14737 (N_14737,N_14653,N_14455);
xor U14738 (N_14738,N_14577,N_14566);
xnor U14739 (N_14739,N_14441,N_14665);
xor U14740 (N_14740,N_14589,N_14503);
nand U14741 (N_14741,N_14562,N_14412);
or U14742 (N_14742,N_14631,N_14555);
nand U14743 (N_14743,N_14477,N_14620);
or U14744 (N_14744,N_14418,N_14539);
nor U14745 (N_14745,N_14426,N_14406);
and U14746 (N_14746,N_14581,N_14567);
nor U14747 (N_14747,N_14505,N_14532);
or U14748 (N_14748,N_14676,N_14682);
and U14749 (N_14749,N_14671,N_14542);
nor U14750 (N_14750,N_14448,N_14636);
nor U14751 (N_14751,N_14568,N_14528);
xnor U14752 (N_14752,N_14487,N_14556);
xor U14753 (N_14753,N_14440,N_14456);
xnor U14754 (N_14754,N_14694,N_14496);
and U14755 (N_14755,N_14611,N_14575);
nor U14756 (N_14756,N_14516,N_14450);
xor U14757 (N_14757,N_14439,N_14404);
nand U14758 (N_14758,N_14624,N_14633);
or U14759 (N_14759,N_14425,N_14606);
nor U14760 (N_14760,N_14443,N_14600);
nand U14761 (N_14761,N_14504,N_14634);
and U14762 (N_14762,N_14409,N_14402);
nand U14763 (N_14763,N_14420,N_14569);
and U14764 (N_14764,N_14642,N_14407);
nor U14765 (N_14765,N_14580,N_14623);
nand U14766 (N_14766,N_14405,N_14697);
xnor U14767 (N_14767,N_14563,N_14527);
or U14768 (N_14768,N_14605,N_14558);
xnor U14769 (N_14769,N_14510,N_14582);
and U14770 (N_14770,N_14533,N_14649);
nand U14771 (N_14771,N_14552,N_14518);
or U14772 (N_14772,N_14464,N_14559);
nor U14773 (N_14773,N_14540,N_14433);
nor U14774 (N_14774,N_14491,N_14414);
nor U14775 (N_14775,N_14413,N_14594);
nor U14776 (N_14776,N_14423,N_14537);
and U14777 (N_14777,N_14459,N_14529);
or U14778 (N_14778,N_14578,N_14436);
nand U14779 (N_14779,N_14638,N_14557);
and U14780 (N_14780,N_14574,N_14651);
nand U14781 (N_14781,N_14644,N_14628);
nor U14782 (N_14782,N_14512,N_14639);
and U14783 (N_14783,N_14630,N_14506);
nand U14784 (N_14784,N_14509,N_14488);
nor U14785 (N_14785,N_14400,N_14660);
and U14786 (N_14786,N_14507,N_14690);
nand U14787 (N_14787,N_14403,N_14517);
or U14788 (N_14788,N_14538,N_14667);
or U14789 (N_14789,N_14545,N_14514);
and U14790 (N_14790,N_14622,N_14618);
nor U14791 (N_14791,N_14590,N_14596);
nand U14792 (N_14792,N_14658,N_14696);
nor U14793 (N_14793,N_14493,N_14560);
and U14794 (N_14794,N_14449,N_14657);
nor U14795 (N_14795,N_14673,N_14482);
or U14796 (N_14796,N_14430,N_14597);
xnor U14797 (N_14797,N_14457,N_14601);
and U14798 (N_14798,N_14677,N_14598);
and U14799 (N_14799,N_14463,N_14536);
nand U14800 (N_14800,N_14501,N_14591);
or U14801 (N_14801,N_14693,N_14454);
or U14802 (N_14802,N_14429,N_14415);
or U14803 (N_14803,N_14541,N_14519);
or U14804 (N_14804,N_14473,N_14663);
xor U14805 (N_14805,N_14662,N_14616);
nor U14806 (N_14806,N_14643,N_14640);
nor U14807 (N_14807,N_14551,N_14683);
or U14808 (N_14808,N_14474,N_14699);
and U14809 (N_14809,N_14452,N_14587);
nand U14810 (N_14810,N_14610,N_14437);
or U14811 (N_14811,N_14655,N_14410);
nand U14812 (N_14812,N_14523,N_14648);
or U14813 (N_14813,N_14458,N_14466);
or U14814 (N_14814,N_14679,N_14508);
nor U14815 (N_14815,N_14550,N_14576);
or U14816 (N_14816,N_14680,N_14419);
or U14817 (N_14817,N_14434,N_14554);
nand U14818 (N_14818,N_14465,N_14674);
nor U14819 (N_14819,N_14489,N_14647);
nor U14820 (N_14820,N_14656,N_14592);
xor U14821 (N_14821,N_14650,N_14586);
xnor U14822 (N_14822,N_14695,N_14534);
and U14823 (N_14823,N_14564,N_14530);
nand U14824 (N_14824,N_14585,N_14570);
and U14825 (N_14825,N_14531,N_14607);
or U14826 (N_14826,N_14588,N_14612);
nand U14827 (N_14827,N_14645,N_14561);
nor U14828 (N_14828,N_14608,N_14626);
xnor U14829 (N_14829,N_14471,N_14614);
and U14830 (N_14830,N_14522,N_14609);
or U14831 (N_14831,N_14421,N_14668);
or U14832 (N_14832,N_14483,N_14547);
and U14833 (N_14833,N_14635,N_14497);
nand U14834 (N_14834,N_14548,N_14478);
or U14835 (N_14835,N_14625,N_14681);
or U14836 (N_14836,N_14684,N_14401);
or U14837 (N_14837,N_14486,N_14461);
nor U14838 (N_14838,N_14670,N_14521);
and U14839 (N_14839,N_14513,N_14476);
or U14840 (N_14840,N_14408,N_14494);
or U14841 (N_14841,N_14447,N_14688);
or U14842 (N_14842,N_14535,N_14515);
or U14843 (N_14843,N_14422,N_14451);
nor U14844 (N_14844,N_14490,N_14432);
xnor U14845 (N_14845,N_14470,N_14543);
and U14846 (N_14846,N_14565,N_14613);
or U14847 (N_14847,N_14428,N_14511);
and U14848 (N_14848,N_14687,N_14444);
nor U14849 (N_14849,N_14617,N_14467);
or U14850 (N_14850,N_14420,N_14419);
nand U14851 (N_14851,N_14437,N_14535);
or U14852 (N_14852,N_14401,N_14607);
nor U14853 (N_14853,N_14462,N_14489);
or U14854 (N_14854,N_14697,N_14497);
and U14855 (N_14855,N_14534,N_14594);
or U14856 (N_14856,N_14667,N_14606);
xnor U14857 (N_14857,N_14434,N_14452);
nand U14858 (N_14858,N_14598,N_14649);
nor U14859 (N_14859,N_14677,N_14488);
or U14860 (N_14860,N_14611,N_14426);
xor U14861 (N_14861,N_14438,N_14571);
nor U14862 (N_14862,N_14619,N_14631);
or U14863 (N_14863,N_14618,N_14692);
nand U14864 (N_14864,N_14474,N_14666);
and U14865 (N_14865,N_14545,N_14401);
xnor U14866 (N_14866,N_14635,N_14468);
nand U14867 (N_14867,N_14594,N_14549);
or U14868 (N_14868,N_14482,N_14631);
nor U14869 (N_14869,N_14449,N_14607);
xor U14870 (N_14870,N_14546,N_14591);
nand U14871 (N_14871,N_14549,N_14677);
and U14872 (N_14872,N_14419,N_14551);
and U14873 (N_14873,N_14593,N_14423);
xor U14874 (N_14874,N_14490,N_14658);
xnor U14875 (N_14875,N_14507,N_14601);
or U14876 (N_14876,N_14653,N_14618);
or U14877 (N_14877,N_14514,N_14605);
or U14878 (N_14878,N_14517,N_14614);
and U14879 (N_14879,N_14653,N_14406);
or U14880 (N_14880,N_14519,N_14682);
nand U14881 (N_14881,N_14602,N_14670);
nor U14882 (N_14882,N_14407,N_14604);
or U14883 (N_14883,N_14547,N_14553);
or U14884 (N_14884,N_14520,N_14521);
nor U14885 (N_14885,N_14665,N_14655);
xnor U14886 (N_14886,N_14444,N_14460);
or U14887 (N_14887,N_14445,N_14412);
nor U14888 (N_14888,N_14444,N_14619);
nand U14889 (N_14889,N_14418,N_14564);
or U14890 (N_14890,N_14422,N_14494);
and U14891 (N_14891,N_14628,N_14680);
and U14892 (N_14892,N_14664,N_14510);
nor U14893 (N_14893,N_14423,N_14601);
xor U14894 (N_14894,N_14552,N_14620);
nand U14895 (N_14895,N_14468,N_14456);
and U14896 (N_14896,N_14674,N_14592);
nor U14897 (N_14897,N_14587,N_14423);
nor U14898 (N_14898,N_14503,N_14406);
nand U14899 (N_14899,N_14513,N_14468);
nor U14900 (N_14900,N_14682,N_14667);
nand U14901 (N_14901,N_14619,N_14560);
nor U14902 (N_14902,N_14609,N_14666);
nand U14903 (N_14903,N_14440,N_14642);
xor U14904 (N_14904,N_14401,N_14417);
nand U14905 (N_14905,N_14546,N_14517);
and U14906 (N_14906,N_14423,N_14461);
or U14907 (N_14907,N_14461,N_14552);
xnor U14908 (N_14908,N_14643,N_14611);
nand U14909 (N_14909,N_14683,N_14446);
xnor U14910 (N_14910,N_14521,N_14559);
or U14911 (N_14911,N_14572,N_14590);
and U14912 (N_14912,N_14588,N_14428);
and U14913 (N_14913,N_14433,N_14441);
and U14914 (N_14914,N_14689,N_14605);
or U14915 (N_14915,N_14650,N_14462);
nor U14916 (N_14916,N_14454,N_14402);
xnor U14917 (N_14917,N_14402,N_14406);
xnor U14918 (N_14918,N_14557,N_14593);
nor U14919 (N_14919,N_14580,N_14512);
nor U14920 (N_14920,N_14662,N_14602);
nor U14921 (N_14921,N_14606,N_14666);
nor U14922 (N_14922,N_14637,N_14467);
nand U14923 (N_14923,N_14690,N_14474);
or U14924 (N_14924,N_14429,N_14591);
nand U14925 (N_14925,N_14542,N_14654);
xnor U14926 (N_14926,N_14536,N_14546);
and U14927 (N_14927,N_14557,N_14625);
xor U14928 (N_14928,N_14513,N_14633);
nand U14929 (N_14929,N_14523,N_14565);
or U14930 (N_14930,N_14489,N_14600);
and U14931 (N_14931,N_14559,N_14645);
and U14932 (N_14932,N_14578,N_14406);
xnor U14933 (N_14933,N_14440,N_14446);
and U14934 (N_14934,N_14621,N_14591);
xnor U14935 (N_14935,N_14533,N_14549);
xor U14936 (N_14936,N_14642,N_14510);
xor U14937 (N_14937,N_14496,N_14553);
nor U14938 (N_14938,N_14682,N_14653);
nand U14939 (N_14939,N_14425,N_14659);
xor U14940 (N_14940,N_14467,N_14478);
or U14941 (N_14941,N_14558,N_14489);
or U14942 (N_14942,N_14641,N_14446);
nand U14943 (N_14943,N_14416,N_14481);
nor U14944 (N_14944,N_14475,N_14698);
or U14945 (N_14945,N_14582,N_14571);
nand U14946 (N_14946,N_14564,N_14561);
xor U14947 (N_14947,N_14578,N_14522);
xor U14948 (N_14948,N_14662,N_14456);
xnor U14949 (N_14949,N_14516,N_14467);
nor U14950 (N_14950,N_14537,N_14503);
nand U14951 (N_14951,N_14518,N_14697);
nand U14952 (N_14952,N_14690,N_14578);
xor U14953 (N_14953,N_14646,N_14501);
nor U14954 (N_14954,N_14559,N_14634);
nor U14955 (N_14955,N_14457,N_14563);
nor U14956 (N_14956,N_14494,N_14519);
xor U14957 (N_14957,N_14466,N_14468);
nand U14958 (N_14958,N_14486,N_14695);
or U14959 (N_14959,N_14522,N_14628);
or U14960 (N_14960,N_14629,N_14435);
or U14961 (N_14961,N_14470,N_14549);
nand U14962 (N_14962,N_14653,N_14622);
or U14963 (N_14963,N_14408,N_14402);
or U14964 (N_14964,N_14489,N_14546);
xnor U14965 (N_14965,N_14635,N_14634);
xnor U14966 (N_14966,N_14524,N_14569);
and U14967 (N_14967,N_14678,N_14610);
or U14968 (N_14968,N_14632,N_14676);
xor U14969 (N_14969,N_14626,N_14678);
nor U14970 (N_14970,N_14469,N_14523);
and U14971 (N_14971,N_14518,N_14473);
and U14972 (N_14972,N_14559,N_14529);
nor U14973 (N_14973,N_14519,N_14572);
nand U14974 (N_14974,N_14634,N_14582);
nand U14975 (N_14975,N_14475,N_14497);
nand U14976 (N_14976,N_14613,N_14697);
or U14977 (N_14977,N_14553,N_14458);
nor U14978 (N_14978,N_14463,N_14480);
nor U14979 (N_14979,N_14460,N_14497);
nand U14980 (N_14980,N_14429,N_14582);
and U14981 (N_14981,N_14446,N_14558);
nand U14982 (N_14982,N_14659,N_14690);
nand U14983 (N_14983,N_14430,N_14470);
xor U14984 (N_14984,N_14512,N_14564);
or U14985 (N_14985,N_14620,N_14476);
or U14986 (N_14986,N_14585,N_14697);
nand U14987 (N_14987,N_14596,N_14465);
xor U14988 (N_14988,N_14401,N_14531);
and U14989 (N_14989,N_14497,N_14485);
nor U14990 (N_14990,N_14645,N_14653);
xor U14991 (N_14991,N_14646,N_14671);
or U14992 (N_14992,N_14442,N_14511);
or U14993 (N_14993,N_14599,N_14537);
and U14994 (N_14994,N_14520,N_14603);
and U14995 (N_14995,N_14435,N_14590);
nand U14996 (N_14996,N_14476,N_14497);
or U14997 (N_14997,N_14464,N_14521);
or U14998 (N_14998,N_14579,N_14559);
nor U14999 (N_14999,N_14637,N_14542);
nand U15000 (N_15000,N_14979,N_14735);
nand U15001 (N_15001,N_14954,N_14950);
xnor U15002 (N_15002,N_14899,N_14888);
nand U15003 (N_15003,N_14732,N_14929);
xnor U15004 (N_15004,N_14860,N_14771);
nand U15005 (N_15005,N_14824,N_14997);
nor U15006 (N_15006,N_14706,N_14948);
nor U15007 (N_15007,N_14985,N_14809);
nand U15008 (N_15008,N_14741,N_14769);
nor U15009 (N_15009,N_14705,N_14756);
nand U15010 (N_15010,N_14907,N_14834);
or U15011 (N_15011,N_14919,N_14920);
nand U15012 (N_15012,N_14845,N_14891);
nor U15013 (N_15013,N_14835,N_14838);
xnor U15014 (N_15014,N_14825,N_14830);
nand U15015 (N_15015,N_14710,N_14990);
nor U15016 (N_15016,N_14731,N_14763);
or U15017 (N_15017,N_14795,N_14962);
nor U15018 (N_15018,N_14799,N_14761);
and U15019 (N_15019,N_14848,N_14903);
and U15020 (N_15020,N_14849,N_14715);
or U15021 (N_15021,N_14945,N_14890);
xor U15022 (N_15022,N_14775,N_14999);
and U15023 (N_15023,N_14952,N_14892);
xnor U15024 (N_15024,N_14882,N_14783);
nand U15025 (N_15025,N_14749,N_14908);
or U15026 (N_15026,N_14802,N_14752);
and U15027 (N_15027,N_14918,N_14730);
xnor U15028 (N_15028,N_14851,N_14955);
and U15029 (N_15029,N_14947,N_14886);
nand U15030 (N_15030,N_14869,N_14837);
nor U15031 (N_15031,N_14737,N_14703);
xnor U15032 (N_15032,N_14711,N_14836);
and U15033 (N_15033,N_14727,N_14844);
nand U15034 (N_15034,N_14957,N_14717);
xnor U15035 (N_15035,N_14826,N_14956);
xnor U15036 (N_15036,N_14906,N_14745);
xor U15037 (N_15037,N_14941,N_14785);
nor U15038 (N_15038,N_14762,N_14718);
or U15039 (N_15039,N_14719,N_14974);
and U15040 (N_15040,N_14966,N_14912);
or U15041 (N_15041,N_14724,N_14819);
nor U15042 (N_15042,N_14855,N_14787);
nor U15043 (N_15043,N_14904,N_14992);
nor U15044 (N_15044,N_14812,N_14884);
xor U15045 (N_15045,N_14807,N_14770);
and U15046 (N_15046,N_14988,N_14782);
or U15047 (N_15047,N_14972,N_14777);
nor U15048 (N_15048,N_14922,N_14895);
or U15049 (N_15049,N_14935,N_14729);
nor U15050 (N_15050,N_14772,N_14924);
nand U15051 (N_15051,N_14900,N_14726);
nor U15052 (N_15052,N_14789,N_14839);
or U15053 (N_15053,N_14712,N_14857);
nand U15054 (N_15054,N_14931,N_14880);
and U15055 (N_15055,N_14949,N_14842);
or U15056 (N_15056,N_14847,N_14934);
xnor U15057 (N_15057,N_14822,N_14865);
or U15058 (N_15058,N_14773,N_14746);
xnor U15059 (N_15059,N_14791,N_14866);
or U15060 (N_15060,N_14821,N_14998);
nand U15061 (N_15061,N_14964,N_14827);
xnor U15062 (N_15062,N_14973,N_14816);
xnor U15063 (N_15063,N_14863,N_14790);
nor U15064 (N_15064,N_14840,N_14722);
and U15065 (N_15065,N_14740,N_14800);
and U15066 (N_15066,N_14960,N_14959);
and U15067 (N_15067,N_14823,N_14833);
and U15068 (N_15068,N_14818,N_14725);
nor U15069 (N_15069,N_14776,N_14905);
xnor U15070 (N_15070,N_14728,N_14750);
xnor U15071 (N_15071,N_14716,N_14971);
or U15072 (N_15072,N_14794,N_14803);
nand U15073 (N_15073,N_14942,N_14909);
xor U15074 (N_15074,N_14798,N_14805);
xor U15075 (N_15075,N_14765,N_14958);
and U15076 (N_15076,N_14780,N_14867);
or U15077 (N_15077,N_14859,N_14961);
and U15078 (N_15078,N_14943,N_14989);
or U15079 (N_15079,N_14792,N_14994);
nand U15080 (N_15080,N_14864,N_14754);
nor U15081 (N_15081,N_14874,N_14878);
nand U15082 (N_15082,N_14829,N_14793);
xor U15083 (N_15083,N_14846,N_14978);
or U15084 (N_15084,N_14817,N_14747);
and U15085 (N_15085,N_14786,N_14877);
nor U15086 (N_15086,N_14797,N_14981);
xor U15087 (N_15087,N_14991,N_14707);
nand U15088 (N_15088,N_14708,N_14963);
nand U15089 (N_15089,N_14755,N_14748);
nor U15090 (N_15090,N_14868,N_14914);
xor U15091 (N_15091,N_14831,N_14781);
and U15092 (N_15092,N_14987,N_14910);
nand U15093 (N_15093,N_14939,N_14977);
xor U15094 (N_15094,N_14744,N_14764);
nand U15095 (N_15095,N_14810,N_14870);
nor U15096 (N_15096,N_14937,N_14925);
xor U15097 (N_15097,N_14739,N_14702);
and U15098 (N_15098,N_14879,N_14940);
nand U15099 (N_15099,N_14967,N_14927);
or U15100 (N_15100,N_14759,N_14933);
or U15101 (N_15101,N_14883,N_14806);
nor U15102 (N_15102,N_14856,N_14861);
or U15103 (N_15103,N_14723,N_14736);
xor U15104 (N_15104,N_14926,N_14928);
or U15105 (N_15105,N_14938,N_14915);
xor U15106 (N_15106,N_14811,N_14815);
nand U15107 (N_15107,N_14982,N_14758);
or U15108 (N_15108,N_14872,N_14862);
nand U15109 (N_15109,N_14808,N_14893);
nand U15110 (N_15110,N_14788,N_14923);
or U15111 (N_15111,N_14841,N_14704);
and U15112 (N_15112,N_14778,N_14986);
or U15113 (N_15113,N_14901,N_14734);
and U15114 (N_15114,N_14995,N_14932);
xnor U15115 (N_15115,N_14944,N_14983);
nand U15116 (N_15116,N_14767,N_14801);
nor U15117 (N_15117,N_14854,N_14733);
and U15118 (N_15118,N_14984,N_14970);
xnor U15119 (N_15119,N_14968,N_14760);
nand U15120 (N_15120,N_14832,N_14738);
nor U15121 (N_15121,N_14796,N_14813);
and U15122 (N_15122,N_14993,N_14898);
and U15123 (N_15123,N_14720,N_14701);
and U15124 (N_15124,N_14743,N_14896);
or U15125 (N_15125,N_14897,N_14885);
and U15126 (N_15126,N_14996,N_14930);
nor U15127 (N_15127,N_14936,N_14881);
or U15128 (N_15128,N_14887,N_14921);
and U15129 (N_15129,N_14875,N_14779);
xor U15130 (N_15130,N_14766,N_14873);
xor U15131 (N_15131,N_14976,N_14913);
and U15132 (N_15132,N_14843,N_14852);
xnor U15133 (N_15133,N_14871,N_14858);
or U15134 (N_15134,N_14853,N_14753);
xor U15135 (N_15135,N_14889,N_14916);
xnor U15136 (N_15136,N_14946,N_14774);
and U15137 (N_15137,N_14804,N_14768);
or U15138 (N_15138,N_14714,N_14700);
nor U15139 (N_15139,N_14721,N_14784);
nor U15140 (N_15140,N_14911,N_14951);
nor U15141 (N_15141,N_14876,N_14980);
and U15142 (N_15142,N_14709,N_14953);
xnor U15143 (N_15143,N_14902,N_14894);
xnor U15144 (N_15144,N_14850,N_14975);
nand U15145 (N_15145,N_14742,N_14828);
nor U15146 (N_15146,N_14713,N_14969);
or U15147 (N_15147,N_14757,N_14965);
nor U15148 (N_15148,N_14917,N_14751);
xor U15149 (N_15149,N_14814,N_14820);
nand U15150 (N_15150,N_14935,N_14841);
nor U15151 (N_15151,N_14970,N_14961);
or U15152 (N_15152,N_14820,N_14733);
nor U15153 (N_15153,N_14729,N_14865);
nand U15154 (N_15154,N_14704,N_14927);
or U15155 (N_15155,N_14767,N_14831);
xnor U15156 (N_15156,N_14917,N_14919);
nor U15157 (N_15157,N_14889,N_14988);
xor U15158 (N_15158,N_14764,N_14858);
nor U15159 (N_15159,N_14722,N_14702);
and U15160 (N_15160,N_14798,N_14833);
nor U15161 (N_15161,N_14895,N_14872);
nand U15162 (N_15162,N_14891,N_14894);
xor U15163 (N_15163,N_14917,N_14958);
xor U15164 (N_15164,N_14811,N_14849);
and U15165 (N_15165,N_14851,N_14735);
nor U15166 (N_15166,N_14962,N_14952);
nor U15167 (N_15167,N_14791,N_14995);
nor U15168 (N_15168,N_14914,N_14940);
or U15169 (N_15169,N_14723,N_14968);
nor U15170 (N_15170,N_14955,N_14945);
nor U15171 (N_15171,N_14803,N_14768);
nand U15172 (N_15172,N_14861,N_14969);
or U15173 (N_15173,N_14879,N_14812);
xor U15174 (N_15174,N_14748,N_14708);
nand U15175 (N_15175,N_14738,N_14877);
xnor U15176 (N_15176,N_14705,N_14807);
nand U15177 (N_15177,N_14857,N_14913);
and U15178 (N_15178,N_14919,N_14735);
or U15179 (N_15179,N_14805,N_14741);
nor U15180 (N_15180,N_14874,N_14908);
nor U15181 (N_15181,N_14882,N_14819);
and U15182 (N_15182,N_14922,N_14882);
or U15183 (N_15183,N_14723,N_14977);
or U15184 (N_15184,N_14795,N_14924);
and U15185 (N_15185,N_14712,N_14764);
nor U15186 (N_15186,N_14735,N_14881);
or U15187 (N_15187,N_14906,N_14782);
or U15188 (N_15188,N_14962,N_14981);
or U15189 (N_15189,N_14916,N_14956);
nor U15190 (N_15190,N_14873,N_14965);
nand U15191 (N_15191,N_14741,N_14772);
nand U15192 (N_15192,N_14702,N_14830);
xnor U15193 (N_15193,N_14950,N_14896);
nor U15194 (N_15194,N_14703,N_14883);
nor U15195 (N_15195,N_14833,N_14723);
nor U15196 (N_15196,N_14855,N_14836);
nand U15197 (N_15197,N_14839,N_14960);
and U15198 (N_15198,N_14961,N_14936);
xor U15199 (N_15199,N_14961,N_14751);
xor U15200 (N_15200,N_14861,N_14821);
and U15201 (N_15201,N_14739,N_14991);
or U15202 (N_15202,N_14974,N_14910);
nand U15203 (N_15203,N_14968,N_14925);
nor U15204 (N_15204,N_14854,N_14895);
or U15205 (N_15205,N_14756,N_14972);
or U15206 (N_15206,N_14834,N_14731);
or U15207 (N_15207,N_14866,N_14749);
and U15208 (N_15208,N_14954,N_14707);
nor U15209 (N_15209,N_14967,N_14892);
or U15210 (N_15210,N_14924,N_14763);
nor U15211 (N_15211,N_14841,N_14967);
nor U15212 (N_15212,N_14879,N_14739);
nor U15213 (N_15213,N_14759,N_14997);
xnor U15214 (N_15214,N_14808,N_14944);
nor U15215 (N_15215,N_14790,N_14779);
nor U15216 (N_15216,N_14918,N_14810);
nor U15217 (N_15217,N_14946,N_14920);
or U15218 (N_15218,N_14843,N_14993);
and U15219 (N_15219,N_14918,N_14716);
nor U15220 (N_15220,N_14800,N_14761);
nor U15221 (N_15221,N_14884,N_14824);
nor U15222 (N_15222,N_14824,N_14748);
nor U15223 (N_15223,N_14998,N_14829);
xnor U15224 (N_15224,N_14780,N_14869);
nor U15225 (N_15225,N_14840,N_14828);
nand U15226 (N_15226,N_14929,N_14968);
xor U15227 (N_15227,N_14788,N_14939);
and U15228 (N_15228,N_14959,N_14833);
or U15229 (N_15229,N_14944,N_14707);
and U15230 (N_15230,N_14994,N_14703);
or U15231 (N_15231,N_14975,N_14961);
nor U15232 (N_15232,N_14872,N_14917);
nand U15233 (N_15233,N_14932,N_14832);
and U15234 (N_15234,N_14939,N_14774);
nand U15235 (N_15235,N_14756,N_14741);
nor U15236 (N_15236,N_14895,N_14765);
nand U15237 (N_15237,N_14979,N_14967);
or U15238 (N_15238,N_14843,N_14913);
and U15239 (N_15239,N_14875,N_14909);
xnor U15240 (N_15240,N_14796,N_14823);
and U15241 (N_15241,N_14919,N_14734);
xor U15242 (N_15242,N_14811,N_14892);
nor U15243 (N_15243,N_14904,N_14729);
xor U15244 (N_15244,N_14704,N_14871);
nor U15245 (N_15245,N_14943,N_14792);
and U15246 (N_15246,N_14956,N_14796);
or U15247 (N_15247,N_14755,N_14818);
and U15248 (N_15248,N_14821,N_14700);
nor U15249 (N_15249,N_14728,N_14710);
and U15250 (N_15250,N_14949,N_14804);
nor U15251 (N_15251,N_14888,N_14802);
nor U15252 (N_15252,N_14984,N_14852);
nand U15253 (N_15253,N_14978,N_14794);
nand U15254 (N_15254,N_14791,N_14794);
xor U15255 (N_15255,N_14919,N_14954);
xor U15256 (N_15256,N_14864,N_14866);
or U15257 (N_15257,N_14956,N_14729);
nand U15258 (N_15258,N_14783,N_14842);
nand U15259 (N_15259,N_14898,N_14906);
or U15260 (N_15260,N_14710,N_14821);
nor U15261 (N_15261,N_14900,N_14791);
xor U15262 (N_15262,N_14988,N_14906);
and U15263 (N_15263,N_14943,N_14912);
or U15264 (N_15264,N_14960,N_14730);
or U15265 (N_15265,N_14997,N_14833);
xor U15266 (N_15266,N_14818,N_14809);
xor U15267 (N_15267,N_14816,N_14969);
nor U15268 (N_15268,N_14908,N_14921);
or U15269 (N_15269,N_14948,N_14789);
and U15270 (N_15270,N_14997,N_14725);
nand U15271 (N_15271,N_14945,N_14970);
xnor U15272 (N_15272,N_14839,N_14761);
nand U15273 (N_15273,N_14768,N_14767);
nor U15274 (N_15274,N_14820,N_14830);
and U15275 (N_15275,N_14885,N_14874);
nand U15276 (N_15276,N_14904,N_14974);
and U15277 (N_15277,N_14857,N_14819);
and U15278 (N_15278,N_14927,N_14847);
xnor U15279 (N_15279,N_14956,N_14752);
nand U15280 (N_15280,N_14794,N_14936);
nand U15281 (N_15281,N_14942,N_14887);
xor U15282 (N_15282,N_14767,N_14808);
and U15283 (N_15283,N_14779,N_14887);
or U15284 (N_15284,N_14969,N_14806);
xnor U15285 (N_15285,N_14964,N_14982);
or U15286 (N_15286,N_14853,N_14914);
and U15287 (N_15287,N_14859,N_14918);
nor U15288 (N_15288,N_14816,N_14925);
and U15289 (N_15289,N_14885,N_14816);
nand U15290 (N_15290,N_14763,N_14971);
or U15291 (N_15291,N_14805,N_14996);
nand U15292 (N_15292,N_14829,N_14894);
nor U15293 (N_15293,N_14755,N_14996);
and U15294 (N_15294,N_14847,N_14911);
nor U15295 (N_15295,N_14809,N_14794);
nand U15296 (N_15296,N_14973,N_14782);
xnor U15297 (N_15297,N_14867,N_14984);
nor U15298 (N_15298,N_14991,N_14839);
nor U15299 (N_15299,N_14890,N_14750);
and U15300 (N_15300,N_15137,N_15130);
xor U15301 (N_15301,N_15049,N_15093);
nor U15302 (N_15302,N_15138,N_15239);
nor U15303 (N_15303,N_15105,N_15293);
and U15304 (N_15304,N_15210,N_15025);
nand U15305 (N_15305,N_15221,N_15023);
and U15306 (N_15306,N_15046,N_15186);
or U15307 (N_15307,N_15296,N_15043);
nor U15308 (N_15308,N_15042,N_15298);
and U15309 (N_15309,N_15036,N_15124);
or U15310 (N_15310,N_15035,N_15057);
and U15311 (N_15311,N_15151,N_15041);
xor U15312 (N_15312,N_15085,N_15242);
nor U15313 (N_15313,N_15155,N_15224);
nor U15314 (N_15314,N_15121,N_15022);
xnor U15315 (N_15315,N_15034,N_15095);
nand U15316 (N_15316,N_15084,N_15238);
and U15317 (N_15317,N_15040,N_15149);
xor U15318 (N_15318,N_15012,N_15253);
nor U15319 (N_15319,N_15286,N_15191);
nor U15320 (N_15320,N_15166,N_15249);
and U15321 (N_15321,N_15052,N_15164);
nor U15322 (N_15322,N_15099,N_15157);
or U15323 (N_15323,N_15182,N_15258);
and U15324 (N_15324,N_15010,N_15196);
xor U15325 (N_15325,N_15156,N_15181);
nor U15326 (N_15326,N_15113,N_15280);
or U15327 (N_15327,N_15171,N_15047);
xor U15328 (N_15328,N_15063,N_15014);
nand U15329 (N_15329,N_15226,N_15159);
nor U15330 (N_15330,N_15100,N_15172);
nand U15331 (N_15331,N_15220,N_15015);
and U15332 (N_15332,N_15295,N_15208);
and U15333 (N_15333,N_15020,N_15179);
or U15334 (N_15334,N_15077,N_15021);
nand U15335 (N_15335,N_15068,N_15125);
and U15336 (N_15336,N_15118,N_15045);
nand U15337 (N_15337,N_15053,N_15235);
and U15338 (N_15338,N_15076,N_15120);
or U15339 (N_15339,N_15061,N_15292);
nand U15340 (N_15340,N_15225,N_15051);
nor U15341 (N_15341,N_15204,N_15203);
nand U15342 (N_15342,N_15176,N_15227);
and U15343 (N_15343,N_15122,N_15002);
nor U15344 (N_15344,N_15223,N_15097);
xor U15345 (N_15345,N_15163,N_15001);
xor U15346 (N_15346,N_15038,N_15144);
nand U15347 (N_15347,N_15107,N_15200);
or U15348 (N_15348,N_15029,N_15205);
nor U15349 (N_15349,N_15216,N_15008);
nand U15350 (N_15350,N_15165,N_15028);
nor U15351 (N_15351,N_15202,N_15212);
xnor U15352 (N_15352,N_15073,N_15246);
and U15353 (N_15353,N_15274,N_15044);
nor U15354 (N_15354,N_15116,N_15005);
xor U15355 (N_15355,N_15148,N_15050);
nand U15356 (N_15356,N_15269,N_15267);
xor U15357 (N_15357,N_15161,N_15016);
nand U15358 (N_15358,N_15090,N_15132);
xor U15359 (N_15359,N_15140,N_15263);
nor U15360 (N_15360,N_15079,N_15187);
or U15361 (N_15361,N_15290,N_15078);
xnor U15362 (N_15362,N_15135,N_15234);
nand U15363 (N_15363,N_15072,N_15070);
nor U15364 (N_15364,N_15123,N_15217);
nor U15365 (N_15365,N_15129,N_15284);
or U15366 (N_15366,N_15056,N_15260);
nor U15367 (N_15367,N_15106,N_15201);
and U15368 (N_15368,N_15244,N_15141);
nor U15369 (N_15369,N_15257,N_15154);
or U15370 (N_15370,N_15261,N_15011);
nand U15371 (N_15371,N_15169,N_15145);
or U15372 (N_15372,N_15264,N_15188);
xnor U15373 (N_15373,N_15207,N_15000);
nand U15374 (N_15374,N_15102,N_15117);
nand U15375 (N_15375,N_15229,N_15233);
nor U15376 (N_15376,N_15126,N_15180);
nor U15377 (N_15377,N_15013,N_15215);
nand U15378 (N_15378,N_15174,N_15031);
and U15379 (N_15379,N_15143,N_15197);
xnor U15380 (N_15380,N_15009,N_15218);
nand U15381 (N_15381,N_15237,N_15245);
or U15382 (N_15382,N_15066,N_15147);
xnor U15383 (N_15383,N_15259,N_15199);
xnor U15384 (N_15384,N_15092,N_15183);
xor U15385 (N_15385,N_15003,N_15048);
nor U15386 (N_15386,N_15167,N_15252);
nand U15387 (N_15387,N_15030,N_15110);
and U15388 (N_15388,N_15243,N_15065);
nand U15389 (N_15389,N_15026,N_15168);
xor U15390 (N_15390,N_15039,N_15024);
nand U15391 (N_15391,N_15091,N_15089);
or U15392 (N_15392,N_15146,N_15104);
xnor U15393 (N_15393,N_15254,N_15268);
nor U15394 (N_15394,N_15271,N_15185);
nor U15395 (N_15395,N_15279,N_15094);
xor U15396 (N_15396,N_15081,N_15131);
nand U15397 (N_15397,N_15178,N_15230);
and U15398 (N_15398,N_15037,N_15285);
or U15399 (N_15399,N_15228,N_15236);
nand U15400 (N_15400,N_15266,N_15272);
nor U15401 (N_15401,N_15004,N_15251);
xnor U15402 (N_15402,N_15075,N_15289);
nor U15403 (N_15403,N_15069,N_15067);
nor U15404 (N_15404,N_15294,N_15017);
or U15405 (N_15405,N_15192,N_15250);
nand U15406 (N_15406,N_15139,N_15096);
and U15407 (N_15407,N_15111,N_15153);
nand U15408 (N_15408,N_15101,N_15214);
nor U15409 (N_15409,N_15232,N_15195);
or U15410 (N_15410,N_15219,N_15086);
and U15411 (N_15411,N_15006,N_15276);
and U15412 (N_15412,N_15241,N_15060);
xor U15413 (N_15413,N_15150,N_15213);
nor U15414 (N_15414,N_15198,N_15128);
nand U15415 (N_15415,N_15184,N_15209);
or U15416 (N_15416,N_15082,N_15206);
and U15417 (N_15417,N_15055,N_15278);
nor U15418 (N_15418,N_15062,N_15297);
nand U15419 (N_15419,N_15032,N_15098);
and U15420 (N_15420,N_15288,N_15064);
xnor U15421 (N_15421,N_15287,N_15255);
xnor U15422 (N_15422,N_15087,N_15194);
and U15423 (N_15423,N_15019,N_15283);
nand U15424 (N_15424,N_15222,N_15054);
nand U15425 (N_15425,N_15231,N_15136);
nor U15426 (N_15426,N_15127,N_15211);
and U15427 (N_15427,N_15262,N_15265);
nor U15428 (N_15428,N_15281,N_15248);
xor U15429 (N_15429,N_15173,N_15175);
or U15430 (N_15430,N_15119,N_15299);
xnor U15431 (N_15431,N_15074,N_15112);
nor U15432 (N_15432,N_15088,N_15142);
or U15433 (N_15433,N_15058,N_15115);
and U15434 (N_15434,N_15160,N_15275);
or U15435 (N_15435,N_15133,N_15162);
or U15436 (N_15436,N_15273,N_15193);
and U15437 (N_15437,N_15270,N_15018);
xnor U15438 (N_15438,N_15134,N_15083);
and U15439 (N_15439,N_15033,N_15007);
xnor U15440 (N_15440,N_15109,N_15108);
nor U15441 (N_15441,N_15152,N_15170);
and U15442 (N_15442,N_15158,N_15059);
nor U15443 (N_15443,N_15247,N_15071);
or U15444 (N_15444,N_15114,N_15282);
or U15445 (N_15445,N_15291,N_15190);
xor U15446 (N_15446,N_15080,N_15027);
nor U15447 (N_15447,N_15177,N_15240);
and U15448 (N_15448,N_15256,N_15277);
xnor U15449 (N_15449,N_15189,N_15103);
nor U15450 (N_15450,N_15016,N_15285);
and U15451 (N_15451,N_15001,N_15222);
or U15452 (N_15452,N_15220,N_15144);
and U15453 (N_15453,N_15013,N_15107);
or U15454 (N_15454,N_15287,N_15177);
and U15455 (N_15455,N_15223,N_15273);
nand U15456 (N_15456,N_15209,N_15201);
nor U15457 (N_15457,N_15148,N_15062);
or U15458 (N_15458,N_15038,N_15181);
nor U15459 (N_15459,N_15006,N_15102);
xor U15460 (N_15460,N_15129,N_15204);
or U15461 (N_15461,N_15057,N_15013);
nor U15462 (N_15462,N_15205,N_15145);
or U15463 (N_15463,N_15170,N_15109);
nand U15464 (N_15464,N_15248,N_15159);
and U15465 (N_15465,N_15046,N_15229);
xor U15466 (N_15466,N_15217,N_15269);
xnor U15467 (N_15467,N_15098,N_15058);
or U15468 (N_15468,N_15129,N_15159);
nand U15469 (N_15469,N_15130,N_15064);
nand U15470 (N_15470,N_15027,N_15111);
and U15471 (N_15471,N_15236,N_15208);
xnor U15472 (N_15472,N_15257,N_15049);
xnor U15473 (N_15473,N_15151,N_15093);
or U15474 (N_15474,N_15222,N_15152);
xor U15475 (N_15475,N_15006,N_15047);
nor U15476 (N_15476,N_15045,N_15088);
nand U15477 (N_15477,N_15172,N_15010);
or U15478 (N_15478,N_15278,N_15033);
and U15479 (N_15479,N_15298,N_15017);
xnor U15480 (N_15480,N_15035,N_15124);
nand U15481 (N_15481,N_15262,N_15289);
xnor U15482 (N_15482,N_15137,N_15003);
and U15483 (N_15483,N_15274,N_15105);
or U15484 (N_15484,N_15289,N_15217);
and U15485 (N_15485,N_15011,N_15259);
nor U15486 (N_15486,N_15277,N_15163);
and U15487 (N_15487,N_15032,N_15183);
xnor U15488 (N_15488,N_15231,N_15236);
nand U15489 (N_15489,N_15265,N_15016);
xnor U15490 (N_15490,N_15032,N_15071);
xor U15491 (N_15491,N_15015,N_15073);
nor U15492 (N_15492,N_15069,N_15164);
or U15493 (N_15493,N_15141,N_15053);
or U15494 (N_15494,N_15005,N_15000);
nor U15495 (N_15495,N_15035,N_15157);
xor U15496 (N_15496,N_15212,N_15222);
xnor U15497 (N_15497,N_15064,N_15052);
and U15498 (N_15498,N_15094,N_15026);
nand U15499 (N_15499,N_15032,N_15087);
nor U15500 (N_15500,N_15243,N_15091);
and U15501 (N_15501,N_15272,N_15275);
xor U15502 (N_15502,N_15142,N_15117);
nor U15503 (N_15503,N_15257,N_15040);
and U15504 (N_15504,N_15249,N_15093);
or U15505 (N_15505,N_15239,N_15036);
and U15506 (N_15506,N_15195,N_15127);
or U15507 (N_15507,N_15207,N_15113);
or U15508 (N_15508,N_15006,N_15148);
nor U15509 (N_15509,N_15071,N_15078);
or U15510 (N_15510,N_15106,N_15046);
or U15511 (N_15511,N_15013,N_15182);
nor U15512 (N_15512,N_15273,N_15136);
nand U15513 (N_15513,N_15135,N_15047);
or U15514 (N_15514,N_15261,N_15236);
xnor U15515 (N_15515,N_15130,N_15089);
and U15516 (N_15516,N_15173,N_15259);
nor U15517 (N_15517,N_15195,N_15125);
nand U15518 (N_15518,N_15019,N_15095);
nand U15519 (N_15519,N_15224,N_15241);
or U15520 (N_15520,N_15157,N_15160);
or U15521 (N_15521,N_15227,N_15107);
and U15522 (N_15522,N_15157,N_15240);
and U15523 (N_15523,N_15249,N_15042);
nand U15524 (N_15524,N_15168,N_15240);
xor U15525 (N_15525,N_15055,N_15051);
nand U15526 (N_15526,N_15266,N_15146);
nand U15527 (N_15527,N_15013,N_15117);
or U15528 (N_15528,N_15199,N_15072);
xor U15529 (N_15529,N_15073,N_15112);
or U15530 (N_15530,N_15115,N_15214);
nor U15531 (N_15531,N_15296,N_15107);
xor U15532 (N_15532,N_15237,N_15214);
and U15533 (N_15533,N_15277,N_15071);
nor U15534 (N_15534,N_15082,N_15248);
xor U15535 (N_15535,N_15143,N_15080);
and U15536 (N_15536,N_15087,N_15176);
or U15537 (N_15537,N_15251,N_15034);
nand U15538 (N_15538,N_15158,N_15090);
and U15539 (N_15539,N_15205,N_15287);
and U15540 (N_15540,N_15160,N_15056);
nand U15541 (N_15541,N_15023,N_15197);
nand U15542 (N_15542,N_15116,N_15014);
xnor U15543 (N_15543,N_15052,N_15115);
nand U15544 (N_15544,N_15105,N_15199);
or U15545 (N_15545,N_15210,N_15202);
nand U15546 (N_15546,N_15114,N_15039);
xor U15547 (N_15547,N_15261,N_15170);
nand U15548 (N_15548,N_15014,N_15195);
nor U15549 (N_15549,N_15184,N_15119);
xnor U15550 (N_15550,N_15136,N_15024);
or U15551 (N_15551,N_15187,N_15006);
xor U15552 (N_15552,N_15142,N_15091);
nand U15553 (N_15553,N_15070,N_15058);
and U15554 (N_15554,N_15056,N_15077);
nor U15555 (N_15555,N_15008,N_15255);
nand U15556 (N_15556,N_15115,N_15109);
and U15557 (N_15557,N_15056,N_15154);
nand U15558 (N_15558,N_15069,N_15024);
or U15559 (N_15559,N_15148,N_15048);
nand U15560 (N_15560,N_15105,N_15092);
xor U15561 (N_15561,N_15268,N_15150);
or U15562 (N_15562,N_15050,N_15291);
xor U15563 (N_15563,N_15176,N_15085);
and U15564 (N_15564,N_15032,N_15113);
or U15565 (N_15565,N_15233,N_15012);
or U15566 (N_15566,N_15193,N_15261);
nand U15567 (N_15567,N_15290,N_15136);
and U15568 (N_15568,N_15209,N_15137);
nand U15569 (N_15569,N_15207,N_15293);
nor U15570 (N_15570,N_15260,N_15022);
and U15571 (N_15571,N_15154,N_15222);
and U15572 (N_15572,N_15299,N_15232);
and U15573 (N_15573,N_15078,N_15052);
nor U15574 (N_15574,N_15083,N_15228);
nand U15575 (N_15575,N_15278,N_15035);
and U15576 (N_15576,N_15041,N_15244);
and U15577 (N_15577,N_15073,N_15250);
or U15578 (N_15578,N_15264,N_15000);
nor U15579 (N_15579,N_15240,N_15211);
xor U15580 (N_15580,N_15152,N_15025);
and U15581 (N_15581,N_15254,N_15067);
nand U15582 (N_15582,N_15250,N_15075);
nor U15583 (N_15583,N_15087,N_15156);
and U15584 (N_15584,N_15016,N_15296);
nor U15585 (N_15585,N_15263,N_15111);
and U15586 (N_15586,N_15080,N_15147);
nor U15587 (N_15587,N_15113,N_15205);
nand U15588 (N_15588,N_15210,N_15178);
nor U15589 (N_15589,N_15246,N_15227);
nor U15590 (N_15590,N_15237,N_15117);
and U15591 (N_15591,N_15263,N_15240);
and U15592 (N_15592,N_15130,N_15097);
xor U15593 (N_15593,N_15089,N_15251);
xor U15594 (N_15594,N_15054,N_15269);
or U15595 (N_15595,N_15176,N_15196);
or U15596 (N_15596,N_15077,N_15146);
nor U15597 (N_15597,N_15091,N_15057);
xor U15598 (N_15598,N_15166,N_15065);
xor U15599 (N_15599,N_15162,N_15243);
xnor U15600 (N_15600,N_15570,N_15358);
nand U15601 (N_15601,N_15306,N_15557);
xor U15602 (N_15602,N_15443,N_15513);
or U15603 (N_15603,N_15559,N_15548);
xnor U15604 (N_15604,N_15477,N_15446);
and U15605 (N_15605,N_15307,N_15410);
or U15606 (N_15606,N_15532,N_15414);
nand U15607 (N_15607,N_15480,N_15310);
nand U15608 (N_15608,N_15500,N_15497);
nor U15609 (N_15609,N_15552,N_15555);
and U15610 (N_15610,N_15538,N_15567);
xor U15611 (N_15611,N_15541,N_15531);
xnor U15612 (N_15612,N_15578,N_15479);
or U15613 (N_15613,N_15396,N_15471);
xor U15614 (N_15614,N_15543,N_15346);
and U15615 (N_15615,N_15515,N_15335);
nand U15616 (N_15616,N_15388,N_15330);
or U15617 (N_15617,N_15431,N_15326);
nand U15618 (N_15618,N_15438,N_15361);
and U15619 (N_15619,N_15577,N_15353);
xor U15620 (N_15620,N_15485,N_15405);
or U15621 (N_15621,N_15328,N_15572);
nor U15622 (N_15622,N_15490,N_15436);
or U15623 (N_15623,N_15394,N_15322);
xor U15624 (N_15624,N_15305,N_15539);
nand U15625 (N_15625,N_15544,N_15599);
and U15626 (N_15626,N_15375,N_15434);
nor U15627 (N_15627,N_15586,N_15393);
xor U15628 (N_15628,N_15558,N_15579);
nand U15629 (N_15629,N_15366,N_15426);
nand U15630 (N_15630,N_15549,N_15516);
and U15631 (N_15631,N_15424,N_15568);
xor U15632 (N_15632,N_15491,N_15444);
xnor U15633 (N_15633,N_15342,N_15464);
nand U15634 (N_15634,N_15536,N_15598);
nand U15635 (N_15635,N_15506,N_15311);
nand U15636 (N_15636,N_15360,N_15593);
nor U15637 (N_15637,N_15364,N_15576);
and U15638 (N_15638,N_15380,N_15357);
nand U15639 (N_15639,N_15560,N_15537);
or U15640 (N_15640,N_15404,N_15408);
and U15641 (N_15641,N_15507,N_15574);
and U15642 (N_15642,N_15407,N_15439);
nand U15643 (N_15643,N_15460,N_15527);
or U15644 (N_15644,N_15587,N_15419);
xor U15645 (N_15645,N_15300,N_15590);
or U15646 (N_15646,N_15522,N_15533);
and U15647 (N_15647,N_15502,N_15542);
and U15648 (N_15648,N_15376,N_15337);
xnor U15649 (N_15649,N_15331,N_15417);
nand U15650 (N_15650,N_15525,N_15403);
nand U15651 (N_15651,N_15445,N_15463);
nor U15652 (N_15652,N_15535,N_15324);
and U15653 (N_15653,N_15496,N_15428);
xnor U15654 (N_15654,N_15315,N_15321);
nor U15655 (N_15655,N_15546,N_15530);
xor U15656 (N_15656,N_15588,N_15529);
xnor U15657 (N_15657,N_15571,N_15447);
nor U15658 (N_15658,N_15493,N_15453);
xor U15659 (N_15659,N_15523,N_15488);
nor U15660 (N_15660,N_15483,N_15473);
and U15661 (N_15661,N_15442,N_15482);
and U15662 (N_15662,N_15378,N_15427);
or U15663 (N_15663,N_15470,N_15458);
nor U15664 (N_15664,N_15467,N_15333);
and U15665 (N_15665,N_15459,N_15401);
nor U15666 (N_15666,N_15309,N_15341);
nand U15667 (N_15667,N_15468,N_15524);
nor U15668 (N_15668,N_15416,N_15415);
or U15669 (N_15669,N_15429,N_15499);
nand U15670 (N_15670,N_15316,N_15301);
and U15671 (N_15671,N_15484,N_15303);
nand U15672 (N_15672,N_15320,N_15374);
or U15673 (N_15673,N_15583,N_15481);
xnor U15674 (N_15674,N_15349,N_15440);
nor U15675 (N_15675,N_15503,N_15461);
nand U15676 (N_15676,N_15457,N_15319);
and U15677 (N_15677,N_15462,N_15545);
or U15678 (N_15678,N_15494,N_15505);
nor U15679 (N_15679,N_15356,N_15379);
or U15680 (N_15680,N_15421,N_15489);
and U15681 (N_15681,N_15314,N_15413);
or U15682 (N_15682,N_15465,N_15399);
xnor U15683 (N_15683,N_15302,N_15308);
or U15684 (N_15684,N_15504,N_15352);
and U15685 (N_15685,N_15372,N_15580);
nand U15686 (N_15686,N_15382,N_15350);
xor U15687 (N_15687,N_15359,N_15565);
nor U15688 (N_15688,N_15562,N_15492);
xnor U15689 (N_15689,N_15486,N_15400);
or U15690 (N_15690,N_15345,N_15534);
nand U15691 (N_15691,N_15581,N_15566);
nor U15692 (N_15692,N_15435,N_15540);
or U15693 (N_15693,N_15390,N_15386);
xnor U15694 (N_15694,N_15433,N_15367);
or U15695 (N_15695,N_15449,N_15550);
nand U15696 (N_15696,N_15441,N_15409);
and U15697 (N_15697,N_15547,N_15313);
nand U15698 (N_15698,N_15348,N_15595);
and U15699 (N_15699,N_15475,N_15430);
nor U15700 (N_15700,N_15343,N_15591);
nor U15701 (N_15701,N_15383,N_15519);
xnor U15702 (N_15702,N_15406,N_15354);
nand U15703 (N_15703,N_15392,N_15318);
xor U15704 (N_15704,N_15385,N_15371);
and U15705 (N_15705,N_15355,N_15312);
nor U15706 (N_15706,N_15338,N_15368);
and U15707 (N_15707,N_15423,N_15365);
nor U15708 (N_15708,N_15323,N_15336);
and U15709 (N_15709,N_15589,N_15594);
or U15710 (N_15710,N_15554,N_15329);
or U15711 (N_15711,N_15373,N_15450);
nor U15712 (N_15712,N_15437,N_15397);
and U15713 (N_15713,N_15597,N_15425);
or U15714 (N_15714,N_15569,N_15452);
nand U15715 (N_15715,N_15448,N_15454);
nor U15716 (N_15716,N_15398,N_15487);
nor U15717 (N_15717,N_15528,N_15432);
nand U15718 (N_15718,N_15317,N_15402);
or U15719 (N_15719,N_15327,N_15469);
nand U15720 (N_15720,N_15512,N_15521);
nor U15721 (N_15721,N_15381,N_15478);
nand U15722 (N_15722,N_15418,N_15575);
or U15723 (N_15723,N_15395,N_15369);
or U15724 (N_15724,N_15377,N_15564);
nand U15725 (N_15725,N_15455,N_15362);
and U15726 (N_15726,N_15514,N_15476);
xor U15727 (N_15727,N_15551,N_15518);
nand U15728 (N_15728,N_15553,N_15420);
and U15729 (N_15729,N_15340,N_15495);
nand U15730 (N_15730,N_15501,N_15389);
and U15731 (N_15731,N_15384,N_15509);
or U15732 (N_15732,N_15474,N_15344);
nand U15733 (N_15733,N_15582,N_15387);
and U15734 (N_15734,N_15584,N_15466);
or U15735 (N_15735,N_15573,N_15370);
and U15736 (N_15736,N_15561,N_15325);
and U15737 (N_15737,N_15510,N_15391);
nor U15738 (N_15738,N_15334,N_15556);
or U15739 (N_15739,N_15347,N_15451);
and U15740 (N_15740,N_15472,N_15339);
nor U15741 (N_15741,N_15563,N_15332);
and U15742 (N_15742,N_15526,N_15596);
nor U15743 (N_15743,N_15363,N_15592);
or U15744 (N_15744,N_15517,N_15456);
nand U15745 (N_15745,N_15304,N_15351);
and U15746 (N_15746,N_15422,N_15508);
xor U15747 (N_15747,N_15520,N_15585);
and U15748 (N_15748,N_15412,N_15498);
xnor U15749 (N_15749,N_15411,N_15511);
and U15750 (N_15750,N_15331,N_15518);
or U15751 (N_15751,N_15557,N_15552);
xnor U15752 (N_15752,N_15445,N_15594);
or U15753 (N_15753,N_15517,N_15349);
nor U15754 (N_15754,N_15508,N_15386);
xor U15755 (N_15755,N_15567,N_15395);
nor U15756 (N_15756,N_15489,N_15525);
or U15757 (N_15757,N_15569,N_15559);
and U15758 (N_15758,N_15304,N_15332);
nor U15759 (N_15759,N_15583,N_15360);
and U15760 (N_15760,N_15446,N_15343);
nand U15761 (N_15761,N_15335,N_15398);
nor U15762 (N_15762,N_15324,N_15311);
nor U15763 (N_15763,N_15424,N_15552);
and U15764 (N_15764,N_15415,N_15322);
and U15765 (N_15765,N_15559,N_15570);
and U15766 (N_15766,N_15447,N_15360);
nand U15767 (N_15767,N_15318,N_15477);
nor U15768 (N_15768,N_15570,N_15496);
xnor U15769 (N_15769,N_15311,N_15352);
and U15770 (N_15770,N_15539,N_15495);
nor U15771 (N_15771,N_15343,N_15482);
xor U15772 (N_15772,N_15487,N_15515);
or U15773 (N_15773,N_15426,N_15494);
or U15774 (N_15774,N_15516,N_15384);
nand U15775 (N_15775,N_15512,N_15427);
xnor U15776 (N_15776,N_15407,N_15370);
xor U15777 (N_15777,N_15533,N_15458);
nor U15778 (N_15778,N_15488,N_15412);
nor U15779 (N_15779,N_15566,N_15543);
xor U15780 (N_15780,N_15537,N_15596);
or U15781 (N_15781,N_15531,N_15413);
nand U15782 (N_15782,N_15327,N_15426);
nor U15783 (N_15783,N_15309,N_15586);
nand U15784 (N_15784,N_15329,N_15330);
xnor U15785 (N_15785,N_15485,N_15458);
nand U15786 (N_15786,N_15411,N_15545);
or U15787 (N_15787,N_15447,N_15490);
nor U15788 (N_15788,N_15320,N_15400);
nand U15789 (N_15789,N_15456,N_15447);
xor U15790 (N_15790,N_15308,N_15566);
nor U15791 (N_15791,N_15373,N_15370);
nand U15792 (N_15792,N_15307,N_15543);
nor U15793 (N_15793,N_15535,N_15454);
xnor U15794 (N_15794,N_15535,N_15493);
xor U15795 (N_15795,N_15441,N_15430);
xnor U15796 (N_15796,N_15346,N_15541);
xor U15797 (N_15797,N_15504,N_15518);
nand U15798 (N_15798,N_15554,N_15305);
nand U15799 (N_15799,N_15441,N_15540);
nor U15800 (N_15800,N_15346,N_15556);
nor U15801 (N_15801,N_15332,N_15493);
and U15802 (N_15802,N_15498,N_15416);
nor U15803 (N_15803,N_15368,N_15599);
nor U15804 (N_15804,N_15434,N_15566);
or U15805 (N_15805,N_15395,N_15451);
or U15806 (N_15806,N_15346,N_15517);
nor U15807 (N_15807,N_15306,N_15438);
and U15808 (N_15808,N_15546,N_15488);
nand U15809 (N_15809,N_15543,N_15460);
or U15810 (N_15810,N_15307,N_15596);
xor U15811 (N_15811,N_15488,N_15365);
xnor U15812 (N_15812,N_15406,N_15421);
xnor U15813 (N_15813,N_15574,N_15321);
xor U15814 (N_15814,N_15588,N_15330);
and U15815 (N_15815,N_15346,N_15398);
xnor U15816 (N_15816,N_15538,N_15464);
nor U15817 (N_15817,N_15340,N_15380);
and U15818 (N_15818,N_15445,N_15501);
or U15819 (N_15819,N_15401,N_15325);
and U15820 (N_15820,N_15491,N_15495);
or U15821 (N_15821,N_15434,N_15447);
nor U15822 (N_15822,N_15530,N_15541);
or U15823 (N_15823,N_15546,N_15315);
and U15824 (N_15824,N_15389,N_15506);
and U15825 (N_15825,N_15412,N_15532);
or U15826 (N_15826,N_15360,N_15557);
nor U15827 (N_15827,N_15356,N_15344);
nor U15828 (N_15828,N_15322,N_15476);
xor U15829 (N_15829,N_15445,N_15576);
nand U15830 (N_15830,N_15530,N_15599);
or U15831 (N_15831,N_15511,N_15549);
and U15832 (N_15832,N_15432,N_15533);
and U15833 (N_15833,N_15355,N_15526);
and U15834 (N_15834,N_15416,N_15402);
or U15835 (N_15835,N_15452,N_15456);
and U15836 (N_15836,N_15564,N_15306);
and U15837 (N_15837,N_15556,N_15406);
or U15838 (N_15838,N_15453,N_15310);
nand U15839 (N_15839,N_15353,N_15536);
nor U15840 (N_15840,N_15502,N_15482);
and U15841 (N_15841,N_15337,N_15357);
and U15842 (N_15842,N_15534,N_15586);
or U15843 (N_15843,N_15578,N_15583);
nor U15844 (N_15844,N_15580,N_15549);
or U15845 (N_15845,N_15582,N_15550);
nor U15846 (N_15846,N_15310,N_15334);
and U15847 (N_15847,N_15329,N_15539);
and U15848 (N_15848,N_15490,N_15316);
or U15849 (N_15849,N_15525,N_15576);
nand U15850 (N_15850,N_15420,N_15361);
nor U15851 (N_15851,N_15578,N_15334);
nor U15852 (N_15852,N_15310,N_15405);
xnor U15853 (N_15853,N_15525,N_15436);
and U15854 (N_15854,N_15378,N_15314);
nor U15855 (N_15855,N_15411,N_15392);
or U15856 (N_15856,N_15436,N_15460);
or U15857 (N_15857,N_15398,N_15498);
and U15858 (N_15858,N_15522,N_15423);
nand U15859 (N_15859,N_15596,N_15336);
xor U15860 (N_15860,N_15589,N_15495);
nand U15861 (N_15861,N_15542,N_15448);
and U15862 (N_15862,N_15544,N_15582);
and U15863 (N_15863,N_15483,N_15561);
nor U15864 (N_15864,N_15490,N_15391);
nand U15865 (N_15865,N_15546,N_15469);
xnor U15866 (N_15866,N_15493,N_15597);
and U15867 (N_15867,N_15438,N_15407);
or U15868 (N_15868,N_15508,N_15526);
nor U15869 (N_15869,N_15387,N_15515);
nand U15870 (N_15870,N_15542,N_15534);
nand U15871 (N_15871,N_15328,N_15591);
nand U15872 (N_15872,N_15323,N_15348);
or U15873 (N_15873,N_15310,N_15516);
xnor U15874 (N_15874,N_15317,N_15596);
and U15875 (N_15875,N_15446,N_15573);
or U15876 (N_15876,N_15599,N_15510);
or U15877 (N_15877,N_15403,N_15493);
or U15878 (N_15878,N_15578,N_15441);
nand U15879 (N_15879,N_15314,N_15483);
xnor U15880 (N_15880,N_15425,N_15346);
xnor U15881 (N_15881,N_15599,N_15433);
xor U15882 (N_15882,N_15471,N_15495);
nand U15883 (N_15883,N_15590,N_15536);
or U15884 (N_15884,N_15357,N_15411);
nand U15885 (N_15885,N_15463,N_15550);
and U15886 (N_15886,N_15342,N_15576);
xnor U15887 (N_15887,N_15415,N_15484);
nand U15888 (N_15888,N_15373,N_15494);
or U15889 (N_15889,N_15306,N_15560);
and U15890 (N_15890,N_15529,N_15331);
and U15891 (N_15891,N_15576,N_15509);
nand U15892 (N_15892,N_15535,N_15380);
nand U15893 (N_15893,N_15365,N_15529);
and U15894 (N_15894,N_15313,N_15469);
nand U15895 (N_15895,N_15400,N_15480);
xor U15896 (N_15896,N_15573,N_15428);
nor U15897 (N_15897,N_15385,N_15538);
nand U15898 (N_15898,N_15314,N_15388);
nand U15899 (N_15899,N_15528,N_15356);
or U15900 (N_15900,N_15683,N_15728);
or U15901 (N_15901,N_15676,N_15871);
or U15902 (N_15902,N_15874,N_15673);
xnor U15903 (N_15903,N_15843,N_15801);
nand U15904 (N_15904,N_15609,N_15691);
nand U15905 (N_15905,N_15678,N_15734);
nand U15906 (N_15906,N_15739,N_15600);
or U15907 (N_15907,N_15857,N_15898);
and U15908 (N_15908,N_15767,N_15668);
nor U15909 (N_15909,N_15613,N_15817);
nand U15910 (N_15910,N_15657,N_15677);
nor U15911 (N_15911,N_15698,N_15794);
and U15912 (N_15912,N_15674,N_15730);
nand U15913 (N_15913,N_15792,N_15731);
nand U15914 (N_15914,N_15760,N_15768);
nand U15915 (N_15915,N_15895,N_15861);
nor U15916 (N_15916,N_15814,N_15772);
nor U15917 (N_15917,N_15686,N_15833);
nand U15918 (N_15918,N_15836,N_15816);
nor U15919 (N_15919,N_15650,N_15709);
nor U15920 (N_15920,N_15696,N_15882);
xor U15921 (N_15921,N_15884,N_15702);
xor U15922 (N_15922,N_15758,N_15839);
and U15923 (N_15923,N_15626,N_15873);
nand U15924 (N_15924,N_15813,N_15659);
and U15925 (N_15925,N_15829,N_15822);
or U15926 (N_15926,N_15893,N_15685);
or U15927 (N_15927,N_15705,N_15740);
nor U15928 (N_15928,N_15791,N_15615);
nand U15929 (N_15929,N_15879,N_15812);
or U15930 (N_15930,N_15846,N_15638);
and U15931 (N_15931,N_15679,N_15856);
and U15932 (N_15932,N_15820,N_15680);
or U15933 (N_15933,N_15756,N_15749);
and U15934 (N_15934,N_15798,N_15867);
and U15935 (N_15935,N_15865,N_15703);
nor U15936 (N_15936,N_15722,N_15644);
xor U15937 (N_15937,N_15635,N_15704);
xnor U15938 (N_15938,N_15684,N_15888);
xnor U15939 (N_15939,N_15751,N_15866);
nor U15940 (N_15940,N_15853,N_15773);
nand U15941 (N_15941,N_15629,N_15776);
nor U15942 (N_15942,N_15640,N_15639);
nor U15943 (N_15943,N_15819,N_15782);
and U15944 (N_15944,N_15706,N_15786);
or U15945 (N_15945,N_15724,N_15634);
nand U15946 (N_15946,N_15618,N_15779);
or U15947 (N_15947,N_15682,N_15752);
or U15948 (N_15948,N_15723,N_15654);
and U15949 (N_15949,N_15642,N_15842);
nor U15950 (N_15950,N_15669,N_15780);
nand U15951 (N_15951,N_15652,N_15745);
nor U15952 (N_15952,N_15851,N_15736);
nor U15953 (N_15953,N_15793,N_15738);
or U15954 (N_15954,N_15818,N_15777);
nand U15955 (N_15955,N_15850,N_15651);
and U15956 (N_15956,N_15789,N_15810);
and U15957 (N_15957,N_15837,N_15627);
or U15958 (N_15958,N_15800,N_15687);
and U15959 (N_15959,N_15887,N_15648);
xnor U15960 (N_15960,N_15719,N_15649);
and U15961 (N_15961,N_15708,N_15746);
nor U15962 (N_15962,N_15774,N_15855);
or U15963 (N_15963,N_15766,N_15610);
xor U15964 (N_15964,N_15718,N_15670);
and U15965 (N_15965,N_15628,N_15690);
or U15966 (N_15966,N_15616,N_15747);
or U15967 (N_15967,N_15844,N_15623);
or U15968 (N_15968,N_15605,N_15869);
nor U15969 (N_15969,N_15636,N_15604);
xnor U15970 (N_15970,N_15894,N_15735);
xnor U15971 (N_15971,N_15707,N_15602);
or U15972 (N_15972,N_15781,N_15611);
and U15973 (N_15973,N_15715,N_15761);
and U15974 (N_15974,N_15872,N_15714);
nand U15975 (N_15975,N_15647,N_15890);
xnor U15976 (N_15976,N_15664,N_15787);
xor U15977 (N_15977,N_15631,N_15625);
nand U15978 (N_15978,N_15838,N_15721);
xor U15979 (N_15979,N_15716,N_15880);
nand U15980 (N_15980,N_15797,N_15886);
and U15981 (N_15981,N_15830,N_15725);
xor U15982 (N_15982,N_15614,N_15630);
xor U15983 (N_15983,N_15675,N_15808);
nand U15984 (N_15984,N_15825,N_15859);
xnor U15985 (N_15985,N_15753,N_15729);
or U15986 (N_15986,N_15784,N_15883);
and U15987 (N_15987,N_15633,N_15821);
or U15988 (N_15988,N_15854,N_15658);
and U15989 (N_15989,N_15617,N_15665);
xnor U15990 (N_15990,N_15732,N_15827);
nor U15991 (N_15991,N_15622,N_15763);
or U15992 (N_15992,N_15845,N_15770);
or U15993 (N_15993,N_15858,N_15620);
and U15994 (N_15994,N_15663,N_15655);
and U15995 (N_15995,N_15726,N_15619);
nand U15996 (N_15996,N_15868,N_15878);
nor U15997 (N_15997,N_15860,N_15656);
xnor U15998 (N_15998,N_15662,N_15764);
and U15999 (N_15999,N_15834,N_15637);
nor U16000 (N_16000,N_15612,N_15896);
nor U16001 (N_16001,N_15828,N_15840);
nor U16002 (N_16002,N_15835,N_15757);
nand U16003 (N_16003,N_15742,N_15778);
or U16004 (N_16004,N_15826,N_15823);
nor U16005 (N_16005,N_15653,N_15688);
xnor U16006 (N_16006,N_15755,N_15892);
nand U16007 (N_16007,N_15645,N_15885);
nand U16008 (N_16008,N_15807,N_15671);
or U16009 (N_16009,N_15775,N_15712);
or U16010 (N_16010,N_15802,N_15841);
or U16011 (N_16011,N_15891,N_15720);
nand U16012 (N_16012,N_15831,N_15788);
nand U16013 (N_16013,N_15899,N_15711);
nor U16014 (N_16014,N_15805,N_15632);
nor U16015 (N_16015,N_15815,N_15697);
nor U16016 (N_16016,N_15769,N_15641);
and U16017 (N_16017,N_15783,N_15660);
nor U16018 (N_16018,N_15881,N_15759);
nand U16019 (N_16019,N_15710,N_15608);
nor U16020 (N_16020,N_15824,N_15795);
and U16021 (N_16021,N_15701,N_15876);
and U16022 (N_16022,N_15607,N_15750);
and U16023 (N_16023,N_15681,N_15877);
and U16024 (N_16024,N_15646,N_15771);
or U16025 (N_16025,N_15695,N_15727);
and U16026 (N_16026,N_15743,N_15744);
or U16027 (N_16027,N_15848,N_15692);
nor U16028 (N_16028,N_15693,N_15803);
or U16029 (N_16029,N_15852,N_15667);
or U16030 (N_16030,N_15741,N_15785);
xor U16031 (N_16031,N_15862,N_15806);
nor U16032 (N_16032,N_15811,N_15694);
or U16033 (N_16033,N_15700,N_15870);
xor U16034 (N_16034,N_15889,N_15733);
nand U16035 (N_16035,N_15621,N_15643);
nand U16036 (N_16036,N_15606,N_15603);
nor U16037 (N_16037,N_15737,N_15601);
nor U16038 (N_16038,N_15748,N_15804);
nand U16039 (N_16039,N_15809,N_15847);
nand U16040 (N_16040,N_15799,N_15713);
or U16041 (N_16041,N_15699,N_15863);
and U16042 (N_16042,N_15717,N_15666);
nand U16043 (N_16043,N_15765,N_15672);
xnor U16044 (N_16044,N_15762,N_15849);
xor U16045 (N_16045,N_15790,N_15689);
or U16046 (N_16046,N_15832,N_15754);
nand U16047 (N_16047,N_15796,N_15661);
nand U16048 (N_16048,N_15624,N_15875);
nor U16049 (N_16049,N_15864,N_15897);
nand U16050 (N_16050,N_15750,N_15884);
and U16051 (N_16051,N_15616,N_15600);
or U16052 (N_16052,N_15674,N_15812);
or U16053 (N_16053,N_15867,N_15839);
or U16054 (N_16054,N_15670,N_15665);
or U16055 (N_16055,N_15669,N_15759);
and U16056 (N_16056,N_15729,N_15831);
nor U16057 (N_16057,N_15884,N_15793);
nor U16058 (N_16058,N_15703,N_15807);
and U16059 (N_16059,N_15668,N_15631);
and U16060 (N_16060,N_15750,N_15746);
nor U16061 (N_16061,N_15686,N_15719);
nor U16062 (N_16062,N_15661,N_15634);
nand U16063 (N_16063,N_15648,N_15743);
or U16064 (N_16064,N_15726,N_15709);
nand U16065 (N_16065,N_15830,N_15896);
nand U16066 (N_16066,N_15837,N_15656);
xnor U16067 (N_16067,N_15897,N_15835);
xnor U16068 (N_16068,N_15714,N_15602);
nand U16069 (N_16069,N_15728,N_15609);
and U16070 (N_16070,N_15680,N_15756);
and U16071 (N_16071,N_15636,N_15698);
or U16072 (N_16072,N_15848,N_15754);
nor U16073 (N_16073,N_15835,N_15772);
or U16074 (N_16074,N_15686,N_15794);
nand U16075 (N_16075,N_15700,N_15640);
nor U16076 (N_16076,N_15671,N_15754);
nor U16077 (N_16077,N_15636,N_15659);
nor U16078 (N_16078,N_15705,N_15881);
nor U16079 (N_16079,N_15852,N_15750);
xnor U16080 (N_16080,N_15898,N_15689);
or U16081 (N_16081,N_15899,N_15710);
nor U16082 (N_16082,N_15850,N_15876);
or U16083 (N_16083,N_15635,N_15816);
or U16084 (N_16084,N_15765,N_15893);
or U16085 (N_16085,N_15665,N_15676);
nand U16086 (N_16086,N_15756,N_15802);
and U16087 (N_16087,N_15601,N_15649);
xnor U16088 (N_16088,N_15719,N_15735);
or U16089 (N_16089,N_15728,N_15778);
and U16090 (N_16090,N_15786,N_15721);
xnor U16091 (N_16091,N_15769,N_15755);
xnor U16092 (N_16092,N_15605,N_15767);
nor U16093 (N_16093,N_15816,N_15770);
and U16094 (N_16094,N_15734,N_15628);
nand U16095 (N_16095,N_15605,N_15799);
nand U16096 (N_16096,N_15787,N_15860);
nand U16097 (N_16097,N_15672,N_15737);
xor U16098 (N_16098,N_15868,N_15708);
xor U16099 (N_16099,N_15746,N_15688);
nand U16100 (N_16100,N_15676,N_15664);
xnor U16101 (N_16101,N_15615,N_15716);
nor U16102 (N_16102,N_15661,N_15650);
and U16103 (N_16103,N_15766,N_15832);
nand U16104 (N_16104,N_15874,N_15873);
and U16105 (N_16105,N_15781,N_15664);
or U16106 (N_16106,N_15613,N_15642);
nor U16107 (N_16107,N_15871,N_15782);
nor U16108 (N_16108,N_15617,N_15835);
nand U16109 (N_16109,N_15855,N_15614);
nand U16110 (N_16110,N_15646,N_15809);
or U16111 (N_16111,N_15690,N_15668);
nand U16112 (N_16112,N_15629,N_15813);
nor U16113 (N_16113,N_15702,N_15603);
and U16114 (N_16114,N_15685,N_15622);
nor U16115 (N_16115,N_15766,N_15746);
or U16116 (N_16116,N_15645,N_15652);
nor U16117 (N_16117,N_15788,N_15812);
and U16118 (N_16118,N_15842,N_15841);
nand U16119 (N_16119,N_15836,N_15802);
nand U16120 (N_16120,N_15816,N_15808);
nor U16121 (N_16121,N_15733,N_15806);
xor U16122 (N_16122,N_15723,N_15871);
nand U16123 (N_16123,N_15665,N_15737);
and U16124 (N_16124,N_15836,N_15745);
nand U16125 (N_16125,N_15863,N_15757);
and U16126 (N_16126,N_15708,N_15870);
nor U16127 (N_16127,N_15746,N_15894);
and U16128 (N_16128,N_15694,N_15852);
xnor U16129 (N_16129,N_15828,N_15792);
nor U16130 (N_16130,N_15883,N_15793);
nand U16131 (N_16131,N_15717,N_15766);
nand U16132 (N_16132,N_15661,N_15898);
xnor U16133 (N_16133,N_15731,N_15773);
or U16134 (N_16134,N_15894,N_15621);
xor U16135 (N_16135,N_15705,N_15843);
and U16136 (N_16136,N_15764,N_15872);
nand U16137 (N_16137,N_15710,N_15637);
nor U16138 (N_16138,N_15719,N_15842);
nor U16139 (N_16139,N_15798,N_15645);
nand U16140 (N_16140,N_15644,N_15810);
and U16141 (N_16141,N_15674,N_15733);
nand U16142 (N_16142,N_15881,N_15792);
xor U16143 (N_16143,N_15767,N_15875);
or U16144 (N_16144,N_15808,N_15831);
xor U16145 (N_16145,N_15789,N_15725);
nor U16146 (N_16146,N_15684,N_15606);
xnor U16147 (N_16147,N_15689,N_15713);
and U16148 (N_16148,N_15856,N_15697);
and U16149 (N_16149,N_15756,N_15729);
or U16150 (N_16150,N_15774,N_15729);
or U16151 (N_16151,N_15864,N_15814);
and U16152 (N_16152,N_15747,N_15824);
nor U16153 (N_16153,N_15762,N_15789);
xor U16154 (N_16154,N_15704,N_15641);
nor U16155 (N_16155,N_15739,N_15840);
and U16156 (N_16156,N_15748,N_15832);
nor U16157 (N_16157,N_15658,N_15613);
nand U16158 (N_16158,N_15781,N_15677);
nand U16159 (N_16159,N_15707,N_15865);
nand U16160 (N_16160,N_15713,N_15607);
nand U16161 (N_16161,N_15773,N_15651);
xnor U16162 (N_16162,N_15749,N_15824);
nand U16163 (N_16163,N_15654,N_15819);
nand U16164 (N_16164,N_15779,N_15704);
xnor U16165 (N_16165,N_15625,N_15607);
xnor U16166 (N_16166,N_15653,N_15610);
or U16167 (N_16167,N_15847,N_15762);
or U16168 (N_16168,N_15700,N_15860);
and U16169 (N_16169,N_15897,N_15838);
nand U16170 (N_16170,N_15746,N_15805);
nor U16171 (N_16171,N_15819,N_15638);
xor U16172 (N_16172,N_15803,N_15887);
and U16173 (N_16173,N_15896,N_15680);
and U16174 (N_16174,N_15684,N_15726);
xnor U16175 (N_16175,N_15750,N_15757);
nand U16176 (N_16176,N_15823,N_15742);
nor U16177 (N_16177,N_15696,N_15828);
nand U16178 (N_16178,N_15871,N_15881);
or U16179 (N_16179,N_15658,N_15791);
and U16180 (N_16180,N_15798,N_15776);
xnor U16181 (N_16181,N_15870,N_15885);
xor U16182 (N_16182,N_15738,N_15884);
and U16183 (N_16183,N_15669,N_15673);
xnor U16184 (N_16184,N_15701,N_15633);
xnor U16185 (N_16185,N_15658,N_15674);
nor U16186 (N_16186,N_15765,N_15701);
nand U16187 (N_16187,N_15873,N_15601);
or U16188 (N_16188,N_15729,N_15653);
or U16189 (N_16189,N_15645,N_15657);
nand U16190 (N_16190,N_15867,N_15893);
xor U16191 (N_16191,N_15698,N_15762);
and U16192 (N_16192,N_15838,N_15697);
nand U16193 (N_16193,N_15769,N_15791);
nand U16194 (N_16194,N_15633,N_15663);
xnor U16195 (N_16195,N_15679,N_15835);
nand U16196 (N_16196,N_15843,N_15759);
nor U16197 (N_16197,N_15867,N_15788);
nor U16198 (N_16198,N_15602,N_15734);
nor U16199 (N_16199,N_15829,N_15617);
nor U16200 (N_16200,N_16087,N_16188);
or U16201 (N_16201,N_16195,N_15926);
nand U16202 (N_16202,N_16059,N_16128);
xor U16203 (N_16203,N_16036,N_15948);
and U16204 (N_16204,N_16082,N_16072);
nand U16205 (N_16205,N_16190,N_16143);
and U16206 (N_16206,N_16056,N_15979);
nand U16207 (N_16207,N_16000,N_16020);
or U16208 (N_16208,N_15917,N_16158);
and U16209 (N_16209,N_16193,N_16064);
or U16210 (N_16210,N_16052,N_15970);
xnor U16211 (N_16211,N_16006,N_15906);
nand U16212 (N_16212,N_15955,N_16119);
nor U16213 (N_16213,N_15943,N_16029);
xnor U16214 (N_16214,N_16102,N_16108);
xnor U16215 (N_16215,N_15976,N_15984);
nor U16216 (N_16216,N_15945,N_16018);
and U16217 (N_16217,N_15944,N_15916);
and U16218 (N_16218,N_16152,N_16041);
xor U16219 (N_16219,N_15909,N_16010);
or U16220 (N_16220,N_16167,N_16185);
or U16221 (N_16221,N_15957,N_16155);
and U16222 (N_16222,N_15932,N_16177);
nor U16223 (N_16223,N_15923,N_15967);
nor U16224 (N_16224,N_15949,N_16025);
xor U16225 (N_16225,N_15975,N_16042);
nand U16226 (N_16226,N_16031,N_16109);
or U16227 (N_16227,N_15969,N_15966);
and U16228 (N_16228,N_15954,N_15958);
and U16229 (N_16229,N_16071,N_16138);
or U16230 (N_16230,N_15902,N_15935);
nand U16231 (N_16231,N_15900,N_16089);
or U16232 (N_16232,N_15939,N_16165);
xnor U16233 (N_16233,N_16101,N_16121);
nor U16234 (N_16234,N_16054,N_16049);
xnor U16235 (N_16235,N_16024,N_16032);
or U16236 (N_16236,N_15997,N_15946);
and U16237 (N_16237,N_16053,N_16160);
and U16238 (N_16238,N_16170,N_16171);
xor U16239 (N_16239,N_15993,N_16065);
nor U16240 (N_16240,N_16081,N_15907);
nor U16241 (N_16241,N_16113,N_16034);
nand U16242 (N_16242,N_15901,N_16043);
or U16243 (N_16243,N_15910,N_15994);
xnor U16244 (N_16244,N_16086,N_16107);
nand U16245 (N_16245,N_16001,N_16186);
nor U16246 (N_16246,N_15942,N_15947);
or U16247 (N_16247,N_16146,N_15922);
or U16248 (N_16248,N_16033,N_15929);
nor U16249 (N_16249,N_16077,N_16110);
and U16250 (N_16250,N_16123,N_16048);
xor U16251 (N_16251,N_16004,N_16106);
nor U16252 (N_16252,N_16046,N_15905);
nor U16253 (N_16253,N_16194,N_16061);
nand U16254 (N_16254,N_16088,N_16080);
nand U16255 (N_16255,N_15987,N_15940);
or U16256 (N_16256,N_16150,N_16192);
xor U16257 (N_16257,N_16181,N_16125);
nor U16258 (N_16258,N_16124,N_16168);
xor U16259 (N_16259,N_16091,N_16189);
nand U16260 (N_16260,N_16069,N_16131);
xor U16261 (N_16261,N_16013,N_16094);
nand U16262 (N_16262,N_16093,N_15952);
and U16263 (N_16263,N_16074,N_16015);
nor U16264 (N_16264,N_16176,N_15982);
nand U16265 (N_16265,N_15915,N_16178);
nor U16266 (N_16266,N_16162,N_16067);
or U16267 (N_16267,N_16005,N_16161);
and U16268 (N_16268,N_15903,N_16130);
nor U16269 (N_16269,N_15988,N_16122);
xnor U16270 (N_16270,N_15904,N_16112);
nor U16271 (N_16271,N_16085,N_15931);
or U16272 (N_16272,N_15963,N_16133);
nor U16273 (N_16273,N_16154,N_16066);
nand U16274 (N_16274,N_15983,N_16145);
xnor U16275 (N_16275,N_16100,N_16179);
nand U16276 (N_16276,N_16076,N_16023);
nand U16277 (N_16277,N_15934,N_16047);
xnor U16278 (N_16278,N_16092,N_16103);
or U16279 (N_16279,N_16037,N_16180);
nand U16280 (N_16280,N_16009,N_16026);
nand U16281 (N_16281,N_16051,N_16058);
xnor U16282 (N_16282,N_16135,N_15930);
nor U16283 (N_16283,N_15919,N_16014);
nor U16284 (N_16284,N_16172,N_16079);
nor U16285 (N_16285,N_16017,N_15924);
and U16286 (N_16286,N_15990,N_16073);
nor U16287 (N_16287,N_15991,N_16097);
and U16288 (N_16288,N_16039,N_16127);
or U16289 (N_16289,N_16012,N_15965);
or U16290 (N_16290,N_15920,N_16175);
xnor U16291 (N_16291,N_16044,N_16104);
or U16292 (N_16292,N_16030,N_16111);
xor U16293 (N_16293,N_15999,N_16011);
and U16294 (N_16294,N_16027,N_16045);
xnor U16295 (N_16295,N_16070,N_16096);
and U16296 (N_16296,N_16166,N_16182);
or U16297 (N_16297,N_15953,N_15996);
nor U16298 (N_16298,N_16114,N_16126);
and U16299 (N_16299,N_16144,N_15960);
and U16300 (N_16300,N_16149,N_16173);
nor U16301 (N_16301,N_16038,N_15992);
or U16302 (N_16302,N_15913,N_16084);
and U16303 (N_16303,N_16140,N_15956);
xnor U16304 (N_16304,N_16118,N_16156);
and U16305 (N_16305,N_15998,N_16083);
and U16306 (N_16306,N_15980,N_16147);
nand U16307 (N_16307,N_15918,N_15914);
nor U16308 (N_16308,N_15962,N_16022);
or U16309 (N_16309,N_16078,N_16068);
nor U16310 (N_16310,N_16134,N_16187);
nor U16311 (N_16311,N_16019,N_16184);
or U16312 (N_16312,N_15911,N_16002);
nor U16313 (N_16313,N_16063,N_15964);
nand U16314 (N_16314,N_15925,N_15927);
nor U16315 (N_16315,N_16115,N_16008);
nor U16316 (N_16316,N_15908,N_16136);
nand U16317 (N_16317,N_15973,N_16164);
nand U16318 (N_16318,N_15968,N_15950);
xor U16319 (N_16319,N_16095,N_16117);
xnor U16320 (N_16320,N_15936,N_15989);
nor U16321 (N_16321,N_16196,N_16120);
or U16322 (N_16322,N_15938,N_16151);
and U16323 (N_16323,N_16159,N_15971);
xnor U16324 (N_16324,N_16132,N_16141);
nand U16325 (N_16325,N_15972,N_15937);
or U16326 (N_16326,N_16060,N_15986);
nand U16327 (N_16327,N_16003,N_15977);
xor U16328 (N_16328,N_16148,N_15912);
or U16329 (N_16329,N_16090,N_16028);
and U16330 (N_16330,N_15985,N_15981);
nor U16331 (N_16331,N_16040,N_16191);
nand U16332 (N_16332,N_16129,N_16142);
xor U16333 (N_16333,N_16197,N_16198);
and U16334 (N_16334,N_16099,N_16007);
nand U16335 (N_16335,N_16035,N_16098);
and U16336 (N_16336,N_16075,N_16139);
or U16337 (N_16337,N_16174,N_15933);
or U16338 (N_16338,N_16116,N_16153);
xor U16339 (N_16339,N_16055,N_15951);
and U16340 (N_16340,N_16050,N_15995);
xor U16341 (N_16341,N_16157,N_16105);
nor U16342 (N_16342,N_16169,N_16199);
or U16343 (N_16343,N_16016,N_15961);
nor U16344 (N_16344,N_16163,N_15941);
xor U16345 (N_16345,N_16062,N_15928);
nor U16346 (N_16346,N_16057,N_15974);
or U16347 (N_16347,N_15978,N_15921);
nor U16348 (N_16348,N_16183,N_15959);
nand U16349 (N_16349,N_16021,N_16137);
nor U16350 (N_16350,N_16099,N_15959);
nor U16351 (N_16351,N_15916,N_15976);
nor U16352 (N_16352,N_15952,N_16110);
or U16353 (N_16353,N_16136,N_16121);
nand U16354 (N_16354,N_15974,N_16105);
nor U16355 (N_16355,N_15994,N_16071);
and U16356 (N_16356,N_16073,N_16055);
xor U16357 (N_16357,N_15936,N_16087);
nor U16358 (N_16358,N_15917,N_15960);
xor U16359 (N_16359,N_16115,N_16013);
and U16360 (N_16360,N_16177,N_16012);
nand U16361 (N_16361,N_16177,N_15917);
nor U16362 (N_16362,N_16126,N_15980);
nand U16363 (N_16363,N_16142,N_16119);
nand U16364 (N_16364,N_16146,N_15909);
xor U16365 (N_16365,N_16089,N_16106);
nor U16366 (N_16366,N_16154,N_15990);
or U16367 (N_16367,N_16167,N_15916);
and U16368 (N_16368,N_16127,N_16012);
or U16369 (N_16369,N_15945,N_16006);
and U16370 (N_16370,N_16143,N_15941);
nand U16371 (N_16371,N_15993,N_16133);
nand U16372 (N_16372,N_16052,N_16016);
nand U16373 (N_16373,N_15937,N_15925);
or U16374 (N_16374,N_15995,N_16002);
nand U16375 (N_16375,N_16136,N_16169);
nor U16376 (N_16376,N_16066,N_15903);
nor U16377 (N_16377,N_15916,N_16081);
xnor U16378 (N_16378,N_15973,N_16121);
nor U16379 (N_16379,N_16089,N_15998);
and U16380 (N_16380,N_15916,N_15973);
and U16381 (N_16381,N_16013,N_16075);
xnor U16382 (N_16382,N_16164,N_15933);
nor U16383 (N_16383,N_16118,N_16187);
nor U16384 (N_16384,N_16094,N_15992);
nand U16385 (N_16385,N_16181,N_15904);
xnor U16386 (N_16386,N_16082,N_15983);
nand U16387 (N_16387,N_15977,N_15997);
and U16388 (N_16388,N_15907,N_16099);
xor U16389 (N_16389,N_15915,N_16164);
or U16390 (N_16390,N_16191,N_15970);
or U16391 (N_16391,N_15923,N_16018);
xnor U16392 (N_16392,N_15971,N_15949);
and U16393 (N_16393,N_15927,N_16083);
nand U16394 (N_16394,N_15960,N_15950);
xnor U16395 (N_16395,N_15974,N_16038);
and U16396 (N_16396,N_16115,N_15994);
nor U16397 (N_16397,N_16042,N_16084);
nor U16398 (N_16398,N_15972,N_16014);
nor U16399 (N_16399,N_16010,N_15997);
nand U16400 (N_16400,N_16073,N_16138);
nand U16401 (N_16401,N_15940,N_16157);
nand U16402 (N_16402,N_15993,N_15967);
xnor U16403 (N_16403,N_15942,N_16198);
or U16404 (N_16404,N_15904,N_15920);
nand U16405 (N_16405,N_16128,N_16145);
xor U16406 (N_16406,N_16115,N_16030);
and U16407 (N_16407,N_15997,N_16007);
xnor U16408 (N_16408,N_16186,N_16016);
and U16409 (N_16409,N_15924,N_16143);
nand U16410 (N_16410,N_16167,N_16005);
nand U16411 (N_16411,N_16011,N_16143);
or U16412 (N_16412,N_16063,N_16054);
xnor U16413 (N_16413,N_16171,N_16025);
nor U16414 (N_16414,N_16088,N_15990);
and U16415 (N_16415,N_16148,N_15918);
or U16416 (N_16416,N_15976,N_15985);
nand U16417 (N_16417,N_15940,N_16158);
or U16418 (N_16418,N_15996,N_16091);
nor U16419 (N_16419,N_15940,N_16123);
nand U16420 (N_16420,N_16072,N_15992);
nor U16421 (N_16421,N_16052,N_16195);
nand U16422 (N_16422,N_16025,N_15921);
and U16423 (N_16423,N_16117,N_15918);
nor U16424 (N_16424,N_15958,N_16046);
nor U16425 (N_16425,N_16199,N_16175);
and U16426 (N_16426,N_16097,N_16052);
and U16427 (N_16427,N_16139,N_15911);
or U16428 (N_16428,N_15906,N_15996);
nor U16429 (N_16429,N_16197,N_16145);
xnor U16430 (N_16430,N_15984,N_16051);
xor U16431 (N_16431,N_15995,N_15901);
or U16432 (N_16432,N_16131,N_16163);
nand U16433 (N_16433,N_16020,N_15945);
nand U16434 (N_16434,N_16121,N_15907);
nor U16435 (N_16435,N_16132,N_16035);
nand U16436 (N_16436,N_16067,N_16091);
xor U16437 (N_16437,N_16192,N_15985);
nor U16438 (N_16438,N_16081,N_16163);
and U16439 (N_16439,N_16089,N_16080);
and U16440 (N_16440,N_16081,N_16074);
nand U16441 (N_16441,N_16124,N_16181);
nor U16442 (N_16442,N_16102,N_15909);
nand U16443 (N_16443,N_16131,N_16070);
or U16444 (N_16444,N_16126,N_16089);
nor U16445 (N_16445,N_16166,N_15928);
and U16446 (N_16446,N_16122,N_16038);
nor U16447 (N_16447,N_16187,N_15943);
and U16448 (N_16448,N_16061,N_15984);
xnor U16449 (N_16449,N_15962,N_16004);
nand U16450 (N_16450,N_15945,N_15966);
or U16451 (N_16451,N_16193,N_16058);
and U16452 (N_16452,N_16117,N_16115);
nor U16453 (N_16453,N_16139,N_16098);
nor U16454 (N_16454,N_15979,N_15943);
nand U16455 (N_16455,N_16065,N_15951);
nor U16456 (N_16456,N_16127,N_16040);
xnor U16457 (N_16457,N_16023,N_16012);
and U16458 (N_16458,N_15994,N_15944);
and U16459 (N_16459,N_15988,N_16030);
and U16460 (N_16460,N_15921,N_16073);
nor U16461 (N_16461,N_15956,N_15986);
or U16462 (N_16462,N_16001,N_16039);
xor U16463 (N_16463,N_15932,N_16164);
and U16464 (N_16464,N_16098,N_16038);
xnor U16465 (N_16465,N_15981,N_15901);
or U16466 (N_16466,N_15918,N_16199);
nor U16467 (N_16467,N_16101,N_15948);
nand U16468 (N_16468,N_15961,N_15989);
and U16469 (N_16469,N_15935,N_15989);
nor U16470 (N_16470,N_16102,N_16183);
nor U16471 (N_16471,N_16068,N_16080);
and U16472 (N_16472,N_16017,N_15921);
nand U16473 (N_16473,N_15900,N_15950);
or U16474 (N_16474,N_15919,N_16034);
or U16475 (N_16475,N_16016,N_15924);
nand U16476 (N_16476,N_16041,N_16052);
xor U16477 (N_16477,N_15930,N_15938);
xor U16478 (N_16478,N_15908,N_16160);
or U16479 (N_16479,N_16114,N_16040);
nand U16480 (N_16480,N_16161,N_16186);
xnor U16481 (N_16481,N_16199,N_15920);
nand U16482 (N_16482,N_16136,N_16026);
and U16483 (N_16483,N_15999,N_16050);
nand U16484 (N_16484,N_15906,N_15930);
nand U16485 (N_16485,N_15904,N_15944);
and U16486 (N_16486,N_15966,N_16114);
nor U16487 (N_16487,N_16065,N_15975);
or U16488 (N_16488,N_15929,N_16198);
and U16489 (N_16489,N_15912,N_16143);
xor U16490 (N_16490,N_15933,N_16047);
nand U16491 (N_16491,N_16107,N_16134);
or U16492 (N_16492,N_16077,N_15951);
and U16493 (N_16493,N_15926,N_15982);
nand U16494 (N_16494,N_15956,N_15984);
xnor U16495 (N_16495,N_16132,N_16106);
and U16496 (N_16496,N_16109,N_16186);
nor U16497 (N_16497,N_16196,N_16082);
nor U16498 (N_16498,N_16131,N_16012);
or U16499 (N_16499,N_16062,N_16044);
or U16500 (N_16500,N_16279,N_16448);
xor U16501 (N_16501,N_16364,N_16404);
or U16502 (N_16502,N_16320,N_16234);
nor U16503 (N_16503,N_16486,N_16491);
and U16504 (N_16504,N_16362,N_16460);
xor U16505 (N_16505,N_16309,N_16451);
nand U16506 (N_16506,N_16218,N_16205);
nand U16507 (N_16507,N_16222,N_16314);
nor U16508 (N_16508,N_16271,N_16267);
or U16509 (N_16509,N_16417,N_16414);
nor U16510 (N_16510,N_16256,N_16418);
nand U16511 (N_16511,N_16359,N_16265);
nand U16512 (N_16512,N_16254,N_16400);
and U16513 (N_16513,N_16423,N_16432);
nor U16514 (N_16514,N_16365,N_16431);
nand U16515 (N_16515,N_16384,N_16268);
nand U16516 (N_16516,N_16356,N_16280);
nand U16517 (N_16517,N_16285,N_16416);
and U16518 (N_16518,N_16250,N_16210);
xnor U16519 (N_16519,N_16380,N_16485);
nor U16520 (N_16520,N_16338,N_16442);
nor U16521 (N_16521,N_16312,N_16288);
nand U16522 (N_16522,N_16408,N_16284);
nand U16523 (N_16523,N_16372,N_16494);
and U16524 (N_16524,N_16323,N_16229);
and U16525 (N_16525,N_16388,N_16335);
and U16526 (N_16526,N_16469,N_16238);
nand U16527 (N_16527,N_16450,N_16459);
xor U16528 (N_16528,N_16353,N_16211);
xor U16529 (N_16529,N_16350,N_16403);
nand U16530 (N_16530,N_16330,N_16474);
xor U16531 (N_16531,N_16440,N_16214);
nor U16532 (N_16532,N_16344,N_16420);
nor U16533 (N_16533,N_16468,N_16382);
or U16534 (N_16534,N_16467,N_16297);
and U16535 (N_16535,N_16274,N_16370);
xor U16536 (N_16536,N_16429,N_16419);
xor U16537 (N_16537,N_16225,N_16295);
xor U16538 (N_16538,N_16224,N_16375);
and U16539 (N_16539,N_16262,N_16347);
nor U16540 (N_16540,N_16345,N_16426);
nor U16541 (N_16541,N_16243,N_16379);
or U16542 (N_16542,N_16464,N_16277);
nor U16543 (N_16543,N_16435,N_16478);
and U16544 (N_16544,N_16292,N_16251);
and U16545 (N_16545,N_16318,N_16287);
nor U16546 (N_16546,N_16480,N_16298);
nor U16547 (N_16547,N_16305,N_16354);
and U16548 (N_16548,N_16294,N_16260);
nor U16549 (N_16549,N_16477,N_16303);
xor U16550 (N_16550,N_16204,N_16289);
and U16551 (N_16551,N_16456,N_16319);
xor U16552 (N_16552,N_16282,N_16249);
nand U16553 (N_16553,N_16449,N_16393);
or U16554 (N_16554,N_16296,N_16278);
and U16555 (N_16555,N_16357,N_16465);
nor U16556 (N_16556,N_16358,N_16458);
nand U16557 (N_16557,N_16377,N_16482);
and U16558 (N_16558,N_16231,N_16471);
nand U16559 (N_16559,N_16457,N_16293);
nor U16560 (N_16560,N_16493,N_16237);
or U16561 (N_16561,N_16240,N_16261);
nor U16562 (N_16562,N_16488,N_16433);
and U16563 (N_16563,N_16302,N_16304);
and U16564 (N_16564,N_16438,N_16409);
nand U16565 (N_16565,N_16290,N_16259);
nor U16566 (N_16566,N_16349,N_16226);
nand U16567 (N_16567,N_16301,N_16483);
and U16568 (N_16568,N_16361,N_16383);
and U16569 (N_16569,N_16373,N_16228);
nand U16570 (N_16570,N_16444,N_16461);
and U16571 (N_16571,N_16208,N_16241);
nor U16572 (N_16572,N_16484,N_16466);
and U16573 (N_16573,N_16317,N_16326);
xnor U16574 (N_16574,N_16399,N_16266);
and U16575 (N_16575,N_16264,N_16328);
or U16576 (N_16576,N_16217,N_16331);
nor U16577 (N_16577,N_16252,N_16415);
and U16578 (N_16578,N_16443,N_16369);
or U16579 (N_16579,N_16425,N_16385);
nor U16580 (N_16580,N_16235,N_16248);
nor U16581 (N_16581,N_16207,N_16233);
xor U16582 (N_16582,N_16454,N_16463);
nand U16583 (N_16583,N_16495,N_16340);
nand U16584 (N_16584,N_16421,N_16275);
xnor U16585 (N_16585,N_16498,N_16230);
nand U16586 (N_16586,N_16339,N_16315);
nand U16587 (N_16587,N_16487,N_16430);
and U16588 (N_16588,N_16216,N_16360);
or U16589 (N_16589,N_16263,N_16223);
nand U16590 (N_16590,N_16321,N_16475);
and U16591 (N_16591,N_16499,N_16201);
and U16592 (N_16592,N_16300,N_16255);
nand U16593 (N_16593,N_16281,N_16401);
nor U16594 (N_16594,N_16424,N_16452);
or U16595 (N_16595,N_16363,N_16367);
nor U16596 (N_16596,N_16283,N_16479);
nand U16597 (N_16597,N_16439,N_16291);
and U16598 (N_16598,N_16376,N_16473);
nand U16599 (N_16599,N_16286,N_16428);
xnor U16600 (N_16600,N_16413,N_16387);
nand U16601 (N_16601,N_16236,N_16206);
or U16602 (N_16602,N_16272,N_16366);
xnor U16603 (N_16603,N_16446,N_16394);
or U16604 (N_16604,N_16476,N_16389);
xnor U16605 (N_16605,N_16246,N_16397);
nand U16606 (N_16606,N_16253,N_16410);
or U16607 (N_16607,N_16244,N_16405);
nand U16608 (N_16608,N_16242,N_16322);
xor U16609 (N_16609,N_16355,N_16332);
nand U16610 (N_16610,N_16386,N_16402);
and U16611 (N_16611,N_16209,N_16313);
or U16612 (N_16612,N_16239,N_16310);
nor U16613 (N_16613,N_16316,N_16348);
nand U16614 (N_16614,N_16490,N_16219);
nor U16615 (N_16615,N_16269,N_16374);
xnor U16616 (N_16616,N_16422,N_16270);
xnor U16617 (N_16617,N_16220,N_16258);
xnor U16618 (N_16618,N_16245,N_16455);
or U16619 (N_16619,N_16329,N_16343);
or U16620 (N_16620,N_16427,N_16337);
xnor U16621 (N_16621,N_16227,N_16247);
or U16622 (N_16622,N_16342,N_16200);
nor U16623 (N_16623,N_16447,N_16437);
xnor U16624 (N_16624,N_16232,N_16327);
xor U16625 (N_16625,N_16436,N_16398);
nor U16626 (N_16626,N_16407,N_16273);
nand U16627 (N_16627,N_16346,N_16202);
or U16628 (N_16628,N_16368,N_16215);
and U16629 (N_16629,N_16470,N_16390);
nor U16630 (N_16630,N_16352,N_16351);
nand U16631 (N_16631,N_16213,N_16391);
nand U16632 (N_16632,N_16333,N_16299);
and U16633 (N_16633,N_16392,N_16325);
and U16634 (N_16634,N_16306,N_16396);
nand U16635 (N_16635,N_16341,N_16445);
nand U16636 (N_16636,N_16307,N_16378);
xnor U16637 (N_16637,N_16412,N_16336);
xnor U16638 (N_16638,N_16276,N_16212);
and U16639 (N_16639,N_16472,N_16221);
nor U16640 (N_16640,N_16497,N_16441);
nor U16641 (N_16641,N_16334,N_16434);
xnor U16642 (N_16642,N_16492,N_16381);
nand U16643 (N_16643,N_16311,N_16406);
nand U16644 (N_16644,N_16324,N_16257);
nand U16645 (N_16645,N_16411,N_16496);
xor U16646 (N_16646,N_16203,N_16462);
or U16647 (N_16647,N_16481,N_16395);
and U16648 (N_16648,N_16371,N_16453);
xor U16649 (N_16649,N_16308,N_16489);
xor U16650 (N_16650,N_16218,N_16220);
or U16651 (N_16651,N_16214,N_16317);
xor U16652 (N_16652,N_16477,N_16467);
and U16653 (N_16653,N_16261,N_16337);
xnor U16654 (N_16654,N_16339,N_16233);
and U16655 (N_16655,N_16207,N_16296);
nor U16656 (N_16656,N_16335,N_16295);
nor U16657 (N_16657,N_16424,N_16242);
and U16658 (N_16658,N_16455,N_16473);
xor U16659 (N_16659,N_16460,N_16325);
nand U16660 (N_16660,N_16477,N_16485);
xnor U16661 (N_16661,N_16481,N_16381);
and U16662 (N_16662,N_16363,N_16220);
nand U16663 (N_16663,N_16381,N_16288);
xnor U16664 (N_16664,N_16371,N_16490);
xor U16665 (N_16665,N_16435,N_16282);
and U16666 (N_16666,N_16422,N_16314);
or U16667 (N_16667,N_16498,N_16415);
nor U16668 (N_16668,N_16463,N_16455);
xnor U16669 (N_16669,N_16377,N_16280);
xor U16670 (N_16670,N_16462,N_16314);
nand U16671 (N_16671,N_16495,N_16330);
or U16672 (N_16672,N_16296,N_16418);
or U16673 (N_16673,N_16340,N_16281);
and U16674 (N_16674,N_16436,N_16409);
nand U16675 (N_16675,N_16446,N_16276);
nand U16676 (N_16676,N_16360,N_16256);
and U16677 (N_16677,N_16475,N_16417);
and U16678 (N_16678,N_16320,N_16305);
xnor U16679 (N_16679,N_16487,N_16479);
nor U16680 (N_16680,N_16394,N_16271);
nand U16681 (N_16681,N_16207,N_16208);
nor U16682 (N_16682,N_16453,N_16251);
or U16683 (N_16683,N_16246,N_16261);
xnor U16684 (N_16684,N_16489,N_16474);
nor U16685 (N_16685,N_16426,N_16270);
or U16686 (N_16686,N_16264,N_16400);
xnor U16687 (N_16687,N_16322,N_16250);
and U16688 (N_16688,N_16482,N_16342);
nand U16689 (N_16689,N_16494,N_16328);
nand U16690 (N_16690,N_16283,N_16384);
nand U16691 (N_16691,N_16224,N_16275);
nand U16692 (N_16692,N_16418,N_16419);
xnor U16693 (N_16693,N_16433,N_16357);
nand U16694 (N_16694,N_16465,N_16243);
nor U16695 (N_16695,N_16300,N_16386);
nor U16696 (N_16696,N_16271,N_16402);
and U16697 (N_16697,N_16402,N_16420);
or U16698 (N_16698,N_16480,N_16437);
or U16699 (N_16699,N_16345,N_16366);
and U16700 (N_16700,N_16462,N_16442);
and U16701 (N_16701,N_16200,N_16316);
nor U16702 (N_16702,N_16298,N_16291);
or U16703 (N_16703,N_16321,N_16414);
nor U16704 (N_16704,N_16456,N_16264);
and U16705 (N_16705,N_16347,N_16489);
nand U16706 (N_16706,N_16310,N_16480);
or U16707 (N_16707,N_16246,N_16355);
nand U16708 (N_16708,N_16396,N_16219);
nand U16709 (N_16709,N_16266,N_16226);
xor U16710 (N_16710,N_16408,N_16333);
and U16711 (N_16711,N_16264,N_16378);
xnor U16712 (N_16712,N_16466,N_16375);
or U16713 (N_16713,N_16405,N_16318);
xor U16714 (N_16714,N_16250,N_16326);
and U16715 (N_16715,N_16245,N_16299);
nand U16716 (N_16716,N_16271,N_16330);
nand U16717 (N_16717,N_16263,N_16348);
and U16718 (N_16718,N_16340,N_16410);
xnor U16719 (N_16719,N_16235,N_16384);
nand U16720 (N_16720,N_16419,N_16323);
nor U16721 (N_16721,N_16413,N_16369);
nand U16722 (N_16722,N_16322,N_16423);
nand U16723 (N_16723,N_16453,N_16327);
nor U16724 (N_16724,N_16423,N_16375);
nand U16725 (N_16725,N_16204,N_16497);
nand U16726 (N_16726,N_16228,N_16305);
and U16727 (N_16727,N_16379,N_16246);
or U16728 (N_16728,N_16466,N_16225);
nor U16729 (N_16729,N_16396,N_16356);
and U16730 (N_16730,N_16203,N_16439);
and U16731 (N_16731,N_16238,N_16218);
nand U16732 (N_16732,N_16450,N_16442);
nand U16733 (N_16733,N_16278,N_16267);
nor U16734 (N_16734,N_16256,N_16300);
and U16735 (N_16735,N_16375,N_16492);
nor U16736 (N_16736,N_16276,N_16224);
nor U16737 (N_16737,N_16488,N_16286);
and U16738 (N_16738,N_16448,N_16225);
nor U16739 (N_16739,N_16346,N_16488);
and U16740 (N_16740,N_16263,N_16407);
and U16741 (N_16741,N_16285,N_16454);
and U16742 (N_16742,N_16314,N_16495);
nor U16743 (N_16743,N_16225,N_16477);
nand U16744 (N_16744,N_16202,N_16409);
or U16745 (N_16745,N_16290,N_16262);
and U16746 (N_16746,N_16241,N_16430);
or U16747 (N_16747,N_16218,N_16257);
xnor U16748 (N_16748,N_16343,N_16361);
xor U16749 (N_16749,N_16299,N_16273);
and U16750 (N_16750,N_16210,N_16234);
nor U16751 (N_16751,N_16386,N_16248);
or U16752 (N_16752,N_16314,N_16369);
nor U16753 (N_16753,N_16469,N_16333);
or U16754 (N_16754,N_16279,N_16236);
nand U16755 (N_16755,N_16395,N_16273);
nor U16756 (N_16756,N_16464,N_16478);
and U16757 (N_16757,N_16455,N_16449);
xor U16758 (N_16758,N_16252,N_16450);
nand U16759 (N_16759,N_16397,N_16446);
xor U16760 (N_16760,N_16247,N_16455);
nor U16761 (N_16761,N_16467,N_16445);
nor U16762 (N_16762,N_16241,N_16234);
and U16763 (N_16763,N_16309,N_16352);
and U16764 (N_16764,N_16216,N_16468);
nand U16765 (N_16765,N_16231,N_16295);
or U16766 (N_16766,N_16495,N_16341);
xnor U16767 (N_16767,N_16466,N_16232);
nor U16768 (N_16768,N_16416,N_16244);
xor U16769 (N_16769,N_16326,N_16214);
nand U16770 (N_16770,N_16317,N_16279);
xor U16771 (N_16771,N_16309,N_16368);
nor U16772 (N_16772,N_16201,N_16236);
nor U16773 (N_16773,N_16468,N_16423);
or U16774 (N_16774,N_16232,N_16258);
nor U16775 (N_16775,N_16468,N_16433);
nand U16776 (N_16776,N_16343,N_16250);
nor U16777 (N_16777,N_16318,N_16242);
nand U16778 (N_16778,N_16414,N_16388);
nor U16779 (N_16779,N_16230,N_16456);
or U16780 (N_16780,N_16273,N_16202);
nand U16781 (N_16781,N_16374,N_16308);
xnor U16782 (N_16782,N_16270,N_16421);
and U16783 (N_16783,N_16469,N_16404);
nor U16784 (N_16784,N_16271,N_16373);
nand U16785 (N_16785,N_16320,N_16222);
or U16786 (N_16786,N_16495,N_16411);
xnor U16787 (N_16787,N_16359,N_16283);
xor U16788 (N_16788,N_16370,N_16438);
nand U16789 (N_16789,N_16445,N_16499);
nand U16790 (N_16790,N_16298,N_16251);
or U16791 (N_16791,N_16223,N_16244);
nor U16792 (N_16792,N_16491,N_16470);
and U16793 (N_16793,N_16442,N_16484);
and U16794 (N_16794,N_16427,N_16256);
nand U16795 (N_16795,N_16206,N_16357);
nor U16796 (N_16796,N_16303,N_16294);
xor U16797 (N_16797,N_16240,N_16370);
xnor U16798 (N_16798,N_16484,N_16235);
nand U16799 (N_16799,N_16236,N_16273);
or U16800 (N_16800,N_16782,N_16624);
and U16801 (N_16801,N_16709,N_16763);
xnor U16802 (N_16802,N_16730,N_16649);
nand U16803 (N_16803,N_16643,N_16510);
and U16804 (N_16804,N_16592,N_16740);
or U16805 (N_16805,N_16717,N_16613);
or U16806 (N_16806,N_16533,N_16580);
xor U16807 (N_16807,N_16634,N_16647);
nor U16808 (N_16808,N_16750,N_16758);
and U16809 (N_16809,N_16625,N_16705);
nor U16810 (N_16810,N_16681,N_16632);
and U16811 (N_16811,N_16517,N_16527);
xnor U16812 (N_16812,N_16711,N_16699);
or U16813 (N_16813,N_16623,N_16574);
nor U16814 (N_16814,N_16668,N_16637);
and U16815 (N_16815,N_16511,N_16566);
xnor U16816 (N_16816,N_16621,N_16604);
and U16817 (N_16817,N_16701,N_16713);
xor U16818 (N_16818,N_16551,N_16596);
nand U16819 (N_16819,N_16591,N_16691);
nor U16820 (N_16820,N_16789,N_16718);
nor U16821 (N_16821,N_16757,N_16512);
or U16822 (N_16822,N_16546,N_16519);
or U16823 (N_16823,N_16531,N_16535);
or U16824 (N_16824,N_16728,N_16619);
and U16825 (N_16825,N_16693,N_16640);
and U16826 (N_16826,N_16501,N_16635);
nor U16827 (N_16827,N_16725,N_16781);
or U16828 (N_16828,N_16651,N_16542);
and U16829 (N_16829,N_16714,N_16582);
nor U16830 (N_16830,N_16570,N_16552);
xor U16831 (N_16831,N_16617,N_16532);
nor U16832 (N_16832,N_16667,N_16661);
xnor U16833 (N_16833,N_16553,N_16684);
nor U16834 (N_16834,N_16727,N_16583);
or U16835 (N_16835,N_16769,N_16572);
or U16836 (N_16836,N_16610,N_16694);
xor U16837 (N_16837,N_16504,N_16629);
or U16838 (N_16838,N_16521,N_16639);
and U16839 (N_16839,N_16520,N_16739);
and U16840 (N_16840,N_16587,N_16584);
nand U16841 (N_16841,N_16654,N_16518);
and U16842 (N_16842,N_16522,N_16579);
nor U16843 (N_16843,N_16503,N_16611);
nand U16844 (N_16844,N_16607,N_16773);
or U16845 (N_16845,N_16720,N_16628);
and U16846 (N_16846,N_16581,N_16799);
and U16847 (N_16847,N_16779,N_16686);
nand U16848 (N_16848,N_16687,N_16790);
nand U16849 (N_16849,N_16756,N_16703);
or U16850 (N_16850,N_16753,N_16509);
xnor U16851 (N_16851,N_16588,N_16704);
xnor U16852 (N_16852,N_16762,N_16768);
and U16853 (N_16853,N_16692,N_16741);
and U16854 (N_16854,N_16657,N_16658);
nand U16855 (N_16855,N_16601,N_16759);
xnor U16856 (N_16856,N_16672,N_16733);
nand U16857 (N_16857,N_16645,N_16752);
or U16858 (N_16858,N_16760,N_16612);
or U16859 (N_16859,N_16547,N_16770);
nand U16860 (N_16860,N_16502,N_16615);
xnor U16861 (N_16861,N_16751,N_16538);
nor U16862 (N_16862,N_16543,N_16630);
nor U16863 (N_16863,N_16641,N_16797);
or U16864 (N_16864,N_16721,N_16598);
nand U16865 (N_16865,N_16743,N_16794);
or U16866 (N_16866,N_16563,N_16669);
nand U16867 (N_16867,N_16676,N_16549);
nor U16868 (N_16868,N_16695,N_16710);
nand U16869 (N_16869,N_16515,N_16576);
nand U16870 (N_16870,N_16569,N_16608);
or U16871 (N_16871,N_16698,N_16772);
nand U16872 (N_16872,N_16568,N_16586);
nand U16873 (N_16873,N_16792,N_16594);
nor U16874 (N_16874,N_16787,N_16665);
nor U16875 (N_16875,N_16674,N_16774);
and U16876 (N_16876,N_16545,N_16777);
and U16877 (N_16877,N_16791,N_16724);
nor U16878 (N_16878,N_16735,N_16776);
xor U16879 (N_16879,N_16622,N_16675);
nand U16880 (N_16880,N_16561,N_16648);
nor U16881 (N_16881,N_16761,N_16633);
nor U16882 (N_16882,N_16614,N_16706);
xnor U16883 (N_16883,N_16644,N_16508);
nand U16884 (N_16884,N_16567,N_16620);
nor U16885 (N_16885,N_16631,N_16626);
or U16886 (N_16886,N_16559,N_16529);
xor U16887 (N_16887,N_16775,N_16603);
and U16888 (N_16888,N_16593,N_16537);
nand U16889 (N_16889,N_16742,N_16793);
nor U16890 (N_16890,N_16573,N_16500);
nand U16891 (N_16891,N_16784,N_16700);
nand U16892 (N_16892,N_16578,N_16778);
nor U16893 (N_16893,N_16764,N_16548);
and U16894 (N_16894,N_16738,N_16534);
and U16895 (N_16895,N_16564,N_16719);
nand U16896 (N_16896,N_16562,N_16679);
nor U16897 (N_16897,N_16526,N_16677);
or U16898 (N_16898,N_16732,N_16663);
xnor U16899 (N_16899,N_16715,N_16656);
nor U16900 (N_16900,N_16590,N_16506);
and U16901 (N_16901,N_16540,N_16530);
nor U16902 (N_16902,N_16688,N_16744);
or U16903 (N_16903,N_16748,N_16765);
and U16904 (N_16904,N_16507,N_16541);
xor U16905 (N_16905,N_16731,N_16666);
nand U16906 (N_16906,N_16655,N_16505);
xnor U16907 (N_16907,N_16659,N_16771);
xnor U16908 (N_16908,N_16514,N_16606);
xor U16909 (N_16909,N_16716,N_16729);
or U16910 (N_16910,N_16571,N_16660);
nand U16911 (N_16911,N_16600,N_16638);
nor U16912 (N_16912,N_16642,N_16746);
nand U16913 (N_16913,N_16798,N_16755);
and U16914 (N_16914,N_16577,N_16708);
and U16915 (N_16915,N_16736,N_16682);
nor U16916 (N_16916,N_16585,N_16653);
nand U16917 (N_16917,N_16550,N_16780);
xor U16918 (N_16918,N_16595,N_16618);
nand U16919 (N_16919,N_16523,N_16767);
nand U16920 (N_16920,N_16680,N_16513);
nor U16921 (N_16921,N_16599,N_16516);
nor U16922 (N_16922,N_16690,N_16670);
xor U16923 (N_16923,N_16722,N_16560);
or U16924 (N_16924,N_16597,N_16747);
and U16925 (N_16925,N_16734,N_16528);
nor U16926 (N_16926,N_16685,N_16652);
and U16927 (N_16927,N_16795,N_16605);
and U16928 (N_16928,N_16602,N_16783);
and U16929 (N_16929,N_16671,N_16627);
nor U16930 (N_16930,N_16737,N_16689);
nor U16931 (N_16931,N_16749,N_16678);
xnor U16932 (N_16932,N_16558,N_16726);
and U16933 (N_16933,N_16650,N_16556);
or U16934 (N_16934,N_16664,N_16589);
or U16935 (N_16935,N_16555,N_16707);
nor U16936 (N_16936,N_16565,N_16723);
nand U16937 (N_16937,N_16683,N_16796);
nor U16938 (N_16938,N_16524,N_16646);
nand U16939 (N_16939,N_16544,N_16673);
nor U16940 (N_16940,N_16662,N_16616);
or U16941 (N_16941,N_16636,N_16754);
nand U16942 (N_16942,N_16745,N_16609);
and U16943 (N_16943,N_16712,N_16788);
and U16944 (N_16944,N_16697,N_16539);
and U16945 (N_16945,N_16554,N_16575);
nor U16946 (N_16946,N_16786,N_16536);
nand U16947 (N_16947,N_16525,N_16696);
xnor U16948 (N_16948,N_16557,N_16702);
xor U16949 (N_16949,N_16766,N_16785);
xnor U16950 (N_16950,N_16630,N_16679);
and U16951 (N_16951,N_16633,N_16591);
nand U16952 (N_16952,N_16754,N_16542);
or U16953 (N_16953,N_16657,N_16798);
nor U16954 (N_16954,N_16789,N_16647);
and U16955 (N_16955,N_16733,N_16665);
nand U16956 (N_16956,N_16605,N_16602);
nand U16957 (N_16957,N_16569,N_16642);
nand U16958 (N_16958,N_16600,N_16582);
and U16959 (N_16959,N_16763,N_16711);
nand U16960 (N_16960,N_16758,N_16794);
nor U16961 (N_16961,N_16702,N_16634);
xnor U16962 (N_16962,N_16507,N_16759);
and U16963 (N_16963,N_16602,N_16653);
nor U16964 (N_16964,N_16559,N_16632);
or U16965 (N_16965,N_16727,N_16531);
or U16966 (N_16966,N_16799,N_16718);
and U16967 (N_16967,N_16500,N_16567);
or U16968 (N_16968,N_16718,N_16563);
xor U16969 (N_16969,N_16753,N_16554);
xor U16970 (N_16970,N_16614,N_16529);
nor U16971 (N_16971,N_16537,N_16705);
nor U16972 (N_16972,N_16583,N_16590);
nor U16973 (N_16973,N_16564,N_16591);
and U16974 (N_16974,N_16777,N_16770);
xor U16975 (N_16975,N_16627,N_16587);
nand U16976 (N_16976,N_16617,N_16527);
xnor U16977 (N_16977,N_16595,N_16737);
xnor U16978 (N_16978,N_16549,N_16527);
or U16979 (N_16979,N_16790,N_16556);
or U16980 (N_16980,N_16516,N_16512);
or U16981 (N_16981,N_16644,N_16623);
or U16982 (N_16982,N_16687,N_16583);
or U16983 (N_16983,N_16533,N_16546);
nor U16984 (N_16984,N_16514,N_16588);
xnor U16985 (N_16985,N_16544,N_16614);
nand U16986 (N_16986,N_16548,N_16606);
or U16987 (N_16987,N_16580,N_16646);
nand U16988 (N_16988,N_16689,N_16783);
xnor U16989 (N_16989,N_16667,N_16556);
xor U16990 (N_16990,N_16676,N_16736);
nand U16991 (N_16991,N_16679,N_16585);
nor U16992 (N_16992,N_16694,N_16707);
nand U16993 (N_16993,N_16761,N_16714);
xnor U16994 (N_16994,N_16611,N_16567);
nand U16995 (N_16995,N_16628,N_16502);
and U16996 (N_16996,N_16549,N_16627);
or U16997 (N_16997,N_16734,N_16673);
nand U16998 (N_16998,N_16609,N_16533);
and U16999 (N_16999,N_16702,N_16539);
nand U17000 (N_17000,N_16651,N_16591);
nor U17001 (N_17001,N_16677,N_16533);
nor U17002 (N_17002,N_16745,N_16787);
or U17003 (N_17003,N_16573,N_16710);
nand U17004 (N_17004,N_16747,N_16662);
nand U17005 (N_17005,N_16701,N_16750);
and U17006 (N_17006,N_16760,N_16595);
nor U17007 (N_17007,N_16689,N_16747);
nor U17008 (N_17008,N_16552,N_16778);
and U17009 (N_17009,N_16733,N_16683);
nor U17010 (N_17010,N_16778,N_16772);
and U17011 (N_17011,N_16617,N_16518);
nor U17012 (N_17012,N_16514,N_16752);
and U17013 (N_17013,N_16700,N_16516);
xnor U17014 (N_17014,N_16618,N_16701);
xor U17015 (N_17015,N_16683,N_16602);
xor U17016 (N_17016,N_16524,N_16656);
nand U17017 (N_17017,N_16787,N_16509);
and U17018 (N_17018,N_16737,N_16784);
nand U17019 (N_17019,N_16790,N_16696);
nand U17020 (N_17020,N_16672,N_16533);
and U17021 (N_17021,N_16555,N_16574);
nor U17022 (N_17022,N_16510,N_16616);
and U17023 (N_17023,N_16503,N_16705);
nand U17024 (N_17024,N_16789,N_16537);
or U17025 (N_17025,N_16670,N_16774);
nand U17026 (N_17026,N_16791,N_16780);
nand U17027 (N_17027,N_16671,N_16769);
nand U17028 (N_17028,N_16597,N_16726);
and U17029 (N_17029,N_16500,N_16730);
nor U17030 (N_17030,N_16618,N_16655);
xor U17031 (N_17031,N_16731,N_16611);
or U17032 (N_17032,N_16761,N_16573);
or U17033 (N_17033,N_16655,N_16753);
or U17034 (N_17034,N_16501,N_16741);
nor U17035 (N_17035,N_16686,N_16652);
xnor U17036 (N_17036,N_16523,N_16718);
nor U17037 (N_17037,N_16562,N_16709);
and U17038 (N_17038,N_16703,N_16622);
or U17039 (N_17039,N_16673,N_16644);
or U17040 (N_17040,N_16711,N_16709);
and U17041 (N_17041,N_16767,N_16527);
nand U17042 (N_17042,N_16501,N_16648);
and U17043 (N_17043,N_16632,N_16512);
xnor U17044 (N_17044,N_16541,N_16769);
or U17045 (N_17045,N_16782,N_16612);
nor U17046 (N_17046,N_16546,N_16700);
or U17047 (N_17047,N_16696,N_16737);
nor U17048 (N_17048,N_16605,N_16785);
xor U17049 (N_17049,N_16794,N_16723);
or U17050 (N_17050,N_16629,N_16718);
nand U17051 (N_17051,N_16500,N_16557);
nor U17052 (N_17052,N_16740,N_16695);
xor U17053 (N_17053,N_16555,N_16549);
nand U17054 (N_17054,N_16774,N_16565);
nor U17055 (N_17055,N_16537,N_16613);
and U17056 (N_17056,N_16758,N_16760);
xnor U17057 (N_17057,N_16729,N_16712);
xor U17058 (N_17058,N_16627,N_16748);
or U17059 (N_17059,N_16524,N_16739);
or U17060 (N_17060,N_16668,N_16725);
nor U17061 (N_17061,N_16618,N_16585);
nand U17062 (N_17062,N_16531,N_16728);
nor U17063 (N_17063,N_16678,N_16515);
or U17064 (N_17064,N_16693,N_16601);
xnor U17065 (N_17065,N_16546,N_16670);
or U17066 (N_17066,N_16729,N_16500);
xor U17067 (N_17067,N_16736,N_16653);
xnor U17068 (N_17068,N_16792,N_16616);
or U17069 (N_17069,N_16730,N_16509);
nand U17070 (N_17070,N_16752,N_16565);
and U17071 (N_17071,N_16684,N_16518);
xor U17072 (N_17072,N_16549,N_16591);
xor U17073 (N_17073,N_16720,N_16699);
nand U17074 (N_17074,N_16648,N_16693);
or U17075 (N_17075,N_16669,N_16547);
or U17076 (N_17076,N_16580,N_16523);
and U17077 (N_17077,N_16530,N_16754);
nand U17078 (N_17078,N_16739,N_16615);
and U17079 (N_17079,N_16562,N_16545);
and U17080 (N_17080,N_16650,N_16586);
or U17081 (N_17081,N_16642,N_16602);
xnor U17082 (N_17082,N_16655,N_16578);
xnor U17083 (N_17083,N_16539,N_16753);
nand U17084 (N_17084,N_16686,N_16726);
and U17085 (N_17085,N_16529,N_16762);
xnor U17086 (N_17086,N_16590,N_16576);
or U17087 (N_17087,N_16642,N_16781);
or U17088 (N_17088,N_16529,N_16672);
nor U17089 (N_17089,N_16657,N_16683);
nand U17090 (N_17090,N_16745,N_16554);
xor U17091 (N_17091,N_16505,N_16568);
and U17092 (N_17092,N_16727,N_16685);
or U17093 (N_17093,N_16624,N_16512);
nand U17094 (N_17094,N_16669,N_16740);
or U17095 (N_17095,N_16660,N_16710);
nor U17096 (N_17096,N_16631,N_16646);
and U17097 (N_17097,N_16559,N_16570);
or U17098 (N_17098,N_16791,N_16541);
nand U17099 (N_17099,N_16508,N_16711);
xnor U17100 (N_17100,N_17038,N_16852);
and U17101 (N_17101,N_16854,N_16889);
or U17102 (N_17102,N_16943,N_16935);
and U17103 (N_17103,N_16842,N_17016);
or U17104 (N_17104,N_16834,N_16932);
nor U17105 (N_17105,N_17014,N_17015);
and U17106 (N_17106,N_17059,N_17075);
nand U17107 (N_17107,N_16989,N_17000);
or U17108 (N_17108,N_16976,N_16864);
xnor U17109 (N_17109,N_16964,N_16924);
and U17110 (N_17110,N_17008,N_17006);
nand U17111 (N_17111,N_17087,N_16868);
xnor U17112 (N_17112,N_16961,N_17001);
and U17113 (N_17113,N_16907,N_16917);
nor U17114 (N_17114,N_16826,N_16905);
or U17115 (N_17115,N_16914,N_16890);
nor U17116 (N_17116,N_16936,N_16880);
and U17117 (N_17117,N_16911,N_17035);
xor U17118 (N_17118,N_17093,N_16993);
nor U17119 (N_17119,N_16865,N_17071);
xor U17120 (N_17120,N_16982,N_16830);
nand U17121 (N_17121,N_16903,N_16853);
or U17122 (N_17122,N_17081,N_17041);
and U17123 (N_17123,N_17026,N_16920);
xor U17124 (N_17124,N_16828,N_16848);
nor U17125 (N_17125,N_16887,N_16840);
or U17126 (N_17126,N_17094,N_16858);
or U17127 (N_17127,N_17031,N_17002);
nand U17128 (N_17128,N_17019,N_16838);
nor U17129 (N_17129,N_16994,N_16856);
or U17130 (N_17130,N_16869,N_16958);
nand U17131 (N_17131,N_16908,N_16851);
nand U17132 (N_17132,N_16934,N_16845);
xnor U17133 (N_17133,N_17078,N_16921);
nand U17134 (N_17134,N_17052,N_16849);
nor U17135 (N_17135,N_16997,N_17063);
nor U17136 (N_17136,N_16983,N_16813);
nor U17137 (N_17137,N_16876,N_16872);
and U17138 (N_17138,N_17057,N_16954);
xor U17139 (N_17139,N_16843,N_16927);
nor U17140 (N_17140,N_16901,N_16896);
xnor U17141 (N_17141,N_16817,N_16801);
or U17142 (N_17142,N_16839,N_16945);
or U17143 (N_17143,N_17045,N_16923);
xnor U17144 (N_17144,N_16915,N_17089);
nor U17145 (N_17145,N_16850,N_16892);
nand U17146 (N_17146,N_16803,N_16971);
or U17147 (N_17147,N_16871,N_16878);
xor U17148 (N_17148,N_16944,N_16991);
nor U17149 (N_17149,N_16916,N_16968);
nand U17150 (N_17150,N_16940,N_16855);
xnor U17151 (N_17151,N_16884,N_16955);
xor U17152 (N_17152,N_17090,N_17027);
xnor U17153 (N_17153,N_17053,N_16980);
and U17154 (N_17154,N_17049,N_16926);
nor U17155 (N_17155,N_17009,N_16898);
or U17156 (N_17156,N_16981,N_16918);
xnor U17157 (N_17157,N_16912,N_16883);
xor U17158 (N_17158,N_16930,N_17036);
and U17159 (N_17159,N_17065,N_16816);
nand U17160 (N_17160,N_17047,N_17091);
nor U17161 (N_17161,N_16992,N_16860);
and U17162 (N_17162,N_17097,N_16942);
xor U17163 (N_17163,N_16806,N_16904);
nand U17164 (N_17164,N_16891,N_17029);
xnor U17165 (N_17165,N_16861,N_16953);
xor U17166 (N_17166,N_16900,N_16802);
xnor U17167 (N_17167,N_16928,N_17018);
xnor U17168 (N_17168,N_16881,N_17099);
and U17169 (N_17169,N_16822,N_16846);
xor U17170 (N_17170,N_16824,N_16882);
and U17171 (N_17171,N_17066,N_16913);
xnor U17172 (N_17172,N_17060,N_17023);
or U17173 (N_17173,N_16974,N_16835);
and U17174 (N_17174,N_16873,N_16877);
or U17175 (N_17175,N_17054,N_16949);
nand U17176 (N_17176,N_16965,N_16844);
xor U17177 (N_17177,N_17025,N_16823);
xor U17178 (N_17178,N_16922,N_16885);
xnor U17179 (N_17179,N_16893,N_17042);
xor U17180 (N_17180,N_17077,N_17044);
xnor U17181 (N_17181,N_16899,N_16820);
xor U17182 (N_17182,N_17068,N_16888);
nor U17183 (N_17183,N_17088,N_17048);
or U17184 (N_17184,N_17061,N_17004);
xnor U17185 (N_17185,N_16959,N_16939);
nand U17186 (N_17186,N_16807,N_16967);
and U17187 (N_17187,N_16894,N_16919);
and U17188 (N_17188,N_17074,N_16951);
xor U17189 (N_17189,N_16812,N_16870);
nand U17190 (N_17190,N_17076,N_17095);
or U17191 (N_17191,N_16875,N_17032);
or U17192 (N_17192,N_17092,N_16978);
nand U17193 (N_17193,N_16909,N_16833);
or U17194 (N_17194,N_16947,N_16975);
nor U17195 (N_17195,N_16941,N_17080);
xnor U17196 (N_17196,N_17067,N_16809);
or U17197 (N_17197,N_16979,N_17050);
xnor U17198 (N_17198,N_17013,N_16929);
nand U17199 (N_17199,N_17024,N_16847);
nor U17200 (N_17200,N_17098,N_16952);
xnor U17201 (N_17201,N_16910,N_17096);
xor U17202 (N_17202,N_16886,N_16999);
and U17203 (N_17203,N_16973,N_16966);
or U17204 (N_17204,N_17010,N_16859);
and U17205 (N_17205,N_16977,N_16819);
nor U17206 (N_17206,N_17058,N_16831);
and U17207 (N_17207,N_17073,N_16810);
and U17208 (N_17208,N_16879,N_16933);
or U17209 (N_17209,N_16874,N_17028);
or U17210 (N_17210,N_16837,N_16946);
and U17211 (N_17211,N_17034,N_16825);
nand U17212 (N_17212,N_16985,N_16948);
nand U17213 (N_17213,N_17084,N_16937);
nand U17214 (N_17214,N_16962,N_17082);
and U17215 (N_17215,N_17017,N_16800);
xnor U17216 (N_17216,N_16987,N_17085);
xnor U17217 (N_17217,N_16957,N_16897);
xnor U17218 (N_17218,N_17037,N_16938);
xor U17219 (N_17219,N_16827,N_16986);
nor U17220 (N_17220,N_16867,N_17007);
nand U17221 (N_17221,N_17064,N_16990);
nand U17222 (N_17222,N_16969,N_17062);
or U17223 (N_17223,N_17069,N_17003);
nand U17224 (N_17224,N_16862,N_16970);
or U17225 (N_17225,N_17079,N_17040);
nand U17226 (N_17226,N_16821,N_17020);
xor U17227 (N_17227,N_16906,N_16857);
xnor U17228 (N_17228,N_16895,N_17022);
and U17229 (N_17229,N_16811,N_16984);
xnor U17230 (N_17230,N_16960,N_16995);
nor U17231 (N_17231,N_17046,N_16902);
or U17232 (N_17232,N_17005,N_16815);
or U17233 (N_17233,N_16836,N_17043);
or U17234 (N_17234,N_17083,N_16988);
or U17235 (N_17235,N_17021,N_16832);
nand U17236 (N_17236,N_16863,N_17055);
nor U17237 (N_17237,N_16804,N_17039);
nand U17238 (N_17238,N_16866,N_16805);
nand U17239 (N_17239,N_16925,N_16956);
nor U17240 (N_17240,N_16808,N_16829);
xnor U17241 (N_17241,N_16814,N_17051);
or U17242 (N_17242,N_16998,N_17072);
and U17243 (N_17243,N_17011,N_17030);
or U17244 (N_17244,N_16996,N_17070);
xor U17245 (N_17245,N_16963,N_17012);
or U17246 (N_17246,N_16818,N_17086);
nand U17247 (N_17247,N_16950,N_16972);
nand U17248 (N_17248,N_17056,N_16931);
xnor U17249 (N_17249,N_17033,N_16841);
and U17250 (N_17250,N_17088,N_16944);
nand U17251 (N_17251,N_17045,N_16812);
and U17252 (N_17252,N_16803,N_16924);
xnor U17253 (N_17253,N_17057,N_17050);
nor U17254 (N_17254,N_16891,N_17068);
or U17255 (N_17255,N_16879,N_17098);
and U17256 (N_17256,N_17034,N_17023);
nand U17257 (N_17257,N_16969,N_16880);
or U17258 (N_17258,N_16850,N_17002);
nor U17259 (N_17259,N_17088,N_16979);
or U17260 (N_17260,N_17000,N_16997);
nor U17261 (N_17261,N_16957,N_16931);
or U17262 (N_17262,N_17058,N_16983);
and U17263 (N_17263,N_17045,N_16974);
xor U17264 (N_17264,N_16894,N_16809);
or U17265 (N_17265,N_16965,N_16827);
nand U17266 (N_17266,N_16955,N_16948);
nor U17267 (N_17267,N_16988,N_16922);
and U17268 (N_17268,N_16861,N_16854);
nor U17269 (N_17269,N_16814,N_16948);
xor U17270 (N_17270,N_16902,N_16941);
nor U17271 (N_17271,N_16887,N_16832);
nor U17272 (N_17272,N_16948,N_16820);
xnor U17273 (N_17273,N_16987,N_16941);
and U17274 (N_17274,N_16821,N_16903);
nand U17275 (N_17275,N_16854,N_16943);
xnor U17276 (N_17276,N_16810,N_17068);
or U17277 (N_17277,N_16981,N_16978);
xor U17278 (N_17278,N_17021,N_16805);
or U17279 (N_17279,N_17038,N_17058);
nor U17280 (N_17280,N_16804,N_17060);
or U17281 (N_17281,N_16893,N_16978);
nand U17282 (N_17282,N_17082,N_17032);
nor U17283 (N_17283,N_17019,N_17021);
nor U17284 (N_17284,N_16954,N_17046);
xnor U17285 (N_17285,N_16851,N_16961);
nor U17286 (N_17286,N_16865,N_17023);
nand U17287 (N_17287,N_16928,N_16847);
nand U17288 (N_17288,N_16852,N_16974);
or U17289 (N_17289,N_16850,N_16877);
and U17290 (N_17290,N_17081,N_17075);
xnor U17291 (N_17291,N_17072,N_16991);
xnor U17292 (N_17292,N_16966,N_17028);
xor U17293 (N_17293,N_16893,N_16953);
nand U17294 (N_17294,N_17059,N_16809);
or U17295 (N_17295,N_16836,N_16834);
or U17296 (N_17296,N_16866,N_17066);
nor U17297 (N_17297,N_16892,N_17047);
or U17298 (N_17298,N_17075,N_16806);
xor U17299 (N_17299,N_17021,N_17037);
nor U17300 (N_17300,N_16961,N_16812);
and U17301 (N_17301,N_16915,N_16919);
or U17302 (N_17302,N_16997,N_17087);
nand U17303 (N_17303,N_17026,N_17028);
xnor U17304 (N_17304,N_16849,N_16902);
nor U17305 (N_17305,N_17043,N_17049);
and U17306 (N_17306,N_16954,N_17073);
and U17307 (N_17307,N_16874,N_16825);
nand U17308 (N_17308,N_16830,N_17051);
xnor U17309 (N_17309,N_16999,N_16918);
nand U17310 (N_17310,N_16849,N_16900);
or U17311 (N_17311,N_17010,N_17086);
or U17312 (N_17312,N_16899,N_17076);
nor U17313 (N_17313,N_17092,N_17076);
xor U17314 (N_17314,N_17068,N_16952);
nor U17315 (N_17315,N_17087,N_16817);
xor U17316 (N_17316,N_17052,N_16800);
nor U17317 (N_17317,N_16885,N_16824);
nand U17318 (N_17318,N_16931,N_16956);
and U17319 (N_17319,N_16985,N_16879);
and U17320 (N_17320,N_17051,N_17033);
xnor U17321 (N_17321,N_17004,N_16949);
xor U17322 (N_17322,N_16887,N_16907);
xor U17323 (N_17323,N_16991,N_16850);
xnor U17324 (N_17324,N_16872,N_16855);
and U17325 (N_17325,N_17067,N_17063);
xnor U17326 (N_17326,N_17091,N_17096);
nor U17327 (N_17327,N_17037,N_17065);
or U17328 (N_17328,N_16840,N_17058);
or U17329 (N_17329,N_17008,N_17060);
and U17330 (N_17330,N_16908,N_17005);
and U17331 (N_17331,N_16894,N_17095);
nor U17332 (N_17332,N_16853,N_16812);
xor U17333 (N_17333,N_16967,N_16892);
xnor U17334 (N_17334,N_16942,N_17035);
or U17335 (N_17335,N_17078,N_16995);
nor U17336 (N_17336,N_16946,N_17009);
nand U17337 (N_17337,N_16897,N_17079);
or U17338 (N_17338,N_17088,N_16958);
and U17339 (N_17339,N_16898,N_16879);
xnor U17340 (N_17340,N_16811,N_17056);
nand U17341 (N_17341,N_16855,N_16917);
nand U17342 (N_17342,N_16824,N_17041);
or U17343 (N_17343,N_16827,N_16993);
xor U17344 (N_17344,N_16966,N_17070);
and U17345 (N_17345,N_16825,N_16881);
or U17346 (N_17346,N_17042,N_16853);
nor U17347 (N_17347,N_16941,N_16934);
and U17348 (N_17348,N_16937,N_16924);
and U17349 (N_17349,N_16802,N_17037);
and U17350 (N_17350,N_16938,N_16990);
xor U17351 (N_17351,N_16832,N_17027);
nor U17352 (N_17352,N_16849,N_16997);
or U17353 (N_17353,N_16808,N_16904);
nand U17354 (N_17354,N_16967,N_17031);
and U17355 (N_17355,N_16857,N_16890);
or U17356 (N_17356,N_16983,N_17027);
nor U17357 (N_17357,N_16902,N_16938);
nand U17358 (N_17358,N_17085,N_16917);
nor U17359 (N_17359,N_16828,N_16900);
xnor U17360 (N_17360,N_16859,N_16875);
nand U17361 (N_17361,N_16873,N_16986);
or U17362 (N_17362,N_16948,N_16861);
xnor U17363 (N_17363,N_16865,N_16889);
and U17364 (N_17364,N_16834,N_16853);
nand U17365 (N_17365,N_16988,N_16967);
nand U17366 (N_17366,N_16818,N_16862);
xor U17367 (N_17367,N_16834,N_16974);
xnor U17368 (N_17368,N_16886,N_16889);
nor U17369 (N_17369,N_17081,N_16803);
and U17370 (N_17370,N_16836,N_16980);
nor U17371 (N_17371,N_17082,N_16895);
nor U17372 (N_17372,N_16986,N_16837);
xnor U17373 (N_17373,N_16834,N_16965);
or U17374 (N_17374,N_16831,N_17084);
or U17375 (N_17375,N_16909,N_16992);
nor U17376 (N_17376,N_17069,N_17008);
or U17377 (N_17377,N_17058,N_16981);
nand U17378 (N_17378,N_16929,N_16996);
nand U17379 (N_17379,N_16997,N_16879);
xnor U17380 (N_17380,N_16987,N_16839);
nand U17381 (N_17381,N_16887,N_16818);
nand U17382 (N_17382,N_16872,N_17026);
or U17383 (N_17383,N_16877,N_16931);
or U17384 (N_17384,N_16890,N_17034);
nand U17385 (N_17385,N_17023,N_16894);
nand U17386 (N_17386,N_17046,N_16889);
and U17387 (N_17387,N_16823,N_17031);
or U17388 (N_17388,N_16931,N_16991);
and U17389 (N_17389,N_16989,N_17094);
and U17390 (N_17390,N_16860,N_17052);
xnor U17391 (N_17391,N_16991,N_17055);
nor U17392 (N_17392,N_17071,N_16979);
nor U17393 (N_17393,N_17029,N_17051);
nor U17394 (N_17394,N_17033,N_16955);
nand U17395 (N_17395,N_16800,N_16860);
or U17396 (N_17396,N_17002,N_17056);
or U17397 (N_17397,N_17019,N_16809);
or U17398 (N_17398,N_16894,N_16823);
xor U17399 (N_17399,N_17086,N_17009);
xor U17400 (N_17400,N_17214,N_17266);
xnor U17401 (N_17401,N_17257,N_17207);
nand U17402 (N_17402,N_17305,N_17116);
xnor U17403 (N_17403,N_17195,N_17221);
and U17404 (N_17404,N_17242,N_17275);
and U17405 (N_17405,N_17182,N_17322);
and U17406 (N_17406,N_17291,N_17357);
nor U17407 (N_17407,N_17235,N_17294);
nand U17408 (N_17408,N_17329,N_17339);
nor U17409 (N_17409,N_17303,N_17215);
xor U17410 (N_17410,N_17114,N_17184);
nand U17411 (N_17411,N_17300,N_17175);
and U17412 (N_17412,N_17335,N_17281);
nor U17413 (N_17413,N_17364,N_17171);
or U17414 (N_17414,N_17234,N_17302);
nand U17415 (N_17415,N_17177,N_17192);
xnor U17416 (N_17416,N_17336,N_17133);
xnor U17417 (N_17417,N_17129,N_17155);
and U17418 (N_17418,N_17220,N_17157);
xor U17419 (N_17419,N_17280,N_17118);
nor U17420 (N_17420,N_17377,N_17333);
and U17421 (N_17421,N_17135,N_17397);
nor U17422 (N_17422,N_17272,N_17313);
nand U17423 (N_17423,N_17340,N_17354);
nand U17424 (N_17424,N_17131,N_17104);
xnor U17425 (N_17425,N_17251,N_17295);
nand U17426 (N_17426,N_17117,N_17170);
and U17427 (N_17427,N_17122,N_17359);
or U17428 (N_17428,N_17211,N_17209);
xor U17429 (N_17429,N_17230,N_17350);
and U17430 (N_17430,N_17115,N_17130);
or U17431 (N_17431,N_17186,N_17226);
and U17432 (N_17432,N_17102,N_17173);
xnor U17433 (N_17433,N_17347,N_17101);
nor U17434 (N_17434,N_17153,N_17236);
and U17435 (N_17435,N_17199,N_17316);
and U17436 (N_17436,N_17204,N_17373);
nor U17437 (N_17437,N_17306,N_17341);
and U17438 (N_17438,N_17140,N_17298);
and U17439 (N_17439,N_17189,N_17164);
and U17440 (N_17440,N_17197,N_17273);
and U17441 (N_17441,N_17307,N_17308);
nand U17442 (N_17442,N_17151,N_17371);
xnor U17443 (N_17443,N_17290,N_17139);
nand U17444 (N_17444,N_17161,N_17391);
nand U17445 (N_17445,N_17282,N_17386);
and U17446 (N_17446,N_17363,N_17247);
nor U17447 (N_17447,N_17200,N_17375);
and U17448 (N_17448,N_17178,N_17198);
and U17449 (N_17449,N_17240,N_17310);
or U17450 (N_17450,N_17219,N_17194);
nor U17451 (N_17451,N_17345,N_17202);
nand U17452 (N_17452,N_17121,N_17278);
nand U17453 (N_17453,N_17224,N_17119);
nor U17454 (N_17454,N_17260,N_17123);
nand U17455 (N_17455,N_17255,N_17328);
or U17456 (N_17456,N_17206,N_17398);
and U17457 (N_17457,N_17293,N_17387);
xnor U17458 (N_17458,N_17250,N_17396);
or U17459 (N_17459,N_17283,N_17180);
xor U17460 (N_17460,N_17124,N_17370);
nand U17461 (N_17461,N_17205,N_17355);
and U17462 (N_17462,N_17254,N_17261);
xnor U17463 (N_17463,N_17393,N_17154);
nor U17464 (N_17464,N_17143,N_17392);
and U17465 (N_17465,N_17125,N_17176);
xnor U17466 (N_17466,N_17120,N_17212);
xnor U17467 (N_17467,N_17142,N_17227);
and U17468 (N_17468,N_17188,N_17362);
and U17469 (N_17469,N_17208,N_17344);
xor U17470 (N_17470,N_17162,N_17150);
or U17471 (N_17471,N_17376,N_17323);
nor U17472 (N_17472,N_17286,N_17337);
xor U17473 (N_17473,N_17331,N_17243);
nor U17474 (N_17474,N_17353,N_17141);
or U17475 (N_17475,N_17320,N_17166);
and U17476 (N_17476,N_17126,N_17193);
or U17477 (N_17477,N_17265,N_17284);
nand U17478 (N_17478,N_17225,N_17379);
or U17479 (N_17479,N_17201,N_17338);
or U17480 (N_17480,N_17348,N_17128);
or U17481 (N_17481,N_17378,N_17145);
nor U17482 (N_17482,N_17304,N_17107);
or U17483 (N_17483,N_17366,N_17259);
xor U17484 (N_17484,N_17394,N_17358);
and U17485 (N_17485,N_17311,N_17105);
xnor U17486 (N_17486,N_17346,N_17382);
nand U17487 (N_17487,N_17203,N_17187);
and U17488 (N_17488,N_17269,N_17244);
nand U17489 (N_17489,N_17361,N_17268);
xnor U17490 (N_17490,N_17190,N_17314);
nand U17491 (N_17491,N_17390,N_17222);
xor U17492 (N_17492,N_17256,N_17174);
xor U17493 (N_17493,N_17330,N_17152);
or U17494 (N_17494,N_17301,N_17276);
nand U17495 (N_17495,N_17223,N_17318);
and U17496 (N_17496,N_17399,N_17110);
nand U17497 (N_17497,N_17332,N_17108);
nor U17498 (N_17498,N_17146,N_17299);
nand U17499 (N_17499,N_17309,N_17381);
nand U17500 (N_17500,N_17389,N_17137);
nor U17501 (N_17501,N_17132,N_17183);
nand U17502 (N_17502,N_17380,N_17279);
or U17503 (N_17503,N_17383,N_17109);
and U17504 (N_17504,N_17317,N_17384);
and U17505 (N_17505,N_17292,N_17385);
or U17506 (N_17506,N_17100,N_17232);
nand U17507 (N_17507,N_17315,N_17267);
and U17508 (N_17508,N_17271,N_17111);
xor U17509 (N_17509,N_17369,N_17325);
xnor U17510 (N_17510,N_17112,N_17165);
xnor U17511 (N_17511,N_17185,N_17368);
xor U17512 (N_17512,N_17210,N_17327);
and U17513 (N_17513,N_17274,N_17228);
and U17514 (N_17514,N_17253,N_17246);
or U17515 (N_17515,N_17106,N_17388);
nor U17516 (N_17516,N_17372,N_17277);
or U17517 (N_17517,N_17169,N_17245);
nand U17518 (N_17518,N_17326,N_17233);
and U17519 (N_17519,N_17365,N_17343);
nor U17520 (N_17520,N_17262,N_17156);
and U17521 (N_17521,N_17113,N_17296);
and U17522 (N_17522,N_17216,N_17231);
nand U17523 (N_17523,N_17168,N_17103);
nand U17524 (N_17524,N_17297,N_17264);
xor U17525 (N_17525,N_17351,N_17321);
or U17526 (N_17526,N_17312,N_17148);
xor U17527 (N_17527,N_17241,N_17229);
or U17528 (N_17528,N_17263,N_17319);
and U17529 (N_17529,N_17367,N_17342);
or U17530 (N_17530,N_17237,N_17158);
nand U17531 (N_17531,N_17352,N_17213);
and U17532 (N_17532,N_17196,N_17356);
xor U17533 (N_17533,N_17252,N_17149);
nand U17534 (N_17534,N_17172,N_17163);
nor U17535 (N_17535,N_17349,N_17249);
xnor U17536 (N_17536,N_17334,N_17167);
nor U17537 (N_17537,N_17134,N_17360);
xor U17538 (N_17538,N_17147,N_17288);
nand U17539 (N_17539,N_17144,N_17238);
nand U17540 (N_17540,N_17248,N_17239);
nand U17541 (N_17541,N_17285,N_17191);
nand U17542 (N_17542,N_17289,N_17218);
and U17543 (N_17543,N_17159,N_17395);
or U17544 (N_17544,N_17179,N_17374);
nor U17545 (N_17545,N_17127,N_17324);
xnor U17546 (N_17546,N_17160,N_17136);
or U17547 (N_17547,N_17287,N_17138);
xor U17548 (N_17548,N_17181,N_17270);
or U17549 (N_17549,N_17217,N_17258);
nor U17550 (N_17550,N_17294,N_17128);
xnor U17551 (N_17551,N_17275,N_17215);
xor U17552 (N_17552,N_17305,N_17169);
nand U17553 (N_17553,N_17134,N_17206);
or U17554 (N_17554,N_17128,N_17133);
xor U17555 (N_17555,N_17196,N_17116);
or U17556 (N_17556,N_17229,N_17342);
nor U17557 (N_17557,N_17132,N_17241);
xor U17558 (N_17558,N_17185,N_17367);
and U17559 (N_17559,N_17284,N_17129);
nand U17560 (N_17560,N_17129,N_17287);
nor U17561 (N_17561,N_17188,N_17293);
and U17562 (N_17562,N_17252,N_17208);
and U17563 (N_17563,N_17157,N_17375);
or U17564 (N_17564,N_17184,N_17282);
xor U17565 (N_17565,N_17212,N_17128);
or U17566 (N_17566,N_17303,N_17181);
and U17567 (N_17567,N_17286,N_17159);
xor U17568 (N_17568,N_17366,N_17315);
nand U17569 (N_17569,N_17261,N_17320);
or U17570 (N_17570,N_17191,N_17114);
nand U17571 (N_17571,N_17273,N_17188);
or U17572 (N_17572,N_17227,N_17298);
and U17573 (N_17573,N_17387,N_17238);
xor U17574 (N_17574,N_17223,N_17340);
nand U17575 (N_17575,N_17381,N_17310);
and U17576 (N_17576,N_17340,N_17375);
xnor U17577 (N_17577,N_17363,N_17368);
nand U17578 (N_17578,N_17116,N_17391);
and U17579 (N_17579,N_17117,N_17347);
nand U17580 (N_17580,N_17191,N_17345);
xnor U17581 (N_17581,N_17147,N_17304);
nor U17582 (N_17582,N_17220,N_17225);
xnor U17583 (N_17583,N_17180,N_17219);
or U17584 (N_17584,N_17106,N_17182);
nor U17585 (N_17585,N_17162,N_17240);
nand U17586 (N_17586,N_17197,N_17343);
and U17587 (N_17587,N_17135,N_17388);
or U17588 (N_17588,N_17221,N_17181);
xor U17589 (N_17589,N_17212,N_17147);
nand U17590 (N_17590,N_17300,N_17289);
and U17591 (N_17591,N_17165,N_17226);
nor U17592 (N_17592,N_17173,N_17344);
nand U17593 (N_17593,N_17263,N_17254);
nor U17594 (N_17594,N_17244,N_17295);
nand U17595 (N_17595,N_17350,N_17326);
xor U17596 (N_17596,N_17264,N_17191);
xnor U17597 (N_17597,N_17301,N_17302);
and U17598 (N_17598,N_17250,N_17355);
or U17599 (N_17599,N_17223,N_17300);
nor U17600 (N_17600,N_17240,N_17152);
nor U17601 (N_17601,N_17207,N_17287);
nor U17602 (N_17602,N_17234,N_17171);
nor U17603 (N_17603,N_17267,N_17230);
and U17604 (N_17604,N_17285,N_17271);
or U17605 (N_17605,N_17266,N_17391);
nor U17606 (N_17606,N_17129,N_17279);
nor U17607 (N_17607,N_17207,N_17302);
or U17608 (N_17608,N_17356,N_17114);
nor U17609 (N_17609,N_17253,N_17210);
or U17610 (N_17610,N_17306,N_17343);
or U17611 (N_17611,N_17230,N_17264);
and U17612 (N_17612,N_17131,N_17300);
nor U17613 (N_17613,N_17303,N_17378);
and U17614 (N_17614,N_17203,N_17160);
nand U17615 (N_17615,N_17275,N_17394);
nor U17616 (N_17616,N_17375,N_17213);
nor U17617 (N_17617,N_17302,N_17229);
xor U17618 (N_17618,N_17316,N_17379);
nand U17619 (N_17619,N_17380,N_17249);
nand U17620 (N_17620,N_17270,N_17290);
xnor U17621 (N_17621,N_17309,N_17278);
nand U17622 (N_17622,N_17273,N_17186);
nor U17623 (N_17623,N_17128,N_17330);
nand U17624 (N_17624,N_17264,N_17327);
nor U17625 (N_17625,N_17208,N_17121);
xor U17626 (N_17626,N_17398,N_17369);
and U17627 (N_17627,N_17155,N_17387);
or U17628 (N_17628,N_17313,N_17201);
nor U17629 (N_17629,N_17331,N_17237);
xor U17630 (N_17630,N_17247,N_17231);
nand U17631 (N_17631,N_17301,N_17345);
or U17632 (N_17632,N_17167,N_17263);
and U17633 (N_17633,N_17337,N_17352);
or U17634 (N_17634,N_17289,N_17179);
nand U17635 (N_17635,N_17213,N_17143);
and U17636 (N_17636,N_17146,N_17303);
xor U17637 (N_17637,N_17386,N_17263);
or U17638 (N_17638,N_17254,N_17265);
or U17639 (N_17639,N_17371,N_17126);
nand U17640 (N_17640,N_17343,N_17318);
nor U17641 (N_17641,N_17300,N_17297);
and U17642 (N_17642,N_17178,N_17347);
and U17643 (N_17643,N_17327,N_17325);
or U17644 (N_17644,N_17121,N_17318);
nor U17645 (N_17645,N_17376,N_17360);
nor U17646 (N_17646,N_17356,N_17299);
nand U17647 (N_17647,N_17186,N_17301);
nand U17648 (N_17648,N_17252,N_17128);
nor U17649 (N_17649,N_17248,N_17360);
xor U17650 (N_17650,N_17394,N_17292);
nor U17651 (N_17651,N_17241,N_17130);
or U17652 (N_17652,N_17294,N_17315);
nor U17653 (N_17653,N_17156,N_17243);
and U17654 (N_17654,N_17332,N_17282);
or U17655 (N_17655,N_17149,N_17266);
nor U17656 (N_17656,N_17212,N_17168);
or U17657 (N_17657,N_17381,N_17215);
or U17658 (N_17658,N_17251,N_17389);
nor U17659 (N_17659,N_17222,N_17283);
and U17660 (N_17660,N_17163,N_17318);
or U17661 (N_17661,N_17381,N_17253);
xor U17662 (N_17662,N_17375,N_17186);
or U17663 (N_17663,N_17124,N_17287);
and U17664 (N_17664,N_17111,N_17338);
or U17665 (N_17665,N_17221,N_17360);
and U17666 (N_17666,N_17229,N_17164);
nor U17667 (N_17667,N_17208,N_17375);
xor U17668 (N_17668,N_17191,N_17177);
and U17669 (N_17669,N_17392,N_17261);
nand U17670 (N_17670,N_17123,N_17180);
nand U17671 (N_17671,N_17302,N_17279);
and U17672 (N_17672,N_17218,N_17352);
nand U17673 (N_17673,N_17132,N_17209);
nor U17674 (N_17674,N_17165,N_17369);
or U17675 (N_17675,N_17275,N_17158);
xnor U17676 (N_17676,N_17199,N_17248);
and U17677 (N_17677,N_17293,N_17305);
xnor U17678 (N_17678,N_17239,N_17258);
nand U17679 (N_17679,N_17118,N_17379);
nor U17680 (N_17680,N_17144,N_17166);
and U17681 (N_17681,N_17123,N_17330);
nor U17682 (N_17682,N_17212,N_17230);
or U17683 (N_17683,N_17322,N_17126);
xor U17684 (N_17684,N_17184,N_17207);
nand U17685 (N_17685,N_17392,N_17346);
nand U17686 (N_17686,N_17122,N_17194);
and U17687 (N_17687,N_17393,N_17388);
nor U17688 (N_17688,N_17260,N_17194);
nand U17689 (N_17689,N_17185,N_17197);
xnor U17690 (N_17690,N_17357,N_17155);
nand U17691 (N_17691,N_17187,N_17270);
xor U17692 (N_17692,N_17189,N_17149);
xnor U17693 (N_17693,N_17271,N_17221);
nor U17694 (N_17694,N_17231,N_17186);
nor U17695 (N_17695,N_17105,N_17200);
nand U17696 (N_17696,N_17122,N_17319);
and U17697 (N_17697,N_17336,N_17152);
xnor U17698 (N_17698,N_17119,N_17322);
nand U17699 (N_17699,N_17272,N_17215);
and U17700 (N_17700,N_17697,N_17599);
nor U17701 (N_17701,N_17550,N_17416);
nor U17702 (N_17702,N_17598,N_17431);
xnor U17703 (N_17703,N_17661,N_17443);
or U17704 (N_17704,N_17514,N_17473);
nand U17705 (N_17705,N_17636,N_17666);
and U17706 (N_17706,N_17466,N_17492);
nand U17707 (N_17707,N_17604,N_17423);
or U17708 (N_17708,N_17678,N_17688);
or U17709 (N_17709,N_17699,N_17607);
nor U17710 (N_17710,N_17617,N_17642);
or U17711 (N_17711,N_17516,N_17451);
or U17712 (N_17712,N_17519,N_17408);
nor U17713 (N_17713,N_17583,N_17430);
nand U17714 (N_17714,N_17437,N_17694);
or U17715 (N_17715,N_17579,N_17648);
and U17716 (N_17716,N_17503,N_17655);
xor U17717 (N_17717,N_17439,N_17621);
or U17718 (N_17718,N_17400,N_17596);
xor U17719 (N_17719,N_17682,N_17549);
xnor U17720 (N_17720,N_17614,N_17402);
xnor U17721 (N_17721,N_17671,N_17421);
or U17722 (N_17722,N_17528,N_17662);
nor U17723 (N_17723,N_17411,N_17651);
nand U17724 (N_17724,N_17667,N_17649);
or U17725 (N_17725,N_17438,N_17568);
nand U17726 (N_17726,N_17417,N_17418);
or U17727 (N_17727,N_17446,N_17577);
or U17728 (N_17728,N_17447,N_17689);
nand U17729 (N_17729,N_17461,N_17687);
nor U17730 (N_17730,N_17640,N_17628);
or U17731 (N_17731,N_17660,N_17618);
or U17732 (N_17732,N_17581,N_17572);
nor U17733 (N_17733,N_17458,N_17523);
and U17734 (N_17734,N_17482,N_17542);
nand U17735 (N_17735,N_17559,N_17606);
nand U17736 (N_17736,N_17463,N_17454);
xnor U17737 (N_17737,N_17506,N_17683);
xor U17738 (N_17738,N_17448,N_17453);
xor U17739 (N_17739,N_17487,N_17539);
nor U17740 (N_17740,N_17459,N_17429);
xnor U17741 (N_17741,N_17403,N_17632);
or U17742 (N_17742,N_17610,N_17691);
xnor U17743 (N_17743,N_17603,N_17479);
and U17744 (N_17744,N_17543,N_17481);
or U17745 (N_17745,N_17552,N_17605);
nor U17746 (N_17746,N_17509,N_17538);
or U17747 (N_17747,N_17677,N_17452);
nor U17748 (N_17748,N_17582,N_17566);
nand U17749 (N_17749,N_17586,N_17483);
or U17750 (N_17750,N_17597,N_17450);
and U17751 (N_17751,N_17435,N_17609);
nand U17752 (N_17752,N_17695,N_17673);
xnor U17753 (N_17753,N_17544,N_17600);
xnor U17754 (N_17754,N_17415,N_17445);
and U17755 (N_17755,N_17536,N_17557);
nor U17756 (N_17756,N_17444,N_17647);
and U17757 (N_17757,N_17637,N_17626);
xnor U17758 (N_17758,N_17546,N_17629);
xnor U17759 (N_17759,N_17668,N_17410);
xnor U17760 (N_17760,N_17476,N_17526);
or U17761 (N_17761,N_17489,N_17571);
nor U17762 (N_17762,N_17592,N_17664);
and U17763 (N_17763,N_17434,N_17643);
or U17764 (N_17764,N_17422,N_17502);
nor U17765 (N_17765,N_17585,N_17471);
or U17766 (N_17766,N_17634,N_17513);
nor U17767 (N_17767,N_17404,N_17501);
xor U17768 (N_17768,N_17527,N_17558);
or U17769 (N_17769,N_17591,N_17428);
xor U17770 (N_17770,N_17669,N_17409);
and U17771 (N_17771,N_17407,N_17474);
xor U17772 (N_17772,N_17653,N_17674);
xor U17773 (N_17773,N_17574,N_17654);
or U17774 (N_17774,N_17525,N_17644);
xor U17775 (N_17775,N_17499,N_17573);
and U17776 (N_17776,N_17505,N_17681);
nand U17777 (N_17777,N_17455,N_17567);
nor U17778 (N_17778,N_17521,N_17560);
nand U17779 (N_17779,N_17530,N_17698);
and U17780 (N_17780,N_17493,N_17534);
and U17781 (N_17781,N_17464,N_17593);
nand U17782 (N_17782,N_17622,N_17612);
nor U17783 (N_17783,N_17569,N_17555);
and U17784 (N_17784,N_17531,N_17633);
and U17785 (N_17785,N_17401,N_17623);
or U17786 (N_17786,N_17627,N_17656);
and U17787 (N_17787,N_17578,N_17427);
nor U17788 (N_17788,N_17646,N_17684);
nand U17789 (N_17789,N_17672,N_17512);
nand U17790 (N_17790,N_17529,N_17561);
and U17791 (N_17791,N_17570,N_17497);
nor U17792 (N_17792,N_17545,N_17562);
and U17793 (N_17793,N_17470,N_17449);
or U17794 (N_17794,N_17620,N_17405);
xnor U17795 (N_17795,N_17520,N_17696);
xor U17796 (N_17796,N_17663,N_17426);
nand U17797 (N_17797,N_17680,N_17630);
or U17798 (N_17798,N_17478,N_17619);
or U17799 (N_17799,N_17495,N_17517);
or U17800 (N_17800,N_17485,N_17556);
xnor U17801 (N_17801,N_17608,N_17511);
nor U17802 (N_17802,N_17584,N_17413);
nor U17803 (N_17803,N_17486,N_17456);
or U17804 (N_17804,N_17522,N_17548);
nand U17805 (N_17805,N_17638,N_17679);
and U17806 (N_17806,N_17419,N_17665);
nand U17807 (N_17807,N_17554,N_17635);
nor U17808 (N_17808,N_17467,N_17564);
xnor U17809 (N_17809,N_17551,N_17650);
and U17810 (N_17810,N_17639,N_17686);
nand U17811 (N_17811,N_17657,N_17692);
nor U17812 (N_17812,N_17533,N_17414);
nand U17813 (N_17813,N_17504,N_17496);
nand U17814 (N_17814,N_17524,N_17468);
and U17815 (N_17815,N_17685,N_17424);
nor U17816 (N_17816,N_17469,N_17693);
nand U17817 (N_17817,N_17433,N_17675);
or U17818 (N_17818,N_17624,N_17477);
xor U17819 (N_17819,N_17588,N_17594);
xor U17820 (N_17820,N_17670,N_17540);
nor U17821 (N_17821,N_17537,N_17472);
xor U17822 (N_17822,N_17565,N_17484);
or U17823 (N_17823,N_17515,N_17535);
nor U17824 (N_17824,N_17518,N_17659);
nor U17825 (N_17825,N_17480,N_17420);
nor U17826 (N_17826,N_17595,N_17602);
and U17827 (N_17827,N_17645,N_17580);
and U17828 (N_17828,N_17460,N_17462);
nand U17829 (N_17829,N_17587,N_17475);
nand U17830 (N_17830,N_17658,N_17488);
nor U17831 (N_17831,N_17575,N_17406);
and U17832 (N_17832,N_17631,N_17690);
and U17833 (N_17833,N_17498,N_17457);
or U17834 (N_17834,N_17611,N_17425);
and U17835 (N_17835,N_17491,N_17590);
and U17836 (N_17836,N_17432,N_17508);
and U17837 (N_17837,N_17500,N_17494);
nand U17838 (N_17838,N_17436,N_17652);
nand U17839 (N_17839,N_17553,N_17613);
and U17840 (N_17840,N_17589,N_17616);
nand U17841 (N_17841,N_17563,N_17532);
or U17842 (N_17842,N_17541,N_17547);
nor U17843 (N_17843,N_17490,N_17625);
nor U17844 (N_17844,N_17442,N_17615);
and U17845 (N_17845,N_17641,N_17576);
xor U17846 (N_17846,N_17465,N_17676);
nand U17847 (N_17847,N_17412,N_17507);
or U17848 (N_17848,N_17440,N_17510);
and U17849 (N_17849,N_17601,N_17441);
nor U17850 (N_17850,N_17567,N_17603);
xnor U17851 (N_17851,N_17627,N_17654);
and U17852 (N_17852,N_17667,N_17509);
nand U17853 (N_17853,N_17600,N_17624);
and U17854 (N_17854,N_17526,N_17449);
or U17855 (N_17855,N_17530,N_17496);
and U17856 (N_17856,N_17412,N_17628);
xnor U17857 (N_17857,N_17497,N_17404);
or U17858 (N_17858,N_17643,N_17636);
and U17859 (N_17859,N_17439,N_17421);
nand U17860 (N_17860,N_17496,N_17416);
nand U17861 (N_17861,N_17545,N_17593);
xnor U17862 (N_17862,N_17557,N_17670);
or U17863 (N_17863,N_17621,N_17685);
or U17864 (N_17864,N_17431,N_17488);
xor U17865 (N_17865,N_17436,N_17416);
nand U17866 (N_17866,N_17465,N_17505);
and U17867 (N_17867,N_17600,N_17425);
xor U17868 (N_17868,N_17480,N_17436);
nor U17869 (N_17869,N_17439,N_17423);
or U17870 (N_17870,N_17463,N_17550);
nand U17871 (N_17871,N_17698,N_17553);
nor U17872 (N_17872,N_17671,N_17501);
nand U17873 (N_17873,N_17443,N_17685);
nor U17874 (N_17874,N_17497,N_17456);
nor U17875 (N_17875,N_17502,N_17614);
nor U17876 (N_17876,N_17612,N_17478);
and U17877 (N_17877,N_17591,N_17573);
xnor U17878 (N_17878,N_17551,N_17553);
or U17879 (N_17879,N_17422,N_17537);
nand U17880 (N_17880,N_17577,N_17619);
xor U17881 (N_17881,N_17426,N_17502);
nor U17882 (N_17882,N_17493,N_17506);
nand U17883 (N_17883,N_17482,N_17490);
and U17884 (N_17884,N_17629,N_17523);
nor U17885 (N_17885,N_17542,N_17543);
or U17886 (N_17886,N_17491,N_17609);
nor U17887 (N_17887,N_17408,N_17422);
and U17888 (N_17888,N_17564,N_17462);
nor U17889 (N_17889,N_17490,N_17518);
and U17890 (N_17890,N_17582,N_17609);
nor U17891 (N_17891,N_17503,N_17652);
nor U17892 (N_17892,N_17510,N_17578);
or U17893 (N_17893,N_17462,N_17519);
nor U17894 (N_17894,N_17487,N_17603);
and U17895 (N_17895,N_17579,N_17459);
or U17896 (N_17896,N_17476,N_17581);
nand U17897 (N_17897,N_17606,N_17574);
and U17898 (N_17898,N_17463,N_17435);
nor U17899 (N_17899,N_17406,N_17589);
nor U17900 (N_17900,N_17504,N_17455);
nand U17901 (N_17901,N_17516,N_17603);
nor U17902 (N_17902,N_17415,N_17532);
nor U17903 (N_17903,N_17669,N_17649);
or U17904 (N_17904,N_17480,N_17516);
nor U17905 (N_17905,N_17511,N_17467);
nand U17906 (N_17906,N_17564,N_17667);
and U17907 (N_17907,N_17673,N_17422);
nand U17908 (N_17908,N_17672,N_17595);
and U17909 (N_17909,N_17697,N_17539);
nor U17910 (N_17910,N_17540,N_17459);
and U17911 (N_17911,N_17621,N_17637);
nor U17912 (N_17912,N_17564,N_17638);
nand U17913 (N_17913,N_17633,N_17682);
xnor U17914 (N_17914,N_17410,N_17579);
xor U17915 (N_17915,N_17490,N_17475);
or U17916 (N_17916,N_17575,N_17668);
xor U17917 (N_17917,N_17512,N_17500);
xnor U17918 (N_17918,N_17641,N_17671);
nor U17919 (N_17919,N_17518,N_17440);
nor U17920 (N_17920,N_17605,N_17571);
xnor U17921 (N_17921,N_17698,N_17604);
or U17922 (N_17922,N_17414,N_17688);
nand U17923 (N_17923,N_17606,N_17492);
nand U17924 (N_17924,N_17514,N_17485);
or U17925 (N_17925,N_17428,N_17500);
or U17926 (N_17926,N_17444,N_17649);
nor U17927 (N_17927,N_17499,N_17661);
xnor U17928 (N_17928,N_17414,N_17696);
nand U17929 (N_17929,N_17610,N_17553);
nor U17930 (N_17930,N_17475,N_17519);
xor U17931 (N_17931,N_17480,N_17444);
nand U17932 (N_17932,N_17673,N_17621);
xnor U17933 (N_17933,N_17444,N_17498);
and U17934 (N_17934,N_17594,N_17496);
xor U17935 (N_17935,N_17536,N_17612);
xor U17936 (N_17936,N_17435,N_17580);
nor U17937 (N_17937,N_17661,N_17470);
or U17938 (N_17938,N_17419,N_17560);
nand U17939 (N_17939,N_17549,N_17582);
nor U17940 (N_17940,N_17601,N_17453);
xor U17941 (N_17941,N_17644,N_17683);
and U17942 (N_17942,N_17618,N_17488);
nand U17943 (N_17943,N_17590,N_17525);
or U17944 (N_17944,N_17536,N_17448);
nor U17945 (N_17945,N_17669,N_17468);
nor U17946 (N_17946,N_17694,N_17515);
and U17947 (N_17947,N_17614,N_17601);
xor U17948 (N_17948,N_17572,N_17464);
nor U17949 (N_17949,N_17538,N_17560);
xor U17950 (N_17950,N_17457,N_17639);
xor U17951 (N_17951,N_17608,N_17497);
and U17952 (N_17952,N_17555,N_17442);
nor U17953 (N_17953,N_17526,N_17411);
and U17954 (N_17954,N_17695,N_17644);
xnor U17955 (N_17955,N_17421,N_17677);
xnor U17956 (N_17956,N_17407,N_17466);
nand U17957 (N_17957,N_17580,N_17460);
xnor U17958 (N_17958,N_17689,N_17592);
xnor U17959 (N_17959,N_17444,N_17534);
xnor U17960 (N_17960,N_17655,N_17428);
xnor U17961 (N_17961,N_17557,N_17515);
xor U17962 (N_17962,N_17410,N_17417);
and U17963 (N_17963,N_17432,N_17474);
or U17964 (N_17964,N_17551,N_17439);
nor U17965 (N_17965,N_17689,N_17436);
or U17966 (N_17966,N_17693,N_17496);
and U17967 (N_17967,N_17621,N_17421);
nor U17968 (N_17968,N_17600,N_17667);
nand U17969 (N_17969,N_17430,N_17686);
nor U17970 (N_17970,N_17656,N_17583);
nor U17971 (N_17971,N_17555,N_17583);
nor U17972 (N_17972,N_17478,N_17511);
nor U17973 (N_17973,N_17674,N_17602);
and U17974 (N_17974,N_17557,N_17626);
or U17975 (N_17975,N_17453,N_17553);
and U17976 (N_17976,N_17575,N_17444);
nor U17977 (N_17977,N_17630,N_17580);
nor U17978 (N_17978,N_17421,N_17605);
and U17979 (N_17979,N_17694,N_17574);
nor U17980 (N_17980,N_17433,N_17522);
nor U17981 (N_17981,N_17586,N_17475);
and U17982 (N_17982,N_17697,N_17448);
or U17983 (N_17983,N_17610,N_17539);
nor U17984 (N_17984,N_17495,N_17677);
or U17985 (N_17985,N_17569,N_17522);
or U17986 (N_17986,N_17540,N_17512);
and U17987 (N_17987,N_17468,N_17600);
nor U17988 (N_17988,N_17599,N_17640);
or U17989 (N_17989,N_17658,N_17557);
and U17990 (N_17990,N_17639,N_17572);
xor U17991 (N_17991,N_17434,N_17455);
or U17992 (N_17992,N_17527,N_17548);
nand U17993 (N_17993,N_17571,N_17460);
xnor U17994 (N_17994,N_17469,N_17558);
nor U17995 (N_17995,N_17596,N_17566);
nor U17996 (N_17996,N_17484,N_17434);
or U17997 (N_17997,N_17627,N_17563);
xnor U17998 (N_17998,N_17645,N_17522);
and U17999 (N_17999,N_17469,N_17568);
or U18000 (N_18000,N_17759,N_17845);
nand U18001 (N_18001,N_17826,N_17886);
nor U18002 (N_18002,N_17933,N_17930);
nor U18003 (N_18003,N_17770,N_17916);
or U18004 (N_18004,N_17832,N_17965);
nor U18005 (N_18005,N_17912,N_17911);
or U18006 (N_18006,N_17902,N_17821);
or U18007 (N_18007,N_17811,N_17846);
or U18008 (N_18008,N_17769,N_17949);
or U18009 (N_18009,N_17996,N_17828);
nor U18010 (N_18010,N_17987,N_17748);
xor U18011 (N_18011,N_17918,N_17941);
or U18012 (N_18012,N_17973,N_17755);
nand U18013 (N_18013,N_17749,N_17808);
or U18014 (N_18014,N_17839,N_17815);
xor U18015 (N_18015,N_17950,N_17931);
or U18016 (N_18016,N_17715,N_17750);
nand U18017 (N_18017,N_17724,N_17817);
nand U18018 (N_18018,N_17919,N_17752);
nand U18019 (N_18019,N_17897,N_17745);
or U18020 (N_18020,N_17823,N_17709);
nor U18021 (N_18021,N_17977,N_17969);
nor U18022 (N_18022,N_17865,N_17863);
xor U18023 (N_18023,N_17867,N_17746);
or U18024 (N_18024,N_17877,N_17940);
and U18025 (N_18025,N_17705,N_17922);
nand U18026 (N_18026,N_17850,N_17766);
xnor U18027 (N_18027,N_17801,N_17730);
nor U18028 (N_18028,N_17790,N_17925);
nand U18029 (N_18029,N_17860,N_17953);
xor U18030 (N_18030,N_17726,N_17926);
nor U18031 (N_18031,N_17921,N_17777);
nand U18032 (N_18032,N_17804,N_17783);
nor U18033 (N_18033,N_17714,N_17989);
nor U18034 (N_18034,N_17871,N_17982);
nand U18035 (N_18035,N_17961,N_17947);
nor U18036 (N_18036,N_17741,N_17731);
nand U18037 (N_18037,N_17791,N_17957);
or U18038 (N_18038,N_17798,N_17797);
and U18039 (N_18039,N_17906,N_17924);
nand U18040 (N_18040,N_17888,N_17814);
xnor U18041 (N_18041,N_17787,N_17717);
and U18042 (N_18042,N_17773,N_17822);
and U18043 (N_18043,N_17778,N_17838);
or U18044 (N_18044,N_17937,N_17908);
xor U18045 (N_18045,N_17994,N_17722);
or U18046 (N_18046,N_17895,N_17818);
xor U18047 (N_18047,N_17934,N_17824);
nor U18048 (N_18048,N_17964,N_17756);
or U18049 (N_18049,N_17927,N_17729);
xor U18050 (N_18050,N_17972,N_17768);
nor U18051 (N_18051,N_17904,N_17707);
nor U18052 (N_18052,N_17760,N_17803);
and U18053 (N_18053,N_17842,N_17998);
xor U18054 (N_18054,N_17767,N_17960);
nor U18055 (N_18055,N_17857,N_17988);
or U18056 (N_18056,N_17843,N_17829);
or U18057 (N_18057,N_17868,N_17742);
xnor U18058 (N_18058,N_17866,N_17898);
or U18059 (N_18059,N_17913,N_17862);
nand U18060 (N_18060,N_17851,N_17728);
nand U18061 (N_18061,N_17971,N_17956);
nand U18062 (N_18062,N_17983,N_17990);
and U18063 (N_18063,N_17735,N_17970);
and U18064 (N_18064,N_17847,N_17880);
nor U18065 (N_18065,N_17747,N_17786);
and U18066 (N_18066,N_17825,N_17951);
xnor U18067 (N_18067,N_17890,N_17819);
xnor U18068 (N_18068,N_17809,N_17720);
or U18069 (N_18069,N_17837,N_17946);
or U18070 (N_18070,N_17872,N_17995);
or U18071 (N_18071,N_17751,N_17810);
and U18072 (N_18072,N_17999,N_17993);
and U18073 (N_18073,N_17974,N_17792);
nor U18074 (N_18074,N_17870,N_17772);
xnor U18075 (N_18075,N_17844,N_17775);
nand U18076 (N_18076,N_17781,N_17892);
nand U18077 (N_18077,N_17859,N_17738);
xnor U18078 (N_18078,N_17861,N_17841);
nor U18079 (N_18079,N_17901,N_17997);
xor U18080 (N_18080,N_17725,N_17780);
or U18081 (N_18081,N_17952,N_17986);
nand U18082 (N_18082,N_17894,N_17736);
xnor U18083 (N_18083,N_17854,N_17807);
xnor U18084 (N_18084,N_17794,N_17849);
nor U18085 (N_18085,N_17882,N_17878);
or U18086 (N_18086,N_17727,N_17789);
and U18087 (N_18087,N_17938,N_17903);
xnor U18088 (N_18088,N_17876,N_17706);
and U18089 (N_18089,N_17856,N_17806);
and U18090 (N_18090,N_17785,N_17761);
and U18091 (N_18091,N_17985,N_17733);
nand U18092 (N_18092,N_17932,N_17732);
or U18093 (N_18093,N_17981,N_17836);
xnor U18094 (N_18094,N_17968,N_17833);
or U18095 (N_18095,N_17914,N_17884);
nor U18096 (N_18096,N_17753,N_17827);
xor U18097 (N_18097,N_17848,N_17928);
or U18098 (N_18098,N_17840,N_17885);
xor U18099 (N_18099,N_17874,N_17723);
nand U18100 (N_18100,N_17853,N_17936);
nor U18101 (N_18101,N_17887,N_17975);
xor U18102 (N_18102,N_17955,N_17943);
xor U18103 (N_18103,N_17805,N_17939);
and U18104 (N_18104,N_17812,N_17784);
xnor U18105 (N_18105,N_17879,N_17793);
nor U18106 (N_18106,N_17702,N_17744);
and U18107 (N_18107,N_17923,N_17883);
xor U18108 (N_18108,N_17800,N_17734);
nor U18109 (N_18109,N_17963,N_17976);
and U18110 (N_18110,N_17782,N_17762);
nor U18111 (N_18111,N_17992,N_17942);
xor U18112 (N_18112,N_17948,N_17855);
nand U18113 (N_18113,N_17891,N_17802);
nand U18114 (N_18114,N_17966,N_17959);
nor U18115 (N_18115,N_17905,N_17774);
or U18116 (N_18116,N_17710,N_17858);
nand U18117 (N_18117,N_17764,N_17889);
and U18118 (N_18118,N_17763,N_17917);
xor U18119 (N_18119,N_17743,N_17737);
and U18120 (N_18120,N_17967,N_17788);
or U18121 (N_18121,N_17719,N_17711);
xnor U18122 (N_18122,N_17765,N_17991);
or U18123 (N_18123,N_17831,N_17962);
or U18124 (N_18124,N_17896,N_17954);
or U18125 (N_18125,N_17779,N_17754);
nand U18126 (N_18126,N_17795,N_17757);
xnor U18127 (N_18127,N_17893,N_17958);
xnor U18128 (N_18128,N_17771,N_17716);
xnor U18129 (N_18129,N_17978,N_17873);
nor U18130 (N_18130,N_17799,N_17910);
nand U18131 (N_18131,N_17813,N_17835);
nor U18132 (N_18132,N_17718,N_17776);
or U18133 (N_18133,N_17920,N_17830);
and U18134 (N_18134,N_17915,N_17701);
or U18135 (N_18135,N_17909,N_17820);
or U18136 (N_18136,N_17796,N_17708);
nand U18137 (N_18137,N_17864,N_17700);
nor U18138 (N_18138,N_17984,N_17980);
xnor U18139 (N_18139,N_17944,N_17900);
xnor U18140 (N_18140,N_17899,N_17712);
nor U18141 (N_18141,N_17907,N_17852);
xnor U18142 (N_18142,N_17935,N_17713);
or U18143 (N_18143,N_17869,N_17721);
or U18144 (N_18144,N_17816,N_17704);
nand U18145 (N_18145,N_17881,N_17929);
and U18146 (N_18146,N_17834,N_17703);
xor U18147 (N_18147,N_17875,N_17758);
or U18148 (N_18148,N_17945,N_17740);
nor U18149 (N_18149,N_17739,N_17979);
nand U18150 (N_18150,N_17869,N_17824);
nand U18151 (N_18151,N_17792,N_17975);
nor U18152 (N_18152,N_17743,N_17968);
nor U18153 (N_18153,N_17990,N_17701);
nand U18154 (N_18154,N_17806,N_17849);
xor U18155 (N_18155,N_17753,N_17904);
or U18156 (N_18156,N_17820,N_17819);
nor U18157 (N_18157,N_17842,N_17919);
nand U18158 (N_18158,N_17884,N_17732);
or U18159 (N_18159,N_17731,N_17987);
and U18160 (N_18160,N_17929,N_17882);
nor U18161 (N_18161,N_17991,N_17718);
or U18162 (N_18162,N_17741,N_17831);
or U18163 (N_18163,N_17944,N_17941);
nand U18164 (N_18164,N_17778,N_17938);
nor U18165 (N_18165,N_17773,N_17849);
and U18166 (N_18166,N_17954,N_17823);
and U18167 (N_18167,N_17954,N_17824);
nor U18168 (N_18168,N_17804,N_17714);
or U18169 (N_18169,N_17916,N_17791);
xor U18170 (N_18170,N_17728,N_17711);
or U18171 (N_18171,N_17702,N_17796);
nand U18172 (N_18172,N_17948,N_17753);
xnor U18173 (N_18173,N_17987,N_17822);
nor U18174 (N_18174,N_17808,N_17842);
nand U18175 (N_18175,N_17776,N_17726);
or U18176 (N_18176,N_17917,N_17740);
and U18177 (N_18177,N_17920,N_17862);
nor U18178 (N_18178,N_17991,N_17938);
xor U18179 (N_18179,N_17739,N_17758);
and U18180 (N_18180,N_17945,N_17909);
nor U18181 (N_18181,N_17970,N_17960);
and U18182 (N_18182,N_17839,N_17924);
or U18183 (N_18183,N_17832,N_17807);
and U18184 (N_18184,N_17886,N_17890);
xor U18185 (N_18185,N_17783,N_17994);
xor U18186 (N_18186,N_17832,N_17814);
nand U18187 (N_18187,N_17994,N_17919);
xor U18188 (N_18188,N_17998,N_17978);
or U18189 (N_18189,N_17925,N_17828);
nand U18190 (N_18190,N_17758,N_17750);
xor U18191 (N_18191,N_17964,N_17837);
or U18192 (N_18192,N_17824,N_17970);
or U18193 (N_18193,N_17777,N_17780);
or U18194 (N_18194,N_17728,N_17782);
or U18195 (N_18195,N_17877,N_17701);
nand U18196 (N_18196,N_17946,N_17857);
xor U18197 (N_18197,N_17904,N_17775);
xnor U18198 (N_18198,N_17720,N_17723);
nor U18199 (N_18199,N_17944,N_17976);
xor U18200 (N_18200,N_17867,N_17717);
or U18201 (N_18201,N_17934,N_17985);
and U18202 (N_18202,N_17921,N_17865);
and U18203 (N_18203,N_17913,N_17780);
nand U18204 (N_18204,N_17990,N_17935);
or U18205 (N_18205,N_17955,N_17804);
xor U18206 (N_18206,N_17938,N_17964);
xnor U18207 (N_18207,N_17913,N_17872);
xor U18208 (N_18208,N_17860,N_17911);
nand U18209 (N_18209,N_17833,N_17701);
xnor U18210 (N_18210,N_17944,N_17918);
nor U18211 (N_18211,N_17755,N_17709);
nand U18212 (N_18212,N_17724,N_17728);
nor U18213 (N_18213,N_17857,N_17721);
xor U18214 (N_18214,N_17835,N_17773);
and U18215 (N_18215,N_17833,N_17759);
or U18216 (N_18216,N_17968,N_17938);
xnor U18217 (N_18217,N_17804,N_17950);
nor U18218 (N_18218,N_17719,N_17923);
and U18219 (N_18219,N_17943,N_17707);
nand U18220 (N_18220,N_17994,N_17876);
nor U18221 (N_18221,N_17940,N_17845);
nor U18222 (N_18222,N_17869,N_17850);
xor U18223 (N_18223,N_17815,N_17946);
and U18224 (N_18224,N_17800,N_17803);
nand U18225 (N_18225,N_17806,N_17752);
xnor U18226 (N_18226,N_17920,N_17797);
nor U18227 (N_18227,N_17801,N_17956);
nor U18228 (N_18228,N_17866,N_17779);
and U18229 (N_18229,N_17790,N_17971);
or U18230 (N_18230,N_17942,N_17703);
or U18231 (N_18231,N_17868,N_17895);
nor U18232 (N_18232,N_17990,N_17814);
and U18233 (N_18233,N_17830,N_17821);
xnor U18234 (N_18234,N_17777,N_17946);
nor U18235 (N_18235,N_17898,N_17721);
nand U18236 (N_18236,N_17872,N_17942);
or U18237 (N_18237,N_17857,N_17758);
xnor U18238 (N_18238,N_17944,N_17915);
nand U18239 (N_18239,N_17725,N_17729);
nand U18240 (N_18240,N_17919,N_17700);
or U18241 (N_18241,N_17745,N_17816);
or U18242 (N_18242,N_17889,N_17728);
nand U18243 (N_18243,N_17838,N_17979);
xnor U18244 (N_18244,N_17857,N_17831);
nand U18245 (N_18245,N_17866,N_17719);
nor U18246 (N_18246,N_17713,N_17743);
xor U18247 (N_18247,N_17895,N_17923);
or U18248 (N_18248,N_17902,N_17905);
nand U18249 (N_18249,N_17912,N_17813);
xnor U18250 (N_18250,N_17731,N_17883);
and U18251 (N_18251,N_17770,N_17868);
nor U18252 (N_18252,N_17903,N_17750);
xnor U18253 (N_18253,N_17834,N_17906);
and U18254 (N_18254,N_17984,N_17953);
nor U18255 (N_18255,N_17740,N_17729);
nand U18256 (N_18256,N_17837,N_17839);
or U18257 (N_18257,N_17754,N_17856);
xnor U18258 (N_18258,N_17916,N_17725);
and U18259 (N_18259,N_17944,N_17709);
nand U18260 (N_18260,N_17816,N_17773);
xnor U18261 (N_18261,N_17819,N_17907);
xor U18262 (N_18262,N_17958,N_17765);
nor U18263 (N_18263,N_17903,N_17769);
nor U18264 (N_18264,N_17804,N_17978);
and U18265 (N_18265,N_17860,N_17735);
xor U18266 (N_18266,N_17920,N_17984);
nand U18267 (N_18267,N_17724,N_17823);
and U18268 (N_18268,N_17753,N_17777);
nor U18269 (N_18269,N_17867,N_17702);
nor U18270 (N_18270,N_17961,N_17778);
nand U18271 (N_18271,N_17724,N_17953);
nand U18272 (N_18272,N_17940,N_17985);
xnor U18273 (N_18273,N_17978,N_17830);
or U18274 (N_18274,N_17751,N_17760);
and U18275 (N_18275,N_17725,N_17883);
xor U18276 (N_18276,N_17842,N_17755);
xor U18277 (N_18277,N_17979,N_17759);
nand U18278 (N_18278,N_17939,N_17933);
nor U18279 (N_18279,N_17743,N_17868);
nand U18280 (N_18280,N_17999,N_17714);
xnor U18281 (N_18281,N_17904,N_17722);
nor U18282 (N_18282,N_17779,N_17713);
or U18283 (N_18283,N_17744,N_17848);
and U18284 (N_18284,N_17769,N_17952);
and U18285 (N_18285,N_17959,N_17748);
or U18286 (N_18286,N_17958,N_17998);
nor U18287 (N_18287,N_17838,N_17815);
nor U18288 (N_18288,N_17944,N_17913);
and U18289 (N_18289,N_17787,N_17926);
nand U18290 (N_18290,N_17953,N_17706);
nand U18291 (N_18291,N_17951,N_17872);
or U18292 (N_18292,N_17734,N_17992);
nor U18293 (N_18293,N_17868,N_17753);
xnor U18294 (N_18294,N_17925,N_17936);
and U18295 (N_18295,N_17935,N_17718);
and U18296 (N_18296,N_17933,N_17805);
nor U18297 (N_18297,N_17723,N_17876);
xor U18298 (N_18298,N_17809,N_17894);
and U18299 (N_18299,N_17860,N_17881);
nand U18300 (N_18300,N_18296,N_18295);
or U18301 (N_18301,N_18096,N_18161);
nand U18302 (N_18302,N_18159,N_18240);
nor U18303 (N_18303,N_18139,N_18219);
or U18304 (N_18304,N_18110,N_18225);
or U18305 (N_18305,N_18049,N_18250);
or U18306 (N_18306,N_18007,N_18029);
or U18307 (N_18307,N_18232,N_18061);
and U18308 (N_18308,N_18059,N_18179);
nor U18309 (N_18309,N_18209,N_18235);
nor U18310 (N_18310,N_18208,N_18068);
nor U18311 (N_18311,N_18255,N_18268);
nand U18312 (N_18312,N_18281,N_18223);
or U18313 (N_18313,N_18163,N_18089);
xnor U18314 (N_18314,N_18211,N_18118);
or U18315 (N_18315,N_18273,N_18189);
xnor U18316 (N_18316,N_18270,N_18041);
or U18317 (N_18317,N_18093,N_18272);
xor U18318 (N_18318,N_18002,N_18030);
nor U18319 (N_18319,N_18063,N_18231);
xnor U18320 (N_18320,N_18199,N_18238);
nand U18321 (N_18321,N_18220,N_18138);
nand U18322 (N_18322,N_18203,N_18056);
nand U18323 (N_18323,N_18197,N_18187);
nand U18324 (N_18324,N_18018,N_18120);
xor U18325 (N_18325,N_18224,N_18131);
nor U18326 (N_18326,N_18191,N_18115);
and U18327 (N_18327,N_18137,N_18155);
and U18328 (N_18328,N_18025,N_18129);
or U18329 (N_18329,N_18124,N_18175);
nand U18330 (N_18330,N_18011,N_18294);
nor U18331 (N_18331,N_18153,N_18198);
nor U18332 (N_18332,N_18290,N_18264);
and U18333 (N_18333,N_18094,N_18257);
nand U18334 (N_18334,N_18230,N_18146);
xor U18335 (N_18335,N_18259,N_18228);
nand U18336 (N_18336,N_18109,N_18183);
and U18337 (N_18337,N_18044,N_18077);
and U18338 (N_18338,N_18251,N_18116);
nor U18339 (N_18339,N_18031,N_18222);
nor U18340 (N_18340,N_18072,N_18165);
nand U18341 (N_18341,N_18121,N_18286);
nor U18342 (N_18342,N_18239,N_18001);
nor U18343 (N_18343,N_18256,N_18026);
xor U18344 (N_18344,N_18032,N_18285);
and U18345 (N_18345,N_18288,N_18095);
nor U18346 (N_18346,N_18054,N_18143);
nand U18347 (N_18347,N_18057,N_18111);
xor U18348 (N_18348,N_18253,N_18252);
xnor U18349 (N_18349,N_18136,N_18112);
nor U18350 (N_18350,N_18174,N_18104);
nor U18351 (N_18351,N_18201,N_18132);
or U18352 (N_18352,N_18069,N_18040);
or U18353 (N_18353,N_18008,N_18035);
xor U18354 (N_18354,N_18188,N_18178);
or U18355 (N_18355,N_18123,N_18051);
nand U18356 (N_18356,N_18090,N_18243);
nand U18357 (N_18357,N_18108,N_18130);
or U18358 (N_18358,N_18176,N_18217);
xnor U18359 (N_18359,N_18145,N_18022);
xnor U18360 (N_18360,N_18084,N_18042);
xnor U18361 (N_18361,N_18043,N_18134);
nor U18362 (N_18362,N_18019,N_18245);
xnor U18363 (N_18363,N_18292,N_18128);
xnor U18364 (N_18364,N_18164,N_18046);
nand U18365 (N_18365,N_18287,N_18086);
nor U18366 (N_18366,N_18169,N_18218);
or U18367 (N_18367,N_18236,N_18140);
xnor U18368 (N_18368,N_18039,N_18027);
nor U18369 (N_18369,N_18216,N_18037);
or U18370 (N_18370,N_18293,N_18014);
nor U18371 (N_18371,N_18122,N_18065);
nand U18372 (N_18372,N_18071,N_18254);
or U18373 (N_18373,N_18221,N_18087);
nor U18374 (N_18374,N_18113,N_18213);
nand U18375 (N_18375,N_18023,N_18249);
nor U18376 (N_18376,N_18280,N_18004);
or U18377 (N_18377,N_18067,N_18227);
and U18378 (N_18378,N_18229,N_18241);
nand U18379 (N_18379,N_18156,N_18015);
xor U18380 (N_18380,N_18000,N_18263);
xnor U18381 (N_18381,N_18180,N_18073);
nand U18382 (N_18382,N_18291,N_18196);
nand U18383 (N_18383,N_18081,N_18016);
and U18384 (N_18384,N_18152,N_18012);
nand U18385 (N_18385,N_18091,N_18184);
nor U18386 (N_18386,N_18101,N_18075);
or U18387 (N_18387,N_18207,N_18050);
and U18388 (N_18388,N_18119,N_18234);
xnor U18389 (N_18389,N_18078,N_18149);
xnor U18390 (N_18390,N_18277,N_18171);
xnor U18391 (N_18391,N_18157,N_18092);
or U18392 (N_18392,N_18233,N_18076);
nor U18393 (N_18393,N_18062,N_18258);
xor U18394 (N_18394,N_18058,N_18009);
nand U18395 (N_18395,N_18060,N_18276);
nor U18396 (N_18396,N_18085,N_18013);
nand U18397 (N_18397,N_18248,N_18275);
xnor U18398 (N_18398,N_18168,N_18055);
nor U18399 (N_18399,N_18126,N_18142);
xor U18400 (N_18400,N_18202,N_18166);
nand U18401 (N_18401,N_18284,N_18262);
xor U18402 (N_18402,N_18210,N_18162);
xor U18403 (N_18403,N_18005,N_18079);
xnor U18404 (N_18404,N_18080,N_18271);
and U18405 (N_18405,N_18088,N_18246);
nand U18406 (N_18406,N_18215,N_18265);
nor U18407 (N_18407,N_18267,N_18100);
or U18408 (N_18408,N_18148,N_18117);
nand U18409 (N_18409,N_18151,N_18024);
or U18410 (N_18410,N_18150,N_18190);
and U18411 (N_18411,N_18177,N_18212);
xor U18412 (N_18412,N_18003,N_18127);
and U18413 (N_18413,N_18070,N_18298);
xor U18414 (N_18414,N_18028,N_18045);
or U18415 (N_18415,N_18102,N_18200);
and U18416 (N_18416,N_18182,N_18226);
and U18417 (N_18417,N_18097,N_18173);
nor U18418 (N_18418,N_18269,N_18106);
nor U18419 (N_18419,N_18237,N_18195);
and U18420 (N_18420,N_18020,N_18034);
or U18421 (N_18421,N_18204,N_18064);
and U18422 (N_18422,N_18141,N_18242);
xnor U18423 (N_18423,N_18021,N_18193);
and U18424 (N_18424,N_18099,N_18147);
nor U18425 (N_18425,N_18033,N_18036);
or U18426 (N_18426,N_18266,N_18299);
and U18427 (N_18427,N_18160,N_18074);
nor U18428 (N_18428,N_18214,N_18260);
or U18429 (N_18429,N_18066,N_18186);
nand U18430 (N_18430,N_18185,N_18052);
or U18431 (N_18431,N_18098,N_18107);
nand U18432 (N_18432,N_18283,N_18181);
and U18433 (N_18433,N_18278,N_18172);
and U18434 (N_18434,N_18133,N_18289);
nor U18435 (N_18435,N_18205,N_18158);
or U18436 (N_18436,N_18247,N_18194);
nor U18437 (N_18437,N_18274,N_18206);
nand U18438 (N_18438,N_18297,N_18154);
and U18439 (N_18439,N_18125,N_18135);
nor U18440 (N_18440,N_18006,N_18144);
or U18441 (N_18441,N_18170,N_18048);
or U18442 (N_18442,N_18279,N_18053);
and U18443 (N_18443,N_18083,N_18105);
nand U18444 (N_18444,N_18082,N_18282);
xnor U18445 (N_18445,N_18038,N_18192);
xnor U18446 (N_18446,N_18103,N_18261);
nor U18447 (N_18447,N_18114,N_18244);
nand U18448 (N_18448,N_18167,N_18017);
or U18449 (N_18449,N_18010,N_18047);
nand U18450 (N_18450,N_18238,N_18122);
nand U18451 (N_18451,N_18157,N_18071);
nand U18452 (N_18452,N_18266,N_18060);
or U18453 (N_18453,N_18052,N_18126);
nand U18454 (N_18454,N_18224,N_18014);
xor U18455 (N_18455,N_18256,N_18070);
or U18456 (N_18456,N_18280,N_18165);
nand U18457 (N_18457,N_18156,N_18293);
xor U18458 (N_18458,N_18227,N_18017);
and U18459 (N_18459,N_18142,N_18145);
xor U18460 (N_18460,N_18257,N_18078);
nand U18461 (N_18461,N_18202,N_18081);
and U18462 (N_18462,N_18154,N_18050);
nor U18463 (N_18463,N_18075,N_18095);
and U18464 (N_18464,N_18240,N_18000);
nor U18465 (N_18465,N_18154,N_18226);
nand U18466 (N_18466,N_18097,N_18284);
or U18467 (N_18467,N_18012,N_18019);
or U18468 (N_18468,N_18089,N_18234);
xnor U18469 (N_18469,N_18131,N_18281);
nand U18470 (N_18470,N_18287,N_18087);
nand U18471 (N_18471,N_18278,N_18050);
or U18472 (N_18472,N_18206,N_18227);
nand U18473 (N_18473,N_18067,N_18109);
and U18474 (N_18474,N_18258,N_18199);
or U18475 (N_18475,N_18032,N_18045);
xnor U18476 (N_18476,N_18254,N_18236);
or U18477 (N_18477,N_18215,N_18290);
xnor U18478 (N_18478,N_18014,N_18130);
and U18479 (N_18479,N_18243,N_18033);
xnor U18480 (N_18480,N_18149,N_18297);
xnor U18481 (N_18481,N_18255,N_18275);
or U18482 (N_18482,N_18136,N_18213);
or U18483 (N_18483,N_18009,N_18176);
and U18484 (N_18484,N_18000,N_18048);
and U18485 (N_18485,N_18175,N_18108);
nand U18486 (N_18486,N_18120,N_18268);
and U18487 (N_18487,N_18128,N_18240);
and U18488 (N_18488,N_18229,N_18219);
and U18489 (N_18489,N_18287,N_18050);
nor U18490 (N_18490,N_18108,N_18093);
and U18491 (N_18491,N_18251,N_18189);
nor U18492 (N_18492,N_18013,N_18029);
nand U18493 (N_18493,N_18054,N_18150);
nand U18494 (N_18494,N_18007,N_18166);
nand U18495 (N_18495,N_18207,N_18189);
nor U18496 (N_18496,N_18107,N_18217);
and U18497 (N_18497,N_18099,N_18158);
nand U18498 (N_18498,N_18077,N_18013);
xor U18499 (N_18499,N_18062,N_18031);
nor U18500 (N_18500,N_18245,N_18190);
nand U18501 (N_18501,N_18094,N_18147);
xor U18502 (N_18502,N_18279,N_18287);
nand U18503 (N_18503,N_18254,N_18105);
nand U18504 (N_18504,N_18139,N_18085);
nand U18505 (N_18505,N_18092,N_18179);
nor U18506 (N_18506,N_18103,N_18122);
xor U18507 (N_18507,N_18022,N_18057);
or U18508 (N_18508,N_18204,N_18109);
and U18509 (N_18509,N_18113,N_18299);
nor U18510 (N_18510,N_18085,N_18253);
or U18511 (N_18511,N_18015,N_18104);
or U18512 (N_18512,N_18002,N_18045);
and U18513 (N_18513,N_18174,N_18170);
nand U18514 (N_18514,N_18016,N_18293);
and U18515 (N_18515,N_18018,N_18037);
xor U18516 (N_18516,N_18114,N_18292);
xor U18517 (N_18517,N_18042,N_18166);
nor U18518 (N_18518,N_18009,N_18130);
and U18519 (N_18519,N_18292,N_18222);
or U18520 (N_18520,N_18294,N_18076);
xnor U18521 (N_18521,N_18245,N_18169);
xnor U18522 (N_18522,N_18016,N_18087);
nand U18523 (N_18523,N_18168,N_18129);
nand U18524 (N_18524,N_18061,N_18102);
or U18525 (N_18525,N_18089,N_18180);
or U18526 (N_18526,N_18180,N_18001);
or U18527 (N_18527,N_18165,N_18160);
or U18528 (N_18528,N_18194,N_18210);
nand U18529 (N_18529,N_18121,N_18071);
or U18530 (N_18530,N_18091,N_18205);
xnor U18531 (N_18531,N_18274,N_18250);
xnor U18532 (N_18532,N_18229,N_18242);
nor U18533 (N_18533,N_18263,N_18203);
nand U18534 (N_18534,N_18284,N_18033);
xor U18535 (N_18535,N_18232,N_18179);
nand U18536 (N_18536,N_18003,N_18265);
nand U18537 (N_18537,N_18020,N_18298);
nand U18538 (N_18538,N_18232,N_18131);
xnor U18539 (N_18539,N_18180,N_18152);
nor U18540 (N_18540,N_18267,N_18207);
nor U18541 (N_18541,N_18154,N_18219);
xnor U18542 (N_18542,N_18018,N_18072);
xor U18543 (N_18543,N_18236,N_18144);
or U18544 (N_18544,N_18131,N_18032);
nor U18545 (N_18545,N_18050,N_18274);
xnor U18546 (N_18546,N_18148,N_18247);
and U18547 (N_18547,N_18001,N_18245);
xor U18548 (N_18548,N_18130,N_18065);
nand U18549 (N_18549,N_18017,N_18244);
nor U18550 (N_18550,N_18159,N_18275);
xnor U18551 (N_18551,N_18253,N_18047);
and U18552 (N_18552,N_18094,N_18260);
and U18553 (N_18553,N_18087,N_18153);
nand U18554 (N_18554,N_18102,N_18035);
nand U18555 (N_18555,N_18052,N_18042);
and U18556 (N_18556,N_18186,N_18076);
nand U18557 (N_18557,N_18008,N_18048);
or U18558 (N_18558,N_18245,N_18003);
xnor U18559 (N_18559,N_18276,N_18120);
xor U18560 (N_18560,N_18175,N_18065);
nand U18561 (N_18561,N_18294,N_18265);
nand U18562 (N_18562,N_18087,N_18253);
xnor U18563 (N_18563,N_18297,N_18133);
and U18564 (N_18564,N_18018,N_18195);
or U18565 (N_18565,N_18141,N_18011);
nand U18566 (N_18566,N_18170,N_18032);
xor U18567 (N_18567,N_18264,N_18020);
or U18568 (N_18568,N_18215,N_18175);
xor U18569 (N_18569,N_18046,N_18032);
nand U18570 (N_18570,N_18051,N_18275);
xor U18571 (N_18571,N_18245,N_18073);
xor U18572 (N_18572,N_18120,N_18090);
or U18573 (N_18573,N_18104,N_18270);
nand U18574 (N_18574,N_18051,N_18212);
xnor U18575 (N_18575,N_18116,N_18128);
xnor U18576 (N_18576,N_18066,N_18058);
nor U18577 (N_18577,N_18180,N_18247);
nor U18578 (N_18578,N_18262,N_18083);
or U18579 (N_18579,N_18270,N_18105);
or U18580 (N_18580,N_18226,N_18080);
nand U18581 (N_18581,N_18045,N_18025);
nor U18582 (N_18582,N_18108,N_18137);
or U18583 (N_18583,N_18034,N_18246);
xnor U18584 (N_18584,N_18030,N_18259);
or U18585 (N_18585,N_18014,N_18123);
nand U18586 (N_18586,N_18269,N_18048);
or U18587 (N_18587,N_18265,N_18005);
or U18588 (N_18588,N_18011,N_18150);
and U18589 (N_18589,N_18124,N_18103);
and U18590 (N_18590,N_18147,N_18052);
nor U18591 (N_18591,N_18029,N_18173);
nor U18592 (N_18592,N_18123,N_18258);
and U18593 (N_18593,N_18189,N_18077);
xnor U18594 (N_18594,N_18173,N_18081);
nor U18595 (N_18595,N_18055,N_18052);
xnor U18596 (N_18596,N_18202,N_18180);
or U18597 (N_18597,N_18024,N_18052);
nand U18598 (N_18598,N_18112,N_18132);
nor U18599 (N_18599,N_18221,N_18282);
or U18600 (N_18600,N_18386,N_18573);
nand U18601 (N_18601,N_18378,N_18466);
nor U18602 (N_18602,N_18479,N_18308);
nor U18603 (N_18603,N_18531,N_18395);
xnor U18604 (N_18604,N_18348,N_18577);
and U18605 (N_18605,N_18400,N_18593);
or U18606 (N_18606,N_18484,N_18338);
or U18607 (N_18607,N_18473,N_18527);
xnor U18608 (N_18608,N_18568,N_18530);
nor U18609 (N_18609,N_18397,N_18320);
nor U18610 (N_18610,N_18476,N_18506);
nor U18611 (N_18611,N_18356,N_18342);
xor U18612 (N_18612,N_18553,N_18350);
or U18613 (N_18613,N_18425,N_18450);
xnor U18614 (N_18614,N_18319,N_18368);
nor U18615 (N_18615,N_18528,N_18539);
nand U18616 (N_18616,N_18599,N_18475);
nor U18617 (N_18617,N_18303,N_18410);
or U18618 (N_18618,N_18351,N_18534);
nor U18619 (N_18619,N_18501,N_18477);
or U18620 (N_18620,N_18487,N_18361);
xor U18621 (N_18621,N_18459,N_18417);
and U18622 (N_18622,N_18566,N_18495);
nor U18623 (N_18623,N_18586,N_18327);
nor U18624 (N_18624,N_18471,N_18366);
nor U18625 (N_18625,N_18565,N_18596);
nand U18626 (N_18626,N_18365,N_18381);
and U18627 (N_18627,N_18310,N_18579);
nor U18628 (N_18628,N_18541,N_18441);
nand U18629 (N_18629,N_18480,N_18333);
and U18630 (N_18630,N_18517,N_18353);
xnor U18631 (N_18631,N_18411,N_18325);
nor U18632 (N_18632,N_18391,N_18556);
nor U18633 (N_18633,N_18312,N_18420);
or U18634 (N_18634,N_18521,N_18555);
xnor U18635 (N_18635,N_18465,N_18551);
and U18636 (N_18636,N_18546,N_18409);
nand U18637 (N_18637,N_18537,N_18500);
nand U18638 (N_18638,N_18520,N_18529);
nor U18639 (N_18639,N_18499,N_18445);
and U18640 (N_18640,N_18560,N_18505);
or U18641 (N_18641,N_18550,N_18526);
xnor U18642 (N_18642,N_18340,N_18403);
nor U18643 (N_18643,N_18592,N_18416);
xnor U18644 (N_18644,N_18371,N_18414);
and U18645 (N_18645,N_18434,N_18494);
or U18646 (N_18646,N_18357,N_18374);
nand U18647 (N_18647,N_18571,N_18516);
xor U18648 (N_18648,N_18582,N_18455);
nand U18649 (N_18649,N_18511,N_18444);
nor U18650 (N_18650,N_18522,N_18405);
and U18651 (N_18651,N_18399,N_18418);
xor U18652 (N_18652,N_18502,N_18438);
and U18653 (N_18653,N_18488,N_18329);
nor U18654 (N_18654,N_18581,N_18321);
and U18655 (N_18655,N_18392,N_18382);
and U18656 (N_18656,N_18362,N_18557);
and U18657 (N_18657,N_18359,N_18481);
nand U18658 (N_18658,N_18326,N_18423);
xor U18659 (N_18659,N_18304,N_18360);
or U18660 (N_18660,N_18585,N_18363);
nor U18661 (N_18661,N_18478,N_18563);
nor U18662 (N_18662,N_18454,N_18462);
nand U18663 (N_18663,N_18460,N_18404);
nand U18664 (N_18664,N_18583,N_18548);
nor U18665 (N_18665,N_18393,N_18370);
nor U18666 (N_18666,N_18496,N_18503);
xor U18667 (N_18667,N_18514,N_18588);
xnor U18668 (N_18668,N_18492,N_18376);
nand U18669 (N_18669,N_18597,N_18334);
or U18670 (N_18670,N_18323,N_18430);
nor U18671 (N_18671,N_18464,N_18515);
xnor U18672 (N_18672,N_18598,N_18307);
xor U18673 (N_18673,N_18578,N_18358);
nand U18674 (N_18674,N_18564,N_18379);
nand U18675 (N_18675,N_18347,N_18383);
or U18676 (N_18676,N_18543,N_18524);
nand U18677 (N_18677,N_18375,N_18387);
xor U18678 (N_18678,N_18349,N_18318);
xor U18679 (N_18679,N_18401,N_18332);
or U18680 (N_18680,N_18335,N_18470);
or U18681 (N_18681,N_18498,N_18372);
and U18682 (N_18682,N_18497,N_18324);
nand U18683 (N_18683,N_18549,N_18384);
and U18684 (N_18684,N_18408,N_18587);
nor U18685 (N_18685,N_18493,N_18309);
xnor U18686 (N_18686,N_18355,N_18453);
nand U18687 (N_18687,N_18429,N_18552);
nand U18688 (N_18688,N_18576,N_18535);
nand U18689 (N_18689,N_18316,N_18431);
nand U18690 (N_18690,N_18390,N_18364);
nor U18691 (N_18691,N_18483,N_18584);
or U18692 (N_18692,N_18377,N_18433);
or U18693 (N_18693,N_18305,N_18437);
nand U18694 (N_18694,N_18426,N_18336);
and U18695 (N_18695,N_18538,N_18467);
nand U18696 (N_18696,N_18512,N_18562);
and U18697 (N_18697,N_18513,N_18570);
nand U18698 (N_18698,N_18407,N_18508);
and U18699 (N_18699,N_18533,N_18567);
nor U18700 (N_18700,N_18373,N_18532);
xnor U18701 (N_18701,N_18415,N_18339);
nand U18702 (N_18702,N_18354,N_18472);
or U18703 (N_18703,N_18561,N_18435);
xnor U18704 (N_18704,N_18545,N_18419);
nor U18705 (N_18705,N_18440,N_18485);
and U18706 (N_18706,N_18306,N_18490);
or U18707 (N_18707,N_18591,N_18428);
and U18708 (N_18708,N_18406,N_18486);
or U18709 (N_18709,N_18525,N_18595);
or U18710 (N_18710,N_18317,N_18542);
nor U18711 (N_18711,N_18482,N_18412);
nand U18712 (N_18712,N_18432,N_18452);
or U18713 (N_18713,N_18507,N_18396);
nand U18714 (N_18714,N_18367,N_18344);
nor U18715 (N_18715,N_18580,N_18523);
or U18716 (N_18716,N_18504,N_18590);
xor U18717 (N_18717,N_18446,N_18300);
nand U18718 (N_18718,N_18463,N_18343);
xor U18719 (N_18719,N_18448,N_18447);
xnor U18720 (N_18720,N_18443,N_18345);
nand U18721 (N_18721,N_18589,N_18544);
nand U18722 (N_18722,N_18540,N_18509);
or U18723 (N_18723,N_18594,N_18451);
and U18724 (N_18724,N_18489,N_18547);
nand U18725 (N_18725,N_18394,N_18559);
or U18726 (N_18726,N_18574,N_18341);
nand U18727 (N_18727,N_18313,N_18331);
xor U18728 (N_18728,N_18337,N_18461);
and U18729 (N_18729,N_18398,N_18468);
xor U18730 (N_18730,N_18424,N_18352);
or U18731 (N_18731,N_18572,N_18554);
xnor U18732 (N_18732,N_18301,N_18569);
nand U18733 (N_18733,N_18575,N_18474);
xnor U18734 (N_18734,N_18449,N_18380);
xnor U18735 (N_18735,N_18402,N_18458);
xnor U18736 (N_18736,N_18442,N_18314);
nand U18737 (N_18737,N_18436,N_18518);
or U18738 (N_18738,N_18536,N_18388);
nor U18739 (N_18739,N_18385,N_18469);
nand U18740 (N_18740,N_18302,N_18413);
nand U18741 (N_18741,N_18330,N_18519);
nor U18742 (N_18742,N_18510,N_18311);
nand U18743 (N_18743,N_18369,N_18328);
nand U18744 (N_18744,N_18346,N_18421);
xnor U18745 (N_18745,N_18491,N_18457);
nor U18746 (N_18746,N_18389,N_18558);
nand U18747 (N_18747,N_18439,N_18322);
and U18748 (N_18748,N_18427,N_18315);
nand U18749 (N_18749,N_18422,N_18456);
nand U18750 (N_18750,N_18415,N_18567);
and U18751 (N_18751,N_18588,N_18535);
and U18752 (N_18752,N_18387,N_18450);
nor U18753 (N_18753,N_18443,N_18469);
xnor U18754 (N_18754,N_18503,N_18529);
nor U18755 (N_18755,N_18598,N_18449);
xnor U18756 (N_18756,N_18414,N_18392);
nand U18757 (N_18757,N_18302,N_18547);
or U18758 (N_18758,N_18386,N_18570);
or U18759 (N_18759,N_18475,N_18458);
and U18760 (N_18760,N_18597,N_18421);
and U18761 (N_18761,N_18557,N_18444);
xor U18762 (N_18762,N_18485,N_18314);
nand U18763 (N_18763,N_18461,N_18391);
nor U18764 (N_18764,N_18505,N_18467);
xnor U18765 (N_18765,N_18584,N_18438);
nand U18766 (N_18766,N_18425,N_18490);
xor U18767 (N_18767,N_18557,N_18524);
xor U18768 (N_18768,N_18497,N_18457);
or U18769 (N_18769,N_18356,N_18574);
or U18770 (N_18770,N_18325,N_18581);
nand U18771 (N_18771,N_18404,N_18335);
nor U18772 (N_18772,N_18422,N_18334);
nor U18773 (N_18773,N_18462,N_18466);
xnor U18774 (N_18774,N_18333,N_18449);
or U18775 (N_18775,N_18319,N_18435);
nand U18776 (N_18776,N_18532,N_18394);
nand U18777 (N_18777,N_18540,N_18357);
xnor U18778 (N_18778,N_18404,N_18334);
nor U18779 (N_18779,N_18388,N_18512);
nand U18780 (N_18780,N_18408,N_18359);
or U18781 (N_18781,N_18439,N_18526);
xnor U18782 (N_18782,N_18439,N_18431);
and U18783 (N_18783,N_18564,N_18301);
nor U18784 (N_18784,N_18581,N_18542);
and U18785 (N_18785,N_18307,N_18327);
nor U18786 (N_18786,N_18360,N_18527);
xnor U18787 (N_18787,N_18470,N_18534);
or U18788 (N_18788,N_18475,N_18333);
nor U18789 (N_18789,N_18328,N_18429);
nand U18790 (N_18790,N_18439,N_18458);
and U18791 (N_18791,N_18485,N_18369);
nand U18792 (N_18792,N_18443,N_18478);
nor U18793 (N_18793,N_18393,N_18305);
nand U18794 (N_18794,N_18470,N_18591);
and U18795 (N_18795,N_18412,N_18302);
xor U18796 (N_18796,N_18405,N_18510);
or U18797 (N_18797,N_18511,N_18566);
and U18798 (N_18798,N_18475,N_18450);
nand U18799 (N_18799,N_18537,N_18491);
nand U18800 (N_18800,N_18546,N_18442);
xor U18801 (N_18801,N_18501,N_18442);
nand U18802 (N_18802,N_18449,N_18441);
and U18803 (N_18803,N_18303,N_18449);
xor U18804 (N_18804,N_18355,N_18482);
xnor U18805 (N_18805,N_18534,N_18449);
nand U18806 (N_18806,N_18515,N_18401);
and U18807 (N_18807,N_18446,N_18450);
xnor U18808 (N_18808,N_18419,N_18540);
nand U18809 (N_18809,N_18465,N_18594);
nor U18810 (N_18810,N_18482,N_18312);
xor U18811 (N_18811,N_18506,N_18438);
nand U18812 (N_18812,N_18308,N_18543);
xor U18813 (N_18813,N_18583,N_18549);
and U18814 (N_18814,N_18319,N_18318);
xnor U18815 (N_18815,N_18568,N_18598);
nor U18816 (N_18816,N_18367,N_18513);
or U18817 (N_18817,N_18390,N_18355);
xor U18818 (N_18818,N_18592,N_18368);
xor U18819 (N_18819,N_18302,N_18415);
and U18820 (N_18820,N_18396,N_18573);
xnor U18821 (N_18821,N_18471,N_18445);
nor U18822 (N_18822,N_18371,N_18339);
xnor U18823 (N_18823,N_18320,N_18332);
nand U18824 (N_18824,N_18444,N_18526);
and U18825 (N_18825,N_18535,N_18383);
and U18826 (N_18826,N_18569,N_18420);
nand U18827 (N_18827,N_18561,N_18316);
nand U18828 (N_18828,N_18313,N_18435);
and U18829 (N_18829,N_18460,N_18410);
and U18830 (N_18830,N_18406,N_18385);
or U18831 (N_18831,N_18454,N_18347);
and U18832 (N_18832,N_18504,N_18333);
xor U18833 (N_18833,N_18372,N_18464);
nand U18834 (N_18834,N_18581,N_18526);
nand U18835 (N_18835,N_18510,N_18550);
xor U18836 (N_18836,N_18387,N_18582);
nor U18837 (N_18837,N_18570,N_18331);
and U18838 (N_18838,N_18391,N_18312);
nand U18839 (N_18839,N_18336,N_18374);
or U18840 (N_18840,N_18384,N_18319);
nand U18841 (N_18841,N_18438,N_18433);
or U18842 (N_18842,N_18542,N_18427);
or U18843 (N_18843,N_18393,N_18365);
or U18844 (N_18844,N_18560,N_18366);
and U18845 (N_18845,N_18540,N_18379);
xor U18846 (N_18846,N_18522,N_18381);
nor U18847 (N_18847,N_18402,N_18307);
xnor U18848 (N_18848,N_18349,N_18432);
or U18849 (N_18849,N_18357,N_18513);
xnor U18850 (N_18850,N_18455,N_18599);
nand U18851 (N_18851,N_18577,N_18404);
xnor U18852 (N_18852,N_18420,N_18413);
and U18853 (N_18853,N_18500,N_18385);
or U18854 (N_18854,N_18416,N_18302);
xnor U18855 (N_18855,N_18597,N_18425);
nor U18856 (N_18856,N_18380,N_18320);
xor U18857 (N_18857,N_18364,N_18587);
and U18858 (N_18858,N_18361,N_18551);
nor U18859 (N_18859,N_18379,N_18480);
nand U18860 (N_18860,N_18418,N_18543);
and U18861 (N_18861,N_18389,N_18432);
nand U18862 (N_18862,N_18560,N_18354);
nor U18863 (N_18863,N_18561,N_18401);
or U18864 (N_18864,N_18305,N_18572);
nand U18865 (N_18865,N_18389,N_18355);
xnor U18866 (N_18866,N_18438,N_18371);
xnor U18867 (N_18867,N_18566,N_18363);
nor U18868 (N_18868,N_18365,N_18435);
nor U18869 (N_18869,N_18543,N_18591);
and U18870 (N_18870,N_18486,N_18322);
and U18871 (N_18871,N_18592,N_18462);
nor U18872 (N_18872,N_18448,N_18487);
nor U18873 (N_18873,N_18504,N_18365);
and U18874 (N_18874,N_18405,N_18545);
nor U18875 (N_18875,N_18416,N_18346);
nor U18876 (N_18876,N_18578,N_18548);
nand U18877 (N_18877,N_18440,N_18537);
and U18878 (N_18878,N_18430,N_18368);
nand U18879 (N_18879,N_18457,N_18429);
or U18880 (N_18880,N_18427,N_18571);
or U18881 (N_18881,N_18444,N_18401);
nand U18882 (N_18882,N_18396,N_18568);
nor U18883 (N_18883,N_18589,N_18440);
nor U18884 (N_18884,N_18357,N_18529);
xnor U18885 (N_18885,N_18343,N_18533);
or U18886 (N_18886,N_18404,N_18391);
nor U18887 (N_18887,N_18497,N_18395);
and U18888 (N_18888,N_18531,N_18495);
nor U18889 (N_18889,N_18415,N_18542);
xor U18890 (N_18890,N_18378,N_18482);
nor U18891 (N_18891,N_18534,N_18393);
and U18892 (N_18892,N_18521,N_18477);
and U18893 (N_18893,N_18365,N_18428);
and U18894 (N_18894,N_18410,N_18386);
or U18895 (N_18895,N_18449,N_18588);
and U18896 (N_18896,N_18384,N_18493);
nand U18897 (N_18897,N_18491,N_18353);
and U18898 (N_18898,N_18468,N_18456);
xor U18899 (N_18899,N_18374,N_18310);
or U18900 (N_18900,N_18838,N_18814);
xnor U18901 (N_18901,N_18613,N_18740);
xnor U18902 (N_18902,N_18705,N_18631);
nand U18903 (N_18903,N_18617,N_18707);
nand U18904 (N_18904,N_18717,N_18702);
xnor U18905 (N_18905,N_18723,N_18605);
and U18906 (N_18906,N_18662,N_18777);
nor U18907 (N_18907,N_18804,N_18810);
or U18908 (N_18908,N_18762,N_18763);
and U18909 (N_18909,N_18749,N_18610);
nand U18910 (N_18910,N_18863,N_18868);
or U18911 (N_18911,N_18837,N_18855);
and U18912 (N_18912,N_18722,N_18649);
and U18913 (N_18913,N_18888,N_18826);
nand U18914 (N_18914,N_18630,N_18690);
and U18915 (N_18915,N_18845,N_18758);
and U18916 (N_18916,N_18780,N_18643);
xor U18917 (N_18917,N_18852,N_18601);
xnor U18918 (N_18918,N_18694,N_18715);
xnor U18919 (N_18919,N_18825,N_18755);
nor U18920 (N_18920,N_18625,N_18672);
nand U18921 (N_18921,N_18618,N_18875);
nand U18922 (N_18922,N_18791,N_18693);
and U18923 (N_18923,N_18830,N_18734);
nor U18924 (N_18924,N_18853,N_18834);
or U18925 (N_18925,N_18687,N_18840);
and U18926 (N_18926,N_18829,N_18872);
xnor U18927 (N_18927,N_18882,N_18709);
nor U18928 (N_18928,N_18698,N_18787);
xnor U18929 (N_18929,N_18768,N_18896);
nor U18930 (N_18930,N_18761,N_18874);
or U18931 (N_18931,N_18674,N_18860);
nor U18932 (N_18932,N_18629,N_18750);
or U18933 (N_18933,N_18833,N_18799);
nand U18934 (N_18934,N_18894,N_18769);
xnor U18935 (N_18935,N_18710,N_18696);
nor U18936 (N_18936,N_18771,N_18623);
nand U18937 (N_18937,N_18607,N_18899);
and U18938 (N_18938,N_18773,N_18671);
nor U18939 (N_18939,N_18800,N_18858);
or U18940 (N_18940,N_18602,N_18893);
or U18941 (N_18941,N_18667,N_18898);
and U18942 (N_18942,N_18747,N_18752);
and U18943 (N_18943,N_18640,N_18684);
nor U18944 (N_18944,N_18759,N_18801);
nor U18945 (N_18945,N_18745,N_18859);
nor U18946 (N_18946,N_18879,N_18876);
nor U18947 (N_18947,N_18712,N_18721);
nand U18948 (N_18948,N_18827,N_18654);
or U18949 (N_18949,N_18781,N_18843);
or U18950 (N_18950,N_18685,N_18600);
nor U18951 (N_18951,N_18831,N_18611);
xor U18952 (N_18952,N_18638,N_18848);
nand U18953 (N_18953,N_18619,N_18603);
xor U18954 (N_18954,N_18641,N_18849);
xnor U18955 (N_18955,N_18784,N_18790);
nand U18956 (N_18956,N_18636,N_18708);
and U18957 (N_18957,N_18627,N_18776);
or U18958 (N_18958,N_18760,N_18862);
nand U18959 (N_18959,N_18884,N_18866);
xnor U18960 (N_18960,N_18892,N_18754);
and U18961 (N_18961,N_18701,N_18828);
nor U18962 (N_18962,N_18819,N_18659);
or U18963 (N_18963,N_18656,N_18714);
xnor U18964 (N_18964,N_18616,N_18737);
nand U18965 (N_18965,N_18748,N_18691);
or U18966 (N_18966,N_18802,N_18620);
xor U18967 (N_18967,N_18869,N_18806);
nand U18968 (N_18968,N_18835,N_18741);
xor U18969 (N_18969,N_18706,N_18670);
nor U18970 (N_18970,N_18779,N_18854);
nor U18971 (N_18971,N_18628,N_18883);
and U18972 (N_18972,N_18655,N_18661);
nand U18973 (N_18973,N_18724,N_18676);
nor U18974 (N_18974,N_18811,N_18728);
nand U18975 (N_18975,N_18744,N_18839);
nand U18976 (N_18976,N_18797,N_18842);
nor U18977 (N_18977,N_18870,N_18635);
xnor U18978 (N_18978,N_18632,N_18716);
or U18979 (N_18979,N_18891,N_18644);
xnor U18980 (N_18980,N_18673,N_18666);
xnor U18981 (N_18981,N_18703,N_18880);
or U18982 (N_18982,N_18699,N_18704);
nand U18983 (N_18983,N_18815,N_18772);
xor U18984 (N_18984,N_18633,N_18788);
and U18985 (N_18985,N_18615,N_18648);
nand U18986 (N_18986,N_18789,N_18794);
or U18987 (N_18987,N_18844,N_18682);
or U18988 (N_18988,N_18805,N_18756);
and U18989 (N_18989,N_18897,N_18887);
nor U18990 (N_18990,N_18680,N_18812);
nand U18991 (N_18991,N_18689,N_18792);
and U18992 (N_18992,N_18720,N_18889);
xnor U18993 (N_18993,N_18808,N_18622);
xor U18994 (N_18994,N_18871,N_18785);
nand U18995 (N_18995,N_18751,N_18621);
and U18996 (N_18996,N_18798,N_18816);
and U18997 (N_18997,N_18864,N_18668);
xnor U18998 (N_18998,N_18700,N_18626);
nand U18999 (N_18999,N_18757,N_18778);
and U19000 (N_19000,N_18824,N_18647);
xor U19001 (N_19001,N_18695,N_18770);
nor U19002 (N_19002,N_18735,N_18807);
and U19003 (N_19003,N_18786,N_18664);
xnor U19004 (N_19004,N_18823,N_18719);
nand U19005 (N_19005,N_18669,N_18642);
or U19006 (N_19006,N_18665,N_18637);
nand U19007 (N_19007,N_18767,N_18742);
nor U19008 (N_19008,N_18678,N_18609);
or U19009 (N_19009,N_18658,N_18624);
xor U19010 (N_19010,N_18832,N_18730);
xor U19011 (N_19011,N_18732,N_18729);
nand U19012 (N_19012,N_18736,N_18686);
nand U19013 (N_19013,N_18713,N_18604);
nor U19014 (N_19014,N_18820,N_18857);
and U19015 (N_19015,N_18877,N_18765);
and U19016 (N_19016,N_18681,N_18856);
xnor U19017 (N_19017,N_18821,N_18675);
nor U19018 (N_19018,N_18606,N_18692);
or U19019 (N_19019,N_18865,N_18688);
or U19020 (N_19020,N_18809,N_18614);
nor U19021 (N_19021,N_18775,N_18646);
xor U19022 (N_19022,N_18841,N_18612);
or U19023 (N_19023,N_18645,N_18651);
and U19024 (N_19024,N_18861,N_18774);
nor U19025 (N_19025,N_18727,N_18634);
nand U19026 (N_19026,N_18782,N_18697);
nand U19027 (N_19027,N_18679,N_18677);
nand U19028 (N_19028,N_18867,N_18847);
nor U19029 (N_19029,N_18895,N_18660);
xnor U19030 (N_19030,N_18881,N_18873);
nand U19031 (N_19031,N_18878,N_18711);
nand U19032 (N_19032,N_18738,N_18813);
nand U19033 (N_19033,N_18733,N_18793);
nand U19034 (N_19034,N_18836,N_18683);
and U19035 (N_19035,N_18851,N_18639);
nand U19036 (N_19036,N_18731,N_18885);
or U19037 (N_19037,N_18795,N_18818);
xor U19038 (N_19038,N_18796,N_18726);
nor U19039 (N_19039,N_18803,N_18608);
or U19040 (N_19040,N_18846,N_18725);
nor U19041 (N_19041,N_18718,N_18822);
nand U19042 (N_19042,N_18753,N_18739);
and U19043 (N_19043,N_18746,N_18766);
nand U19044 (N_19044,N_18850,N_18663);
nor U19045 (N_19045,N_18783,N_18890);
and U19046 (N_19046,N_18653,N_18886);
nand U19047 (N_19047,N_18650,N_18652);
or U19048 (N_19048,N_18743,N_18657);
nand U19049 (N_19049,N_18817,N_18764);
and U19050 (N_19050,N_18859,N_18763);
nand U19051 (N_19051,N_18848,N_18831);
and U19052 (N_19052,N_18649,N_18761);
and U19053 (N_19053,N_18689,N_18757);
and U19054 (N_19054,N_18621,N_18828);
nand U19055 (N_19055,N_18867,N_18749);
and U19056 (N_19056,N_18801,N_18601);
nand U19057 (N_19057,N_18638,N_18602);
and U19058 (N_19058,N_18686,N_18676);
or U19059 (N_19059,N_18792,N_18835);
nand U19060 (N_19060,N_18658,N_18604);
nand U19061 (N_19061,N_18614,N_18833);
and U19062 (N_19062,N_18844,N_18895);
nand U19063 (N_19063,N_18897,N_18708);
nor U19064 (N_19064,N_18786,N_18898);
nand U19065 (N_19065,N_18748,N_18605);
nor U19066 (N_19066,N_18676,N_18839);
nand U19067 (N_19067,N_18726,N_18884);
nor U19068 (N_19068,N_18678,N_18814);
and U19069 (N_19069,N_18633,N_18879);
nor U19070 (N_19070,N_18707,N_18794);
or U19071 (N_19071,N_18638,N_18623);
nand U19072 (N_19072,N_18683,N_18776);
nand U19073 (N_19073,N_18819,N_18690);
or U19074 (N_19074,N_18685,N_18721);
and U19075 (N_19075,N_18620,N_18656);
xnor U19076 (N_19076,N_18699,N_18604);
and U19077 (N_19077,N_18821,N_18878);
nand U19078 (N_19078,N_18667,N_18619);
xnor U19079 (N_19079,N_18732,N_18698);
or U19080 (N_19080,N_18761,N_18738);
and U19081 (N_19081,N_18622,N_18852);
or U19082 (N_19082,N_18600,N_18771);
and U19083 (N_19083,N_18781,N_18897);
nand U19084 (N_19084,N_18772,N_18812);
nor U19085 (N_19085,N_18767,N_18741);
nand U19086 (N_19086,N_18652,N_18625);
nand U19087 (N_19087,N_18809,N_18774);
nand U19088 (N_19088,N_18692,N_18869);
and U19089 (N_19089,N_18848,N_18660);
nand U19090 (N_19090,N_18729,N_18890);
nor U19091 (N_19091,N_18790,N_18698);
and U19092 (N_19092,N_18829,N_18727);
nor U19093 (N_19093,N_18808,N_18603);
or U19094 (N_19094,N_18867,N_18844);
nand U19095 (N_19095,N_18831,N_18637);
nand U19096 (N_19096,N_18714,N_18731);
nor U19097 (N_19097,N_18603,N_18741);
or U19098 (N_19098,N_18686,N_18734);
and U19099 (N_19099,N_18629,N_18838);
nand U19100 (N_19100,N_18830,N_18726);
or U19101 (N_19101,N_18876,N_18720);
or U19102 (N_19102,N_18811,N_18671);
and U19103 (N_19103,N_18621,N_18673);
nand U19104 (N_19104,N_18795,N_18723);
or U19105 (N_19105,N_18863,N_18740);
nor U19106 (N_19106,N_18892,N_18788);
or U19107 (N_19107,N_18865,N_18644);
or U19108 (N_19108,N_18746,N_18892);
or U19109 (N_19109,N_18617,N_18757);
xnor U19110 (N_19110,N_18826,N_18733);
or U19111 (N_19111,N_18791,N_18713);
nor U19112 (N_19112,N_18896,N_18644);
xor U19113 (N_19113,N_18817,N_18667);
xor U19114 (N_19114,N_18764,N_18890);
nand U19115 (N_19115,N_18641,N_18773);
nor U19116 (N_19116,N_18878,N_18814);
or U19117 (N_19117,N_18841,N_18798);
nor U19118 (N_19118,N_18723,N_18811);
or U19119 (N_19119,N_18788,N_18790);
xor U19120 (N_19120,N_18820,N_18754);
and U19121 (N_19121,N_18658,N_18640);
nor U19122 (N_19122,N_18677,N_18649);
nor U19123 (N_19123,N_18863,N_18803);
and U19124 (N_19124,N_18630,N_18767);
and U19125 (N_19125,N_18732,N_18875);
xor U19126 (N_19126,N_18659,N_18891);
nor U19127 (N_19127,N_18736,N_18833);
and U19128 (N_19128,N_18855,N_18815);
xnor U19129 (N_19129,N_18670,N_18680);
and U19130 (N_19130,N_18859,N_18621);
nor U19131 (N_19131,N_18723,N_18879);
xor U19132 (N_19132,N_18741,N_18807);
or U19133 (N_19133,N_18753,N_18698);
nor U19134 (N_19134,N_18718,N_18686);
or U19135 (N_19135,N_18779,N_18788);
xnor U19136 (N_19136,N_18892,N_18755);
and U19137 (N_19137,N_18888,N_18847);
xor U19138 (N_19138,N_18800,N_18848);
nor U19139 (N_19139,N_18782,N_18855);
xor U19140 (N_19140,N_18840,N_18877);
or U19141 (N_19141,N_18607,N_18853);
xnor U19142 (N_19142,N_18863,N_18708);
xnor U19143 (N_19143,N_18811,N_18749);
and U19144 (N_19144,N_18837,N_18821);
and U19145 (N_19145,N_18850,N_18698);
or U19146 (N_19146,N_18611,N_18769);
nand U19147 (N_19147,N_18790,N_18744);
nor U19148 (N_19148,N_18851,N_18813);
and U19149 (N_19149,N_18840,N_18885);
and U19150 (N_19150,N_18855,N_18820);
nor U19151 (N_19151,N_18793,N_18622);
or U19152 (N_19152,N_18835,N_18803);
and U19153 (N_19153,N_18895,N_18869);
or U19154 (N_19154,N_18775,N_18741);
xnor U19155 (N_19155,N_18814,N_18604);
nor U19156 (N_19156,N_18775,N_18721);
or U19157 (N_19157,N_18827,N_18814);
nand U19158 (N_19158,N_18779,N_18774);
xor U19159 (N_19159,N_18790,N_18604);
nand U19160 (N_19160,N_18669,N_18629);
nor U19161 (N_19161,N_18760,N_18810);
xor U19162 (N_19162,N_18760,N_18780);
nor U19163 (N_19163,N_18726,N_18814);
nand U19164 (N_19164,N_18673,N_18793);
or U19165 (N_19165,N_18664,N_18791);
nor U19166 (N_19166,N_18606,N_18612);
nor U19167 (N_19167,N_18871,N_18846);
xor U19168 (N_19168,N_18786,N_18725);
xnor U19169 (N_19169,N_18625,N_18822);
nor U19170 (N_19170,N_18815,N_18754);
nand U19171 (N_19171,N_18603,N_18881);
nand U19172 (N_19172,N_18658,N_18600);
nor U19173 (N_19173,N_18810,N_18776);
nand U19174 (N_19174,N_18857,N_18664);
or U19175 (N_19175,N_18763,N_18824);
or U19176 (N_19176,N_18782,N_18713);
or U19177 (N_19177,N_18734,N_18642);
and U19178 (N_19178,N_18872,N_18623);
and U19179 (N_19179,N_18720,N_18727);
and U19180 (N_19180,N_18755,N_18626);
nor U19181 (N_19181,N_18676,N_18682);
and U19182 (N_19182,N_18726,N_18860);
nand U19183 (N_19183,N_18746,N_18888);
and U19184 (N_19184,N_18659,N_18828);
and U19185 (N_19185,N_18805,N_18897);
or U19186 (N_19186,N_18841,N_18821);
or U19187 (N_19187,N_18677,N_18850);
nor U19188 (N_19188,N_18819,N_18893);
nand U19189 (N_19189,N_18714,N_18602);
or U19190 (N_19190,N_18601,N_18894);
or U19191 (N_19191,N_18612,N_18787);
and U19192 (N_19192,N_18618,N_18655);
or U19193 (N_19193,N_18660,N_18770);
and U19194 (N_19194,N_18836,N_18811);
or U19195 (N_19195,N_18626,N_18776);
xnor U19196 (N_19196,N_18726,N_18815);
xor U19197 (N_19197,N_18864,N_18710);
nor U19198 (N_19198,N_18646,N_18797);
nor U19199 (N_19199,N_18660,N_18705);
nor U19200 (N_19200,N_19196,N_19142);
and U19201 (N_19201,N_19011,N_19190);
nand U19202 (N_19202,N_18923,N_19038);
and U19203 (N_19203,N_19008,N_19080);
xnor U19204 (N_19204,N_18904,N_19000);
nand U19205 (N_19205,N_18921,N_18924);
xor U19206 (N_19206,N_18930,N_18978);
nor U19207 (N_19207,N_19108,N_18999);
xor U19208 (N_19208,N_19040,N_19115);
or U19209 (N_19209,N_18900,N_18986);
and U19210 (N_19210,N_19199,N_18960);
and U19211 (N_19211,N_19092,N_19068);
nor U19212 (N_19212,N_19197,N_19022);
nor U19213 (N_19213,N_19042,N_19153);
xor U19214 (N_19214,N_18984,N_19044);
or U19215 (N_19215,N_19017,N_19159);
nor U19216 (N_19216,N_19103,N_18997);
nor U19217 (N_19217,N_19039,N_18935);
nand U19218 (N_19218,N_18909,N_19111);
xor U19219 (N_19219,N_19057,N_18929);
nor U19220 (N_19220,N_19001,N_19123);
and U19221 (N_19221,N_18952,N_18977);
and U19222 (N_19222,N_19032,N_19051);
and U19223 (N_19223,N_19157,N_19192);
xor U19224 (N_19224,N_18969,N_19064);
nand U19225 (N_19225,N_19113,N_19061);
nand U19226 (N_19226,N_19110,N_18927);
and U19227 (N_19227,N_19094,N_19020);
xnor U19228 (N_19228,N_19066,N_19134);
or U19229 (N_19229,N_19125,N_18936);
xor U19230 (N_19230,N_19075,N_19100);
xnor U19231 (N_19231,N_18988,N_19118);
nor U19232 (N_19232,N_19127,N_18903);
nand U19233 (N_19233,N_19161,N_18948);
and U19234 (N_19234,N_19099,N_19165);
nand U19235 (N_19235,N_19049,N_19023);
or U19236 (N_19236,N_19045,N_18970);
xnor U19237 (N_19237,N_19174,N_18990);
nand U19238 (N_19238,N_19102,N_18908);
nor U19239 (N_19239,N_19137,N_19183);
or U19240 (N_19240,N_19116,N_19193);
and U19241 (N_19241,N_18902,N_19025);
nand U19242 (N_19242,N_18901,N_19139);
nor U19243 (N_19243,N_18995,N_19194);
and U19244 (N_19244,N_19097,N_19135);
nand U19245 (N_19245,N_18931,N_19091);
or U19246 (N_19246,N_18979,N_19005);
or U19247 (N_19247,N_18905,N_19069);
nand U19248 (N_19248,N_19033,N_19055);
or U19249 (N_19249,N_18932,N_18920);
xnor U19250 (N_19250,N_18994,N_18943);
and U19251 (N_19251,N_18926,N_18951);
nor U19252 (N_19252,N_19088,N_19004);
xnor U19253 (N_19253,N_19114,N_19019);
or U19254 (N_19254,N_19106,N_19084);
and U19255 (N_19255,N_19074,N_19098);
nor U19256 (N_19256,N_18992,N_19083);
nor U19257 (N_19257,N_19101,N_19180);
nand U19258 (N_19258,N_19043,N_19187);
and U19259 (N_19259,N_18906,N_18945);
nor U19260 (N_19260,N_19041,N_19067);
and U19261 (N_19261,N_19024,N_18940);
or U19262 (N_19262,N_19046,N_19141);
nor U19263 (N_19263,N_19050,N_18982);
and U19264 (N_19264,N_18962,N_19037);
nand U19265 (N_19265,N_19147,N_18938);
or U19266 (N_19266,N_19031,N_18987);
nor U19267 (N_19267,N_19130,N_19184);
xnor U19268 (N_19268,N_19076,N_19027);
xnor U19269 (N_19269,N_18983,N_19009);
nor U19270 (N_19270,N_19126,N_18950);
or U19271 (N_19271,N_18966,N_18974);
and U19272 (N_19272,N_19035,N_18918);
nor U19273 (N_19273,N_18973,N_19168);
or U19274 (N_19274,N_18947,N_19186);
or U19275 (N_19275,N_19185,N_19145);
xnor U19276 (N_19276,N_18912,N_19006);
nand U19277 (N_19277,N_18981,N_18961);
nor U19278 (N_19278,N_18937,N_19007);
nand U19279 (N_19279,N_19052,N_18907);
or U19280 (N_19280,N_19063,N_19117);
and U19281 (N_19281,N_19104,N_19029);
and U19282 (N_19282,N_19003,N_19162);
or U19283 (N_19283,N_19133,N_18910);
nand U19284 (N_19284,N_18913,N_19166);
and U19285 (N_19285,N_19138,N_19169);
nand U19286 (N_19286,N_19175,N_19121);
xor U19287 (N_19287,N_19177,N_19073);
nor U19288 (N_19288,N_19086,N_19191);
nand U19289 (N_19289,N_18959,N_19034);
or U19290 (N_19290,N_19176,N_19013);
or U19291 (N_19291,N_19060,N_19156);
and U19292 (N_19292,N_19058,N_19143);
nor U19293 (N_19293,N_19182,N_19078);
or U19294 (N_19294,N_19164,N_18946);
xor U19295 (N_19295,N_19077,N_19129);
nor U19296 (N_19296,N_19105,N_18916);
xnor U19297 (N_19297,N_18955,N_19171);
and U19298 (N_19298,N_18954,N_19195);
nand U19299 (N_19299,N_18925,N_18965);
or U19300 (N_19300,N_18917,N_19155);
or U19301 (N_19301,N_19163,N_18949);
nor U19302 (N_19302,N_19059,N_18915);
nand U19303 (N_19303,N_19128,N_19122);
and U19304 (N_19304,N_19015,N_18980);
or U19305 (N_19305,N_18958,N_19093);
or U19306 (N_19306,N_19018,N_19198);
nor U19307 (N_19307,N_19026,N_18934);
or U19308 (N_19308,N_18928,N_19150);
nand U19309 (N_19309,N_19132,N_19030);
or U19310 (N_19310,N_18963,N_19065);
xor U19311 (N_19311,N_19179,N_19012);
nor U19312 (N_19312,N_18971,N_19054);
nand U19313 (N_19313,N_18967,N_19124);
or U19314 (N_19314,N_19172,N_19167);
nand U19315 (N_19315,N_19095,N_19071);
and U19316 (N_19316,N_19072,N_19160);
or U19317 (N_19317,N_18939,N_19070);
and U19318 (N_19318,N_18968,N_18922);
nor U19319 (N_19319,N_19010,N_19120);
xor U19320 (N_19320,N_19090,N_19131);
nor U19321 (N_19321,N_19140,N_19158);
nand U19322 (N_19322,N_19014,N_19096);
or U19323 (N_19323,N_19107,N_19181);
xnor U19324 (N_19324,N_19136,N_19188);
xnor U19325 (N_19325,N_18998,N_18996);
or U19326 (N_19326,N_19119,N_19087);
xnor U19327 (N_19327,N_19154,N_18919);
or U19328 (N_19328,N_19112,N_18941);
and U19329 (N_19329,N_19144,N_19178);
or U19330 (N_19330,N_19189,N_19081);
xor U19331 (N_19331,N_19021,N_18944);
and U19332 (N_19332,N_18975,N_18914);
or U19333 (N_19333,N_19062,N_19085);
and U19334 (N_19334,N_19149,N_19089);
and U19335 (N_19335,N_18976,N_19053);
xor U19336 (N_19336,N_18989,N_19170);
nand U19337 (N_19337,N_18942,N_18911);
or U19338 (N_19338,N_19047,N_19002);
xnor U19339 (N_19339,N_18933,N_18991);
nor U19340 (N_19340,N_18956,N_19028);
nor U19341 (N_19341,N_19173,N_18972);
nor U19342 (N_19342,N_19148,N_19036);
xnor U19343 (N_19343,N_19151,N_19109);
nand U19344 (N_19344,N_19079,N_18953);
and U19345 (N_19345,N_19016,N_19082);
nor U19346 (N_19346,N_18964,N_18993);
nor U19347 (N_19347,N_19056,N_18985);
xor U19348 (N_19348,N_19146,N_19048);
and U19349 (N_19349,N_18957,N_19152);
nand U19350 (N_19350,N_18906,N_18939);
xor U19351 (N_19351,N_19127,N_19136);
and U19352 (N_19352,N_19104,N_19004);
and U19353 (N_19353,N_19003,N_19131);
xnor U19354 (N_19354,N_19078,N_19044);
and U19355 (N_19355,N_18971,N_19033);
or U19356 (N_19356,N_19006,N_18987);
nand U19357 (N_19357,N_18984,N_19043);
nor U19358 (N_19358,N_19026,N_19005);
nor U19359 (N_19359,N_19118,N_19072);
xor U19360 (N_19360,N_19031,N_18994);
nor U19361 (N_19361,N_19050,N_19189);
and U19362 (N_19362,N_19047,N_19092);
and U19363 (N_19363,N_18996,N_19007);
nand U19364 (N_19364,N_19073,N_19050);
nor U19365 (N_19365,N_18960,N_18958);
xnor U19366 (N_19366,N_19130,N_18957);
nand U19367 (N_19367,N_19108,N_19192);
nor U19368 (N_19368,N_19143,N_19163);
nor U19369 (N_19369,N_18937,N_18993);
nor U19370 (N_19370,N_19093,N_18954);
or U19371 (N_19371,N_19054,N_18946);
or U19372 (N_19372,N_19130,N_19150);
and U19373 (N_19373,N_19007,N_18951);
nand U19374 (N_19374,N_19046,N_18973);
nand U19375 (N_19375,N_18976,N_18940);
or U19376 (N_19376,N_19026,N_19051);
and U19377 (N_19377,N_19190,N_18999);
or U19378 (N_19378,N_19141,N_18929);
or U19379 (N_19379,N_18901,N_18931);
and U19380 (N_19380,N_18967,N_19191);
nor U19381 (N_19381,N_19155,N_19010);
xor U19382 (N_19382,N_19185,N_18921);
xnor U19383 (N_19383,N_19171,N_18986);
xnor U19384 (N_19384,N_18931,N_18953);
nand U19385 (N_19385,N_19102,N_19127);
and U19386 (N_19386,N_18921,N_19045);
nand U19387 (N_19387,N_18974,N_19169);
or U19388 (N_19388,N_19137,N_18975);
xnor U19389 (N_19389,N_18950,N_19038);
and U19390 (N_19390,N_19186,N_19167);
xnor U19391 (N_19391,N_19068,N_19186);
and U19392 (N_19392,N_18983,N_19114);
and U19393 (N_19393,N_19164,N_19167);
or U19394 (N_19394,N_19003,N_18996);
xnor U19395 (N_19395,N_19069,N_18957);
xnor U19396 (N_19396,N_19006,N_19023);
and U19397 (N_19397,N_19085,N_18907);
and U19398 (N_19398,N_19198,N_19058);
nand U19399 (N_19399,N_19148,N_19058);
and U19400 (N_19400,N_19185,N_18917);
nor U19401 (N_19401,N_19112,N_18975);
or U19402 (N_19402,N_18925,N_19141);
nand U19403 (N_19403,N_19110,N_18920);
and U19404 (N_19404,N_19173,N_18913);
and U19405 (N_19405,N_19122,N_18913);
xor U19406 (N_19406,N_19133,N_19159);
or U19407 (N_19407,N_19103,N_19183);
and U19408 (N_19408,N_19106,N_18922);
nor U19409 (N_19409,N_19087,N_19054);
xor U19410 (N_19410,N_18937,N_18939);
or U19411 (N_19411,N_19056,N_19171);
nand U19412 (N_19412,N_19151,N_18903);
or U19413 (N_19413,N_19157,N_18943);
nand U19414 (N_19414,N_19167,N_19108);
nand U19415 (N_19415,N_19174,N_19068);
and U19416 (N_19416,N_18955,N_19087);
and U19417 (N_19417,N_18931,N_18949);
nand U19418 (N_19418,N_19187,N_19117);
or U19419 (N_19419,N_19087,N_18919);
nor U19420 (N_19420,N_19004,N_19028);
xnor U19421 (N_19421,N_19049,N_19110);
nand U19422 (N_19422,N_18927,N_19061);
xnor U19423 (N_19423,N_19076,N_19192);
and U19424 (N_19424,N_19083,N_18931);
nand U19425 (N_19425,N_18993,N_18994);
xnor U19426 (N_19426,N_19167,N_18992);
and U19427 (N_19427,N_18968,N_19113);
xor U19428 (N_19428,N_19001,N_19045);
xor U19429 (N_19429,N_18905,N_19096);
nand U19430 (N_19430,N_18969,N_18940);
nor U19431 (N_19431,N_19057,N_19122);
or U19432 (N_19432,N_19097,N_18979);
nor U19433 (N_19433,N_18939,N_19021);
and U19434 (N_19434,N_19084,N_18961);
nand U19435 (N_19435,N_18916,N_18944);
xnor U19436 (N_19436,N_18926,N_19108);
nand U19437 (N_19437,N_19002,N_19056);
or U19438 (N_19438,N_19073,N_19137);
or U19439 (N_19439,N_19096,N_19086);
nand U19440 (N_19440,N_19072,N_19068);
xor U19441 (N_19441,N_19161,N_19076);
and U19442 (N_19442,N_19181,N_18901);
xnor U19443 (N_19443,N_19118,N_19070);
and U19444 (N_19444,N_19149,N_19190);
nand U19445 (N_19445,N_19052,N_19176);
nand U19446 (N_19446,N_18976,N_19021);
xnor U19447 (N_19447,N_18986,N_18966);
nand U19448 (N_19448,N_19069,N_19032);
xnor U19449 (N_19449,N_19094,N_19016);
xnor U19450 (N_19450,N_18933,N_19142);
xnor U19451 (N_19451,N_19135,N_18931);
and U19452 (N_19452,N_19143,N_19066);
nor U19453 (N_19453,N_19115,N_18956);
nand U19454 (N_19454,N_19103,N_19047);
or U19455 (N_19455,N_19120,N_19023);
and U19456 (N_19456,N_18906,N_19109);
nor U19457 (N_19457,N_19067,N_18928);
xnor U19458 (N_19458,N_19042,N_18973);
xnor U19459 (N_19459,N_19185,N_19020);
xnor U19460 (N_19460,N_19056,N_19165);
xnor U19461 (N_19461,N_19088,N_18936);
nor U19462 (N_19462,N_19064,N_19029);
nand U19463 (N_19463,N_18935,N_19048);
xor U19464 (N_19464,N_19043,N_18948);
or U19465 (N_19465,N_19028,N_18998);
xor U19466 (N_19466,N_18964,N_19065);
nand U19467 (N_19467,N_19013,N_19162);
and U19468 (N_19468,N_19107,N_19087);
nor U19469 (N_19469,N_19176,N_19102);
and U19470 (N_19470,N_18965,N_18988);
xor U19471 (N_19471,N_19185,N_19006);
and U19472 (N_19472,N_18952,N_19079);
and U19473 (N_19473,N_19095,N_19083);
nand U19474 (N_19474,N_19070,N_18970);
xnor U19475 (N_19475,N_18988,N_19089);
or U19476 (N_19476,N_19012,N_19062);
nand U19477 (N_19477,N_19184,N_19011);
nor U19478 (N_19478,N_19047,N_19191);
nand U19479 (N_19479,N_19033,N_18906);
xor U19480 (N_19480,N_18914,N_18957);
xor U19481 (N_19481,N_19085,N_19001);
or U19482 (N_19482,N_19025,N_19189);
and U19483 (N_19483,N_19145,N_19105);
nand U19484 (N_19484,N_19057,N_18946);
xnor U19485 (N_19485,N_18928,N_19037);
nand U19486 (N_19486,N_19082,N_18902);
and U19487 (N_19487,N_18998,N_18972);
and U19488 (N_19488,N_18984,N_19134);
nor U19489 (N_19489,N_19054,N_18907);
and U19490 (N_19490,N_19183,N_19021);
nand U19491 (N_19491,N_19162,N_18904);
xor U19492 (N_19492,N_19010,N_18964);
nor U19493 (N_19493,N_18955,N_18936);
nor U19494 (N_19494,N_19089,N_19114);
and U19495 (N_19495,N_19146,N_19057);
nand U19496 (N_19496,N_18982,N_18945);
xor U19497 (N_19497,N_18910,N_19032);
xnor U19498 (N_19498,N_19181,N_19028);
nor U19499 (N_19499,N_19069,N_19182);
nor U19500 (N_19500,N_19372,N_19499);
nand U19501 (N_19501,N_19436,N_19345);
nand U19502 (N_19502,N_19321,N_19323);
nor U19503 (N_19503,N_19248,N_19466);
and U19504 (N_19504,N_19231,N_19277);
nand U19505 (N_19505,N_19244,N_19452);
or U19506 (N_19506,N_19293,N_19402);
nor U19507 (N_19507,N_19457,N_19341);
nor U19508 (N_19508,N_19413,N_19219);
and U19509 (N_19509,N_19268,N_19291);
and U19510 (N_19510,N_19428,N_19458);
or U19511 (N_19511,N_19467,N_19403);
or U19512 (N_19512,N_19300,N_19253);
xnor U19513 (N_19513,N_19234,N_19303);
nand U19514 (N_19514,N_19265,N_19232);
and U19515 (N_19515,N_19239,N_19358);
nand U19516 (N_19516,N_19274,N_19371);
and U19517 (N_19517,N_19410,N_19242);
xor U19518 (N_19518,N_19495,N_19355);
xor U19519 (N_19519,N_19204,N_19250);
or U19520 (N_19520,N_19456,N_19370);
xor U19521 (N_19521,N_19289,N_19388);
nand U19522 (N_19522,N_19263,N_19241);
nor U19523 (N_19523,N_19415,N_19337);
or U19524 (N_19524,N_19475,N_19399);
nor U19525 (N_19525,N_19258,N_19423);
nand U19526 (N_19526,N_19366,N_19471);
and U19527 (N_19527,N_19276,N_19243);
xor U19528 (N_19528,N_19492,N_19412);
xnor U19529 (N_19529,N_19275,N_19405);
nor U19530 (N_19530,N_19297,N_19351);
nor U19531 (N_19531,N_19352,N_19472);
xor U19532 (N_19532,N_19357,N_19331);
and U19533 (N_19533,N_19335,N_19319);
nand U19534 (N_19534,N_19272,N_19392);
xor U19535 (N_19535,N_19236,N_19356);
or U19536 (N_19536,N_19486,N_19223);
or U19537 (N_19537,N_19271,N_19266);
xnor U19538 (N_19538,N_19498,N_19430);
xor U19539 (N_19539,N_19483,N_19365);
xnor U19540 (N_19540,N_19391,N_19210);
nand U19541 (N_19541,N_19380,N_19340);
nor U19542 (N_19542,N_19346,N_19469);
xnor U19543 (N_19543,N_19262,N_19247);
nor U19544 (N_19544,N_19240,N_19447);
or U19545 (N_19545,N_19317,N_19453);
xor U19546 (N_19546,N_19427,N_19269);
and U19547 (N_19547,N_19259,N_19406);
xnor U19548 (N_19548,N_19254,N_19398);
xnor U19549 (N_19549,N_19316,N_19480);
or U19550 (N_19550,N_19360,N_19379);
nand U19551 (N_19551,N_19260,N_19455);
and U19552 (N_19552,N_19494,N_19414);
and U19553 (N_19553,N_19228,N_19216);
nor U19554 (N_19554,N_19464,N_19279);
xor U19555 (N_19555,N_19327,N_19238);
or U19556 (N_19556,N_19387,N_19382);
and U19557 (N_19557,N_19426,N_19446);
xnor U19558 (N_19558,N_19218,N_19349);
xor U19559 (N_19559,N_19220,N_19377);
nand U19560 (N_19560,N_19417,N_19201);
nor U19561 (N_19561,N_19282,N_19255);
or U19562 (N_19562,N_19318,N_19288);
nor U19563 (N_19563,N_19299,N_19313);
nand U19564 (N_19564,N_19373,N_19336);
nor U19565 (N_19565,N_19226,N_19344);
xor U19566 (N_19566,N_19257,N_19381);
xnor U19567 (N_19567,N_19322,N_19347);
xor U19568 (N_19568,N_19407,N_19361);
nand U19569 (N_19569,N_19315,N_19296);
xor U19570 (N_19570,N_19330,N_19487);
nand U19571 (N_19571,N_19229,N_19252);
xnor U19572 (N_19572,N_19261,N_19310);
nand U19573 (N_19573,N_19353,N_19444);
and U19574 (N_19574,N_19302,N_19488);
or U19575 (N_19575,N_19249,N_19207);
xnor U19576 (N_19576,N_19376,N_19217);
or U19577 (N_19577,N_19235,N_19450);
and U19578 (N_19578,N_19443,N_19211);
xor U19579 (N_19579,N_19431,N_19369);
xnor U19580 (N_19580,N_19230,N_19460);
nor U19581 (N_19581,N_19437,N_19213);
nor U19582 (N_19582,N_19292,N_19237);
xor U19583 (N_19583,N_19485,N_19203);
or U19584 (N_19584,N_19484,N_19440);
xnor U19585 (N_19585,N_19280,N_19301);
nor U19586 (N_19586,N_19393,N_19468);
nor U19587 (N_19587,N_19332,N_19489);
or U19588 (N_19588,N_19283,N_19215);
nor U19589 (N_19589,N_19429,N_19294);
xnor U19590 (N_19590,N_19422,N_19325);
or U19591 (N_19591,N_19342,N_19481);
or U19592 (N_19592,N_19390,N_19295);
nor U19593 (N_19593,N_19290,N_19224);
nor U19594 (N_19594,N_19368,N_19432);
nor U19595 (N_19595,N_19497,N_19383);
or U19596 (N_19596,N_19202,N_19397);
or U19597 (N_19597,N_19386,N_19479);
or U19598 (N_19598,N_19478,N_19298);
xor U19599 (N_19599,N_19212,N_19438);
nor U19600 (N_19600,N_19419,N_19307);
nand U19601 (N_19601,N_19490,N_19278);
and U19602 (N_19602,N_19264,N_19451);
nor U19603 (N_19603,N_19306,N_19328);
nor U19604 (N_19604,N_19362,N_19320);
xor U19605 (N_19605,N_19374,N_19401);
nand U19606 (N_19606,N_19214,N_19395);
nand U19607 (N_19607,N_19359,N_19225);
or U19608 (N_19608,N_19420,N_19364);
nand U19609 (N_19609,N_19245,N_19461);
or U19610 (N_19610,N_19465,N_19334);
nor U19611 (N_19611,N_19348,N_19363);
or U19612 (N_19612,N_19389,N_19433);
nor U19613 (N_19613,N_19286,N_19445);
and U19614 (N_19614,N_19408,N_19384);
xnor U19615 (N_19615,N_19256,N_19281);
nand U19616 (N_19616,N_19425,N_19270);
or U19617 (N_19617,N_19350,N_19404);
or U19618 (N_19618,N_19434,N_19339);
xor U19619 (N_19619,N_19308,N_19208);
or U19620 (N_19620,N_19209,N_19354);
nor U19621 (N_19621,N_19396,N_19329);
and U19622 (N_19622,N_19375,N_19439);
and U19623 (N_19623,N_19462,N_19273);
nand U19624 (N_19624,N_19206,N_19400);
xor U19625 (N_19625,N_19285,N_19476);
or U19626 (N_19626,N_19251,N_19304);
xor U19627 (N_19627,N_19200,N_19287);
nor U19628 (N_19628,N_19416,N_19378);
and U19629 (N_19629,N_19421,N_19333);
nand U19630 (N_19630,N_19314,N_19482);
or U19631 (N_19631,N_19435,N_19409);
and U19632 (N_19632,N_19470,N_19454);
xor U19633 (N_19633,N_19338,N_19459);
nor U19634 (N_19634,N_19418,N_19312);
or U19635 (N_19635,N_19343,N_19474);
nor U19636 (N_19636,N_19385,N_19367);
nand U19637 (N_19637,N_19491,N_19493);
nand U19638 (N_19638,N_19411,N_19233);
nand U19639 (N_19639,N_19227,N_19473);
or U19640 (N_19640,N_19477,N_19442);
and U19641 (N_19641,N_19267,N_19448);
xnor U19642 (N_19642,N_19311,N_19424);
or U19643 (N_19643,N_19463,N_19326);
xnor U19644 (N_19644,N_19222,N_19246);
or U19645 (N_19645,N_19324,N_19205);
and U19646 (N_19646,N_19305,N_19394);
and U19647 (N_19647,N_19449,N_19441);
and U19648 (N_19648,N_19221,N_19284);
xnor U19649 (N_19649,N_19309,N_19496);
xor U19650 (N_19650,N_19396,N_19376);
and U19651 (N_19651,N_19345,N_19224);
and U19652 (N_19652,N_19387,N_19443);
or U19653 (N_19653,N_19209,N_19385);
or U19654 (N_19654,N_19497,N_19396);
or U19655 (N_19655,N_19403,N_19229);
and U19656 (N_19656,N_19227,N_19424);
nand U19657 (N_19657,N_19389,N_19282);
nand U19658 (N_19658,N_19248,N_19278);
or U19659 (N_19659,N_19215,N_19450);
xnor U19660 (N_19660,N_19232,N_19326);
nand U19661 (N_19661,N_19225,N_19258);
nor U19662 (N_19662,N_19254,N_19331);
xor U19663 (N_19663,N_19374,N_19209);
and U19664 (N_19664,N_19206,N_19482);
or U19665 (N_19665,N_19312,N_19476);
nand U19666 (N_19666,N_19249,N_19416);
xnor U19667 (N_19667,N_19385,N_19348);
and U19668 (N_19668,N_19319,N_19395);
xnor U19669 (N_19669,N_19448,N_19383);
or U19670 (N_19670,N_19414,N_19391);
nor U19671 (N_19671,N_19243,N_19286);
and U19672 (N_19672,N_19350,N_19491);
xnor U19673 (N_19673,N_19229,N_19492);
nor U19674 (N_19674,N_19267,N_19347);
xnor U19675 (N_19675,N_19455,N_19424);
nor U19676 (N_19676,N_19429,N_19200);
or U19677 (N_19677,N_19245,N_19346);
and U19678 (N_19678,N_19384,N_19498);
and U19679 (N_19679,N_19463,N_19433);
or U19680 (N_19680,N_19348,N_19334);
xnor U19681 (N_19681,N_19356,N_19200);
and U19682 (N_19682,N_19349,N_19229);
or U19683 (N_19683,N_19409,N_19322);
xor U19684 (N_19684,N_19328,N_19480);
or U19685 (N_19685,N_19441,N_19207);
or U19686 (N_19686,N_19413,N_19221);
nand U19687 (N_19687,N_19245,N_19384);
xor U19688 (N_19688,N_19254,N_19351);
or U19689 (N_19689,N_19464,N_19477);
nor U19690 (N_19690,N_19463,N_19452);
xor U19691 (N_19691,N_19207,N_19293);
xnor U19692 (N_19692,N_19384,N_19219);
nor U19693 (N_19693,N_19257,N_19316);
nor U19694 (N_19694,N_19458,N_19208);
and U19695 (N_19695,N_19424,N_19325);
xor U19696 (N_19696,N_19454,N_19304);
nor U19697 (N_19697,N_19297,N_19204);
nor U19698 (N_19698,N_19217,N_19280);
or U19699 (N_19699,N_19339,N_19480);
nand U19700 (N_19700,N_19315,N_19233);
nand U19701 (N_19701,N_19477,N_19380);
xnor U19702 (N_19702,N_19316,N_19454);
or U19703 (N_19703,N_19280,N_19287);
nor U19704 (N_19704,N_19315,N_19328);
nor U19705 (N_19705,N_19386,N_19257);
nor U19706 (N_19706,N_19434,N_19479);
and U19707 (N_19707,N_19445,N_19308);
and U19708 (N_19708,N_19258,N_19382);
or U19709 (N_19709,N_19355,N_19456);
or U19710 (N_19710,N_19389,N_19437);
and U19711 (N_19711,N_19257,N_19213);
nor U19712 (N_19712,N_19445,N_19407);
and U19713 (N_19713,N_19485,N_19307);
or U19714 (N_19714,N_19264,N_19305);
or U19715 (N_19715,N_19285,N_19499);
nand U19716 (N_19716,N_19429,N_19479);
xor U19717 (N_19717,N_19424,N_19310);
xnor U19718 (N_19718,N_19264,N_19335);
nand U19719 (N_19719,N_19201,N_19299);
and U19720 (N_19720,N_19366,N_19447);
or U19721 (N_19721,N_19405,N_19443);
xor U19722 (N_19722,N_19212,N_19273);
or U19723 (N_19723,N_19377,N_19331);
and U19724 (N_19724,N_19466,N_19294);
nor U19725 (N_19725,N_19333,N_19452);
and U19726 (N_19726,N_19232,N_19249);
xor U19727 (N_19727,N_19332,N_19295);
nor U19728 (N_19728,N_19327,N_19219);
or U19729 (N_19729,N_19343,N_19323);
nor U19730 (N_19730,N_19271,N_19236);
or U19731 (N_19731,N_19469,N_19233);
nor U19732 (N_19732,N_19200,N_19286);
nand U19733 (N_19733,N_19474,N_19476);
xnor U19734 (N_19734,N_19275,N_19290);
nand U19735 (N_19735,N_19233,N_19322);
nand U19736 (N_19736,N_19403,N_19243);
nand U19737 (N_19737,N_19285,N_19400);
or U19738 (N_19738,N_19343,N_19391);
nor U19739 (N_19739,N_19476,N_19302);
nand U19740 (N_19740,N_19398,N_19343);
nand U19741 (N_19741,N_19399,N_19272);
nor U19742 (N_19742,N_19227,N_19323);
nor U19743 (N_19743,N_19427,N_19487);
or U19744 (N_19744,N_19388,N_19433);
nand U19745 (N_19745,N_19271,N_19333);
xnor U19746 (N_19746,N_19451,N_19274);
xor U19747 (N_19747,N_19380,N_19496);
nor U19748 (N_19748,N_19376,N_19210);
nor U19749 (N_19749,N_19289,N_19411);
xnor U19750 (N_19750,N_19495,N_19466);
nand U19751 (N_19751,N_19243,N_19419);
xnor U19752 (N_19752,N_19474,N_19302);
and U19753 (N_19753,N_19355,N_19257);
nand U19754 (N_19754,N_19349,N_19406);
xnor U19755 (N_19755,N_19376,N_19466);
nand U19756 (N_19756,N_19312,N_19336);
xor U19757 (N_19757,N_19201,N_19414);
or U19758 (N_19758,N_19319,N_19445);
nor U19759 (N_19759,N_19483,N_19403);
and U19760 (N_19760,N_19297,N_19370);
and U19761 (N_19761,N_19443,N_19288);
or U19762 (N_19762,N_19469,N_19396);
or U19763 (N_19763,N_19458,N_19299);
and U19764 (N_19764,N_19204,N_19277);
nor U19765 (N_19765,N_19221,N_19315);
and U19766 (N_19766,N_19215,N_19471);
or U19767 (N_19767,N_19470,N_19363);
xnor U19768 (N_19768,N_19382,N_19211);
and U19769 (N_19769,N_19205,N_19371);
or U19770 (N_19770,N_19281,N_19398);
nand U19771 (N_19771,N_19400,N_19460);
or U19772 (N_19772,N_19424,N_19316);
or U19773 (N_19773,N_19317,N_19266);
nor U19774 (N_19774,N_19371,N_19321);
or U19775 (N_19775,N_19406,N_19378);
and U19776 (N_19776,N_19449,N_19387);
xor U19777 (N_19777,N_19404,N_19390);
xor U19778 (N_19778,N_19280,N_19481);
xor U19779 (N_19779,N_19384,N_19222);
and U19780 (N_19780,N_19487,N_19470);
and U19781 (N_19781,N_19295,N_19396);
nand U19782 (N_19782,N_19334,N_19323);
and U19783 (N_19783,N_19411,N_19319);
nand U19784 (N_19784,N_19282,N_19310);
or U19785 (N_19785,N_19389,N_19355);
nand U19786 (N_19786,N_19404,N_19274);
nand U19787 (N_19787,N_19339,N_19383);
nor U19788 (N_19788,N_19419,N_19388);
or U19789 (N_19789,N_19219,N_19392);
nand U19790 (N_19790,N_19341,N_19368);
or U19791 (N_19791,N_19466,N_19448);
or U19792 (N_19792,N_19316,N_19248);
and U19793 (N_19793,N_19256,N_19427);
and U19794 (N_19794,N_19204,N_19256);
or U19795 (N_19795,N_19499,N_19270);
nand U19796 (N_19796,N_19458,N_19230);
or U19797 (N_19797,N_19345,N_19256);
xnor U19798 (N_19798,N_19446,N_19332);
and U19799 (N_19799,N_19411,N_19210);
nand U19800 (N_19800,N_19553,N_19547);
and U19801 (N_19801,N_19719,N_19577);
and U19802 (N_19802,N_19520,N_19578);
and U19803 (N_19803,N_19586,N_19512);
xor U19804 (N_19804,N_19660,N_19678);
xor U19805 (N_19805,N_19721,N_19510);
or U19806 (N_19806,N_19528,N_19761);
nand U19807 (N_19807,N_19789,N_19613);
and U19808 (N_19808,N_19693,N_19692);
nand U19809 (N_19809,N_19662,N_19772);
xor U19810 (N_19810,N_19738,N_19582);
nand U19811 (N_19811,N_19786,N_19597);
and U19812 (N_19812,N_19783,N_19709);
xor U19813 (N_19813,N_19515,N_19680);
nand U19814 (N_19814,N_19667,N_19734);
and U19815 (N_19815,N_19538,N_19595);
nand U19816 (N_19816,N_19691,N_19712);
or U19817 (N_19817,N_19747,N_19634);
xor U19818 (N_19818,N_19689,N_19537);
or U19819 (N_19819,N_19707,N_19697);
nand U19820 (N_19820,N_19599,N_19509);
xnor U19821 (N_19821,N_19529,N_19548);
or U19822 (N_19822,N_19778,N_19521);
or U19823 (N_19823,N_19612,N_19505);
xnor U19824 (N_19824,N_19592,N_19640);
or U19825 (N_19825,N_19675,N_19581);
and U19826 (N_19826,N_19506,N_19642);
or U19827 (N_19827,N_19618,N_19768);
xor U19828 (N_19828,N_19589,N_19793);
or U19829 (N_19829,N_19552,N_19610);
nand U19830 (N_19830,N_19777,N_19731);
and U19831 (N_19831,N_19523,N_19751);
xor U19832 (N_19832,N_19795,N_19729);
and U19833 (N_19833,N_19790,N_19704);
xnor U19834 (N_19834,N_19759,N_19755);
xor U19835 (N_19835,N_19514,N_19666);
nand U19836 (N_19836,N_19658,N_19767);
and U19837 (N_19837,N_19573,N_19636);
or U19838 (N_19838,N_19614,N_19574);
xor U19839 (N_19839,N_19593,N_19530);
xor U19840 (N_19840,N_19564,N_19715);
xnor U19841 (N_19841,N_19796,N_19594);
nor U19842 (N_19842,N_19798,N_19742);
xnor U19843 (N_19843,N_19611,N_19519);
xnor U19844 (N_19844,N_19779,N_19566);
or U19845 (N_19845,N_19503,N_19671);
xor U19846 (N_19846,N_19763,N_19744);
nor U19847 (N_19847,N_19797,N_19532);
or U19848 (N_19848,N_19765,N_19621);
nand U19849 (N_19849,N_19739,N_19769);
nand U19850 (N_19850,N_19746,N_19639);
nand U19851 (N_19851,N_19668,N_19588);
and U19852 (N_19852,N_19624,N_19665);
nor U19853 (N_19853,N_19708,N_19590);
nor U19854 (N_19854,N_19560,N_19698);
nand U19855 (N_19855,N_19683,N_19717);
xnor U19856 (N_19856,N_19638,N_19569);
xor U19857 (N_19857,N_19679,N_19794);
nor U19858 (N_19858,N_19622,N_19605);
nor U19859 (N_19859,N_19511,N_19733);
or U19860 (N_19860,N_19602,N_19688);
xor U19861 (N_19861,N_19664,N_19785);
nor U19862 (N_19862,N_19587,N_19631);
xor U19863 (N_19863,N_19730,N_19549);
nor U19864 (N_19864,N_19702,N_19722);
or U19865 (N_19865,N_19727,N_19791);
and U19866 (N_19866,N_19782,N_19655);
or U19867 (N_19867,N_19726,N_19661);
nand U19868 (N_19868,N_19645,N_19695);
or U19869 (N_19869,N_19572,N_19585);
and U19870 (N_19870,N_19652,N_19559);
xor U19871 (N_19871,N_19555,N_19705);
nand U19872 (N_19872,N_19720,N_19780);
nor U19873 (N_19873,N_19539,N_19659);
xor U19874 (N_19874,N_19648,N_19604);
nand U19875 (N_19875,N_19654,N_19762);
xor U19876 (N_19876,N_19771,N_19644);
xnor U19877 (N_19877,N_19699,N_19627);
xor U19878 (N_19878,N_19682,N_19686);
or U19879 (N_19879,N_19651,N_19724);
nand U19880 (N_19880,N_19629,N_19637);
xnor U19881 (N_19881,N_19646,N_19580);
xnor U19882 (N_19882,N_19542,N_19556);
or U19883 (N_19883,N_19653,N_19567);
or U19884 (N_19884,N_19562,N_19632);
and U19885 (N_19885,N_19770,N_19527);
nor U19886 (N_19886,N_19756,N_19576);
nor U19887 (N_19887,N_19608,N_19526);
or U19888 (N_19888,N_19754,N_19656);
nand U19889 (N_19889,N_19570,N_19601);
nor U19890 (N_19890,N_19536,N_19535);
xnor U19891 (N_19891,N_19623,N_19540);
or U19892 (N_19892,N_19740,N_19554);
nor U19893 (N_19893,N_19513,N_19748);
xor U19894 (N_19894,N_19728,N_19713);
nor U19895 (N_19895,N_19617,N_19706);
nor U19896 (N_19896,N_19534,N_19591);
and U19897 (N_19897,N_19716,N_19545);
xor U19898 (N_19898,N_19524,N_19663);
and U19899 (N_19899,N_19583,N_19753);
nand U19900 (N_19900,N_19781,N_19694);
and U19901 (N_19901,N_19701,N_19558);
nand U19902 (N_19902,N_19619,N_19557);
nand U19903 (N_19903,N_19544,N_19690);
nand U19904 (N_19904,N_19792,N_19714);
or U19905 (N_19905,N_19518,N_19745);
or U19906 (N_19906,N_19672,N_19635);
xnor U19907 (N_19907,N_19626,N_19500);
or U19908 (N_19908,N_19504,N_19741);
xor U19909 (N_19909,N_19649,N_19776);
xnor U19910 (N_19910,N_19643,N_19673);
xnor U19911 (N_19911,N_19696,N_19579);
nor U19912 (N_19912,N_19757,N_19609);
nand U19913 (N_19913,N_19710,N_19773);
or U19914 (N_19914,N_19723,N_19516);
xor U19915 (N_19915,N_19799,N_19522);
xnor U19916 (N_19916,N_19507,N_19568);
or U19917 (N_19917,N_19766,N_19685);
and U19918 (N_19918,N_19775,N_19517);
nor U19919 (N_19919,N_19758,N_19647);
nand U19920 (N_19920,N_19703,N_19502);
nand U19921 (N_19921,N_19681,N_19737);
and U19922 (N_19922,N_19684,N_19508);
nor U19923 (N_19923,N_19606,N_19687);
nor U19924 (N_19924,N_19732,N_19501);
and U19925 (N_19925,N_19711,N_19561);
or U19926 (N_19926,N_19633,N_19764);
nand U19927 (N_19927,N_19630,N_19735);
or U19928 (N_19928,N_19546,N_19750);
and U19929 (N_19929,N_19575,N_19603);
or U19930 (N_19930,N_19787,N_19736);
nand U19931 (N_19931,N_19628,N_19657);
xnor U19932 (N_19932,N_19774,N_19615);
or U19933 (N_19933,N_19788,N_19525);
nor U19934 (N_19934,N_19718,N_19669);
xor U19935 (N_19935,N_19620,N_19700);
xor U19936 (N_19936,N_19752,N_19543);
nor U19937 (N_19937,N_19650,N_19743);
xnor U19938 (N_19938,N_19749,N_19598);
or U19939 (N_19939,N_19784,N_19565);
nor U19940 (N_19940,N_19551,N_19616);
or U19941 (N_19941,N_19760,N_19725);
xor U19942 (N_19942,N_19674,N_19641);
nor U19943 (N_19943,N_19550,N_19563);
xor U19944 (N_19944,N_19571,N_19607);
and U19945 (N_19945,N_19670,N_19676);
and U19946 (N_19946,N_19584,N_19533);
and U19947 (N_19947,N_19600,N_19596);
and U19948 (N_19948,N_19625,N_19541);
and U19949 (N_19949,N_19531,N_19677);
nor U19950 (N_19950,N_19657,N_19712);
nand U19951 (N_19951,N_19718,N_19644);
xor U19952 (N_19952,N_19572,N_19765);
nand U19953 (N_19953,N_19674,N_19548);
nor U19954 (N_19954,N_19755,N_19574);
or U19955 (N_19955,N_19774,N_19632);
xnor U19956 (N_19956,N_19692,N_19723);
or U19957 (N_19957,N_19782,N_19549);
nor U19958 (N_19958,N_19742,N_19603);
or U19959 (N_19959,N_19672,N_19725);
nor U19960 (N_19960,N_19524,N_19690);
and U19961 (N_19961,N_19641,N_19602);
or U19962 (N_19962,N_19774,N_19511);
xnor U19963 (N_19963,N_19568,N_19616);
and U19964 (N_19964,N_19639,N_19575);
nand U19965 (N_19965,N_19651,N_19580);
xnor U19966 (N_19966,N_19575,N_19791);
nand U19967 (N_19967,N_19792,N_19603);
nand U19968 (N_19968,N_19646,N_19683);
nand U19969 (N_19969,N_19664,N_19610);
and U19970 (N_19970,N_19578,N_19508);
xnor U19971 (N_19971,N_19675,N_19624);
or U19972 (N_19972,N_19709,N_19669);
nor U19973 (N_19973,N_19693,N_19581);
nand U19974 (N_19974,N_19557,N_19582);
nand U19975 (N_19975,N_19629,N_19781);
nor U19976 (N_19976,N_19598,N_19739);
nor U19977 (N_19977,N_19520,N_19787);
nor U19978 (N_19978,N_19725,N_19776);
or U19979 (N_19979,N_19709,N_19595);
xnor U19980 (N_19980,N_19777,N_19624);
xor U19981 (N_19981,N_19704,N_19706);
nand U19982 (N_19982,N_19520,N_19549);
nor U19983 (N_19983,N_19669,N_19654);
xnor U19984 (N_19984,N_19502,N_19673);
nand U19985 (N_19985,N_19518,N_19729);
and U19986 (N_19986,N_19585,N_19529);
nand U19987 (N_19987,N_19597,N_19695);
and U19988 (N_19988,N_19526,N_19679);
xor U19989 (N_19989,N_19512,N_19771);
xor U19990 (N_19990,N_19728,N_19778);
or U19991 (N_19991,N_19791,N_19721);
nand U19992 (N_19992,N_19564,N_19648);
nand U19993 (N_19993,N_19641,N_19606);
nor U19994 (N_19994,N_19596,N_19685);
nor U19995 (N_19995,N_19724,N_19535);
nor U19996 (N_19996,N_19748,N_19793);
xor U19997 (N_19997,N_19755,N_19655);
nand U19998 (N_19998,N_19687,N_19719);
and U19999 (N_19999,N_19729,N_19730);
xor U20000 (N_20000,N_19736,N_19512);
or U20001 (N_20001,N_19741,N_19556);
or U20002 (N_20002,N_19703,N_19782);
nand U20003 (N_20003,N_19543,N_19640);
nand U20004 (N_20004,N_19725,N_19554);
and U20005 (N_20005,N_19576,N_19644);
or U20006 (N_20006,N_19544,N_19624);
nor U20007 (N_20007,N_19697,N_19758);
nor U20008 (N_20008,N_19596,N_19576);
or U20009 (N_20009,N_19642,N_19668);
nand U20010 (N_20010,N_19527,N_19746);
or U20011 (N_20011,N_19659,N_19797);
or U20012 (N_20012,N_19599,N_19789);
or U20013 (N_20013,N_19510,N_19727);
nand U20014 (N_20014,N_19623,N_19782);
nand U20015 (N_20015,N_19711,N_19575);
nor U20016 (N_20016,N_19759,N_19746);
or U20017 (N_20017,N_19706,N_19707);
xnor U20018 (N_20018,N_19768,N_19711);
nand U20019 (N_20019,N_19729,N_19516);
nand U20020 (N_20020,N_19547,N_19613);
nand U20021 (N_20021,N_19543,N_19665);
and U20022 (N_20022,N_19613,N_19581);
or U20023 (N_20023,N_19541,N_19739);
nand U20024 (N_20024,N_19554,N_19737);
or U20025 (N_20025,N_19752,N_19791);
nand U20026 (N_20026,N_19744,N_19796);
xnor U20027 (N_20027,N_19596,N_19505);
and U20028 (N_20028,N_19708,N_19666);
xnor U20029 (N_20029,N_19670,N_19792);
nand U20030 (N_20030,N_19711,N_19715);
or U20031 (N_20031,N_19534,N_19541);
and U20032 (N_20032,N_19620,N_19609);
xnor U20033 (N_20033,N_19665,N_19690);
nand U20034 (N_20034,N_19678,N_19771);
xnor U20035 (N_20035,N_19724,N_19599);
nor U20036 (N_20036,N_19560,N_19737);
xnor U20037 (N_20037,N_19641,N_19592);
nor U20038 (N_20038,N_19657,N_19582);
xor U20039 (N_20039,N_19659,N_19683);
nand U20040 (N_20040,N_19792,N_19709);
nor U20041 (N_20041,N_19571,N_19623);
and U20042 (N_20042,N_19577,N_19681);
or U20043 (N_20043,N_19515,N_19779);
and U20044 (N_20044,N_19632,N_19531);
nand U20045 (N_20045,N_19556,N_19746);
xor U20046 (N_20046,N_19620,N_19554);
nor U20047 (N_20047,N_19656,N_19773);
and U20048 (N_20048,N_19728,N_19539);
xnor U20049 (N_20049,N_19606,N_19744);
nor U20050 (N_20050,N_19547,N_19610);
nor U20051 (N_20051,N_19544,N_19676);
nand U20052 (N_20052,N_19681,N_19580);
and U20053 (N_20053,N_19767,N_19508);
xnor U20054 (N_20054,N_19784,N_19753);
nand U20055 (N_20055,N_19576,N_19725);
nand U20056 (N_20056,N_19625,N_19515);
nand U20057 (N_20057,N_19788,N_19613);
xor U20058 (N_20058,N_19638,N_19630);
or U20059 (N_20059,N_19565,N_19664);
nor U20060 (N_20060,N_19698,N_19795);
and U20061 (N_20061,N_19685,N_19617);
and U20062 (N_20062,N_19714,N_19578);
or U20063 (N_20063,N_19525,N_19612);
nand U20064 (N_20064,N_19520,N_19673);
or U20065 (N_20065,N_19556,N_19611);
and U20066 (N_20066,N_19677,N_19500);
xor U20067 (N_20067,N_19776,N_19525);
xor U20068 (N_20068,N_19536,N_19646);
nor U20069 (N_20069,N_19600,N_19518);
nand U20070 (N_20070,N_19638,N_19501);
or U20071 (N_20071,N_19547,N_19672);
xnor U20072 (N_20072,N_19628,N_19663);
or U20073 (N_20073,N_19560,N_19568);
or U20074 (N_20074,N_19750,N_19669);
and U20075 (N_20075,N_19757,N_19720);
xnor U20076 (N_20076,N_19545,N_19651);
or U20077 (N_20077,N_19598,N_19621);
nand U20078 (N_20078,N_19604,N_19714);
nor U20079 (N_20079,N_19738,N_19606);
or U20080 (N_20080,N_19734,N_19719);
nand U20081 (N_20081,N_19514,N_19747);
xnor U20082 (N_20082,N_19542,N_19723);
or U20083 (N_20083,N_19509,N_19510);
nor U20084 (N_20084,N_19780,N_19644);
xnor U20085 (N_20085,N_19769,N_19637);
or U20086 (N_20086,N_19757,N_19583);
nand U20087 (N_20087,N_19611,N_19558);
xor U20088 (N_20088,N_19724,N_19646);
or U20089 (N_20089,N_19662,N_19716);
nor U20090 (N_20090,N_19703,N_19528);
nor U20091 (N_20091,N_19680,N_19519);
and U20092 (N_20092,N_19573,N_19671);
nor U20093 (N_20093,N_19595,N_19781);
nor U20094 (N_20094,N_19655,N_19596);
or U20095 (N_20095,N_19603,N_19576);
and U20096 (N_20096,N_19544,N_19761);
and U20097 (N_20097,N_19704,N_19559);
nor U20098 (N_20098,N_19588,N_19622);
or U20099 (N_20099,N_19791,N_19756);
xor U20100 (N_20100,N_19891,N_20044);
xnor U20101 (N_20101,N_19965,N_19812);
nor U20102 (N_20102,N_19807,N_20094);
or U20103 (N_20103,N_20018,N_20052);
or U20104 (N_20104,N_19810,N_19843);
xor U20105 (N_20105,N_19992,N_19951);
or U20106 (N_20106,N_20092,N_20078);
or U20107 (N_20107,N_20096,N_20083);
or U20108 (N_20108,N_19800,N_20025);
or U20109 (N_20109,N_19929,N_19892);
and U20110 (N_20110,N_19957,N_19846);
xnor U20111 (N_20111,N_19837,N_19808);
or U20112 (N_20112,N_19913,N_19968);
nor U20113 (N_20113,N_20088,N_19805);
or U20114 (N_20114,N_19956,N_19982);
xor U20115 (N_20115,N_19912,N_19860);
xnor U20116 (N_20116,N_20007,N_20039);
xor U20117 (N_20117,N_20010,N_20000);
xnor U20118 (N_20118,N_19842,N_19854);
nand U20119 (N_20119,N_20089,N_19889);
or U20120 (N_20120,N_19910,N_20066);
nor U20121 (N_20121,N_20059,N_20035);
xnor U20122 (N_20122,N_20067,N_20060);
nand U20123 (N_20123,N_19878,N_20081);
xnor U20124 (N_20124,N_19987,N_20051);
nand U20125 (N_20125,N_20040,N_20054);
nand U20126 (N_20126,N_20061,N_20056);
nor U20127 (N_20127,N_20047,N_19893);
and U20128 (N_20128,N_19950,N_20079);
or U20129 (N_20129,N_20042,N_19949);
or U20130 (N_20130,N_20012,N_19997);
or U20131 (N_20131,N_19820,N_19827);
and U20132 (N_20132,N_19862,N_19919);
nor U20133 (N_20133,N_19826,N_19848);
or U20134 (N_20134,N_19849,N_20020);
nand U20135 (N_20135,N_19993,N_19817);
nor U20136 (N_20136,N_19954,N_20053);
and U20137 (N_20137,N_19969,N_20099);
nand U20138 (N_20138,N_19888,N_19815);
nor U20139 (N_20139,N_19803,N_20085);
xnor U20140 (N_20140,N_20076,N_19941);
nand U20141 (N_20141,N_19962,N_20095);
nand U20142 (N_20142,N_20026,N_19847);
or U20143 (N_20143,N_19818,N_19911);
nand U20144 (N_20144,N_19833,N_19973);
and U20145 (N_20145,N_19813,N_19963);
nand U20146 (N_20146,N_20005,N_20086);
xnor U20147 (N_20147,N_19924,N_19985);
nand U20148 (N_20148,N_19885,N_19830);
nor U20149 (N_20149,N_20070,N_20055);
nor U20150 (N_20150,N_19852,N_19980);
or U20151 (N_20151,N_19900,N_19948);
nand U20152 (N_20152,N_19958,N_19850);
or U20153 (N_20153,N_19930,N_19974);
and U20154 (N_20154,N_19906,N_20038);
nand U20155 (N_20155,N_19864,N_19907);
nand U20156 (N_20156,N_19943,N_19855);
and U20157 (N_20157,N_20084,N_19867);
nor U20158 (N_20158,N_19875,N_19884);
nor U20159 (N_20159,N_20030,N_19880);
and U20160 (N_20160,N_19942,N_19981);
nand U20161 (N_20161,N_19845,N_20045);
nor U20162 (N_20162,N_19904,N_19897);
xor U20163 (N_20163,N_20090,N_19883);
nor U20164 (N_20164,N_19918,N_19881);
nor U20165 (N_20165,N_20082,N_19895);
and U20166 (N_20166,N_19866,N_19856);
and U20167 (N_20167,N_20062,N_20065);
nand U20168 (N_20168,N_19936,N_20075);
and U20169 (N_20169,N_20009,N_19931);
and U20170 (N_20170,N_19937,N_19976);
or U20171 (N_20171,N_20029,N_20036);
xnor U20172 (N_20172,N_19857,N_19814);
nor U20173 (N_20173,N_19841,N_19960);
xor U20174 (N_20174,N_19865,N_19986);
or U20175 (N_20175,N_20087,N_19995);
nand U20176 (N_20176,N_20023,N_19984);
xnor U20177 (N_20177,N_19970,N_20080);
nand U20178 (N_20178,N_19839,N_20073);
nand U20179 (N_20179,N_19999,N_20064);
or U20180 (N_20180,N_19945,N_19903);
nor U20181 (N_20181,N_19851,N_19834);
xor U20182 (N_20182,N_20046,N_20097);
or U20183 (N_20183,N_19836,N_19990);
and U20184 (N_20184,N_19994,N_19806);
xor U20185 (N_20185,N_20072,N_19923);
and U20186 (N_20186,N_19953,N_19894);
xnor U20187 (N_20187,N_19802,N_19838);
or U20188 (N_20188,N_19859,N_19868);
nor U20189 (N_20189,N_19955,N_19983);
nor U20190 (N_20190,N_19944,N_19917);
or U20191 (N_20191,N_19979,N_19873);
and U20192 (N_20192,N_19964,N_19946);
or U20193 (N_20193,N_19932,N_19840);
nand U20194 (N_20194,N_19832,N_20003);
nor U20195 (N_20195,N_19863,N_19988);
or U20196 (N_20196,N_19939,N_20011);
and U20197 (N_20197,N_19938,N_20071);
xor U20198 (N_20198,N_20063,N_19952);
nand U20199 (N_20199,N_20050,N_19921);
xor U20200 (N_20200,N_19972,N_19935);
xnor U20201 (N_20201,N_19804,N_19914);
xnor U20202 (N_20202,N_20033,N_20016);
xnor U20203 (N_20203,N_20037,N_19882);
nor U20204 (N_20204,N_20034,N_19801);
xnor U20205 (N_20205,N_19975,N_19966);
nand U20206 (N_20206,N_20002,N_20074);
or U20207 (N_20207,N_19874,N_20057);
xnor U20208 (N_20208,N_19824,N_19890);
nand U20209 (N_20209,N_19915,N_20006);
and U20210 (N_20210,N_20015,N_19821);
nor U20211 (N_20211,N_19896,N_19828);
xor U20212 (N_20212,N_19844,N_20017);
and U20213 (N_20213,N_19961,N_19901);
nand U20214 (N_20214,N_20098,N_19925);
xor U20215 (N_20215,N_19998,N_20058);
nor U20216 (N_20216,N_19927,N_19829);
nor U20217 (N_20217,N_20027,N_20014);
nand U20218 (N_20218,N_20019,N_19876);
xnor U20219 (N_20219,N_19899,N_20013);
xor U20220 (N_20220,N_19835,N_19928);
nor U20221 (N_20221,N_19869,N_19816);
nor U20222 (N_20222,N_19940,N_20004);
and U20223 (N_20223,N_20068,N_19991);
xor U20224 (N_20224,N_19861,N_19902);
and U20225 (N_20225,N_19916,N_19809);
nor U20226 (N_20226,N_20049,N_20048);
and U20227 (N_20227,N_19853,N_19967);
nor U20228 (N_20228,N_20043,N_19831);
nand U20229 (N_20229,N_20022,N_19823);
xnor U20230 (N_20230,N_20008,N_19870);
nand U20231 (N_20231,N_19871,N_20024);
nand U20232 (N_20232,N_19872,N_19977);
nand U20233 (N_20233,N_20032,N_20091);
and U20234 (N_20234,N_19922,N_20077);
or U20235 (N_20235,N_19822,N_20031);
nor U20236 (N_20236,N_20093,N_19971);
nand U20237 (N_20237,N_19825,N_20028);
or U20238 (N_20238,N_19877,N_19926);
nand U20239 (N_20239,N_19879,N_19858);
nor U20240 (N_20240,N_19898,N_20069);
and U20241 (N_20241,N_19887,N_19905);
nand U20242 (N_20242,N_19978,N_19908);
nand U20243 (N_20243,N_19811,N_19909);
nor U20244 (N_20244,N_19947,N_19920);
nor U20245 (N_20245,N_20041,N_19989);
and U20246 (N_20246,N_19819,N_20021);
or U20247 (N_20247,N_19996,N_19886);
and U20248 (N_20248,N_20001,N_19934);
nand U20249 (N_20249,N_19933,N_19959);
nor U20250 (N_20250,N_19820,N_20072);
nand U20251 (N_20251,N_20034,N_20066);
xor U20252 (N_20252,N_19862,N_20000);
nand U20253 (N_20253,N_19980,N_19836);
and U20254 (N_20254,N_19804,N_19991);
nand U20255 (N_20255,N_20046,N_19965);
or U20256 (N_20256,N_19871,N_20078);
or U20257 (N_20257,N_19986,N_20022);
xor U20258 (N_20258,N_19925,N_19951);
nand U20259 (N_20259,N_19915,N_19975);
or U20260 (N_20260,N_19922,N_19985);
nor U20261 (N_20261,N_19837,N_19872);
nand U20262 (N_20262,N_19960,N_20055);
xnor U20263 (N_20263,N_19851,N_19993);
nor U20264 (N_20264,N_20034,N_19910);
nand U20265 (N_20265,N_19874,N_19987);
and U20266 (N_20266,N_19928,N_20082);
nor U20267 (N_20267,N_20071,N_20076);
nand U20268 (N_20268,N_19892,N_20081);
and U20269 (N_20269,N_20010,N_19820);
and U20270 (N_20270,N_19802,N_19812);
nor U20271 (N_20271,N_19831,N_20077);
or U20272 (N_20272,N_20065,N_20024);
nand U20273 (N_20273,N_19919,N_20093);
nor U20274 (N_20274,N_19852,N_20024);
nor U20275 (N_20275,N_19883,N_20052);
and U20276 (N_20276,N_19953,N_19825);
xor U20277 (N_20277,N_20041,N_20048);
nor U20278 (N_20278,N_20089,N_19912);
or U20279 (N_20279,N_19987,N_20035);
nor U20280 (N_20280,N_19944,N_19992);
nor U20281 (N_20281,N_20078,N_20004);
or U20282 (N_20282,N_19869,N_19856);
and U20283 (N_20283,N_19965,N_19868);
or U20284 (N_20284,N_20067,N_20076);
or U20285 (N_20285,N_19912,N_19994);
nand U20286 (N_20286,N_19977,N_19973);
or U20287 (N_20287,N_20038,N_20018);
nand U20288 (N_20288,N_20053,N_20025);
or U20289 (N_20289,N_19879,N_19968);
nor U20290 (N_20290,N_19864,N_19961);
or U20291 (N_20291,N_20097,N_19854);
nor U20292 (N_20292,N_20013,N_20070);
or U20293 (N_20293,N_19846,N_19900);
nor U20294 (N_20294,N_19848,N_19999);
nand U20295 (N_20295,N_19869,N_19868);
nand U20296 (N_20296,N_19863,N_19981);
or U20297 (N_20297,N_19916,N_20054);
or U20298 (N_20298,N_19883,N_19947);
nor U20299 (N_20299,N_19995,N_19845);
xnor U20300 (N_20300,N_20057,N_19897);
or U20301 (N_20301,N_20030,N_19858);
nor U20302 (N_20302,N_20000,N_19993);
nand U20303 (N_20303,N_19904,N_19979);
and U20304 (N_20304,N_20011,N_20095);
nand U20305 (N_20305,N_19860,N_19837);
and U20306 (N_20306,N_19842,N_19906);
xnor U20307 (N_20307,N_19845,N_19896);
or U20308 (N_20308,N_20012,N_19950);
nand U20309 (N_20309,N_19923,N_19820);
nor U20310 (N_20310,N_19965,N_19809);
xor U20311 (N_20311,N_20099,N_19810);
xor U20312 (N_20312,N_19975,N_20080);
nand U20313 (N_20313,N_20046,N_20079);
xnor U20314 (N_20314,N_19862,N_20066);
nor U20315 (N_20315,N_19821,N_19848);
xnor U20316 (N_20316,N_20078,N_19949);
nand U20317 (N_20317,N_19918,N_19940);
and U20318 (N_20318,N_19922,N_20017);
nand U20319 (N_20319,N_19937,N_19939);
nor U20320 (N_20320,N_19802,N_19915);
nor U20321 (N_20321,N_19918,N_20010);
xnor U20322 (N_20322,N_19817,N_20034);
xor U20323 (N_20323,N_19933,N_19848);
and U20324 (N_20324,N_20051,N_19855);
nand U20325 (N_20325,N_19840,N_19875);
or U20326 (N_20326,N_19977,N_19941);
nand U20327 (N_20327,N_19986,N_20099);
nor U20328 (N_20328,N_19955,N_20057);
or U20329 (N_20329,N_19875,N_20071);
and U20330 (N_20330,N_19859,N_19867);
and U20331 (N_20331,N_19851,N_20021);
xnor U20332 (N_20332,N_19885,N_19948);
or U20333 (N_20333,N_20000,N_20062);
or U20334 (N_20334,N_19921,N_20011);
and U20335 (N_20335,N_19848,N_19931);
nor U20336 (N_20336,N_19966,N_20080);
nor U20337 (N_20337,N_19945,N_19994);
xor U20338 (N_20338,N_20017,N_19962);
xor U20339 (N_20339,N_20069,N_20002);
nand U20340 (N_20340,N_19910,N_20069);
or U20341 (N_20341,N_19836,N_19965);
or U20342 (N_20342,N_19888,N_19979);
nor U20343 (N_20343,N_19962,N_20005);
and U20344 (N_20344,N_20042,N_20048);
or U20345 (N_20345,N_19849,N_19992);
and U20346 (N_20346,N_19963,N_19907);
xnor U20347 (N_20347,N_19905,N_19826);
nor U20348 (N_20348,N_19980,N_19865);
and U20349 (N_20349,N_19857,N_19844);
xnor U20350 (N_20350,N_19873,N_20062);
nand U20351 (N_20351,N_20098,N_20010);
nor U20352 (N_20352,N_19891,N_19941);
or U20353 (N_20353,N_19828,N_20039);
and U20354 (N_20354,N_20029,N_19920);
and U20355 (N_20355,N_19942,N_19972);
xor U20356 (N_20356,N_19956,N_20057);
xor U20357 (N_20357,N_19807,N_19970);
and U20358 (N_20358,N_20073,N_19833);
or U20359 (N_20359,N_19872,N_19904);
nor U20360 (N_20360,N_19863,N_20075);
or U20361 (N_20361,N_19989,N_19943);
xor U20362 (N_20362,N_19995,N_19889);
xor U20363 (N_20363,N_19994,N_19876);
nand U20364 (N_20364,N_19818,N_19870);
or U20365 (N_20365,N_19876,N_19992);
and U20366 (N_20366,N_20026,N_19958);
nor U20367 (N_20367,N_19884,N_20066);
and U20368 (N_20368,N_19958,N_19937);
xnor U20369 (N_20369,N_19970,N_19963);
nand U20370 (N_20370,N_19877,N_19864);
nor U20371 (N_20371,N_19820,N_19860);
xnor U20372 (N_20372,N_19802,N_19834);
nand U20373 (N_20373,N_20080,N_19817);
nor U20374 (N_20374,N_19839,N_19855);
nand U20375 (N_20375,N_20066,N_19904);
or U20376 (N_20376,N_19968,N_20005);
nor U20377 (N_20377,N_19862,N_19910);
and U20378 (N_20378,N_19957,N_19848);
or U20379 (N_20379,N_20086,N_19912);
nand U20380 (N_20380,N_19934,N_19851);
xnor U20381 (N_20381,N_19969,N_20030);
nor U20382 (N_20382,N_19954,N_20068);
and U20383 (N_20383,N_20098,N_19817);
nand U20384 (N_20384,N_19987,N_19814);
nor U20385 (N_20385,N_19906,N_19952);
or U20386 (N_20386,N_19997,N_19822);
nand U20387 (N_20387,N_19953,N_19913);
nor U20388 (N_20388,N_19866,N_19858);
nand U20389 (N_20389,N_20064,N_19963);
nor U20390 (N_20390,N_19876,N_19803);
nand U20391 (N_20391,N_19921,N_19838);
xnor U20392 (N_20392,N_19856,N_20084);
or U20393 (N_20393,N_19969,N_19928);
nand U20394 (N_20394,N_20041,N_20007);
xnor U20395 (N_20395,N_19983,N_19956);
or U20396 (N_20396,N_19939,N_19912);
and U20397 (N_20397,N_19899,N_19938);
xnor U20398 (N_20398,N_19968,N_20078);
xor U20399 (N_20399,N_19989,N_19893);
or U20400 (N_20400,N_20200,N_20114);
nand U20401 (N_20401,N_20327,N_20180);
xnor U20402 (N_20402,N_20208,N_20108);
nor U20403 (N_20403,N_20139,N_20230);
xnor U20404 (N_20404,N_20357,N_20132);
xor U20405 (N_20405,N_20294,N_20118);
and U20406 (N_20406,N_20287,N_20104);
nor U20407 (N_20407,N_20315,N_20383);
and U20408 (N_20408,N_20236,N_20381);
or U20409 (N_20409,N_20159,N_20189);
and U20410 (N_20410,N_20188,N_20356);
nand U20411 (N_20411,N_20152,N_20196);
or U20412 (N_20412,N_20319,N_20329);
or U20413 (N_20413,N_20325,N_20115);
xor U20414 (N_20414,N_20359,N_20273);
xor U20415 (N_20415,N_20182,N_20295);
and U20416 (N_20416,N_20238,N_20246);
or U20417 (N_20417,N_20202,N_20393);
nor U20418 (N_20418,N_20312,N_20235);
and U20419 (N_20419,N_20268,N_20318);
nor U20420 (N_20420,N_20392,N_20142);
xor U20421 (N_20421,N_20293,N_20353);
nor U20422 (N_20422,N_20258,N_20223);
nand U20423 (N_20423,N_20323,N_20289);
xnor U20424 (N_20424,N_20270,N_20128);
xnor U20425 (N_20425,N_20156,N_20351);
nor U20426 (N_20426,N_20167,N_20212);
nand U20427 (N_20427,N_20251,N_20390);
nor U20428 (N_20428,N_20234,N_20121);
nor U20429 (N_20429,N_20310,N_20131);
xor U20430 (N_20430,N_20185,N_20197);
and U20431 (N_20431,N_20225,N_20346);
xor U20432 (N_20432,N_20370,N_20360);
nor U20433 (N_20433,N_20168,N_20333);
and U20434 (N_20434,N_20164,N_20116);
xnor U20435 (N_20435,N_20304,N_20307);
xor U20436 (N_20436,N_20379,N_20378);
or U20437 (N_20437,N_20240,N_20394);
or U20438 (N_20438,N_20317,N_20321);
xor U20439 (N_20439,N_20284,N_20369);
or U20440 (N_20440,N_20101,N_20338);
nor U20441 (N_20441,N_20179,N_20229);
xnor U20442 (N_20442,N_20172,N_20166);
nor U20443 (N_20443,N_20291,N_20146);
or U20444 (N_20444,N_20303,N_20178);
or U20445 (N_20445,N_20169,N_20140);
or U20446 (N_20446,N_20190,N_20395);
nand U20447 (N_20447,N_20271,N_20306);
or U20448 (N_20448,N_20122,N_20339);
nor U20449 (N_20449,N_20399,N_20102);
nor U20450 (N_20450,N_20385,N_20331);
or U20451 (N_20451,N_20214,N_20309);
and U20452 (N_20452,N_20382,N_20137);
xnor U20453 (N_20453,N_20123,N_20264);
and U20454 (N_20454,N_20100,N_20398);
nand U20455 (N_20455,N_20345,N_20361);
and U20456 (N_20456,N_20239,N_20124);
nor U20457 (N_20457,N_20285,N_20199);
nor U20458 (N_20458,N_20194,N_20191);
nor U20459 (N_20459,N_20371,N_20337);
nand U20460 (N_20460,N_20184,N_20155);
xnor U20461 (N_20461,N_20355,N_20372);
nand U20462 (N_20462,N_20219,N_20298);
nor U20463 (N_20463,N_20316,N_20389);
and U20464 (N_20464,N_20343,N_20396);
xor U20465 (N_20465,N_20148,N_20161);
or U20466 (N_20466,N_20244,N_20340);
nor U20467 (N_20467,N_20375,N_20320);
xor U20468 (N_20468,N_20377,N_20272);
or U20469 (N_20469,N_20130,N_20157);
nand U20470 (N_20470,N_20126,N_20133);
nor U20471 (N_20471,N_20233,N_20301);
or U20472 (N_20472,N_20231,N_20120);
xnor U20473 (N_20473,N_20143,N_20170);
and U20474 (N_20474,N_20109,N_20368);
xnor U20475 (N_20475,N_20342,N_20267);
xor U20476 (N_20476,N_20232,N_20127);
nor U20477 (N_20477,N_20335,N_20311);
nand U20478 (N_20478,N_20165,N_20313);
nor U20479 (N_20479,N_20384,N_20141);
and U20480 (N_20480,N_20218,N_20300);
and U20481 (N_20481,N_20162,N_20112);
xor U20482 (N_20482,N_20203,N_20247);
xnor U20483 (N_20483,N_20111,N_20220);
or U20484 (N_20484,N_20193,N_20269);
nand U20485 (N_20485,N_20279,N_20248);
or U20486 (N_20486,N_20263,N_20265);
nand U20487 (N_20487,N_20347,N_20243);
or U20488 (N_20488,N_20376,N_20228);
nor U20489 (N_20489,N_20107,N_20171);
and U20490 (N_20490,N_20255,N_20241);
and U20491 (N_20491,N_20158,N_20147);
nand U20492 (N_20492,N_20328,N_20217);
xnor U20493 (N_20493,N_20281,N_20282);
xor U20494 (N_20494,N_20324,N_20154);
or U20495 (N_20495,N_20245,N_20388);
nor U20496 (N_20496,N_20149,N_20174);
or U20497 (N_20497,N_20195,N_20129);
nand U20498 (N_20498,N_20134,N_20326);
nor U20499 (N_20499,N_20106,N_20297);
and U20500 (N_20500,N_20119,N_20397);
xnor U20501 (N_20501,N_20209,N_20144);
and U20502 (N_20502,N_20201,N_20103);
nor U20503 (N_20503,N_20286,N_20367);
or U20504 (N_20504,N_20322,N_20192);
xor U20505 (N_20505,N_20205,N_20387);
nand U20506 (N_20506,N_20253,N_20373);
or U20507 (N_20507,N_20336,N_20186);
nand U20508 (N_20508,N_20374,N_20183);
nand U20509 (N_20509,N_20177,N_20187);
and U20510 (N_20510,N_20283,N_20296);
nor U20511 (N_20511,N_20222,N_20262);
nor U20512 (N_20512,N_20150,N_20207);
xor U20513 (N_20513,N_20366,N_20237);
and U20514 (N_20514,N_20221,N_20135);
xnor U20515 (N_20515,N_20288,N_20341);
nor U20516 (N_20516,N_20254,N_20292);
xnor U20517 (N_20517,N_20198,N_20278);
nor U20518 (N_20518,N_20257,N_20176);
nor U20519 (N_20519,N_20227,N_20365);
nand U20520 (N_20520,N_20386,N_20117);
or U20521 (N_20521,N_20349,N_20216);
nand U20522 (N_20522,N_20210,N_20259);
nand U20523 (N_20523,N_20163,N_20277);
xnor U20524 (N_20524,N_20110,N_20354);
or U20525 (N_20525,N_20256,N_20334);
nor U20526 (N_20526,N_20260,N_20145);
xnor U20527 (N_20527,N_20364,N_20350);
or U20528 (N_20528,N_20160,N_20151);
xnor U20529 (N_20529,N_20249,N_20362);
xnor U20530 (N_20530,N_20358,N_20224);
nor U20531 (N_20531,N_20211,N_20274);
nand U20532 (N_20532,N_20363,N_20344);
nor U20533 (N_20533,N_20136,N_20276);
nor U20534 (N_20534,N_20242,N_20352);
nor U20535 (N_20535,N_20261,N_20275);
or U20536 (N_20536,N_20380,N_20252);
and U20537 (N_20537,N_20204,N_20302);
nand U20538 (N_20538,N_20215,N_20206);
and U20539 (N_20539,N_20308,N_20181);
nand U20540 (N_20540,N_20153,N_20250);
nor U20541 (N_20541,N_20330,N_20290);
xor U20542 (N_20542,N_20173,N_20213);
xnor U20543 (N_20543,N_20266,N_20175);
xor U20544 (N_20544,N_20138,N_20332);
nand U20545 (N_20545,N_20314,N_20105);
nand U20546 (N_20546,N_20113,N_20280);
nand U20547 (N_20547,N_20391,N_20226);
nand U20548 (N_20548,N_20125,N_20305);
and U20549 (N_20549,N_20299,N_20348);
or U20550 (N_20550,N_20342,N_20338);
or U20551 (N_20551,N_20319,N_20247);
nor U20552 (N_20552,N_20232,N_20396);
or U20553 (N_20553,N_20193,N_20189);
xnor U20554 (N_20554,N_20242,N_20374);
xor U20555 (N_20555,N_20238,N_20205);
nand U20556 (N_20556,N_20186,N_20256);
nor U20557 (N_20557,N_20324,N_20264);
and U20558 (N_20558,N_20365,N_20111);
xnor U20559 (N_20559,N_20278,N_20144);
nand U20560 (N_20560,N_20139,N_20278);
nand U20561 (N_20561,N_20140,N_20167);
and U20562 (N_20562,N_20156,N_20246);
nor U20563 (N_20563,N_20301,N_20236);
or U20564 (N_20564,N_20349,N_20176);
xor U20565 (N_20565,N_20210,N_20240);
or U20566 (N_20566,N_20338,N_20138);
or U20567 (N_20567,N_20214,N_20169);
xor U20568 (N_20568,N_20343,N_20137);
xnor U20569 (N_20569,N_20136,N_20105);
and U20570 (N_20570,N_20337,N_20206);
nor U20571 (N_20571,N_20272,N_20371);
and U20572 (N_20572,N_20317,N_20261);
and U20573 (N_20573,N_20370,N_20210);
and U20574 (N_20574,N_20198,N_20207);
xnor U20575 (N_20575,N_20204,N_20293);
nor U20576 (N_20576,N_20374,N_20241);
xor U20577 (N_20577,N_20171,N_20386);
or U20578 (N_20578,N_20391,N_20255);
and U20579 (N_20579,N_20254,N_20191);
xnor U20580 (N_20580,N_20290,N_20283);
nand U20581 (N_20581,N_20146,N_20223);
xnor U20582 (N_20582,N_20348,N_20289);
and U20583 (N_20583,N_20169,N_20125);
or U20584 (N_20584,N_20372,N_20228);
and U20585 (N_20585,N_20246,N_20197);
or U20586 (N_20586,N_20296,N_20298);
xnor U20587 (N_20587,N_20355,N_20239);
and U20588 (N_20588,N_20292,N_20223);
and U20589 (N_20589,N_20318,N_20360);
xor U20590 (N_20590,N_20242,N_20390);
nand U20591 (N_20591,N_20105,N_20177);
nand U20592 (N_20592,N_20113,N_20251);
nor U20593 (N_20593,N_20399,N_20101);
or U20594 (N_20594,N_20386,N_20193);
nor U20595 (N_20595,N_20264,N_20204);
xnor U20596 (N_20596,N_20111,N_20376);
xor U20597 (N_20597,N_20376,N_20147);
nor U20598 (N_20598,N_20361,N_20170);
or U20599 (N_20599,N_20122,N_20116);
or U20600 (N_20600,N_20198,N_20240);
and U20601 (N_20601,N_20339,N_20257);
and U20602 (N_20602,N_20112,N_20174);
or U20603 (N_20603,N_20397,N_20202);
nor U20604 (N_20604,N_20307,N_20255);
xor U20605 (N_20605,N_20313,N_20124);
and U20606 (N_20606,N_20272,N_20326);
or U20607 (N_20607,N_20216,N_20163);
or U20608 (N_20608,N_20374,N_20255);
nor U20609 (N_20609,N_20324,N_20131);
nor U20610 (N_20610,N_20269,N_20274);
nor U20611 (N_20611,N_20138,N_20346);
or U20612 (N_20612,N_20124,N_20310);
and U20613 (N_20613,N_20217,N_20123);
xor U20614 (N_20614,N_20303,N_20193);
nor U20615 (N_20615,N_20325,N_20355);
xor U20616 (N_20616,N_20339,N_20285);
nor U20617 (N_20617,N_20305,N_20136);
and U20618 (N_20618,N_20277,N_20109);
nor U20619 (N_20619,N_20367,N_20176);
nand U20620 (N_20620,N_20246,N_20161);
and U20621 (N_20621,N_20140,N_20161);
xor U20622 (N_20622,N_20105,N_20228);
xnor U20623 (N_20623,N_20261,N_20168);
xnor U20624 (N_20624,N_20151,N_20378);
nand U20625 (N_20625,N_20195,N_20180);
nor U20626 (N_20626,N_20156,N_20184);
nor U20627 (N_20627,N_20102,N_20283);
or U20628 (N_20628,N_20157,N_20383);
nand U20629 (N_20629,N_20303,N_20384);
or U20630 (N_20630,N_20396,N_20259);
nor U20631 (N_20631,N_20187,N_20366);
nand U20632 (N_20632,N_20291,N_20290);
xor U20633 (N_20633,N_20220,N_20201);
and U20634 (N_20634,N_20247,N_20186);
or U20635 (N_20635,N_20199,N_20203);
nand U20636 (N_20636,N_20176,N_20196);
and U20637 (N_20637,N_20359,N_20226);
nor U20638 (N_20638,N_20173,N_20291);
or U20639 (N_20639,N_20346,N_20243);
nor U20640 (N_20640,N_20112,N_20171);
or U20641 (N_20641,N_20327,N_20319);
nand U20642 (N_20642,N_20387,N_20190);
nor U20643 (N_20643,N_20381,N_20316);
and U20644 (N_20644,N_20173,N_20319);
and U20645 (N_20645,N_20164,N_20125);
xor U20646 (N_20646,N_20137,N_20109);
nand U20647 (N_20647,N_20317,N_20379);
nand U20648 (N_20648,N_20102,N_20327);
or U20649 (N_20649,N_20185,N_20189);
nor U20650 (N_20650,N_20238,N_20323);
and U20651 (N_20651,N_20323,N_20321);
xor U20652 (N_20652,N_20277,N_20215);
and U20653 (N_20653,N_20254,N_20323);
nand U20654 (N_20654,N_20164,N_20250);
nor U20655 (N_20655,N_20215,N_20230);
xnor U20656 (N_20656,N_20175,N_20261);
nor U20657 (N_20657,N_20284,N_20140);
or U20658 (N_20658,N_20221,N_20206);
nor U20659 (N_20659,N_20182,N_20342);
nor U20660 (N_20660,N_20358,N_20278);
and U20661 (N_20661,N_20223,N_20204);
or U20662 (N_20662,N_20234,N_20231);
and U20663 (N_20663,N_20376,N_20140);
or U20664 (N_20664,N_20328,N_20148);
nor U20665 (N_20665,N_20362,N_20224);
and U20666 (N_20666,N_20175,N_20134);
and U20667 (N_20667,N_20144,N_20399);
xor U20668 (N_20668,N_20303,N_20274);
or U20669 (N_20669,N_20255,N_20233);
nand U20670 (N_20670,N_20205,N_20341);
nor U20671 (N_20671,N_20199,N_20220);
or U20672 (N_20672,N_20387,N_20312);
and U20673 (N_20673,N_20141,N_20394);
nand U20674 (N_20674,N_20399,N_20308);
xor U20675 (N_20675,N_20393,N_20268);
or U20676 (N_20676,N_20275,N_20131);
nor U20677 (N_20677,N_20162,N_20208);
nor U20678 (N_20678,N_20205,N_20111);
nand U20679 (N_20679,N_20199,N_20146);
xor U20680 (N_20680,N_20171,N_20173);
and U20681 (N_20681,N_20136,N_20144);
nor U20682 (N_20682,N_20241,N_20171);
nor U20683 (N_20683,N_20122,N_20117);
nand U20684 (N_20684,N_20213,N_20165);
or U20685 (N_20685,N_20148,N_20108);
or U20686 (N_20686,N_20277,N_20328);
nand U20687 (N_20687,N_20344,N_20314);
nor U20688 (N_20688,N_20296,N_20174);
nand U20689 (N_20689,N_20271,N_20370);
or U20690 (N_20690,N_20247,N_20365);
or U20691 (N_20691,N_20206,N_20263);
xor U20692 (N_20692,N_20308,N_20149);
xor U20693 (N_20693,N_20241,N_20100);
and U20694 (N_20694,N_20273,N_20315);
or U20695 (N_20695,N_20200,N_20345);
or U20696 (N_20696,N_20173,N_20121);
nand U20697 (N_20697,N_20177,N_20291);
nand U20698 (N_20698,N_20360,N_20159);
nand U20699 (N_20699,N_20260,N_20215);
or U20700 (N_20700,N_20579,N_20633);
nand U20701 (N_20701,N_20447,N_20611);
and U20702 (N_20702,N_20471,N_20427);
nand U20703 (N_20703,N_20487,N_20689);
and U20704 (N_20704,N_20522,N_20478);
and U20705 (N_20705,N_20669,N_20465);
and U20706 (N_20706,N_20430,N_20652);
or U20707 (N_20707,N_20693,N_20437);
nor U20708 (N_20708,N_20537,N_20670);
xnor U20709 (N_20709,N_20668,N_20542);
nand U20710 (N_20710,N_20593,N_20483);
or U20711 (N_20711,N_20540,N_20557);
nor U20712 (N_20712,N_20494,N_20492);
and U20713 (N_20713,N_20495,N_20421);
and U20714 (N_20714,N_20516,N_20684);
and U20715 (N_20715,N_20449,N_20520);
and U20716 (N_20716,N_20418,N_20507);
nand U20717 (N_20717,N_20416,N_20550);
or U20718 (N_20718,N_20463,N_20554);
or U20719 (N_20719,N_20612,N_20588);
and U20720 (N_20720,N_20490,N_20543);
and U20721 (N_20721,N_20628,N_20451);
xor U20722 (N_20722,N_20691,N_20544);
xor U20723 (N_20723,N_20657,N_20622);
nor U20724 (N_20724,N_20623,N_20672);
nor U20725 (N_20725,N_20469,N_20577);
and U20726 (N_20726,N_20553,N_20667);
nand U20727 (N_20727,N_20545,N_20555);
xor U20728 (N_20728,N_20493,N_20404);
or U20729 (N_20729,N_20631,N_20400);
xnor U20730 (N_20730,N_20435,N_20629);
xor U20731 (N_20731,N_20662,N_20424);
xor U20732 (N_20732,N_20605,N_20444);
or U20733 (N_20733,N_20403,N_20582);
nand U20734 (N_20734,N_20446,N_20461);
and U20735 (N_20735,N_20408,N_20531);
or U20736 (N_20736,N_20517,N_20406);
nor U20737 (N_20737,N_20692,N_20674);
xnor U20738 (N_20738,N_20642,N_20509);
nand U20739 (N_20739,N_20431,N_20417);
and U20740 (N_20740,N_20491,N_20632);
nand U20741 (N_20741,N_20506,N_20534);
and U20742 (N_20742,N_20578,N_20666);
xor U20743 (N_20743,N_20499,N_20671);
nor U20744 (N_20744,N_20432,N_20525);
and U20745 (N_20745,N_20616,N_20586);
xnor U20746 (N_20746,N_20473,N_20502);
nor U20747 (N_20747,N_20414,N_20585);
nand U20748 (N_20748,N_20519,N_20452);
or U20749 (N_20749,N_20647,N_20618);
nor U20750 (N_20750,N_20590,N_20556);
nand U20751 (N_20751,N_20640,N_20453);
or U20752 (N_20752,N_20575,N_20485);
or U20753 (N_20753,N_20568,N_20475);
nand U20754 (N_20754,N_20570,N_20497);
nor U20755 (N_20755,N_20551,N_20442);
nor U20756 (N_20756,N_20694,N_20646);
or U20757 (N_20757,N_20619,N_20676);
nor U20758 (N_20758,N_20659,N_20466);
xnor U20759 (N_20759,N_20462,N_20472);
or U20760 (N_20760,N_20470,N_20594);
nor U20761 (N_20761,N_20539,N_20597);
or U20762 (N_20762,N_20614,N_20467);
and U20763 (N_20763,N_20411,N_20690);
nor U20764 (N_20764,N_20604,N_20439);
nor U20765 (N_20765,N_20602,N_20603);
nand U20766 (N_20766,N_20562,N_20501);
nor U20767 (N_20767,N_20533,N_20607);
and U20768 (N_20768,N_20587,N_20613);
and U20769 (N_20769,N_20455,N_20436);
nand U20770 (N_20770,N_20620,N_20584);
nand U20771 (N_20771,N_20675,N_20610);
nand U20772 (N_20772,N_20571,N_20630);
xnor U20773 (N_20773,N_20626,N_20526);
nor U20774 (N_20774,N_20569,N_20512);
xnor U20775 (N_20775,N_20634,N_20565);
or U20776 (N_20776,N_20420,N_20650);
nor U20777 (N_20777,N_20527,N_20637);
and U20778 (N_20778,N_20482,N_20655);
nand U20779 (N_20779,N_20589,N_20481);
and U20780 (N_20780,N_20649,N_20488);
and U20781 (N_20781,N_20425,N_20617);
nor U20782 (N_20782,N_20558,N_20687);
nor U20783 (N_20783,N_20561,N_20698);
and U20784 (N_20784,N_20643,N_20468);
xor U20785 (N_20785,N_20627,N_20685);
nand U20786 (N_20786,N_20592,N_20508);
xor U20787 (N_20787,N_20567,N_20529);
xor U20788 (N_20788,N_20412,N_20433);
nor U20789 (N_20789,N_20456,N_20673);
nor U20790 (N_20790,N_20479,N_20663);
nand U20791 (N_20791,N_20680,N_20625);
xor U20792 (N_20792,N_20688,N_20434);
or U20793 (N_20793,N_20648,N_20504);
and U20794 (N_20794,N_20496,N_20401);
and U20795 (N_20795,N_20598,N_20600);
or U20796 (N_20796,N_20419,N_20644);
xnor U20797 (N_20797,N_20665,N_20682);
or U20798 (N_20798,N_20615,N_20500);
xor U20799 (N_20799,N_20521,N_20679);
nor U20800 (N_20800,N_20523,N_20653);
nand U20801 (N_20801,N_20581,N_20503);
nor U20802 (N_20802,N_20528,N_20477);
xor U20803 (N_20803,N_20547,N_20515);
nand U20804 (N_20804,N_20664,N_20489);
nor U20805 (N_20805,N_20474,N_20450);
and U20806 (N_20806,N_20426,N_20410);
nor U20807 (N_20807,N_20448,N_20415);
nand U20808 (N_20808,N_20505,N_20660);
or U20809 (N_20809,N_20639,N_20645);
nor U20810 (N_20810,N_20651,N_20428);
or U20811 (N_20811,N_20566,N_20530);
or U20812 (N_20812,N_20596,N_20683);
and U20813 (N_20813,N_20443,N_20699);
nor U20814 (N_20814,N_20438,N_20697);
or U20815 (N_20815,N_20552,N_20641);
nor U20816 (N_20816,N_20514,N_20656);
and U20817 (N_20817,N_20621,N_20457);
nor U20818 (N_20818,N_20661,N_20548);
or U20819 (N_20819,N_20636,N_20572);
and U20820 (N_20820,N_20445,N_20638);
nor U20821 (N_20821,N_20624,N_20518);
or U20822 (N_20822,N_20599,N_20677);
nor U20823 (N_20823,N_20654,N_20460);
nand U20824 (N_20824,N_20429,N_20681);
nand U20825 (N_20825,N_20583,N_20459);
and U20826 (N_20826,N_20608,N_20484);
and U20827 (N_20827,N_20696,N_20532);
and U20828 (N_20828,N_20476,N_20409);
and U20829 (N_20829,N_20658,N_20536);
nand U20830 (N_20830,N_20511,N_20524);
nor U20831 (N_20831,N_20441,N_20458);
and U20832 (N_20832,N_20405,N_20498);
xor U20833 (N_20833,N_20606,N_20563);
or U20834 (N_20834,N_20573,N_20695);
nand U20835 (N_20835,N_20480,N_20546);
and U20836 (N_20836,N_20422,N_20609);
xnor U20837 (N_20837,N_20440,N_20564);
xnor U20838 (N_20838,N_20686,N_20464);
nor U20839 (N_20839,N_20591,N_20601);
and U20840 (N_20840,N_20486,N_20535);
nor U20841 (N_20841,N_20549,N_20513);
and U20842 (N_20842,N_20576,N_20423);
xor U20843 (N_20843,N_20580,N_20510);
nor U20844 (N_20844,N_20678,N_20413);
nor U20845 (N_20845,N_20635,N_20454);
and U20846 (N_20846,N_20560,N_20574);
nand U20847 (N_20847,N_20595,N_20402);
xor U20848 (N_20848,N_20541,N_20538);
or U20849 (N_20849,N_20407,N_20559);
and U20850 (N_20850,N_20615,N_20603);
xnor U20851 (N_20851,N_20442,N_20685);
xor U20852 (N_20852,N_20687,N_20544);
and U20853 (N_20853,N_20650,N_20563);
xor U20854 (N_20854,N_20671,N_20596);
nand U20855 (N_20855,N_20535,N_20426);
nor U20856 (N_20856,N_20628,N_20658);
and U20857 (N_20857,N_20464,N_20579);
or U20858 (N_20858,N_20428,N_20443);
xnor U20859 (N_20859,N_20631,N_20628);
nor U20860 (N_20860,N_20469,N_20573);
nand U20861 (N_20861,N_20595,N_20689);
and U20862 (N_20862,N_20452,N_20489);
xnor U20863 (N_20863,N_20630,N_20621);
or U20864 (N_20864,N_20534,N_20661);
and U20865 (N_20865,N_20435,N_20455);
and U20866 (N_20866,N_20659,N_20627);
or U20867 (N_20867,N_20600,N_20645);
nand U20868 (N_20868,N_20419,N_20688);
or U20869 (N_20869,N_20410,N_20584);
xnor U20870 (N_20870,N_20599,N_20681);
nor U20871 (N_20871,N_20550,N_20409);
and U20872 (N_20872,N_20666,N_20560);
and U20873 (N_20873,N_20548,N_20649);
xnor U20874 (N_20874,N_20408,N_20546);
and U20875 (N_20875,N_20443,N_20637);
and U20876 (N_20876,N_20413,N_20637);
and U20877 (N_20877,N_20427,N_20619);
nor U20878 (N_20878,N_20653,N_20502);
nor U20879 (N_20879,N_20665,N_20541);
nor U20880 (N_20880,N_20604,N_20424);
and U20881 (N_20881,N_20665,N_20510);
xor U20882 (N_20882,N_20546,N_20530);
nor U20883 (N_20883,N_20446,N_20517);
nand U20884 (N_20884,N_20520,N_20514);
xnor U20885 (N_20885,N_20456,N_20451);
and U20886 (N_20886,N_20506,N_20484);
xor U20887 (N_20887,N_20561,N_20443);
xor U20888 (N_20888,N_20582,N_20662);
or U20889 (N_20889,N_20590,N_20646);
xnor U20890 (N_20890,N_20405,N_20522);
xnor U20891 (N_20891,N_20679,N_20443);
xor U20892 (N_20892,N_20685,N_20416);
nor U20893 (N_20893,N_20656,N_20693);
nand U20894 (N_20894,N_20603,N_20675);
or U20895 (N_20895,N_20594,N_20634);
and U20896 (N_20896,N_20660,N_20417);
or U20897 (N_20897,N_20402,N_20464);
or U20898 (N_20898,N_20413,N_20407);
nor U20899 (N_20899,N_20437,N_20679);
nand U20900 (N_20900,N_20645,N_20411);
or U20901 (N_20901,N_20584,N_20456);
nand U20902 (N_20902,N_20585,N_20512);
or U20903 (N_20903,N_20620,N_20604);
xnor U20904 (N_20904,N_20645,N_20417);
nor U20905 (N_20905,N_20497,N_20615);
xnor U20906 (N_20906,N_20608,N_20420);
nor U20907 (N_20907,N_20474,N_20467);
nor U20908 (N_20908,N_20526,N_20462);
nand U20909 (N_20909,N_20415,N_20483);
nor U20910 (N_20910,N_20406,N_20443);
and U20911 (N_20911,N_20557,N_20488);
nor U20912 (N_20912,N_20516,N_20505);
nand U20913 (N_20913,N_20638,N_20628);
xor U20914 (N_20914,N_20412,N_20424);
nor U20915 (N_20915,N_20554,N_20541);
nand U20916 (N_20916,N_20476,N_20662);
nor U20917 (N_20917,N_20419,N_20694);
xor U20918 (N_20918,N_20527,N_20538);
xor U20919 (N_20919,N_20471,N_20498);
nand U20920 (N_20920,N_20651,N_20575);
and U20921 (N_20921,N_20508,N_20404);
and U20922 (N_20922,N_20663,N_20623);
and U20923 (N_20923,N_20572,N_20545);
xor U20924 (N_20924,N_20618,N_20555);
nor U20925 (N_20925,N_20480,N_20511);
xnor U20926 (N_20926,N_20697,N_20699);
nor U20927 (N_20927,N_20415,N_20547);
xnor U20928 (N_20928,N_20589,N_20511);
or U20929 (N_20929,N_20606,N_20480);
nor U20930 (N_20930,N_20555,N_20659);
or U20931 (N_20931,N_20696,N_20568);
nor U20932 (N_20932,N_20553,N_20610);
nor U20933 (N_20933,N_20600,N_20543);
xnor U20934 (N_20934,N_20412,N_20576);
xnor U20935 (N_20935,N_20406,N_20482);
nand U20936 (N_20936,N_20654,N_20502);
and U20937 (N_20937,N_20612,N_20691);
and U20938 (N_20938,N_20635,N_20642);
or U20939 (N_20939,N_20631,N_20472);
nand U20940 (N_20940,N_20680,N_20639);
or U20941 (N_20941,N_20688,N_20682);
nand U20942 (N_20942,N_20458,N_20424);
and U20943 (N_20943,N_20686,N_20671);
nor U20944 (N_20944,N_20688,N_20454);
xnor U20945 (N_20945,N_20465,N_20534);
nand U20946 (N_20946,N_20416,N_20483);
and U20947 (N_20947,N_20408,N_20459);
or U20948 (N_20948,N_20693,N_20580);
nand U20949 (N_20949,N_20487,N_20679);
xor U20950 (N_20950,N_20419,N_20611);
or U20951 (N_20951,N_20563,N_20490);
and U20952 (N_20952,N_20648,N_20507);
or U20953 (N_20953,N_20423,N_20521);
or U20954 (N_20954,N_20668,N_20657);
or U20955 (N_20955,N_20618,N_20419);
and U20956 (N_20956,N_20496,N_20406);
nand U20957 (N_20957,N_20678,N_20516);
or U20958 (N_20958,N_20545,N_20551);
nand U20959 (N_20959,N_20695,N_20565);
xnor U20960 (N_20960,N_20456,N_20644);
nor U20961 (N_20961,N_20639,N_20575);
and U20962 (N_20962,N_20562,N_20413);
and U20963 (N_20963,N_20678,N_20485);
and U20964 (N_20964,N_20603,N_20424);
or U20965 (N_20965,N_20454,N_20460);
and U20966 (N_20966,N_20625,N_20668);
nand U20967 (N_20967,N_20617,N_20599);
nand U20968 (N_20968,N_20563,N_20657);
and U20969 (N_20969,N_20623,N_20456);
nor U20970 (N_20970,N_20594,N_20674);
xnor U20971 (N_20971,N_20697,N_20633);
or U20972 (N_20972,N_20476,N_20612);
nand U20973 (N_20973,N_20487,N_20698);
and U20974 (N_20974,N_20672,N_20593);
or U20975 (N_20975,N_20418,N_20405);
xor U20976 (N_20976,N_20686,N_20609);
or U20977 (N_20977,N_20629,N_20505);
or U20978 (N_20978,N_20425,N_20653);
nand U20979 (N_20979,N_20691,N_20412);
xnor U20980 (N_20980,N_20508,N_20532);
xnor U20981 (N_20981,N_20627,N_20658);
and U20982 (N_20982,N_20584,N_20415);
and U20983 (N_20983,N_20453,N_20561);
nand U20984 (N_20984,N_20562,N_20478);
nor U20985 (N_20985,N_20585,N_20570);
nand U20986 (N_20986,N_20594,N_20602);
nand U20987 (N_20987,N_20692,N_20625);
or U20988 (N_20988,N_20557,N_20442);
or U20989 (N_20989,N_20581,N_20572);
xor U20990 (N_20990,N_20548,N_20645);
and U20991 (N_20991,N_20535,N_20694);
xnor U20992 (N_20992,N_20647,N_20514);
nor U20993 (N_20993,N_20616,N_20486);
nor U20994 (N_20994,N_20555,N_20559);
nand U20995 (N_20995,N_20691,N_20487);
xnor U20996 (N_20996,N_20562,N_20634);
or U20997 (N_20997,N_20556,N_20400);
or U20998 (N_20998,N_20574,N_20644);
nand U20999 (N_20999,N_20497,N_20660);
or U21000 (N_21000,N_20949,N_20890);
nor U21001 (N_21001,N_20700,N_20917);
nor U21002 (N_21002,N_20730,N_20825);
and U21003 (N_21003,N_20791,N_20860);
xor U21004 (N_21004,N_20862,N_20938);
nand U21005 (N_21005,N_20896,N_20839);
or U21006 (N_21006,N_20741,N_20876);
or U21007 (N_21007,N_20918,N_20882);
and U21008 (N_21008,N_20905,N_20824);
nand U21009 (N_21009,N_20924,N_20929);
and U21010 (N_21010,N_20992,N_20734);
and U21011 (N_21011,N_20977,N_20758);
xnor U21012 (N_21012,N_20980,N_20775);
nor U21013 (N_21013,N_20845,N_20806);
nand U21014 (N_21014,N_20897,N_20947);
nand U21015 (N_21015,N_20751,N_20837);
xnor U21016 (N_21016,N_20969,N_20927);
or U21017 (N_21017,N_20941,N_20979);
xnor U21018 (N_21018,N_20809,N_20867);
nor U21019 (N_21019,N_20945,N_20827);
nor U21020 (N_21020,N_20994,N_20735);
xnor U21021 (N_21021,N_20701,N_20963);
nor U21022 (N_21022,N_20884,N_20930);
xor U21023 (N_21023,N_20970,N_20871);
nand U21024 (N_21024,N_20966,N_20750);
and U21025 (N_21025,N_20936,N_20742);
nor U21026 (N_21026,N_20861,N_20712);
nand U21027 (N_21027,N_20747,N_20802);
nor U21028 (N_21028,N_20767,N_20740);
nand U21029 (N_21029,N_20958,N_20797);
and U21030 (N_21030,N_20965,N_20946);
nor U21031 (N_21031,N_20996,N_20810);
or U21032 (N_21032,N_20726,N_20848);
and U21033 (N_21033,N_20879,N_20940);
and U21034 (N_21034,N_20779,N_20836);
nor U21035 (N_21035,N_20989,N_20722);
nor U21036 (N_21036,N_20752,N_20816);
and U21037 (N_21037,N_20978,N_20898);
and U21038 (N_21038,N_20834,N_20826);
nand U21039 (N_21039,N_20737,N_20803);
nor U21040 (N_21040,N_20921,N_20983);
nand U21041 (N_21041,N_20870,N_20736);
and U21042 (N_21042,N_20909,N_20844);
nor U21043 (N_21043,N_20908,N_20768);
nand U21044 (N_21044,N_20894,N_20944);
nand U21045 (N_21045,N_20817,N_20785);
or U21046 (N_21046,N_20863,N_20888);
nor U21047 (N_21047,N_20968,N_20997);
nand U21048 (N_21048,N_20828,N_20832);
nand U21049 (N_21049,N_20986,N_20838);
nor U21050 (N_21050,N_20885,N_20973);
or U21051 (N_21051,N_20893,N_20928);
or U21052 (N_21052,N_20932,N_20985);
xnor U21053 (N_21053,N_20781,N_20998);
nor U21054 (N_21054,N_20960,N_20962);
and U21055 (N_21055,N_20883,N_20956);
xor U21056 (N_21056,N_20780,N_20759);
nor U21057 (N_21057,N_20872,N_20716);
and U21058 (N_21058,N_20784,N_20711);
nand U21059 (N_21059,N_20811,N_20991);
or U21060 (N_21060,N_20721,N_20895);
or U21061 (N_21061,N_20739,N_20913);
or U21062 (N_21062,N_20729,N_20774);
or U21063 (N_21063,N_20748,N_20934);
nand U21064 (N_21064,N_20902,N_20987);
xor U21065 (N_21065,N_20939,N_20813);
nor U21066 (N_21066,N_20812,N_20766);
and U21067 (N_21067,N_20852,N_20731);
nor U21068 (N_21068,N_20880,N_20942);
nand U21069 (N_21069,N_20818,N_20926);
or U21070 (N_21070,N_20807,N_20709);
or U21071 (N_21071,N_20822,N_20714);
nor U21072 (N_21072,N_20961,N_20795);
and U21073 (N_21073,N_20952,N_20821);
and U21074 (N_21074,N_20903,N_20976);
and U21075 (N_21075,N_20725,N_20702);
and U21076 (N_21076,N_20851,N_20873);
nor U21077 (N_21077,N_20793,N_20988);
nor U21078 (N_21078,N_20887,N_20910);
or U21079 (N_21079,N_20788,N_20866);
nand U21080 (N_21080,N_20943,N_20923);
or U21081 (N_21081,N_20857,N_20771);
and U21082 (N_21082,N_20981,N_20819);
nand U21083 (N_21083,N_20829,N_20972);
xnor U21084 (N_21084,N_20841,N_20782);
nor U21085 (N_21085,N_20899,N_20744);
and U21086 (N_21086,N_20990,N_20886);
or U21087 (N_21087,N_20764,N_20787);
xor U21088 (N_21088,N_20790,N_20765);
or U21089 (N_21089,N_20906,N_20763);
and U21090 (N_21090,N_20756,N_20911);
nand U21091 (N_21091,N_20877,N_20776);
and U21092 (N_21092,N_20955,N_20749);
and U21093 (N_21093,N_20892,N_20773);
xnor U21094 (N_21094,N_20935,N_20904);
xor U21095 (N_21095,N_20783,N_20874);
or U21096 (N_21096,N_20720,N_20717);
or U21097 (N_21097,N_20907,N_20919);
xor U21098 (N_21098,N_20953,N_20931);
xnor U21099 (N_21099,N_20761,N_20869);
xor U21100 (N_21100,N_20846,N_20833);
xor U21101 (N_21101,N_20933,N_20850);
or U21102 (N_21102,N_20772,N_20891);
nor U21103 (N_21103,N_20724,N_20999);
or U21104 (N_21104,N_20743,N_20964);
xor U21105 (N_21105,N_20814,N_20732);
or U21106 (N_21106,N_20753,N_20728);
nand U21107 (N_21107,N_20993,N_20937);
xnor U21108 (N_21108,N_20868,N_20796);
or U21109 (N_21109,N_20975,N_20995);
or U21110 (N_21110,N_20859,N_20733);
nand U21111 (N_21111,N_20912,N_20842);
and U21112 (N_21112,N_20875,N_20984);
and U21113 (N_21113,N_20957,N_20754);
nor U21114 (N_21114,N_20705,N_20914);
nor U21115 (N_21115,N_20703,N_20704);
or U21116 (N_21116,N_20715,N_20786);
or U21117 (N_21117,N_20755,N_20830);
nand U21118 (N_21118,N_20738,N_20922);
or U21119 (N_21119,N_20718,N_20770);
and U21120 (N_21120,N_20849,N_20878);
or U21121 (N_21121,N_20815,N_20920);
or U21122 (N_21122,N_20865,N_20925);
nor U21123 (N_21123,N_20881,N_20789);
xor U21124 (N_21124,N_20847,N_20727);
nor U21125 (N_21125,N_20982,N_20794);
nor U21126 (N_21126,N_20864,N_20915);
and U21127 (N_21127,N_20808,N_20954);
nand U21128 (N_21128,N_20719,N_20713);
or U21129 (N_21129,N_20799,N_20831);
and U21130 (N_21130,N_20801,N_20805);
nand U21131 (N_21131,N_20820,N_20757);
xor U21132 (N_21132,N_20835,N_20974);
nor U21133 (N_21133,N_20798,N_20948);
or U21134 (N_21134,N_20959,N_20708);
nor U21135 (N_21135,N_20777,N_20967);
or U21136 (N_21136,N_20823,N_20792);
nand U21137 (N_21137,N_20707,N_20745);
or U21138 (N_21138,N_20723,N_20800);
nand U21139 (N_21139,N_20706,N_20916);
nor U21140 (N_21140,N_20858,N_20971);
nand U21141 (N_21141,N_20843,N_20855);
and U21142 (N_21142,N_20760,N_20710);
nand U21143 (N_21143,N_20889,N_20854);
and U21144 (N_21144,N_20951,N_20900);
nor U21145 (N_21145,N_20901,N_20804);
or U21146 (N_21146,N_20762,N_20746);
xnor U21147 (N_21147,N_20856,N_20950);
xnor U21148 (N_21148,N_20778,N_20840);
nor U21149 (N_21149,N_20769,N_20853);
or U21150 (N_21150,N_20977,N_20801);
xnor U21151 (N_21151,N_20975,N_20953);
nand U21152 (N_21152,N_20818,N_20968);
nor U21153 (N_21153,N_20888,N_20809);
and U21154 (N_21154,N_20757,N_20911);
nand U21155 (N_21155,N_20724,N_20745);
nor U21156 (N_21156,N_20768,N_20819);
nor U21157 (N_21157,N_20979,N_20901);
nor U21158 (N_21158,N_20872,N_20869);
and U21159 (N_21159,N_20802,N_20735);
nand U21160 (N_21160,N_20725,N_20718);
nand U21161 (N_21161,N_20884,N_20955);
or U21162 (N_21162,N_20815,N_20821);
and U21163 (N_21163,N_20965,N_20800);
xnor U21164 (N_21164,N_20831,N_20996);
and U21165 (N_21165,N_20979,N_20706);
or U21166 (N_21166,N_20721,N_20889);
or U21167 (N_21167,N_20909,N_20772);
and U21168 (N_21168,N_20959,N_20817);
xor U21169 (N_21169,N_20723,N_20782);
and U21170 (N_21170,N_20891,N_20844);
nor U21171 (N_21171,N_20944,N_20942);
xor U21172 (N_21172,N_20742,N_20807);
nand U21173 (N_21173,N_20827,N_20954);
and U21174 (N_21174,N_20849,N_20999);
and U21175 (N_21175,N_20860,N_20777);
xor U21176 (N_21176,N_20790,N_20822);
or U21177 (N_21177,N_20763,N_20742);
xor U21178 (N_21178,N_20759,N_20945);
and U21179 (N_21179,N_20910,N_20727);
nor U21180 (N_21180,N_20742,N_20908);
and U21181 (N_21181,N_20767,N_20915);
nand U21182 (N_21182,N_20778,N_20724);
or U21183 (N_21183,N_20836,N_20979);
nand U21184 (N_21184,N_20741,N_20770);
nor U21185 (N_21185,N_20765,N_20835);
and U21186 (N_21186,N_20837,N_20729);
xor U21187 (N_21187,N_20990,N_20747);
or U21188 (N_21188,N_20888,N_20958);
or U21189 (N_21189,N_20838,N_20765);
and U21190 (N_21190,N_20926,N_20763);
or U21191 (N_21191,N_20906,N_20792);
or U21192 (N_21192,N_20701,N_20736);
xnor U21193 (N_21193,N_20712,N_20964);
xnor U21194 (N_21194,N_20904,N_20707);
and U21195 (N_21195,N_20843,N_20999);
nor U21196 (N_21196,N_20818,N_20701);
nand U21197 (N_21197,N_20889,N_20991);
nor U21198 (N_21198,N_20968,N_20994);
nor U21199 (N_21199,N_20922,N_20712);
and U21200 (N_21200,N_20719,N_20745);
nor U21201 (N_21201,N_20795,N_20820);
nor U21202 (N_21202,N_20829,N_20712);
nor U21203 (N_21203,N_20762,N_20728);
nor U21204 (N_21204,N_20980,N_20766);
nor U21205 (N_21205,N_20756,N_20775);
nor U21206 (N_21206,N_20898,N_20739);
and U21207 (N_21207,N_20871,N_20805);
and U21208 (N_21208,N_20839,N_20824);
nand U21209 (N_21209,N_20870,N_20778);
nor U21210 (N_21210,N_20933,N_20718);
xnor U21211 (N_21211,N_20998,N_20877);
xnor U21212 (N_21212,N_20963,N_20721);
and U21213 (N_21213,N_20941,N_20839);
nand U21214 (N_21214,N_20934,N_20792);
nand U21215 (N_21215,N_20713,N_20748);
nand U21216 (N_21216,N_20910,N_20886);
nor U21217 (N_21217,N_20813,N_20973);
and U21218 (N_21218,N_20734,N_20722);
or U21219 (N_21219,N_20721,N_20965);
nand U21220 (N_21220,N_20772,N_20738);
nand U21221 (N_21221,N_20709,N_20953);
and U21222 (N_21222,N_20985,N_20777);
xor U21223 (N_21223,N_20936,N_20976);
or U21224 (N_21224,N_20965,N_20932);
nand U21225 (N_21225,N_20903,N_20722);
xor U21226 (N_21226,N_20817,N_20793);
xor U21227 (N_21227,N_20855,N_20984);
or U21228 (N_21228,N_20712,N_20702);
or U21229 (N_21229,N_20923,N_20712);
and U21230 (N_21230,N_20882,N_20791);
xnor U21231 (N_21231,N_20977,N_20867);
nand U21232 (N_21232,N_20851,N_20842);
and U21233 (N_21233,N_20812,N_20794);
nor U21234 (N_21234,N_20871,N_20761);
and U21235 (N_21235,N_20829,N_20775);
xor U21236 (N_21236,N_20941,N_20921);
nor U21237 (N_21237,N_20901,N_20807);
or U21238 (N_21238,N_20785,N_20953);
nand U21239 (N_21239,N_20741,N_20897);
xor U21240 (N_21240,N_20951,N_20911);
nand U21241 (N_21241,N_20918,N_20800);
and U21242 (N_21242,N_20772,N_20870);
xor U21243 (N_21243,N_20836,N_20937);
or U21244 (N_21244,N_20794,N_20855);
nand U21245 (N_21245,N_20906,N_20825);
nor U21246 (N_21246,N_20727,N_20938);
and U21247 (N_21247,N_20781,N_20715);
xor U21248 (N_21248,N_20879,N_20846);
nor U21249 (N_21249,N_20991,N_20984);
nor U21250 (N_21250,N_20952,N_20788);
or U21251 (N_21251,N_20748,N_20774);
xor U21252 (N_21252,N_20736,N_20837);
nand U21253 (N_21253,N_20968,N_20923);
nor U21254 (N_21254,N_20782,N_20925);
nand U21255 (N_21255,N_20857,N_20846);
nor U21256 (N_21256,N_20869,N_20747);
xor U21257 (N_21257,N_20795,N_20756);
or U21258 (N_21258,N_20777,N_20788);
and U21259 (N_21259,N_20761,N_20812);
nand U21260 (N_21260,N_20786,N_20971);
xor U21261 (N_21261,N_20781,N_20828);
nor U21262 (N_21262,N_20787,N_20989);
nor U21263 (N_21263,N_20710,N_20749);
or U21264 (N_21264,N_20755,N_20883);
nor U21265 (N_21265,N_20779,N_20847);
or U21266 (N_21266,N_20904,N_20997);
or U21267 (N_21267,N_20976,N_20728);
and U21268 (N_21268,N_20858,N_20820);
xor U21269 (N_21269,N_20832,N_20901);
nor U21270 (N_21270,N_20984,N_20781);
nor U21271 (N_21271,N_20811,N_20877);
nor U21272 (N_21272,N_20714,N_20989);
nor U21273 (N_21273,N_20722,N_20716);
xor U21274 (N_21274,N_20720,N_20864);
xor U21275 (N_21275,N_20798,N_20926);
or U21276 (N_21276,N_20956,N_20869);
or U21277 (N_21277,N_20896,N_20993);
xor U21278 (N_21278,N_20787,N_20727);
xor U21279 (N_21279,N_20860,N_20864);
nand U21280 (N_21280,N_20993,N_20736);
nand U21281 (N_21281,N_20737,N_20702);
nor U21282 (N_21282,N_20851,N_20794);
nor U21283 (N_21283,N_20866,N_20895);
or U21284 (N_21284,N_20721,N_20799);
xnor U21285 (N_21285,N_20901,N_20894);
or U21286 (N_21286,N_20722,N_20781);
nor U21287 (N_21287,N_20773,N_20821);
and U21288 (N_21288,N_20924,N_20856);
or U21289 (N_21289,N_20895,N_20953);
xor U21290 (N_21290,N_20953,N_20980);
xor U21291 (N_21291,N_20775,N_20839);
nand U21292 (N_21292,N_20713,N_20722);
and U21293 (N_21293,N_20810,N_20825);
and U21294 (N_21294,N_20751,N_20771);
xnor U21295 (N_21295,N_20982,N_20986);
or U21296 (N_21296,N_20819,N_20887);
nor U21297 (N_21297,N_20996,N_20904);
nor U21298 (N_21298,N_20785,N_20759);
nor U21299 (N_21299,N_20911,N_20896);
and U21300 (N_21300,N_21121,N_21198);
nor U21301 (N_21301,N_21129,N_21107);
nor U21302 (N_21302,N_21002,N_21089);
nand U21303 (N_21303,N_21049,N_21112);
nor U21304 (N_21304,N_21061,N_21267);
nor U21305 (N_21305,N_21269,N_21152);
nor U21306 (N_21306,N_21035,N_21164);
xnor U21307 (N_21307,N_21253,N_21133);
and U21308 (N_21308,N_21060,N_21171);
xor U21309 (N_21309,N_21087,N_21252);
and U21310 (N_21310,N_21259,N_21230);
nor U21311 (N_21311,N_21177,N_21190);
nand U21312 (N_21312,N_21176,N_21038);
nor U21313 (N_21313,N_21104,N_21001);
nand U21314 (N_21314,N_21010,N_21017);
xnor U21315 (N_21315,N_21026,N_21231);
nor U21316 (N_21316,N_21139,N_21282);
xnor U21317 (N_21317,N_21195,N_21221);
nand U21318 (N_21318,N_21170,N_21039);
nand U21319 (N_21319,N_21042,N_21130);
xnor U21320 (N_21320,N_21100,N_21291);
xnor U21321 (N_21321,N_21288,N_21268);
nor U21322 (N_21322,N_21157,N_21261);
and U21323 (N_21323,N_21216,N_21080);
nand U21324 (N_21324,N_21147,N_21086);
nor U21325 (N_21325,N_21225,N_21120);
or U21326 (N_21326,N_21289,N_21169);
nor U21327 (N_21327,N_21296,N_21155);
nor U21328 (N_21328,N_21191,N_21223);
and U21329 (N_21329,N_21202,N_21141);
nand U21330 (N_21330,N_21031,N_21124);
or U21331 (N_21331,N_21123,N_21159);
xor U21332 (N_21332,N_21207,N_21209);
or U21333 (N_21333,N_21092,N_21197);
nor U21334 (N_21334,N_21113,N_21078);
nand U21335 (N_21335,N_21256,N_21237);
and U21336 (N_21336,N_21040,N_21236);
nand U21337 (N_21337,N_21199,N_21240);
xor U21338 (N_21338,N_21227,N_21137);
nor U21339 (N_21339,N_21142,N_21204);
or U21340 (N_21340,N_21229,N_21116);
xnor U21341 (N_21341,N_21108,N_21262);
and U21342 (N_21342,N_21166,N_21165);
xnor U21343 (N_21343,N_21295,N_21097);
nand U21344 (N_21344,N_21154,N_21136);
xnor U21345 (N_21345,N_21036,N_21016);
and U21346 (N_21346,N_21299,N_21298);
and U21347 (N_21347,N_21180,N_21072);
and U21348 (N_21348,N_21109,N_21075);
and U21349 (N_21349,N_21125,N_21009);
and U21350 (N_21350,N_21074,N_21015);
nand U21351 (N_21351,N_21096,N_21059);
and U21352 (N_21352,N_21069,N_21008);
xnor U21353 (N_21353,N_21029,N_21156);
nand U21354 (N_21354,N_21068,N_21127);
nand U21355 (N_21355,N_21064,N_21174);
nand U21356 (N_21356,N_21067,N_21255);
and U21357 (N_21357,N_21234,N_21258);
xnor U21358 (N_21358,N_21012,N_21247);
nor U21359 (N_21359,N_21119,N_21149);
nor U21360 (N_21360,N_21027,N_21297);
or U21361 (N_21361,N_21014,N_21025);
and U21362 (N_21362,N_21250,N_21224);
xnor U21363 (N_21363,N_21161,N_21238);
or U21364 (N_21364,N_21251,N_21030);
nor U21365 (N_21365,N_21028,N_21128);
or U21366 (N_21366,N_21287,N_21079);
and U21367 (N_21367,N_21265,N_21076);
and U21368 (N_21368,N_21126,N_21057);
and U21369 (N_21369,N_21274,N_21004);
xnor U21370 (N_21370,N_21150,N_21090);
or U21371 (N_21371,N_21219,N_21019);
nor U21372 (N_21372,N_21048,N_21056);
nor U21373 (N_21373,N_21117,N_21037);
nor U21374 (N_21374,N_21254,N_21003);
or U21375 (N_21375,N_21091,N_21073);
or U21376 (N_21376,N_21132,N_21077);
xnor U21377 (N_21377,N_21148,N_21228);
nand U21378 (N_21378,N_21110,N_21214);
nor U21379 (N_21379,N_21168,N_21115);
or U21380 (N_21380,N_21290,N_21145);
nor U21381 (N_21381,N_21275,N_21058);
or U21382 (N_21382,N_21102,N_21196);
nor U21383 (N_21383,N_21099,N_21245);
nand U21384 (N_21384,N_21182,N_21034);
nand U21385 (N_21385,N_21144,N_21217);
or U21386 (N_21386,N_21022,N_21242);
or U21387 (N_21387,N_21052,N_21140);
nor U21388 (N_21388,N_21101,N_21260);
nand U21389 (N_21389,N_21248,N_21095);
nor U21390 (N_21390,N_21226,N_21205);
or U21391 (N_21391,N_21283,N_21111);
nand U21392 (N_21392,N_21257,N_21071);
nor U21393 (N_21393,N_21000,N_21013);
or U21394 (N_21394,N_21206,N_21181);
and U21395 (N_21395,N_21044,N_21055);
and U21396 (N_21396,N_21193,N_21285);
and U21397 (N_21397,N_21280,N_21232);
or U21398 (N_21398,N_21188,N_21184);
or U21399 (N_21399,N_21246,N_21187);
xor U21400 (N_21400,N_21118,N_21192);
and U21401 (N_21401,N_21239,N_21098);
xor U21402 (N_21402,N_21281,N_21054);
nor U21403 (N_21403,N_21211,N_21158);
nand U21404 (N_21404,N_21050,N_21163);
and U21405 (N_21405,N_21011,N_21063);
xnor U21406 (N_21406,N_21143,N_21167);
nand U21407 (N_21407,N_21135,N_21083);
nor U21408 (N_21408,N_21006,N_21005);
nor U21409 (N_21409,N_21062,N_21183);
and U21410 (N_21410,N_21194,N_21189);
nor U21411 (N_21411,N_21277,N_21047);
nor U21412 (N_21412,N_21185,N_21200);
nand U21413 (N_21413,N_21160,N_21272);
nand U21414 (N_21414,N_21105,N_21276);
or U21415 (N_21415,N_21045,N_21210);
nand U21416 (N_21416,N_21203,N_21106);
xnor U21417 (N_21417,N_21131,N_21088);
nor U21418 (N_21418,N_21215,N_21093);
and U21419 (N_21419,N_21220,N_21235);
and U21420 (N_21420,N_21094,N_21294);
or U21421 (N_21421,N_21243,N_21208);
nand U21422 (N_21422,N_21271,N_21018);
xor U21423 (N_21423,N_21020,N_21046);
nor U21424 (N_21424,N_21053,N_21033);
xor U21425 (N_21425,N_21082,N_21043);
and U21426 (N_21426,N_21284,N_21172);
xor U21427 (N_21427,N_21293,N_21178);
nand U21428 (N_21428,N_21218,N_21233);
xor U21429 (N_21429,N_21153,N_21146);
or U21430 (N_21430,N_21024,N_21278);
or U21431 (N_21431,N_21270,N_21023);
xor U21432 (N_21432,N_21213,N_21175);
nand U21433 (N_21433,N_21292,N_21266);
or U21434 (N_21434,N_21279,N_21212);
or U21435 (N_21435,N_21273,N_21070);
nand U21436 (N_21436,N_21114,N_21032);
or U21437 (N_21437,N_21249,N_21007);
xnor U21438 (N_21438,N_21084,N_21241);
nand U21439 (N_21439,N_21138,N_21081);
xor U21440 (N_21440,N_21244,N_21286);
xor U21441 (N_21441,N_21103,N_21134);
or U21442 (N_21442,N_21122,N_21066);
nand U21443 (N_21443,N_21264,N_21162);
xor U21444 (N_21444,N_21085,N_21051);
and U21445 (N_21445,N_21222,N_21263);
xnor U21446 (N_21446,N_21201,N_21173);
xnor U21447 (N_21447,N_21151,N_21021);
nand U21448 (N_21448,N_21186,N_21179);
or U21449 (N_21449,N_21065,N_21041);
nor U21450 (N_21450,N_21110,N_21061);
nor U21451 (N_21451,N_21026,N_21200);
nor U21452 (N_21452,N_21086,N_21016);
nand U21453 (N_21453,N_21088,N_21176);
nor U21454 (N_21454,N_21131,N_21020);
and U21455 (N_21455,N_21235,N_21149);
and U21456 (N_21456,N_21061,N_21095);
nor U21457 (N_21457,N_21041,N_21040);
nand U21458 (N_21458,N_21099,N_21078);
or U21459 (N_21459,N_21004,N_21173);
and U21460 (N_21460,N_21163,N_21086);
and U21461 (N_21461,N_21152,N_21099);
nor U21462 (N_21462,N_21185,N_21155);
xor U21463 (N_21463,N_21289,N_21291);
and U21464 (N_21464,N_21160,N_21199);
xnor U21465 (N_21465,N_21250,N_21102);
nand U21466 (N_21466,N_21203,N_21162);
nand U21467 (N_21467,N_21188,N_21031);
nor U21468 (N_21468,N_21106,N_21130);
or U21469 (N_21469,N_21007,N_21216);
xor U21470 (N_21470,N_21157,N_21246);
nand U21471 (N_21471,N_21253,N_21098);
nor U21472 (N_21472,N_21161,N_21289);
xnor U21473 (N_21473,N_21268,N_21298);
or U21474 (N_21474,N_21053,N_21105);
nor U21475 (N_21475,N_21061,N_21283);
and U21476 (N_21476,N_21163,N_21085);
nand U21477 (N_21477,N_21010,N_21013);
and U21478 (N_21478,N_21189,N_21278);
nor U21479 (N_21479,N_21014,N_21209);
and U21480 (N_21480,N_21085,N_21036);
nor U21481 (N_21481,N_21242,N_21037);
nor U21482 (N_21482,N_21053,N_21226);
xor U21483 (N_21483,N_21075,N_21038);
nand U21484 (N_21484,N_21072,N_21148);
or U21485 (N_21485,N_21211,N_21112);
and U21486 (N_21486,N_21255,N_21230);
or U21487 (N_21487,N_21140,N_21165);
or U21488 (N_21488,N_21237,N_21147);
nor U21489 (N_21489,N_21040,N_21023);
nand U21490 (N_21490,N_21265,N_21060);
xnor U21491 (N_21491,N_21023,N_21279);
nor U21492 (N_21492,N_21227,N_21256);
and U21493 (N_21493,N_21114,N_21015);
or U21494 (N_21494,N_21298,N_21022);
nand U21495 (N_21495,N_21283,N_21293);
nand U21496 (N_21496,N_21050,N_21086);
xor U21497 (N_21497,N_21007,N_21058);
xor U21498 (N_21498,N_21030,N_21203);
or U21499 (N_21499,N_21050,N_21176);
nand U21500 (N_21500,N_21070,N_21279);
xor U21501 (N_21501,N_21224,N_21009);
xor U21502 (N_21502,N_21112,N_21185);
xnor U21503 (N_21503,N_21023,N_21277);
xor U21504 (N_21504,N_21003,N_21245);
or U21505 (N_21505,N_21063,N_21128);
and U21506 (N_21506,N_21207,N_21167);
and U21507 (N_21507,N_21146,N_21264);
or U21508 (N_21508,N_21186,N_21212);
xor U21509 (N_21509,N_21274,N_21220);
xor U21510 (N_21510,N_21206,N_21049);
and U21511 (N_21511,N_21283,N_21074);
xnor U21512 (N_21512,N_21146,N_21260);
or U21513 (N_21513,N_21148,N_21023);
or U21514 (N_21514,N_21005,N_21025);
and U21515 (N_21515,N_21145,N_21058);
nand U21516 (N_21516,N_21237,N_21253);
xnor U21517 (N_21517,N_21105,N_21130);
and U21518 (N_21518,N_21138,N_21076);
nand U21519 (N_21519,N_21145,N_21143);
xor U21520 (N_21520,N_21138,N_21034);
xnor U21521 (N_21521,N_21008,N_21107);
nand U21522 (N_21522,N_21149,N_21023);
nor U21523 (N_21523,N_21092,N_21142);
and U21524 (N_21524,N_21017,N_21283);
xor U21525 (N_21525,N_21022,N_21189);
xnor U21526 (N_21526,N_21149,N_21255);
and U21527 (N_21527,N_21257,N_21164);
nor U21528 (N_21528,N_21016,N_21261);
nand U21529 (N_21529,N_21078,N_21217);
and U21530 (N_21530,N_21252,N_21073);
xnor U21531 (N_21531,N_21228,N_21035);
nand U21532 (N_21532,N_21092,N_21042);
nand U21533 (N_21533,N_21226,N_21092);
nor U21534 (N_21534,N_21277,N_21100);
and U21535 (N_21535,N_21242,N_21175);
nand U21536 (N_21536,N_21106,N_21078);
or U21537 (N_21537,N_21169,N_21024);
or U21538 (N_21538,N_21002,N_21087);
nor U21539 (N_21539,N_21143,N_21189);
or U21540 (N_21540,N_21229,N_21188);
nor U21541 (N_21541,N_21199,N_21181);
nand U21542 (N_21542,N_21040,N_21047);
and U21543 (N_21543,N_21189,N_21003);
nor U21544 (N_21544,N_21163,N_21156);
and U21545 (N_21545,N_21008,N_21028);
nand U21546 (N_21546,N_21169,N_21050);
xnor U21547 (N_21547,N_21086,N_21125);
xor U21548 (N_21548,N_21036,N_21206);
and U21549 (N_21549,N_21007,N_21122);
nand U21550 (N_21550,N_21068,N_21096);
nand U21551 (N_21551,N_21137,N_21292);
or U21552 (N_21552,N_21010,N_21135);
xnor U21553 (N_21553,N_21030,N_21047);
nand U21554 (N_21554,N_21230,N_21241);
xor U21555 (N_21555,N_21049,N_21001);
or U21556 (N_21556,N_21051,N_21092);
nand U21557 (N_21557,N_21140,N_21085);
nand U21558 (N_21558,N_21117,N_21008);
nand U21559 (N_21559,N_21230,N_21164);
and U21560 (N_21560,N_21116,N_21259);
or U21561 (N_21561,N_21243,N_21034);
or U21562 (N_21562,N_21247,N_21279);
and U21563 (N_21563,N_21092,N_21060);
or U21564 (N_21564,N_21296,N_21126);
nor U21565 (N_21565,N_21146,N_21035);
nor U21566 (N_21566,N_21284,N_21105);
xnor U21567 (N_21567,N_21183,N_21299);
and U21568 (N_21568,N_21065,N_21058);
or U21569 (N_21569,N_21073,N_21044);
nor U21570 (N_21570,N_21119,N_21188);
nor U21571 (N_21571,N_21282,N_21197);
xnor U21572 (N_21572,N_21128,N_21209);
nor U21573 (N_21573,N_21270,N_21225);
nand U21574 (N_21574,N_21124,N_21241);
or U21575 (N_21575,N_21268,N_21231);
nand U21576 (N_21576,N_21063,N_21202);
nand U21577 (N_21577,N_21275,N_21037);
and U21578 (N_21578,N_21205,N_21249);
nor U21579 (N_21579,N_21212,N_21235);
and U21580 (N_21580,N_21129,N_21143);
or U21581 (N_21581,N_21221,N_21046);
xor U21582 (N_21582,N_21105,N_21242);
nor U21583 (N_21583,N_21103,N_21117);
nor U21584 (N_21584,N_21138,N_21024);
xor U21585 (N_21585,N_21247,N_21278);
nor U21586 (N_21586,N_21055,N_21274);
nor U21587 (N_21587,N_21149,N_21062);
nand U21588 (N_21588,N_21124,N_21105);
xnor U21589 (N_21589,N_21228,N_21144);
and U21590 (N_21590,N_21214,N_21177);
xor U21591 (N_21591,N_21016,N_21298);
and U21592 (N_21592,N_21153,N_21004);
nand U21593 (N_21593,N_21198,N_21046);
nor U21594 (N_21594,N_21006,N_21128);
xnor U21595 (N_21595,N_21220,N_21198);
xnor U21596 (N_21596,N_21222,N_21285);
xnor U21597 (N_21597,N_21086,N_21272);
and U21598 (N_21598,N_21070,N_21064);
nor U21599 (N_21599,N_21131,N_21009);
xnor U21600 (N_21600,N_21491,N_21469);
nor U21601 (N_21601,N_21407,N_21429);
and U21602 (N_21602,N_21340,N_21401);
and U21603 (N_21603,N_21310,N_21346);
nor U21604 (N_21604,N_21410,N_21446);
nand U21605 (N_21605,N_21355,N_21348);
and U21606 (N_21606,N_21363,N_21399);
xor U21607 (N_21607,N_21513,N_21328);
or U21608 (N_21608,N_21305,N_21307);
xnor U21609 (N_21609,N_21406,N_21441);
xnor U21610 (N_21610,N_21501,N_21336);
or U21611 (N_21611,N_21338,N_21487);
nand U21612 (N_21612,N_21524,N_21466);
nand U21613 (N_21613,N_21594,N_21538);
nand U21614 (N_21614,N_21558,N_21312);
nor U21615 (N_21615,N_21499,N_21376);
or U21616 (N_21616,N_21511,N_21489);
nor U21617 (N_21617,N_21564,N_21563);
nor U21618 (N_21618,N_21554,N_21368);
xor U21619 (N_21619,N_21536,N_21395);
nand U21620 (N_21620,N_21521,N_21349);
nor U21621 (N_21621,N_21303,N_21381);
xor U21622 (N_21622,N_21343,N_21560);
or U21623 (N_21623,N_21551,N_21337);
xor U21624 (N_21624,N_21448,N_21315);
xnor U21625 (N_21625,N_21475,N_21582);
and U21626 (N_21626,N_21514,N_21530);
nand U21627 (N_21627,N_21393,N_21592);
nand U21628 (N_21628,N_21414,N_21552);
or U21629 (N_21629,N_21413,N_21300);
nand U21630 (N_21630,N_21484,N_21308);
nand U21631 (N_21631,N_21492,N_21557);
and U21632 (N_21632,N_21588,N_21593);
xnor U21633 (N_21633,N_21463,N_21423);
nor U21634 (N_21634,N_21540,N_21474);
or U21635 (N_21635,N_21544,N_21498);
xnor U21636 (N_21636,N_21431,N_21546);
nand U21637 (N_21637,N_21437,N_21462);
xnor U21638 (N_21638,N_21411,N_21573);
or U21639 (N_21639,N_21380,N_21311);
nand U21640 (N_21640,N_21433,N_21365);
nand U21641 (N_21641,N_21319,N_21317);
xnor U21642 (N_21642,N_21476,N_21589);
nor U21643 (N_21643,N_21427,N_21494);
xnor U21644 (N_21644,N_21534,N_21358);
nand U21645 (N_21645,N_21532,N_21364);
or U21646 (N_21646,N_21458,N_21331);
nor U21647 (N_21647,N_21506,N_21374);
nor U21648 (N_21648,N_21559,N_21490);
or U21649 (N_21649,N_21528,N_21581);
xor U21650 (N_21650,N_21412,N_21516);
nor U21651 (N_21651,N_21525,N_21339);
and U21652 (N_21652,N_21424,N_21495);
nor U21653 (N_21653,N_21415,N_21493);
nand U21654 (N_21654,N_21370,N_21366);
xor U21655 (N_21655,N_21353,N_21596);
and U21656 (N_21656,N_21527,N_21359);
nand U21657 (N_21657,N_21396,N_21575);
xnor U21658 (N_21658,N_21464,N_21459);
xnor U21659 (N_21659,N_21488,N_21599);
nand U21660 (N_21660,N_21425,N_21426);
nand U21661 (N_21661,N_21482,N_21480);
and U21662 (N_21662,N_21377,N_21409);
xor U21663 (N_21663,N_21422,N_21379);
or U21664 (N_21664,N_21361,N_21390);
xnor U21665 (N_21665,N_21419,N_21435);
xor U21666 (N_21666,N_21460,N_21496);
or U21667 (N_21667,N_21590,N_21509);
xnor U21668 (N_21668,N_21510,N_21342);
xnor U21669 (N_21669,N_21391,N_21595);
or U21670 (N_21670,N_21321,N_21545);
nor U21671 (N_21671,N_21354,N_21447);
nor U21672 (N_21672,N_21565,N_21372);
nand U21673 (N_21673,N_21392,N_21486);
and U21674 (N_21674,N_21378,N_21522);
nor U21675 (N_21675,N_21455,N_21541);
and U21676 (N_21676,N_21316,N_21485);
and U21677 (N_21677,N_21301,N_21576);
or U21678 (N_21678,N_21334,N_21497);
or U21679 (N_21679,N_21443,N_21386);
xor U21680 (N_21680,N_21345,N_21335);
and U21681 (N_21681,N_21561,N_21539);
or U21682 (N_21682,N_21453,N_21542);
or U21683 (N_21683,N_21397,N_21318);
nor U21684 (N_21684,N_21577,N_21529);
nand U21685 (N_21685,N_21327,N_21450);
nand U21686 (N_21686,N_21531,N_21304);
nor U21687 (N_21687,N_21325,N_21333);
nor U21688 (N_21688,N_21585,N_21535);
or U21689 (N_21689,N_21389,N_21385);
and U21690 (N_21690,N_21436,N_21357);
nand U21691 (N_21691,N_21313,N_21580);
and U21692 (N_21692,N_21508,N_21445);
nand U21693 (N_21693,N_21512,N_21586);
xor U21694 (N_21694,N_21356,N_21418);
nand U21695 (N_21695,N_21550,N_21571);
nand U21696 (N_21696,N_21520,N_21519);
and U21697 (N_21697,N_21449,N_21347);
nand U21698 (N_21698,N_21440,N_21421);
and U21699 (N_21699,N_21382,N_21387);
or U21700 (N_21700,N_21481,N_21583);
xnor U21701 (N_21701,N_21587,N_21434);
nor U21702 (N_21702,N_21457,N_21362);
nor U21703 (N_21703,N_21574,N_21330);
nor U21704 (N_21704,N_21504,N_21373);
xnor U21705 (N_21705,N_21537,N_21526);
and U21706 (N_21706,N_21548,N_21430);
and U21707 (N_21707,N_21302,N_21444);
xnor U21708 (N_21708,N_21470,N_21468);
or U21709 (N_21709,N_21405,N_21329);
xnor U21710 (N_21710,N_21523,N_21420);
xor U21711 (N_21711,N_21597,N_21467);
xor U21712 (N_21712,N_21322,N_21326);
nor U21713 (N_21713,N_21473,N_21478);
or U21714 (N_21714,N_21432,N_21360);
nand U21715 (N_21715,N_21454,N_21567);
and U21716 (N_21716,N_21394,N_21584);
and U21717 (N_21717,N_21344,N_21384);
nand U21718 (N_21718,N_21369,N_21533);
nor U21719 (N_21719,N_21598,N_21518);
or U21720 (N_21720,N_21483,N_21439);
or U21721 (N_21721,N_21579,N_21416);
xnor U21722 (N_21722,N_21309,N_21549);
xnor U21723 (N_21723,N_21367,N_21479);
or U21724 (N_21724,N_21403,N_21591);
xnor U21725 (N_21725,N_21562,N_21351);
or U21726 (N_21726,N_21383,N_21438);
or U21727 (N_21727,N_21572,N_21507);
and U21728 (N_21728,N_21569,N_21461);
and U21729 (N_21729,N_21400,N_21332);
nand U21730 (N_21730,N_21428,N_21408);
and U21731 (N_21731,N_21556,N_21388);
and U21732 (N_21732,N_21472,N_21352);
or U21733 (N_21733,N_21503,N_21375);
nor U21734 (N_21734,N_21341,N_21477);
nand U21735 (N_21735,N_21417,N_21555);
xnor U21736 (N_21736,N_21324,N_21500);
or U21737 (N_21737,N_21320,N_21505);
nand U21738 (N_21738,N_21456,N_21465);
nor U21739 (N_21739,N_21502,N_21547);
or U21740 (N_21740,N_21471,N_21566);
nand U21741 (N_21741,N_21570,N_21553);
and U21742 (N_21742,N_21451,N_21323);
xnor U21743 (N_21743,N_21398,N_21578);
nand U21744 (N_21744,N_21350,N_21402);
and U21745 (N_21745,N_21371,N_21452);
nor U21746 (N_21746,N_21306,N_21404);
and U21747 (N_21747,N_21515,N_21543);
and U21748 (N_21748,N_21442,N_21568);
nor U21749 (N_21749,N_21314,N_21517);
nor U21750 (N_21750,N_21429,N_21589);
or U21751 (N_21751,N_21513,N_21379);
xnor U21752 (N_21752,N_21563,N_21335);
xnor U21753 (N_21753,N_21396,N_21519);
or U21754 (N_21754,N_21535,N_21374);
nand U21755 (N_21755,N_21596,N_21457);
or U21756 (N_21756,N_21312,N_21448);
nor U21757 (N_21757,N_21417,N_21590);
xnor U21758 (N_21758,N_21532,N_21497);
nor U21759 (N_21759,N_21489,N_21405);
and U21760 (N_21760,N_21420,N_21392);
xor U21761 (N_21761,N_21409,N_21473);
nor U21762 (N_21762,N_21358,N_21498);
xor U21763 (N_21763,N_21408,N_21480);
xnor U21764 (N_21764,N_21320,N_21350);
and U21765 (N_21765,N_21483,N_21539);
and U21766 (N_21766,N_21467,N_21439);
nor U21767 (N_21767,N_21369,N_21465);
nand U21768 (N_21768,N_21564,N_21320);
and U21769 (N_21769,N_21331,N_21375);
nor U21770 (N_21770,N_21317,N_21562);
nor U21771 (N_21771,N_21549,N_21349);
xor U21772 (N_21772,N_21566,N_21362);
xnor U21773 (N_21773,N_21507,N_21464);
xor U21774 (N_21774,N_21490,N_21393);
and U21775 (N_21775,N_21377,N_21558);
and U21776 (N_21776,N_21370,N_21456);
nor U21777 (N_21777,N_21573,N_21498);
nand U21778 (N_21778,N_21540,N_21321);
or U21779 (N_21779,N_21460,N_21560);
or U21780 (N_21780,N_21345,N_21523);
or U21781 (N_21781,N_21461,N_21578);
xor U21782 (N_21782,N_21313,N_21309);
xor U21783 (N_21783,N_21380,N_21385);
nor U21784 (N_21784,N_21424,N_21381);
nand U21785 (N_21785,N_21445,N_21571);
or U21786 (N_21786,N_21380,N_21475);
or U21787 (N_21787,N_21451,N_21581);
xor U21788 (N_21788,N_21541,N_21397);
xor U21789 (N_21789,N_21570,N_21488);
and U21790 (N_21790,N_21516,N_21337);
and U21791 (N_21791,N_21443,N_21545);
xnor U21792 (N_21792,N_21564,N_21457);
nor U21793 (N_21793,N_21573,N_21307);
or U21794 (N_21794,N_21393,N_21404);
nand U21795 (N_21795,N_21401,N_21582);
and U21796 (N_21796,N_21523,N_21542);
xor U21797 (N_21797,N_21548,N_21449);
xor U21798 (N_21798,N_21361,N_21332);
nand U21799 (N_21799,N_21446,N_21303);
xor U21800 (N_21800,N_21380,N_21592);
and U21801 (N_21801,N_21497,N_21389);
nor U21802 (N_21802,N_21492,N_21523);
or U21803 (N_21803,N_21481,N_21448);
and U21804 (N_21804,N_21598,N_21371);
or U21805 (N_21805,N_21593,N_21314);
nor U21806 (N_21806,N_21599,N_21437);
xor U21807 (N_21807,N_21564,N_21423);
nor U21808 (N_21808,N_21383,N_21409);
and U21809 (N_21809,N_21414,N_21472);
xor U21810 (N_21810,N_21441,N_21575);
xnor U21811 (N_21811,N_21403,N_21466);
and U21812 (N_21812,N_21442,N_21528);
nor U21813 (N_21813,N_21341,N_21594);
or U21814 (N_21814,N_21470,N_21521);
or U21815 (N_21815,N_21383,N_21379);
and U21816 (N_21816,N_21480,N_21575);
xor U21817 (N_21817,N_21374,N_21554);
xor U21818 (N_21818,N_21366,N_21308);
xnor U21819 (N_21819,N_21496,N_21349);
xnor U21820 (N_21820,N_21432,N_21410);
xor U21821 (N_21821,N_21356,N_21511);
nor U21822 (N_21822,N_21577,N_21588);
nor U21823 (N_21823,N_21513,N_21308);
and U21824 (N_21824,N_21354,N_21514);
nor U21825 (N_21825,N_21504,N_21524);
or U21826 (N_21826,N_21502,N_21348);
or U21827 (N_21827,N_21548,N_21518);
or U21828 (N_21828,N_21440,N_21573);
nor U21829 (N_21829,N_21565,N_21395);
nor U21830 (N_21830,N_21333,N_21393);
xor U21831 (N_21831,N_21399,N_21377);
and U21832 (N_21832,N_21358,N_21373);
and U21833 (N_21833,N_21528,N_21579);
nand U21834 (N_21834,N_21571,N_21584);
nand U21835 (N_21835,N_21509,N_21501);
or U21836 (N_21836,N_21356,N_21408);
xnor U21837 (N_21837,N_21565,N_21437);
and U21838 (N_21838,N_21497,N_21508);
or U21839 (N_21839,N_21308,N_21390);
or U21840 (N_21840,N_21561,N_21501);
xnor U21841 (N_21841,N_21440,N_21337);
xor U21842 (N_21842,N_21480,N_21471);
and U21843 (N_21843,N_21595,N_21465);
and U21844 (N_21844,N_21545,N_21502);
and U21845 (N_21845,N_21593,N_21478);
and U21846 (N_21846,N_21412,N_21464);
or U21847 (N_21847,N_21310,N_21590);
nor U21848 (N_21848,N_21317,N_21434);
or U21849 (N_21849,N_21566,N_21572);
xor U21850 (N_21850,N_21497,N_21383);
or U21851 (N_21851,N_21368,N_21418);
nand U21852 (N_21852,N_21309,N_21444);
nor U21853 (N_21853,N_21317,N_21467);
nor U21854 (N_21854,N_21507,N_21380);
nor U21855 (N_21855,N_21425,N_21569);
xnor U21856 (N_21856,N_21560,N_21443);
or U21857 (N_21857,N_21577,N_21336);
xnor U21858 (N_21858,N_21542,N_21310);
nand U21859 (N_21859,N_21555,N_21575);
nand U21860 (N_21860,N_21328,N_21450);
xor U21861 (N_21861,N_21349,N_21403);
nand U21862 (N_21862,N_21401,N_21502);
nand U21863 (N_21863,N_21525,N_21388);
nor U21864 (N_21864,N_21582,N_21489);
nor U21865 (N_21865,N_21306,N_21439);
nor U21866 (N_21866,N_21325,N_21597);
and U21867 (N_21867,N_21321,N_21426);
or U21868 (N_21868,N_21523,N_21336);
and U21869 (N_21869,N_21311,N_21525);
nor U21870 (N_21870,N_21432,N_21389);
nor U21871 (N_21871,N_21410,N_21407);
and U21872 (N_21872,N_21336,N_21375);
and U21873 (N_21873,N_21395,N_21433);
and U21874 (N_21874,N_21562,N_21441);
or U21875 (N_21875,N_21326,N_21462);
xnor U21876 (N_21876,N_21303,N_21413);
xor U21877 (N_21877,N_21421,N_21523);
nand U21878 (N_21878,N_21357,N_21419);
and U21879 (N_21879,N_21557,N_21549);
and U21880 (N_21880,N_21306,N_21414);
nand U21881 (N_21881,N_21363,N_21469);
nand U21882 (N_21882,N_21349,N_21437);
xnor U21883 (N_21883,N_21485,N_21536);
or U21884 (N_21884,N_21381,N_21473);
or U21885 (N_21885,N_21372,N_21465);
and U21886 (N_21886,N_21536,N_21554);
xnor U21887 (N_21887,N_21471,N_21339);
nor U21888 (N_21888,N_21406,N_21411);
nand U21889 (N_21889,N_21541,N_21426);
and U21890 (N_21890,N_21334,N_21397);
nor U21891 (N_21891,N_21335,N_21504);
or U21892 (N_21892,N_21519,N_21590);
nor U21893 (N_21893,N_21441,N_21311);
or U21894 (N_21894,N_21354,N_21310);
xor U21895 (N_21895,N_21480,N_21497);
xor U21896 (N_21896,N_21474,N_21584);
or U21897 (N_21897,N_21455,N_21568);
and U21898 (N_21898,N_21360,N_21353);
and U21899 (N_21899,N_21365,N_21554);
and U21900 (N_21900,N_21796,N_21860);
xor U21901 (N_21901,N_21638,N_21609);
nand U21902 (N_21902,N_21733,N_21771);
xor U21903 (N_21903,N_21842,N_21728);
nor U21904 (N_21904,N_21780,N_21741);
or U21905 (N_21905,N_21727,N_21642);
and U21906 (N_21906,N_21847,N_21615);
nand U21907 (N_21907,N_21817,N_21608);
or U21908 (N_21908,N_21677,N_21600);
nor U21909 (N_21909,N_21791,N_21603);
nor U21910 (N_21910,N_21878,N_21686);
and U21911 (N_21911,N_21678,N_21862);
nor U21912 (N_21912,N_21711,N_21648);
nand U21913 (N_21913,N_21782,N_21719);
nand U21914 (N_21914,N_21866,N_21879);
and U21915 (N_21915,N_21849,N_21655);
nand U21916 (N_21916,N_21896,N_21649);
and U21917 (N_21917,N_21641,N_21645);
nand U21918 (N_21918,N_21831,N_21852);
nand U21919 (N_21919,N_21848,N_21833);
nor U21920 (N_21920,N_21869,N_21807);
or U21921 (N_21921,N_21787,N_21809);
and U21922 (N_21922,N_21716,N_21836);
nor U21923 (N_21923,N_21701,N_21799);
xnor U21924 (N_21924,N_21626,N_21822);
nor U21925 (N_21925,N_21895,N_21762);
nor U21926 (N_21926,N_21816,N_21653);
or U21927 (N_21927,N_21758,N_21739);
or U21928 (N_21928,N_21684,N_21851);
nor U21929 (N_21929,N_21613,N_21802);
and U21930 (N_21930,N_21614,N_21611);
and U21931 (N_21931,N_21618,N_21650);
nor U21932 (N_21932,N_21874,N_21804);
xnor U21933 (N_21933,N_21743,N_21738);
and U21934 (N_21934,N_21685,N_21897);
or U21935 (N_21935,N_21661,N_21763);
or U21936 (N_21936,N_21721,N_21769);
xnor U21937 (N_21937,N_21681,N_21643);
and U21938 (N_21938,N_21752,N_21773);
nor U21939 (N_21939,N_21607,N_21774);
and U21940 (N_21940,N_21835,N_21764);
xnor U21941 (N_21941,N_21737,N_21759);
nor U21942 (N_21942,N_21644,N_21631);
or U21943 (N_21943,N_21620,N_21765);
nand U21944 (N_21944,N_21646,N_21659);
and U21945 (N_21945,N_21825,N_21781);
or U21946 (N_21946,N_21829,N_21656);
xnor U21947 (N_21947,N_21756,N_21899);
xor U21948 (N_21948,N_21875,N_21841);
xnor U21949 (N_21949,N_21725,N_21814);
nand U21950 (N_21950,N_21669,N_21663);
and U21951 (N_21951,N_21657,N_21637);
nand U21952 (N_21952,N_21894,N_21710);
xor U21953 (N_21953,N_21838,N_21694);
and U21954 (N_21954,N_21754,N_21667);
and U21955 (N_21955,N_21610,N_21888);
and U21956 (N_21956,N_21749,N_21766);
and U21957 (N_21957,N_21827,N_21867);
xor U21958 (N_21958,N_21664,N_21673);
and U21959 (N_21959,N_21772,N_21666);
nand U21960 (N_21960,N_21660,N_21709);
xor U21961 (N_21961,N_21883,N_21820);
nor U21962 (N_21962,N_21884,N_21806);
and U21963 (N_21963,N_21753,N_21813);
or U21964 (N_21964,N_21744,N_21689);
or U21965 (N_21965,N_21751,N_21794);
and U21966 (N_21966,N_21880,N_21887);
or U21967 (N_21967,N_21675,N_21882);
xnor U21968 (N_21968,N_21605,N_21691);
nand U21969 (N_21969,N_21635,N_21826);
or U21970 (N_21970,N_21837,N_21870);
nor U21971 (N_21971,N_21636,N_21602);
or U21972 (N_21972,N_21624,N_21778);
or U21973 (N_21973,N_21857,N_21606);
nor U21974 (N_21974,N_21750,N_21695);
and U21975 (N_21975,N_21844,N_21865);
nor U21976 (N_21976,N_21670,N_21748);
nand U21977 (N_21977,N_21877,N_21784);
nor U21978 (N_21978,N_21705,N_21617);
or U21979 (N_21979,N_21714,N_21858);
and U21980 (N_21980,N_21698,N_21793);
nand U21981 (N_21981,N_21770,N_21843);
nor U21982 (N_21982,N_21658,N_21652);
xor U21983 (N_21983,N_21651,N_21682);
and U21984 (N_21984,N_21604,N_21619);
xor U21985 (N_21985,N_21824,N_21706);
nand U21986 (N_21986,N_21881,N_21855);
or U21987 (N_21987,N_21742,N_21811);
nor U21988 (N_21988,N_21795,N_21768);
and U21989 (N_21989,N_21779,N_21789);
nand U21990 (N_21990,N_21747,N_21828);
and U21991 (N_21991,N_21845,N_21730);
nor U21992 (N_21992,N_21854,N_21783);
or U21993 (N_21993,N_21654,N_21693);
nor U21994 (N_21994,N_21680,N_21746);
xor U21995 (N_21995,N_21801,N_21785);
or U21996 (N_21996,N_21731,N_21699);
xor U21997 (N_21997,N_21622,N_21621);
xnor U21998 (N_21998,N_21776,N_21671);
nor U21999 (N_21999,N_21775,N_21616);
nand U22000 (N_22000,N_21839,N_21868);
and U22001 (N_22001,N_21672,N_21700);
nand U22002 (N_22002,N_21740,N_21832);
or U22003 (N_22003,N_21676,N_21729);
or U22004 (N_22004,N_21788,N_21859);
nand U22005 (N_22005,N_21668,N_21715);
nor U22006 (N_22006,N_21885,N_21856);
nor U22007 (N_22007,N_21818,N_21892);
nand U22008 (N_22008,N_21629,N_21732);
nor U22009 (N_22009,N_21761,N_21688);
or U22010 (N_22010,N_21679,N_21755);
xor U22011 (N_22011,N_21723,N_21601);
nor U22012 (N_22012,N_21718,N_21713);
and U22013 (N_22013,N_21726,N_21861);
nor U22014 (N_22014,N_21840,N_21639);
xnor U22015 (N_22015,N_21808,N_21815);
and U22016 (N_22016,N_21893,N_21760);
xnor U22017 (N_22017,N_21690,N_21708);
nor U22018 (N_22018,N_21797,N_21798);
nor U22019 (N_22019,N_21876,N_21623);
and U22020 (N_22020,N_21792,N_21786);
nand U22021 (N_22021,N_21805,N_21735);
or U22022 (N_22022,N_21830,N_21630);
nand U22023 (N_22023,N_21665,N_21898);
nor U22024 (N_22024,N_21800,N_21819);
and U22025 (N_22025,N_21890,N_21717);
or U22026 (N_22026,N_21628,N_21702);
xnor U22027 (N_22027,N_21712,N_21757);
xor U22028 (N_22028,N_21707,N_21886);
nand U22029 (N_22029,N_21625,N_21872);
nor U22030 (N_22030,N_21889,N_21627);
nand U22031 (N_22031,N_21734,N_21803);
or U22032 (N_22032,N_21846,N_21634);
nand U22033 (N_22033,N_21687,N_21722);
xnor U22034 (N_22034,N_21871,N_21863);
nand U22035 (N_22035,N_21703,N_21683);
xnor U22036 (N_22036,N_21873,N_21834);
nand U22037 (N_22037,N_21720,N_21674);
nor U22038 (N_22038,N_21853,N_21821);
nand U22039 (N_22039,N_21724,N_21810);
and U22040 (N_22040,N_21704,N_21891);
and U22041 (N_22041,N_21745,N_21692);
nand U22042 (N_22042,N_21697,N_21633);
nor U22043 (N_22043,N_21736,N_21612);
or U22044 (N_22044,N_21767,N_21640);
or U22045 (N_22045,N_21696,N_21850);
nor U22046 (N_22046,N_21812,N_21632);
or U22047 (N_22047,N_21647,N_21864);
nor U22048 (N_22048,N_21777,N_21662);
and U22049 (N_22049,N_21790,N_21823);
xnor U22050 (N_22050,N_21647,N_21790);
and U22051 (N_22051,N_21633,N_21622);
xor U22052 (N_22052,N_21841,N_21857);
or U22053 (N_22053,N_21665,N_21714);
xor U22054 (N_22054,N_21743,N_21797);
nand U22055 (N_22055,N_21713,N_21624);
and U22056 (N_22056,N_21644,N_21699);
xnor U22057 (N_22057,N_21776,N_21716);
and U22058 (N_22058,N_21846,N_21643);
nand U22059 (N_22059,N_21643,N_21741);
nand U22060 (N_22060,N_21719,N_21706);
or U22061 (N_22061,N_21851,N_21795);
and U22062 (N_22062,N_21842,N_21724);
nand U22063 (N_22063,N_21713,N_21652);
nor U22064 (N_22064,N_21671,N_21833);
xnor U22065 (N_22065,N_21661,N_21665);
nor U22066 (N_22066,N_21651,N_21692);
nand U22067 (N_22067,N_21842,N_21798);
and U22068 (N_22068,N_21671,N_21855);
nor U22069 (N_22069,N_21843,N_21762);
nor U22070 (N_22070,N_21859,N_21627);
and U22071 (N_22071,N_21887,N_21676);
nand U22072 (N_22072,N_21781,N_21759);
nand U22073 (N_22073,N_21762,N_21860);
xnor U22074 (N_22074,N_21849,N_21666);
xnor U22075 (N_22075,N_21669,N_21861);
nor U22076 (N_22076,N_21641,N_21617);
nor U22077 (N_22077,N_21668,N_21760);
nand U22078 (N_22078,N_21671,N_21755);
nand U22079 (N_22079,N_21894,N_21722);
nand U22080 (N_22080,N_21864,N_21680);
nor U22081 (N_22081,N_21638,N_21775);
nand U22082 (N_22082,N_21804,N_21849);
xor U22083 (N_22083,N_21691,N_21659);
and U22084 (N_22084,N_21690,N_21843);
and U22085 (N_22085,N_21814,N_21657);
and U22086 (N_22086,N_21785,N_21874);
nand U22087 (N_22087,N_21757,N_21649);
nand U22088 (N_22088,N_21629,N_21780);
nor U22089 (N_22089,N_21695,N_21674);
nor U22090 (N_22090,N_21823,N_21760);
and U22091 (N_22091,N_21779,N_21745);
xor U22092 (N_22092,N_21833,N_21636);
nand U22093 (N_22093,N_21786,N_21808);
and U22094 (N_22094,N_21773,N_21674);
xor U22095 (N_22095,N_21655,N_21678);
xor U22096 (N_22096,N_21789,N_21619);
nor U22097 (N_22097,N_21644,N_21657);
nand U22098 (N_22098,N_21630,N_21869);
nor U22099 (N_22099,N_21615,N_21713);
nand U22100 (N_22100,N_21864,N_21851);
nor U22101 (N_22101,N_21810,N_21631);
and U22102 (N_22102,N_21891,N_21794);
nor U22103 (N_22103,N_21826,N_21728);
or U22104 (N_22104,N_21666,N_21846);
nand U22105 (N_22105,N_21786,N_21700);
xor U22106 (N_22106,N_21875,N_21717);
and U22107 (N_22107,N_21786,N_21788);
and U22108 (N_22108,N_21854,N_21837);
xnor U22109 (N_22109,N_21695,N_21740);
nor U22110 (N_22110,N_21698,N_21622);
or U22111 (N_22111,N_21773,N_21790);
xnor U22112 (N_22112,N_21833,N_21633);
nor U22113 (N_22113,N_21758,N_21852);
or U22114 (N_22114,N_21747,N_21883);
and U22115 (N_22115,N_21606,N_21814);
or U22116 (N_22116,N_21656,N_21713);
or U22117 (N_22117,N_21794,N_21843);
xor U22118 (N_22118,N_21725,N_21811);
xnor U22119 (N_22119,N_21706,N_21895);
nor U22120 (N_22120,N_21850,N_21806);
or U22121 (N_22121,N_21713,N_21709);
xor U22122 (N_22122,N_21687,N_21855);
and U22123 (N_22123,N_21718,N_21647);
xnor U22124 (N_22124,N_21722,N_21724);
nand U22125 (N_22125,N_21858,N_21806);
nor U22126 (N_22126,N_21637,N_21848);
or U22127 (N_22127,N_21656,N_21668);
and U22128 (N_22128,N_21761,N_21605);
nand U22129 (N_22129,N_21724,N_21723);
or U22130 (N_22130,N_21884,N_21852);
nor U22131 (N_22131,N_21744,N_21872);
nand U22132 (N_22132,N_21888,N_21631);
nor U22133 (N_22133,N_21737,N_21868);
xnor U22134 (N_22134,N_21779,N_21710);
or U22135 (N_22135,N_21691,N_21888);
or U22136 (N_22136,N_21668,N_21884);
or U22137 (N_22137,N_21654,N_21747);
xor U22138 (N_22138,N_21756,N_21613);
or U22139 (N_22139,N_21743,N_21811);
or U22140 (N_22140,N_21782,N_21629);
nor U22141 (N_22141,N_21630,N_21718);
nor U22142 (N_22142,N_21866,N_21701);
nor U22143 (N_22143,N_21668,N_21683);
nand U22144 (N_22144,N_21698,N_21794);
nor U22145 (N_22145,N_21674,N_21721);
or U22146 (N_22146,N_21844,N_21605);
or U22147 (N_22147,N_21668,N_21738);
nor U22148 (N_22148,N_21717,N_21705);
and U22149 (N_22149,N_21819,N_21602);
and U22150 (N_22150,N_21880,N_21600);
nand U22151 (N_22151,N_21727,N_21725);
nand U22152 (N_22152,N_21637,N_21787);
or U22153 (N_22153,N_21713,N_21884);
xnor U22154 (N_22154,N_21765,N_21894);
and U22155 (N_22155,N_21775,N_21889);
nand U22156 (N_22156,N_21783,N_21632);
xnor U22157 (N_22157,N_21701,N_21643);
nand U22158 (N_22158,N_21619,N_21874);
nor U22159 (N_22159,N_21669,N_21851);
xnor U22160 (N_22160,N_21805,N_21730);
and U22161 (N_22161,N_21815,N_21746);
xnor U22162 (N_22162,N_21691,N_21896);
xnor U22163 (N_22163,N_21804,N_21637);
nand U22164 (N_22164,N_21618,N_21672);
and U22165 (N_22165,N_21844,N_21613);
nor U22166 (N_22166,N_21677,N_21662);
nor U22167 (N_22167,N_21710,N_21658);
or U22168 (N_22168,N_21844,N_21654);
nor U22169 (N_22169,N_21837,N_21629);
or U22170 (N_22170,N_21838,N_21606);
or U22171 (N_22171,N_21762,N_21685);
or U22172 (N_22172,N_21695,N_21793);
nand U22173 (N_22173,N_21652,N_21773);
or U22174 (N_22174,N_21899,N_21698);
and U22175 (N_22175,N_21753,N_21884);
nand U22176 (N_22176,N_21616,N_21733);
or U22177 (N_22177,N_21862,N_21666);
nand U22178 (N_22178,N_21884,N_21748);
nand U22179 (N_22179,N_21745,N_21740);
or U22180 (N_22180,N_21730,N_21800);
nand U22181 (N_22181,N_21802,N_21805);
and U22182 (N_22182,N_21655,N_21870);
xnor U22183 (N_22183,N_21600,N_21851);
nor U22184 (N_22184,N_21645,N_21866);
xnor U22185 (N_22185,N_21688,N_21704);
or U22186 (N_22186,N_21715,N_21633);
nor U22187 (N_22187,N_21707,N_21754);
or U22188 (N_22188,N_21649,N_21762);
and U22189 (N_22189,N_21666,N_21842);
xnor U22190 (N_22190,N_21642,N_21647);
nor U22191 (N_22191,N_21856,N_21742);
and U22192 (N_22192,N_21619,N_21768);
and U22193 (N_22193,N_21820,N_21683);
nor U22194 (N_22194,N_21872,N_21887);
and U22195 (N_22195,N_21631,N_21710);
nor U22196 (N_22196,N_21808,N_21895);
nand U22197 (N_22197,N_21727,N_21647);
xor U22198 (N_22198,N_21876,N_21712);
nor U22199 (N_22199,N_21676,N_21693);
and U22200 (N_22200,N_22179,N_22188);
or U22201 (N_22201,N_22024,N_22084);
xnor U22202 (N_22202,N_21933,N_21919);
or U22203 (N_22203,N_21926,N_22071);
xnor U22204 (N_22204,N_21987,N_22182);
xor U22205 (N_22205,N_22064,N_21930);
and U22206 (N_22206,N_22055,N_22126);
nand U22207 (N_22207,N_21931,N_21904);
nor U22208 (N_22208,N_22073,N_22120);
xnor U22209 (N_22209,N_22093,N_22173);
nand U22210 (N_22210,N_22152,N_22144);
nor U22211 (N_22211,N_21922,N_22147);
nand U22212 (N_22212,N_21984,N_22197);
and U22213 (N_22213,N_21932,N_22072);
nand U22214 (N_22214,N_22165,N_22170);
nand U22215 (N_22215,N_21953,N_21927);
nor U22216 (N_22216,N_22074,N_22159);
xor U22217 (N_22217,N_22135,N_22088);
nand U22218 (N_22218,N_21972,N_22061);
and U22219 (N_22219,N_22114,N_22008);
nor U22220 (N_22220,N_21974,N_22195);
nor U22221 (N_22221,N_22062,N_22103);
nor U22222 (N_22222,N_22017,N_22151);
or U22223 (N_22223,N_22056,N_22112);
nand U22224 (N_22224,N_21925,N_22106);
xnor U22225 (N_22225,N_22022,N_21979);
and U22226 (N_22226,N_21910,N_22154);
nor U22227 (N_22227,N_22115,N_22164);
and U22228 (N_22228,N_21907,N_22142);
or U22229 (N_22229,N_22044,N_22092);
nand U22230 (N_22230,N_22030,N_22014);
or U22231 (N_22231,N_22079,N_21939);
nand U22232 (N_22232,N_22032,N_22052);
xnor U22233 (N_22233,N_22155,N_22026);
nor U22234 (N_22234,N_21971,N_21911);
xor U22235 (N_22235,N_22053,N_21999);
xor U22236 (N_22236,N_22190,N_22192);
nand U22237 (N_22237,N_22015,N_21952);
nor U22238 (N_22238,N_22162,N_22133);
xor U22239 (N_22239,N_22117,N_21900);
xnor U22240 (N_22240,N_22012,N_22006);
and U22241 (N_22241,N_22123,N_22127);
nor U22242 (N_22242,N_22002,N_21929);
nand U22243 (N_22243,N_21981,N_21975);
nor U22244 (N_22244,N_21909,N_22047);
nor U22245 (N_22245,N_22175,N_22167);
nor U22246 (N_22246,N_22119,N_22045);
or U22247 (N_22247,N_22153,N_22004);
xor U22248 (N_22248,N_22134,N_21982);
and U22249 (N_22249,N_22187,N_22196);
or U22250 (N_22250,N_22007,N_22057);
nand U22251 (N_22251,N_22149,N_21958);
or U22252 (N_22252,N_21954,N_22086);
nor U22253 (N_22253,N_21948,N_21912);
nand U22254 (N_22254,N_21998,N_22099);
and U22255 (N_22255,N_21980,N_22011);
and U22256 (N_22256,N_21943,N_21915);
or U22257 (N_22257,N_21951,N_22129);
nand U22258 (N_22258,N_22068,N_22122);
nor U22259 (N_22259,N_21965,N_21937);
xnor U22260 (N_22260,N_22128,N_21983);
nand U22261 (N_22261,N_21989,N_22183);
nor U22262 (N_22262,N_22090,N_22033);
or U22263 (N_22263,N_21905,N_22043);
xnor U22264 (N_22264,N_22036,N_22040);
xor U22265 (N_22265,N_22029,N_22141);
nor U22266 (N_22266,N_21938,N_21977);
and U22267 (N_22267,N_21985,N_21923);
xnor U22268 (N_22268,N_22186,N_22146);
or U22269 (N_22269,N_22027,N_22091);
or U22270 (N_22270,N_22009,N_22003);
nor U22271 (N_22271,N_22189,N_22077);
and U22272 (N_22272,N_21957,N_22070);
xnor U22273 (N_22273,N_22028,N_22160);
xor U22274 (N_22274,N_21959,N_22176);
or U22275 (N_22275,N_21906,N_22100);
nor U22276 (N_22276,N_22080,N_22016);
xnor U22277 (N_22277,N_21973,N_21993);
nor U22278 (N_22278,N_22124,N_22191);
xnor U22279 (N_22279,N_22021,N_22156);
xor U22280 (N_22280,N_22050,N_21936);
nor U22281 (N_22281,N_22082,N_21963);
and U22282 (N_22282,N_22038,N_22095);
nand U22283 (N_22283,N_22000,N_21916);
nor U22284 (N_22284,N_22125,N_21961);
nand U22285 (N_22285,N_22018,N_22069);
nand U22286 (N_22286,N_21902,N_22181);
nand U22287 (N_22287,N_22054,N_22121);
and U22288 (N_22288,N_22098,N_21913);
nand U22289 (N_22289,N_22136,N_22194);
xor U22290 (N_22290,N_22039,N_22111);
or U22291 (N_22291,N_22148,N_22174);
nand U22292 (N_22292,N_22116,N_22118);
and U22293 (N_22293,N_22065,N_21924);
nor U22294 (N_22294,N_22101,N_21944);
nand U22295 (N_22295,N_22169,N_21967);
or U22296 (N_22296,N_21914,N_22198);
or U22297 (N_22297,N_22042,N_21908);
xor U22298 (N_22298,N_22051,N_22087);
and U22299 (N_22299,N_22166,N_22059);
or U22300 (N_22300,N_22178,N_21968);
nor U22301 (N_22301,N_22137,N_22102);
nor U22302 (N_22302,N_22107,N_22089);
nand U22303 (N_22303,N_21945,N_22048);
and U22304 (N_22304,N_22110,N_22096);
or U22305 (N_22305,N_22143,N_21995);
or U22306 (N_22306,N_21960,N_22037);
nor U22307 (N_22307,N_22013,N_22105);
nand U22308 (N_22308,N_21947,N_22060);
nand U22309 (N_22309,N_22049,N_21956);
xor U22310 (N_22310,N_22031,N_21942);
and U22311 (N_22311,N_22010,N_22177);
nand U22312 (N_22312,N_21941,N_22019);
nand U22313 (N_22313,N_22108,N_22058);
nand U22314 (N_22314,N_22076,N_21997);
and U22315 (N_22315,N_22023,N_22078);
or U22316 (N_22316,N_22168,N_21921);
xor U22317 (N_22317,N_21978,N_21986);
or U22318 (N_22318,N_21955,N_21917);
nor U22319 (N_22319,N_22140,N_22131);
nor U22320 (N_22320,N_22138,N_21903);
xnor U22321 (N_22321,N_22180,N_22066);
nand U22322 (N_22322,N_22193,N_22139);
xor U22323 (N_22323,N_21918,N_22157);
or U22324 (N_22324,N_21934,N_21949);
nand U22325 (N_22325,N_22104,N_21901);
or U22326 (N_22326,N_22085,N_21946);
or U22327 (N_22327,N_21964,N_22067);
nand U22328 (N_22328,N_22109,N_22163);
nor U22329 (N_22329,N_22161,N_22075);
nor U22330 (N_22330,N_22041,N_21996);
xnor U22331 (N_22331,N_21966,N_21950);
and U22332 (N_22332,N_22025,N_21994);
xnor U22333 (N_22333,N_21988,N_22020);
xor U22334 (N_22334,N_22094,N_22130);
xor U22335 (N_22335,N_21970,N_22001);
and U22336 (N_22336,N_22132,N_22046);
nor U22337 (N_22337,N_21928,N_21990);
nand U22338 (N_22338,N_22005,N_21991);
nor U22339 (N_22339,N_22199,N_22063);
or U22340 (N_22340,N_21920,N_21962);
xor U22341 (N_22341,N_22185,N_22150);
or U22342 (N_22342,N_22184,N_22097);
nor U22343 (N_22343,N_22034,N_22158);
and U22344 (N_22344,N_21969,N_22035);
nand U22345 (N_22345,N_22081,N_22113);
and U22346 (N_22346,N_21992,N_21976);
nand U22347 (N_22347,N_22171,N_21935);
xnor U22348 (N_22348,N_22145,N_22083);
or U22349 (N_22349,N_22172,N_21940);
xor U22350 (N_22350,N_21989,N_22145);
and U22351 (N_22351,N_22028,N_21958);
and U22352 (N_22352,N_22152,N_22171);
xnor U22353 (N_22353,N_22173,N_22070);
nor U22354 (N_22354,N_21923,N_22046);
and U22355 (N_22355,N_22123,N_22111);
nor U22356 (N_22356,N_22157,N_21969);
xor U22357 (N_22357,N_21979,N_22143);
xnor U22358 (N_22358,N_21926,N_21945);
or U22359 (N_22359,N_21960,N_21994);
or U22360 (N_22360,N_22159,N_21999);
nor U22361 (N_22361,N_21979,N_22127);
and U22362 (N_22362,N_22093,N_22083);
xnor U22363 (N_22363,N_22088,N_22148);
or U22364 (N_22364,N_22093,N_22023);
xnor U22365 (N_22365,N_21903,N_21935);
nor U22366 (N_22366,N_22109,N_22130);
nand U22367 (N_22367,N_21950,N_22020);
nor U22368 (N_22368,N_21981,N_22159);
xor U22369 (N_22369,N_21917,N_21913);
nor U22370 (N_22370,N_22004,N_21961);
nand U22371 (N_22371,N_22007,N_22073);
nor U22372 (N_22372,N_21935,N_22161);
xor U22373 (N_22373,N_22161,N_22186);
and U22374 (N_22374,N_22039,N_22043);
and U22375 (N_22375,N_22162,N_22059);
xor U22376 (N_22376,N_22140,N_21981);
or U22377 (N_22377,N_22136,N_22052);
nand U22378 (N_22378,N_22177,N_22098);
nor U22379 (N_22379,N_21961,N_22118);
nor U22380 (N_22380,N_22152,N_22128);
nand U22381 (N_22381,N_21958,N_21988);
or U22382 (N_22382,N_21986,N_22169);
nand U22383 (N_22383,N_22072,N_21906);
or U22384 (N_22384,N_22143,N_22052);
nand U22385 (N_22385,N_22076,N_22083);
xnor U22386 (N_22386,N_22142,N_22082);
and U22387 (N_22387,N_22149,N_21944);
nand U22388 (N_22388,N_22121,N_22068);
or U22389 (N_22389,N_22085,N_22108);
xor U22390 (N_22390,N_22123,N_22178);
nand U22391 (N_22391,N_22125,N_22164);
nand U22392 (N_22392,N_22051,N_22194);
nand U22393 (N_22393,N_22012,N_21962);
xnor U22394 (N_22394,N_21924,N_22012);
nand U22395 (N_22395,N_21986,N_22000);
or U22396 (N_22396,N_21981,N_21962);
xnor U22397 (N_22397,N_21924,N_22061);
and U22398 (N_22398,N_22144,N_22064);
or U22399 (N_22399,N_22070,N_22014);
nor U22400 (N_22400,N_22187,N_22096);
xnor U22401 (N_22401,N_22000,N_22158);
and U22402 (N_22402,N_21972,N_22125);
xnor U22403 (N_22403,N_22141,N_22140);
xor U22404 (N_22404,N_21916,N_22104);
nor U22405 (N_22405,N_22050,N_22081);
nand U22406 (N_22406,N_21994,N_22028);
nor U22407 (N_22407,N_21941,N_21914);
nand U22408 (N_22408,N_21960,N_22130);
xnor U22409 (N_22409,N_22092,N_22095);
nand U22410 (N_22410,N_21952,N_21917);
xnor U22411 (N_22411,N_22199,N_22185);
nand U22412 (N_22412,N_21990,N_22081);
nor U22413 (N_22413,N_22078,N_22194);
xor U22414 (N_22414,N_21941,N_22036);
and U22415 (N_22415,N_22179,N_22062);
xnor U22416 (N_22416,N_21929,N_22018);
nor U22417 (N_22417,N_22190,N_22032);
nor U22418 (N_22418,N_22055,N_22170);
nor U22419 (N_22419,N_22135,N_22093);
nand U22420 (N_22420,N_21971,N_22010);
nor U22421 (N_22421,N_21968,N_21975);
nor U22422 (N_22422,N_22172,N_22190);
nand U22423 (N_22423,N_21915,N_22188);
and U22424 (N_22424,N_22023,N_22055);
xnor U22425 (N_22425,N_22126,N_22024);
nand U22426 (N_22426,N_22176,N_21967);
nand U22427 (N_22427,N_21907,N_22192);
or U22428 (N_22428,N_21998,N_21900);
and U22429 (N_22429,N_22074,N_21976);
nor U22430 (N_22430,N_22045,N_21945);
nand U22431 (N_22431,N_22009,N_21998);
and U22432 (N_22432,N_21900,N_22111);
or U22433 (N_22433,N_22106,N_22198);
nand U22434 (N_22434,N_21990,N_22102);
xnor U22435 (N_22435,N_22190,N_21916);
and U22436 (N_22436,N_22189,N_22033);
nor U22437 (N_22437,N_22097,N_21979);
or U22438 (N_22438,N_22046,N_21990);
nand U22439 (N_22439,N_21982,N_21957);
xnor U22440 (N_22440,N_22054,N_22099);
nor U22441 (N_22441,N_22006,N_22072);
nor U22442 (N_22442,N_22158,N_22070);
and U22443 (N_22443,N_22119,N_22139);
nand U22444 (N_22444,N_22192,N_21996);
and U22445 (N_22445,N_21938,N_22071);
xor U22446 (N_22446,N_22022,N_22083);
and U22447 (N_22447,N_22098,N_21916);
and U22448 (N_22448,N_21906,N_22090);
nor U22449 (N_22449,N_22033,N_22065);
nand U22450 (N_22450,N_21929,N_21966);
or U22451 (N_22451,N_22122,N_21915);
or U22452 (N_22452,N_22169,N_22116);
xnor U22453 (N_22453,N_22183,N_22109);
nor U22454 (N_22454,N_22169,N_22129);
and U22455 (N_22455,N_22029,N_21918);
nand U22456 (N_22456,N_22145,N_21987);
nand U22457 (N_22457,N_22104,N_21930);
and U22458 (N_22458,N_22110,N_22151);
and U22459 (N_22459,N_22179,N_21910);
and U22460 (N_22460,N_22093,N_21965);
and U22461 (N_22461,N_22176,N_21940);
or U22462 (N_22462,N_22044,N_21998);
nor U22463 (N_22463,N_22039,N_22134);
nor U22464 (N_22464,N_21945,N_21940);
xor U22465 (N_22465,N_22138,N_21957);
xor U22466 (N_22466,N_22120,N_22105);
nand U22467 (N_22467,N_21952,N_22069);
nor U22468 (N_22468,N_21915,N_22131);
nand U22469 (N_22469,N_21994,N_22194);
or U22470 (N_22470,N_22106,N_22014);
or U22471 (N_22471,N_22041,N_22053);
nor U22472 (N_22472,N_22149,N_21970);
or U22473 (N_22473,N_22188,N_22003);
and U22474 (N_22474,N_21927,N_22026);
nand U22475 (N_22475,N_22101,N_22190);
or U22476 (N_22476,N_21984,N_21945);
xor U22477 (N_22477,N_21977,N_21974);
and U22478 (N_22478,N_22158,N_22020);
and U22479 (N_22479,N_22020,N_21955);
and U22480 (N_22480,N_21984,N_22121);
and U22481 (N_22481,N_22157,N_22119);
or U22482 (N_22482,N_22062,N_22034);
nor U22483 (N_22483,N_21961,N_22055);
xor U22484 (N_22484,N_22066,N_22140);
xor U22485 (N_22485,N_22138,N_22196);
or U22486 (N_22486,N_22144,N_21940);
nand U22487 (N_22487,N_22079,N_22147);
nand U22488 (N_22488,N_21902,N_22053);
xor U22489 (N_22489,N_22015,N_21995);
or U22490 (N_22490,N_22026,N_21903);
xor U22491 (N_22491,N_22177,N_22093);
nor U22492 (N_22492,N_22127,N_21908);
nor U22493 (N_22493,N_22015,N_21988);
or U22494 (N_22494,N_22011,N_21929);
xor U22495 (N_22495,N_22106,N_21987);
xnor U22496 (N_22496,N_22171,N_22055);
xor U22497 (N_22497,N_22006,N_22134);
nor U22498 (N_22498,N_22040,N_22142);
and U22499 (N_22499,N_21996,N_21942);
or U22500 (N_22500,N_22442,N_22201);
or U22501 (N_22501,N_22317,N_22335);
nor U22502 (N_22502,N_22203,N_22233);
or U22503 (N_22503,N_22347,N_22221);
nor U22504 (N_22504,N_22300,N_22456);
xor U22505 (N_22505,N_22436,N_22467);
xor U22506 (N_22506,N_22338,N_22278);
and U22507 (N_22507,N_22396,N_22411);
nor U22508 (N_22508,N_22390,N_22357);
nor U22509 (N_22509,N_22315,N_22471);
nor U22510 (N_22510,N_22325,N_22382);
nor U22511 (N_22511,N_22407,N_22206);
nor U22512 (N_22512,N_22298,N_22288);
nor U22513 (N_22513,N_22336,N_22324);
nand U22514 (N_22514,N_22220,N_22277);
or U22515 (N_22515,N_22341,N_22214);
nand U22516 (N_22516,N_22469,N_22374);
and U22517 (N_22517,N_22303,N_22497);
and U22518 (N_22518,N_22440,N_22474);
xor U22519 (N_22519,N_22496,N_22438);
or U22520 (N_22520,N_22406,N_22398);
and U22521 (N_22521,N_22250,N_22448);
nand U22522 (N_22522,N_22275,N_22416);
xor U22523 (N_22523,N_22358,N_22413);
or U22524 (N_22524,N_22232,N_22356);
or U22525 (N_22525,N_22224,N_22421);
nand U22526 (N_22526,N_22395,N_22366);
or U22527 (N_22527,N_22238,N_22423);
or U22528 (N_22528,N_22443,N_22302);
xor U22529 (N_22529,N_22241,N_22293);
nor U22530 (N_22530,N_22375,N_22237);
xnor U22531 (N_22531,N_22263,N_22260);
nand U22532 (N_22532,N_22269,N_22309);
or U22533 (N_22533,N_22249,N_22242);
xnor U22534 (N_22534,N_22267,N_22428);
and U22535 (N_22535,N_22222,N_22259);
nor U22536 (N_22536,N_22449,N_22344);
xor U22537 (N_22537,N_22240,N_22393);
nor U22538 (N_22538,N_22454,N_22257);
and U22539 (N_22539,N_22297,N_22294);
and U22540 (N_22540,N_22280,N_22472);
and U22541 (N_22541,N_22330,N_22494);
and U22542 (N_22542,N_22306,N_22296);
xnor U22543 (N_22543,N_22468,N_22234);
xnor U22544 (N_22544,N_22386,N_22482);
nor U22545 (N_22545,N_22483,N_22248);
nor U22546 (N_22546,N_22384,N_22349);
xor U22547 (N_22547,N_22350,N_22400);
nand U22548 (N_22548,N_22217,N_22245);
or U22549 (N_22549,N_22334,N_22289);
or U22550 (N_22550,N_22422,N_22353);
xnor U22551 (N_22551,N_22337,N_22210);
or U22552 (N_22552,N_22355,N_22343);
and U22553 (N_22553,N_22307,N_22333);
nand U22554 (N_22554,N_22464,N_22476);
and U22555 (N_22555,N_22435,N_22273);
and U22556 (N_22556,N_22322,N_22447);
or U22557 (N_22557,N_22418,N_22320);
xnor U22558 (N_22558,N_22256,N_22433);
xor U22559 (N_22559,N_22485,N_22208);
or U22560 (N_22560,N_22488,N_22419);
or U22561 (N_22561,N_22254,N_22424);
and U22562 (N_22562,N_22463,N_22265);
and U22563 (N_22563,N_22239,N_22215);
nand U22564 (N_22564,N_22364,N_22351);
or U22565 (N_22565,N_22229,N_22342);
nand U22566 (N_22566,N_22498,N_22369);
or U22567 (N_22567,N_22445,N_22481);
and U22568 (N_22568,N_22420,N_22432);
and U22569 (N_22569,N_22427,N_22409);
and U22570 (N_22570,N_22453,N_22284);
nor U22571 (N_22571,N_22270,N_22410);
and U22572 (N_22572,N_22332,N_22415);
nand U22573 (N_22573,N_22389,N_22323);
nand U22574 (N_22574,N_22354,N_22276);
or U22575 (N_22575,N_22262,N_22408);
xor U22576 (N_22576,N_22328,N_22499);
or U22577 (N_22577,N_22441,N_22253);
nor U22578 (N_22578,N_22279,N_22271);
and U22579 (N_22579,N_22491,N_22379);
and U22580 (N_22580,N_22377,N_22236);
xnor U22581 (N_22581,N_22360,N_22425);
nand U22582 (N_22582,N_22200,N_22230);
xor U22583 (N_22583,N_22402,N_22479);
nand U22584 (N_22584,N_22255,N_22380);
nor U22585 (N_22585,N_22295,N_22429);
xor U22586 (N_22586,N_22216,N_22414);
nor U22587 (N_22587,N_22391,N_22223);
or U22588 (N_22588,N_22251,N_22339);
xor U22589 (N_22589,N_22412,N_22202);
nor U22590 (N_22590,N_22281,N_22444);
and U22591 (N_22591,N_22478,N_22345);
or U22592 (N_22592,N_22305,N_22274);
xor U22593 (N_22593,N_22458,N_22460);
and U22594 (N_22594,N_22348,N_22247);
xnor U22595 (N_22595,N_22213,N_22401);
xnor U22596 (N_22596,N_22363,N_22286);
and U22597 (N_22597,N_22211,N_22312);
xnor U22598 (N_22598,N_22327,N_22283);
and U22599 (N_22599,N_22475,N_22462);
and U22600 (N_22600,N_22207,N_22218);
and U22601 (N_22601,N_22311,N_22272);
nor U22602 (N_22602,N_22266,N_22227);
nor U22603 (N_22603,N_22461,N_22431);
or U22604 (N_22604,N_22319,N_22361);
xor U22605 (N_22605,N_22403,N_22466);
and U22606 (N_22606,N_22235,N_22313);
or U22607 (N_22607,N_22326,N_22434);
or U22608 (N_22608,N_22484,N_22290);
and U22609 (N_22609,N_22437,N_22314);
and U22610 (N_22610,N_22291,N_22261);
xnor U22611 (N_22611,N_22228,N_22209);
xnor U22612 (N_22612,N_22219,N_22470);
nand U22613 (N_22613,N_22205,N_22490);
and U22614 (N_22614,N_22489,N_22310);
xnor U22615 (N_22615,N_22362,N_22459);
nor U22616 (N_22616,N_22455,N_22321);
nor U22617 (N_22617,N_22473,N_22225);
and U22618 (N_22618,N_22397,N_22367);
nor U22619 (N_22619,N_22299,N_22495);
nor U22620 (N_22620,N_22352,N_22226);
nor U22621 (N_22621,N_22388,N_22264);
nand U22622 (N_22622,N_22308,N_22246);
nand U22623 (N_22623,N_22292,N_22426);
nand U22624 (N_22624,N_22331,N_22450);
nand U22625 (N_22625,N_22282,N_22477);
nand U22626 (N_22626,N_22370,N_22457);
xor U22627 (N_22627,N_22394,N_22439);
nor U22628 (N_22628,N_22381,N_22365);
xor U22629 (N_22629,N_22204,N_22417);
xnor U22630 (N_22630,N_22383,N_22492);
and U22631 (N_22631,N_22285,N_22404);
and U22632 (N_22632,N_22244,N_22212);
nand U22633 (N_22633,N_22451,N_22318);
nor U22634 (N_22634,N_22493,N_22430);
xor U22635 (N_22635,N_22392,N_22399);
xnor U22636 (N_22636,N_22231,N_22243);
nand U22637 (N_22637,N_22465,N_22373);
nand U22638 (N_22638,N_22405,N_22376);
nand U22639 (N_22639,N_22378,N_22329);
or U22640 (N_22640,N_22340,N_22372);
or U22641 (N_22641,N_22359,N_22385);
and U22642 (N_22642,N_22387,N_22252);
nor U22643 (N_22643,N_22287,N_22316);
xnor U22644 (N_22644,N_22371,N_22346);
xor U22645 (N_22645,N_22487,N_22446);
or U22646 (N_22646,N_22301,N_22486);
xnor U22647 (N_22647,N_22268,N_22258);
and U22648 (N_22648,N_22452,N_22480);
or U22649 (N_22649,N_22304,N_22368);
nand U22650 (N_22650,N_22443,N_22448);
nor U22651 (N_22651,N_22414,N_22345);
nor U22652 (N_22652,N_22427,N_22469);
nand U22653 (N_22653,N_22224,N_22360);
xnor U22654 (N_22654,N_22472,N_22438);
nand U22655 (N_22655,N_22231,N_22359);
nor U22656 (N_22656,N_22295,N_22320);
and U22657 (N_22657,N_22451,N_22292);
nand U22658 (N_22658,N_22385,N_22261);
and U22659 (N_22659,N_22348,N_22340);
nand U22660 (N_22660,N_22258,N_22359);
xnor U22661 (N_22661,N_22234,N_22348);
nor U22662 (N_22662,N_22341,N_22471);
xnor U22663 (N_22663,N_22443,N_22493);
nand U22664 (N_22664,N_22211,N_22237);
xnor U22665 (N_22665,N_22283,N_22487);
nor U22666 (N_22666,N_22332,N_22392);
nor U22667 (N_22667,N_22323,N_22393);
or U22668 (N_22668,N_22289,N_22389);
xnor U22669 (N_22669,N_22233,N_22369);
nor U22670 (N_22670,N_22229,N_22320);
nor U22671 (N_22671,N_22450,N_22342);
xor U22672 (N_22672,N_22358,N_22429);
xor U22673 (N_22673,N_22315,N_22307);
and U22674 (N_22674,N_22304,N_22343);
nor U22675 (N_22675,N_22264,N_22428);
nor U22676 (N_22676,N_22355,N_22426);
nand U22677 (N_22677,N_22236,N_22340);
xnor U22678 (N_22678,N_22317,N_22355);
and U22679 (N_22679,N_22217,N_22253);
nor U22680 (N_22680,N_22203,N_22355);
or U22681 (N_22681,N_22202,N_22288);
nand U22682 (N_22682,N_22493,N_22349);
nand U22683 (N_22683,N_22204,N_22329);
nand U22684 (N_22684,N_22312,N_22495);
xnor U22685 (N_22685,N_22335,N_22405);
and U22686 (N_22686,N_22460,N_22362);
xor U22687 (N_22687,N_22297,N_22447);
or U22688 (N_22688,N_22330,N_22282);
nor U22689 (N_22689,N_22253,N_22367);
nor U22690 (N_22690,N_22470,N_22421);
or U22691 (N_22691,N_22416,N_22293);
and U22692 (N_22692,N_22226,N_22460);
xnor U22693 (N_22693,N_22403,N_22404);
and U22694 (N_22694,N_22373,N_22440);
xor U22695 (N_22695,N_22249,N_22299);
and U22696 (N_22696,N_22449,N_22473);
or U22697 (N_22697,N_22272,N_22470);
nor U22698 (N_22698,N_22287,N_22358);
and U22699 (N_22699,N_22433,N_22328);
nor U22700 (N_22700,N_22316,N_22262);
or U22701 (N_22701,N_22269,N_22408);
or U22702 (N_22702,N_22278,N_22234);
and U22703 (N_22703,N_22230,N_22441);
xnor U22704 (N_22704,N_22211,N_22305);
nor U22705 (N_22705,N_22218,N_22374);
nor U22706 (N_22706,N_22278,N_22365);
or U22707 (N_22707,N_22479,N_22410);
nand U22708 (N_22708,N_22273,N_22229);
and U22709 (N_22709,N_22213,N_22490);
or U22710 (N_22710,N_22389,N_22436);
and U22711 (N_22711,N_22273,N_22250);
xnor U22712 (N_22712,N_22353,N_22376);
nor U22713 (N_22713,N_22323,N_22410);
xnor U22714 (N_22714,N_22286,N_22395);
nand U22715 (N_22715,N_22271,N_22274);
xor U22716 (N_22716,N_22263,N_22268);
xnor U22717 (N_22717,N_22225,N_22380);
or U22718 (N_22718,N_22487,N_22383);
and U22719 (N_22719,N_22445,N_22277);
nand U22720 (N_22720,N_22295,N_22275);
or U22721 (N_22721,N_22262,N_22272);
or U22722 (N_22722,N_22202,N_22447);
xnor U22723 (N_22723,N_22324,N_22360);
and U22724 (N_22724,N_22384,N_22325);
nor U22725 (N_22725,N_22276,N_22399);
or U22726 (N_22726,N_22416,N_22453);
nand U22727 (N_22727,N_22451,N_22395);
and U22728 (N_22728,N_22205,N_22215);
nor U22729 (N_22729,N_22369,N_22205);
nor U22730 (N_22730,N_22321,N_22393);
nand U22731 (N_22731,N_22271,N_22269);
and U22732 (N_22732,N_22426,N_22259);
nand U22733 (N_22733,N_22252,N_22309);
and U22734 (N_22734,N_22376,N_22342);
or U22735 (N_22735,N_22380,N_22373);
nand U22736 (N_22736,N_22404,N_22448);
or U22737 (N_22737,N_22421,N_22475);
nor U22738 (N_22738,N_22299,N_22239);
nor U22739 (N_22739,N_22359,N_22338);
nor U22740 (N_22740,N_22280,N_22453);
and U22741 (N_22741,N_22217,N_22333);
nand U22742 (N_22742,N_22478,N_22395);
nor U22743 (N_22743,N_22207,N_22489);
nand U22744 (N_22744,N_22417,N_22446);
or U22745 (N_22745,N_22353,N_22234);
nor U22746 (N_22746,N_22484,N_22415);
nand U22747 (N_22747,N_22312,N_22208);
or U22748 (N_22748,N_22374,N_22473);
and U22749 (N_22749,N_22302,N_22453);
xnor U22750 (N_22750,N_22402,N_22442);
or U22751 (N_22751,N_22461,N_22337);
nand U22752 (N_22752,N_22286,N_22411);
nand U22753 (N_22753,N_22402,N_22470);
nand U22754 (N_22754,N_22393,N_22497);
nor U22755 (N_22755,N_22378,N_22350);
nand U22756 (N_22756,N_22278,N_22448);
nor U22757 (N_22757,N_22387,N_22328);
nor U22758 (N_22758,N_22473,N_22357);
or U22759 (N_22759,N_22208,N_22478);
and U22760 (N_22760,N_22258,N_22345);
nand U22761 (N_22761,N_22470,N_22333);
nor U22762 (N_22762,N_22458,N_22382);
and U22763 (N_22763,N_22212,N_22347);
and U22764 (N_22764,N_22274,N_22477);
and U22765 (N_22765,N_22330,N_22339);
nand U22766 (N_22766,N_22380,N_22341);
nor U22767 (N_22767,N_22428,N_22444);
nor U22768 (N_22768,N_22482,N_22251);
nor U22769 (N_22769,N_22378,N_22411);
nand U22770 (N_22770,N_22462,N_22317);
nand U22771 (N_22771,N_22314,N_22269);
nand U22772 (N_22772,N_22241,N_22414);
and U22773 (N_22773,N_22233,N_22412);
and U22774 (N_22774,N_22235,N_22316);
nor U22775 (N_22775,N_22492,N_22244);
nand U22776 (N_22776,N_22218,N_22371);
xor U22777 (N_22777,N_22324,N_22256);
and U22778 (N_22778,N_22223,N_22421);
nor U22779 (N_22779,N_22394,N_22418);
xor U22780 (N_22780,N_22454,N_22308);
xor U22781 (N_22781,N_22208,N_22499);
nor U22782 (N_22782,N_22285,N_22338);
or U22783 (N_22783,N_22331,N_22243);
nor U22784 (N_22784,N_22420,N_22342);
or U22785 (N_22785,N_22488,N_22212);
or U22786 (N_22786,N_22262,N_22201);
and U22787 (N_22787,N_22450,N_22297);
or U22788 (N_22788,N_22235,N_22256);
and U22789 (N_22789,N_22208,N_22328);
xnor U22790 (N_22790,N_22273,N_22279);
nand U22791 (N_22791,N_22258,N_22288);
nand U22792 (N_22792,N_22398,N_22258);
nand U22793 (N_22793,N_22450,N_22214);
nand U22794 (N_22794,N_22390,N_22422);
or U22795 (N_22795,N_22210,N_22357);
nand U22796 (N_22796,N_22219,N_22403);
and U22797 (N_22797,N_22212,N_22278);
xnor U22798 (N_22798,N_22297,N_22283);
and U22799 (N_22799,N_22319,N_22402);
or U22800 (N_22800,N_22799,N_22755);
and U22801 (N_22801,N_22708,N_22631);
nand U22802 (N_22802,N_22795,N_22734);
or U22803 (N_22803,N_22528,N_22653);
nor U22804 (N_22804,N_22591,N_22738);
and U22805 (N_22805,N_22730,N_22683);
or U22806 (N_22806,N_22772,N_22507);
nor U22807 (N_22807,N_22583,N_22532);
nor U22808 (N_22808,N_22557,N_22508);
xor U22809 (N_22809,N_22668,N_22787);
nand U22810 (N_22810,N_22602,N_22779);
nor U22811 (N_22811,N_22530,N_22641);
nor U22812 (N_22812,N_22605,N_22661);
nand U22813 (N_22813,N_22623,N_22770);
or U22814 (N_22814,N_22526,N_22645);
and U22815 (N_22815,N_22617,N_22614);
xor U22816 (N_22816,N_22718,N_22757);
nand U22817 (N_22817,N_22639,N_22760);
nor U22818 (N_22818,N_22626,N_22759);
nor U22819 (N_22819,N_22548,N_22589);
xor U22820 (N_22820,N_22769,N_22776);
xor U22821 (N_22821,N_22505,N_22567);
or U22822 (N_22822,N_22585,N_22588);
xor U22823 (N_22823,N_22731,N_22594);
or U22824 (N_22824,N_22727,N_22774);
xor U22825 (N_22825,N_22549,N_22612);
nand U22826 (N_22826,N_22579,N_22762);
nand U22827 (N_22827,N_22790,N_22761);
xor U22828 (N_22828,N_22542,N_22563);
nor U22829 (N_22829,N_22729,N_22522);
and U22830 (N_22830,N_22705,N_22561);
nand U22831 (N_22831,N_22552,N_22573);
nor U22832 (N_22832,N_22722,N_22611);
nor U22833 (N_22833,N_22741,N_22778);
or U22834 (N_22834,N_22655,N_22686);
nand U22835 (N_22835,N_22749,N_22527);
nor U22836 (N_22836,N_22764,N_22572);
nand U22837 (N_22837,N_22791,N_22740);
nor U22838 (N_22838,N_22581,N_22745);
or U22839 (N_22839,N_22514,N_22712);
nand U22840 (N_22840,N_22586,N_22679);
nand U22841 (N_22841,N_22562,N_22553);
and U22842 (N_22842,N_22644,N_22750);
xor U22843 (N_22843,N_22606,N_22698);
and U22844 (N_22844,N_22502,N_22516);
or U22845 (N_22845,N_22540,N_22656);
nor U22846 (N_22846,N_22580,N_22650);
xor U22847 (N_22847,N_22765,N_22739);
or U22848 (N_22848,N_22674,N_22696);
or U22849 (N_22849,N_22569,N_22638);
or U22850 (N_22850,N_22733,N_22637);
nor U22851 (N_22851,N_22609,N_22578);
or U22852 (N_22852,N_22535,N_22700);
or U22853 (N_22853,N_22667,N_22719);
nor U22854 (N_22854,N_22664,N_22780);
xor U22855 (N_22855,N_22701,N_22517);
xnor U22856 (N_22856,N_22649,N_22775);
nand U22857 (N_22857,N_22554,N_22789);
nand U22858 (N_22858,N_22681,N_22544);
nor U22859 (N_22859,N_22682,N_22666);
xnor U22860 (N_22860,N_22736,N_22720);
nor U22861 (N_22861,N_22545,N_22515);
nand U22862 (N_22862,N_22537,N_22788);
xnor U22863 (N_22863,N_22642,N_22504);
nand U22864 (N_22864,N_22782,N_22794);
xnor U22865 (N_22865,N_22568,N_22500);
xnor U22866 (N_22866,N_22771,N_22630);
xnor U22867 (N_22867,N_22798,N_22703);
and U22868 (N_22868,N_22640,N_22747);
and U22869 (N_22869,N_22506,N_22744);
or U22870 (N_22870,N_22558,N_22556);
and U22871 (N_22871,N_22533,N_22793);
nand U22872 (N_22872,N_22582,N_22726);
nor U22873 (N_22873,N_22543,N_22797);
xor U22874 (N_22874,N_22518,N_22783);
nor U22875 (N_22875,N_22601,N_22560);
and U22876 (N_22876,N_22695,N_22675);
and U22877 (N_22877,N_22574,N_22538);
nor U22878 (N_22878,N_22657,N_22627);
nor U22879 (N_22879,N_22732,N_22636);
or U22880 (N_22880,N_22559,N_22531);
and U22881 (N_22881,N_22629,N_22704);
or U22882 (N_22882,N_22723,N_22711);
and U22883 (N_22883,N_22691,N_22539);
nand U22884 (N_22884,N_22633,N_22746);
or U22885 (N_22885,N_22785,N_22714);
xnor U22886 (N_22886,N_22587,N_22784);
nand U22887 (N_22887,N_22752,N_22669);
or U22888 (N_22888,N_22680,N_22520);
nand U22889 (N_22889,N_22768,N_22743);
or U22890 (N_22890,N_22763,N_22707);
nand U22891 (N_22891,N_22616,N_22503);
xnor U22892 (N_22892,N_22603,N_22725);
nor U22893 (N_22893,N_22519,N_22600);
and U22894 (N_22894,N_22754,N_22748);
nor U22895 (N_22895,N_22510,N_22724);
or U22896 (N_22896,N_22575,N_22786);
or U22897 (N_22897,N_22628,N_22570);
or U22898 (N_22898,N_22524,N_22697);
and U22899 (N_22899,N_22792,N_22521);
nand U22900 (N_22900,N_22756,N_22663);
nand U22901 (N_22901,N_22670,N_22654);
nand U22902 (N_22902,N_22576,N_22721);
and U22903 (N_22903,N_22662,N_22608);
nand U22904 (N_22904,N_22687,N_22742);
xnor U22905 (N_22905,N_22547,N_22607);
xnor U22906 (N_22906,N_22692,N_22584);
xor U22907 (N_22907,N_22676,N_22753);
and U22908 (N_22908,N_22737,N_22660);
xor U22909 (N_22909,N_22541,N_22777);
or U22910 (N_22910,N_22672,N_22716);
or U22911 (N_22911,N_22566,N_22647);
nor U22912 (N_22912,N_22525,N_22643);
nor U22913 (N_22913,N_22796,N_22595);
xor U22914 (N_22914,N_22685,N_22625);
or U22915 (N_22915,N_22599,N_22717);
nand U22916 (N_22916,N_22593,N_22635);
or U22917 (N_22917,N_22546,N_22615);
xor U22918 (N_22918,N_22702,N_22551);
nand U22919 (N_22919,N_22671,N_22565);
nor U22920 (N_22920,N_22690,N_22673);
nor U22921 (N_22921,N_22513,N_22598);
and U22922 (N_22922,N_22651,N_22597);
nand U22923 (N_22923,N_22693,N_22699);
xnor U22924 (N_22924,N_22501,N_22632);
nand U22925 (N_22925,N_22646,N_22622);
xor U22926 (N_22926,N_22689,N_22659);
or U22927 (N_22927,N_22652,N_22592);
nand U22928 (N_22928,N_22710,N_22610);
or U22929 (N_22929,N_22735,N_22590);
nand U22930 (N_22930,N_22534,N_22677);
and U22931 (N_22931,N_22781,N_22758);
xor U22932 (N_22932,N_22613,N_22596);
nand U22933 (N_22933,N_22751,N_22709);
xor U22934 (N_22934,N_22713,N_22529);
nand U22935 (N_22935,N_22767,N_22536);
nand U22936 (N_22936,N_22509,N_22523);
xnor U22937 (N_22937,N_22634,N_22773);
xnor U22938 (N_22938,N_22706,N_22624);
or U22939 (N_22939,N_22648,N_22577);
and U22940 (N_22940,N_22550,N_22694);
nand U22941 (N_22941,N_22618,N_22555);
nand U22942 (N_22942,N_22511,N_22619);
or U22943 (N_22943,N_22715,N_22512);
nand U22944 (N_22944,N_22665,N_22658);
and U22945 (N_22945,N_22688,N_22684);
or U22946 (N_22946,N_22604,N_22620);
nand U22947 (N_22947,N_22728,N_22766);
nor U22948 (N_22948,N_22571,N_22564);
or U22949 (N_22949,N_22678,N_22621);
nand U22950 (N_22950,N_22668,N_22518);
xor U22951 (N_22951,N_22532,N_22589);
or U22952 (N_22952,N_22555,N_22617);
nand U22953 (N_22953,N_22796,N_22750);
xnor U22954 (N_22954,N_22790,N_22647);
or U22955 (N_22955,N_22616,N_22701);
and U22956 (N_22956,N_22587,N_22701);
and U22957 (N_22957,N_22727,N_22618);
xor U22958 (N_22958,N_22545,N_22691);
nor U22959 (N_22959,N_22679,N_22558);
or U22960 (N_22960,N_22592,N_22744);
or U22961 (N_22961,N_22545,N_22625);
nor U22962 (N_22962,N_22782,N_22563);
or U22963 (N_22963,N_22656,N_22581);
and U22964 (N_22964,N_22628,N_22625);
nor U22965 (N_22965,N_22552,N_22584);
nor U22966 (N_22966,N_22568,N_22660);
or U22967 (N_22967,N_22674,N_22584);
nand U22968 (N_22968,N_22791,N_22595);
nor U22969 (N_22969,N_22617,N_22708);
xnor U22970 (N_22970,N_22531,N_22751);
or U22971 (N_22971,N_22691,N_22648);
and U22972 (N_22972,N_22766,N_22537);
and U22973 (N_22973,N_22769,N_22532);
xnor U22974 (N_22974,N_22576,N_22551);
nor U22975 (N_22975,N_22673,N_22732);
or U22976 (N_22976,N_22738,N_22613);
and U22977 (N_22977,N_22517,N_22620);
xor U22978 (N_22978,N_22728,N_22648);
nand U22979 (N_22979,N_22645,N_22523);
or U22980 (N_22980,N_22737,N_22761);
nor U22981 (N_22981,N_22560,N_22731);
xor U22982 (N_22982,N_22644,N_22589);
nor U22983 (N_22983,N_22528,N_22763);
xor U22984 (N_22984,N_22764,N_22654);
nand U22985 (N_22985,N_22731,N_22523);
nor U22986 (N_22986,N_22526,N_22527);
xnor U22987 (N_22987,N_22632,N_22680);
nor U22988 (N_22988,N_22573,N_22536);
nand U22989 (N_22989,N_22569,N_22712);
xnor U22990 (N_22990,N_22525,N_22758);
and U22991 (N_22991,N_22669,N_22736);
xor U22992 (N_22992,N_22601,N_22765);
or U22993 (N_22993,N_22710,N_22537);
xor U22994 (N_22994,N_22784,N_22726);
and U22995 (N_22995,N_22677,N_22667);
nor U22996 (N_22996,N_22508,N_22541);
and U22997 (N_22997,N_22572,N_22510);
or U22998 (N_22998,N_22596,N_22733);
or U22999 (N_22999,N_22750,N_22558);
or U23000 (N_23000,N_22519,N_22645);
nand U23001 (N_23001,N_22599,N_22788);
or U23002 (N_23002,N_22730,N_22692);
nor U23003 (N_23003,N_22530,N_22580);
xor U23004 (N_23004,N_22695,N_22571);
xnor U23005 (N_23005,N_22685,N_22660);
nor U23006 (N_23006,N_22515,N_22522);
nand U23007 (N_23007,N_22715,N_22526);
xor U23008 (N_23008,N_22756,N_22689);
or U23009 (N_23009,N_22526,N_22531);
nand U23010 (N_23010,N_22525,N_22620);
nand U23011 (N_23011,N_22587,N_22697);
xnor U23012 (N_23012,N_22710,N_22647);
xnor U23013 (N_23013,N_22555,N_22577);
or U23014 (N_23014,N_22522,N_22630);
nor U23015 (N_23015,N_22720,N_22758);
and U23016 (N_23016,N_22542,N_22590);
and U23017 (N_23017,N_22535,N_22616);
or U23018 (N_23018,N_22614,N_22735);
xor U23019 (N_23019,N_22685,N_22520);
or U23020 (N_23020,N_22791,N_22519);
nand U23021 (N_23021,N_22569,N_22764);
xor U23022 (N_23022,N_22596,N_22790);
and U23023 (N_23023,N_22590,N_22642);
nand U23024 (N_23024,N_22743,N_22632);
nor U23025 (N_23025,N_22622,N_22743);
or U23026 (N_23026,N_22686,N_22615);
or U23027 (N_23027,N_22542,N_22627);
nand U23028 (N_23028,N_22672,N_22770);
xnor U23029 (N_23029,N_22595,N_22554);
xor U23030 (N_23030,N_22544,N_22638);
nor U23031 (N_23031,N_22595,N_22633);
nand U23032 (N_23032,N_22578,N_22659);
nand U23033 (N_23033,N_22711,N_22630);
nor U23034 (N_23034,N_22698,N_22701);
nor U23035 (N_23035,N_22667,N_22781);
or U23036 (N_23036,N_22718,N_22753);
nor U23037 (N_23037,N_22501,N_22773);
and U23038 (N_23038,N_22552,N_22647);
xor U23039 (N_23039,N_22505,N_22557);
and U23040 (N_23040,N_22567,N_22771);
xnor U23041 (N_23041,N_22735,N_22524);
nor U23042 (N_23042,N_22575,N_22571);
or U23043 (N_23043,N_22518,N_22728);
and U23044 (N_23044,N_22590,N_22555);
xor U23045 (N_23045,N_22502,N_22694);
nor U23046 (N_23046,N_22632,N_22635);
nor U23047 (N_23047,N_22671,N_22709);
xor U23048 (N_23048,N_22687,N_22641);
or U23049 (N_23049,N_22798,N_22630);
or U23050 (N_23050,N_22547,N_22646);
or U23051 (N_23051,N_22638,N_22750);
nor U23052 (N_23052,N_22745,N_22714);
or U23053 (N_23053,N_22534,N_22744);
and U23054 (N_23054,N_22738,N_22731);
nor U23055 (N_23055,N_22558,N_22521);
nand U23056 (N_23056,N_22681,N_22690);
nand U23057 (N_23057,N_22742,N_22795);
and U23058 (N_23058,N_22533,N_22643);
nor U23059 (N_23059,N_22755,N_22666);
nand U23060 (N_23060,N_22705,N_22587);
xor U23061 (N_23061,N_22614,N_22509);
nor U23062 (N_23062,N_22697,N_22718);
nand U23063 (N_23063,N_22674,N_22614);
or U23064 (N_23064,N_22549,N_22637);
nor U23065 (N_23065,N_22557,N_22751);
xor U23066 (N_23066,N_22523,N_22605);
or U23067 (N_23067,N_22644,N_22656);
and U23068 (N_23068,N_22787,N_22786);
nor U23069 (N_23069,N_22673,N_22753);
or U23070 (N_23070,N_22715,N_22586);
or U23071 (N_23071,N_22663,N_22583);
nand U23072 (N_23072,N_22510,N_22520);
or U23073 (N_23073,N_22656,N_22516);
or U23074 (N_23074,N_22590,N_22643);
and U23075 (N_23075,N_22704,N_22757);
xor U23076 (N_23076,N_22659,N_22534);
and U23077 (N_23077,N_22573,N_22788);
xnor U23078 (N_23078,N_22584,N_22724);
xnor U23079 (N_23079,N_22535,N_22546);
xor U23080 (N_23080,N_22563,N_22663);
nor U23081 (N_23081,N_22768,N_22748);
and U23082 (N_23082,N_22604,N_22627);
nor U23083 (N_23083,N_22553,N_22699);
xnor U23084 (N_23084,N_22665,N_22709);
nand U23085 (N_23085,N_22754,N_22578);
and U23086 (N_23086,N_22675,N_22793);
or U23087 (N_23087,N_22792,N_22566);
or U23088 (N_23088,N_22768,N_22564);
or U23089 (N_23089,N_22770,N_22710);
xor U23090 (N_23090,N_22573,N_22775);
and U23091 (N_23091,N_22768,N_22628);
nor U23092 (N_23092,N_22600,N_22763);
and U23093 (N_23093,N_22557,N_22791);
xor U23094 (N_23094,N_22670,N_22761);
and U23095 (N_23095,N_22585,N_22720);
or U23096 (N_23096,N_22593,N_22554);
nor U23097 (N_23097,N_22578,N_22591);
xor U23098 (N_23098,N_22553,N_22703);
nor U23099 (N_23099,N_22701,N_22775);
xor U23100 (N_23100,N_22825,N_23054);
or U23101 (N_23101,N_22883,N_22894);
xor U23102 (N_23102,N_22882,N_22927);
or U23103 (N_23103,N_22975,N_23050);
xnor U23104 (N_23104,N_23027,N_22807);
or U23105 (N_23105,N_23097,N_22818);
and U23106 (N_23106,N_23007,N_22897);
nand U23107 (N_23107,N_22913,N_23089);
xor U23108 (N_23108,N_22892,N_23049);
nor U23109 (N_23109,N_23074,N_22817);
nor U23110 (N_23110,N_22843,N_22877);
and U23111 (N_23111,N_22985,N_22865);
and U23112 (N_23112,N_22950,N_22961);
xor U23113 (N_23113,N_22871,N_22858);
and U23114 (N_23114,N_22964,N_22845);
xnor U23115 (N_23115,N_23009,N_23099);
nand U23116 (N_23116,N_22984,N_22988);
xnor U23117 (N_23117,N_23069,N_23016);
nor U23118 (N_23118,N_22889,N_23033);
and U23119 (N_23119,N_22943,N_23055);
nor U23120 (N_23120,N_22827,N_22955);
and U23121 (N_23121,N_22886,N_22868);
and U23122 (N_23122,N_23066,N_23026);
nor U23123 (N_23123,N_22954,N_22905);
nor U23124 (N_23124,N_23085,N_22936);
or U23125 (N_23125,N_23041,N_22866);
xnor U23126 (N_23126,N_22924,N_23096);
nand U23127 (N_23127,N_22930,N_23025);
nand U23128 (N_23128,N_22801,N_22862);
or U23129 (N_23129,N_23048,N_22947);
or U23130 (N_23130,N_22829,N_22931);
or U23131 (N_23131,N_23019,N_23042);
xnor U23132 (N_23132,N_22802,N_22884);
nand U23133 (N_23133,N_22870,N_22838);
nand U23134 (N_23134,N_22828,N_22980);
nor U23135 (N_23135,N_22855,N_22847);
nor U23136 (N_23136,N_22902,N_22903);
nor U23137 (N_23137,N_22959,N_23056);
and U23138 (N_23138,N_23031,N_22813);
xor U23139 (N_23139,N_23084,N_22873);
or U23140 (N_23140,N_23006,N_23030);
nor U23141 (N_23141,N_23024,N_22990);
nor U23142 (N_23142,N_22850,N_22876);
nand U23143 (N_23143,N_22932,N_22972);
and U23144 (N_23144,N_22812,N_22803);
nor U23145 (N_23145,N_23008,N_22916);
xnor U23146 (N_23146,N_22965,N_22987);
nand U23147 (N_23147,N_22944,N_23010);
nand U23148 (N_23148,N_22998,N_22928);
nor U23149 (N_23149,N_22842,N_23004);
nand U23150 (N_23150,N_22839,N_22929);
nand U23151 (N_23151,N_22983,N_22923);
nand U23152 (N_23152,N_22914,N_22821);
and U23153 (N_23153,N_22958,N_22853);
xor U23154 (N_23154,N_23076,N_23022);
nor U23155 (N_23155,N_23045,N_23072);
nand U23156 (N_23156,N_23018,N_22901);
xnor U23157 (N_23157,N_22835,N_22997);
nand U23158 (N_23158,N_22945,N_22860);
and U23159 (N_23159,N_22887,N_23040);
xor U23160 (N_23160,N_22826,N_22977);
xor U23161 (N_23161,N_22879,N_22906);
xnor U23162 (N_23162,N_22808,N_23094);
or U23163 (N_23163,N_22859,N_22974);
and U23164 (N_23164,N_23095,N_22836);
and U23165 (N_23165,N_23032,N_23086);
nand U23166 (N_23166,N_23017,N_22819);
xor U23167 (N_23167,N_23090,N_22957);
xor U23168 (N_23168,N_22895,N_23063);
and U23169 (N_23169,N_23080,N_22992);
xnor U23170 (N_23170,N_22814,N_22949);
and U23171 (N_23171,N_23020,N_22849);
nand U23172 (N_23172,N_23021,N_22934);
or U23173 (N_23173,N_23064,N_22996);
and U23174 (N_23174,N_22846,N_23082);
xor U23175 (N_23175,N_23060,N_22976);
or U23176 (N_23176,N_23029,N_22854);
and U23177 (N_23177,N_22926,N_23057);
nand U23178 (N_23178,N_22938,N_22874);
or U23179 (N_23179,N_22844,N_22922);
nand U23180 (N_23180,N_23077,N_22952);
xor U23181 (N_23181,N_22920,N_22937);
xnor U23182 (N_23182,N_22811,N_23071);
nor U23183 (N_23183,N_23075,N_23014);
and U23184 (N_23184,N_22810,N_22890);
nand U23185 (N_23185,N_23002,N_22933);
nor U23186 (N_23186,N_22994,N_22872);
nand U23187 (N_23187,N_22939,N_22917);
and U23188 (N_23188,N_23051,N_23015);
xor U23189 (N_23189,N_22912,N_22848);
nand U23190 (N_23190,N_22951,N_23039);
xor U23191 (N_23191,N_22898,N_22935);
xnor U23192 (N_23192,N_22918,N_23065);
nor U23193 (N_23193,N_23034,N_23028);
and U23194 (N_23194,N_22911,N_22875);
nor U23195 (N_23195,N_23043,N_23038);
nand U23196 (N_23196,N_22900,N_23037);
nor U23197 (N_23197,N_22910,N_22820);
nand U23198 (N_23198,N_22981,N_22968);
or U23199 (N_23199,N_23011,N_22856);
and U23200 (N_23200,N_23052,N_23036);
xnor U23201 (N_23201,N_22971,N_23023);
xnor U23202 (N_23202,N_22999,N_23083);
or U23203 (N_23203,N_22940,N_22960);
and U23204 (N_23204,N_22919,N_23079);
or U23205 (N_23205,N_22925,N_22823);
nor U23206 (N_23206,N_23073,N_23046);
xnor U23207 (N_23207,N_22824,N_22963);
or U23208 (N_23208,N_22837,N_22982);
nor U23209 (N_23209,N_22851,N_22948);
and U23210 (N_23210,N_22881,N_22816);
nand U23211 (N_23211,N_22832,N_22840);
nand U23212 (N_23212,N_23005,N_22921);
nand U23213 (N_23213,N_22809,N_22831);
nand U23214 (N_23214,N_22908,N_23091);
or U23215 (N_23215,N_22888,N_22893);
nand U23216 (N_23216,N_22899,N_23068);
or U23217 (N_23217,N_22969,N_22993);
nor U23218 (N_23218,N_23067,N_22942);
nor U23219 (N_23219,N_23088,N_22857);
or U23220 (N_23220,N_23003,N_22953);
xnor U23221 (N_23221,N_22979,N_22864);
xnor U23222 (N_23222,N_22946,N_22891);
nand U23223 (N_23223,N_22907,N_22804);
nand U23224 (N_23224,N_22991,N_22880);
and U23225 (N_23225,N_22941,N_22878);
nand U23226 (N_23226,N_22967,N_22805);
or U23227 (N_23227,N_23012,N_22852);
nand U23228 (N_23228,N_22830,N_22989);
nand U23229 (N_23229,N_22863,N_23058);
nor U23230 (N_23230,N_22896,N_22861);
xor U23231 (N_23231,N_22978,N_23093);
and U23232 (N_23232,N_22833,N_22904);
nand U23233 (N_23233,N_22956,N_22867);
nand U23234 (N_23234,N_22973,N_23081);
and U23235 (N_23235,N_22995,N_23044);
nor U23236 (N_23236,N_23059,N_23053);
xnor U23237 (N_23237,N_23047,N_22885);
and U23238 (N_23238,N_23000,N_23078);
xor U23239 (N_23239,N_22909,N_22966);
nor U23240 (N_23240,N_23035,N_22834);
and U23241 (N_23241,N_23013,N_22970);
nor U23242 (N_23242,N_23061,N_22800);
nor U23243 (N_23243,N_23092,N_22986);
nor U23244 (N_23244,N_22869,N_22915);
and U23245 (N_23245,N_22822,N_22815);
nand U23246 (N_23246,N_22962,N_23001);
xor U23247 (N_23247,N_23087,N_23070);
xnor U23248 (N_23248,N_22806,N_23098);
nand U23249 (N_23249,N_22841,N_23062);
nor U23250 (N_23250,N_23051,N_22928);
xor U23251 (N_23251,N_22810,N_22831);
nand U23252 (N_23252,N_22971,N_23082);
and U23253 (N_23253,N_22942,N_22907);
and U23254 (N_23254,N_22862,N_22836);
xor U23255 (N_23255,N_22988,N_22803);
and U23256 (N_23256,N_23066,N_23098);
xor U23257 (N_23257,N_22917,N_23003);
or U23258 (N_23258,N_23093,N_22874);
nor U23259 (N_23259,N_22806,N_23068);
xnor U23260 (N_23260,N_23054,N_22837);
nand U23261 (N_23261,N_22800,N_22990);
nor U23262 (N_23262,N_22836,N_22989);
nor U23263 (N_23263,N_22865,N_22893);
nor U23264 (N_23264,N_22975,N_22819);
nor U23265 (N_23265,N_23099,N_23068);
or U23266 (N_23266,N_22804,N_23062);
and U23267 (N_23267,N_22878,N_22975);
or U23268 (N_23268,N_22919,N_23091);
nor U23269 (N_23269,N_22835,N_22839);
xor U23270 (N_23270,N_22965,N_22839);
nand U23271 (N_23271,N_22845,N_23069);
nand U23272 (N_23272,N_22822,N_23025);
or U23273 (N_23273,N_23044,N_22866);
or U23274 (N_23274,N_23097,N_22833);
xor U23275 (N_23275,N_22972,N_23056);
and U23276 (N_23276,N_22850,N_22890);
nor U23277 (N_23277,N_23031,N_22919);
xor U23278 (N_23278,N_22932,N_22822);
nand U23279 (N_23279,N_22928,N_23039);
nor U23280 (N_23280,N_22946,N_22817);
nor U23281 (N_23281,N_23057,N_22909);
xnor U23282 (N_23282,N_23048,N_23061);
and U23283 (N_23283,N_22834,N_23054);
nor U23284 (N_23284,N_23019,N_23014);
nor U23285 (N_23285,N_23086,N_22990);
and U23286 (N_23286,N_23089,N_23002);
nand U23287 (N_23287,N_23081,N_23089);
nor U23288 (N_23288,N_22858,N_22992);
xor U23289 (N_23289,N_23030,N_22994);
and U23290 (N_23290,N_22877,N_22995);
xor U23291 (N_23291,N_22991,N_23062);
or U23292 (N_23292,N_22866,N_22921);
nor U23293 (N_23293,N_22966,N_22981);
nand U23294 (N_23294,N_22858,N_23022);
and U23295 (N_23295,N_23025,N_23047);
and U23296 (N_23296,N_22986,N_23086);
nor U23297 (N_23297,N_23049,N_23061);
nand U23298 (N_23298,N_23079,N_22849);
and U23299 (N_23299,N_22836,N_23059);
nand U23300 (N_23300,N_22971,N_22837);
or U23301 (N_23301,N_22934,N_23015);
nor U23302 (N_23302,N_23073,N_22928);
nor U23303 (N_23303,N_22803,N_23028);
and U23304 (N_23304,N_22930,N_22959);
nand U23305 (N_23305,N_22946,N_23034);
nor U23306 (N_23306,N_22807,N_23067);
xor U23307 (N_23307,N_23082,N_22849);
xor U23308 (N_23308,N_23002,N_22872);
xor U23309 (N_23309,N_23031,N_23083);
and U23310 (N_23310,N_22885,N_23018);
or U23311 (N_23311,N_22983,N_23064);
or U23312 (N_23312,N_22925,N_22988);
and U23313 (N_23313,N_22993,N_23024);
or U23314 (N_23314,N_22927,N_23037);
and U23315 (N_23315,N_22983,N_23055);
or U23316 (N_23316,N_22950,N_23047);
or U23317 (N_23317,N_23084,N_23041);
and U23318 (N_23318,N_22921,N_22909);
or U23319 (N_23319,N_22882,N_22982);
or U23320 (N_23320,N_22975,N_22974);
nor U23321 (N_23321,N_22932,N_22987);
xnor U23322 (N_23322,N_22929,N_22986);
nor U23323 (N_23323,N_22907,N_22994);
and U23324 (N_23324,N_22808,N_22906);
and U23325 (N_23325,N_22994,N_22810);
and U23326 (N_23326,N_23033,N_22917);
nand U23327 (N_23327,N_23033,N_23071);
xor U23328 (N_23328,N_23063,N_22841);
xor U23329 (N_23329,N_22837,N_22820);
xnor U23330 (N_23330,N_22900,N_23069);
or U23331 (N_23331,N_22982,N_22818);
or U23332 (N_23332,N_22833,N_23060);
xnor U23333 (N_23333,N_22812,N_22901);
and U23334 (N_23334,N_22972,N_22976);
nand U23335 (N_23335,N_22868,N_23080);
or U23336 (N_23336,N_22991,N_22994);
and U23337 (N_23337,N_23067,N_22936);
or U23338 (N_23338,N_23060,N_22942);
nand U23339 (N_23339,N_23002,N_23048);
or U23340 (N_23340,N_22975,N_22991);
xnor U23341 (N_23341,N_22921,N_22820);
or U23342 (N_23342,N_23087,N_23063);
xor U23343 (N_23343,N_23003,N_23086);
nor U23344 (N_23344,N_22940,N_23070);
nand U23345 (N_23345,N_22816,N_23025);
xnor U23346 (N_23346,N_22914,N_22822);
or U23347 (N_23347,N_23024,N_22896);
or U23348 (N_23348,N_22840,N_23079);
xor U23349 (N_23349,N_22964,N_23022);
or U23350 (N_23350,N_23056,N_22843);
and U23351 (N_23351,N_23037,N_23080);
or U23352 (N_23352,N_22803,N_22895);
or U23353 (N_23353,N_22914,N_22855);
xor U23354 (N_23354,N_22959,N_23075);
nand U23355 (N_23355,N_22904,N_22991);
nand U23356 (N_23356,N_23051,N_22914);
xnor U23357 (N_23357,N_22996,N_22860);
xor U23358 (N_23358,N_22957,N_23076);
xor U23359 (N_23359,N_22827,N_23003);
xnor U23360 (N_23360,N_22875,N_22889);
nor U23361 (N_23361,N_22924,N_22984);
xnor U23362 (N_23362,N_23087,N_22979);
or U23363 (N_23363,N_22848,N_23030);
or U23364 (N_23364,N_22944,N_23068);
nand U23365 (N_23365,N_22921,N_22972);
nand U23366 (N_23366,N_22895,N_22848);
and U23367 (N_23367,N_23052,N_23019);
or U23368 (N_23368,N_23058,N_22810);
nor U23369 (N_23369,N_22814,N_22810);
xnor U23370 (N_23370,N_22855,N_22944);
nand U23371 (N_23371,N_22801,N_23033);
nand U23372 (N_23372,N_22811,N_23094);
or U23373 (N_23373,N_22982,N_22966);
nor U23374 (N_23374,N_22930,N_23062);
and U23375 (N_23375,N_22832,N_22849);
xor U23376 (N_23376,N_22839,N_22856);
nor U23377 (N_23377,N_22823,N_22953);
or U23378 (N_23378,N_22968,N_22842);
xnor U23379 (N_23379,N_22861,N_22818);
nor U23380 (N_23380,N_22899,N_23071);
and U23381 (N_23381,N_23015,N_22858);
or U23382 (N_23382,N_23084,N_22931);
and U23383 (N_23383,N_22975,N_22856);
or U23384 (N_23384,N_23097,N_22995);
nand U23385 (N_23385,N_23009,N_22981);
or U23386 (N_23386,N_23093,N_22817);
and U23387 (N_23387,N_22910,N_22995);
and U23388 (N_23388,N_23047,N_22917);
or U23389 (N_23389,N_22857,N_23007);
and U23390 (N_23390,N_22847,N_23012);
nand U23391 (N_23391,N_22891,N_22858);
nor U23392 (N_23392,N_23080,N_22949);
nand U23393 (N_23393,N_22882,N_22826);
or U23394 (N_23394,N_23093,N_22968);
nand U23395 (N_23395,N_23000,N_22803);
and U23396 (N_23396,N_22808,N_22889);
or U23397 (N_23397,N_22839,N_22937);
nor U23398 (N_23398,N_22945,N_23055);
or U23399 (N_23399,N_22870,N_23030);
xnor U23400 (N_23400,N_23239,N_23177);
or U23401 (N_23401,N_23197,N_23158);
nor U23402 (N_23402,N_23272,N_23243);
and U23403 (N_23403,N_23331,N_23136);
and U23404 (N_23404,N_23351,N_23325);
and U23405 (N_23405,N_23375,N_23286);
nor U23406 (N_23406,N_23297,N_23104);
nand U23407 (N_23407,N_23121,N_23291);
nor U23408 (N_23408,N_23112,N_23228);
nand U23409 (N_23409,N_23192,N_23357);
or U23410 (N_23410,N_23203,N_23361);
xor U23411 (N_23411,N_23290,N_23316);
and U23412 (N_23412,N_23358,N_23265);
or U23413 (N_23413,N_23380,N_23269);
and U23414 (N_23414,N_23343,N_23374);
nor U23415 (N_23415,N_23248,N_23370);
or U23416 (N_23416,N_23268,N_23339);
xor U23417 (N_23417,N_23308,N_23394);
nor U23418 (N_23418,N_23313,N_23212);
nor U23419 (N_23419,N_23242,N_23186);
or U23420 (N_23420,N_23392,N_23257);
xor U23421 (N_23421,N_23143,N_23173);
nand U23422 (N_23422,N_23205,N_23307);
and U23423 (N_23423,N_23170,N_23200);
xnor U23424 (N_23424,N_23145,N_23167);
xor U23425 (N_23425,N_23383,N_23367);
and U23426 (N_23426,N_23311,N_23235);
and U23427 (N_23427,N_23139,N_23151);
and U23428 (N_23428,N_23246,N_23127);
nand U23429 (N_23429,N_23169,N_23253);
and U23430 (N_23430,N_23211,N_23349);
nor U23431 (N_23431,N_23163,N_23260);
nand U23432 (N_23432,N_23126,N_23198);
or U23433 (N_23433,N_23189,N_23110);
nor U23434 (N_23434,N_23237,N_23280);
or U23435 (N_23435,N_23301,N_23363);
or U23436 (N_23436,N_23334,N_23319);
xnor U23437 (N_23437,N_23354,N_23346);
nor U23438 (N_23438,N_23174,N_23284);
nand U23439 (N_23439,N_23149,N_23382);
nor U23440 (N_23440,N_23111,N_23210);
xor U23441 (N_23441,N_23344,N_23310);
xnor U23442 (N_23442,N_23222,N_23241);
xnor U23443 (N_23443,N_23254,N_23296);
and U23444 (N_23444,N_23160,N_23350);
and U23445 (N_23445,N_23276,N_23259);
nor U23446 (N_23446,N_23196,N_23214);
xnor U23447 (N_23447,N_23152,N_23266);
and U23448 (N_23448,N_23336,N_23236);
nor U23449 (N_23449,N_23378,N_23396);
nand U23450 (N_23450,N_23220,N_23289);
xor U23451 (N_23451,N_23180,N_23226);
or U23452 (N_23452,N_23154,N_23326);
nand U23453 (N_23453,N_23399,N_23223);
nand U23454 (N_23454,N_23285,N_23251);
and U23455 (N_23455,N_23391,N_23373);
and U23456 (N_23456,N_23395,N_23352);
or U23457 (N_23457,N_23328,N_23318);
xnor U23458 (N_23458,N_23314,N_23356);
and U23459 (N_23459,N_23106,N_23309);
and U23460 (N_23460,N_23155,N_23130);
or U23461 (N_23461,N_23217,N_23172);
or U23462 (N_23462,N_23287,N_23142);
xor U23463 (N_23463,N_23338,N_23122);
nand U23464 (N_23464,N_23113,N_23381);
and U23465 (N_23465,N_23162,N_23333);
nand U23466 (N_23466,N_23204,N_23393);
nor U23467 (N_23467,N_23277,N_23137);
xor U23468 (N_23468,N_23267,N_23201);
nand U23469 (N_23469,N_23207,N_23138);
and U23470 (N_23470,N_23182,N_23215);
and U23471 (N_23471,N_23337,N_23181);
nand U23472 (N_23472,N_23305,N_23332);
and U23473 (N_23473,N_23195,N_23190);
xor U23474 (N_23474,N_23238,N_23366);
or U23475 (N_23475,N_23250,N_23258);
or U23476 (N_23476,N_23295,N_23321);
and U23477 (N_23477,N_23304,N_23281);
and U23478 (N_23478,N_23398,N_23369);
nor U23479 (N_23479,N_23379,N_23168);
nand U23480 (N_23480,N_23179,N_23191);
xor U23481 (N_23481,N_23324,N_23178);
nor U23482 (N_23482,N_23194,N_23146);
nor U23483 (N_23483,N_23225,N_23109);
and U23484 (N_23484,N_23107,N_23302);
and U23485 (N_23485,N_23329,N_23124);
nor U23486 (N_23486,N_23119,N_23244);
nor U23487 (N_23487,N_23218,N_23252);
nand U23488 (N_23488,N_23219,N_23262);
nor U23489 (N_23489,N_23264,N_23274);
or U23490 (N_23490,N_23131,N_23340);
xnor U23491 (N_23491,N_23213,N_23231);
and U23492 (N_23492,N_23273,N_23105);
nand U23493 (N_23493,N_23271,N_23125);
nor U23494 (N_23494,N_23232,N_23345);
nor U23495 (N_23495,N_23157,N_23123);
or U23496 (N_23496,N_23323,N_23193);
xnor U23497 (N_23497,N_23279,N_23135);
nand U23498 (N_23498,N_23115,N_23114);
nor U23499 (N_23499,N_23306,N_23233);
xnor U23500 (N_23500,N_23288,N_23188);
nand U23501 (N_23501,N_23300,N_23385);
nor U23502 (N_23502,N_23368,N_23322);
xor U23503 (N_23503,N_23245,N_23372);
or U23504 (N_23504,N_23208,N_23298);
xor U23505 (N_23505,N_23156,N_23390);
and U23506 (N_23506,N_23282,N_23227);
nand U23507 (N_23507,N_23240,N_23101);
and U23508 (N_23508,N_23102,N_23317);
nand U23509 (N_23509,N_23256,N_23270);
and U23510 (N_23510,N_23221,N_23360);
xor U23511 (N_23511,N_23159,N_23161);
and U23512 (N_23512,N_23320,N_23355);
xor U23513 (N_23513,N_23128,N_23183);
nor U23514 (N_23514,N_23150,N_23342);
nor U23515 (N_23515,N_23299,N_23224);
xnor U23516 (N_23516,N_23348,N_23377);
xor U23517 (N_23517,N_23175,N_23315);
or U23518 (N_23518,N_23388,N_23364);
xor U23519 (N_23519,N_23327,N_23247);
xnor U23520 (N_23520,N_23303,N_23120);
and U23521 (N_23521,N_23216,N_23129);
nor U23522 (N_23522,N_23206,N_23376);
nor U23523 (N_23523,N_23362,N_23209);
and U23524 (N_23524,N_23359,N_23353);
nand U23525 (N_23525,N_23199,N_23292);
nor U23526 (N_23526,N_23255,N_23144);
nor U23527 (N_23527,N_23341,N_23118);
nand U23528 (N_23528,N_23347,N_23330);
nor U23529 (N_23529,N_23389,N_23386);
nand U23530 (N_23530,N_23294,N_23261);
nand U23531 (N_23531,N_23249,N_23153);
and U23532 (N_23532,N_23229,N_23365);
and U23533 (N_23533,N_23134,N_23140);
xnor U23534 (N_23534,N_23132,N_23117);
xor U23535 (N_23535,N_23147,N_23275);
nand U23536 (N_23536,N_23187,N_23166);
and U23537 (N_23537,N_23397,N_23116);
xnor U23538 (N_23538,N_23133,N_23148);
and U23539 (N_23539,N_23164,N_23234);
nand U23540 (N_23540,N_23263,N_23384);
nor U23541 (N_23541,N_23371,N_23165);
nor U23542 (N_23542,N_23100,N_23171);
or U23543 (N_23543,N_23230,N_23283);
nor U23544 (N_23544,N_23108,N_23103);
nand U23545 (N_23545,N_23312,N_23184);
nor U23546 (N_23546,N_23293,N_23278);
or U23547 (N_23547,N_23176,N_23185);
nor U23548 (N_23548,N_23387,N_23335);
xor U23549 (N_23549,N_23141,N_23202);
and U23550 (N_23550,N_23139,N_23258);
nor U23551 (N_23551,N_23295,N_23115);
nand U23552 (N_23552,N_23275,N_23177);
nor U23553 (N_23553,N_23381,N_23239);
nor U23554 (N_23554,N_23269,N_23195);
and U23555 (N_23555,N_23302,N_23339);
nor U23556 (N_23556,N_23116,N_23321);
nor U23557 (N_23557,N_23157,N_23140);
or U23558 (N_23558,N_23314,N_23150);
or U23559 (N_23559,N_23174,N_23163);
and U23560 (N_23560,N_23204,N_23146);
or U23561 (N_23561,N_23142,N_23199);
nand U23562 (N_23562,N_23293,N_23272);
and U23563 (N_23563,N_23227,N_23329);
xor U23564 (N_23564,N_23164,N_23110);
or U23565 (N_23565,N_23241,N_23391);
nand U23566 (N_23566,N_23335,N_23141);
and U23567 (N_23567,N_23369,N_23197);
xor U23568 (N_23568,N_23382,N_23244);
nand U23569 (N_23569,N_23186,N_23382);
nand U23570 (N_23570,N_23174,N_23188);
or U23571 (N_23571,N_23337,N_23216);
xnor U23572 (N_23572,N_23285,N_23103);
xor U23573 (N_23573,N_23328,N_23134);
nor U23574 (N_23574,N_23323,N_23139);
and U23575 (N_23575,N_23358,N_23381);
and U23576 (N_23576,N_23368,N_23115);
nor U23577 (N_23577,N_23181,N_23343);
nand U23578 (N_23578,N_23182,N_23201);
and U23579 (N_23579,N_23351,N_23187);
nor U23580 (N_23580,N_23121,N_23207);
nand U23581 (N_23581,N_23265,N_23337);
nand U23582 (N_23582,N_23296,N_23152);
and U23583 (N_23583,N_23212,N_23255);
xnor U23584 (N_23584,N_23261,N_23127);
nor U23585 (N_23585,N_23361,N_23324);
nor U23586 (N_23586,N_23150,N_23369);
nor U23587 (N_23587,N_23303,N_23341);
nand U23588 (N_23588,N_23296,N_23330);
and U23589 (N_23589,N_23283,N_23126);
nor U23590 (N_23590,N_23343,N_23272);
xor U23591 (N_23591,N_23385,N_23180);
and U23592 (N_23592,N_23255,N_23233);
nor U23593 (N_23593,N_23292,N_23373);
nor U23594 (N_23594,N_23335,N_23346);
nand U23595 (N_23595,N_23374,N_23199);
or U23596 (N_23596,N_23161,N_23235);
and U23597 (N_23597,N_23309,N_23128);
nor U23598 (N_23598,N_23223,N_23135);
nor U23599 (N_23599,N_23310,N_23140);
nor U23600 (N_23600,N_23283,N_23181);
xnor U23601 (N_23601,N_23202,N_23110);
nor U23602 (N_23602,N_23385,N_23264);
nor U23603 (N_23603,N_23126,N_23337);
nor U23604 (N_23604,N_23392,N_23147);
or U23605 (N_23605,N_23323,N_23303);
or U23606 (N_23606,N_23368,N_23117);
and U23607 (N_23607,N_23130,N_23246);
or U23608 (N_23608,N_23347,N_23154);
and U23609 (N_23609,N_23122,N_23253);
and U23610 (N_23610,N_23259,N_23122);
nand U23611 (N_23611,N_23104,N_23293);
nand U23612 (N_23612,N_23217,N_23215);
and U23613 (N_23613,N_23210,N_23130);
xor U23614 (N_23614,N_23220,N_23122);
nor U23615 (N_23615,N_23203,N_23281);
xnor U23616 (N_23616,N_23363,N_23332);
or U23617 (N_23617,N_23279,N_23116);
xnor U23618 (N_23618,N_23378,N_23373);
nand U23619 (N_23619,N_23360,N_23158);
or U23620 (N_23620,N_23326,N_23103);
nor U23621 (N_23621,N_23134,N_23301);
xor U23622 (N_23622,N_23275,N_23392);
and U23623 (N_23623,N_23242,N_23340);
or U23624 (N_23624,N_23298,N_23234);
xnor U23625 (N_23625,N_23209,N_23264);
and U23626 (N_23626,N_23360,N_23288);
and U23627 (N_23627,N_23165,N_23261);
and U23628 (N_23628,N_23196,N_23392);
and U23629 (N_23629,N_23337,N_23253);
and U23630 (N_23630,N_23147,N_23360);
nand U23631 (N_23631,N_23270,N_23319);
nor U23632 (N_23632,N_23213,N_23286);
and U23633 (N_23633,N_23164,N_23190);
or U23634 (N_23634,N_23291,N_23113);
xor U23635 (N_23635,N_23278,N_23167);
xor U23636 (N_23636,N_23141,N_23111);
nand U23637 (N_23637,N_23197,N_23378);
xnor U23638 (N_23638,N_23202,N_23337);
and U23639 (N_23639,N_23345,N_23284);
xnor U23640 (N_23640,N_23234,N_23374);
xor U23641 (N_23641,N_23368,N_23304);
nand U23642 (N_23642,N_23183,N_23323);
xnor U23643 (N_23643,N_23242,N_23381);
or U23644 (N_23644,N_23294,N_23104);
nand U23645 (N_23645,N_23200,N_23224);
nor U23646 (N_23646,N_23379,N_23132);
nor U23647 (N_23647,N_23198,N_23145);
or U23648 (N_23648,N_23364,N_23181);
or U23649 (N_23649,N_23182,N_23234);
nand U23650 (N_23650,N_23211,N_23289);
xor U23651 (N_23651,N_23310,N_23184);
and U23652 (N_23652,N_23117,N_23309);
or U23653 (N_23653,N_23147,N_23140);
nand U23654 (N_23654,N_23327,N_23113);
or U23655 (N_23655,N_23329,N_23396);
nand U23656 (N_23656,N_23122,N_23245);
nand U23657 (N_23657,N_23366,N_23290);
and U23658 (N_23658,N_23223,N_23341);
nand U23659 (N_23659,N_23175,N_23114);
nor U23660 (N_23660,N_23167,N_23251);
nand U23661 (N_23661,N_23387,N_23158);
nor U23662 (N_23662,N_23279,N_23167);
nor U23663 (N_23663,N_23395,N_23131);
nor U23664 (N_23664,N_23328,N_23289);
xnor U23665 (N_23665,N_23158,N_23103);
and U23666 (N_23666,N_23110,N_23185);
nand U23667 (N_23667,N_23329,N_23226);
nor U23668 (N_23668,N_23116,N_23395);
or U23669 (N_23669,N_23345,N_23177);
or U23670 (N_23670,N_23140,N_23197);
and U23671 (N_23671,N_23213,N_23118);
nor U23672 (N_23672,N_23182,N_23250);
and U23673 (N_23673,N_23321,N_23177);
nor U23674 (N_23674,N_23377,N_23235);
nor U23675 (N_23675,N_23196,N_23127);
xnor U23676 (N_23676,N_23385,N_23374);
xor U23677 (N_23677,N_23246,N_23311);
nand U23678 (N_23678,N_23321,N_23194);
xnor U23679 (N_23679,N_23225,N_23391);
and U23680 (N_23680,N_23156,N_23323);
nand U23681 (N_23681,N_23299,N_23264);
nor U23682 (N_23682,N_23187,N_23392);
nor U23683 (N_23683,N_23111,N_23311);
and U23684 (N_23684,N_23336,N_23191);
nor U23685 (N_23685,N_23223,N_23209);
nand U23686 (N_23686,N_23245,N_23271);
nand U23687 (N_23687,N_23196,N_23136);
xnor U23688 (N_23688,N_23325,N_23289);
and U23689 (N_23689,N_23292,N_23164);
nand U23690 (N_23690,N_23243,N_23269);
xnor U23691 (N_23691,N_23396,N_23323);
xor U23692 (N_23692,N_23377,N_23257);
nand U23693 (N_23693,N_23381,N_23225);
nor U23694 (N_23694,N_23311,N_23268);
or U23695 (N_23695,N_23189,N_23315);
xnor U23696 (N_23696,N_23388,N_23133);
xnor U23697 (N_23697,N_23113,N_23282);
and U23698 (N_23698,N_23207,N_23338);
xnor U23699 (N_23699,N_23311,N_23121);
nand U23700 (N_23700,N_23669,N_23584);
or U23701 (N_23701,N_23526,N_23574);
and U23702 (N_23702,N_23514,N_23573);
nor U23703 (N_23703,N_23458,N_23529);
xor U23704 (N_23704,N_23568,N_23619);
nand U23705 (N_23705,N_23682,N_23400);
and U23706 (N_23706,N_23547,N_23549);
nand U23707 (N_23707,N_23532,N_23634);
nor U23708 (N_23708,N_23658,N_23615);
xnor U23709 (N_23709,N_23531,N_23425);
nor U23710 (N_23710,N_23606,N_23626);
nor U23711 (N_23711,N_23578,N_23496);
or U23712 (N_23712,N_23510,N_23672);
xor U23713 (N_23713,N_23689,N_23567);
nor U23714 (N_23714,N_23404,N_23687);
nand U23715 (N_23715,N_23632,N_23685);
and U23716 (N_23716,N_23644,N_23421);
nor U23717 (N_23717,N_23412,N_23469);
and U23718 (N_23718,N_23663,N_23671);
xor U23719 (N_23719,N_23661,N_23419);
nand U23720 (N_23720,N_23456,N_23442);
nand U23721 (N_23721,N_23471,N_23544);
nand U23722 (N_23722,N_23603,N_23478);
xnor U23723 (N_23723,N_23543,N_23409);
nor U23724 (N_23724,N_23487,N_23569);
or U23725 (N_23725,N_23534,N_23683);
xor U23726 (N_23726,N_23556,N_23473);
and U23727 (N_23727,N_23472,N_23608);
and U23728 (N_23728,N_23620,N_23630);
or U23729 (N_23729,N_23449,N_23485);
xor U23730 (N_23730,N_23506,N_23403);
or U23731 (N_23731,N_23596,N_23503);
and U23732 (N_23732,N_23410,N_23509);
nor U23733 (N_23733,N_23560,N_23686);
or U23734 (N_23734,N_23646,N_23435);
nand U23735 (N_23735,N_23645,N_23538);
xor U23736 (N_23736,N_23428,N_23657);
xor U23737 (N_23737,N_23414,N_23426);
nand U23738 (N_23738,N_23495,N_23621);
xnor U23739 (N_23739,N_23464,N_23440);
and U23740 (N_23740,N_23612,N_23670);
and U23741 (N_23741,N_23515,N_23443);
and U23742 (N_23742,N_23470,N_23633);
nand U23743 (N_23743,N_23447,N_23659);
nand U23744 (N_23744,N_23548,N_23642);
and U23745 (N_23745,N_23500,N_23511);
or U23746 (N_23746,N_23656,N_23616);
nor U23747 (N_23747,N_23681,N_23519);
xnor U23748 (N_23748,N_23488,N_23591);
nand U23749 (N_23749,N_23589,N_23635);
nor U23750 (N_23750,N_23597,N_23627);
or U23751 (N_23751,N_23486,N_23406);
xor U23752 (N_23752,N_23451,N_23494);
xnor U23753 (N_23753,N_23434,N_23655);
or U23754 (N_23754,N_23674,N_23609);
xor U23755 (N_23755,N_23423,N_23680);
nor U23756 (N_23756,N_23628,N_23643);
and U23757 (N_23757,N_23459,N_23429);
xor U23758 (N_23758,N_23542,N_23594);
nor U23759 (N_23759,N_23629,N_23614);
xor U23760 (N_23760,N_23579,N_23582);
nor U23761 (N_23761,N_23483,N_23581);
nand U23762 (N_23762,N_23557,N_23554);
xnor U23763 (N_23763,N_23453,N_23572);
and U23764 (N_23764,N_23516,N_23651);
nand U23765 (N_23765,N_23518,N_23610);
and U23766 (N_23766,N_23507,N_23580);
and U23767 (N_23767,N_23536,N_23601);
or U23768 (N_23768,N_23576,N_23438);
xor U23769 (N_23769,N_23521,N_23690);
nor U23770 (N_23770,N_23537,N_23545);
xnor U23771 (N_23771,N_23679,N_23476);
xor U23772 (N_23772,N_23617,N_23505);
nor U23773 (N_23773,N_23437,N_23457);
xnor U23774 (N_23774,N_23401,N_23513);
nand U23775 (N_23775,N_23698,N_23420);
nand U23776 (N_23776,N_23415,N_23583);
or U23777 (N_23777,N_23636,N_23413);
xor U23778 (N_23778,N_23575,N_23402);
nand U23779 (N_23779,N_23431,N_23462);
xor U23780 (N_23780,N_23558,N_23481);
nand U23781 (N_23781,N_23696,N_23436);
and U23782 (N_23782,N_23502,N_23444);
nor U23783 (N_23783,N_23571,N_23525);
xor U23784 (N_23784,N_23650,N_23699);
nand U23785 (N_23785,N_23607,N_23647);
nor U23786 (N_23786,N_23664,N_23605);
nor U23787 (N_23787,N_23676,N_23416);
and U23788 (N_23788,N_23551,N_23499);
xnor U23789 (N_23789,N_23504,N_23563);
nand U23790 (N_23790,N_23463,N_23535);
and U23791 (N_23791,N_23695,N_23441);
xnor U23792 (N_23792,N_23520,N_23477);
nor U23793 (N_23793,N_23692,N_23562);
or U23794 (N_23794,N_23565,N_23461);
nand U23795 (N_23795,N_23446,N_23675);
nand U23796 (N_23796,N_23524,N_23455);
nor U23797 (N_23797,N_23624,N_23587);
or U23798 (N_23798,N_23673,N_23522);
xor U23799 (N_23799,N_23640,N_23490);
nand U23800 (N_23800,N_23595,N_23497);
xnor U23801 (N_23801,N_23475,N_23454);
xor U23802 (N_23802,N_23652,N_23540);
nand U23803 (N_23803,N_23460,N_23561);
nor U23804 (N_23804,N_23598,N_23489);
nor U23805 (N_23805,N_23622,N_23508);
and U23806 (N_23806,N_23492,N_23694);
nand U23807 (N_23807,N_23452,N_23604);
nand U23808 (N_23808,N_23530,N_23450);
and U23809 (N_23809,N_23611,N_23411);
or U23810 (N_23810,N_23592,N_23527);
and U23811 (N_23811,N_23528,N_23566);
nand U23812 (N_23812,N_23641,N_23448);
and U23813 (N_23813,N_23480,N_23466);
xnor U23814 (N_23814,N_23407,N_23555);
nor U23815 (N_23815,N_23427,N_23599);
or U23816 (N_23816,N_23465,N_23593);
xor U23817 (N_23817,N_23418,N_23552);
and U23818 (N_23818,N_23662,N_23533);
xor U23819 (N_23819,N_23445,N_23653);
nor U23820 (N_23820,N_23479,N_23631);
and U23821 (N_23821,N_23590,N_23660);
and U23822 (N_23822,N_23550,N_23498);
and U23823 (N_23823,N_23439,N_23546);
nor U23824 (N_23824,N_23678,N_23405);
nor U23825 (N_23825,N_23417,N_23433);
and U23826 (N_23826,N_23408,N_23613);
nor U23827 (N_23827,N_23625,N_23570);
or U23828 (N_23828,N_23484,N_23693);
and U23829 (N_23829,N_23517,N_23654);
nand U23830 (N_23830,N_23577,N_23422);
xor U23831 (N_23831,N_23665,N_23585);
nand U23832 (N_23832,N_23677,N_23623);
xor U23833 (N_23833,N_23424,N_23668);
and U23834 (N_23834,N_23649,N_23697);
or U23835 (N_23835,N_23467,N_23553);
or U23836 (N_23836,N_23684,N_23688);
nand U23837 (N_23837,N_23602,N_23474);
nor U23838 (N_23838,N_23618,N_23639);
nor U23839 (N_23839,N_23468,N_23586);
and U23840 (N_23840,N_23648,N_23667);
and U23841 (N_23841,N_23637,N_23482);
or U23842 (N_23842,N_23430,N_23638);
and U23843 (N_23843,N_23564,N_23491);
and U23844 (N_23844,N_23666,N_23588);
or U23845 (N_23845,N_23691,N_23493);
and U23846 (N_23846,N_23432,N_23600);
and U23847 (N_23847,N_23523,N_23559);
nor U23848 (N_23848,N_23512,N_23539);
and U23849 (N_23849,N_23501,N_23541);
nand U23850 (N_23850,N_23511,N_23680);
nand U23851 (N_23851,N_23677,N_23574);
nand U23852 (N_23852,N_23411,N_23598);
and U23853 (N_23853,N_23576,N_23631);
or U23854 (N_23854,N_23605,N_23442);
nand U23855 (N_23855,N_23640,N_23521);
or U23856 (N_23856,N_23411,N_23579);
nor U23857 (N_23857,N_23642,N_23535);
xor U23858 (N_23858,N_23466,N_23441);
nor U23859 (N_23859,N_23685,N_23583);
nand U23860 (N_23860,N_23569,N_23441);
nand U23861 (N_23861,N_23424,N_23452);
nand U23862 (N_23862,N_23442,N_23487);
and U23863 (N_23863,N_23660,N_23656);
nor U23864 (N_23864,N_23448,N_23687);
or U23865 (N_23865,N_23430,N_23667);
and U23866 (N_23866,N_23635,N_23685);
nand U23867 (N_23867,N_23575,N_23498);
xnor U23868 (N_23868,N_23631,N_23535);
or U23869 (N_23869,N_23467,N_23691);
nor U23870 (N_23870,N_23532,N_23418);
nand U23871 (N_23871,N_23488,N_23611);
nor U23872 (N_23872,N_23690,N_23447);
or U23873 (N_23873,N_23467,N_23502);
xor U23874 (N_23874,N_23424,N_23608);
or U23875 (N_23875,N_23549,N_23490);
nor U23876 (N_23876,N_23428,N_23599);
and U23877 (N_23877,N_23658,N_23438);
or U23878 (N_23878,N_23564,N_23469);
and U23879 (N_23879,N_23566,N_23485);
and U23880 (N_23880,N_23410,N_23565);
nand U23881 (N_23881,N_23567,N_23524);
nand U23882 (N_23882,N_23672,N_23631);
nor U23883 (N_23883,N_23684,N_23653);
nand U23884 (N_23884,N_23556,N_23634);
xor U23885 (N_23885,N_23593,N_23405);
xor U23886 (N_23886,N_23613,N_23524);
and U23887 (N_23887,N_23688,N_23463);
nor U23888 (N_23888,N_23424,N_23599);
nor U23889 (N_23889,N_23457,N_23444);
or U23890 (N_23890,N_23441,N_23624);
xor U23891 (N_23891,N_23659,N_23637);
xnor U23892 (N_23892,N_23605,N_23597);
nand U23893 (N_23893,N_23609,N_23400);
or U23894 (N_23894,N_23474,N_23619);
nand U23895 (N_23895,N_23621,N_23559);
xnor U23896 (N_23896,N_23425,N_23505);
xnor U23897 (N_23897,N_23637,N_23653);
xor U23898 (N_23898,N_23622,N_23497);
nand U23899 (N_23899,N_23513,N_23403);
xnor U23900 (N_23900,N_23428,N_23677);
xnor U23901 (N_23901,N_23582,N_23613);
or U23902 (N_23902,N_23697,N_23541);
nor U23903 (N_23903,N_23496,N_23685);
or U23904 (N_23904,N_23696,N_23577);
xnor U23905 (N_23905,N_23537,N_23655);
and U23906 (N_23906,N_23614,N_23504);
nor U23907 (N_23907,N_23522,N_23473);
or U23908 (N_23908,N_23637,N_23516);
nor U23909 (N_23909,N_23449,N_23400);
nand U23910 (N_23910,N_23556,N_23439);
nor U23911 (N_23911,N_23609,N_23415);
and U23912 (N_23912,N_23520,N_23469);
and U23913 (N_23913,N_23567,N_23451);
or U23914 (N_23914,N_23405,N_23565);
or U23915 (N_23915,N_23402,N_23621);
or U23916 (N_23916,N_23543,N_23490);
xnor U23917 (N_23917,N_23526,N_23444);
xor U23918 (N_23918,N_23440,N_23638);
and U23919 (N_23919,N_23636,N_23446);
and U23920 (N_23920,N_23463,N_23573);
or U23921 (N_23921,N_23682,N_23491);
nand U23922 (N_23922,N_23491,N_23483);
or U23923 (N_23923,N_23475,N_23543);
nand U23924 (N_23924,N_23552,N_23485);
nor U23925 (N_23925,N_23567,N_23656);
and U23926 (N_23926,N_23626,N_23657);
and U23927 (N_23927,N_23688,N_23443);
and U23928 (N_23928,N_23459,N_23625);
nand U23929 (N_23929,N_23478,N_23529);
xnor U23930 (N_23930,N_23444,N_23567);
nand U23931 (N_23931,N_23417,N_23533);
nor U23932 (N_23932,N_23578,N_23611);
nand U23933 (N_23933,N_23678,N_23559);
or U23934 (N_23934,N_23668,N_23562);
and U23935 (N_23935,N_23609,N_23529);
xor U23936 (N_23936,N_23697,N_23569);
nor U23937 (N_23937,N_23499,N_23659);
nor U23938 (N_23938,N_23519,N_23625);
or U23939 (N_23939,N_23618,N_23603);
or U23940 (N_23940,N_23570,N_23626);
nor U23941 (N_23941,N_23404,N_23639);
and U23942 (N_23942,N_23442,N_23424);
and U23943 (N_23943,N_23475,N_23638);
or U23944 (N_23944,N_23551,N_23603);
and U23945 (N_23945,N_23510,N_23689);
or U23946 (N_23946,N_23677,N_23583);
nand U23947 (N_23947,N_23578,N_23401);
or U23948 (N_23948,N_23476,N_23442);
nand U23949 (N_23949,N_23631,N_23533);
or U23950 (N_23950,N_23594,N_23690);
and U23951 (N_23951,N_23572,N_23439);
and U23952 (N_23952,N_23569,N_23664);
or U23953 (N_23953,N_23687,N_23677);
or U23954 (N_23954,N_23484,N_23559);
xor U23955 (N_23955,N_23501,N_23638);
and U23956 (N_23956,N_23478,N_23669);
and U23957 (N_23957,N_23472,N_23488);
nand U23958 (N_23958,N_23637,N_23527);
nand U23959 (N_23959,N_23479,N_23550);
nand U23960 (N_23960,N_23670,N_23632);
nor U23961 (N_23961,N_23541,N_23602);
or U23962 (N_23962,N_23470,N_23408);
nor U23963 (N_23963,N_23539,N_23466);
and U23964 (N_23964,N_23471,N_23482);
or U23965 (N_23965,N_23594,N_23645);
or U23966 (N_23966,N_23653,N_23572);
xnor U23967 (N_23967,N_23599,N_23558);
and U23968 (N_23968,N_23491,N_23460);
nor U23969 (N_23969,N_23505,N_23578);
nand U23970 (N_23970,N_23661,N_23589);
nor U23971 (N_23971,N_23564,N_23508);
or U23972 (N_23972,N_23668,N_23468);
nor U23973 (N_23973,N_23644,N_23691);
nor U23974 (N_23974,N_23477,N_23671);
and U23975 (N_23975,N_23514,N_23576);
and U23976 (N_23976,N_23580,N_23626);
and U23977 (N_23977,N_23682,N_23647);
nand U23978 (N_23978,N_23419,N_23547);
xor U23979 (N_23979,N_23547,N_23578);
nor U23980 (N_23980,N_23415,N_23645);
xnor U23981 (N_23981,N_23661,N_23663);
nand U23982 (N_23982,N_23665,N_23434);
xnor U23983 (N_23983,N_23472,N_23652);
or U23984 (N_23984,N_23544,N_23626);
nor U23985 (N_23985,N_23457,N_23433);
xor U23986 (N_23986,N_23453,N_23401);
xor U23987 (N_23987,N_23525,N_23547);
and U23988 (N_23988,N_23471,N_23666);
nand U23989 (N_23989,N_23677,N_23542);
nand U23990 (N_23990,N_23688,N_23403);
xor U23991 (N_23991,N_23512,N_23622);
or U23992 (N_23992,N_23403,N_23481);
xnor U23993 (N_23993,N_23681,N_23545);
nor U23994 (N_23994,N_23596,N_23436);
nor U23995 (N_23995,N_23444,N_23462);
and U23996 (N_23996,N_23420,N_23638);
xnor U23997 (N_23997,N_23527,N_23426);
nor U23998 (N_23998,N_23595,N_23420);
xor U23999 (N_23999,N_23666,N_23614);
and U24000 (N_24000,N_23819,N_23786);
or U24001 (N_24001,N_23937,N_23709);
nor U24002 (N_24002,N_23813,N_23815);
and U24003 (N_24003,N_23993,N_23836);
nor U24004 (N_24004,N_23857,N_23715);
and U24005 (N_24005,N_23753,N_23979);
xnor U24006 (N_24006,N_23833,N_23773);
xor U24007 (N_24007,N_23822,N_23884);
or U24008 (N_24008,N_23821,N_23835);
nand U24009 (N_24009,N_23919,N_23917);
nor U24010 (N_24010,N_23708,N_23714);
nand U24011 (N_24011,N_23970,N_23814);
nand U24012 (N_24012,N_23781,N_23712);
nor U24013 (N_24013,N_23971,N_23905);
nand U24014 (N_24014,N_23757,N_23872);
nand U24015 (N_24015,N_23855,N_23901);
nor U24016 (N_24016,N_23796,N_23774);
and U24017 (N_24017,N_23903,N_23828);
or U24018 (N_24018,N_23939,N_23703);
nand U24019 (N_24019,N_23930,N_23824);
xor U24020 (N_24020,N_23826,N_23870);
and U24021 (N_24021,N_23910,N_23951);
and U24022 (N_24022,N_23927,N_23888);
and U24023 (N_24023,N_23705,N_23793);
nor U24024 (N_24024,N_23916,N_23854);
and U24025 (N_24025,N_23876,N_23874);
nor U24026 (N_24026,N_23920,N_23850);
xor U24027 (N_24027,N_23984,N_23805);
or U24028 (N_24028,N_23952,N_23840);
nand U24029 (N_24029,N_23767,N_23856);
and U24030 (N_24030,N_23766,N_23871);
nor U24031 (N_24031,N_23740,N_23889);
or U24032 (N_24032,N_23776,N_23724);
xnor U24033 (N_24033,N_23769,N_23780);
xor U24034 (N_24034,N_23926,N_23700);
and U24035 (N_24035,N_23990,N_23895);
and U24036 (N_24036,N_23862,N_23883);
nand U24037 (N_24037,N_23987,N_23898);
or U24038 (N_24038,N_23710,N_23974);
or U24039 (N_24039,N_23754,N_23839);
or U24040 (N_24040,N_23962,N_23750);
nand U24041 (N_24041,N_23906,N_23860);
xor U24042 (N_24042,N_23879,N_23795);
nor U24043 (N_24043,N_23789,N_23823);
nand U24044 (N_24044,N_23859,N_23798);
and U24045 (N_24045,N_23999,N_23932);
nand U24046 (N_24046,N_23729,N_23950);
xor U24047 (N_24047,N_23954,N_23972);
nand U24048 (N_24048,N_23734,N_23717);
and U24049 (N_24049,N_23858,N_23790);
nand U24050 (N_24050,N_23845,N_23728);
nor U24051 (N_24051,N_23785,N_23985);
and U24052 (N_24052,N_23940,N_23763);
or U24053 (N_24053,N_23991,N_23912);
or U24054 (N_24054,N_23818,N_23816);
and U24055 (N_24055,N_23849,N_23820);
nor U24056 (N_24056,N_23738,N_23977);
nor U24057 (N_24057,N_23743,N_23961);
xor U24058 (N_24058,N_23936,N_23934);
or U24059 (N_24059,N_23944,N_23844);
and U24060 (N_24060,N_23810,N_23706);
nand U24061 (N_24061,N_23960,N_23865);
nor U24062 (N_24062,N_23739,N_23707);
xnor U24063 (N_24063,N_23748,N_23949);
xnor U24064 (N_24064,N_23878,N_23834);
or U24065 (N_24065,N_23908,N_23921);
nand U24066 (N_24066,N_23770,N_23959);
xnor U24067 (N_24067,N_23981,N_23782);
nor U24068 (N_24068,N_23742,N_23745);
nor U24069 (N_24069,N_23812,N_23722);
and U24070 (N_24070,N_23846,N_23827);
or U24071 (N_24071,N_23802,N_23966);
and U24072 (N_24072,N_23913,N_23777);
nor U24073 (N_24073,N_23877,N_23727);
nor U24074 (N_24074,N_23851,N_23807);
nand U24075 (N_24075,N_23825,N_23762);
nor U24076 (N_24076,N_23843,N_23914);
or U24077 (N_24077,N_23732,N_23736);
or U24078 (N_24078,N_23980,N_23829);
and U24079 (N_24079,N_23718,N_23783);
nor U24080 (N_24080,N_23923,N_23744);
and U24081 (N_24081,N_23969,N_23867);
and U24082 (N_24082,N_23830,N_23968);
nand U24083 (N_24083,N_23925,N_23842);
nor U24084 (N_24084,N_23702,N_23947);
nand U24085 (N_24085,N_23792,N_23994);
and U24086 (N_24086,N_23946,N_23978);
or U24087 (N_24087,N_23896,N_23933);
and U24088 (N_24088,N_23853,N_23806);
xnor U24089 (N_24089,N_23760,N_23751);
nor U24090 (N_24090,N_23887,N_23797);
xor U24091 (N_24091,N_23938,N_23869);
xor U24092 (N_24092,N_23801,N_23701);
nor U24093 (N_24093,N_23747,N_23746);
nand U24094 (N_24094,N_23873,N_23964);
nand U24095 (N_24095,N_23922,N_23953);
nand U24096 (N_24096,N_23880,N_23737);
nor U24097 (N_24097,N_23809,N_23899);
nor U24098 (N_24098,N_23749,N_23918);
or U24099 (N_24099,N_23931,N_23787);
nand U24100 (N_24100,N_23723,N_23988);
or U24101 (N_24101,N_23861,N_23758);
nor U24102 (N_24102,N_23771,N_23982);
nand U24103 (N_24103,N_23800,N_23995);
or U24104 (N_24104,N_23778,N_23764);
or U24105 (N_24105,N_23928,N_23721);
nand U24106 (N_24106,N_23892,N_23956);
nand U24107 (N_24107,N_23791,N_23719);
or U24108 (N_24108,N_23772,N_23756);
nand U24109 (N_24109,N_23866,N_23886);
xnor U24110 (N_24110,N_23831,N_23811);
nor U24111 (N_24111,N_23983,N_23929);
nand U24112 (N_24112,N_23837,N_23963);
or U24113 (N_24113,N_23752,N_23726);
and U24114 (N_24114,N_23881,N_23768);
and U24115 (N_24115,N_23967,N_23909);
nor U24116 (N_24116,N_23942,N_23882);
nand U24117 (N_24117,N_23848,N_23832);
or U24118 (N_24118,N_23894,N_23808);
xor U24119 (N_24119,N_23904,N_23817);
or U24120 (N_24120,N_23911,N_23875);
or U24121 (N_24121,N_23885,N_23711);
nor U24122 (N_24122,N_23868,N_23733);
and U24123 (N_24123,N_23976,N_23716);
nand U24124 (N_24124,N_23713,N_23863);
and U24125 (N_24125,N_23759,N_23945);
nor U24126 (N_24126,N_23890,N_23897);
nand U24127 (N_24127,N_23730,N_23948);
and U24128 (N_24128,N_23989,N_23847);
or U24129 (N_24129,N_23986,N_23997);
nor U24130 (N_24130,N_23841,N_23975);
xnor U24131 (N_24131,N_23891,N_23735);
or U24132 (N_24132,N_23996,N_23761);
nand U24133 (N_24133,N_23799,N_23704);
or U24134 (N_24134,N_23958,N_23924);
or U24135 (N_24135,N_23973,N_23965);
xnor U24136 (N_24136,N_23957,N_23852);
and U24137 (N_24137,N_23915,N_23941);
nor U24138 (N_24138,N_23992,N_23779);
xor U24139 (N_24139,N_23741,N_23907);
xor U24140 (N_24140,N_23720,N_23998);
or U24141 (N_24141,N_23803,N_23794);
xor U24142 (N_24142,N_23893,N_23838);
nor U24143 (N_24143,N_23955,N_23935);
or U24144 (N_24144,N_23788,N_23755);
nand U24145 (N_24145,N_23731,N_23725);
and U24146 (N_24146,N_23775,N_23900);
nor U24147 (N_24147,N_23864,N_23804);
nor U24148 (N_24148,N_23765,N_23943);
xor U24149 (N_24149,N_23784,N_23902);
and U24150 (N_24150,N_23772,N_23979);
or U24151 (N_24151,N_23838,N_23924);
nor U24152 (N_24152,N_23939,N_23729);
xor U24153 (N_24153,N_23766,N_23985);
nor U24154 (N_24154,N_23927,N_23846);
and U24155 (N_24155,N_23777,N_23976);
xnor U24156 (N_24156,N_23813,N_23772);
and U24157 (N_24157,N_23898,N_23965);
nor U24158 (N_24158,N_23812,N_23769);
nand U24159 (N_24159,N_23885,N_23909);
nand U24160 (N_24160,N_23838,N_23987);
nand U24161 (N_24161,N_23986,N_23926);
or U24162 (N_24162,N_23704,N_23713);
xor U24163 (N_24163,N_23817,N_23783);
or U24164 (N_24164,N_23790,N_23777);
nand U24165 (N_24165,N_23701,N_23749);
or U24166 (N_24166,N_23728,N_23759);
xnor U24167 (N_24167,N_23817,N_23885);
xnor U24168 (N_24168,N_23861,N_23713);
nand U24169 (N_24169,N_23862,N_23714);
or U24170 (N_24170,N_23841,N_23955);
or U24171 (N_24171,N_23919,N_23859);
nand U24172 (N_24172,N_23877,N_23816);
or U24173 (N_24173,N_23973,N_23707);
nor U24174 (N_24174,N_23906,N_23849);
nand U24175 (N_24175,N_23902,N_23831);
nand U24176 (N_24176,N_23807,N_23768);
nor U24177 (N_24177,N_23944,N_23946);
xor U24178 (N_24178,N_23768,N_23928);
nand U24179 (N_24179,N_23706,N_23790);
and U24180 (N_24180,N_23873,N_23909);
nor U24181 (N_24181,N_23935,N_23909);
xor U24182 (N_24182,N_23959,N_23853);
nand U24183 (N_24183,N_23952,N_23953);
xnor U24184 (N_24184,N_23998,N_23749);
nor U24185 (N_24185,N_23726,N_23858);
and U24186 (N_24186,N_23985,N_23825);
nand U24187 (N_24187,N_23875,N_23990);
or U24188 (N_24188,N_23901,N_23946);
and U24189 (N_24189,N_23785,N_23869);
nor U24190 (N_24190,N_23992,N_23723);
and U24191 (N_24191,N_23711,N_23888);
and U24192 (N_24192,N_23870,N_23835);
nor U24193 (N_24193,N_23815,N_23825);
nand U24194 (N_24194,N_23905,N_23805);
xor U24195 (N_24195,N_23817,N_23834);
nand U24196 (N_24196,N_23723,N_23995);
and U24197 (N_24197,N_23756,N_23820);
nand U24198 (N_24198,N_23867,N_23768);
nand U24199 (N_24199,N_23786,N_23923);
or U24200 (N_24200,N_23924,N_23836);
nand U24201 (N_24201,N_23808,N_23858);
or U24202 (N_24202,N_23840,N_23782);
nor U24203 (N_24203,N_23736,N_23730);
or U24204 (N_24204,N_23739,N_23741);
nor U24205 (N_24205,N_23813,N_23774);
xor U24206 (N_24206,N_23779,N_23835);
and U24207 (N_24207,N_23728,N_23902);
nand U24208 (N_24208,N_23827,N_23985);
xnor U24209 (N_24209,N_23775,N_23903);
or U24210 (N_24210,N_23943,N_23839);
or U24211 (N_24211,N_23746,N_23817);
and U24212 (N_24212,N_23891,N_23807);
nand U24213 (N_24213,N_23851,N_23908);
and U24214 (N_24214,N_23850,N_23782);
xnor U24215 (N_24215,N_23872,N_23860);
and U24216 (N_24216,N_23736,N_23762);
xnor U24217 (N_24217,N_23758,N_23723);
and U24218 (N_24218,N_23858,N_23995);
xor U24219 (N_24219,N_23848,N_23833);
and U24220 (N_24220,N_23891,N_23701);
and U24221 (N_24221,N_23871,N_23997);
and U24222 (N_24222,N_23800,N_23750);
xnor U24223 (N_24223,N_23786,N_23741);
and U24224 (N_24224,N_23759,N_23807);
nor U24225 (N_24225,N_23712,N_23973);
nor U24226 (N_24226,N_23766,N_23757);
xnor U24227 (N_24227,N_23753,N_23744);
nor U24228 (N_24228,N_23988,N_23892);
and U24229 (N_24229,N_23735,N_23970);
or U24230 (N_24230,N_23725,N_23931);
xnor U24231 (N_24231,N_23887,N_23878);
nand U24232 (N_24232,N_23960,N_23762);
xor U24233 (N_24233,N_23795,N_23709);
nand U24234 (N_24234,N_23724,N_23885);
nor U24235 (N_24235,N_23738,N_23959);
xor U24236 (N_24236,N_23836,N_23709);
or U24237 (N_24237,N_23860,N_23836);
nor U24238 (N_24238,N_23971,N_23997);
and U24239 (N_24239,N_23819,N_23856);
and U24240 (N_24240,N_23876,N_23802);
xnor U24241 (N_24241,N_23875,N_23822);
xnor U24242 (N_24242,N_23707,N_23873);
and U24243 (N_24243,N_23901,N_23930);
nand U24244 (N_24244,N_23901,N_23779);
xor U24245 (N_24245,N_23802,N_23875);
xor U24246 (N_24246,N_23714,N_23950);
xor U24247 (N_24247,N_23736,N_23779);
nor U24248 (N_24248,N_23865,N_23896);
nand U24249 (N_24249,N_23742,N_23717);
or U24250 (N_24250,N_23900,N_23968);
xnor U24251 (N_24251,N_23800,N_23862);
or U24252 (N_24252,N_23776,N_23779);
or U24253 (N_24253,N_23970,N_23810);
xor U24254 (N_24254,N_23744,N_23946);
xnor U24255 (N_24255,N_23839,N_23808);
xor U24256 (N_24256,N_23850,N_23795);
and U24257 (N_24257,N_23731,N_23802);
nand U24258 (N_24258,N_23937,N_23824);
and U24259 (N_24259,N_23863,N_23810);
nor U24260 (N_24260,N_23791,N_23787);
or U24261 (N_24261,N_23710,N_23789);
or U24262 (N_24262,N_23851,N_23823);
nor U24263 (N_24263,N_23981,N_23933);
nor U24264 (N_24264,N_23924,N_23912);
xnor U24265 (N_24265,N_23978,N_23711);
nor U24266 (N_24266,N_23887,N_23739);
and U24267 (N_24267,N_23778,N_23892);
or U24268 (N_24268,N_23850,N_23845);
and U24269 (N_24269,N_23846,N_23881);
and U24270 (N_24270,N_23922,N_23968);
xor U24271 (N_24271,N_23741,N_23740);
nand U24272 (N_24272,N_23711,N_23730);
nor U24273 (N_24273,N_23905,N_23874);
nand U24274 (N_24274,N_23943,N_23998);
xnor U24275 (N_24275,N_23993,N_23743);
nor U24276 (N_24276,N_23894,N_23780);
nand U24277 (N_24277,N_23853,N_23701);
or U24278 (N_24278,N_23958,N_23841);
xor U24279 (N_24279,N_23725,N_23735);
nor U24280 (N_24280,N_23797,N_23763);
and U24281 (N_24281,N_23809,N_23790);
xnor U24282 (N_24282,N_23815,N_23976);
xnor U24283 (N_24283,N_23705,N_23903);
or U24284 (N_24284,N_23921,N_23929);
or U24285 (N_24285,N_23814,N_23815);
nor U24286 (N_24286,N_23980,N_23866);
and U24287 (N_24287,N_23753,N_23997);
xnor U24288 (N_24288,N_23874,N_23760);
nand U24289 (N_24289,N_23839,N_23938);
nor U24290 (N_24290,N_23773,N_23728);
nor U24291 (N_24291,N_23724,N_23832);
and U24292 (N_24292,N_23761,N_23799);
xor U24293 (N_24293,N_23881,N_23824);
nand U24294 (N_24294,N_23719,N_23704);
and U24295 (N_24295,N_23855,N_23823);
or U24296 (N_24296,N_23991,N_23824);
and U24297 (N_24297,N_23866,N_23958);
nand U24298 (N_24298,N_23890,N_23909);
and U24299 (N_24299,N_23829,N_23819);
nand U24300 (N_24300,N_24065,N_24116);
nor U24301 (N_24301,N_24062,N_24269);
nor U24302 (N_24302,N_24255,N_24216);
nand U24303 (N_24303,N_24289,N_24097);
nand U24304 (N_24304,N_24106,N_24279);
xnor U24305 (N_24305,N_24205,N_24090);
xor U24306 (N_24306,N_24144,N_24112);
or U24307 (N_24307,N_24247,N_24037);
or U24308 (N_24308,N_24108,N_24230);
or U24309 (N_24309,N_24231,N_24174);
nor U24310 (N_24310,N_24163,N_24023);
or U24311 (N_24311,N_24058,N_24249);
nor U24312 (N_24312,N_24122,N_24011);
nor U24313 (N_24313,N_24118,N_24137);
or U24314 (N_24314,N_24153,N_24089);
and U24315 (N_24315,N_24151,N_24043);
xor U24316 (N_24316,N_24154,N_24055);
xor U24317 (N_24317,N_24236,N_24213);
or U24318 (N_24318,N_24202,N_24141);
nand U24319 (N_24319,N_24189,N_24028);
and U24320 (N_24320,N_24282,N_24197);
and U24321 (N_24321,N_24050,N_24179);
xnor U24322 (N_24322,N_24059,N_24252);
nor U24323 (N_24323,N_24192,N_24152);
and U24324 (N_24324,N_24207,N_24087);
and U24325 (N_24325,N_24265,N_24000);
xnor U24326 (N_24326,N_24256,N_24027);
and U24327 (N_24327,N_24067,N_24100);
or U24328 (N_24328,N_24226,N_24129);
xor U24329 (N_24329,N_24267,N_24096);
xnor U24330 (N_24330,N_24042,N_24015);
nor U24331 (N_24331,N_24271,N_24009);
or U24332 (N_24332,N_24227,N_24283);
nand U24333 (N_24333,N_24101,N_24168);
and U24334 (N_24334,N_24007,N_24035);
xor U24335 (N_24335,N_24121,N_24166);
xnor U24336 (N_24336,N_24177,N_24054);
nor U24337 (N_24337,N_24159,N_24048);
nand U24338 (N_24338,N_24240,N_24068);
xor U24339 (N_24339,N_24260,N_24248);
xor U24340 (N_24340,N_24261,N_24085);
or U24341 (N_24341,N_24243,N_24204);
and U24342 (N_24342,N_24018,N_24084);
nor U24343 (N_24343,N_24298,N_24071);
nor U24344 (N_24344,N_24195,N_24276);
or U24345 (N_24345,N_24002,N_24194);
or U24346 (N_24346,N_24031,N_24294);
or U24347 (N_24347,N_24024,N_24286);
xor U24348 (N_24348,N_24081,N_24187);
xor U24349 (N_24349,N_24079,N_24008);
nor U24350 (N_24350,N_24056,N_24244);
and U24351 (N_24351,N_24201,N_24171);
and U24352 (N_24352,N_24257,N_24045);
and U24353 (N_24353,N_24099,N_24128);
nand U24354 (N_24354,N_24188,N_24274);
nor U24355 (N_24355,N_24039,N_24021);
and U24356 (N_24356,N_24093,N_24033);
nand U24357 (N_24357,N_24125,N_24262);
nor U24358 (N_24358,N_24281,N_24223);
xnor U24359 (N_24359,N_24047,N_24113);
nand U24360 (N_24360,N_24211,N_24044);
or U24361 (N_24361,N_24228,N_24117);
or U24362 (N_24362,N_24155,N_24135);
xnor U24363 (N_24363,N_24025,N_24127);
xor U24364 (N_24364,N_24217,N_24026);
or U24365 (N_24365,N_24221,N_24190);
nand U24366 (N_24366,N_24268,N_24126);
or U24367 (N_24367,N_24034,N_24086);
or U24368 (N_24368,N_24158,N_24091);
nand U24369 (N_24369,N_24246,N_24291);
xor U24370 (N_24370,N_24242,N_24070);
and U24371 (N_24371,N_24077,N_24133);
nor U24372 (N_24372,N_24280,N_24094);
nand U24373 (N_24373,N_24212,N_24175);
xor U24374 (N_24374,N_24098,N_24156);
xnor U24375 (N_24375,N_24235,N_24075);
xor U24376 (N_24376,N_24073,N_24001);
nor U24377 (N_24377,N_24131,N_24209);
or U24378 (N_24378,N_24191,N_24147);
or U24379 (N_24379,N_24234,N_24016);
or U24380 (N_24380,N_24210,N_24132);
or U24381 (N_24381,N_24064,N_24134);
xnor U24382 (N_24382,N_24287,N_24119);
nor U24383 (N_24383,N_24299,N_24130);
nor U24384 (N_24384,N_24005,N_24264);
nor U24385 (N_24385,N_24104,N_24046);
and U24386 (N_24386,N_24275,N_24105);
nor U24387 (N_24387,N_24273,N_24297);
and U24388 (N_24388,N_24120,N_24167);
xnor U24389 (N_24389,N_24038,N_24136);
nand U24390 (N_24390,N_24111,N_24143);
or U24391 (N_24391,N_24010,N_24115);
nor U24392 (N_24392,N_24258,N_24041);
or U24393 (N_24393,N_24245,N_24170);
nor U24394 (N_24394,N_24040,N_24102);
and U24395 (N_24395,N_24032,N_24150);
xor U24396 (N_24396,N_24083,N_24030);
nor U24397 (N_24397,N_24003,N_24270);
nand U24398 (N_24398,N_24263,N_24004);
nor U24399 (N_24399,N_24251,N_24186);
or U24400 (N_24400,N_24161,N_24165);
xor U24401 (N_24401,N_24013,N_24053);
and U24402 (N_24402,N_24285,N_24239);
or U24403 (N_24403,N_24214,N_24019);
nand U24404 (N_24404,N_24149,N_24061);
xnor U24405 (N_24405,N_24200,N_24220);
nand U24406 (N_24406,N_24254,N_24082);
xor U24407 (N_24407,N_24052,N_24215);
xnor U24408 (N_24408,N_24172,N_24088);
xnor U24409 (N_24409,N_24014,N_24225);
nor U24410 (N_24410,N_24145,N_24057);
nor U24411 (N_24411,N_24066,N_24290);
xor U24412 (N_24412,N_24138,N_24266);
nand U24413 (N_24413,N_24110,N_24160);
and U24414 (N_24414,N_24006,N_24095);
nor U24415 (N_24415,N_24080,N_24241);
nand U24416 (N_24416,N_24278,N_24185);
xor U24417 (N_24417,N_24193,N_24277);
xnor U24418 (N_24418,N_24284,N_24076);
or U24419 (N_24419,N_24253,N_24103);
or U24420 (N_24420,N_24029,N_24199);
xor U24421 (N_24421,N_24222,N_24139);
xnor U24422 (N_24422,N_24022,N_24229);
nor U24423 (N_24423,N_24036,N_24292);
and U24424 (N_24424,N_24178,N_24224);
nor U24425 (N_24425,N_24164,N_24293);
nor U24426 (N_24426,N_24232,N_24107);
and U24427 (N_24427,N_24272,N_24020);
and U24428 (N_24428,N_24233,N_24173);
nor U24429 (N_24429,N_24060,N_24296);
or U24430 (N_24430,N_24051,N_24157);
and U24431 (N_24431,N_24238,N_24295);
or U24432 (N_24432,N_24148,N_24017);
xnor U24433 (N_24433,N_24074,N_24069);
nor U24434 (N_24434,N_24072,N_24012);
xor U24435 (N_24435,N_24218,N_24181);
and U24436 (N_24436,N_24196,N_24049);
or U24437 (N_24437,N_24063,N_24109);
nand U24438 (N_24438,N_24176,N_24124);
nand U24439 (N_24439,N_24114,N_24288);
and U24440 (N_24440,N_24184,N_24169);
or U24441 (N_24441,N_24219,N_24208);
xnor U24442 (N_24442,N_24078,N_24123);
nor U24443 (N_24443,N_24237,N_24146);
nor U24444 (N_24444,N_24142,N_24198);
and U24445 (N_24445,N_24182,N_24250);
or U24446 (N_24446,N_24162,N_24259);
nor U24447 (N_24447,N_24203,N_24183);
nand U24448 (N_24448,N_24140,N_24092);
nor U24449 (N_24449,N_24180,N_24206);
or U24450 (N_24450,N_24283,N_24202);
and U24451 (N_24451,N_24243,N_24130);
nand U24452 (N_24452,N_24157,N_24175);
nor U24453 (N_24453,N_24151,N_24259);
nand U24454 (N_24454,N_24030,N_24050);
nand U24455 (N_24455,N_24077,N_24249);
xnor U24456 (N_24456,N_24200,N_24265);
and U24457 (N_24457,N_24084,N_24035);
or U24458 (N_24458,N_24005,N_24245);
nor U24459 (N_24459,N_24299,N_24150);
nand U24460 (N_24460,N_24256,N_24107);
nand U24461 (N_24461,N_24074,N_24166);
xor U24462 (N_24462,N_24181,N_24071);
nor U24463 (N_24463,N_24167,N_24210);
xnor U24464 (N_24464,N_24267,N_24280);
or U24465 (N_24465,N_24027,N_24074);
nand U24466 (N_24466,N_24282,N_24297);
or U24467 (N_24467,N_24178,N_24072);
nor U24468 (N_24468,N_24078,N_24193);
or U24469 (N_24469,N_24183,N_24065);
nor U24470 (N_24470,N_24047,N_24270);
nand U24471 (N_24471,N_24020,N_24112);
and U24472 (N_24472,N_24245,N_24270);
nor U24473 (N_24473,N_24240,N_24236);
nor U24474 (N_24474,N_24037,N_24226);
and U24475 (N_24475,N_24294,N_24004);
xor U24476 (N_24476,N_24290,N_24294);
and U24477 (N_24477,N_24082,N_24184);
nand U24478 (N_24478,N_24167,N_24048);
nor U24479 (N_24479,N_24090,N_24069);
nand U24480 (N_24480,N_24240,N_24046);
and U24481 (N_24481,N_24116,N_24238);
or U24482 (N_24482,N_24290,N_24266);
nor U24483 (N_24483,N_24004,N_24057);
nand U24484 (N_24484,N_24189,N_24050);
nand U24485 (N_24485,N_24117,N_24077);
or U24486 (N_24486,N_24232,N_24255);
xnor U24487 (N_24487,N_24259,N_24200);
or U24488 (N_24488,N_24001,N_24017);
nor U24489 (N_24489,N_24151,N_24029);
or U24490 (N_24490,N_24091,N_24131);
nand U24491 (N_24491,N_24202,N_24002);
nand U24492 (N_24492,N_24135,N_24186);
or U24493 (N_24493,N_24185,N_24013);
nor U24494 (N_24494,N_24057,N_24021);
nand U24495 (N_24495,N_24130,N_24151);
and U24496 (N_24496,N_24199,N_24259);
nor U24497 (N_24497,N_24127,N_24179);
or U24498 (N_24498,N_24247,N_24021);
nand U24499 (N_24499,N_24087,N_24220);
or U24500 (N_24500,N_24118,N_24291);
xnor U24501 (N_24501,N_24038,N_24278);
nor U24502 (N_24502,N_24177,N_24215);
nor U24503 (N_24503,N_24211,N_24128);
nor U24504 (N_24504,N_24046,N_24015);
xor U24505 (N_24505,N_24013,N_24007);
or U24506 (N_24506,N_24229,N_24269);
and U24507 (N_24507,N_24078,N_24051);
and U24508 (N_24508,N_24053,N_24237);
xnor U24509 (N_24509,N_24272,N_24029);
nor U24510 (N_24510,N_24236,N_24196);
xor U24511 (N_24511,N_24055,N_24011);
nand U24512 (N_24512,N_24234,N_24137);
nor U24513 (N_24513,N_24213,N_24078);
nor U24514 (N_24514,N_24248,N_24056);
or U24515 (N_24515,N_24097,N_24176);
nor U24516 (N_24516,N_24124,N_24040);
or U24517 (N_24517,N_24100,N_24296);
or U24518 (N_24518,N_24069,N_24150);
nand U24519 (N_24519,N_24045,N_24198);
nand U24520 (N_24520,N_24025,N_24141);
nand U24521 (N_24521,N_24215,N_24121);
or U24522 (N_24522,N_24272,N_24175);
and U24523 (N_24523,N_24088,N_24020);
xor U24524 (N_24524,N_24182,N_24049);
nor U24525 (N_24525,N_24260,N_24241);
nand U24526 (N_24526,N_24170,N_24263);
xnor U24527 (N_24527,N_24104,N_24283);
nand U24528 (N_24528,N_24298,N_24203);
nor U24529 (N_24529,N_24236,N_24280);
xnor U24530 (N_24530,N_24068,N_24002);
xnor U24531 (N_24531,N_24281,N_24133);
xor U24532 (N_24532,N_24295,N_24239);
nand U24533 (N_24533,N_24283,N_24076);
nand U24534 (N_24534,N_24248,N_24129);
xnor U24535 (N_24535,N_24164,N_24037);
nor U24536 (N_24536,N_24275,N_24139);
xor U24537 (N_24537,N_24062,N_24019);
xor U24538 (N_24538,N_24126,N_24243);
nor U24539 (N_24539,N_24174,N_24049);
or U24540 (N_24540,N_24204,N_24053);
or U24541 (N_24541,N_24173,N_24024);
nor U24542 (N_24542,N_24291,N_24230);
xor U24543 (N_24543,N_24180,N_24080);
and U24544 (N_24544,N_24208,N_24225);
or U24545 (N_24545,N_24127,N_24122);
nand U24546 (N_24546,N_24050,N_24017);
nor U24547 (N_24547,N_24286,N_24219);
and U24548 (N_24548,N_24047,N_24122);
and U24549 (N_24549,N_24067,N_24011);
nor U24550 (N_24550,N_24104,N_24058);
and U24551 (N_24551,N_24164,N_24031);
nor U24552 (N_24552,N_24239,N_24206);
xnor U24553 (N_24553,N_24216,N_24262);
nand U24554 (N_24554,N_24130,N_24185);
xnor U24555 (N_24555,N_24231,N_24238);
and U24556 (N_24556,N_24206,N_24234);
and U24557 (N_24557,N_24058,N_24196);
xor U24558 (N_24558,N_24283,N_24171);
xnor U24559 (N_24559,N_24150,N_24114);
or U24560 (N_24560,N_24163,N_24052);
nand U24561 (N_24561,N_24261,N_24184);
nor U24562 (N_24562,N_24233,N_24263);
and U24563 (N_24563,N_24051,N_24249);
and U24564 (N_24564,N_24121,N_24081);
nand U24565 (N_24565,N_24181,N_24299);
or U24566 (N_24566,N_24111,N_24271);
and U24567 (N_24567,N_24007,N_24131);
and U24568 (N_24568,N_24264,N_24106);
xnor U24569 (N_24569,N_24228,N_24279);
xor U24570 (N_24570,N_24272,N_24088);
or U24571 (N_24571,N_24011,N_24212);
nor U24572 (N_24572,N_24133,N_24093);
and U24573 (N_24573,N_24233,N_24006);
or U24574 (N_24574,N_24126,N_24178);
and U24575 (N_24575,N_24266,N_24171);
nor U24576 (N_24576,N_24118,N_24010);
nor U24577 (N_24577,N_24201,N_24108);
and U24578 (N_24578,N_24165,N_24033);
xnor U24579 (N_24579,N_24206,N_24062);
nor U24580 (N_24580,N_24056,N_24049);
and U24581 (N_24581,N_24176,N_24090);
nor U24582 (N_24582,N_24003,N_24170);
nor U24583 (N_24583,N_24135,N_24193);
nor U24584 (N_24584,N_24238,N_24249);
or U24585 (N_24585,N_24259,N_24266);
nand U24586 (N_24586,N_24010,N_24178);
nor U24587 (N_24587,N_24036,N_24233);
and U24588 (N_24588,N_24172,N_24061);
or U24589 (N_24589,N_24197,N_24259);
nor U24590 (N_24590,N_24041,N_24234);
nand U24591 (N_24591,N_24196,N_24095);
xnor U24592 (N_24592,N_24160,N_24101);
nand U24593 (N_24593,N_24145,N_24206);
nor U24594 (N_24594,N_24284,N_24100);
or U24595 (N_24595,N_24120,N_24062);
xor U24596 (N_24596,N_24044,N_24189);
and U24597 (N_24597,N_24166,N_24087);
nor U24598 (N_24598,N_24143,N_24126);
nor U24599 (N_24599,N_24140,N_24141);
and U24600 (N_24600,N_24403,N_24356);
nor U24601 (N_24601,N_24332,N_24420);
xor U24602 (N_24602,N_24490,N_24351);
xnor U24603 (N_24603,N_24474,N_24331);
and U24604 (N_24604,N_24410,N_24461);
nor U24605 (N_24605,N_24498,N_24556);
and U24606 (N_24606,N_24486,N_24530);
xor U24607 (N_24607,N_24585,N_24427);
xor U24608 (N_24608,N_24570,N_24496);
nor U24609 (N_24609,N_24590,N_24405);
nand U24610 (N_24610,N_24528,N_24564);
nor U24611 (N_24611,N_24416,N_24449);
or U24612 (N_24612,N_24598,N_24436);
xnor U24613 (N_24613,N_24561,N_24434);
xor U24614 (N_24614,N_24450,N_24360);
xor U24615 (N_24615,N_24300,N_24574);
xor U24616 (N_24616,N_24318,N_24509);
xor U24617 (N_24617,N_24479,N_24518);
and U24618 (N_24618,N_24302,N_24320);
and U24619 (N_24619,N_24525,N_24371);
and U24620 (N_24620,N_24488,N_24435);
and U24621 (N_24621,N_24539,N_24306);
and U24622 (N_24622,N_24563,N_24358);
xor U24623 (N_24623,N_24465,N_24557);
nand U24624 (N_24624,N_24534,N_24549);
or U24625 (N_24625,N_24388,N_24417);
or U24626 (N_24626,N_24505,N_24552);
or U24627 (N_24627,N_24357,N_24473);
nor U24628 (N_24628,N_24596,N_24385);
and U24629 (N_24629,N_24425,N_24307);
and U24630 (N_24630,N_24431,N_24379);
and U24631 (N_24631,N_24487,N_24433);
and U24632 (N_24632,N_24338,N_24316);
and U24633 (N_24633,N_24482,N_24391);
nor U24634 (N_24634,N_24418,N_24346);
or U24635 (N_24635,N_24322,N_24523);
nor U24636 (N_24636,N_24312,N_24430);
xor U24637 (N_24637,N_24339,N_24581);
nor U24638 (N_24638,N_24377,N_24462);
xor U24639 (N_24639,N_24454,N_24582);
nor U24640 (N_24640,N_24413,N_24527);
xor U24641 (N_24641,N_24368,N_24345);
or U24642 (N_24642,N_24389,N_24476);
nand U24643 (N_24643,N_24484,N_24458);
or U24644 (N_24644,N_24562,N_24508);
nor U24645 (N_24645,N_24426,N_24513);
nand U24646 (N_24646,N_24411,N_24392);
nand U24647 (N_24647,N_24369,N_24439);
nand U24648 (N_24648,N_24515,N_24538);
nor U24649 (N_24649,N_24429,N_24399);
nor U24650 (N_24650,N_24492,N_24468);
xor U24651 (N_24651,N_24572,N_24423);
nor U24652 (N_24652,N_24397,N_24576);
nor U24653 (N_24653,N_24412,N_24567);
or U24654 (N_24654,N_24308,N_24344);
nor U24655 (N_24655,N_24526,N_24355);
or U24656 (N_24656,N_24553,N_24428);
or U24657 (N_24657,N_24510,N_24521);
nand U24658 (N_24658,N_24342,N_24364);
or U24659 (N_24659,N_24540,N_24375);
and U24660 (N_24660,N_24363,N_24470);
nor U24661 (N_24661,N_24575,N_24500);
nor U24662 (N_24662,N_24477,N_24578);
nand U24663 (N_24663,N_24489,N_24566);
xor U24664 (N_24664,N_24361,N_24592);
and U24665 (N_24665,N_24336,N_24466);
nand U24666 (N_24666,N_24464,N_24475);
or U24667 (N_24667,N_24373,N_24365);
or U24668 (N_24668,N_24579,N_24343);
nor U24669 (N_24669,N_24536,N_24478);
xnor U24670 (N_24670,N_24506,N_24401);
nor U24671 (N_24671,N_24400,N_24502);
xnor U24672 (N_24672,N_24384,N_24447);
and U24673 (N_24673,N_24547,N_24531);
or U24674 (N_24674,N_24443,N_24376);
nor U24675 (N_24675,N_24512,N_24594);
or U24676 (N_24676,N_24471,N_24324);
and U24677 (N_24677,N_24480,N_24551);
nand U24678 (N_24678,N_24472,N_24370);
nor U24679 (N_24679,N_24352,N_24587);
xor U24680 (N_24680,N_24390,N_24593);
nor U24681 (N_24681,N_24548,N_24366);
nor U24682 (N_24682,N_24440,N_24387);
and U24683 (N_24683,N_24481,N_24541);
nand U24684 (N_24684,N_24348,N_24441);
nand U24685 (N_24685,N_24334,N_24325);
nand U24686 (N_24686,N_24558,N_24337);
nor U24687 (N_24687,N_24532,N_24381);
nor U24688 (N_24688,N_24414,N_24577);
nor U24689 (N_24689,N_24595,N_24326);
nand U24690 (N_24690,N_24341,N_24437);
nand U24691 (N_24691,N_24565,N_24580);
or U24692 (N_24692,N_24304,N_24503);
nand U24693 (N_24693,N_24455,N_24395);
and U24694 (N_24694,N_24559,N_24485);
nor U24695 (N_24695,N_24599,N_24330);
xnor U24696 (N_24696,N_24483,N_24408);
nand U24697 (N_24697,N_24327,N_24317);
xor U24698 (N_24698,N_24347,N_24545);
nor U24699 (N_24699,N_24374,N_24456);
and U24700 (N_24700,N_24448,N_24340);
or U24701 (N_24701,N_24367,N_24444);
and U24702 (N_24702,N_24323,N_24314);
nand U24703 (N_24703,N_24386,N_24380);
nor U24704 (N_24704,N_24402,N_24504);
or U24705 (N_24705,N_24584,N_24573);
or U24706 (N_24706,N_24451,N_24511);
nand U24707 (N_24707,N_24383,N_24514);
nand U24708 (N_24708,N_24544,N_24537);
xor U24709 (N_24709,N_24409,N_24305);
nand U24710 (N_24710,N_24522,N_24493);
xnor U24711 (N_24711,N_24546,N_24315);
nor U24712 (N_24712,N_24394,N_24560);
or U24713 (N_24713,N_24497,N_24469);
xor U24714 (N_24714,N_24350,N_24353);
nor U24715 (N_24715,N_24311,N_24533);
and U24716 (N_24716,N_24393,N_24589);
and U24717 (N_24717,N_24419,N_24378);
and U24718 (N_24718,N_24398,N_24349);
or U24719 (N_24719,N_24586,N_24501);
and U24720 (N_24720,N_24467,N_24591);
xor U24721 (N_24721,N_24568,N_24404);
and U24722 (N_24722,N_24309,N_24588);
nor U24723 (N_24723,N_24571,N_24438);
nand U24724 (N_24724,N_24446,N_24457);
or U24725 (N_24725,N_24445,N_24335);
nand U24726 (N_24726,N_24460,N_24421);
nand U24727 (N_24727,N_24301,N_24303);
or U24728 (N_24728,N_24362,N_24396);
nand U24729 (N_24729,N_24550,N_24569);
and U24730 (N_24730,N_24597,N_24313);
nand U24731 (N_24731,N_24422,N_24310);
or U24732 (N_24732,N_24407,N_24507);
xor U24733 (N_24733,N_24328,N_24453);
or U24734 (N_24734,N_24542,N_24491);
or U24735 (N_24735,N_24406,N_24529);
nand U24736 (N_24736,N_24463,N_24333);
or U24737 (N_24737,N_24354,N_24516);
and U24738 (N_24738,N_24499,N_24554);
xnor U24739 (N_24739,N_24321,N_24535);
nor U24740 (N_24740,N_24424,N_24329);
nand U24741 (N_24741,N_24543,N_24432);
nor U24742 (N_24742,N_24524,N_24494);
nand U24743 (N_24743,N_24415,N_24555);
and U24744 (N_24744,N_24459,N_24517);
and U24745 (N_24745,N_24372,N_24382);
nand U24746 (N_24746,N_24319,N_24442);
or U24747 (N_24747,N_24520,N_24519);
or U24748 (N_24748,N_24495,N_24359);
and U24749 (N_24749,N_24583,N_24452);
nand U24750 (N_24750,N_24542,N_24593);
xor U24751 (N_24751,N_24478,N_24573);
and U24752 (N_24752,N_24305,N_24456);
xnor U24753 (N_24753,N_24349,N_24418);
xor U24754 (N_24754,N_24551,N_24421);
and U24755 (N_24755,N_24483,N_24543);
xnor U24756 (N_24756,N_24367,N_24438);
nor U24757 (N_24757,N_24412,N_24548);
xnor U24758 (N_24758,N_24430,N_24538);
or U24759 (N_24759,N_24354,N_24577);
and U24760 (N_24760,N_24566,N_24585);
xor U24761 (N_24761,N_24473,N_24599);
and U24762 (N_24762,N_24544,N_24402);
nand U24763 (N_24763,N_24458,N_24435);
xor U24764 (N_24764,N_24458,N_24437);
and U24765 (N_24765,N_24551,N_24314);
nand U24766 (N_24766,N_24539,N_24465);
nor U24767 (N_24767,N_24575,N_24493);
or U24768 (N_24768,N_24509,N_24565);
nor U24769 (N_24769,N_24567,N_24337);
nand U24770 (N_24770,N_24325,N_24422);
nor U24771 (N_24771,N_24421,N_24585);
nor U24772 (N_24772,N_24581,N_24485);
xnor U24773 (N_24773,N_24498,N_24518);
nand U24774 (N_24774,N_24403,N_24361);
and U24775 (N_24775,N_24561,N_24533);
nor U24776 (N_24776,N_24358,N_24483);
and U24777 (N_24777,N_24311,N_24549);
xnor U24778 (N_24778,N_24561,N_24473);
xor U24779 (N_24779,N_24489,N_24482);
nor U24780 (N_24780,N_24539,N_24542);
and U24781 (N_24781,N_24403,N_24576);
nand U24782 (N_24782,N_24505,N_24347);
xnor U24783 (N_24783,N_24324,N_24434);
xnor U24784 (N_24784,N_24487,N_24556);
xnor U24785 (N_24785,N_24597,N_24505);
nor U24786 (N_24786,N_24533,N_24356);
and U24787 (N_24787,N_24362,N_24402);
or U24788 (N_24788,N_24488,N_24554);
and U24789 (N_24789,N_24394,N_24365);
and U24790 (N_24790,N_24467,N_24520);
xor U24791 (N_24791,N_24582,N_24435);
and U24792 (N_24792,N_24312,N_24528);
or U24793 (N_24793,N_24525,N_24383);
and U24794 (N_24794,N_24372,N_24424);
nor U24795 (N_24795,N_24304,N_24517);
xnor U24796 (N_24796,N_24473,N_24534);
and U24797 (N_24797,N_24454,N_24353);
and U24798 (N_24798,N_24570,N_24384);
nand U24799 (N_24799,N_24475,N_24461);
nor U24800 (N_24800,N_24433,N_24376);
nor U24801 (N_24801,N_24499,N_24550);
nand U24802 (N_24802,N_24304,N_24451);
or U24803 (N_24803,N_24476,N_24431);
xor U24804 (N_24804,N_24467,N_24327);
and U24805 (N_24805,N_24582,N_24429);
xnor U24806 (N_24806,N_24592,N_24305);
and U24807 (N_24807,N_24322,N_24535);
nor U24808 (N_24808,N_24338,N_24328);
nor U24809 (N_24809,N_24571,N_24325);
nand U24810 (N_24810,N_24549,N_24440);
or U24811 (N_24811,N_24446,N_24330);
nand U24812 (N_24812,N_24579,N_24440);
nand U24813 (N_24813,N_24369,N_24543);
or U24814 (N_24814,N_24444,N_24538);
and U24815 (N_24815,N_24326,N_24410);
or U24816 (N_24816,N_24406,N_24434);
nor U24817 (N_24817,N_24593,N_24421);
nand U24818 (N_24818,N_24392,N_24584);
or U24819 (N_24819,N_24478,N_24408);
nand U24820 (N_24820,N_24594,N_24493);
xnor U24821 (N_24821,N_24472,N_24588);
or U24822 (N_24822,N_24522,N_24354);
xor U24823 (N_24823,N_24591,N_24374);
or U24824 (N_24824,N_24573,N_24339);
nor U24825 (N_24825,N_24501,N_24417);
nor U24826 (N_24826,N_24478,N_24402);
nor U24827 (N_24827,N_24425,N_24555);
or U24828 (N_24828,N_24403,N_24368);
xor U24829 (N_24829,N_24327,N_24590);
xor U24830 (N_24830,N_24550,N_24544);
and U24831 (N_24831,N_24385,N_24548);
nor U24832 (N_24832,N_24454,N_24563);
or U24833 (N_24833,N_24431,N_24316);
nor U24834 (N_24834,N_24596,N_24383);
nand U24835 (N_24835,N_24561,N_24343);
or U24836 (N_24836,N_24317,N_24370);
and U24837 (N_24837,N_24342,N_24546);
nor U24838 (N_24838,N_24592,N_24491);
xnor U24839 (N_24839,N_24356,N_24463);
and U24840 (N_24840,N_24573,N_24574);
or U24841 (N_24841,N_24565,N_24329);
and U24842 (N_24842,N_24433,N_24366);
nor U24843 (N_24843,N_24397,N_24446);
nand U24844 (N_24844,N_24315,N_24471);
nor U24845 (N_24845,N_24410,N_24305);
or U24846 (N_24846,N_24369,N_24413);
and U24847 (N_24847,N_24565,N_24545);
and U24848 (N_24848,N_24596,N_24558);
and U24849 (N_24849,N_24517,N_24434);
xnor U24850 (N_24850,N_24489,N_24461);
and U24851 (N_24851,N_24424,N_24489);
nor U24852 (N_24852,N_24388,N_24475);
or U24853 (N_24853,N_24388,N_24381);
and U24854 (N_24854,N_24376,N_24524);
nor U24855 (N_24855,N_24492,N_24572);
xor U24856 (N_24856,N_24591,N_24565);
and U24857 (N_24857,N_24545,N_24416);
nor U24858 (N_24858,N_24516,N_24495);
xnor U24859 (N_24859,N_24408,N_24514);
nand U24860 (N_24860,N_24535,N_24569);
xnor U24861 (N_24861,N_24372,N_24465);
nor U24862 (N_24862,N_24570,N_24550);
nand U24863 (N_24863,N_24326,N_24574);
xnor U24864 (N_24864,N_24526,N_24579);
xor U24865 (N_24865,N_24465,N_24525);
or U24866 (N_24866,N_24426,N_24347);
xnor U24867 (N_24867,N_24502,N_24459);
nand U24868 (N_24868,N_24366,N_24557);
or U24869 (N_24869,N_24368,N_24432);
and U24870 (N_24870,N_24332,N_24340);
or U24871 (N_24871,N_24309,N_24326);
and U24872 (N_24872,N_24420,N_24438);
or U24873 (N_24873,N_24512,N_24548);
and U24874 (N_24874,N_24315,N_24407);
or U24875 (N_24875,N_24425,N_24466);
and U24876 (N_24876,N_24460,N_24553);
and U24877 (N_24877,N_24337,N_24542);
and U24878 (N_24878,N_24480,N_24396);
nor U24879 (N_24879,N_24461,N_24539);
nand U24880 (N_24880,N_24478,N_24349);
nor U24881 (N_24881,N_24409,N_24362);
xnor U24882 (N_24882,N_24508,N_24585);
xnor U24883 (N_24883,N_24348,N_24485);
and U24884 (N_24884,N_24369,N_24436);
and U24885 (N_24885,N_24372,N_24544);
or U24886 (N_24886,N_24441,N_24304);
or U24887 (N_24887,N_24516,N_24392);
and U24888 (N_24888,N_24548,N_24398);
and U24889 (N_24889,N_24436,N_24463);
xnor U24890 (N_24890,N_24317,N_24435);
nand U24891 (N_24891,N_24597,N_24473);
nor U24892 (N_24892,N_24550,N_24519);
or U24893 (N_24893,N_24399,N_24466);
nand U24894 (N_24894,N_24385,N_24449);
xnor U24895 (N_24895,N_24407,N_24340);
and U24896 (N_24896,N_24538,N_24390);
xnor U24897 (N_24897,N_24569,N_24457);
and U24898 (N_24898,N_24588,N_24580);
nor U24899 (N_24899,N_24380,N_24460);
nand U24900 (N_24900,N_24611,N_24608);
and U24901 (N_24901,N_24613,N_24755);
nand U24902 (N_24902,N_24650,N_24673);
nor U24903 (N_24903,N_24645,N_24668);
or U24904 (N_24904,N_24712,N_24688);
nor U24905 (N_24905,N_24609,N_24617);
nand U24906 (N_24906,N_24797,N_24640);
or U24907 (N_24907,N_24761,N_24666);
or U24908 (N_24908,N_24665,N_24888);
nand U24909 (N_24909,N_24649,N_24777);
xor U24910 (N_24910,N_24618,N_24766);
xor U24911 (N_24911,N_24612,N_24843);
xor U24912 (N_24912,N_24816,N_24678);
xor U24913 (N_24913,N_24760,N_24833);
nand U24914 (N_24914,N_24871,N_24742);
or U24915 (N_24915,N_24628,N_24773);
and U24916 (N_24916,N_24614,N_24890);
nand U24917 (N_24917,N_24895,N_24835);
xor U24918 (N_24918,N_24732,N_24641);
nor U24919 (N_24919,N_24644,N_24824);
and U24920 (N_24920,N_24606,N_24826);
or U24921 (N_24921,N_24892,N_24779);
xnor U24922 (N_24922,N_24686,N_24707);
nand U24923 (N_24923,N_24889,N_24702);
nand U24924 (N_24924,N_24625,N_24872);
or U24925 (N_24925,N_24726,N_24756);
nand U24926 (N_24926,N_24727,N_24848);
or U24927 (N_24927,N_24801,N_24704);
nor U24928 (N_24928,N_24845,N_24720);
xnor U24929 (N_24929,N_24868,N_24854);
nor U24930 (N_24930,N_24894,N_24663);
or U24931 (N_24931,N_24786,N_24714);
xnor U24932 (N_24932,N_24604,N_24775);
xnor U24933 (N_24933,N_24810,N_24631);
or U24934 (N_24934,N_24697,N_24667);
nor U24935 (N_24935,N_24737,N_24881);
and U24936 (N_24936,N_24780,N_24870);
nand U24937 (N_24937,N_24654,N_24770);
or U24938 (N_24938,N_24887,N_24701);
xnor U24939 (N_24939,N_24836,N_24602);
or U24940 (N_24940,N_24800,N_24837);
xnor U24941 (N_24941,N_24627,N_24776);
and U24942 (N_24942,N_24818,N_24684);
nor U24943 (N_24943,N_24869,N_24823);
nand U24944 (N_24944,N_24815,N_24794);
and U24945 (N_24945,N_24600,N_24687);
and U24946 (N_24946,N_24691,N_24656);
nor U24947 (N_24947,N_24693,N_24821);
or U24948 (N_24948,N_24638,N_24763);
or U24949 (N_24949,N_24758,N_24875);
nand U24950 (N_24950,N_24859,N_24730);
and U24951 (N_24951,N_24739,N_24849);
and U24952 (N_24952,N_24879,N_24711);
nand U24953 (N_24953,N_24782,N_24839);
and U24954 (N_24954,N_24657,N_24689);
or U24955 (N_24955,N_24799,N_24675);
or U24956 (N_24956,N_24876,N_24655);
or U24957 (N_24957,N_24743,N_24831);
xor U24958 (N_24958,N_24793,N_24813);
xor U24959 (N_24959,N_24722,N_24741);
or U24960 (N_24960,N_24671,N_24685);
nor U24961 (N_24961,N_24718,N_24851);
and U24962 (N_24962,N_24768,N_24746);
or U24963 (N_24963,N_24808,N_24731);
and U24964 (N_24964,N_24642,N_24857);
nand U24965 (N_24965,N_24661,N_24728);
and U24966 (N_24966,N_24844,N_24652);
and U24967 (N_24967,N_24771,N_24812);
nor U24968 (N_24968,N_24636,N_24862);
nand U24969 (N_24969,N_24736,N_24715);
xor U24970 (N_24970,N_24695,N_24878);
xnor U24971 (N_24971,N_24795,N_24725);
nand U24972 (N_24972,N_24791,N_24694);
nor U24973 (N_24973,N_24807,N_24825);
nor U24974 (N_24974,N_24623,N_24616);
and U24975 (N_24975,N_24789,N_24819);
and U24976 (N_24976,N_24802,N_24670);
or U24977 (N_24977,N_24774,N_24706);
or U24978 (N_24978,N_24863,N_24750);
nor U24979 (N_24979,N_24834,N_24785);
nand U24980 (N_24980,N_24769,N_24877);
nand U24981 (N_24981,N_24767,N_24735);
and U24982 (N_24982,N_24784,N_24709);
xnor U24983 (N_24983,N_24882,N_24713);
and U24984 (N_24984,N_24647,N_24864);
nor U24985 (N_24985,N_24717,N_24703);
and U24986 (N_24986,N_24733,N_24749);
or U24987 (N_24987,N_24753,N_24705);
xnor U24988 (N_24988,N_24886,N_24729);
and U24989 (N_24989,N_24619,N_24865);
and U24990 (N_24990,N_24814,N_24829);
and U24991 (N_24991,N_24610,N_24669);
nor U24992 (N_24992,N_24867,N_24885);
nor U24993 (N_24993,N_24873,N_24621);
or U24994 (N_24994,N_24788,N_24804);
nor U24995 (N_24995,N_24790,N_24620);
nand U24996 (N_24996,N_24603,N_24752);
nor U24997 (N_24997,N_24632,N_24883);
and U24998 (N_24998,N_24806,N_24861);
nand U24999 (N_24999,N_24855,N_24852);
nand U25000 (N_25000,N_24783,N_24624);
and U25001 (N_25001,N_24662,N_24757);
nand U25002 (N_25002,N_24893,N_24842);
xor U25003 (N_25003,N_24762,N_24648);
xnor U25004 (N_25004,N_24630,N_24853);
nor U25005 (N_25005,N_24811,N_24747);
or U25006 (N_25006,N_24723,N_24798);
xnor U25007 (N_25007,N_24751,N_24787);
and U25008 (N_25008,N_24699,N_24828);
xnor U25009 (N_25009,N_24690,N_24692);
nand U25010 (N_25010,N_24772,N_24708);
or U25011 (N_25011,N_24898,N_24734);
nand U25012 (N_25012,N_24817,N_24622);
or U25013 (N_25013,N_24846,N_24827);
xnor U25014 (N_25014,N_24635,N_24880);
and U25015 (N_25015,N_24778,N_24637);
or U25016 (N_25016,N_24601,N_24674);
or U25017 (N_25017,N_24738,N_24803);
nor U25018 (N_25018,N_24626,N_24809);
xor U25019 (N_25019,N_24651,N_24860);
or U25020 (N_25020,N_24719,N_24633);
nor U25021 (N_25021,N_24897,N_24792);
and U25022 (N_25022,N_24639,N_24805);
xnor U25023 (N_25023,N_24677,N_24850);
nor U25024 (N_25024,N_24754,N_24745);
or U25025 (N_25025,N_24679,N_24765);
xor U25026 (N_25026,N_24840,N_24646);
nor U25027 (N_25027,N_24744,N_24820);
nor U25028 (N_25028,N_24615,N_24653);
nor U25029 (N_25029,N_24899,N_24724);
xor U25030 (N_25030,N_24847,N_24607);
or U25031 (N_25031,N_24716,N_24781);
or U25032 (N_25032,N_24710,N_24858);
nor U25033 (N_25033,N_24896,N_24891);
nor U25034 (N_25034,N_24838,N_24796);
nand U25035 (N_25035,N_24721,N_24841);
and U25036 (N_25036,N_24629,N_24698);
and U25037 (N_25037,N_24700,N_24696);
nor U25038 (N_25038,N_24672,N_24856);
or U25039 (N_25039,N_24680,N_24866);
nand U25040 (N_25040,N_24764,N_24643);
nand U25041 (N_25041,N_24676,N_24664);
xnor U25042 (N_25042,N_24681,N_24605);
nor U25043 (N_25043,N_24682,N_24683);
xor U25044 (N_25044,N_24634,N_24740);
nor U25045 (N_25045,N_24748,N_24874);
nor U25046 (N_25046,N_24658,N_24830);
or U25047 (N_25047,N_24759,N_24822);
xor U25048 (N_25048,N_24660,N_24659);
xnor U25049 (N_25049,N_24832,N_24884);
and U25050 (N_25050,N_24735,N_24697);
nand U25051 (N_25051,N_24602,N_24801);
or U25052 (N_25052,N_24643,N_24898);
or U25053 (N_25053,N_24637,N_24638);
or U25054 (N_25054,N_24614,N_24805);
or U25055 (N_25055,N_24890,N_24678);
nor U25056 (N_25056,N_24633,N_24735);
or U25057 (N_25057,N_24755,N_24879);
xor U25058 (N_25058,N_24671,N_24812);
or U25059 (N_25059,N_24697,N_24812);
nand U25060 (N_25060,N_24896,N_24757);
nor U25061 (N_25061,N_24869,N_24604);
and U25062 (N_25062,N_24624,N_24806);
nand U25063 (N_25063,N_24832,N_24690);
nor U25064 (N_25064,N_24687,N_24886);
xor U25065 (N_25065,N_24735,N_24703);
xnor U25066 (N_25066,N_24743,N_24650);
and U25067 (N_25067,N_24671,N_24828);
xnor U25068 (N_25068,N_24691,N_24620);
nor U25069 (N_25069,N_24842,N_24624);
or U25070 (N_25070,N_24861,N_24840);
nand U25071 (N_25071,N_24632,N_24675);
or U25072 (N_25072,N_24826,N_24757);
nand U25073 (N_25073,N_24679,N_24747);
xnor U25074 (N_25074,N_24851,N_24754);
xnor U25075 (N_25075,N_24717,N_24700);
xor U25076 (N_25076,N_24810,N_24720);
and U25077 (N_25077,N_24685,N_24703);
xnor U25078 (N_25078,N_24896,N_24729);
nor U25079 (N_25079,N_24817,N_24838);
xor U25080 (N_25080,N_24699,N_24640);
xor U25081 (N_25081,N_24753,N_24875);
or U25082 (N_25082,N_24660,N_24720);
nand U25083 (N_25083,N_24873,N_24806);
or U25084 (N_25084,N_24756,N_24897);
nand U25085 (N_25085,N_24825,N_24885);
xnor U25086 (N_25086,N_24689,N_24895);
and U25087 (N_25087,N_24707,N_24683);
nor U25088 (N_25088,N_24808,N_24602);
xor U25089 (N_25089,N_24693,N_24791);
or U25090 (N_25090,N_24816,N_24747);
or U25091 (N_25091,N_24817,N_24758);
nor U25092 (N_25092,N_24764,N_24715);
xor U25093 (N_25093,N_24638,N_24694);
nand U25094 (N_25094,N_24609,N_24781);
or U25095 (N_25095,N_24679,N_24754);
xnor U25096 (N_25096,N_24772,N_24705);
nor U25097 (N_25097,N_24623,N_24700);
or U25098 (N_25098,N_24763,N_24841);
nor U25099 (N_25099,N_24604,N_24819);
xnor U25100 (N_25100,N_24723,N_24713);
nor U25101 (N_25101,N_24640,N_24888);
nor U25102 (N_25102,N_24818,N_24638);
and U25103 (N_25103,N_24879,N_24708);
xnor U25104 (N_25104,N_24869,N_24855);
or U25105 (N_25105,N_24687,N_24850);
xor U25106 (N_25106,N_24804,N_24810);
or U25107 (N_25107,N_24837,N_24881);
nor U25108 (N_25108,N_24714,N_24686);
xor U25109 (N_25109,N_24807,N_24746);
nand U25110 (N_25110,N_24856,N_24773);
nand U25111 (N_25111,N_24818,N_24656);
nand U25112 (N_25112,N_24817,N_24803);
or U25113 (N_25113,N_24604,N_24878);
or U25114 (N_25114,N_24866,N_24617);
or U25115 (N_25115,N_24692,N_24831);
nor U25116 (N_25116,N_24732,N_24743);
and U25117 (N_25117,N_24830,N_24612);
xor U25118 (N_25118,N_24631,N_24790);
xor U25119 (N_25119,N_24664,N_24772);
and U25120 (N_25120,N_24674,N_24698);
and U25121 (N_25121,N_24871,N_24686);
and U25122 (N_25122,N_24864,N_24730);
nand U25123 (N_25123,N_24837,N_24742);
xor U25124 (N_25124,N_24856,N_24766);
and U25125 (N_25125,N_24766,N_24657);
nand U25126 (N_25126,N_24685,N_24797);
or U25127 (N_25127,N_24648,N_24647);
or U25128 (N_25128,N_24612,N_24783);
nand U25129 (N_25129,N_24639,N_24738);
or U25130 (N_25130,N_24813,N_24870);
xor U25131 (N_25131,N_24819,N_24834);
nand U25132 (N_25132,N_24674,N_24784);
nand U25133 (N_25133,N_24612,N_24631);
nand U25134 (N_25134,N_24847,N_24616);
or U25135 (N_25135,N_24825,N_24721);
xnor U25136 (N_25136,N_24635,N_24631);
xnor U25137 (N_25137,N_24809,N_24714);
and U25138 (N_25138,N_24611,N_24709);
nor U25139 (N_25139,N_24633,N_24602);
or U25140 (N_25140,N_24747,N_24859);
and U25141 (N_25141,N_24862,N_24638);
nand U25142 (N_25142,N_24892,N_24620);
nor U25143 (N_25143,N_24641,N_24727);
nand U25144 (N_25144,N_24786,N_24875);
and U25145 (N_25145,N_24622,N_24692);
and U25146 (N_25146,N_24809,N_24838);
nand U25147 (N_25147,N_24654,N_24676);
nand U25148 (N_25148,N_24617,N_24786);
nor U25149 (N_25149,N_24866,N_24832);
nand U25150 (N_25150,N_24859,N_24830);
xor U25151 (N_25151,N_24683,N_24781);
xnor U25152 (N_25152,N_24731,N_24670);
nand U25153 (N_25153,N_24873,N_24755);
nor U25154 (N_25154,N_24735,N_24870);
or U25155 (N_25155,N_24654,N_24652);
nand U25156 (N_25156,N_24801,N_24869);
nor U25157 (N_25157,N_24648,N_24712);
xor U25158 (N_25158,N_24887,N_24685);
nor U25159 (N_25159,N_24797,N_24687);
nor U25160 (N_25160,N_24604,N_24694);
nand U25161 (N_25161,N_24768,N_24818);
nor U25162 (N_25162,N_24841,N_24878);
and U25163 (N_25163,N_24665,N_24825);
and U25164 (N_25164,N_24858,N_24867);
and U25165 (N_25165,N_24817,N_24845);
nor U25166 (N_25166,N_24730,N_24734);
xnor U25167 (N_25167,N_24629,N_24838);
or U25168 (N_25168,N_24631,N_24834);
nand U25169 (N_25169,N_24851,N_24600);
or U25170 (N_25170,N_24770,N_24687);
xor U25171 (N_25171,N_24742,N_24763);
nor U25172 (N_25172,N_24755,N_24807);
xor U25173 (N_25173,N_24749,N_24622);
and U25174 (N_25174,N_24688,N_24610);
nand U25175 (N_25175,N_24720,N_24670);
and U25176 (N_25176,N_24873,N_24692);
or U25177 (N_25177,N_24644,N_24630);
nand U25178 (N_25178,N_24808,N_24612);
nor U25179 (N_25179,N_24832,N_24726);
and U25180 (N_25180,N_24753,N_24663);
and U25181 (N_25181,N_24756,N_24777);
and U25182 (N_25182,N_24739,N_24722);
nor U25183 (N_25183,N_24830,N_24812);
and U25184 (N_25184,N_24745,N_24681);
or U25185 (N_25185,N_24793,N_24611);
nor U25186 (N_25186,N_24721,N_24732);
xor U25187 (N_25187,N_24640,N_24610);
and U25188 (N_25188,N_24627,N_24693);
nor U25189 (N_25189,N_24632,N_24829);
or U25190 (N_25190,N_24726,N_24747);
nor U25191 (N_25191,N_24839,N_24811);
nand U25192 (N_25192,N_24816,N_24718);
nand U25193 (N_25193,N_24617,N_24895);
and U25194 (N_25194,N_24624,N_24851);
and U25195 (N_25195,N_24603,N_24775);
or U25196 (N_25196,N_24727,N_24606);
xor U25197 (N_25197,N_24606,N_24781);
or U25198 (N_25198,N_24879,N_24688);
and U25199 (N_25199,N_24766,N_24649);
nand U25200 (N_25200,N_25181,N_24965);
xor U25201 (N_25201,N_25053,N_25014);
and U25202 (N_25202,N_25160,N_25108);
nor U25203 (N_25203,N_24960,N_25119);
or U25204 (N_25204,N_24935,N_25115);
xnor U25205 (N_25205,N_25177,N_24921);
or U25206 (N_25206,N_25086,N_24946);
xor U25207 (N_25207,N_24913,N_24942);
nor U25208 (N_25208,N_24986,N_25010);
and U25209 (N_25209,N_25156,N_25133);
or U25210 (N_25210,N_25045,N_25071);
xnor U25211 (N_25211,N_25138,N_25185);
or U25212 (N_25212,N_25087,N_24971);
or U25213 (N_25213,N_24991,N_25093);
nand U25214 (N_25214,N_25130,N_25064);
nor U25215 (N_25215,N_25150,N_25186);
and U25216 (N_25216,N_25082,N_25025);
xnor U25217 (N_25217,N_25123,N_25166);
and U25218 (N_25218,N_25011,N_25131);
nand U25219 (N_25219,N_24985,N_24927);
nor U25220 (N_25220,N_25190,N_24918);
nor U25221 (N_25221,N_25132,N_24984);
xor U25222 (N_25222,N_24947,N_24926);
xnor U25223 (N_25223,N_25152,N_24988);
nor U25224 (N_25224,N_25089,N_25050);
xor U25225 (N_25225,N_25081,N_24998);
nor U25226 (N_25226,N_25069,N_25032);
or U25227 (N_25227,N_24901,N_24944);
nor U25228 (N_25228,N_24904,N_25111);
and U25229 (N_25229,N_25194,N_25099);
nand U25230 (N_25230,N_24967,N_24900);
nand U25231 (N_25231,N_25068,N_24990);
nand U25232 (N_25232,N_25136,N_25174);
xor U25233 (N_25233,N_25044,N_25148);
nor U25234 (N_25234,N_24914,N_25055);
xnor U25235 (N_25235,N_25172,N_25070);
nor U25236 (N_25236,N_25007,N_25128);
nand U25237 (N_25237,N_25173,N_25134);
and U25238 (N_25238,N_25066,N_25004);
xor U25239 (N_25239,N_24906,N_25059);
nor U25240 (N_25240,N_25153,N_25037);
nor U25241 (N_25241,N_24954,N_25121);
nor U25242 (N_25242,N_25051,N_24994);
nand U25243 (N_25243,N_25000,N_25022);
nand U25244 (N_25244,N_24919,N_25159);
nand U25245 (N_25245,N_25016,N_25164);
nand U25246 (N_25246,N_24977,N_24905);
xor U25247 (N_25247,N_25057,N_25098);
or U25248 (N_25248,N_24989,N_25100);
nor U25249 (N_25249,N_24902,N_24922);
or U25250 (N_25250,N_24973,N_25056);
nor U25251 (N_25251,N_25195,N_25106);
or U25252 (N_25252,N_24974,N_25104);
xor U25253 (N_25253,N_25002,N_24958);
and U25254 (N_25254,N_25033,N_25184);
nor U25255 (N_25255,N_25084,N_25122);
xnor U25256 (N_25256,N_25120,N_24925);
xnor U25257 (N_25257,N_25080,N_24975);
xnor U25258 (N_25258,N_25075,N_25112);
xor U25259 (N_25259,N_24950,N_25171);
or U25260 (N_25260,N_25178,N_25142);
or U25261 (N_25261,N_25030,N_25013);
and U25262 (N_25262,N_25113,N_24936);
nor U25263 (N_25263,N_24980,N_24963);
or U25264 (N_25264,N_24920,N_24964);
nand U25265 (N_25265,N_24953,N_25073);
xor U25266 (N_25266,N_25039,N_24966);
or U25267 (N_25267,N_25143,N_25008);
and U25268 (N_25268,N_25145,N_25180);
nand U25269 (N_25269,N_25097,N_24931);
nor U25270 (N_25270,N_25062,N_25135);
or U25271 (N_25271,N_24907,N_25001);
xor U25272 (N_25272,N_25198,N_25137);
nor U25273 (N_25273,N_24948,N_25091);
xor U25274 (N_25274,N_25157,N_25058);
nor U25275 (N_25275,N_24987,N_25065);
and U25276 (N_25276,N_24959,N_25079);
and U25277 (N_25277,N_25147,N_24915);
nor U25278 (N_25278,N_24909,N_24910);
nand U25279 (N_25279,N_24941,N_25024);
nand U25280 (N_25280,N_24933,N_25012);
xor U25281 (N_25281,N_25036,N_24940);
nand U25282 (N_25282,N_25199,N_25094);
xor U25283 (N_25283,N_25003,N_24916);
nand U25284 (N_25284,N_24912,N_24978);
nand U25285 (N_25285,N_25175,N_24976);
xor U25286 (N_25286,N_25067,N_25102);
or U25287 (N_25287,N_24945,N_24983);
nand U25288 (N_25288,N_24962,N_25074);
or U25289 (N_25289,N_25061,N_24997);
and U25290 (N_25290,N_25126,N_24939);
or U25291 (N_25291,N_25124,N_25018);
and U25292 (N_25292,N_25072,N_25041);
nor U25293 (N_25293,N_25192,N_25103);
or U25294 (N_25294,N_24949,N_25114);
and U25295 (N_25295,N_24917,N_24996);
or U25296 (N_25296,N_25189,N_25034);
or U25297 (N_25297,N_25006,N_25116);
nand U25298 (N_25298,N_25026,N_25049);
nand U25299 (N_25299,N_24928,N_25170);
or U25300 (N_25300,N_24999,N_25188);
xnor U25301 (N_25301,N_25107,N_25060);
xnor U25302 (N_25302,N_25125,N_25168);
or U25303 (N_25303,N_25127,N_25176);
xnor U25304 (N_25304,N_25110,N_24995);
nor U25305 (N_25305,N_24961,N_25031);
or U25306 (N_25306,N_24992,N_25193);
nand U25307 (N_25307,N_25038,N_25179);
xor U25308 (N_25308,N_25191,N_25047);
nand U25309 (N_25309,N_25076,N_25085);
nand U25310 (N_25310,N_25129,N_24923);
nand U25311 (N_25311,N_25139,N_25077);
nand U25312 (N_25312,N_25141,N_24981);
or U25313 (N_25313,N_25144,N_24982);
and U25314 (N_25314,N_25149,N_25109);
nor U25315 (N_25315,N_25187,N_24993);
nand U25316 (N_25316,N_25015,N_25028);
nor U25317 (N_25317,N_24969,N_25161);
and U25318 (N_25318,N_24937,N_24957);
xnor U25319 (N_25319,N_25162,N_25155);
nor U25320 (N_25320,N_25154,N_24908);
and U25321 (N_25321,N_25048,N_25196);
and U25322 (N_25322,N_25083,N_24979);
and U25323 (N_25323,N_25052,N_25197);
and U25324 (N_25324,N_25090,N_25095);
nand U25325 (N_25325,N_25151,N_25035);
nor U25326 (N_25326,N_25078,N_24968);
xor U25327 (N_25327,N_25118,N_25029);
or U25328 (N_25328,N_24955,N_25054);
or U25329 (N_25329,N_25158,N_24924);
or U25330 (N_25330,N_24943,N_25088);
or U25331 (N_25331,N_25046,N_25140);
nor U25332 (N_25332,N_24970,N_25063);
nand U25333 (N_25333,N_24952,N_25101);
and U25334 (N_25334,N_24932,N_25165);
nor U25335 (N_25335,N_25042,N_25009);
or U25336 (N_25336,N_25005,N_25105);
or U25337 (N_25337,N_25092,N_24930);
nor U25338 (N_25338,N_24972,N_25019);
or U25339 (N_25339,N_25182,N_24934);
or U25340 (N_25340,N_25163,N_24938);
xnor U25341 (N_25341,N_25040,N_25023);
nor U25342 (N_25342,N_25146,N_25017);
or U25343 (N_25343,N_25117,N_24903);
or U25344 (N_25344,N_24951,N_24956);
or U25345 (N_25345,N_25169,N_25183);
nor U25346 (N_25346,N_25096,N_24911);
nor U25347 (N_25347,N_25043,N_24929);
nor U25348 (N_25348,N_25021,N_25167);
nor U25349 (N_25349,N_25027,N_25020);
and U25350 (N_25350,N_24974,N_25136);
and U25351 (N_25351,N_24933,N_25118);
nand U25352 (N_25352,N_25069,N_24912);
nand U25353 (N_25353,N_25137,N_25087);
and U25354 (N_25354,N_24974,N_25160);
nor U25355 (N_25355,N_24955,N_25165);
and U25356 (N_25356,N_25131,N_24976);
nor U25357 (N_25357,N_25044,N_25074);
or U25358 (N_25358,N_24954,N_25083);
xor U25359 (N_25359,N_24961,N_25052);
nand U25360 (N_25360,N_25101,N_25094);
nand U25361 (N_25361,N_25141,N_25092);
nand U25362 (N_25362,N_25152,N_25147);
or U25363 (N_25363,N_25139,N_25162);
and U25364 (N_25364,N_25131,N_25184);
or U25365 (N_25365,N_25049,N_24955);
nand U25366 (N_25366,N_25068,N_25139);
xor U25367 (N_25367,N_25066,N_24998);
nor U25368 (N_25368,N_24983,N_25110);
or U25369 (N_25369,N_24991,N_25082);
nor U25370 (N_25370,N_25171,N_24925);
xnor U25371 (N_25371,N_25136,N_25030);
or U25372 (N_25372,N_25047,N_25088);
nand U25373 (N_25373,N_25079,N_25134);
xor U25374 (N_25374,N_25199,N_24929);
and U25375 (N_25375,N_25096,N_24962);
or U25376 (N_25376,N_24925,N_25049);
nor U25377 (N_25377,N_25063,N_24927);
and U25378 (N_25378,N_25178,N_25196);
and U25379 (N_25379,N_24968,N_25012);
nand U25380 (N_25380,N_25047,N_25028);
xor U25381 (N_25381,N_25124,N_25052);
and U25382 (N_25382,N_24952,N_25153);
nand U25383 (N_25383,N_25136,N_25042);
or U25384 (N_25384,N_24943,N_25116);
nor U25385 (N_25385,N_25013,N_25124);
nand U25386 (N_25386,N_25123,N_25165);
or U25387 (N_25387,N_24918,N_24903);
xnor U25388 (N_25388,N_25099,N_25144);
nand U25389 (N_25389,N_24939,N_25015);
or U25390 (N_25390,N_25028,N_25188);
nor U25391 (N_25391,N_25079,N_25031);
nand U25392 (N_25392,N_24942,N_24998);
and U25393 (N_25393,N_24973,N_25064);
nor U25394 (N_25394,N_25103,N_25116);
xnor U25395 (N_25395,N_25121,N_25009);
and U25396 (N_25396,N_25138,N_25088);
and U25397 (N_25397,N_25114,N_24933);
nor U25398 (N_25398,N_25040,N_25086);
nand U25399 (N_25399,N_25082,N_25196);
nor U25400 (N_25400,N_24960,N_24968);
nand U25401 (N_25401,N_25155,N_25164);
and U25402 (N_25402,N_25176,N_24977);
and U25403 (N_25403,N_25073,N_24951);
or U25404 (N_25404,N_25121,N_25150);
nor U25405 (N_25405,N_25162,N_25122);
nand U25406 (N_25406,N_25034,N_24969);
xnor U25407 (N_25407,N_25049,N_24906);
or U25408 (N_25408,N_25102,N_25021);
nand U25409 (N_25409,N_25080,N_25054);
and U25410 (N_25410,N_24995,N_25011);
nor U25411 (N_25411,N_24911,N_24943);
nor U25412 (N_25412,N_25132,N_25107);
nor U25413 (N_25413,N_25105,N_25110);
nor U25414 (N_25414,N_24918,N_25069);
and U25415 (N_25415,N_25105,N_25037);
xnor U25416 (N_25416,N_25002,N_24908);
nor U25417 (N_25417,N_24916,N_25180);
or U25418 (N_25418,N_25048,N_25087);
xnor U25419 (N_25419,N_25044,N_25176);
or U25420 (N_25420,N_24965,N_25189);
and U25421 (N_25421,N_24961,N_25055);
or U25422 (N_25422,N_25103,N_25124);
xor U25423 (N_25423,N_24953,N_25013);
or U25424 (N_25424,N_25105,N_25138);
and U25425 (N_25425,N_25159,N_25058);
and U25426 (N_25426,N_24990,N_24962);
and U25427 (N_25427,N_24978,N_25180);
nor U25428 (N_25428,N_25031,N_25174);
and U25429 (N_25429,N_25107,N_25051);
and U25430 (N_25430,N_25070,N_25170);
nor U25431 (N_25431,N_25080,N_25152);
and U25432 (N_25432,N_24937,N_25032);
xnor U25433 (N_25433,N_25038,N_25108);
xor U25434 (N_25434,N_25076,N_25122);
xnor U25435 (N_25435,N_25162,N_24916);
nor U25436 (N_25436,N_24964,N_25051);
and U25437 (N_25437,N_25025,N_24969);
and U25438 (N_25438,N_25099,N_25058);
or U25439 (N_25439,N_25068,N_24968);
nand U25440 (N_25440,N_24991,N_25068);
nor U25441 (N_25441,N_25019,N_25140);
and U25442 (N_25442,N_25009,N_25075);
and U25443 (N_25443,N_25150,N_25195);
and U25444 (N_25444,N_25162,N_24906);
and U25445 (N_25445,N_24920,N_25156);
xnor U25446 (N_25446,N_25052,N_25068);
nor U25447 (N_25447,N_24957,N_25156);
nand U25448 (N_25448,N_25103,N_25040);
xor U25449 (N_25449,N_25009,N_25104);
or U25450 (N_25450,N_24902,N_25076);
xnor U25451 (N_25451,N_24989,N_25116);
and U25452 (N_25452,N_25004,N_25185);
nand U25453 (N_25453,N_25042,N_25093);
xnor U25454 (N_25454,N_24910,N_25123);
xor U25455 (N_25455,N_25079,N_25032);
or U25456 (N_25456,N_25131,N_25050);
nand U25457 (N_25457,N_25135,N_24939);
nand U25458 (N_25458,N_24947,N_24904);
or U25459 (N_25459,N_25076,N_25091);
or U25460 (N_25460,N_25180,N_25051);
nand U25461 (N_25461,N_25039,N_25000);
xnor U25462 (N_25462,N_25004,N_25138);
or U25463 (N_25463,N_25183,N_25036);
xnor U25464 (N_25464,N_25141,N_25041);
and U25465 (N_25465,N_24903,N_25016);
nand U25466 (N_25466,N_25194,N_25197);
and U25467 (N_25467,N_24905,N_24981);
nand U25468 (N_25468,N_24904,N_25141);
and U25469 (N_25469,N_24921,N_24925);
nand U25470 (N_25470,N_24980,N_25004);
nand U25471 (N_25471,N_24907,N_24948);
or U25472 (N_25472,N_25018,N_24904);
and U25473 (N_25473,N_24966,N_25004);
nor U25474 (N_25474,N_25134,N_25014);
nor U25475 (N_25475,N_24911,N_25006);
nor U25476 (N_25476,N_24985,N_25171);
xnor U25477 (N_25477,N_24977,N_24957);
or U25478 (N_25478,N_25152,N_25063);
and U25479 (N_25479,N_25142,N_25008);
and U25480 (N_25480,N_25158,N_24917);
and U25481 (N_25481,N_25099,N_25039);
xnor U25482 (N_25482,N_25190,N_25176);
nand U25483 (N_25483,N_24927,N_25185);
or U25484 (N_25484,N_25094,N_24981);
nand U25485 (N_25485,N_24974,N_24922);
or U25486 (N_25486,N_25134,N_24962);
or U25487 (N_25487,N_24990,N_24997);
nor U25488 (N_25488,N_25081,N_25003);
nand U25489 (N_25489,N_25098,N_24917);
xor U25490 (N_25490,N_25093,N_24930);
nor U25491 (N_25491,N_25163,N_25183);
nor U25492 (N_25492,N_24963,N_24967);
nand U25493 (N_25493,N_24933,N_25083);
and U25494 (N_25494,N_24974,N_24948);
nand U25495 (N_25495,N_25181,N_24935);
xor U25496 (N_25496,N_25154,N_25143);
nor U25497 (N_25497,N_25024,N_24974);
and U25498 (N_25498,N_24939,N_25003);
or U25499 (N_25499,N_24913,N_25065);
xnor U25500 (N_25500,N_25389,N_25229);
or U25501 (N_25501,N_25412,N_25421);
xor U25502 (N_25502,N_25479,N_25277);
and U25503 (N_25503,N_25330,N_25336);
and U25504 (N_25504,N_25374,N_25423);
and U25505 (N_25505,N_25284,N_25395);
xnor U25506 (N_25506,N_25472,N_25443);
or U25507 (N_25507,N_25205,N_25486);
nor U25508 (N_25508,N_25359,N_25224);
nor U25509 (N_25509,N_25222,N_25351);
and U25510 (N_25510,N_25429,N_25332);
nor U25511 (N_25511,N_25397,N_25470);
nand U25512 (N_25512,N_25202,N_25311);
nor U25513 (N_25513,N_25393,N_25238);
xor U25514 (N_25514,N_25390,N_25244);
and U25515 (N_25515,N_25498,N_25484);
and U25516 (N_25516,N_25442,N_25258);
xnor U25517 (N_25517,N_25362,N_25207);
or U25518 (N_25518,N_25411,N_25296);
nor U25519 (N_25519,N_25360,N_25223);
nor U25520 (N_25520,N_25241,N_25368);
nand U25521 (N_25521,N_25304,N_25408);
xnor U25522 (N_25522,N_25346,N_25438);
and U25523 (N_25523,N_25451,N_25416);
nor U25524 (N_25524,N_25220,N_25444);
xor U25525 (N_25525,N_25335,N_25372);
and U25526 (N_25526,N_25490,N_25385);
or U25527 (N_25527,N_25289,N_25237);
or U25528 (N_25528,N_25495,N_25320);
nor U25529 (N_25529,N_25278,N_25405);
nor U25530 (N_25530,N_25328,N_25268);
and U25531 (N_25531,N_25434,N_25459);
nor U25532 (N_25532,N_25256,N_25483);
xnor U25533 (N_25533,N_25274,N_25373);
and U25534 (N_25534,N_25380,N_25454);
or U25535 (N_25535,N_25428,N_25325);
or U25536 (N_25536,N_25246,N_25457);
xor U25537 (N_25537,N_25489,N_25425);
nor U25538 (N_25538,N_25394,N_25469);
nand U25539 (N_25539,N_25306,N_25365);
xnor U25540 (N_25540,N_25219,N_25384);
or U25541 (N_25541,N_25292,N_25269);
nand U25542 (N_25542,N_25348,N_25303);
nand U25543 (N_25543,N_25300,N_25293);
xnor U25544 (N_25544,N_25485,N_25343);
or U25545 (N_25545,N_25386,N_25427);
and U25546 (N_25546,N_25253,N_25266);
and U25547 (N_25547,N_25354,N_25496);
or U25548 (N_25548,N_25430,N_25420);
nor U25549 (N_25549,N_25271,N_25232);
or U25550 (N_25550,N_25461,N_25298);
xnor U25551 (N_25551,N_25265,N_25295);
xnor U25552 (N_25552,N_25334,N_25497);
or U25553 (N_25553,N_25409,N_25262);
xor U25554 (N_25554,N_25339,N_25305);
and U25555 (N_25555,N_25302,N_25458);
and U25556 (N_25556,N_25214,N_25326);
xnor U25557 (N_25557,N_25249,N_25388);
and U25558 (N_25558,N_25297,N_25445);
nand U25559 (N_25559,N_25406,N_25364);
and U25560 (N_25560,N_25478,N_25281);
or U25561 (N_25561,N_25323,N_25301);
or U25562 (N_25562,N_25236,N_25309);
xor U25563 (N_25563,N_25358,N_25475);
nor U25564 (N_25564,N_25235,N_25337);
or U25565 (N_25565,N_25476,N_25216);
nor U25566 (N_25566,N_25402,N_25452);
and U25567 (N_25567,N_25383,N_25482);
xor U25568 (N_25568,N_25213,N_25234);
nand U25569 (N_25569,N_25401,N_25200);
or U25570 (N_25570,N_25382,N_25436);
xor U25571 (N_25571,N_25288,N_25240);
xor U25572 (N_25572,N_25403,N_25215);
nor U25573 (N_25573,N_25468,N_25313);
and U25574 (N_25574,N_25283,N_25212);
and U25575 (N_25575,N_25464,N_25290);
nor U25576 (N_25576,N_25350,N_25462);
xnor U25577 (N_25577,N_25433,N_25227);
and U25578 (N_25578,N_25487,N_25338);
xnor U25579 (N_25579,N_25419,N_25342);
and U25580 (N_25580,N_25387,N_25280);
nor U25581 (N_25581,N_25327,N_25391);
and U25582 (N_25582,N_25285,N_25321);
nand U25583 (N_25583,N_25398,N_25432);
nand U25584 (N_25584,N_25488,N_25493);
xnor U25585 (N_25585,N_25448,N_25204);
and U25586 (N_25586,N_25463,N_25446);
and U25587 (N_25587,N_25460,N_25480);
nand U25588 (N_25588,N_25435,N_25375);
nor U25589 (N_25589,N_25376,N_25206);
or U25590 (N_25590,N_25286,N_25344);
or U25591 (N_25591,N_25340,N_25261);
and U25592 (N_25592,N_25331,N_25426);
or U25593 (N_25593,N_25294,N_25422);
or U25594 (N_25594,N_25447,N_25228);
or U25595 (N_25595,N_25252,N_25251);
xnor U25596 (N_25596,N_25455,N_25379);
or U25597 (N_25597,N_25415,N_25247);
nand U25598 (N_25598,N_25381,N_25270);
or U25599 (N_25599,N_25471,N_25267);
or U25600 (N_25600,N_25250,N_25257);
and U25601 (N_25601,N_25367,N_25400);
nor U25602 (N_25602,N_25410,N_25314);
xor U25603 (N_25603,N_25453,N_25449);
nand U25604 (N_25604,N_25353,N_25417);
nor U25605 (N_25605,N_25316,N_25441);
or U25606 (N_25606,N_25225,N_25450);
and U25607 (N_25607,N_25371,N_25491);
and U25608 (N_25608,N_25291,N_25259);
or U25609 (N_25609,N_25287,N_25260);
and U25610 (N_25610,N_25254,N_25264);
nand U25611 (N_25611,N_25263,N_25201);
and U25612 (N_25612,N_25345,N_25439);
nor U25613 (N_25613,N_25431,N_25369);
nor U25614 (N_25614,N_25404,N_25355);
nor U25615 (N_25615,N_25465,N_25318);
nor U25616 (N_25616,N_25407,N_25413);
xor U25617 (N_25617,N_25322,N_25312);
nor U25618 (N_25618,N_25473,N_25481);
or U25619 (N_25619,N_25399,N_25230);
nor U25620 (N_25620,N_25324,N_25492);
nand U25621 (N_25621,N_25329,N_25467);
or U25622 (N_25622,N_25272,N_25341);
or U25623 (N_25623,N_25275,N_25424);
xnor U25624 (N_25624,N_25418,N_25203);
nor U25625 (N_25625,N_25377,N_25437);
or U25626 (N_25626,N_25310,N_25349);
and U25627 (N_25627,N_25242,N_25366);
nor U25628 (N_25628,N_25276,N_25352);
nand U25629 (N_25629,N_25357,N_25209);
nand U25630 (N_25630,N_25239,N_25211);
and U25631 (N_25631,N_25218,N_25499);
and U25632 (N_25632,N_25308,N_25456);
nand U25633 (N_25633,N_25273,N_25282);
nand U25634 (N_25634,N_25279,N_25245);
nor U25635 (N_25635,N_25347,N_25307);
and U25636 (N_25636,N_25208,N_25299);
or U25637 (N_25637,N_25363,N_25248);
and U25638 (N_25638,N_25356,N_25494);
nor U25639 (N_25639,N_25317,N_25221);
nand U25640 (N_25640,N_25466,N_25231);
xor U25641 (N_25641,N_25233,N_25361);
nand U25642 (N_25642,N_25226,N_25392);
or U25643 (N_25643,N_25315,N_25217);
or U25644 (N_25644,N_25243,N_25378);
or U25645 (N_25645,N_25414,N_25396);
or U25646 (N_25646,N_25474,N_25440);
and U25647 (N_25647,N_25333,N_25319);
nor U25648 (N_25648,N_25210,N_25370);
xor U25649 (N_25649,N_25255,N_25477);
and U25650 (N_25650,N_25228,N_25252);
xor U25651 (N_25651,N_25236,N_25420);
xor U25652 (N_25652,N_25243,N_25349);
and U25653 (N_25653,N_25278,N_25471);
nor U25654 (N_25654,N_25244,N_25435);
or U25655 (N_25655,N_25203,N_25351);
and U25656 (N_25656,N_25490,N_25240);
or U25657 (N_25657,N_25333,N_25323);
nand U25658 (N_25658,N_25246,N_25354);
and U25659 (N_25659,N_25285,N_25247);
or U25660 (N_25660,N_25271,N_25484);
nand U25661 (N_25661,N_25264,N_25337);
or U25662 (N_25662,N_25383,N_25343);
nor U25663 (N_25663,N_25315,N_25467);
or U25664 (N_25664,N_25440,N_25200);
nor U25665 (N_25665,N_25452,N_25346);
nor U25666 (N_25666,N_25269,N_25420);
nor U25667 (N_25667,N_25361,N_25408);
nor U25668 (N_25668,N_25329,N_25376);
or U25669 (N_25669,N_25445,N_25301);
and U25670 (N_25670,N_25382,N_25234);
nor U25671 (N_25671,N_25313,N_25231);
and U25672 (N_25672,N_25252,N_25303);
nand U25673 (N_25673,N_25495,N_25391);
nand U25674 (N_25674,N_25326,N_25350);
xor U25675 (N_25675,N_25243,N_25306);
xor U25676 (N_25676,N_25377,N_25492);
nor U25677 (N_25677,N_25463,N_25402);
nor U25678 (N_25678,N_25300,N_25317);
and U25679 (N_25679,N_25322,N_25493);
or U25680 (N_25680,N_25440,N_25412);
or U25681 (N_25681,N_25380,N_25204);
nand U25682 (N_25682,N_25475,N_25301);
or U25683 (N_25683,N_25219,N_25246);
or U25684 (N_25684,N_25322,N_25264);
nand U25685 (N_25685,N_25316,N_25256);
and U25686 (N_25686,N_25457,N_25497);
or U25687 (N_25687,N_25373,N_25321);
nand U25688 (N_25688,N_25201,N_25276);
or U25689 (N_25689,N_25295,N_25477);
xor U25690 (N_25690,N_25253,N_25379);
xor U25691 (N_25691,N_25207,N_25445);
nor U25692 (N_25692,N_25476,N_25469);
nor U25693 (N_25693,N_25203,N_25470);
nand U25694 (N_25694,N_25339,N_25455);
nand U25695 (N_25695,N_25479,N_25213);
and U25696 (N_25696,N_25203,N_25347);
and U25697 (N_25697,N_25245,N_25419);
or U25698 (N_25698,N_25250,N_25322);
nor U25699 (N_25699,N_25351,N_25374);
nor U25700 (N_25700,N_25482,N_25381);
or U25701 (N_25701,N_25377,N_25428);
nand U25702 (N_25702,N_25242,N_25340);
nor U25703 (N_25703,N_25452,N_25443);
or U25704 (N_25704,N_25273,N_25488);
and U25705 (N_25705,N_25242,N_25265);
nand U25706 (N_25706,N_25453,N_25332);
nor U25707 (N_25707,N_25363,N_25336);
xnor U25708 (N_25708,N_25356,N_25201);
nor U25709 (N_25709,N_25281,N_25497);
and U25710 (N_25710,N_25388,N_25253);
xor U25711 (N_25711,N_25441,N_25448);
nand U25712 (N_25712,N_25458,N_25276);
or U25713 (N_25713,N_25263,N_25254);
and U25714 (N_25714,N_25372,N_25466);
nand U25715 (N_25715,N_25353,N_25442);
and U25716 (N_25716,N_25319,N_25446);
nor U25717 (N_25717,N_25250,N_25343);
nand U25718 (N_25718,N_25465,N_25441);
or U25719 (N_25719,N_25339,N_25360);
nand U25720 (N_25720,N_25239,N_25232);
nor U25721 (N_25721,N_25314,N_25356);
nand U25722 (N_25722,N_25329,N_25490);
or U25723 (N_25723,N_25372,N_25205);
and U25724 (N_25724,N_25267,N_25480);
xnor U25725 (N_25725,N_25426,N_25335);
xor U25726 (N_25726,N_25203,N_25434);
or U25727 (N_25727,N_25321,N_25303);
nand U25728 (N_25728,N_25368,N_25223);
nand U25729 (N_25729,N_25470,N_25370);
and U25730 (N_25730,N_25361,N_25495);
nor U25731 (N_25731,N_25235,N_25266);
and U25732 (N_25732,N_25489,N_25448);
nor U25733 (N_25733,N_25388,N_25425);
and U25734 (N_25734,N_25382,N_25308);
nor U25735 (N_25735,N_25495,N_25402);
nor U25736 (N_25736,N_25355,N_25346);
and U25737 (N_25737,N_25211,N_25404);
nand U25738 (N_25738,N_25353,N_25333);
and U25739 (N_25739,N_25373,N_25304);
nor U25740 (N_25740,N_25425,N_25226);
xor U25741 (N_25741,N_25337,N_25210);
or U25742 (N_25742,N_25378,N_25463);
xnor U25743 (N_25743,N_25450,N_25271);
or U25744 (N_25744,N_25340,N_25427);
nand U25745 (N_25745,N_25313,N_25385);
xnor U25746 (N_25746,N_25299,N_25206);
nand U25747 (N_25747,N_25356,N_25469);
and U25748 (N_25748,N_25413,N_25302);
xor U25749 (N_25749,N_25326,N_25256);
or U25750 (N_25750,N_25400,N_25426);
and U25751 (N_25751,N_25317,N_25224);
or U25752 (N_25752,N_25299,N_25341);
nor U25753 (N_25753,N_25485,N_25358);
nor U25754 (N_25754,N_25444,N_25410);
and U25755 (N_25755,N_25363,N_25462);
and U25756 (N_25756,N_25457,N_25221);
and U25757 (N_25757,N_25331,N_25215);
and U25758 (N_25758,N_25324,N_25329);
or U25759 (N_25759,N_25405,N_25493);
xor U25760 (N_25760,N_25308,N_25421);
nand U25761 (N_25761,N_25461,N_25212);
nor U25762 (N_25762,N_25249,N_25251);
nor U25763 (N_25763,N_25261,N_25388);
xnor U25764 (N_25764,N_25232,N_25215);
and U25765 (N_25765,N_25440,N_25405);
and U25766 (N_25766,N_25237,N_25441);
or U25767 (N_25767,N_25228,N_25337);
and U25768 (N_25768,N_25206,N_25387);
nand U25769 (N_25769,N_25492,N_25496);
nand U25770 (N_25770,N_25330,N_25443);
and U25771 (N_25771,N_25386,N_25421);
xnor U25772 (N_25772,N_25491,N_25274);
xnor U25773 (N_25773,N_25304,N_25470);
xnor U25774 (N_25774,N_25225,N_25406);
nand U25775 (N_25775,N_25242,N_25395);
or U25776 (N_25776,N_25249,N_25370);
nor U25777 (N_25777,N_25369,N_25237);
nand U25778 (N_25778,N_25261,N_25328);
or U25779 (N_25779,N_25295,N_25298);
or U25780 (N_25780,N_25419,N_25207);
xnor U25781 (N_25781,N_25485,N_25353);
and U25782 (N_25782,N_25285,N_25395);
or U25783 (N_25783,N_25327,N_25267);
xor U25784 (N_25784,N_25272,N_25267);
nor U25785 (N_25785,N_25306,N_25272);
nand U25786 (N_25786,N_25415,N_25399);
nand U25787 (N_25787,N_25251,N_25458);
or U25788 (N_25788,N_25375,N_25441);
nor U25789 (N_25789,N_25347,N_25460);
or U25790 (N_25790,N_25472,N_25221);
nand U25791 (N_25791,N_25224,N_25352);
nand U25792 (N_25792,N_25323,N_25496);
or U25793 (N_25793,N_25202,N_25280);
nand U25794 (N_25794,N_25449,N_25202);
and U25795 (N_25795,N_25442,N_25446);
nand U25796 (N_25796,N_25262,N_25236);
and U25797 (N_25797,N_25223,N_25456);
nor U25798 (N_25798,N_25351,N_25262);
or U25799 (N_25799,N_25368,N_25425);
nand U25800 (N_25800,N_25764,N_25695);
or U25801 (N_25801,N_25520,N_25798);
nand U25802 (N_25802,N_25788,N_25782);
xnor U25803 (N_25803,N_25654,N_25573);
or U25804 (N_25804,N_25688,N_25507);
xor U25805 (N_25805,N_25706,N_25601);
nand U25806 (N_25806,N_25506,N_25754);
and U25807 (N_25807,N_25722,N_25578);
and U25808 (N_25808,N_25748,N_25550);
and U25809 (N_25809,N_25567,N_25770);
nor U25810 (N_25810,N_25576,N_25628);
and U25811 (N_25811,N_25787,N_25681);
or U25812 (N_25812,N_25703,N_25684);
nand U25813 (N_25813,N_25635,N_25715);
or U25814 (N_25814,N_25501,N_25517);
or U25815 (N_25815,N_25526,N_25630);
xor U25816 (N_25816,N_25699,N_25645);
and U25817 (N_25817,N_25707,N_25780);
nand U25818 (N_25818,N_25740,N_25799);
and U25819 (N_25819,N_25647,N_25757);
nor U25820 (N_25820,N_25562,N_25784);
or U25821 (N_25821,N_25708,N_25527);
and U25822 (N_25822,N_25551,N_25587);
nand U25823 (N_25823,N_25514,N_25646);
or U25824 (N_25824,N_25679,N_25563);
nor U25825 (N_25825,N_25687,N_25714);
xor U25826 (N_25826,N_25720,N_25543);
and U25827 (N_25827,N_25656,N_25553);
or U25828 (N_25828,N_25602,N_25653);
nor U25829 (N_25829,N_25540,N_25724);
and U25830 (N_25830,N_25739,N_25505);
xor U25831 (N_25831,N_25579,N_25648);
nor U25832 (N_25832,N_25660,N_25795);
nor U25833 (N_25833,N_25552,N_25618);
xor U25834 (N_25834,N_25600,N_25560);
nor U25835 (N_25835,N_25522,N_25697);
nor U25836 (N_25836,N_25756,N_25556);
xor U25837 (N_25837,N_25592,N_25531);
nor U25838 (N_25838,N_25557,N_25595);
and U25839 (N_25839,N_25629,N_25700);
nand U25840 (N_25840,N_25752,N_25564);
and U25841 (N_25841,N_25512,N_25528);
xor U25842 (N_25842,N_25670,N_25738);
and U25843 (N_25843,N_25554,N_25589);
nor U25844 (N_25844,N_25650,N_25736);
xor U25845 (N_25845,N_25685,N_25741);
or U25846 (N_25846,N_25668,N_25723);
and U25847 (N_25847,N_25755,N_25559);
nand U25848 (N_25848,N_25636,N_25524);
or U25849 (N_25849,N_25642,N_25544);
nor U25850 (N_25850,N_25725,N_25539);
nand U25851 (N_25851,N_25605,N_25521);
and U25852 (N_25852,N_25638,N_25655);
and U25853 (N_25853,N_25581,N_25588);
or U25854 (N_25854,N_25745,N_25504);
or U25855 (N_25855,N_25509,N_25682);
or U25856 (N_25856,N_25769,N_25611);
nand U25857 (N_25857,N_25730,N_25675);
nor U25858 (N_25858,N_25500,N_25713);
or U25859 (N_25859,N_25767,N_25689);
and U25860 (N_25860,N_25674,N_25624);
or U25861 (N_25861,N_25594,N_25606);
or U25862 (N_25862,N_25790,N_25536);
nor U25863 (N_25863,N_25542,N_25758);
and U25864 (N_25864,N_25693,N_25533);
and U25865 (N_25865,N_25572,N_25609);
xnor U25866 (N_25866,N_25603,N_25786);
or U25867 (N_25867,N_25596,N_25510);
nor U25868 (N_25868,N_25623,N_25663);
xnor U25869 (N_25869,N_25515,N_25779);
and U25870 (N_25870,N_25761,N_25791);
or U25871 (N_25871,N_25625,N_25731);
nor U25872 (N_25872,N_25718,N_25537);
or U25873 (N_25873,N_25657,N_25622);
nand U25874 (N_25874,N_25619,N_25793);
nand U25875 (N_25875,N_25705,N_25669);
nor U25876 (N_25876,N_25640,N_25701);
xor U25877 (N_25877,N_25570,N_25667);
xnor U25878 (N_25878,N_25749,N_25532);
and U25879 (N_25879,N_25571,N_25727);
or U25880 (N_25880,N_25734,N_25585);
nor U25881 (N_25881,N_25702,N_25746);
and U25882 (N_25882,N_25565,N_25765);
xnor U25883 (N_25883,N_25677,N_25789);
nor U25884 (N_25884,N_25661,N_25644);
nand U25885 (N_25885,N_25586,N_25781);
and U25886 (N_25886,N_25568,N_25632);
nand U25887 (N_25887,N_25704,N_25709);
and U25888 (N_25888,N_25508,N_25743);
nand U25889 (N_25889,N_25582,N_25538);
and U25890 (N_25890,N_25530,N_25549);
nor U25891 (N_25891,N_25664,N_25523);
and U25892 (N_25892,N_25785,N_25771);
nand U25893 (N_25893,N_25692,N_25658);
nand U25894 (N_25894,N_25759,N_25776);
or U25895 (N_25895,N_25732,N_25691);
nand U25896 (N_25896,N_25659,N_25721);
xnor U25897 (N_25897,N_25607,N_25778);
nand U25898 (N_25898,N_25649,N_25735);
nand U25899 (N_25899,N_25614,N_25729);
or U25900 (N_25900,N_25717,N_25598);
and U25901 (N_25901,N_25604,N_25676);
nand U25902 (N_25902,N_25580,N_25555);
xnor U25903 (N_25903,N_25751,N_25643);
xnor U25904 (N_25904,N_25698,N_25627);
xnor U25905 (N_25905,N_25792,N_25597);
nand U25906 (N_25906,N_25516,N_25615);
and U25907 (N_25907,N_25558,N_25548);
nand U25908 (N_25908,N_25626,N_25513);
nand U25909 (N_25909,N_25584,N_25546);
nor U25910 (N_25910,N_25535,N_25742);
or U25911 (N_25911,N_25719,N_25621);
and U25912 (N_25912,N_25529,N_25613);
nor U25913 (N_25913,N_25577,N_25634);
or U25914 (N_25914,N_25637,N_25561);
and U25915 (N_25915,N_25662,N_25760);
and U25916 (N_25916,N_25690,N_25511);
nand U25917 (N_25917,N_25633,N_25737);
nor U25918 (N_25918,N_25794,N_25616);
or U25919 (N_25919,N_25744,N_25686);
nand U25920 (N_25920,N_25710,N_25566);
and U25921 (N_25921,N_25774,N_25569);
and U25922 (N_25922,N_25620,N_25575);
nor U25923 (N_25923,N_25672,N_25639);
nand U25924 (N_25924,N_25518,N_25651);
and U25925 (N_25925,N_25762,N_25673);
nor U25926 (N_25926,N_25733,N_25631);
nand U25927 (N_25927,N_25753,N_25591);
nand U25928 (N_25928,N_25502,N_25680);
xor U25929 (N_25929,N_25763,N_25750);
or U25930 (N_25930,N_25711,N_25666);
and U25931 (N_25931,N_25590,N_25574);
xor U25932 (N_25932,N_25547,N_25797);
and U25933 (N_25933,N_25503,N_25772);
and U25934 (N_25934,N_25641,N_25777);
nand U25935 (N_25935,N_25652,N_25768);
and U25936 (N_25936,N_25726,N_25747);
xor U25937 (N_25937,N_25696,N_25665);
nor U25938 (N_25938,N_25612,N_25716);
nor U25939 (N_25939,N_25541,N_25519);
nor U25940 (N_25940,N_25617,N_25671);
nor U25941 (N_25941,N_25728,N_25712);
and U25942 (N_25942,N_25783,N_25796);
xnor U25943 (N_25943,N_25599,N_25773);
xnor U25944 (N_25944,N_25683,N_25610);
and U25945 (N_25945,N_25593,N_25583);
xor U25946 (N_25946,N_25766,N_25678);
and U25947 (N_25947,N_25525,N_25694);
and U25948 (N_25948,N_25534,N_25775);
xnor U25949 (N_25949,N_25545,N_25608);
nand U25950 (N_25950,N_25679,N_25764);
xnor U25951 (N_25951,N_25657,N_25710);
and U25952 (N_25952,N_25615,N_25657);
xor U25953 (N_25953,N_25674,N_25504);
nor U25954 (N_25954,N_25754,N_25778);
and U25955 (N_25955,N_25674,N_25511);
xnor U25956 (N_25956,N_25743,N_25632);
and U25957 (N_25957,N_25541,N_25632);
and U25958 (N_25958,N_25555,N_25701);
xnor U25959 (N_25959,N_25653,N_25571);
xnor U25960 (N_25960,N_25686,N_25575);
and U25961 (N_25961,N_25712,N_25595);
nand U25962 (N_25962,N_25705,N_25753);
or U25963 (N_25963,N_25534,N_25637);
nand U25964 (N_25964,N_25613,N_25669);
or U25965 (N_25965,N_25741,N_25523);
and U25966 (N_25966,N_25534,N_25624);
nand U25967 (N_25967,N_25539,N_25661);
nor U25968 (N_25968,N_25786,N_25726);
nand U25969 (N_25969,N_25711,N_25793);
nor U25970 (N_25970,N_25703,N_25719);
nand U25971 (N_25971,N_25526,N_25754);
or U25972 (N_25972,N_25548,N_25557);
xnor U25973 (N_25973,N_25614,N_25526);
nor U25974 (N_25974,N_25769,N_25596);
nand U25975 (N_25975,N_25719,N_25714);
and U25976 (N_25976,N_25576,N_25559);
and U25977 (N_25977,N_25782,N_25583);
xnor U25978 (N_25978,N_25638,N_25544);
and U25979 (N_25979,N_25508,N_25683);
and U25980 (N_25980,N_25763,N_25507);
or U25981 (N_25981,N_25599,N_25537);
nor U25982 (N_25982,N_25646,N_25730);
nand U25983 (N_25983,N_25636,N_25729);
and U25984 (N_25984,N_25646,N_25786);
nand U25985 (N_25985,N_25675,N_25670);
or U25986 (N_25986,N_25587,N_25720);
and U25987 (N_25987,N_25770,N_25602);
and U25988 (N_25988,N_25588,N_25537);
or U25989 (N_25989,N_25645,N_25706);
nor U25990 (N_25990,N_25563,N_25572);
or U25991 (N_25991,N_25584,N_25728);
xor U25992 (N_25992,N_25611,N_25654);
and U25993 (N_25993,N_25631,N_25748);
xor U25994 (N_25994,N_25770,N_25614);
or U25995 (N_25995,N_25623,N_25651);
nand U25996 (N_25996,N_25631,N_25553);
or U25997 (N_25997,N_25662,N_25671);
nor U25998 (N_25998,N_25554,N_25619);
nand U25999 (N_25999,N_25769,N_25556);
nor U26000 (N_26000,N_25775,N_25788);
nand U26001 (N_26001,N_25635,N_25565);
xnor U26002 (N_26002,N_25569,N_25680);
xnor U26003 (N_26003,N_25629,N_25576);
nand U26004 (N_26004,N_25596,N_25793);
or U26005 (N_26005,N_25771,N_25726);
xnor U26006 (N_26006,N_25584,N_25559);
nor U26007 (N_26007,N_25541,N_25716);
xnor U26008 (N_26008,N_25553,N_25596);
nor U26009 (N_26009,N_25754,N_25620);
xor U26010 (N_26010,N_25568,N_25586);
nand U26011 (N_26011,N_25522,N_25601);
nand U26012 (N_26012,N_25702,N_25578);
nand U26013 (N_26013,N_25505,N_25588);
nor U26014 (N_26014,N_25539,N_25593);
and U26015 (N_26015,N_25621,N_25718);
and U26016 (N_26016,N_25703,N_25630);
xor U26017 (N_26017,N_25679,N_25632);
and U26018 (N_26018,N_25686,N_25615);
nor U26019 (N_26019,N_25608,N_25790);
and U26020 (N_26020,N_25551,N_25631);
nand U26021 (N_26021,N_25701,N_25654);
and U26022 (N_26022,N_25769,N_25554);
nor U26023 (N_26023,N_25781,N_25604);
and U26024 (N_26024,N_25588,N_25621);
nor U26025 (N_26025,N_25571,N_25520);
xnor U26026 (N_26026,N_25693,N_25647);
nand U26027 (N_26027,N_25615,N_25585);
nand U26028 (N_26028,N_25636,N_25614);
or U26029 (N_26029,N_25785,N_25676);
xnor U26030 (N_26030,N_25648,N_25541);
and U26031 (N_26031,N_25678,N_25689);
xor U26032 (N_26032,N_25548,N_25755);
nand U26033 (N_26033,N_25658,N_25744);
or U26034 (N_26034,N_25665,N_25611);
or U26035 (N_26035,N_25666,N_25648);
nand U26036 (N_26036,N_25722,N_25690);
xor U26037 (N_26037,N_25658,N_25522);
xor U26038 (N_26038,N_25714,N_25641);
nand U26039 (N_26039,N_25628,N_25600);
or U26040 (N_26040,N_25633,N_25734);
and U26041 (N_26041,N_25585,N_25755);
or U26042 (N_26042,N_25597,N_25736);
or U26043 (N_26043,N_25545,N_25723);
and U26044 (N_26044,N_25539,N_25783);
or U26045 (N_26045,N_25533,N_25528);
nor U26046 (N_26046,N_25795,N_25566);
nor U26047 (N_26047,N_25785,N_25702);
nand U26048 (N_26048,N_25656,N_25731);
nand U26049 (N_26049,N_25530,N_25720);
and U26050 (N_26050,N_25767,N_25749);
xor U26051 (N_26051,N_25567,N_25685);
nor U26052 (N_26052,N_25612,N_25730);
xor U26053 (N_26053,N_25635,N_25606);
or U26054 (N_26054,N_25576,N_25593);
nor U26055 (N_26055,N_25751,N_25648);
xor U26056 (N_26056,N_25797,N_25636);
nand U26057 (N_26057,N_25668,N_25688);
xnor U26058 (N_26058,N_25573,N_25595);
and U26059 (N_26059,N_25799,N_25789);
nor U26060 (N_26060,N_25560,N_25590);
nand U26061 (N_26061,N_25698,N_25686);
xnor U26062 (N_26062,N_25523,N_25520);
or U26063 (N_26063,N_25789,N_25608);
and U26064 (N_26064,N_25556,N_25526);
and U26065 (N_26065,N_25605,N_25714);
and U26066 (N_26066,N_25679,N_25683);
or U26067 (N_26067,N_25568,N_25785);
xor U26068 (N_26068,N_25750,N_25637);
and U26069 (N_26069,N_25788,N_25587);
xnor U26070 (N_26070,N_25518,N_25640);
and U26071 (N_26071,N_25589,N_25624);
or U26072 (N_26072,N_25613,N_25521);
nand U26073 (N_26073,N_25676,N_25731);
xnor U26074 (N_26074,N_25773,N_25784);
and U26075 (N_26075,N_25523,N_25586);
and U26076 (N_26076,N_25761,N_25684);
xnor U26077 (N_26077,N_25737,N_25703);
xor U26078 (N_26078,N_25617,N_25652);
and U26079 (N_26079,N_25581,N_25602);
nor U26080 (N_26080,N_25737,N_25712);
xnor U26081 (N_26081,N_25646,N_25647);
or U26082 (N_26082,N_25740,N_25768);
xor U26083 (N_26083,N_25764,N_25655);
or U26084 (N_26084,N_25688,N_25735);
xnor U26085 (N_26085,N_25736,N_25688);
nand U26086 (N_26086,N_25629,N_25748);
nor U26087 (N_26087,N_25696,N_25630);
nor U26088 (N_26088,N_25585,N_25504);
nor U26089 (N_26089,N_25767,N_25729);
or U26090 (N_26090,N_25584,N_25625);
xnor U26091 (N_26091,N_25664,N_25778);
and U26092 (N_26092,N_25630,N_25796);
or U26093 (N_26093,N_25645,N_25556);
nand U26094 (N_26094,N_25660,N_25631);
nand U26095 (N_26095,N_25714,N_25600);
or U26096 (N_26096,N_25629,N_25631);
xor U26097 (N_26097,N_25532,N_25600);
nor U26098 (N_26098,N_25617,N_25530);
nor U26099 (N_26099,N_25544,N_25509);
xnor U26100 (N_26100,N_25957,N_26008);
xor U26101 (N_26101,N_25917,N_25853);
or U26102 (N_26102,N_25998,N_25982);
nand U26103 (N_26103,N_25800,N_26076);
and U26104 (N_26104,N_25929,N_25989);
nand U26105 (N_26105,N_25805,N_26056);
nor U26106 (N_26106,N_25804,N_25943);
xor U26107 (N_26107,N_26025,N_26071);
nand U26108 (N_26108,N_26005,N_26094);
or U26109 (N_26109,N_26060,N_26037);
xor U26110 (N_26110,N_25988,N_25911);
nand U26111 (N_26111,N_25908,N_25938);
and U26112 (N_26112,N_25833,N_26068);
xnor U26113 (N_26113,N_25986,N_25876);
xor U26114 (N_26114,N_25885,N_25803);
and U26115 (N_26115,N_26041,N_25958);
xnor U26116 (N_26116,N_26012,N_25900);
nor U26117 (N_26117,N_25994,N_26055);
nor U26118 (N_26118,N_26024,N_26023);
nor U26119 (N_26119,N_25874,N_26043);
nor U26120 (N_26120,N_25906,N_26017);
nor U26121 (N_26121,N_26007,N_26011);
and U26122 (N_26122,N_25960,N_25858);
or U26123 (N_26123,N_26001,N_25901);
nand U26124 (N_26124,N_26061,N_26085);
nand U26125 (N_26125,N_25930,N_25813);
nor U26126 (N_26126,N_25879,N_25965);
nand U26127 (N_26127,N_25814,N_26096);
or U26128 (N_26128,N_25851,N_25864);
and U26129 (N_26129,N_26033,N_25822);
nand U26130 (N_26130,N_25875,N_26045);
xor U26131 (N_26131,N_25920,N_26057);
nor U26132 (N_26132,N_25999,N_25831);
and U26133 (N_26133,N_25827,N_26099);
and U26134 (N_26134,N_26042,N_25954);
nor U26135 (N_26135,N_25832,N_26063);
nand U26136 (N_26136,N_25862,N_25997);
nor U26137 (N_26137,N_26079,N_25990);
and U26138 (N_26138,N_25889,N_25870);
nand U26139 (N_26139,N_25896,N_26064);
xnor U26140 (N_26140,N_26020,N_25919);
xnor U26141 (N_26141,N_26031,N_25849);
or U26142 (N_26142,N_25823,N_25860);
xor U26143 (N_26143,N_26027,N_25944);
and U26144 (N_26144,N_25946,N_25970);
xor U26145 (N_26145,N_25809,N_26000);
xor U26146 (N_26146,N_25839,N_25921);
nand U26147 (N_26147,N_26081,N_25909);
nand U26148 (N_26148,N_25941,N_25976);
nand U26149 (N_26149,N_25923,N_26036);
and U26150 (N_26150,N_25977,N_25895);
nor U26151 (N_26151,N_25980,N_26082);
xor U26152 (N_26152,N_26014,N_25955);
nand U26153 (N_26153,N_26016,N_26087);
nand U26154 (N_26154,N_26052,N_26044);
nand U26155 (N_26155,N_25825,N_25968);
xor U26156 (N_26156,N_25863,N_25924);
or U26157 (N_26157,N_26002,N_26003);
nor U26158 (N_26158,N_25956,N_25973);
or U26159 (N_26159,N_25892,N_25835);
nand U26160 (N_26160,N_25945,N_26088);
or U26161 (N_26161,N_25811,N_26073);
nor U26162 (N_26162,N_25869,N_25888);
nor U26163 (N_26163,N_25852,N_25806);
xor U26164 (N_26164,N_25812,N_25848);
and U26165 (N_26165,N_25951,N_25912);
or U26166 (N_26166,N_26010,N_26078);
nand U26167 (N_26167,N_25995,N_26046);
nand U26168 (N_26168,N_25878,N_25850);
xor U26169 (N_26169,N_25873,N_25981);
xor U26170 (N_26170,N_25807,N_25983);
nand U26171 (N_26171,N_25828,N_25926);
or U26172 (N_26172,N_25934,N_26048);
nand U26173 (N_26173,N_25959,N_26026);
and U26174 (N_26174,N_26009,N_25841);
nand U26175 (N_26175,N_25867,N_26067);
nor U26176 (N_26176,N_25872,N_26015);
nor U26177 (N_26177,N_25819,N_25861);
xnor U26178 (N_26178,N_26053,N_25845);
and U26179 (N_26179,N_25836,N_26021);
nand U26180 (N_26180,N_25910,N_25880);
and U26181 (N_26181,N_26098,N_25846);
nand U26182 (N_26182,N_25890,N_26097);
nand U26183 (N_26183,N_26080,N_26075);
xnor U26184 (N_26184,N_26038,N_26059);
xor U26185 (N_26185,N_25843,N_25844);
or U26186 (N_26186,N_25933,N_26047);
and U26187 (N_26187,N_26070,N_25810);
and U26188 (N_26188,N_25935,N_25916);
and U26189 (N_26189,N_25840,N_25979);
xnor U26190 (N_26190,N_26030,N_25991);
and U26191 (N_26191,N_26062,N_25886);
and U26192 (N_26192,N_25818,N_26051);
and U26193 (N_26193,N_25914,N_26049);
xnor U26194 (N_26194,N_26035,N_25975);
nand U26195 (N_26195,N_26066,N_25974);
and U26196 (N_26196,N_25996,N_25838);
or U26197 (N_26197,N_26032,N_25820);
nand U26198 (N_26198,N_25992,N_25928);
or U26199 (N_26199,N_26029,N_25817);
xor U26200 (N_26200,N_26006,N_25834);
xnor U26201 (N_26201,N_25984,N_25902);
nor U26202 (N_26202,N_25855,N_25987);
and U26203 (N_26203,N_25967,N_26091);
nand U26204 (N_26204,N_25932,N_25899);
nor U26205 (N_26205,N_25942,N_25801);
xor U26206 (N_26206,N_25815,N_26054);
xnor U26207 (N_26207,N_25952,N_26074);
nand U26208 (N_26208,N_25925,N_25821);
xor U26209 (N_26209,N_25859,N_26069);
xor U26210 (N_26210,N_25842,N_25830);
or U26211 (N_26211,N_25816,N_26022);
nand U26212 (N_26212,N_25887,N_26058);
and U26213 (N_26213,N_25894,N_25856);
nor U26214 (N_26214,N_26086,N_25918);
and U26215 (N_26215,N_25915,N_25966);
xor U26216 (N_26216,N_25897,N_25883);
xor U26217 (N_26217,N_25950,N_25847);
nor U26218 (N_26218,N_25931,N_26095);
and U26219 (N_26219,N_25907,N_26077);
or U26220 (N_26220,N_25985,N_26004);
xnor U26221 (N_26221,N_25877,N_25882);
nand U26222 (N_26222,N_26083,N_25808);
or U26223 (N_26223,N_25868,N_25940);
nand U26224 (N_26224,N_26039,N_25871);
nor U26225 (N_26225,N_26018,N_25898);
and U26226 (N_26226,N_26028,N_25824);
nor U26227 (N_26227,N_25893,N_25837);
nand U26228 (N_26228,N_26093,N_25962);
and U26229 (N_26229,N_26089,N_25963);
nand U26230 (N_26230,N_26013,N_25971);
xnor U26231 (N_26231,N_26019,N_25826);
nand U26232 (N_26232,N_26040,N_25961);
nor U26233 (N_26233,N_25927,N_25953);
nor U26234 (N_26234,N_25922,N_25993);
and U26235 (N_26235,N_25857,N_25829);
or U26236 (N_26236,N_25913,N_25904);
xnor U26237 (N_26237,N_25936,N_26092);
nor U26238 (N_26238,N_25881,N_25903);
and U26239 (N_26239,N_25972,N_25948);
nor U26240 (N_26240,N_25891,N_25884);
and U26241 (N_26241,N_25969,N_25854);
or U26242 (N_26242,N_26034,N_25949);
or U26243 (N_26243,N_26084,N_25939);
nand U26244 (N_26244,N_26090,N_25978);
nor U26245 (N_26245,N_26065,N_25964);
nand U26246 (N_26246,N_25937,N_25865);
and U26247 (N_26247,N_25947,N_25802);
or U26248 (N_26248,N_25905,N_26072);
nor U26249 (N_26249,N_25866,N_26050);
or U26250 (N_26250,N_26008,N_25814);
nand U26251 (N_26251,N_25804,N_26082);
xnor U26252 (N_26252,N_25800,N_25801);
xor U26253 (N_26253,N_25985,N_25969);
nor U26254 (N_26254,N_25951,N_26003);
and U26255 (N_26255,N_25994,N_25980);
xor U26256 (N_26256,N_25915,N_25874);
xnor U26257 (N_26257,N_26011,N_26017);
and U26258 (N_26258,N_26057,N_25905);
or U26259 (N_26259,N_25835,N_25828);
xnor U26260 (N_26260,N_25802,N_26085);
or U26261 (N_26261,N_25907,N_25864);
nor U26262 (N_26262,N_26022,N_26012);
nor U26263 (N_26263,N_25953,N_25865);
nor U26264 (N_26264,N_25967,N_25915);
xnor U26265 (N_26265,N_25975,N_26022);
or U26266 (N_26266,N_26042,N_25809);
nand U26267 (N_26267,N_26025,N_25860);
and U26268 (N_26268,N_25904,N_25849);
nor U26269 (N_26269,N_25844,N_25939);
xor U26270 (N_26270,N_25838,N_25971);
or U26271 (N_26271,N_25992,N_25929);
nand U26272 (N_26272,N_25887,N_26059);
or U26273 (N_26273,N_26087,N_25854);
nor U26274 (N_26274,N_25872,N_25877);
xor U26275 (N_26275,N_25847,N_26023);
or U26276 (N_26276,N_26015,N_25906);
nor U26277 (N_26277,N_25925,N_25988);
or U26278 (N_26278,N_26099,N_25920);
nor U26279 (N_26279,N_25840,N_25818);
nand U26280 (N_26280,N_25856,N_25958);
or U26281 (N_26281,N_25813,N_25929);
nand U26282 (N_26282,N_25834,N_25981);
xnor U26283 (N_26283,N_25957,N_26058);
nand U26284 (N_26284,N_25954,N_26019);
nand U26285 (N_26285,N_26032,N_26060);
or U26286 (N_26286,N_25815,N_25884);
and U26287 (N_26287,N_26054,N_25854);
nand U26288 (N_26288,N_25911,N_25958);
nor U26289 (N_26289,N_26049,N_25858);
nor U26290 (N_26290,N_25842,N_26057);
and U26291 (N_26291,N_25990,N_25899);
xor U26292 (N_26292,N_25866,N_26033);
or U26293 (N_26293,N_26053,N_25918);
xor U26294 (N_26294,N_26002,N_25850);
xor U26295 (N_26295,N_26021,N_26006);
and U26296 (N_26296,N_25821,N_25951);
or U26297 (N_26297,N_26010,N_25831);
and U26298 (N_26298,N_26008,N_25951);
and U26299 (N_26299,N_25853,N_25902);
or U26300 (N_26300,N_25833,N_26002);
nand U26301 (N_26301,N_25967,N_25987);
or U26302 (N_26302,N_26076,N_26088);
nand U26303 (N_26303,N_25870,N_25935);
nand U26304 (N_26304,N_26009,N_26018);
and U26305 (N_26305,N_25958,N_25814);
or U26306 (N_26306,N_26035,N_25942);
and U26307 (N_26307,N_26025,N_25867);
nand U26308 (N_26308,N_26050,N_26034);
nand U26309 (N_26309,N_26007,N_25969);
nand U26310 (N_26310,N_26061,N_25920);
nand U26311 (N_26311,N_25862,N_26079);
xor U26312 (N_26312,N_25875,N_26068);
nor U26313 (N_26313,N_26014,N_25916);
nor U26314 (N_26314,N_25877,N_26095);
nand U26315 (N_26315,N_25916,N_25901);
nand U26316 (N_26316,N_25919,N_25836);
or U26317 (N_26317,N_26047,N_25815);
nand U26318 (N_26318,N_25933,N_25813);
and U26319 (N_26319,N_26097,N_25961);
xnor U26320 (N_26320,N_26052,N_26013);
nand U26321 (N_26321,N_26085,N_26003);
xnor U26322 (N_26322,N_25892,N_25858);
and U26323 (N_26323,N_25808,N_26008);
nor U26324 (N_26324,N_26005,N_26007);
nor U26325 (N_26325,N_25948,N_25982);
nor U26326 (N_26326,N_26077,N_25847);
or U26327 (N_26327,N_25951,N_26086);
nor U26328 (N_26328,N_25852,N_25894);
and U26329 (N_26329,N_25946,N_25993);
nor U26330 (N_26330,N_25966,N_25800);
nor U26331 (N_26331,N_25954,N_26029);
nor U26332 (N_26332,N_25821,N_26086);
nor U26333 (N_26333,N_25832,N_26018);
nor U26334 (N_26334,N_26020,N_25951);
or U26335 (N_26335,N_26028,N_26029);
nor U26336 (N_26336,N_25905,N_26022);
xnor U26337 (N_26337,N_25810,N_25968);
and U26338 (N_26338,N_25862,N_26092);
nor U26339 (N_26339,N_26029,N_25888);
nand U26340 (N_26340,N_26090,N_25905);
or U26341 (N_26341,N_26021,N_25873);
or U26342 (N_26342,N_26020,N_26036);
nand U26343 (N_26343,N_26090,N_25863);
xor U26344 (N_26344,N_25980,N_26054);
xnor U26345 (N_26345,N_25853,N_26001);
or U26346 (N_26346,N_26039,N_25864);
or U26347 (N_26347,N_25999,N_25855);
or U26348 (N_26348,N_26055,N_26003);
xor U26349 (N_26349,N_25858,N_25871);
nand U26350 (N_26350,N_25988,N_25833);
nor U26351 (N_26351,N_26044,N_25849);
nand U26352 (N_26352,N_26070,N_25884);
nand U26353 (N_26353,N_25899,N_26078);
xor U26354 (N_26354,N_26075,N_25982);
nand U26355 (N_26355,N_25872,N_26072);
nor U26356 (N_26356,N_25915,N_25977);
nor U26357 (N_26357,N_25974,N_26023);
and U26358 (N_26358,N_25837,N_26012);
nor U26359 (N_26359,N_26079,N_26018);
xor U26360 (N_26360,N_25907,N_25836);
and U26361 (N_26361,N_25988,N_25866);
and U26362 (N_26362,N_25804,N_25905);
xnor U26363 (N_26363,N_25872,N_26095);
or U26364 (N_26364,N_25856,N_26076);
nor U26365 (N_26365,N_26095,N_25801);
nand U26366 (N_26366,N_25885,N_26005);
nand U26367 (N_26367,N_25843,N_25879);
or U26368 (N_26368,N_25810,N_26067);
and U26369 (N_26369,N_25881,N_25915);
nand U26370 (N_26370,N_26077,N_26098);
xor U26371 (N_26371,N_25998,N_26056);
xnor U26372 (N_26372,N_25979,N_25973);
or U26373 (N_26373,N_25903,N_25961);
nand U26374 (N_26374,N_25861,N_26039);
or U26375 (N_26375,N_26033,N_26044);
nor U26376 (N_26376,N_25970,N_25841);
or U26377 (N_26377,N_25821,N_25942);
nand U26378 (N_26378,N_25804,N_25888);
nand U26379 (N_26379,N_25845,N_25873);
xnor U26380 (N_26380,N_25939,N_26052);
and U26381 (N_26381,N_25902,N_26042);
and U26382 (N_26382,N_25919,N_26065);
xor U26383 (N_26383,N_25836,N_25964);
nor U26384 (N_26384,N_25916,N_25804);
and U26385 (N_26385,N_26066,N_26002);
nor U26386 (N_26386,N_25968,N_25928);
nand U26387 (N_26387,N_25804,N_26004);
nor U26388 (N_26388,N_25915,N_26038);
xnor U26389 (N_26389,N_25906,N_25867);
xor U26390 (N_26390,N_25859,N_25975);
or U26391 (N_26391,N_26041,N_25886);
and U26392 (N_26392,N_25966,N_25977);
nor U26393 (N_26393,N_25817,N_25906);
nand U26394 (N_26394,N_25827,N_26030);
nor U26395 (N_26395,N_25900,N_26014);
nor U26396 (N_26396,N_25868,N_26093);
nor U26397 (N_26397,N_26014,N_25913);
nor U26398 (N_26398,N_25958,N_25842);
nor U26399 (N_26399,N_26053,N_26019);
xnor U26400 (N_26400,N_26159,N_26323);
nand U26401 (N_26401,N_26372,N_26324);
or U26402 (N_26402,N_26134,N_26359);
xor U26403 (N_26403,N_26137,N_26292);
and U26404 (N_26404,N_26332,N_26100);
and U26405 (N_26405,N_26380,N_26259);
xnor U26406 (N_26406,N_26310,N_26327);
xnor U26407 (N_26407,N_26382,N_26333);
xor U26408 (N_26408,N_26185,N_26144);
and U26409 (N_26409,N_26227,N_26352);
xor U26410 (N_26410,N_26188,N_26308);
and U26411 (N_26411,N_26285,N_26291);
nand U26412 (N_26412,N_26218,N_26373);
and U26413 (N_26413,N_26138,N_26167);
xor U26414 (N_26414,N_26153,N_26349);
or U26415 (N_26415,N_26160,N_26374);
and U26416 (N_26416,N_26395,N_26330);
nor U26417 (N_26417,N_26321,N_26271);
nor U26418 (N_26418,N_26265,N_26340);
xor U26419 (N_26419,N_26354,N_26126);
and U26420 (N_26420,N_26115,N_26216);
or U26421 (N_26421,N_26275,N_26398);
nor U26422 (N_26422,N_26256,N_26389);
xnor U26423 (N_26423,N_26225,N_26318);
nor U26424 (N_26424,N_26262,N_26128);
nand U26425 (N_26425,N_26257,N_26118);
nand U26426 (N_26426,N_26231,N_26127);
xor U26427 (N_26427,N_26252,N_26201);
or U26428 (N_26428,N_26103,N_26350);
and U26429 (N_26429,N_26136,N_26179);
or U26430 (N_26430,N_26379,N_26388);
nand U26431 (N_26431,N_26260,N_26233);
or U26432 (N_26432,N_26325,N_26183);
or U26433 (N_26433,N_26235,N_26375);
or U26434 (N_26434,N_26156,N_26197);
and U26435 (N_26435,N_26255,N_26391);
nand U26436 (N_26436,N_26173,N_26239);
xnor U26437 (N_26437,N_26152,N_26346);
xor U26438 (N_26438,N_26243,N_26345);
nor U26439 (N_26439,N_26151,N_26176);
nand U26440 (N_26440,N_26210,N_26172);
nor U26441 (N_26441,N_26129,N_26119);
or U26442 (N_26442,N_26338,N_26104);
nand U26443 (N_26443,N_26312,N_26224);
and U26444 (N_26444,N_26311,N_26170);
xor U26445 (N_26445,N_26278,N_26108);
nand U26446 (N_26446,N_26246,N_26303);
nand U26447 (N_26447,N_26378,N_26253);
nand U26448 (N_26448,N_26300,N_26288);
xor U26449 (N_26449,N_26133,N_26258);
nand U26450 (N_26450,N_26226,N_26281);
xor U26451 (N_26451,N_26299,N_26106);
and U26452 (N_26452,N_26397,N_26270);
or U26453 (N_26453,N_26229,N_26171);
or U26454 (N_26454,N_26364,N_26301);
and U26455 (N_26455,N_26187,N_26204);
nor U26456 (N_26456,N_26155,N_26272);
or U26457 (N_26457,N_26174,N_26290);
xor U26458 (N_26458,N_26337,N_26169);
xor U26459 (N_26459,N_26162,N_26360);
nor U26460 (N_26460,N_26396,N_26205);
xnor U26461 (N_26461,N_26353,N_26177);
nor U26462 (N_26462,N_26287,N_26390);
nand U26463 (N_26463,N_26236,N_26122);
or U26464 (N_26464,N_26112,N_26120);
and U26465 (N_26465,N_26101,N_26381);
nand U26466 (N_26466,N_26191,N_26211);
and U26467 (N_26467,N_26200,N_26363);
or U26468 (N_26468,N_26297,N_26307);
nand U26469 (N_26469,N_26215,N_26117);
xnor U26470 (N_26470,N_26219,N_26198);
and U26471 (N_26471,N_26322,N_26102);
nand U26472 (N_26472,N_26358,N_26336);
or U26473 (N_26473,N_26277,N_26348);
nand U26474 (N_26474,N_26341,N_26362);
nand U26475 (N_26475,N_26343,N_26139);
and U26476 (N_26476,N_26369,N_26165);
nor U26477 (N_26477,N_26241,N_26130);
xnor U26478 (N_26478,N_26266,N_26295);
nand U26479 (N_26479,N_26182,N_26367);
nor U26480 (N_26480,N_26280,N_26344);
nor U26481 (N_26481,N_26175,N_26304);
nand U26482 (N_26482,N_26357,N_26158);
and U26483 (N_26483,N_26193,N_26387);
or U26484 (N_26484,N_26249,N_26223);
and U26485 (N_26485,N_26315,N_26221);
xnor U26486 (N_26486,N_26161,N_26181);
nor U26487 (N_26487,N_26335,N_26244);
nor U26488 (N_26488,N_26124,N_26282);
xnor U26489 (N_26489,N_26296,N_26355);
and U26490 (N_26490,N_26109,N_26347);
or U26491 (N_26491,N_26157,N_26125);
xnor U26492 (N_26492,N_26196,N_26199);
and U26493 (N_26493,N_26328,N_26254);
and U26494 (N_26494,N_26293,N_26334);
and U26495 (N_26495,N_26248,N_26194);
xnor U26496 (N_26496,N_26356,N_26208);
and U26497 (N_26497,N_26230,N_26351);
and U26498 (N_26498,N_26143,N_26361);
and U26499 (N_26499,N_26142,N_26240);
or U26500 (N_26500,N_26377,N_26195);
nor U26501 (N_26501,N_26276,N_26365);
nor U26502 (N_26502,N_26213,N_26148);
nand U26503 (N_26503,N_26186,N_26393);
nor U26504 (N_26504,N_26313,N_26371);
nor U26505 (N_26505,N_26294,N_26309);
nor U26506 (N_26506,N_26279,N_26329);
nand U26507 (N_26507,N_26384,N_26189);
nand U26508 (N_26508,N_26298,N_26286);
or U26509 (N_26509,N_26146,N_26326);
and U26510 (N_26510,N_26247,N_26222);
nand U26511 (N_26511,N_26131,N_26164);
xor U26512 (N_26512,N_26209,N_26190);
xnor U26513 (N_26513,N_26261,N_26245);
nor U26514 (N_26514,N_26342,N_26132);
nor U26515 (N_26515,N_26386,N_26385);
nand U26516 (N_26516,N_26180,N_26220);
xnor U26517 (N_26517,N_26123,N_26317);
xnor U26518 (N_26518,N_26376,N_26392);
xor U26519 (N_26519,N_26394,N_26192);
nor U26520 (N_26520,N_26366,N_26263);
nor U26521 (N_26521,N_26141,N_26284);
xnor U26522 (N_26522,N_26368,N_26242);
xor U26523 (N_26523,N_26206,N_26163);
xor U26524 (N_26524,N_26203,N_26268);
or U26525 (N_26525,N_26114,N_26269);
xnor U26526 (N_26526,N_26237,N_26145);
xor U26527 (N_26527,N_26228,N_26184);
xor U26528 (N_26528,N_26399,N_26305);
and U26529 (N_26529,N_26154,N_26316);
and U26530 (N_26530,N_26168,N_26238);
nor U26531 (N_26531,N_26110,N_26178);
and U26532 (N_26532,N_26149,N_26302);
nand U26533 (N_26533,N_26207,N_26166);
nand U26534 (N_26534,N_26113,N_26234);
nor U26535 (N_26535,N_26370,N_26250);
xor U26536 (N_26536,N_26306,N_26116);
xor U26537 (N_26537,N_26232,N_26107);
nand U26538 (N_26538,N_26331,N_26217);
or U26539 (N_26539,N_26105,N_26264);
nand U26540 (N_26540,N_26267,N_26140);
nor U26541 (N_26541,N_26283,N_26289);
xnor U26542 (N_26542,N_26274,N_26212);
nand U26543 (N_26543,N_26273,N_26383);
nand U26544 (N_26544,N_26135,N_26150);
xor U26545 (N_26545,N_26202,N_26147);
nor U26546 (N_26546,N_26251,N_26214);
nand U26547 (N_26547,N_26111,N_26339);
nor U26548 (N_26548,N_26121,N_26320);
xnor U26549 (N_26549,N_26314,N_26319);
nor U26550 (N_26550,N_26134,N_26114);
and U26551 (N_26551,N_26234,N_26373);
or U26552 (N_26552,N_26377,N_26366);
nor U26553 (N_26553,N_26166,N_26279);
and U26554 (N_26554,N_26225,N_26102);
nand U26555 (N_26555,N_26201,N_26145);
or U26556 (N_26556,N_26339,N_26120);
xor U26557 (N_26557,N_26177,N_26382);
nand U26558 (N_26558,N_26171,N_26352);
nand U26559 (N_26559,N_26260,N_26333);
nor U26560 (N_26560,N_26248,N_26216);
xor U26561 (N_26561,N_26307,N_26389);
and U26562 (N_26562,N_26349,N_26388);
and U26563 (N_26563,N_26258,N_26176);
xnor U26564 (N_26564,N_26316,N_26226);
nand U26565 (N_26565,N_26349,N_26207);
or U26566 (N_26566,N_26384,N_26223);
nor U26567 (N_26567,N_26321,N_26310);
and U26568 (N_26568,N_26184,N_26298);
nand U26569 (N_26569,N_26348,N_26220);
nor U26570 (N_26570,N_26330,N_26155);
nor U26571 (N_26571,N_26348,N_26135);
xnor U26572 (N_26572,N_26183,N_26179);
or U26573 (N_26573,N_26289,N_26193);
nand U26574 (N_26574,N_26394,N_26214);
nor U26575 (N_26575,N_26166,N_26164);
nand U26576 (N_26576,N_26290,N_26170);
nand U26577 (N_26577,N_26181,N_26307);
and U26578 (N_26578,N_26366,N_26386);
and U26579 (N_26579,N_26126,N_26213);
xnor U26580 (N_26580,N_26189,N_26289);
or U26581 (N_26581,N_26338,N_26127);
nand U26582 (N_26582,N_26125,N_26350);
and U26583 (N_26583,N_26137,N_26395);
xnor U26584 (N_26584,N_26213,N_26243);
nand U26585 (N_26585,N_26257,N_26362);
and U26586 (N_26586,N_26347,N_26121);
and U26587 (N_26587,N_26194,N_26308);
xor U26588 (N_26588,N_26139,N_26163);
or U26589 (N_26589,N_26228,N_26279);
nor U26590 (N_26590,N_26384,N_26353);
and U26591 (N_26591,N_26181,N_26361);
xnor U26592 (N_26592,N_26244,N_26142);
xnor U26593 (N_26593,N_26396,N_26117);
or U26594 (N_26594,N_26320,N_26302);
nand U26595 (N_26595,N_26393,N_26107);
xnor U26596 (N_26596,N_26118,N_26304);
xnor U26597 (N_26597,N_26258,N_26320);
nand U26598 (N_26598,N_26303,N_26238);
or U26599 (N_26599,N_26224,N_26379);
or U26600 (N_26600,N_26366,N_26265);
nor U26601 (N_26601,N_26233,N_26140);
or U26602 (N_26602,N_26322,N_26172);
nand U26603 (N_26603,N_26184,N_26250);
nor U26604 (N_26604,N_26306,N_26372);
nand U26605 (N_26605,N_26304,N_26338);
xnor U26606 (N_26606,N_26266,N_26188);
and U26607 (N_26607,N_26236,N_26240);
xor U26608 (N_26608,N_26276,N_26399);
xnor U26609 (N_26609,N_26297,N_26276);
and U26610 (N_26610,N_26213,N_26256);
xnor U26611 (N_26611,N_26314,N_26174);
xor U26612 (N_26612,N_26113,N_26305);
xnor U26613 (N_26613,N_26347,N_26209);
nor U26614 (N_26614,N_26193,N_26262);
or U26615 (N_26615,N_26232,N_26311);
or U26616 (N_26616,N_26348,N_26182);
and U26617 (N_26617,N_26104,N_26130);
xor U26618 (N_26618,N_26198,N_26166);
nor U26619 (N_26619,N_26210,N_26264);
nand U26620 (N_26620,N_26291,N_26392);
nor U26621 (N_26621,N_26299,N_26136);
xnor U26622 (N_26622,N_26314,N_26335);
or U26623 (N_26623,N_26388,N_26129);
and U26624 (N_26624,N_26372,N_26187);
nor U26625 (N_26625,N_26328,N_26208);
or U26626 (N_26626,N_26180,N_26115);
nand U26627 (N_26627,N_26330,N_26242);
and U26628 (N_26628,N_26248,N_26192);
nor U26629 (N_26629,N_26182,N_26387);
and U26630 (N_26630,N_26199,N_26268);
nor U26631 (N_26631,N_26300,N_26317);
and U26632 (N_26632,N_26212,N_26210);
or U26633 (N_26633,N_26203,N_26271);
nor U26634 (N_26634,N_26190,N_26320);
nand U26635 (N_26635,N_26394,N_26255);
nand U26636 (N_26636,N_26124,N_26219);
xor U26637 (N_26637,N_26336,N_26289);
or U26638 (N_26638,N_26270,N_26367);
and U26639 (N_26639,N_26331,N_26157);
and U26640 (N_26640,N_26339,N_26182);
and U26641 (N_26641,N_26260,N_26112);
nand U26642 (N_26642,N_26231,N_26295);
or U26643 (N_26643,N_26161,N_26204);
xor U26644 (N_26644,N_26201,N_26222);
nand U26645 (N_26645,N_26252,N_26131);
nand U26646 (N_26646,N_26246,N_26164);
nand U26647 (N_26647,N_26157,N_26116);
and U26648 (N_26648,N_26379,N_26209);
and U26649 (N_26649,N_26150,N_26331);
and U26650 (N_26650,N_26175,N_26203);
and U26651 (N_26651,N_26222,N_26162);
or U26652 (N_26652,N_26107,N_26175);
nand U26653 (N_26653,N_26187,N_26173);
or U26654 (N_26654,N_26205,N_26310);
nor U26655 (N_26655,N_26221,N_26374);
or U26656 (N_26656,N_26181,N_26304);
and U26657 (N_26657,N_26141,N_26192);
nor U26658 (N_26658,N_26253,N_26212);
nand U26659 (N_26659,N_26329,N_26197);
nor U26660 (N_26660,N_26164,N_26185);
xnor U26661 (N_26661,N_26125,N_26310);
and U26662 (N_26662,N_26206,N_26232);
and U26663 (N_26663,N_26161,N_26194);
nor U26664 (N_26664,N_26252,N_26354);
and U26665 (N_26665,N_26171,N_26282);
nand U26666 (N_26666,N_26256,N_26148);
xnor U26667 (N_26667,N_26299,N_26263);
xor U26668 (N_26668,N_26331,N_26159);
xnor U26669 (N_26669,N_26183,N_26336);
xnor U26670 (N_26670,N_26201,N_26379);
xor U26671 (N_26671,N_26149,N_26140);
nor U26672 (N_26672,N_26337,N_26317);
and U26673 (N_26673,N_26327,N_26255);
nor U26674 (N_26674,N_26258,N_26315);
or U26675 (N_26675,N_26393,N_26167);
or U26676 (N_26676,N_26306,N_26328);
and U26677 (N_26677,N_26206,N_26198);
or U26678 (N_26678,N_26299,N_26228);
and U26679 (N_26679,N_26255,N_26229);
and U26680 (N_26680,N_26319,N_26126);
and U26681 (N_26681,N_26288,N_26317);
or U26682 (N_26682,N_26398,N_26167);
nand U26683 (N_26683,N_26129,N_26312);
xnor U26684 (N_26684,N_26177,N_26284);
xor U26685 (N_26685,N_26222,N_26281);
nor U26686 (N_26686,N_26257,N_26206);
nand U26687 (N_26687,N_26161,N_26307);
nand U26688 (N_26688,N_26117,N_26236);
and U26689 (N_26689,N_26244,N_26384);
nand U26690 (N_26690,N_26328,N_26131);
nor U26691 (N_26691,N_26201,N_26139);
nand U26692 (N_26692,N_26187,N_26381);
nor U26693 (N_26693,N_26126,N_26203);
or U26694 (N_26694,N_26232,N_26352);
or U26695 (N_26695,N_26226,N_26173);
xnor U26696 (N_26696,N_26128,N_26227);
nor U26697 (N_26697,N_26273,N_26298);
and U26698 (N_26698,N_26372,N_26380);
nand U26699 (N_26699,N_26324,N_26328);
or U26700 (N_26700,N_26682,N_26511);
and U26701 (N_26701,N_26505,N_26450);
xor U26702 (N_26702,N_26673,N_26421);
nand U26703 (N_26703,N_26545,N_26566);
and U26704 (N_26704,N_26423,N_26592);
and U26705 (N_26705,N_26596,N_26419);
or U26706 (N_26706,N_26430,N_26424);
nand U26707 (N_26707,N_26698,N_26409);
or U26708 (N_26708,N_26670,N_26535);
and U26709 (N_26709,N_26520,N_26401);
nand U26710 (N_26710,N_26671,N_26528);
xor U26711 (N_26711,N_26526,N_26668);
or U26712 (N_26712,N_26490,N_26561);
and U26713 (N_26713,N_26620,N_26532);
and U26714 (N_26714,N_26657,N_26597);
nand U26715 (N_26715,N_26694,N_26610);
or U26716 (N_26716,N_26496,N_26576);
and U26717 (N_26717,N_26619,N_26636);
or U26718 (N_26718,N_26529,N_26593);
nor U26719 (N_26719,N_26582,N_26574);
and U26720 (N_26720,N_26674,N_26443);
or U26721 (N_26721,N_26553,N_26590);
nand U26722 (N_26722,N_26500,N_26402);
or U26723 (N_26723,N_26512,N_26541);
xnor U26724 (N_26724,N_26523,N_26513);
xnor U26725 (N_26725,N_26426,N_26436);
and U26726 (N_26726,N_26648,N_26482);
nor U26727 (N_26727,N_26571,N_26570);
nand U26728 (N_26728,N_26493,N_26488);
nor U26729 (N_26729,N_26413,N_26689);
or U26730 (N_26730,N_26417,N_26609);
or U26731 (N_26731,N_26412,N_26525);
or U26732 (N_26732,N_26514,N_26696);
nand U26733 (N_26733,N_26481,N_26699);
or U26734 (N_26734,N_26618,N_26415);
nor U26735 (N_26735,N_26509,N_26400);
xnor U26736 (N_26736,N_26688,N_26598);
and U26737 (N_26737,N_26492,N_26621);
and U26738 (N_26738,N_26644,N_26465);
nand U26739 (N_26739,N_26418,N_26641);
or U26740 (N_26740,N_26558,N_26637);
and U26741 (N_26741,N_26608,N_26538);
or U26742 (N_26742,N_26403,N_26470);
xnor U26743 (N_26743,N_26414,N_26602);
xnor U26744 (N_26744,N_26678,N_26527);
or U26745 (N_26745,N_26647,N_26585);
xnor U26746 (N_26746,N_26444,N_26518);
and U26747 (N_26747,N_26676,N_26662);
nor U26748 (N_26748,N_26447,N_26448);
xnor U26749 (N_26749,N_26642,N_26564);
nor U26750 (N_26750,N_26568,N_26632);
and U26751 (N_26751,N_26587,N_26473);
nand U26752 (N_26752,N_26416,N_26449);
or U26753 (N_26753,N_26633,N_26581);
nand U26754 (N_26754,N_26562,N_26472);
xor U26755 (N_26755,N_26690,N_26476);
and U26756 (N_26756,N_26584,N_26677);
and U26757 (N_26757,N_26652,N_26557);
nor U26758 (N_26758,N_26654,N_26475);
nor U26759 (N_26759,N_26548,N_26517);
nand U26760 (N_26760,N_26580,N_26628);
xor U26761 (N_26761,N_26510,N_26563);
xnor U26762 (N_26762,N_26693,N_26630);
or U26763 (N_26763,N_26603,N_26589);
nor U26764 (N_26764,N_26626,N_26624);
nor U26765 (N_26765,N_26645,N_26604);
and U26766 (N_26766,N_26605,N_26495);
or U26767 (N_26767,N_26466,N_26462);
xnor U26768 (N_26768,N_26441,N_26429);
xor U26769 (N_26769,N_26464,N_26486);
nor U26770 (N_26770,N_26687,N_26600);
or U26771 (N_26771,N_26550,N_26506);
xnor U26772 (N_26772,N_26463,N_26504);
or U26773 (N_26773,N_26681,N_26667);
or U26774 (N_26774,N_26588,N_26404);
xor U26775 (N_26775,N_26573,N_26695);
nand U26776 (N_26776,N_26627,N_26485);
xnor U26777 (N_26777,N_26614,N_26543);
xnor U26778 (N_26778,N_26559,N_26546);
xnor U26779 (N_26779,N_26474,N_26459);
xnor U26780 (N_26780,N_26530,N_26643);
or U26781 (N_26781,N_26613,N_26461);
nor U26782 (N_26782,N_26531,N_26675);
nor U26783 (N_26783,N_26615,N_26544);
nor U26784 (N_26784,N_26640,N_26536);
nor U26785 (N_26785,N_26437,N_26487);
xor U26786 (N_26786,N_26438,N_26458);
xnor U26787 (N_26787,N_26494,N_26468);
or U26788 (N_26788,N_26554,N_26483);
and U26789 (N_26789,N_26623,N_26507);
or U26790 (N_26790,N_26469,N_26524);
or U26791 (N_26791,N_26655,N_26407);
or U26792 (N_26792,N_26425,N_26567);
or U26793 (N_26793,N_26497,N_26501);
and U26794 (N_26794,N_26442,N_26455);
xnor U26795 (N_26795,N_26478,N_26606);
and U26796 (N_26796,N_26622,N_26586);
or U26797 (N_26797,N_26601,N_26428);
or U26798 (N_26798,N_26612,N_26692);
xnor U26799 (N_26799,N_26542,N_26656);
nor U26800 (N_26800,N_26549,N_26499);
nand U26801 (N_26801,N_26491,N_26406);
and U26802 (N_26802,N_26522,N_26638);
or U26803 (N_26803,N_26569,N_26516);
xor U26804 (N_26804,N_26508,N_26467);
and U26805 (N_26805,N_26433,N_26456);
xnor U26806 (N_26806,N_26661,N_26539);
nand U26807 (N_26807,N_26555,N_26515);
nand U26808 (N_26808,N_26686,N_26540);
and U26809 (N_26809,N_26639,N_26680);
xor U26810 (N_26810,N_26471,N_26547);
nand U26811 (N_26811,N_26420,N_26408);
and U26812 (N_26812,N_26479,N_26440);
nor U26813 (N_26813,N_26594,N_26577);
and U26814 (N_26814,N_26669,N_26599);
or U26815 (N_26815,N_26560,N_26659);
and U26816 (N_26816,N_26663,N_26629);
and U26817 (N_26817,N_26651,N_26521);
nand U26818 (N_26818,N_26431,N_26583);
or U26819 (N_26819,N_26480,N_26672);
xor U26820 (N_26820,N_26446,N_26611);
xnor U26821 (N_26821,N_26435,N_26460);
or U26822 (N_26822,N_26405,N_26556);
and U26823 (N_26823,N_26665,N_26537);
or U26824 (N_26824,N_26595,N_26664);
nand U26825 (N_26825,N_26551,N_26650);
xor U26826 (N_26826,N_26533,N_26649);
xnor U26827 (N_26827,N_26578,N_26457);
or U26828 (N_26828,N_26679,N_26634);
nor U26829 (N_26829,N_26519,N_26452);
nor U26830 (N_26830,N_26616,N_26489);
and U26831 (N_26831,N_26411,N_26591);
nor U26832 (N_26832,N_26625,N_26498);
xor U26833 (N_26833,N_26502,N_26410);
or U26834 (N_26834,N_26422,N_26451);
nor U26835 (N_26835,N_26607,N_26660);
and U26836 (N_26836,N_26432,N_26635);
nand U26837 (N_26837,N_26579,N_26685);
nor U26838 (N_26838,N_26646,N_26477);
nor U26839 (N_26839,N_26691,N_26534);
nand U26840 (N_26840,N_26653,N_26658);
and U26841 (N_26841,N_26427,N_26439);
or U26842 (N_26842,N_26445,N_26684);
nor U26843 (N_26843,N_26666,N_26484);
or U26844 (N_26844,N_26575,N_26697);
or U26845 (N_26845,N_26565,N_26572);
xnor U26846 (N_26846,N_26503,N_26434);
nand U26847 (N_26847,N_26453,N_26617);
or U26848 (N_26848,N_26631,N_26552);
and U26849 (N_26849,N_26454,N_26683);
and U26850 (N_26850,N_26421,N_26682);
xor U26851 (N_26851,N_26446,N_26500);
and U26852 (N_26852,N_26485,N_26583);
xor U26853 (N_26853,N_26621,N_26580);
or U26854 (N_26854,N_26409,N_26619);
or U26855 (N_26855,N_26687,N_26672);
nor U26856 (N_26856,N_26505,N_26418);
and U26857 (N_26857,N_26502,N_26624);
or U26858 (N_26858,N_26549,N_26459);
xnor U26859 (N_26859,N_26667,N_26489);
nand U26860 (N_26860,N_26585,N_26571);
or U26861 (N_26861,N_26439,N_26476);
nor U26862 (N_26862,N_26421,N_26627);
nand U26863 (N_26863,N_26403,N_26452);
nand U26864 (N_26864,N_26585,N_26472);
nor U26865 (N_26865,N_26631,N_26411);
or U26866 (N_26866,N_26499,N_26579);
nor U26867 (N_26867,N_26577,N_26609);
nand U26868 (N_26868,N_26443,N_26473);
nand U26869 (N_26869,N_26501,N_26634);
and U26870 (N_26870,N_26495,N_26414);
nor U26871 (N_26871,N_26645,N_26533);
xor U26872 (N_26872,N_26446,N_26573);
or U26873 (N_26873,N_26676,N_26541);
or U26874 (N_26874,N_26456,N_26431);
or U26875 (N_26875,N_26510,N_26622);
and U26876 (N_26876,N_26640,N_26473);
or U26877 (N_26877,N_26412,N_26434);
or U26878 (N_26878,N_26688,N_26680);
xnor U26879 (N_26879,N_26605,N_26459);
xor U26880 (N_26880,N_26575,N_26687);
and U26881 (N_26881,N_26660,N_26487);
and U26882 (N_26882,N_26632,N_26505);
and U26883 (N_26883,N_26484,N_26538);
and U26884 (N_26884,N_26507,N_26654);
xor U26885 (N_26885,N_26641,N_26449);
nor U26886 (N_26886,N_26499,N_26668);
and U26887 (N_26887,N_26566,N_26673);
xnor U26888 (N_26888,N_26468,N_26607);
nand U26889 (N_26889,N_26626,N_26614);
xor U26890 (N_26890,N_26594,N_26507);
nand U26891 (N_26891,N_26557,N_26618);
nand U26892 (N_26892,N_26537,N_26507);
xnor U26893 (N_26893,N_26493,N_26569);
and U26894 (N_26894,N_26404,N_26640);
and U26895 (N_26895,N_26504,N_26578);
nand U26896 (N_26896,N_26545,N_26676);
or U26897 (N_26897,N_26417,N_26629);
or U26898 (N_26898,N_26548,N_26441);
xnor U26899 (N_26899,N_26611,N_26488);
nand U26900 (N_26900,N_26590,N_26610);
nor U26901 (N_26901,N_26553,N_26412);
nand U26902 (N_26902,N_26625,N_26448);
or U26903 (N_26903,N_26662,N_26614);
nand U26904 (N_26904,N_26530,N_26568);
nand U26905 (N_26905,N_26686,N_26541);
and U26906 (N_26906,N_26618,N_26406);
and U26907 (N_26907,N_26677,N_26624);
or U26908 (N_26908,N_26604,N_26476);
nand U26909 (N_26909,N_26562,N_26421);
xor U26910 (N_26910,N_26698,N_26622);
and U26911 (N_26911,N_26687,N_26689);
and U26912 (N_26912,N_26474,N_26648);
and U26913 (N_26913,N_26617,N_26461);
and U26914 (N_26914,N_26545,N_26604);
or U26915 (N_26915,N_26423,N_26571);
nand U26916 (N_26916,N_26476,N_26665);
or U26917 (N_26917,N_26534,N_26619);
and U26918 (N_26918,N_26433,N_26669);
xor U26919 (N_26919,N_26457,N_26608);
nand U26920 (N_26920,N_26620,N_26664);
xor U26921 (N_26921,N_26611,N_26420);
xor U26922 (N_26922,N_26685,N_26694);
xnor U26923 (N_26923,N_26690,N_26600);
nand U26924 (N_26924,N_26567,N_26428);
and U26925 (N_26925,N_26668,N_26437);
or U26926 (N_26926,N_26434,N_26622);
and U26927 (N_26927,N_26660,N_26500);
nand U26928 (N_26928,N_26656,N_26484);
nor U26929 (N_26929,N_26603,N_26610);
and U26930 (N_26930,N_26669,N_26513);
or U26931 (N_26931,N_26481,N_26456);
nor U26932 (N_26932,N_26604,N_26456);
or U26933 (N_26933,N_26445,N_26566);
and U26934 (N_26934,N_26621,N_26480);
or U26935 (N_26935,N_26656,N_26618);
or U26936 (N_26936,N_26545,N_26474);
nand U26937 (N_26937,N_26670,N_26582);
and U26938 (N_26938,N_26520,N_26586);
nor U26939 (N_26939,N_26532,N_26454);
and U26940 (N_26940,N_26467,N_26625);
nor U26941 (N_26941,N_26497,N_26649);
nand U26942 (N_26942,N_26432,N_26522);
and U26943 (N_26943,N_26696,N_26595);
xor U26944 (N_26944,N_26579,N_26633);
and U26945 (N_26945,N_26666,N_26504);
or U26946 (N_26946,N_26567,N_26628);
nor U26947 (N_26947,N_26408,N_26644);
nand U26948 (N_26948,N_26623,N_26497);
nor U26949 (N_26949,N_26481,N_26414);
nand U26950 (N_26950,N_26560,N_26588);
xor U26951 (N_26951,N_26580,N_26412);
or U26952 (N_26952,N_26542,N_26681);
and U26953 (N_26953,N_26499,N_26575);
nor U26954 (N_26954,N_26582,N_26654);
nand U26955 (N_26955,N_26422,N_26505);
or U26956 (N_26956,N_26544,N_26567);
and U26957 (N_26957,N_26495,N_26482);
nand U26958 (N_26958,N_26471,N_26600);
and U26959 (N_26959,N_26537,N_26573);
xnor U26960 (N_26960,N_26416,N_26593);
and U26961 (N_26961,N_26433,N_26656);
nand U26962 (N_26962,N_26540,N_26400);
and U26963 (N_26963,N_26529,N_26508);
nor U26964 (N_26964,N_26412,N_26693);
and U26965 (N_26965,N_26628,N_26493);
xor U26966 (N_26966,N_26696,N_26665);
nor U26967 (N_26967,N_26688,N_26460);
or U26968 (N_26968,N_26581,N_26435);
nand U26969 (N_26969,N_26460,N_26683);
xnor U26970 (N_26970,N_26454,N_26486);
xnor U26971 (N_26971,N_26553,N_26614);
xor U26972 (N_26972,N_26478,N_26437);
nand U26973 (N_26973,N_26480,N_26655);
nor U26974 (N_26974,N_26531,N_26593);
nor U26975 (N_26975,N_26478,N_26567);
nand U26976 (N_26976,N_26549,N_26403);
and U26977 (N_26977,N_26647,N_26464);
nand U26978 (N_26978,N_26559,N_26596);
xnor U26979 (N_26979,N_26430,N_26460);
or U26980 (N_26980,N_26423,N_26400);
xor U26981 (N_26981,N_26477,N_26438);
xor U26982 (N_26982,N_26516,N_26690);
nand U26983 (N_26983,N_26590,N_26693);
and U26984 (N_26984,N_26432,N_26500);
nor U26985 (N_26985,N_26621,N_26517);
or U26986 (N_26986,N_26585,N_26648);
and U26987 (N_26987,N_26655,N_26592);
and U26988 (N_26988,N_26640,N_26665);
or U26989 (N_26989,N_26423,N_26653);
nor U26990 (N_26990,N_26566,N_26525);
nor U26991 (N_26991,N_26533,N_26419);
nand U26992 (N_26992,N_26578,N_26416);
or U26993 (N_26993,N_26600,N_26552);
nor U26994 (N_26994,N_26462,N_26519);
and U26995 (N_26995,N_26596,N_26422);
or U26996 (N_26996,N_26548,N_26426);
or U26997 (N_26997,N_26694,N_26661);
nor U26998 (N_26998,N_26633,N_26697);
xnor U26999 (N_26999,N_26686,N_26414);
xnor U27000 (N_27000,N_26982,N_26950);
xnor U27001 (N_27001,N_26803,N_26776);
nand U27002 (N_27002,N_26866,N_26985);
and U27003 (N_27003,N_26967,N_26744);
or U27004 (N_27004,N_26879,N_26863);
and U27005 (N_27005,N_26867,N_26761);
and U27006 (N_27006,N_26873,N_26981);
nor U27007 (N_27007,N_26984,N_26928);
and U27008 (N_27008,N_26811,N_26785);
nand U27009 (N_27009,N_26860,N_26816);
or U27010 (N_27010,N_26908,N_26876);
or U27011 (N_27011,N_26815,N_26812);
or U27012 (N_27012,N_26729,N_26880);
nand U27013 (N_27013,N_26992,N_26912);
nand U27014 (N_27014,N_26813,N_26870);
and U27015 (N_27015,N_26706,N_26920);
nor U27016 (N_27016,N_26721,N_26995);
and U27017 (N_27017,N_26947,N_26893);
or U27018 (N_27018,N_26805,N_26888);
xnor U27019 (N_27019,N_26709,N_26939);
nand U27020 (N_27020,N_26759,N_26956);
nand U27021 (N_27021,N_26892,N_26977);
xnor U27022 (N_27022,N_26733,N_26951);
or U27023 (N_27023,N_26802,N_26821);
and U27024 (N_27024,N_26897,N_26868);
nor U27025 (N_27025,N_26792,N_26970);
and U27026 (N_27026,N_26701,N_26903);
and U27027 (N_27027,N_26788,N_26865);
and U27028 (N_27028,N_26851,N_26944);
nand U27029 (N_27029,N_26946,N_26971);
nand U27030 (N_27030,N_26760,N_26753);
xor U27031 (N_27031,N_26796,N_26878);
nor U27032 (N_27032,N_26906,N_26714);
and U27033 (N_27033,N_26864,N_26924);
and U27034 (N_27034,N_26933,N_26961);
xnor U27035 (N_27035,N_26728,N_26810);
nand U27036 (N_27036,N_26964,N_26949);
nand U27037 (N_27037,N_26926,N_26998);
or U27038 (N_27038,N_26828,N_26787);
nor U27039 (N_27039,N_26820,N_26835);
nor U27040 (N_27040,N_26739,N_26809);
nand U27041 (N_27041,N_26777,N_26840);
nor U27042 (N_27042,N_26837,N_26713);
and U27043 (N_27043,N_26881,N_26754);
and U27044 (N_27044,N_26742,N_26883);
xor U27045 (N_27045,N_26929,N_26937);
or U27046 (N_27046,N_26849,N_26855);
and U27047 (N_27047,N_26751,N_26853);
nor U27048 (N_27048,N_26889,N_26814);
xnor U27049 (N_27049,N_26996,N_26836);
xnor U27050 (N_27050,N_26755,N_26703);
and U27051 (N_27051,N_26765,N_26915);
xor U27052 (N_27052,N_26769,N_26871);
nand U27053 (N_27053,N_26720,N_26972);
and U27054 (N_27054,N_26983,N_26907);
and U27055 (N_27055,N_26936,N_26749);
nand U27056 (N_27056,N_26752,N_26758);
xor U27057 (N_27057,N_26965,N_26843);
and U27058 (N_27058,N_26770,N_26825);
or U27059 (N_27059,N_26778,N_26979);
and U27060 (N_27060,N_26819,N_26700);
xnor U27061 (N_27061,N_26799,N_26790);
or U27062 (N_27062,N_26845,N_26917);
or U27063 (N_27063,N_26774,N_26757);
nand U27064 (N_27064,N_26842,N_26885);
nand U27065 (N_27065,N_26856,N_26955);
xor U27066 (N_27066,N_26978,N_26730);
and U27067 (N_27067,N_26801,N_26782);
xor U27068 (N_27068,N_26705,N_26891);
nor U27069 (N_27069,N_26962,N_26794);
nand U27070 (N_27070,N_26895,N_26850);
and U27071 (N_27071,N_26740,N_26857);
or U27072 (N_27072,N_26875,N_26807);
nor U27073 (N_27073,N_26966,N_26838);
nand U27074 (N_27074,N_26741,N_26734);
and U27075 (N_27075,N_26991,N_26953);
or U27076 (N_27076,N_26986,N_26909);
nor U27077 (N_27077,N_26710,N_26771);
or U27078 (N_27078,N_26723,N_26960);
or U27079 (N_27079,N_26932,N_26724);
and U27080 (N_27080,N_26922,N_26874);
or U27081 (N_27081,N_26702,N_26784);
and U27082 (N_27082,N_26763,N_26822);
and U27083 (N_27083,N_26725,N_26957);
xnor U27084 (N_27084,N_26904,N_26877);
xnor U27085 (N_27085,N_26898,N_26779);
and U27086 (N_27086,N_26923,N_26743);
and U27087 (N_27087,N_26884,N_26795);
and U27088 (N_27088,N_26839,N_26767);
xor U27089 (N_27089,N_26841,N_26941);
or U27090 (N_27090,N_26833,N_26737);
nor U27091 (N_27091,N_26783,N_26712);
or U27092 (N_27092,N_26791,N_26797);
and U27093 (N_27093,N_26886,N_26900);
and U27094 (N_27094,N_26817,N_26975);
nor U27095 (N_27095,N_26804,N_26832);
xor U27096 (N_27096,N_26704,N_26948);
xor U27097 (N_27097,N_26727,N_26818);
and U27098 (N_27098,N_26859,N_26894);
nand U27099 (N_27099,N_26773,N_26719);
or U27100 (N_27100,N_26764,N_26890);
nor U27101 (N_27101,N_26934,N_26973);
nand U27102 (N_27102,N_26808,N_26916);
nand U27103 (N_27103,N_26980,N_26945);
nor U27104 (N_27104,N_26862,N_26738);
or U27105 (N_27105,N_26899,N_26942);
and U27106 (N_27106,N_26954,N_26988);
and U27107 (N_27107,N_26748,N_26823);
nand U27108 (N_27108,N_26935,N_26708);
and U27109 (N_27109,N_26715,N_26827);
nor U27110 (N_27110,N_26902,N_26974);
xor U27111 (N_27111,N_26989,N_26969);
xnor U27112 (N_27112,N_26913,N_26968);
nand U27113 (N_27113,N_26768,N_26736);
or U27114 (N_27114,N_26844,N_26976);
xor U27115 (N_27115,N_26716,N_26952);
xnor U27116 (N_27116,N_26958,N_26829);
and U27117 (N_27117,N_26756,N_26789);
nor U27118 (N_27118,N_26896,N_26830);
or U27119 (N_27119,N_26780,N_26993);
nor U27120 (N_27120,N_26766,N_26718);
nor U27121 (N_27121,N_26762,N_26750);
xor U27122 (N_27122,N_26834,N_26858);
or U27123 (N_27123,N_26793,N_26806);
or U27124 (N_27124,N_26918,N_26861);
xnor U27125 (N_27125,N_26943,N_26938);
nor U27126 (N_27126,N_26745,N_26911);
nand U27127 (N_27127,N_26910,N_26775);
and U27128 (N_27128,N_26746,N_26786);
and U27129 (N_27129,N_26987,N_26997);
nor U27130 (N_27130,N_26824,N_26990);
or U27131 (N_27131,N_26914,N_26999);
nand U27132 (N_27132,N_26994,N_26959);
xor U27133 (N_27133,N_26732,N_26930);
xor U27134 (N_27134,N_26717,N_26722);
xor U27135 (N_27135,N_26921,N_26905);
nor U27136 (N_27136,N_26831,N_26772);
xnor U27137 (N_27137,N_26852,N_26848);
xnor U27138 (N_27138,N_26872,N_26731);
xor U27139 (N_27139,N_26846,N_26826);
and U27140 (N_27140,N_26927,N_26798);
or U27141 (N_27141,N_26931,N_26887);
or U27142 (N_27142,N_26882,N_26747);
and U27143 (N_27143,N_26707,N_26963);
or U27144 (N_27144,N_26781,N_26901);
nand U27145 (N_27145,N_26726,N_26800);
or U27146 (N_27146,N_26869,N_26711);
nand U27147 (N_27147,N_26925,N_26854);
or U27148 (N_27148,N_26940,N_26847);
xor U27149 (N_27149,N_26919,N_26735);
and U27150 (N_27150,N_26952,N_26874);
nand U27151 (N_27151,N_26708,N_26712);
nand U27152 (N_27152,N_26774,N_26816);
nor U27153 (N_27153,N_26982,N_26906);
or U27154 (N_27154,N_26902,N_26883);
xor U27155 (N_27155,N_26731,N_26984);
xnor U27156 (N_27156,N_26822,N_26736);
xor U27157 (N_27157,N_26827,N_26999);
and U27158 (N_27158,N_26718,N_26762);
and U27159 (N_27159,N_26836,N_26949);
nor U27160 (N_27160,N_26721,N_26792);
or U27161 (N_27161,N_26741,N_26751);
xnor U27162 (N_27162,N_26844,N_26840);
nand U27163 (N_27163,N_26875,N_26730);
nand U27164 (N_27164,N_26933,N_26700);
nand U27165 (N_27165,N_26803,N_26845);
nor U27166 (N_27166,N_26764,N_26729);
nand U27167 (N_27167,N_26917,N_26770);
and U27168 (N_27168,N_26873,N_26979);
nor U27169 (N_27169,N_26809,N_26892);
xor U27170 (N_27170,N_26913,N_26856);
nand U27171 (N_27171,N_26805,N_26718);
nor U27172 (N_27172,N_26864,N_26795);
or U27173 (N_27173,N_26972,N_26789);
nand U27174 (N_27174,N_26727,N_26993);
nand U27175 (N_27175,N_26823,N_26930);
and U27176 (N_27176,N_26886,N_26948);
or U27177 (N_27177,N_26844,N_26796);
and U27178 (N_27178,N_26841,N_26902);
or U27179 (N_27179,N_26713,N_26992);
nor U27180 (N_27180,N_26972,N_26723);
xor U27181 (N_27181,N_26958,N_26782);
and U27182 (N_27182,N_26804,N_26838);
nand U27183 (N_27183,N_26965,N_26835);
nand U27184 (N_27184,N_26953,N_26773);
or U27185 (N_27185,N_26937,N_26909);
nor U27186 (N_27186,N_26706,N_26887);
nor U27187 (N_27187,N_26929,N_26738);
nor U27188 (N_27188,N_26825,N_26798);
xor U27189 (N_27189,N_26952,N_26956);
and U27190 (N_27190,N_26703,N_26807);
nor U27191 (N_27191,N_26955,N_26792);
nand U27192 (N_27192,N_26897,N_26822);
xor U27193 (N_27193,N_26896,N_26876);
xor U27194 (N_27194,N_26820,N_26923);
or U27195 (N_27195,N_26973,N_26935);
nor U27196 (N_27196,N_26940,N_26704);
nand U27197 (N_27197,N_26794,N_26835);
nor U27198 (N_27198,N_26942,N_26975);
and U27199 (N_27199,N_26932,N_26731);
nor U27200 (N_27200,N_26976,N_26761);
and U27201 (N_27201,N_26818,N_26906);
nor U27202 (N_27202,N_26998,N_26806);
nor U27203 (N_27203,N_26998,N_26700);
nand U27204 (N_27204,N_26861,N_26930);
nand U27205 (N_27205,N_26754,N_26845);
nor U27206 (N_27206,N_26704,N_26789);
nor U27207 (N_27207,N_26790,N_26810);
and U27208 (N_27208,N_26846,N_26831);
or U27209 (N_27209,N_26937,N_26891);
nand U27210 (N_27210,N_26796,N_26830);
nor U27211 (N_27211,N_26970,N_26921);
nor U27212 (N_27212,N_26929,N_26717);
and U27213 (N_27213,N_26902,N_26748);
and U27214 (N_27214,N_26926,N_26720);
and U27215 (N_27215,N_26869,N_26707);
nand U27216 (N_27216,N_26885,N_26875);
and U27217 (N_27217,N_26911,N_26849);
or U27218 (N_27218,N_26740,N_26725);
or U27219 (N_27219,N_26832,N_26876);
nor U27220 (N_27220,N_26762,N_26961);
or U27221 (N_27221,N_26763,N_26988);
nor U27222 (N_27222,N_26889,N_26952);
nand U27223 (N_27223,N_26867,N_26721);
nand U27224 (N_27224,N_26907,N_26707);
nor U27225 (N_27225,N_26910,N_26889);
and U27226 (N_27226,N_26913,N_26898);
nand U27227 (N_27227,N_26950,N_26705);
nand U27228 (N_27228,N_26951,N_26742);
nand U27229 (N_27229,N_26777,N_26778);
and U27230 (N_27230,N_26969,N_26735);
nand U27231 (N_27231,N_26774,N_26983);
and U27232 (N_27232,N_26894,N_26941);
xnor U27233 (N_27233,N_26926,N_26710);
and U27234 (N_27234,N_26919,N_26803);
nor U27235 (N_27235,N_26969,N_26997);
nand U27236 (N_27236,N_26795,N_26799);
nand U27237 (N_27237,N_26826,N_26868);
or U27238 (N_27238,N_26757,N_26822);
nor U27239 (N_27239,N_26791,N_26865);
nor U27240 (N_27240,N_26786,N_26815);
nand U27241 (N_27241,N_26802,N_26763);
or U27242 (N_27242,N_26897,N_26824);
nand U27243 (N_27243,N_26789,N_26952);
xnor U27244 (N_27244,N_26799,N_26824);
and U27245 (N_27245,N_26972,N_26874);
nand U27246 (N_27246,N_26905,N_26950);
and U27247 (N_27247,N_26976,N_26848);
and U27248 (N_27248,N_26989,N_26965);
or U27249 (N_27249,N_26820,N_26847);
nor U27250 (N_27250,N_26935,N_26938);
nand U27251 (N_27251,N_26800,N_26803);
nor U27252 (N_27252,N_26885,N_26715);
nand U27253 (N_27253,N_26854,N_26812);
and U27254 (N_27254,N_26765,N_26970);
or U27255 (N_27255,N_26966,N_26979);
xnor U27256 (N_27256,N_26811,N_26934);
and U27257 (N_27257,N_26912,N_26713);
and U27258 (N_27258,N_26757,N_26829);
nor U27259 (N_27259,N_26950,N_26765);
or U27260 (N_27260,N_26897,N_26950);
xnor U27261 (N_27261,N_26766,N_26933);
and U27262 (N_27262,N_26702,N_26851);
xor U27263 (N_27263,N_26730,N_26745);
xnor U27264 (N_27264,N_26884,N_26933);
xor U27265 (N_27265,N_26944,N_26755);
and U27266 (N_27266,N_26957,N_26907);
or U27267 (N_27267,N_26788,N_26767);
nand U27268 (N_27268,N_26968,N_26904);
and U27269 (N_27269,N_26766,N_26832);
xnor U27270 (N_27270,N_26831,N_26836);
nand U27271 (N_27271,N_26936,N_26917);
nor U27272 (N_27272,N_26709,N_26974);
and U27273 (N_27273,N_26984,N_26911);
or U27274 (N_27274,N_26877,N_26829);
xnor U27275 (N_27275,N_26957,N_26852);
nor U27276 (N_27276,N_26887,N_26777);
and U27277 (N_27277,N_26772,N_26996);
or U27278 (N_27278,N_26987,N_26713);
or U27279 (N_27279,N_26809,N_26843);
xor U27280 (N_27280,N_26843,N_26850);
nor U27281 (N_27281,N_26822,N_26787);
nor U27282 (N_27282,N_26757,N_26990);
nor U27283 (N_27283,N_26812,N_26772);
xor U27284 (N_27284,N_26801,N_26910);
nand U27285 (N_27285,N_26732,N_26847);
nor U27286 (N_27286,N_26788,N_26876);
xnor U27287 (N_27287,N_26755,N_26810);
nand U27288 (N_27288,N_26909,N_26762);
nand U27289 (N_27289,N_26931,N_26705);
or U27290 (N_27290,N_26950,N_26923);
nand U27291 (N_27291,N_26700,N_26747);
xor U27292 (N_27292,N_26813,N_26773);
nor U27293 (N_27293,N_26894,N_26851);
nand U27294 (N_27294,N_26864,N_26810);
nand U27295 (N_27295,N_26945,N_26851);
xor U27296 (N_27296,N_26997,N_26756);
xor U27297 (N_27297,N_26809,N_26975);
and U27298 (N_27298,N_26716,N_26987);
or U27299 (N_27299,N_26763,N_26837);
nor U27300 (N_27300,N_27117,N_27190);
or U27301 (N_27301,N_27209,N_27281);
nor U27302 (N_27302,N_27175,N_27155);
nand U27303 (N_27303,N_27044,N_27023);
or U27304 (N_27304,N_27121,N_27021);
nand U27305 (N_27305,N_27148,N_27173);
nor U27306 (N_27306,N_27098,N_27197);
nor U27307 (N_27307,N_27139,N_27081);
and U27308 (N_27308,N_27001,N_27291);
and U27309 (N_27309,N_27034,N_27004);
nand U27310 (N_27310,N_27168,N_27091);
and U27311 (N_27311,N_27035,N_27261);
nor U27312 (N_27312,N_27079,N_27217);
nor U27313 (N_27313,N_27104,N_27052);
nand U27314 (N_27314,N_27051,N_27258);
nand U27315 (N_27315,N_27270,N_27083);
nand U27316 (N_27316,N_27245,N_27212);
nor U27317 (N_27317,N_27187,N_27074);
and U27318 (N_27318,N_27229,N_27237);
xnor U27319 (N_27319,N_27076,N_27150);
nand U27320 (N_27320,N_27191,N_27196);
nor U27321 (N_27321,N_27038,N_27231);
or U27322 (N_27322,N_27131,N_27031);
nand U27323 (N_27323,N_27111,N_27140);
and U27324 (N_27324,N_27183,N_27216);
xor U27325 (N_27325,N_27165,N_27019);
nand U27326 (N_27326,N_27126,N_27127);
xnor U27327 (N_27327,N_27103,N_27100);
xnor U27328 (N_27328,N_27253,N_27124);
and U27329 (N_27329,N_27230,N_27105);
nand U27330 (N_27330,N_27101,N_27295);
xor U27331 (N_27331,N_27028,N_27233);
and U27332 (N_27332,N_27288,N_27254);
xnor U27333 (N_27333,N_27228,N_27055);
nand U27334 (N_27334,N_27181,N_27161);
nor U27335 (N_27335,N_27003,N_27041);
and U27336 (N_27336,N_27136,N_27205);
nor U27337 (N_27337,N_27266,N_27267);
or U27338 (N_27338,N_27172,N_27210);
and U27339 (N_27339,N_27075,N_27241);
xor U27340 (N_27340,N_27146,N_27211);
nor U27341 (N_27341,N_27201,N_27296);
nand U27342 (N_27342,N_27032,N_27027);
nand U27343 (N_27343,N_27043,N_27089);
or U27344 (N_27344,N_27192,N_27221);
and U27345 (N_27345,N_27108,N_27005);
and U27346 (N_27346,N_27132,N_27222);
and U27347 (N_27347,N_27282,N_27274);
or U27348 (N_27348,N_27122,N_27269);
xor U27349 (N_27349,N_27252,N_27234);
or U27350 (N_27350,N_27257,N_27073);
nor U27351 (N_27351,N_27134,N_27153);
nand U27352 (N_27352,N_27239,N_27145);
xnor U27353 (N_27353,N_27260,N_27141);
nor U27354 (N_27354,N_27066,N_27092);
and U27355 (N_27355,N_27093,N_27188);
nand U27356 (N_27356,N_27208,N_27119);
xnor U27357 (N_27357,N_27294,N_27162);
nand U27358 (N_27358,N_27120,N_27290);
or U27359 (N_27359,N_27219,N_27200);
or U27360 (N_27360,N_27275,N_27289);
nand U27361 (N_27361,N_27128,N_27184);
and U27362 (N_27362,N_27068,N_27144);
and U27363 (N_27363,N_27138,N_27226);
and U27364 (N_27364,N_27297,N_27242);
or U27365 (N_27365,N_27036,N_27225);
xnor U27366 (N_27366,N_27143,N_27096);
nor U27367 (N_27367,N_27263,N_27203);
xnor U27368 (N_27368,N_27223,N_27248);
nand U27369 (N_27369,N_27236,N_27195);
nor U27370 (N_27370,N_27189,N_27247);
nor U27371 (N_27371,N_27159,N_27174);
or U27372 (N_27372,N_27067,N_27064);
nand U27373 (N_27373,N_27244,N_27037);
or U27374 (N_27374,N_27271,N_27009);
nand U27375 (N_27375,N_27106,N_27265);
xnor U27376 (N_27376,N_27220,N_27026);
nor U27377 (N_27377,N_27118,N_27163);
xnor U27378 (N_27378,N_27042,N_27099);
xor U27379 (N_27379,N_27206,N_27243);
and U27380 (N_27380,N_27298,N_27273);
nand U27381 (N_27381,N_27213,N_27277);
nor U27382 (N_27382,N_27177,N_27025);
xnor U27383 (N_27383,N_27062,N_27010);
xor U27384 (N_27384,N_27072,N_27137);
nand U27385 (N_27385,N_27017,N_27285);
or U27386 (N_27386,N_27133,N_27193);
or U27387 (N_27387,N_27060,N_27279);
or U27388 (N_27388,N_27115,N_27116);
and U27389 (N_27389,N_27202,N_27147);
and U27390 (N_27390,N_27110,N_27059);
nand U27391 (N_27391,N_27088,N_27033);
nand U27392 (N_27392,N_27204,N_27130);
or U27393 (N_27393,N_27090,N_27286);
nand U27394 (N_27394,N_27158,N_27109);
nor U27395 (N_27395,N_27048,N_27050);
nor U27396 (N_27396,N_27082,N_27077);
xor U27397 (N_27397,N_27056,N_27224);
xnor U27398 (N_27398,N_27293,N_27284);
and U27399 (N_27399,N_27142,N_27250);
nand U27400 (N_27400,N_27084,N_27194);
nand U27401 (N_27401,N_27167,N_27039);
and U27402 (N_27402,N_27272,N_27246);
or U27403 (N_27403,N_27006,N_27014);
nor U27404 (N_27404,N_27264,N_27008);
nor U27405 (N_27405,N_27057,N_27151);
or U27406 (N_27406,N_27182,N_27232);
nand U27407 (N_27407,N_27287,N_27024);
or U27408 (N_27408,N_27094,N_27071);
or U27409 (N_27409,N_27125,N_27102);
nand U27410 (N_27410,N_27235,N_27179);
nor U27411 (N_27411,N_27012,N_27268);
xor U27412 (N_27412,N_27013,N_27070);
xor U27413 (N_27413,N_27018,N_27164);
or U27414 (N_27414,N_27097,N_27107);
xnor U27415 (N_27415,N_27240,N_27086);
or U27416 (N_27416,N_27123,N_27054);
xor U27417 (N_27417,N_27157,N_27283);
and U27418 (N_27418,N_27276,N_27218);
or U27419 (N_27419,N_27049,N_27149);
xnor U27420 (N_27420,N_27045,N_27040);
nand U27421 (N_27421,N_27238,N_27015);
nand U27422 (N_27422,N_27262,N_27095);
nor U27423 (N_27423,N_27047,N_27007);
xor U27424 (N_27424,N_27053,N_27061);
nand U27425 (N_27425,N_27135,N_27112);
nand U27426 (N_27426,N_27046,N_27251);
xnor U27427 (N_27427,N_27198,N_27186);
or U27428 (N_27428,N_27000,N_27080);
nor U27429 (N_27429,N_27215,N_27063);
nand U27430 (N_27430,N_27278,N_27259);
or U27431 (N_27431,N_27207,N_27171);
xnor U27432 (N_27432,N_27249,N_27002);
or U27433 (N_27433,N_27292,N_27280);
nor U27434 (N_27434,N_27020,N_27214);
nor U27435 (N_27435,N_27030,N_27227);
xor U27436 (N_27436,N_27058,N_27199);
nand U27437 (N_27437,N_27160,N_27170);
nor U27438 (N_27438,N_27129,N_27078);
and U27439 (N_27439,N_27299,N_27156);
xnor U27440 (N_27440,N_27166,N_27185);
xor U27441 (N_27441,N_27085,N_27152);
or U27442 (N_27442,N_27180,N_27029);
and U27443 (N_27443,N_27255,N_27169);
xor U27444 (N_27444,N_27176,N_27178);
and U27445 (N_27445,N_27069,N_27256);
and U27446 (N_27446,N_27087,N_27065);
xnor U27447 (N_27447,N_27016,N_27114);
or U27448 (N_27448,N_27022,N_27113);
nor U27449 (N_27449,N_27011,N_27154);
nand U27450 (N_27450,N_27247,N_27241);
nand U27451 (N_27451,N_27012,N_27093);
nor U27452 (N_27452,N_27105,N_27063);
xor U27453 (N_27453,N_27193,N_27136);
or U27454 (N_27454,N_27274,N_27132);
nor U27455 (N_27455,N_27064,N_27189);
xnor U27456 (N_27456,N_27247,N_27005);
or U27457 (N_27457,N_27173,N_27234);
nand U27458 (N_27458,N_27055,N_27285);
xor U27459 (N_27459,N_27127,N_27139);
nor U27460 (N_27460,N_27060,N_27280);
nor U27461 (N_27461,N_27216,N_27234);
xor U27462 (N_27462,N_27217,N_27150);
nand U27463 (N_27463,N_27298,N_27062);
or U27464 (N_27464,N_27108,N_27178);
nand U27465 (N_27465,N_27298,N_27068);
nor U27466 (N_27466,N_27043,N_27098);
xor U27467 (N_27467,N_27298,N_27104);
and U27468 (N_27468,N_27000,N_27082);
xor U27469 (N_27469,N_27147,N_27163);
xor U27470 (N_27470,N_27084,N_27224);
and U27471 (N_27471,N_27206,N_27083);
xor U27472 (N_27472,N_27187,N_27260);
nor U27473 (N_27473,N_27158,N_27011);
and U27474 (N_27474,N_27218,N_27072);
or U27475 (N_27475,N_27145,N_27129);
xnor U27476 (N_27476,N_27230,N_27126);
nor U27477 (N_27477,N_27182,N_27296);
or U27478 (N_27478,N_27285,N_27001);
or U27479 (N_27479,N_27154,N_27035);
and U27480 (N_27480,N_27097,N_27099);
or U27481 (N_27481,N_27172,N_27117);
or U27482 (N_27482,N_27086,N_27088);
xnor U27483 (N_27483,N_27022,N_27197);
nand U27484 (N_27484,N_27126,N_27152);
nand U27485 (N_27485,N_27168,N_27125);
and U27486 (N_27486,N_27288,N_27204);
xnor U27487 (N_27487,N_27027,N_27183);
xnor U27488 (N_27488,N_27120,N_27180);
xnor U27489 (N_27489,N_27240,N_27239);
xor U27490 (N_27490,N_27146,N_27244);
nand U27491 (N_27491,N_27265,N_27211);
nor U27492 (N_27492,N_27082,N_27241);
and U27493 (N_27493,N_27206,N_27099);
nor U27494 (N_27494,N_27149,N_27061);
xnor U27495 (N_27495,N_27096,N_27151);
xor U27496 (N_27496,N_27087,N_27246);
xnor U27497 (N_27497,N_27159,N_27135);
and U27498 (N_27498,N_27168,N_27161);
or U27499 (N_27499,N_27237,N_27128);
nand U27500 (N_27500,N_27078,N_27275);
xor U27501 (N_27501,N_27173,N_27124);
xor U27502 (N_27502,N_27294,N_27228);
and U27503 (N_27503,N_27023,N_27132);
and U27504 (N_27504,N_27070,N_27280);
and U27505 (N_27505,N_27270,N_27040);
xnor U27506 (N_27506,N_27025,N_27201);
and U27507 (N_27507,N_27037,N_27028);
and U27508 (N_27508,N_27068,N_27146);
or U27509 (N_27509,N_27209,N_27260);
nor U27510 (N_27510,N_27002,N_27276);
nand U27511 (N_27511,N_27137,N_27251);
and U27512 (N_27512,N_27211,N_27204);
nor U27513 (N_27513,N_27124,N_27294);
xnor U27514 (N_27514,N_27186,N_27008);
nand U27515 (N_27515,N_27009,N_27112);
nor U27516 (N_27516,N_27005,N_27241);
and U27517 (N_27517,N_27296,N_27172);
and U27518 (N_27518,N_27280,N_27263);
nand U27519 (N_27519,N_27115,N_27245);
nand U27520 (N_27520,N_27161,N_27005);
and U27521 (N_27521,N_27079,N_27245);
and U27522 (N_27522,N_27148,N_27021);
nor U27523 (N_27523,N_27254,N_27226);
nor U27524 (N_27524,N_27160,N_27181);
or U27525 (N_27525,N_27266,N_27015);
and U27526 (N_27526,N_27155,N_27052);
nand U27527 (N_27527,N_27148,N_27099);
xor U27528 (N_27528,N_27190,N_27049);
nand U27529 (N_27529,N_27021,N_27297);
or U27530 (N_27530,N_27202,N_27022);
xor U27531 (N_27531,N_27049,N_27053);
or U27532 (N_27532,N_27218,N_27121);
nor U27533 (N_27533,N_27053,N_27086);
xor U27534 (N_27534,N_27165,N_27174);
xnor U27535 (N_27535,N_27264,N_27131);
and U27536 (N_27536,N_27047,N_27108);
and U27537 (N_27537,N_27006,N_27260);
nand U27538 (N_27538,N_27212,N_27204);
and U27539 (N_27539,N_27245,N_27225);
xor U27540 (N_27540,N_27201,N_27262);
and U27541 (N_27541,N_27093,N_27111);
nor U27542 (N_27542,N_27275,N_27107);
nor U27543 (N_27543,N_27234,N_27126);
nand U27544 (N_27544,N_27238,N_27052);
and U27545 (N_27545,N_27128,N_27272);
or U27546 (N_27546,N_27279,N_27207);
xor U27547 (N_27547,N_27038,N_27102);
or U27548 (N_27548,N_27124,N_27073);
xor U27549 (N_27549,N_27131,N_27227);
or U27550 (N_27550,N_27155,N_27018);
and U27551 (N_27551,N_27085,N_27075);
nand U27552 (N_27552,N_27043,N_27239);
or U27553 (N_27553,N_27295,N_27181);
nand U27554 (N_27554,N_27157,N_27001);
xor U27555 (N_27555,N_27284,N_27198);
or U27556 (N_27556,N_27160,N_27297);
or U27557 (N_27557,N_27086,N_27280);
xnor U27558 (N_27558,N_27281,N_27126);
xnor U27559 (N_27559,N_27236,N_27011);
xor U27560 (N_27560,N_27124,N_27076);
and U27561 (N_27561,N_27237,N_27209);
nand U27562 (N_27562,N_27013,N_27218);
nor U27563 (N_27563,N_27106,N_27287);
nand U27564 (N_27564,N_27053,N_27042);
or U27565 (N_27565,N_27116,N_27142);
and U27566 (N_27566,N_27102,N_27219);
xnor U27567 (N_27567,N_27282,N_27261);
nand U27568 (N_27568,N_27183,N_27170);
nand U27569 (N_27569,N_27174,N_27028);
xor U27570 (N_27570,N_27260,N_27055);
nand U27571 (N_27571,N_27277,N_27051);
nand U27572 (N_27572,N_27063,N_27009);
nand U27573 (N_27573,N_27080,N_27289);
or U27574 (N_27574,N_27086,N_27248);
nor U27575 (N_27575,N_27223,N_27293);
and U27576 (N_27576,N_27078,N_27040);
nor U27577 (N_27577,N_27256,N_27117);
and U27578 (N_27578,N_27006,N_27167);
and U27579 (N_27579,N_27291,N_27048);
xor U27580 (N_27580,N_27242,N_27151);
nand U27581 (N_27581,N_27013,N_27280);
nand U27582 (N_27582,N_27105,N_27029);
nand U27583 (N_27583,N_27166,N_27075);
nor U27584 (N_27584,N_27243,N_27037);
or U27585 (N_27585,N_27009,N_27286);
nand U27586 (N_27586,N_27108,N_27250);
and U27587 (N_27587,N_27205,N_27144);
and U27588 (N_27588,N_27017,N_27137);
xnor U27589 (N_27589,N_27240,N_27210);
and U27590 (N_27590,N_27020,N_27114);
nand U27591 (N_27591,N_27110,N_27145);
or U27592 (N_27592,N_27265,N_27154);
nor U27593 (N_27593,N_27249,N_27055);
nand U27594 (N_27594,N_27060,N_27222);
and U27595 (N_27595,N_27272,N_27038);
nor U27596 (N_27596,N_27241,N_27266);
nor U27597 (N_27597,N_27245,N_27280);
xor U27598 (N_27598,N_27052,N_27245);
xnor U27599 (N_27599,N_27104,N_27087);
or U27600 (N_27600,N_27595,N_27574);
nor U27601 (N_27601,N_27458,N_27355);
nand U27602 (N_27602,N_27411,N_27393);
and U27603 (N_27603,N_27381,N_27456);
nor U27604 (N_27604,N_27489,N_27342);
xnor U27605 (N_27605,N_27597,N_27359);
or U27606 (N_27606,N_27545,N_27395);
nand U27607 (N_27607,N_27539,N_27562);
xnor U27608 (N_27608,N_27441,N_27544);
or U27609 (N_27609,N_27464,N_27498);
or U27610 (N_27610,N_27470,N_27341);
nor U27611 (N_27611,N_27483,N_27344);
xnor U27612 (N_27612,N_27491,N_27587);
or U27613 (N_27613,N_27334,N_27451);
and U27614 (N_27614,N_27372,N_27450);
nor U27615 (N_27615,N_27556,N_27519);
xnor U27616 (N_27616,N_27376,N_27570);
or U27617 (N_27617,N_27346,N_27347);
nand U27618 (N_27618,N_27404,N_27496);
xor U27619 (N_27619,N_27503,N_27412);
or U27620 (N_27620,N_27596,N_27466);
nor U27621 (N_27621,N_27516,N_27429);
or U27622 (N_27622,N_27399,N_27368);
xnor U27623 (N_27623,N_27312,N_27563);
or U27624 (N_27624,N_27364,N_27408);
and U27625 (N_27625,N_27308,N_27529);
xor U27626 (N_27626,N_27388,N_27313);
nor U27627 (N_27627,N_27481,N_27463);
and U27628 (N_27628,N_27379,N_27521);
xor U27629 (N_27629,N_27490,N_27448);
or U27630 (N_27630,N_27367,N_27509);
nand U27631 (N_27631,N_27378,N_27317);
and U27632 (N_27632,N_27440,N_27437);
nor U27633 (N_27633,N_27422,N_27484);
xnor U27634 (N_27634,N_27565,N_27338);
or U27635 (N_27635,N_27599,N_27373);
or U27636 (N_27636,N_27309,N_27366);
nand U27637 (N_27637,N_27428,N_27418);
xnor U27638 (N_27638,N_27377,N_27406);
and U27639 (N_27639,N_27535,N_27573);
nor U27640 (N_27640,N_27485,N_27306);
or U27641 (N_27641,N_27541,N_27527);
nand U27642 (N_27642,N_27575,N_27585);
xnor U27643 (N_27643,N_27319,N_27434);
and U27644 (N_27644,N_27542,N_27580);
or U27645 (N_27645,N_27560,N_27588);
nand U27646 (N_27646,N_27323,N_27325);
nand U27647 (N_27647,N_27537,N_27400);
and U27648 (N_27648,N_27505,N_27326);
nand U27649 (N_27649,N_27474,N_27543);
or U27650 (N_27650,N_27506,N_27592);
xor U27651 (N_27651,N_27522,N_27551);
or U27652 (N_27652,N_27518,N_27532);
nand U27653 (N_27653,N_27510,N_27419);
nor U27654 (N_27654,N_27436,N_27536);
and U27655 (N_27655,N_27321,N_27476);
xor U27656 (N_27656,N_27449,N_27569);
nor U27657 (N_27657,N_27486,N_27546);
nor U27658 (N_27658,N_27593,N_27357);
nor U27659 (N_27659,N_27337,N_27438);
and U27660 (N_27660,N_27443,N_27384);
and U27661 (N_27661,N_27305,N_27502);
or U27662 (N_27662,N_27479,N_27533);
nor U27663 (N_27663,N_27414,N_27314);
xnor U27664 (N_27664,N_27442,N_27307);
or U27665 (N_27665,N_27446,N_27421);
nand U27666 (N_27666,N_27591,N_27469);
or U27667 (N_27667,N_27584,N_27540);
and U27668 (N_27668,N_27457,N_27362);
and U27669 (N_27669,N_27329,N_27335);
or U27670 (N_27670,N_27324,N_27439);
or U27671 (N_27671,N_27396,N_27375);
nor U27672 (N_27672,N_27382,N_27514);
and U27673 (N_27673,N_27475,N_27526);
xor U27674 (N_27674,N_27467,N_27363);
nand U27675 (N_27675,N_27331,N_27311);
or U27676 (N_27676,N_27572,N_27413);
xor U27677 (N_27677,N_27425,N_27327);
and U27678 (N_27678,N_27390,N_27552);
and U27679 (N_27679,N_27555,N_27461);
and U27680 (N_27680,N_27497,N_27530);
nor U27681 (N_27681,N_27332,N_27517);
nor U27682 (N_27682,N_27568,N_27559);
xor U27683 (N_27683,N_27576,N_27330);
nand U27684 (N_27684,N_27548,N_27495);
xor U27685 (N_27685,N_27561,N_27493);
and U27686 (N_27686,N_27547,N_27459);
xor U27687 (N_27687,N_27424,N_27435);
and U27688 (N_27688,N_27369,N_27383);
or U27689 (N_27689,N_27358,N_27582);
nand U27690 (N_27690,N_27586,N_27564);
nor U27691 (N_27691,N_27432,N_27531);
nand U27692 (N_27692,N_27583,N_27389);
nor U27693 (N_27693,N_27310,N_27508);
and U27694 (N_27694,N_27480,N_27352);
or U27695 (N_27695,N_27447,N_27402);
xor U27696 (N_27696,N_27349,N_27303);
and U27697 (N_27697,N_27351,N_27453);
or U27698 (N_27698,N_27520,N_27523);
and U27699 (N_27699,N_27407,N_27482);
nand U27700 (N_27700,N_27524,N_27557);
or U27701 (N_27701,N_27566,N_27445);
and U27702 (N_27702,N_27405,N_27471);
and U27703 (N_27703,N_27410,N_27354);
nor U27704 (N_27704,N_27578,N_27525);
nor U27705 (N_27705,N_27423,N_27558);
nand U27706 (N_27706,N_27433,N_27374);
and U27707 (N_27707,N_27304,N_27473);
xnor U27708 (N_27708,N_27452,N_27488);
and U27709 (N_27709,N_27454,N_27507);
nand U27710 (N_27710,N_27460,N_27420);
nand U27711 (N_27711,N_27528,N_27513);
or U27712 (N_27712,N_27394,N_27538);
nand U27713 (N_27713,N_27511,N_27356);
or U27714 (N_27714,N_27567,N_27397);
and U27715 (N_27715,N_27579,N_27431);
xor U27716 (N_27716,N_27571,N_27426);
xnor U27717 (N_27717,N_27492,N_27343);
and U27718 (N_27718,N_27365,N_27468);
xor U27719 (N_27719,N_27302,N_27478);
or U27720 (N_27720,N_27398,N_27427);
nand U27721 (N_27721,N_27380,N_27415);
nand U27722 (N_27722,N_27328,N_27361);
xnor U27723 (N_27723,N_27577,N_27589);
nand U27724 (N_27724,N_27391,N_27340);
nor U27725 (N_27725,N_27392,N_27549);
xor U27726 (N_27726,N_27316,N_27360);
xor U27727 (N_27727,N_27386,N_27318);
nand U27728 (N_27728,N_27333,N_27345);
or U27729 (N_27729,N_27512,N_27430);
and U27730 (N_27730,N_27387,N_27515);
or U27731 (N_27731,N_27499,N_27500);
nor U27732 (N_27732,N_27320,N_27598);
and U27733 (N_27733,N_27487,N_27370);
and U27734 (N_27734,N_27336,N_27534);
nor U27735 (N_27735,N_27581,N_27300);
or U27736 (N_27736,N_27504,N_27371);
nand U27737 (N_27737,N_27554,N_27550);
and U27738 (N_27738,N_27350,N_27339);
nand U27739 (N_27739,N_27465,N_27444);
or U27740 (N_27740,N_27590,N_27462);
nand U27741 (N_27741,N_27416,N_27385);
nand U27742 (N_27742,N_27455,N_27353);
or U27743 (N_27743,N_27501,N_27348);
and U27744 (N_27744,N_27409,N_27494);
xnor U27745 (N_27745,N_27417,N_27403);
xnor U27746 (N_27746,N_27477,N_27315);
or U27747 (N_27747,N_27401,N_27594);
and U27748 (N_27748,N_27472,N_27553);
or U27749 (N_27749,N_27301,N_27322);
nand U27750 (N_27750,N_27562,N_27565);
nor U27751 (N_27751,N_27327,N_27340);
or U27752 (N_27752,N_27492,N_27524);
and U27753 (N_27753,N_27378,N_27475);
and U27754 (N_27754,N_27597,N_27322);
nor U27755 (N_27755,N_27421,N_27599);
nand U27756 (N_27756,N_27543,N_27512);
nand U27757 (N_27757,N_27535,N_27536);
nor U27758 (N_27758,N_27440,N_27373);
or U27759 (N_27759,N_27474,N_27596);
or U27760 (N_27760,N_27549,N_27490);
xor U27761 (N_27761,N_27483,N_27309);
nand U27762 (N_27762,N_27422,N_27456);
and U27763 (N_27763,N_27448,N_27572);
xor U27764 (N_27764,N_27328,N_27558);
nand U27765 (N_27765,N_27550,N_27577);
or U27766 (N_27766,N_27599,N_27556);
and U27767 (N_27767,N_27385,N_27375);
or U27768 (N_27768,N_27528,N_27300);
nand U27769 (N_27769,N_27571,N_27581);
xor U27770 (N_27770,N_27499,N_27543);
nand U27771 (N_27771,N_27595,N_27335);
xor U27772 (N_27772,N_27308,N_27474);
nor U27773 (N_27773,N_27433,N_27438);
and U27774 (N_27774,N_27523,N_27538);
nor U27775 (N_27775,N_27428,N_27381);
and U27776 (N_27776,N_27438,N_27589);
nor U27777 (N_27777,N_27597,N_27429);
xor U27778 (N_27778,N_27580,N_27328);
xor U27779 (N_27779,N_27483,N_27477);
or U27780 (N_27780,N_27354,N_27477);
xnor U27781 (N_27781,N_27378,N_27489);
nand U27782 (N_27782,N_27467,N_27416);
or U27783 (N_27783,N_27348,N_27505);
and U27784 (N_27784,N_27313,N_27554);
and U27785 (N_27785,N_27392,N_27505);
and U27786 (N_27786,N_27311,N_27598);
and U27787 (N_27787,N_27497,N_27448);
xor U27788 (N_27788,N_27515,N_27360);
or U27789 (N_27789,N_27406,N_27528);
nand U27790 (N_27790,N_27402,N_27446);
and U27791 (N_27791,N_27559,N_27507);
and U27792 (N_27792,N_27559,N_27476);
xor U27793 (N_27793,N_27461,N_27330);
or U27794 (N_27794,N_27455,N_27548);
xor U27795 (N_27795,N_27396,N_27513);
or U27796 (N_27796,N_27548,N_27572);
xnor U27797 (N_27797,N_27387,N_27444);
nor U27798 (N_27798,N_27596,N_27380);
nand U27799 (N_27799,N_27488,N_27454);
nand U27800 (N_27800,N_27550,N_27316);
and U27801 (N_27801,N_27304,N_27550);
or U27802 (N_27802,N_27459,N_27549);
nand U27803 (N_27803,N_27553,N_27456);
or U27804 (N_27804,N_27334,N_27327);
xnor U27805 (N_27805,N_27361,N_27515);
xnor U27806 (N_27806,N_27468,N_27406);
nor U27807 (N_27807,N_27425,N_27401);
nand U27808 (N_27808,N_27509,N_27429);
and U27809 (N_27809,N_27325,N_27381);
or U27810 (N_27810,N_27595,N_27494);
and U27811 (N_27811,N_27410,N_27595);
nand U27812 (N_27812,N_27364,N_27596);
nand U27813 (N_27813,N_27457,N_27494);
nand U27814 (N_27814,N_27527,N_27308);
xnor U27815 (N_27815,N_27314,N_27457);
xor U27816 (N_27816,N_27307,N_27304);
or U27817 (N_27817,N_27427,N_27471);
and U27818 (N_27818,N_27528,N_27353);
nor U27819 (N_27819,N_27319,N_27303);
nor U27820 (N_27820,N_27429,N_27373);
nor U27821 (N_27821,N_27369,N_27519);
nor U27822 (N_27822,N_27409,N_27568);
xnor U27823 (N_27823,N_27307,N_27511);
or U27824 (N_27824,N_27345,N_27464);
and U27825 (N_27825,N_27509,N_27506);
nand U27826 (N_27826,N_27476,N_27598);
nand U27827 (N_27827,N_27418,N_27575);
nor U27828 (N_27828,N_27551,N_27320);
nand U27829 (N_27829,N_27383,N_27555);
xnor U27830 (N_27830,N_27515,N_27444);
nor U27831 (N_27831,N_27548,N_27492);
xnor U27832 (N_27832,N_27561,N_27505);
and U27833 (N_27833,N_27544,N_27510);
nor U27834 (N_27834,N_27584,N_27482);
or U27835 (N_27835,N_27599,N_27310);
nand U27836 (N_27836,N_27440,N_27382);
and U27837 (N_27837,N_27341,N_27466);
and U27838 (N_27838,N_27544,N_27423);
xor U27839 (N_27839,N_27331,N_27560);
or U27840 (N_27840,N_27417,N_27352);
and U27841 (N_27841,N_27465,N_27373);
xnor U27842 (N_27842,N_27488,N_27564);
or U27843 (N_27843,N_27453,N_27568);
and U27844 (N_27844,N_27450,N_27383);
or U27845 (N_27845,N_27485,N_27478);
and U27846 (N_27846,N_27338,N_27355);
xnor U27847 (N_27847,N_27487,N_27572);
and U27848 (N_27848,N_27496,N_27507);
or U27849 (N_27849,N_27305,N_27556);
xnor U27850 (N_27850,N_27401,N_27330);
xor U27851 (N_27851,N_27398,N_27563);
and U27852 (N_27852,N_27512,N_27391);
or U27853 (N_27853,N_27339,N_27357);
nand U27854 (N_27854,N_27458,N_27336);
or U27855 (N_27855,N_27541,N_27581);
or U27856 (N_27856,N_27557,N_27528);
nand U27857 (N_27857,N_27587,N_27591);
nor U27858 (N_27858,N_27469,N_27401);
xor U27859 (N_27859,N_27420,N_27382);
nor U27860 (N_27860,N_27370,N_27396);
nor U27861 (N_27861,N_27530,N_27518);
or U27862 (N_27862,N_27356,N_27527);
xor U27863 (N_27863,N_27426,N_27435);
xor U27864 (N_27864,N_27517,N_27379);
nor U27865 (N_27865,N_27433,N_27462);
nand U27866 (N_27866,N_27494,N_27420);
nor U27867 (N_27867,N_27446,N_27339);
or U27868 (N_27868,N_27409,N_27439);
nor U27869 (N_27869,N_27542,N_27509);
xor U27870 (N_27870,N_27407,N_27516);
or U27871 (N_27871,N_27408,N_27469);
or U27872 (N_27872,N_27542,N_27388);
xnor U27873 (N_27873,N_27482,N_27378);
nor U27874 (N_27874,N_27409,N_27366);
xor U27875 (N_27875,N_27452,N_27341);
nor U27876 (N_27876,N_27454,N_27305);
and U27877 (N_27877,N_27515,N_27321);
xnor U27878 (N_27878,N_27557,N_27576);
nor U27879 (N_27879,N_27452,N_27499);
nand U27880 (N_27880,N_27370,N_27306);
xnor U27881 (N_27881,N_27551,N_27495);
and U27882 (N_27882,N_27589,N_27481);
and U27883 (N_27883,N_27510,N_27558);
xnor U27884 (N_27884,N_27422,N_27494);
xnor U27885 (N_27885,N_27595,N_27461);
and U27886 (N_27886,N_27482,N_27552);
and U27887 (N_27887,N_27433,N_27390);
nand U27888 (N_27888,N_27412,N_27381);
or U27889 (N_27889,N_27313,N_27318);
or U27890 (N_27890,N_27513,N_27442);
nand U27891 (N_27891,N_27450,N_27599);
nor U27892 (N_27892,N_27554,N_27460);
or U27893 (N_27893,N_27347,N_27369);
nor U27894 (N_27894,N_27583,N_27417);
nor U27895 (N_27895,N_27519,N_27500);
and U27896 (N_27896,N_27324,N_27369);
and U27897 (N_27897,N_27414,N_27407);
nor U27898 (N_27898,N_27471,N_27404);
and U27899 (N_27899,N_27430,N_27428);
nand U27900 (N_27900,N_27781,N_27748);
and U27901 (N_27901,N_27634,N_27726);
xnor U27902 (N_27902,N_27868,N_27707);
nor U27903 (N_27903,N_27725,N_27744);
nor U27904 (N_27904,N_27801,N_27700);
or U27905 (N_27905,N_27660,N_27706);
or U27906 (N_27906,N_27762,N_27639);
nand U27907 (N_27907,N_27765,N_27767);
xor U27908 (N_27908,N_27761,N_27784);
nand U27909 (N_27909,N_27740,N_27606);
xnor U27910 (N_27910,N_27642,N_27733);
xor U27911 (N_27911,N_27858,N_27617);
nor U27912 (N_27912,N_27800,N_27861);
xor U27913 (N_27913,N_27711,N_27742);
nand U27914 (N_27914,N_27717,N_27754);
and U27915 (N_27915,N_27689,N_27876);
or U27916 (N_27916,N_27723,N_27890);
or U27917 (N_27917,N_27720,N_27797);
xor U27918 (N_27918,N_27853,N_27758);
and U27919 (N_27919,N_27894,N_27613);
or U27920 (N_27920,N_27786,N_27691);
nor U27921 (N_27921,N_27722,N_27741);
nor U27922 (N_27922,N_27685,N_27701);
or U27923 (N_27923,N_27829,N_27844);
nand U27924 (N_27924,N_27698,N_27734);
or U27925 (N_27925,N_27863,N_27878);
or U27926 (N_27926,N_27806,N_27895);
or U27927 (N_27927,N_27777,N_27735);
and U27928 (N_27928,N_27747,N_27803);
xnor U27929 (N_27929,N_27884,N_27760);
or U27930 (N_27930,N_27752,N_27826);
nor U27931 (N_27931,N_27852,N_27798);
and U27932 (N_27932,N_27886,N_27757);
nand U27933 (N_27933,N_27819,N_27773);
and U27934 (N_27934,N_27710,N_27724);
nor U27935 (N_27935,N_27641,N_27833);
xor U27936 (N_27936,N_27825,N_27790);
and U27937 (N_27937,N_27662,N_27877);
nor U27938 (N_27938,N_27821,N_27843);
nand U27939 (N_27939,N_27675,N_27655);
or U27940 (N_27940,N_27831,N_27632);
nand U27941 (N_27941,N_27705,N_27793);
xor U27942 (N_27942,N_27645,N_27750);
nand U27943 (N_27943,N_27610,N_27630);
nand U27944 (N_27944,N_27648,N_27649);
and U27945 (N_27945,N_27620,N_27749);
nor U27946 (N_27946,N_27622,N_27719);
xnor U27947 (N_27947,N_27860,N_27653);
or U27948 (N_27948,N_27899,N_27772);
and U27949 (N_27949,N_27898,N_27888);
nor U27950 (N_27950,N_27796,N_27864);
nand U27951 (N_27951,N_27680,N_27881);
and U27952 (N_27952,N_27842,N_27817);
and U27953 (N_27953,N_27841,N_27702);
nand U27954 (N_27954,N_27669,N_27805);
nor U27955 (N_27955,N_27654,N_27812);
nor U27956 (N_27956,N_27769,N_27650);
xor U27957 (N_27957,N_27730,N_27775);
nor U27958 (N_27958,N_27739,N_27746);
nor U27959 (N_27959,N_27856,N_27820);
nor U27960 (N_27960,N_27712,N_27727);
and U27961 (N_27961,N_27670,N_27713);
and U27962 (N_27962,N_27804,N_27646);
or U27963 (N_27963,N_27729,N_27647);
or U27964 (N_27964,N_27847,N_27849);
xnor U27965 (N_27965,N_27755,N_27708);
nand U27966 (N_27966,N_27629,N_27663);
or U27967 (N_27967,N_27618,N_27794);
or U27968 (N_27968,N_27893,N_27605);
nand U27969 (N_27969,N_27880,N_27695);
and U27970 (N_27970,N_27840,N_27791);
and U27971 (N_27971,N_27751,N_27872);
nand U27972 (N_27972,N_27745,N_27783);
xnor U27973 (N_27973,N_27846,N_27731);
and U27974 (N_27974,N_27616,N_27871);
xnor U27975 (N_27975,N_27827,N_27756);
nor U27976 (N_27976,N_27736,N_27809);
xnor U27977 (N_27977,N_27792,N_27859);
or U27978 (N_27978,N_27602,N_27683);
nand U27979 (N_27979,N_27811,N_27866);
and U27980 (N_27980,N_27674,N_27694);
xor U27981 (N_27981,N_27766,N_27690);
nor U27982 (N_27982,N_27603,N_27870);
xor U27983 (N_27983,N_27838,N_27823);
nand U27984 (N_27984,N_27788,N_27665);
and U27985 (N_27985,N_27714,N_27633);
nor U27986 (N_27986,N_27728,N_27614);
nor U27987 (N_27987,N_27743,N_27658);
xnor U27988 (N_27988,N_27815,N_27640);
or U27989 (N_27989,N_27676,N_27779);
nand U27990 (N_27990,N_27636,N_27818);
nor U27991 (N_27991,N_27709,N_27774);
nor U27992 (N_27992,N_27810,N_27608);
nand U27993 (N_27993,N_27776,N_27737);
and U27994 (N_27994,N_27609,N_27628);
xnor U27995 (N_27995,N_27703,N_27855);
nand U27996 (N_27996,N_27611,N_27604);
nor U27997 (N_27997,N_27721,N_27850);
nand U27998 (N_27998,N_27824,N_27666);
nand U27999 (N_27999,N_27619,N_27873);
xnor U28000 (N_28000,N_27657,N_27780);
and U28001 (N_28001,N_27857,N_27867);
nor U28002 (N_28002,N_27621,N_27673);
xnor U28003 (N_28003,N_27626,N_27600);
xnor U28004 (N_28004,N_27768,N_27759);
and U28005 (N_28005,N_27764,N_27885);
nor U28006 (N_28006,N_27686,N_27692);
and U28007 (N_28007,N_27638,N_27787);
or U28008 (N_28008,N_27862,N_27715);
nor U28009 (N_28009,N_27808,N_27652);
nand U28010 (N_28010,N_27834,N_27896);
nor U28011 (N_28011,N_27822,N_27718);
xor U28012 (N_28012,N_27732,N_27643);
xor U28013 (N_28013,N_27882,N_27789);
nor U28014 (N_28014,N_27672,N_27854);
nor U28015 (N_28015,N_27631,N_27644);
nand U28016 (N_28016,N_27661,N_27839);
nand U28017 (N_28017,N_27869,N_27623);
xnor U28018 (N_28018,N_27697,N_27696);
nand U28019 (N_28019,N_27688,N_27659);
nor U28020 (N_28020,N_27699,N_27668);
xnor U28021 (N_28021,N_27671,N_27678);
or U28022 (N_28022,N_27874,N_27651);
nand U28023 (N_28023,N_27624,N_27627);
nor U28024 (N_28024,N_27716,N_27656);
and U28025 (N_28025,N_27795,N_27687);
or U28026 (N_28026,N_27770,N_27753);
or U28027 (N_28027,N_27848,N_27738);
or U28028 (N_28028,N_27704,N_27892);
nor U28029 (N_28029,N_27679,N_27681);
and U28030 (N_28030,N_27607,N_27667);
xnor U28031 (N_28031,N_27677,N_27865);
xnor U28032 (N_28032,N_27778,N_27830);
and U28033 (N_28033,N_27837,N_27799);
or U28034 (N_28034,N_27601,N_27832);
and U28035 (N_28035,N_27835,N_27814);
nor U28036 (N_28036,N_27771,N_27615);
xnor U28037 (N_28037,N_27883,N_27807);
xor U28038 (N_28038,N_27891,N_27875);
and U28039 (N_28039,N_27879,N_27637);
nor U28040 (N_28040,N_27802,N_27635);
nand U28041 (N_28041,N_27816,N_27612);
or U28042 (N_28042,N_27828,N_27813);
or U28043 (N_28043,N_27625,N_27682);
and U28044 (N_28044,N_27897,N_27845);
xor U28045 (N_28045,N_27763,N_27887);
or U28046 (N_28046,N_27889,N_27664);
and U28047 (N_28047,N_27851,N_27836);
nand U28048 (N_28048,N_27785,N_27693);
nor U28049 (N_28049,N_27684,N_27782);
or U28050 (N_28050,N_27856,N_27790);
nand U28051 (N_28051,N_27842,N_27611);
or U28052 (N_28052,N_27849,N_27738);
nand U28053 (N_28053,N_27691,N_27866);
nor U28054 (N_28054,N_27825,N_27742);
xnor U28055 (N_28055,N_27776,N_27801);
and U28056 (N_28056,N_27817,N_27888);
and U28057 (N_28057,N_27721,N_27695);
nand U28058 (N_28058,N_27732,N_27729);
nor U28059 (N_28059,N_27861,N_27688);
xnor U28060 (N_28060,N_27838,N_27844);
or U28061 (N_28061,N_27639,N_27858);
or U28062 (N_28062,N_27722,N_27827);
nand U28063 (N_28063,N_27613,N_27697);
or U28064 (N_28064,N_27710,N_27878);
and U28065 (N_28065,N_27602,N_27743);
and U28066 (N_28066,N_27759,N_27647);
nand U28067 (N_28067,N_27779,N_27885);
or U28068 (N_28068,N_27774,N_27691);
xnor U28069 (N_28069,N_27733,N_27819);
nand U28070 (N_28070,N_27691,N_27878);
nor U28071 (N_28071,N_27694,N_27871);
xnor U28072 (N_28072,N_27743,N_27799);
xnor U28073 (N_28073,N_27828,N_27838);
and U28074 (N_28074,N_27734,N_27813);
xor U28075 (N_28075,N_27800,N_27881);
and U28076 (N_28076,N_27647,N_27796);
nand U28077 (N_28077,N_27607,N_27896);
or U28078 (N_28078,N_27894,N_27624);
xnor U28079 (N_28079,N_27809,N_27782);
nand U28080 (N_28080,N_27802,N_27812);
xor U28081 (N_28081,N_27894,N_27707);
and U28082 (N_28082,N_27704,N_27793);
and U28083 (N_28083,N_27647,N_27665);
nor U28084 (N_28084,N_27621,N_27762);
or U28085 (N_28085,N_27746,N_27838);
nor U28086 (N_28086,N_27666,N_27720);
nor U28087 (N_28087,N_27861,N_27895);
and U28088 (N_28088,N_27656,N_27626);
nand U28089 (N_28089,N_27659,N_27714);
nand U28090 (N_28090,N_27708,N_27616);
and U28091 (N_28091,N_27713,N_27628);
and U28092 (N_28092,N_27611,N_27799);
and U28093 (N_28093,N_27775,N_27793);
nand U28094 (N_28094,N_27724,N_27842);
xor U28095 (N_28095,N_27603,N_27745);
xor U28096 (N_28096,N_27608,N_27839);
xor U28097 (N_28097,N_27852,N_27650);
nand U28098 (N_28098,N_27614,N_27814);
nand U28099 (N_28099,N_27673,N_27679);
nor U28100 (N_28100,N_27867,N_27750);
nand U28101 (N_28101,N_27638,N_27840);
or U28102 (N_28102,N_27857,N_27786);
or U28103 (N_28103,N_27808,N_27814);
or U28104 (N_28104,N_27773,N_27783);
xnor U28105 (N_28105,N_27840,N_27874);
nand U28106 (N_28106,N_27857,N_27889);
nand U28107 (N_28107,N_27879,N_27640);
nand U28108 (N_28108,N_27731,N_27627);
xor U28109 (N_28109,N_27708,N_27624);
nand U28110 (N_28110,N_27623,N_27619);
nand U28111 (N_28111,N_27779,N_27823);
and U28112 (N_28112,N_27682,N_27670);
xnor U28113 (N_28113,N_27801,N_27714);
xor U28114 (N_28114,N_27677,N_27815);
nor U28115 (N_28115,N_27635,N_27859);
nand U28116 (N_28116,N_27866,N_27627);
xor U28117 (N_28117,N_27740,N_27811);
or U28118 (N_28118,N_27652,N_27751);
nor U28119 (N_28119,N_27893,N_27850);
xor U28120 (N_28120,N_27622,N_27877);
and U28121 (N_28121,N_27612,N_27624);
and U28122 (N_28122,N_27767,N_27827);
and U28123 (N_28123,N_27782,N_27761);
or U28124 (N_28124,N_27808,N_27655);
xnor U28125 (N_28125,N_27659,N_27831);
nor U28126 (N_28126,N_27706,N_27866);
xnor U28127 (N_28127,N_27652,N_27641);
and U28128 (N_28128,N_27810,N_27627);
nor U28129 (N_28129,N_27610,N_27743);
nand U28130 (N_28130,N_27843,N_27769);
nor U28131 (N_28131,N_27668,N_27859);
nor U28132 (N_28132,N_27600,N_27855);
nor U28133 (N_28133,N_27693,N_27875);
nand U28134 (N_28134,N_27831,N_27607);
and U28135 (N_28135,N_27849,N_27778);
and U28136 (N_28136,N_27600,N_27644);
or U28137 (N_28137,N_27865,N_27681);
and U28138 (N_28138,N_27886,N_27859);
and U28139 (N_28139,N_27850,N_27761);
and U28140 (N_28140,N_27729,N_27814);
or U28141 (N_28141,N_27879,N_27794);
nand U28142 (N_28142,N_27742,N_27721);
nand U28143 (N_28143,N_27654,N_27731);
xor U28144 (N_28144,N_27824,N_27832);
xor U28145 (N_28145,N_27779,N_27867);
or U28146 (N_28146,N_27792,N_27894);
xnor U28147 (N_28147,N_27657,N_27726);
nand U28148 (N_28148,N_27859,N_27835);
or U28149 (N_28149,N_27749,N_27847);
and U28150 (N_28150,N_27748,N_27681);
xnor U28151 (N_28151,N_27759,N_27620);
nand U28152 (N_28152,N_27681,N_27676);
or U28153 (N_28153,N_27818,N_27637);
or U28154 (N_28154,N_27710,N_27708);
xnor U28155 (N_28155,N_27808,N_27888);
and U28156 (N_28156,N_27662,N_27690);
nor U28157 (N_28157,N_27672,N_27781);
nor U28158 (N_28158,N_27796,N_27851);
and U28159 (N_28159,N_27757,N_27804);
or U28160 (N_28160,N_27718,N_27849);
nand U28161 (N_28161,N_27753,N_27667);
nand U28162 (N_28162,N_27821,N_27715);
nor U28163 (N_28163,N_27817,N_27715);
nand U28164 (N_28164,N_27753,N_27804);
nor U28165 (N_28165,N_27873,N_27775);
xnor U28166 (N_28166,N_27729,N_27867);
and U28167 (N_28167,N_27872,N_27668);
xor U28168 (N_28168,N_27716,N_27897);
or U28169 (N_28169,N_27704,N_27801);
and U28170 (N_28170,N_27671,N_27690);
xor U28171 (N_28171,N_27757,N_27700);
xnor U28172 (N_28172,N_27796,N_27789);
nor U28173 (N_28173,N_27600,N_27610);
or U28174 (N_28174,N_27653,N_27606);
nor U28175 (N_28175,N_27778,N_27605);
nand U28176 (N_28176,N_27608,N_27859);
nor U28177 (N_28177,N_27709,N_27830);
nand U28178 (N_28178,N_27751,N_27710);
nor U28179 (N_28179,N_27773,N_27726);
nand U28180 (N_28180,N_27677,N_27810);
or U28181 (N_28181,N_27666,N_27764);
nand U28182 (N_28182,N_27765,N_27813);
nor U28183 (N_28183,N_27687,N_27856);
or U28184 (N_28184,N_27795,N_27605);
or U28185 (N_28185,N_27776,N_27649);
or U28186 (N_28186,N_27809,N_27628);
nor U28187 (N_28187,N_27660,N_27807);
xor U28188 (N_28188,N_27668,N_27729);
or U28189 (N_28189,N_27663,N_27701);
xor U28190 (N_28190,N_27893,N_27675);
xnor U28191 (N_28191,N_27820,N_27741);
nand U28192 (N_28192,N_27774,N_27822);
xnor U28193 (N_28193,N_27776,N_27839);
xor U28194 (N_28194,N_27808,N_27638);
and U28195 (N_28195,N_27823,N_27884);
nor U28196 (N_28196,N_27684,N_27861);
or U28197 (N_28197,N_27625,N_27679);
nand U28198 (N_28198,N_27780,N_27652);
or U28199 (N_28199,N_27768,N_27674);
nor U28200 (N_28200,N_28050,N_27916);
nand U28201 (N_28201,N_28107,N_28097);
nor U28202 (N_28202,N_27931,N_28052);
xor U28203 (N_28203,N_28112,N_28140);
xor U28204 (N_28204,N_28195,N_27935);
xor U28205 (N_28205,N_27929,N_28012);
and U28206 (N_28206,N_27982,N_28000);
xnor U28207 (N_28207,N_28113,N_27912);
xnor U28208 (N_28208,N_28077,N_28082);
xor U28209 (N_28209,N_27998,N_28046);
and U28210 (N_28210,N_28006,N_28119);
xor U28211 (N_28211,N_27960,N_28011);
nor U28212 (N_28212,N_28127,N_28180);
nand U28213 (N_28213,N_28122,N_27942);
and U28214 (N_28214,N_28089,N_27962);
nor U28215 (N_28215,N_28149,N_28146);
and U28216 (N_28216,N_28043,N_28185);
nor U28217 (N_28217,N_28060,N_27946);
xnor U28218 (N_28218,N_28019,N_27965);
xnor U28219 (N_28219,N_27990,N_27996);
and U28220 (N_28220,N_28069,N_27975);
nand U28221 (N_28221,N_28179,N_27902);
nand U28222 (N_28222,N_27988,N_28045);
or U28223 (N_28223,N_28135,N_28166);
or U28224 (N_28224,N_28121,N_28010);
or U28225 (N_28225,N_28198,N_27906);
xor U28226 (N_28226,N_28020,N_28015);
and U28227 (N_28227,N_27903,N_27986);
xnor U28228 (N_28228,N_27955,N_28147);
xnor U28229 (N_28229,N_28068,N_28001);
nand U28230 (N_28230,N_28144,N_27907);
or U28231 (N_28231,N_27980,N_28039);
xnor U28232 (N_28232,N_28062,N_28162);
xor U28233 (N_28233,N_28057,N_28025);
xor U28234 (N_28234,N_28067,N_28183);
nand U28235 (N_28235,N_28129,N_27908);
or U28236 (N_28236,N_27910,N_28114);
xnor U28237 (N_28237,N_28092,N_28111);
xor U28238 (N_28238,N_28037,N_28048);
xnor U28239 (N_28239,N_28073,N_27993);
nor U28240 (N_28240,N_28133,N_28141);
nor U28241 (N_28241,N_28079,N_28199);
or U28242 (N_28242,N_28059,N_27947);
and U28243 (N_28243,N_27969,N_28030);
and U28244 (N_28244,N_27951,N_27945);
xor U28245 (N_28245,N_27964,N_27983);
or U28246 (N_28246,N_28142,N_27926);
xnor U28247 (N_28247,N_27985,N_28017);
nor U28248 (N_28248,N_28053,N_28177);
and U28249 (N_28249,N_28158,N_27905);
xnor U28250 (N_28250,N_27914,N_27909);
nor U28251 (N_28251,N_28138,N_28044);
and U28252 (N_28252,N_28157,N_28153);
and U28253 (N_28253,N_28182,N_27977);
nor U28254 (N_28254,N_27958,N_28087);
and U28255 (N_28255,N_28118,N_27989);
or U28256 (N_28256,N_28194,N_28145);
nand U28257 (N_28257,N_27921,N_28174);
nand U28258 (N_28258,N_28058,N_27941);
or U28259 (N_28259,N_27987,N_28130);
nand U28260 (N_28260,N_27979,N_28120);
xnor U28261 (N_28261,N_27973,N_28086);
xor U28262 (N_28262,N_28131,N_27953);
and U28263 (N_28263,N_28159,N_28192);
nor U28264 (N_28264,N_28186,N_27928);
nor U28265 (N_28265,N_27924,N_28070);
nand U28266 (N_28266,N_28169,N_28190);
or U28267 (N_28267,N_27944,N_27938);
nand U28268 (N_28268,N_28023,N_28165);
or U28269 (N_28269,N_28061,N_28139);
and U28270 (N_28270,N_28102,N_27932);
and U28271 (N_28271,N_28007,N_28074);
nand U28272 (N_28272,N_28032,N_28103);
nand U28273 (N_28273,N_28160,N_27999);
nor U28274 (N_28274,N_28196,N_28066);
or U28275 (N_28275,N_28055,N_27957);
nand U28276 (N_28276,N_28095,N_27948);
or U28277 (N_28277,N_27934,N_28027);
xor U28278 (N_28278,N_28128,N_28108);
nor U28279 (N_28279,N_27963,N_27978);
and U28280 (N_28280,N_28187,N_28109);
or U28281 (N_28281,N_27997,N_28072);
xnor U28282 (N_28282,N_27919,N_28164);
nor U28283 (N_28283,N_28075,N_28099);
nand U28284 (N_28284,N_28167,N_28175);
nor U28285 (N_28285,N_27933,N_28098);
nor U28286 (N_28286,N_28110,N_28134);
nand U28287 (N_28287,N_28197,N_27954);
xnor U28288 (N_28288,N_28029,N_28151);
nand U28289 (N_28289,N_28143,N_28084);
or U28290 (N_28290,N_27995,N_28005);
nor U28291 (N_28291,N_27956,N_27915);
or U28292 (N_28292,N_28155,N_28105);
or U28293 (N_28293,N_28117,N_27991);
or U28294 (N_28294,N_28009,N_27959);
and U28295 (N_28295,N_27952,N_28170);
or U28296 (N_28296,N_27901,N_28085);
and U28297 (N_28297,N_28136,N_28014);
xor U28298 (N_28298,N_28028,N_27930);
nor U28299 (N_28299,N_28181,N_28026);
or U28300 (N_28300,N_28096,N_28191);
and U28301 (N_28301,N_28065,N_28163);
nand U28302 (N_28302,N_27940,N_28004);
xnor U28303 (N_28303,N_28115,N_28041);
nor U28304 (N_28304,N_27922,N_28184);
nand U28305 (N_28305,N_28040,N_27925);
nor U28306 (N_28306,N_28094,N_28063);
nand U28307 (N_28307,N_27970,N_27950);
or U28308 (N_28308,N_27904,N_28008);
nand U28309 (N_28309,N_28002,N_27937);
nand U28310 (N_28310,N_28064,N_28171);
nand U28311 (N_28311,N_27972,N_28154);
nand U28312 (N_28312,N_28080,N_28116);
or U28313 (N_28313,N_28172,N_27976);
and U28314 (N_28314,N_27923,N_28152);
nor U28315 (N_28315,N_27913,N_27936);
xor U28316 (N_28316,N_28056,N_27911);
nor U28317 (N_28317,N_28003,N_28013);
and U28318 (N_28318,N_28161,N_28178);
or U28319 (N_28319,N_27971,N_28137);
nor U28320 (N_28320,N_28071,N_28018);
and U28321 (N_28321,N_27992,N_28104);
xor U28322 (N_28322,N_27939,N_27917);
and U28323 (N_28323,N_28125,N_28173);
and U28324 (N_28324,N_27994,N_27966);
nor U28325 (N_28325,N_28035,N_28036);
nor U28326 (N_28326,N_28022,N_28093);
or U28327 (N_28327,N_27968,N_27961);
xor U28328 (N_28328,N_27981,N_28090);
nor U28329 (N_28329,N_27900,N_27920);
nand U28330 (N_28330,N_28031,N_28126);
xnor U28331 (N_28331,N_28193,N_28189);
xnor U28332 (N_28332,N_28049,N_28168);
nor U28333 (N_28333,N_28054,N_28132);
nand U28334 (N_28334,N_28176,N_28021);
nor U28335 (N_28335,N_28106,N_27984);
and U28336 (N_28336,N_27927,N_27949);
or U28337 (N_28337,N_28076,N_28100);
nand U28338 (N_28338,N_28148,N_28083);
or U28339 (N_28339,N_28124,N_28047);
nand U28340 (N_28340,N_27918,N_28042);
xor U28341 (N_28341,N_28150,N_28156);
and U28342 (N_28342,N_28024,N_28101);
nand U28343 (N_28343,N_27943,N_28088);
or U28344 (N_28344,N_28078,N_28051);
or U28345 (N_28345,N_28188,N_27974);
nand U28346 (N_28346,N_28016,N_28033);
and U28347 (N_28347,N_28038,N_28123);
nand U28348 (N_28348,N_28091,N_28081);
nand U28349 (N_28349,N_28034,N_27967);
xnor U28350 (N_28350,N_28119,N_27958);
nand U28351 (N_28351,N_28071,N_28029);
nor U28352 (N_28352,N_28197,N_28117);
xnor U28353 (N_28353,N_28115,N_28191);
nand U28354 (N_28354,N_28121,N_28132);
xnor U28355 (N_28355,N_28133,N_28152);
nand U28356 (N_28356,N_28131,N_28141);
nand U28357 (N_28357,N_27982,N_28186);
nor U28358 (N_28358,N_27960,N_27932);
xor U28359 (N_28359,N_28142,N_28141);
nor U28360 (N_28360,N_27949,N_28039);
and U28361 (N_28361,N_27934,N_28038);
nor U28362 (N_28362,N_28072,N_28102);
or U28363 (N_28363,N_28022,N_28089);
nor U28364 (N_28364,N_28008,N_27936);
nor U28365 (N_28365,N_27971,N_28120);
nor U28366 (N_28366,N_28149,N_27969);
or U28367 (N_28367,N_28168,N_28035);
nor U28368 (N_28368,N_28180,N_28119);
nand U28369 (N_28369,N_27986,N_28125);
or U28370 (N_28370,N_28051,N_28106);
nor U28371 (N_28371,N_28024,N_28191);
xor U28372 (N_28372,N_28018,N_28182);
or U28373 (N_28373,N_27953,N_28158);
nor U28374 (N_28374,N_28189,N_28183);
nor U28375 (N_28375,N_28070,N_28063);
nor U28376 (N_28376,N_27943,N_28121);
xnor U28377 (N_28377,N_27903,N_28170);
nor U28378 (N_28378,N_28196,N_28167);
nand U28379 (N_28379,N_27979,N_28121);
xor U28380 (N_28380,N_27983,N_27931);
or U28381 (N_28381,N_28119,N_28070);
nor U28382 (N_28382,N_28010,N_27909);
nand U28383 (N_28383,N_28053,N_27979);
and U28384 (N_28384,N_27906,N_27945);
or U28385 (N_28385,N_28017,N_28163);
nor U28386 (N_28386,N_27961,N_28113);
or U28387 (N_28387,N_28109,N_28080);
nand U28388 (N_28388,N_27965,N_27912);
and U28389 (N_28389,N_28136,N_28072);
nand U28390 (N_28390,N_27948,N_28074);
xor U28391 (N_28391,N_28104,N_27962);
nor U28392 (N_28392,N_27943,N_28051);
xnor U28393 (N_28393,N_27914,N_27969);
nor U28394 (N_28394,N_27916,N_27932);
xnor U28395 (N_28395,N_28016,N_28070);
nand U28396 (N_28396,N_27967,N_28066);
nand U28397 (N_28397,N_28079,N_27905);
or U28398 (N_28398,N_27978,N_27959);
or U28399 (N_28399,N_27938,N_27936);
or U28400 (N_28400,N_27936,N_27949);
nand U28401 (N_28401,N_27927,N_28001);
nor U28402 (N_28402,N_27901,N_28197);
and U28403 (N_28403,N_28126,N_27985);
nor U28404 (N_28404,N_27913,N_27941);
or U28405 (N_28405,N_28009,N_27931);
nand U28406 (N_28406,N_28006,N_27909);
nor U28407 (N_28407,N_28106,N_27938);
and U28408 (N_28408,N_27995,N_27937);
nor U28409 (N_28409,N_27941,N_28056);
nand U28410 (N_28410,N_28015,N_27975);
or U28411 (N_28411,N_28103,N_28052);
nor U28412 (N_28412,N_28138,N_27925);
nor U28413 (N_28413,N_28120,N_27914);
or U28414 (N_28414,N_28145,N_28046);
xnor U28415 (N_28415,N_28077,N_28116);
or U28416 (N_28416,N_28101,N_28038);
nand U28417 (N_28417,N_28046,N_27960);
and U28418 (N_28418,N_28115,N_28110);
xor U28419 (N_28419,N_28122,N_28172);
or U28420 (N_28420,N_27970,N_27941);
nor U28421 (N_28421,N_28030,N_27924);
nor U28422 (N_28422,N_27970,N_27918);
nand U28423 (N_28423,N_27965,N_27927);
and U28424 (N_28424,N_27911,N_27999);
or U28425 (N_28425,N_28074,N_28089);
nor U28426 (N_28426,N_28164,N_28002);
xor U28427 (N_28427,N_28068,N_28110);
nor U28428 (N_28428,N_28092,N_27967);
nand U28429 (N_28429,N_28106,N_27988);
or U28430 (N_28430,N_28171,N_27931);
nor U28431 (N_28431,N_28153,N_28174);
nand U28432 (N_28432,N_28172,N_28011);
or U28433 (N_28433,N_27932,N_28058);
nor U28434 (N_28434,N_27918,N_28180);
or U28435 (N_28435,N_28112,N_27915);
nand U28436 (N_28436,N_27999,N_28046);
xnor U28437 (N_28437,N_28185,N_27921);
nor U28438 (N_28438,N_27938,N_28079);
nor U28439 (N_28439,N_28110,N_28052);
nor U28440 (N_28440,N_28180,N_28043);
or U28441 (N_28441,N_27985,N_28184);
xor U28442 (N_28442,N_28183,N_27963);
nor U28443 (N_28443,N_28068,N_28062);
and U28444 (N_28444,N_28110,N_28159);
nor U28445 (N_28445,N_27933,N_28029);
nor U28446 (N_28446,N_28117,N_28151);
or U28447 (N_28447,N_27964,N_28093);
nor U28448 (N_28448,N_27914,N_28000);
nand U28449 (N_28449,N_28132,N_27912);
nand U28450 (N_28450,N_27966,N_27936);
nand U28451 (N_28451,N_28094,N_28120);
or U28452 (N_28452,N_28026,N_28017);
nand U28453 (N_28453,N_28064,N_28030);
and U28454 (N_28454,N_27966,N_28076);
nor U28455 (N_28455,N_27976,N_28006);
or U28456 (N_28456,N_27977,N_28108);
xnor U28457 (N_28457,N_28041,N_28027);
or U28458 (N_28458,N_28184,N_28005);
xor U28459 (N_28459,N_28139,N_28191);
or U28460 (N_28460,N_28014,N_27917);
or U28461 (N_28461,N_28105,N_27980);
and U28462 (N_28462,N_27946,N_28028);
xor U28463 (N_28463,N_28009,N_28027);
nand U28464 (N_28464,N_28157,N_27981);
nand U28465 (N_28465,N_27995,N_28022);
or U28466 (N_28466,N_27914,N_28070);
nor U28467 (N_28467,N_28101,N_27982);
xor U28468 (N_28468,N_28081,N_28072);
and U28469 (N_28469,N_28153,N_28139);
and U28470 (N_28470,N_28127,N_28153);
or U28471 (N_28471,N_28180,N_27937);
xor U28472 (N_28472,N_28070,N_27921);
and U28473 (N_28473,N_28195,N_28181);
xnor U28474 (N_28474,N_28019,N_28078);
and U28475 (N_28475,N_27932,N_28156);
nand U28476 (N_28476,N_28096,N_28126);
xor U28477 (N_28477,N_27947,N_28072);
and U28478 (N_28478,N_28136,N_28086);
and U28479 (N_28479,N_27918,N_27917);
xnor U28480 (N_28480,N_28182,N_28110);
nand U28481 (N_28481,N_28097,N_28106);
xnor U28482 (N_28482,N_28028,N_27989);
or U28483 (N_28483,N_27994,N_27915);
or U28484 (N_28484,N_28085,N_27982);
xnor U28485 (N_28485,N_28158,N_27992);
or U28486 (N_28486,N_28056,N_27996);
nor U28487 (N_28487,N_27907,N_27949);
nor U28488 (N_28488,N_28177,N_27981);
xnor U28489 (N_28489,N_28035,N_28122);
and U28490 (N_28490,N_28138,N_27959);
xor U28491 (N_28491,N_28117,N_28022);
nor U28492 (N_28492,N_28182,N_27998);
xnor U28493 (N_28493,N_28118,N_28030);
nand U28494 (N_28494,N_27998,N_27902);
nor U28495 (N_28495,N_28096,N_28014);
and U28496 (N_28496,N_27985,N_27913);
nand U28497 (N_28497,N_27952,N_28171);
nor U28498 (N_28498,N_28091,N_28117);
nor U28499 (N_28499,N_27989,N_28020);
nor U28500 (N_28500,N_28330,N_28464);
or U28501 (N_28501,N_28429,N_28275);
nand U28502 (N_28502,N_28422,N_28311);
nand U28503 (N_28503,N_28489,N_28231);
nor U28504 (N_28504,N_28423,N_28325);
and U28505 (N_28505,N_28286,N_28200);
nand U28506 (N_28506,N_28449,N_28332);
or U28507 (N_28507,N_28333,N_28425);
or U28508 (N_28508,N_28480,N_28440);
nor U28509 (N_28509,N_28498,N_28383);
and U28510 (N_28510,N_28267,N_28209);
xor U28511 (N_28511,N_28445,N_28379);
or U28512 (N_28512,N_28236,N_28278);
nor U28513 (N_28513,N_28315,N_28321);
nor U28514 (N_28514,N_28309,N_28451);
nand U28515 (N_28515,N_28388,N_28202);
nand U28516 (N_28516,N_28214,N_28443);
xnor U28517 (N_28517,N_28351,N_28326);
nand U28518 (N_28518,N_28446,N_28274);
nand U28519 (N_28519,N_28312,N_28226);
or U28520 (N_28520,N_28413,N_28466);
and U28521 (N_28521,N_28385,N_28428);
and U28522 (N_28522,N_28346,N_28328);
and U28523 (N_28523,N_28320,N_28465);
and U28524 (N_28524,N_28256,N_28453);
xor U28525 (N_28525,N_28387,N_28353);
xnor U28526 (N_28526,N_28350,N_28363);
or U28527 (N_28527,N_28303,N_28481);
xor U28528 (N_28528,N_28486,N_28461);
xnor U28529 (N_28529,N_28241,N_28458);
nor U28530 (N_28530,N_28477,N_28245);
nor U28531 (N_28531,N_28397,N_28239);
nand U28532 (N_28532,N_28225,N_28365);
and U28533 (N_28533,N_28483,N_28374);
or U28534 (N_28534,N_28433,N_28349);
or U28535 (N_28535,N_28475,N_28364);
nor U28536 (N_28536,N_28289,N_28336);
and U28537 (N_28537,N_28487,N_28265);
and U28538 (N_28538,N_28427,N_28484);
or U28539 (N_28539,N_28208,N_28287);
nor U28540 (N_28540,N_28400,N_28248);
nor U28541 (N_28541,N_28213,N_28401);
or U28542 (N_28542,N_28264,N_28409);
or U28543 (N_28543,N_28369,N_28235);
nand U28544 (N_28544,N_28368,N_28493);
nand U28545 (N_28545,N_28244,N_28420);
nand U28546 (N_28546,N_28393,N_28259);
or U28547 (N_28547,N_28292,N_28270);
nand U28548 (N_28548,N_28459,N_28468);
xor U28549 (N_28549,N_28447,N_28436);
or U28550 (N_28550,N_28279,N_28306);
and U28551 (N_28551,N_28347,N_28485);
nor U28552 (N_28552,N_28367,N_28340);
nand U28553 (N_28553,N_28450,N_28492);
nor U28554 (N_28554,N_28419,N_28377);
or U28555 (N_28555,N_28212,N_28405);
or U28556 (N_28556,N_28354,N_28372);
or U28557 (N_28557,N_28271,N_28233);
nand U28558 (N_28558,N_28399,N_28373);
and U28559 (N_28559,N_28358,N_28282);
or U28560 (N_28560,N_28201,N_28253);
and U28561 (N_28561,N_28389,N_28276);
nor U28562 (N_28562,N_28316,N_28403);
or U28563 (N_28563,N_28227,N_28479);
nand U28564 (N_28564,N_28232,N_28307);
nand U28565 (N_28565,N_28293,N_28376);
nand U28566 (N_28566,N_28291,N_28331);
nand U28567 (N_28567,N_28497,N_28421);
nand U28568 (N_28568,N_28207,N_28412);
or U28569 (N_28569,N_28448,N_28476);
and U28570 (N_28570,N_28470,N_28246);
nor U28571 (N_28571,N_28402,N_28426);
xnor U28572 (N_28572,N_28452,N_28215);
or U28573 (N_28573,N_28310,N_28277);
nand U28574 (N_28574,N_28495,N_28472);
or U28575 (N_28575,N_28488,N_28304);
xnor U28576 (N_28576,N_28444,N_28255);
and U28577 (N_28577,N_28318,N_28268);
nor U28578 (N_28578,N_28378,N_28357);
nand U28579 (N_28579,N_28366,N_28273);
or U28580 (N_28580,N_28308,N_28237);
or U28581 (N_28581,N_28414,N_28299);
or U28582 (N_28582,N_28345,N_28352);
and U28583 (N_28583,N_28211,N_28473);
nand U28584 (N_28584,N_28240,N_28348);
and U28585 (N_28585,N_28281,N_28272);
and U28586 (N_28586,N_28329,N_28482);
or U28587 (N_28587,N_28390,N_28242);
nand U28588 (N_28588,N_28437,N_28284);
and U28589 (N_28589,N_28398,N_28324);
nand U28590 (N_28590,N_28362,N_28355);
or U28591 (N_28591,N_28234,N_28218);
nand U28592 (N_28592,N_28294,N_28204);
and U28593 (N_28593,N_28296,N_28463);
and U28594 (N_28594,N_28314,N_28381);
xnor U28595 (N_28595,N_28396,N_28406);
and U28596 (N_28596,N_28408,N_28229);
xor U28597 (N_28597,N_28221,N_28343);
nor U28598 (N_28598,N_28260,N_28471);
nor U28599 (N_28599,N_28300,N_28432);
xor U28600 (N_28600,N_28219,N_28210);
or U28601 (N_28601,N_28417,N_28243);
nand U28602 (N_28602,N_28317,N_28410);
and U28603 (N_28603,N_28261,N_28431);
nor U28604 (N_28604,N_28395,N_28490);
and U28605 (N_28605,N_28462,N_28305);
xor U28606 (N_28606,N_28205,N_28382);
xor U28607 (N_28607,N_28430,N_28418);
nand U28608 (N_28608,N_28356,N_28249);
and U28609 (N_28609,N_28258,N_28337);
or U28610 (N_28610,N_28375,N_28435);
nor U28611 (N_28611,N_28251,N_28335);
nor U28612 (N_28612,N_28301,N_28285);
nand U28613 (N_28613,N_28361,N_28323);
xor U28614 (N_28614,N_28206,N_28220);
nand U28615 (N_28615,N_28460,N_28262);
or U28616 (N_28616,N_28371,N_28384);
and U28617 (N_28617,N_28394,N_28334);
xnor U28618 (N_28618,N_28416,N_28454);
and U28619 (N_28619,N_28288,N_28456);
nand U28620 (N_28620,N_28469,N_28230);
or U28621 (N_28621,N_28467,N_28203);
and U28622 (N_28622,N_28491,N_28341);
nor U28623 (N_28623,N_28359,N_28499);
and U28624 (N_28624,N_28344,N_28302);
nor U28625 (N_28625,N_28455,N_28434);
nand U28626 (N_28626,N_28238,N_28266);
nand U28627 (N_28627,N_28247,N_28338);
nand U28628 (N_28628,N_28250,N_28280);
nor U28629 (N_28629,N_28252,N_28327);
nand U28630 (N_28630,N_28222,N_28339);
nor U28631 (N_28631,N_28342,N_28283);
nor U28632 (N_28632,N_28392,N_28313);
xor U28633 (N_28633,N_28439,N_28415);
nand U28634 (N_28634,N_28297,N_28228);
or U28635 (N_28635,N_28404,N_28263);
nand U28636 (N_28636,N_28223,N_28474);
or U28637 (N_28637,N_28496,N_28424);
and U28638 (N_28638,N_28295,N_28442);
or U28639 (N_28639,N_28254,N_28217);
nand U28640 (N_28640,N_28319,N_28269);
or U28641 (N_28641,N_28386,N_28411);
nand U28642 (N_28642,N_28290,N_28298);
nor U28643 (N_28643,N_28216,N_28380);
xnor U28644 (N_28644,N_28407,N_28257);
nand U28645 (N_28645,N_28224,N_28441);
nand U28646 (N_28646,N_28391,N_28438);
or U28647 (N_28647,N_28322,N_28457);
xor U28648 (N_28648,N_28360,N_28494);
or U28649 (N_28649,N_28370,N_28478);
nor U28650 (N_28650,N_28310,N_28420);
and U28651 (N_28651,N_28481,N_28374);
and U28652 (N_28652,N_28241,N_28237);
nand U28653 (N_28653,N_28200,N_28433);
xor U28654 (N_28654,N_28437,N_28333);
nand U28655 (N_28655,N_28323,N_28248);
and U28656 (N_28656,N_28490,N_28239);
and U28657 (N_28657,N_28221,N_28487);
or U28658 (N_28658,N_28389,N_28349);
and U28659 (N_28659,N_28345,N_28255);
xor U28660 (N_28660,N_28427,N_28486);
xor U28661 (N_28661,N_28485,N_28468);
nand U28662 (N_28662,N_28325,N_28334);
nand U28663 (N_28663,N_28216,N_28264);
nor U28664 (N_28664,N_28351,N_28245);
nor U28665 (N_28665,N_28299,N_28422);
or U28666 (N_28666,N_28452,N_28263);
and U28667 (N_28667,N_28460,N_28231);
and U28668 (N_28668,N_28281,N_28462);
and U28669 (N_28669,N_28434,N_28334);
xnor U28670 (N_28670,N_28461,N_28491);
or U28671 (N_28671,N_28442,N_28471);
nor U28672 (N_28672,N_28254,N_28251);
nand U28673 (N_28673,N_28251,N_28271);
nor U28674 (N_28674,N_28447,N_28218);
or U28675 (N_28675,N_28312,N_28470);
xnor U28676 (N_28676,N_28340,N_28347);
nor U28677 (N_28677,N_28382,N_28294);
nand U28678 (N_28678,N_28474,N_28314);
xnor U28679 (N_28679,N_28359,N_28232);
xnor U28680 (N_28680,N_28417,N_28407);
nor U28681 (N_28681,N_28312,N_28488);
nand U28682 (N_28682,N_28490,N_28274);
nand U28683 (N_28683,N_28463,N_28426);
nor U28684 (N_28684,N_28380,N_28220);
nand U28685 (N_28685,N_28359,N_28282);
xor U28686 (N_28686,N_28261,N_28365);
nand U28687 (N_28687,N_28398,N_28491);
nand U28688 (N_28688,N_28255,N_28342);
xnor U28689 (N_28689,N_28359,N_28368);
xor U28690 (N_28690,N_28493,N_28370);
xor U28691 (N_28691,N_28343,N_28365);
xnor U28692 (N_28692,N_28419,N_28271);
or U28693 (N_28693,N_28437,N_28343);
xor U28694 (N_28694,N_28206,N_28279);
nand U28695 (N_28695,N_28302,N_28326);
nor U28696 (N_28696,N_28368,N_28310);
nor U28697 (N_28697,N_28240,N_28431);
and U28698 (N_28698,N_28475,N_28207);
nand U28699 (N_28699,N_28308,N_28346);
xor U28700 (N_28700,N_28437,N_28424);
nand U28701 (N_28701,N_28357,N_28244);
nand U28702 (N_28702,N_28335,N_28407);
nand U28703 (N_28703,N_28321,N_28403);
xor U28704 (N_28704,N_28419,N_28260);
or U28705 (N_28705,N_28336,N_28234);
nand U28706 (N_28706,N_28411,N_28320);
nor U28707 (N_28707,N_28406,N_28353);
xnor U28708 (N_28708,N_28320,N_28210);
or U28709 (N_28709,N_28341,N_28219);
and U28710 (N_28710,N_28380,N_28474);
nand U28711 (N_28711,N_28315,N_28482);
xor U28712 (N_28712,N_28321,N_28285);
nand U28713 (N_28713,N_28477,N_28463);
xnor U28714 (N_28714,N_28259,N_28476);
nor U28715 (N_28715,N_28271,N_28493);
nor U28716 (N_28716,N_28360,N_28239);
xnor U28717 (N_28717,N_28494,N_28246);
xnor U28718 (N_28718,N_28328,N_28399);
nand U28719 (N_28719,N_28402,N_28363);
xnor U28720 (N_28720,N_28348,N_28443);
and U28721 (N_28721,N_28361,N_28278);
and U28722 (N_28722,N_28428,N_28225);
nand U28723 (N_28723,N_28481,N_28348);
or U28724 (N_28724,N_28256,N_28251);
or U28725 (N_28725,N_28451,N_28333);
xnor U28726 (N_28726,N_28487,N_28485);
xor U28727 (N_28727,N_28483,N_28464);
or U28728 (N_28728,N_28291,N_28250);
xor U28729 (N_28729,N_28302,N_28465);
or U28730 (N_28730,N_28447,N_28349);
and U28731 (N_28731,N_28295,N_28459);
nand U28732 (N_28732,N_28386,N_28272);
or U28733 (N_28733,N_28388,N_28230);
nand U28734 (N_28734,N_28393,N_28403);
nor U28735 (N_28735,N_28267,N_28361);
or U28736 (N_28736,N_28453,N_28396);
nand U28737 (N_28737,N_28390,N_28480);
nand U28738 (N_28738,N_28424,N_28379);
nand U28739 (N_28739,N_28296,N_28397);
nor U28740 (N_28740,N_28237,N_28425);
nor U28741 (N_28741,N_28347,N_28422);
nor U28742 (N_28742,N_28419,N_28270);
or U28743 (N_28743,N_28222,N_28200);
nand U28744 (N_28744,N_28285,N_28235);
xnor U28745 (N_28745,N_28246,N_28407);
and U28746 (N_28746,N_28341,N_28407);
or U28747 (N_28747,N_28464,N_28303);
nand U28748 (N_28748,N_28428,N_28345);
or U28749 (N_28749,N_28386,N_28329);
nand U28750 (N_28750,N_28469,N_28296);
xnor U28751 (N_28751,N_28336,N_28231);
and U28752 (N_28752,N_28218,N_28307);
nand U28753 (N_28753,N_28360,N_28444);
nor U28754 (N_28754,N_28279,N_28357);
and U28755 (N_28755,N_28229,N_28297);
xnor U28756 (N_28756,N_28282,N_28426);
nor U28757 (N_28757,N_28265,N_28240);
nor U28758 (N_28758,N_28330,N_28489);
nand U28759 (N_28759,N_28283,N_28297);
nor U28760 (N_28760,N_28299,N_28214);
xor U28761 (N_28761,N_28356,N_28464);
nand U28762 (N_28762,N_28325,N_28320);
xor U28763 (N_28763,N_28374,N_28275);
nor U28764 (N_28764,N_28267,N_28394);
nand U28765 (N_28765,N_28235,N_28415);
or U28766 (N_28766,N_28466,N_28239);
xor U28767 (N_28767,N_28212,N_28322);
nand U28768 (N_28768,N_28286,N_28444);
xor U28769 (N_28769,N_28201,N_28232);
nor U28770 (N_28770,N_28290,N_28354);
or U28771 (N_28771,N_28456,N_28475);
xor U28772 (N_28772,N_28405,N_28328);
nand U28773 (N_28773,N_28366,N_28491);
and U28774 (N_28774,N_28476,N_28316);
xor U28775 (N_28775,N_28307,N_28256);
or U28776 (N_28776,N_28413,N_28486);
or U28777 (N_28777,N_28357,N_28460);
and U28778 (N_28778,N_28247,N_28402);
or U28779 (N_28779,N_28289,N_28215);
nor U28780 (N_28780,N_28389,N_28330);
nand U28781 (N_28781,N_28423,N_28266);
xnor U28782 (N_28782,N_28249,N_28418);
and U28783 (N_28783,N_28260,N_28323);
nand U28784 (N_28784,N_28467,N_28285);
and U28785 (N_28785,N_28255,N_28295);
nand U28786 (N_28786,N_28245,N_28241);
or U28787 (N_28787,N_28444,N_28248);
nand U28788 (N_28788,N_28327,N_28443);
nor U28789 (N_28789,N_28219,N_28218);
nand U28790 (N_28790,N_28417,N_28481);
xor U28791 (N_28791,N_28368,N_28286);
xnor U28792 (N_28792,N_28461,N_28324);
xor U28793 (N_28793,N_28375,N_28417);
nor U28794 (N_28794,N_28397,N_28499);
xor U28795 (N_28795,N_28287,N_28498);
xnor U28796 (N_28796,N_28243,N_28212);
nor U28797 (N_28797,N_28352,N_28436);
or U28798 (N_28798,N_28414,N_28221);
xor U28799 (N_28799,N_28236,N_28468);
xnor U28800 (N_28800,N_28712,N_28735);
nand U28801 (N_28801,N_28641,N_28761);
xnor U28802 (N_28802,N_28635,N_28640);
and U28803 (N_28803,N_28526,N_28557);
xor U28804 (N_28804,N_28704,N_28611);
or U28805 (N_28805,N_28500,N_28749);
or U28806 (N_28806,N_28779,N_28796);
nor U28807 (N_28807,N_28548,N_28577);
or U28808 (N_28808,N_28503,N_28628);
xnor U28809 (N_28809,N_28709,N_28639);
xnor U28810 (N_28810,N_28703,N_28584);
nand U28811 (N_28811,N_28513,N_28676);
nand U28812 (N_28812,N_28595,N_28520);
or U28813 (N_28813,N_28614,N_28581);
or U28814 (N_28814,N_28666,N_28524);
xor U28815 (N_28815,N_28619,N_28592);
xnor U28816 (N_28816,N_28786,N_28782);
nor U28817 (N_28817,N_28732,N_28508);
nor U28818 (N_28818,N_28522,N_28701);
nand U28819 (N_28819,N_28665,N_28682);
or U28820 (N_28820,N_28776,N_28572);
xnor U28821 (N_28821,N_28751,N_28759);
nand U28822 (N_28822,N_28783,N_28724);
nor U28823 (N_28823,N_28609,N_28693);
nor U28824 (N_28824,N_28564,N_28723);
xor U28825 (N_28825,N_28634,N_28718);
and U28826 (N_28826,N_28604,N_28558);
xor U28827 (N_28827,N_28714,N_28504);
and U28828 (N_28828,N_28578,N_28667);
xor U28829 (N_28829,N_28556,N_28650);
and U28830 (N_28830,N_28729,N_28502);
and U28831 (N_28831,N_28618,N_28711);
and U28832 (N_28832,N_28763,N_28661);
or U28833 (N_28833,N_28744,N_28766);
nand U28834 (N_28834,N_28510,N_28629);
nor U28835 (N_28835,N_28638,N_28659);
nor U28836 (N_28836,N_28683,N_28784);
nor U28837 (N_28837,N_28599,N_28617);
nor U28838 (N_28838,N_28746,N_28725);
nor U28839 (N_28839,N_28575,N_28752);
nor U28840 (N_28840,N_28603,N_28764);
or U28841 (N_28841,N_28625,N_28540);
nand U28842 (N_28842,N_28553,N_28538);
nand U28843 (N_28843,N_28760,N_28535);
xor U28844 (N_28844,N_28602,N_28569);
nor U28845 (N_28845,N_28546,N_28792);
nand U28846 (N_28846,N_28612,N_28598);
nor U28847 (N_28847,N_28663,N_28728);
or U28848 (N_28848,N_28610,N_28527);
nor U28849 (N_28849,N_28621,N_28799);
xnor U28850 (N_28850,N_28547,N_28791);
xor U28851 (N_28851,N_28565,N_28566);
nor U28852 (N_28852,N_28632,N_28669);
xnor U28853 (N_28853,N_28787,N_28793);
nor U28854 (N_28854,N_28652,N_28739);
or U28855 (N_28855,N_28771,N_28530);
nor U28856 (N_28856,N_28798,N_28658);
or U28857 (N_28857,N_28708,N_28631);
nor U28858 (N_28858,N_28644,N_28673);
xnor U28859 (N_28859,N_28685,N_28675);
or U28860 (N_28860,N_28554,N_28509);
and U28861 (N_28861,N_28545,N_28706);
or U28862 (N_28862,N_28608,N_28710);
nand U28863 (N_28863,N_28778,N_28774);
nor U28864 (N_28864,N_28529,N_28506);
nand U28865 (N_28865,N_28576,N_28533);
xnor U28866 (N_28866,N_28742,N_28505);
and U28867 (N_28867,N_28624,N_28660);
nor U28868 (N_28868,N_28767,N_28636);
and U28869 (N_28869,N_28637,N_28551);
nand U28870 (N_28870,N_28594,N_28544);
nand U28871 (N_28871,N_28717,N_28588);
nor U28872 (N_28872,N_28656,N_28626);
nand U28873 (N_28873,N_28720,N_28773);
and U28874 (N_28874,N_28563,N_28597);
xor U28875 (N_28875,N_28668,N_28698);
nand U28876 (N_28876,N_28688,N_28605);
nor U28877 (N_28877,N_28507,N_28737);
or U28878 (N_28878,N_28756,N_28549);
or U28879 (N_28879,N_28573,N_28654);
nand U28880 (N_28880,N_28672,N_28700);
nor U28881 (N_28881,N_28689,N_28516);
or U28882 (N_28882,N_28586,N_28519);
nor U28883 (N_28883,N_28550,N_28757);
and U28884 (N_28884,N_28731,N_28726);
nand U28885 (N_28885,N_28696,N_28517);
and U28886 (N_28886,N_28590,N_28733);
nand U28887 (N_28887,N_28579,N_28679);
and U28888 (N_28888,N_28699,N_28606);
nand U28889 (N_28889,N_28713,N_28562);
and U28890 (N_28890,N_28568,N_28600);
nand U28891 (N_28891,N_28657,N_28531);
nand U28892 (N_28892,N_28738,N_28781);
nand U28893 (N_28893,N_28601,N_28705);
xor U28894 (N_28894,N_28518,N_28747);
nor U28895 (N_28895,N_28677,N_28753);
or U28896 (N_28896,N_28662,N_28647);
nand U28897 (N_28897,N_28559,N_28691);
nor U28898 (N_28898,N_28543,N_28511);
nand U28899 (N_28899,N_28722,N_28697);
nor U28900 (N_28900,N_28646,N_28670);
nand U28901 (N_28901,N_28539,N_28740);
nand U28902 (N_28902,N_28648,N_28620);
nor U28903 (N_28903,N_28580,N_28583);
nand U28904 (N_28904,N_28521,N_28555);
and U28905 (N_28905,N_28643,N_28765);
nor U28906 (N_28906,N_28772,N_28645);
or U28907 (N_28907,N_28552,N_28775);
nand U28908 (N_28908,N_28736,N_28719);
or U28909 (N_28909,N_28541,N_28622);
nor U28910 (N_28910,N_28630,N_28587);
and U28911 (N_28911,N_28748,N_28585);
nor U28912 (N_28912,N_28567,N_28542);
nor U28913 (N_28913,N_28694,N_28750);
and U28914 (N_28914,N_28754,N_28777);
nand U28915 (N_28915,N_28570,N_28741);
and U28916 (N_28916,N_28797,N_28780);
nor U28917 (N_28917,N_28690,N_28616);
or U28918 (N_28918,N_28649,N_28615);
xnor U28919 (N_28919,N_28515,N_28642);
or U28920 (N_28920,N_28655,N_28727);
or U28921 (N_28921,N_28591,N_28523);
and U28922 (N_28922,N_28664,N_28534);
nor U28923 (N_28923,N_28743,N_28790);
or U28924 (N_28924,N_28687,N_28758);
nor U28925 (N_28925,N_28762,N_28755);
nand U28926 (N_28926,N_28536,N_28715);
and U28927 (N_28927,N_28653,N_28627);
nand U28928 (N_28928,N_28528,N_28769);
xor U28929 (N_28929,N_28734,N_28607);
and U28930 (N_28930,N_28692,N_28525);
xnor U28931 (N_28931,N_28671,N_28684);
nand U28932 (N_28932,N_28721,N_28571);
and U28933 (N_28933,N_28561,N_28596);
nand U28934 (N_28934,N_28770,N_28789);
nand U28935 (N_28935,N_28532,N_28651);
nor U28936 (N_28936,N_28681,N_28745);
nor U28937 (N_28937,N_28589,N_28613);
xor U28938 (N_28938,N_28788,N_28707);
and U28939 (N_28939,N_28702,N_28695);
nor U28940 (N_28940,N_28560,N_28501);
xor U28941 (N_28941,N_28680,N_28623);
and U28942 (N_28942,N_28785,N_28768);
nand U28943 (N_28943,N_28674,N_28716);
and U28944 (N_28944,N_28794,N_28574);
nor U28945 (N_28945,N_28593,N_28795);
nand U28946 (N_28946,N_28512,N_28582);
and U28947 (N_28947,N_28537,N_28730);
and U28948 (N_28948,N_28686,N_28633);
nor U28949 (N_28949,N_28678,N_28514);
nand U28950 (N_28950,N_28792,N_28617);
nand U28951 (N_28951,N_28543,N_28555);
xor U28952 (N_28952,N_28652,N_28775);
and U28953 (N_28953,N_28700,N_28663);
and U28954 (N_28954,N_28575,N_28598);
and U28955 (N_28955,N_28790,N_28534);
nand U28956 (N_28956,N_28586,N_28751);
nand U28957 (N_28957,N_28637,N_28728);
nor U28958 (N_28958,N_28624,N_28623);
nor U28959 (N_28959,N_28620,N_28616);
nand U28960 (N_28960,N_28569,N_28653);
nand U28961 (N_28961,N_28607,N_28648);
or U28962 (N_28962,N_28710,N_28556);
or U28963 (N_28963,N_28742,N_28743);
xor U28964 (N_28964,N_28699,N_28679);
or U28965 (N_28965,N_28718,N_28576);
nand U28966 (N_28966,N_28632,N_28750);
xnor U28967 (N_28967,N_28546,N_28731);
and U28968 (N_28968,N_28781,N_28721);
nor U28969 (N_28969,N_28777,N_28514);
nor U28970 (N_28970,N_28671,N_28775);
or U28971 (N_28971,N_28654,N_28627);
xnor U28972 (N_28972,N_28758,N_28786);
and U28973 (N_28973,N_28649,N_28713);
or U28974 (N_28974,N_28753,N_28623);
nand U28975 (N_28975,N_28563,N_28792);
or U28976 (N_28976,N_28788,N_28754);
nand U28977 (N_28977,N_28696,N_28650);
nand U28978 (N_28978,N_28628,N_28773);
or U28979 (N_28979,N_28686,N_28770);
nor U28980 (N_28980,N_28663,N_28584);
or U28981 (N_28981,N_28572,N_28501);
and U28982 (N_28982,N_28773,N_28789);
nand U28983 (N_28983,N_28584,N_28675);
or U28984 (N_28984,N_28565,N_28528);
and U28985 (N_28985,N_28513,N_28604);
xnor U28986 (N_28986,N_28750,N_28690);
or U28987 (N_28987,N_28737,N_28780);
and U28988 (N_28988,N_28508,N_28687);
and U28989 (N_28989,N_28610,N_28514);
and U28990 (N_28990,N_28674,N_28690);
and U28991 (N_28991,N_28560,N_28710);
nand U28992 (N_28992,N_28572,N_28599);
or U28993 (N_28993,N_28654,N_28503);
or U28994 (N_28994,N_28693,N_28596);
and U28995 (N_28995,N_28549,N_28602);
or U28996 (N_28996,N_28755,N_28506);
xnor U28997 (N_28997,N_28644,N_28636);
and U28998 (N_28998,N_28790,N_28501);
or U28999 (N_28999,N_28523,N_28552);
or U29000 (N_29000,N_28567,N_28759);
nor U29001 (N_29001,N_28544,N_28513);
and U29002 (N_29002,N_28718,N_28510);
and U29003 (N_29003,N_28664,N_28574);
nand U29004 (N_29004,N_28553,N_28565);
xnor U29005 (N_29005,N_28751,N_28686);
or U29006 (N_29006,N_28693,N_28681);
and U29007 (N_29007,N_28713,N_28522);
and U29008 (N_29008,N_28717,N_28526);
and U29009 (N_29009,N_28600,N_28748);
and U29010 (N_29010,N_28684,N_28675);
or U29011 (N_29011,N_28574,N_28646);
or U29012 (N_29012,N_28633,N_28678);
nor U29013 (N_29013,N_28725,N_28519);
nand U29014 (N_29014,N_28524,N_28762);
nor U29015 (N_29015,N_28595,N_28687);
nor U29016 (N_29016,N_28656,N_28676);
nand U29017 (N_29017,N_28748,N_28751);
nand U29018 (N_29018,N_28607,N_28529);
nand U29019 (N_29019,N_28598,N_28680);
nand U29020 (N_29020,N_28677,N_28697);
xor U29021 (N_29021,N_28678,N_28723);
nor U29022 (N_29022,N_28723,N_28625);
nor U29023 (N_29023,N_28699,N_28605);
nand U29024 (N_29024,N_28526,N_28507);
and U29025 (N_29025,N_28646,N_28565);
or U29026 (N_29026,N_28512,N_28567);
xor U29027 (N_29027,N_28779,N_28719);
nand U29028 (N_29028,N_28501,N_28547);
and U29029 (N_29029,N_28571,N_28771);
nor U29030 (N_29030,N_28652,N_28640);
and U29031 (N_29031,N_28714,N_28559);
xnor U29032 (N_29032,N_28703,N_28694);
and U29033 (N_29033,N_28623,N_28687);
xor U29034 (N_29034,N_28608,N_28667);
or U29035 (N_29035,N_28574,N_28649);
and U29036 (N_29036,N_28590,N_28793);
nor U29037 (N_29037,N_28596,N_28560);
nor U29038 (N_29038,N_28770,N_28535);
and U29039 (N_29039,N_28668,N_28765);
or U29040 (N_29040,N_28699,N_28592);
nand U29041 (N_29041,N_28585,N_28709);
nand U29042 (N_29042,N_28726,N_28554);
and U29043 (N_29043,N_28779,N_28700);
or U29044 (N_29044,N_28553,N_28508);
nor U29045 (N_29045,N_28624,N_28591);
nor U29046 (N_29046,N_28693,N_28658);
xnor U29047 (N_29047,N_28664,N_28516);
nand U29048 (N_29048,N_28558,N_28687);
or U29049 (N_29049,N_28637,N_28588);
or U29050 (N_29050,N_28758,N_28677);
and U29051 (N_29051,N_28636,N_28774);
or U29052 (N_29052,N_28608,N_28757);
nor U29053 (N_29053,N_28592,N_28796);
or U29054 (N_29054,N_28509,N_28636);
or U29055 (N_29055,N_28651,N_28551);
xor U29056 (N_29056,N_28647,N_28715);
nor U29057 (N_29057,N_28612,N_28670);
xor U29058 (N_29058,N_28793,N_28545);
nand U29059 (N_29059,N_28700,N_28544);
nand U29060 (N_29060,N_28641,N_28544);
and U29061 (N_29061,N_28633,N_28781);
nand U29062 (N_29062,N_28584,N_28727);
and U29063 (N_29063,N_28685,N_28590);
nand U29064 (N_29064,N_28773,N_28646);
and U29065 (N_29065,N_28636,N_28571);
xnor U29066 (N_29066,N_28650,N_28543);
nor U29067 (N_29067,N_28581,N_28593);
nand U29068 (N_29068,N_28589,N_28713);
xor U29069 (N_29069,N_28571,N_28684);
nor U29070 (N_29070,N_28778,N_28515);
nand U29071 (N_29071,N_28655,N_28578);
and U29072 (N_29072,N_28680,N_28545);
or U29073 (N_29073,N_28709,N_28656);
and U29074 (N_29074,N_28627,N_28687);
xor U29075 (N_29075,N_28581,N_28753);
nand U29076 (N_29076,N_28688,N_28547);
xnor U29077 (N_29077,N_28738,N_28662);
and U29078 (N_29078,N_28536,N_28697);
xor U29079 (N_29079,N_28555,N_28580);
or U29080 (N_29080,N_28735,N_28690);
nor U29081 (N_29081,N_28615,N_28593);
and U29082 (N_29082,N_28734,N_28547);
nor U29083 (N_29083,N_28797,N_28728);
nor U29084 (N_29084,N_28741,N_28531);
and U29085 (N_29085,N_28750,N_28770);
nand U29086 (N_29086,N_28701,N_28673);
nor U29087 (N_29087,N_28606,N_28712);
and U29088 (N_29088,N_28701,N_28580);
nand U29089 (N_29089,N_28752,N_28726);
nand U29090 (N_29090,N_28723,N_28500);
nor U29091 (N_29091,N_28622,N_28714);
and U29092 (N_29092,N_28739,N_28577);
nor U29093 (N_29093,N_28605,N_28781);
nor U29094 (N_29094,N_28658,N_28777);
and U29095 (N_29095,N_28787,N_28761);
nor U29096 (N_29096,N_28771,N_28582);
and U29097 (N_29097,N_28542,N_28613);
xnor U29098 (N_29098,N_28703,N_28786);
xnor U29099 (N_29099,N_28767,N_28656);
nand U29100 (N_29100,N_28996,N_28892);
nand U29101 (N_29101,N_28991,N_29035);
nor U29102 (N_29102,N_28984,N_29089);
nand U29103 (N_29103,N_28854,N_28955);
nand U29104 (N_29104,N_28810,N_28868);
and U29105 (N_29105,N_29097,N_29002);
nand U29106 (N_29106,N_28914,N_28869);
xor U29107 (N_29107,N_28846,N_28830);
and U29108 (N_29108,N_29047,N_28938);
nor U29109 (N_29109,N_28989,N_29099);
nand U29110 (N_29110,N_28814,N_28884);
or U29111 (N_29111,N_28905,N_28806);
and U29112 (N_29112,N_29007,N_29005);
xor U29113 (N_29113,N_28852,N_29092);
xor U29114 (N_29114,N_29080,N_28800);
nor U29115 (N_29115,N_29043,N_29029);
nand U29116 (N_29116,N_28944,N_28873);
nand U29117 (N_29117,N_28900,N_28923);
or U29118 (N_29118,N_28913,N_28987);
xor U29119 (N_29119,N_28818,N_28986);
nand U29120 (N_29120,N_28804,N_28942);
or U29121 (N_29121,N_29028,N_28811);
and U29122 (N_29122,N_28994,N_29074);
nor U29123 (N_29123,N_28917,N_28920);
xnor U29124 (N_29124,N_29059,N_29051);
or U29125 (N_29125,N_28916,N_28912);
xnor U29126 (N_29126,N_28896,N_29086);
xnor U29127 (N_29127,N_28845,N_29065);
nand U29128 (N_29128,N_28928,N_28969);
and U29129 (N_29129,N_28995,N_28894);
nor U29130 (N_29130,N_28973,N_28890);
nand U29131 (N_29131,N_29090,N_28831);
and U29132 (N_29132,N_28824,N_28895);
nand U29133 (N_29133,N_28897,N_28977);
or U29134 (N_29134,N_28817,N_29071);
nor U29135 (N_29135,N_28957,N_29046);
nor U29136 (N_29136,N_28975,N_28813);
nand U29137 (N_29137,N_29067,N_28870);
and U29138 (N_29138,N_28933,N_29095);
and U29139 (N_29139,N_28820,N_28825);
and U29140 (N_29140,N_28945,N_28891);
and U29141 (N_29141,N_28956,N_28835);
xor U29142 (N_29142,N_29098,N_29024);
or U29143 (N_29143,N_28823,N_29030);
or U29144 (N_29144,N_28812,N_28861);
xnor U29145 (N_29145,N_28860,N_29032);
xor U29146 (N_29146,N_29066,N_29023);
nor U29147 (N_29147,N_29026,N_29083);
xor U29148 (N_29148,N_28941,N_29039);
nor U29149 (N_29149,N_29048,N_29041);
nand U29150 (N_29150,N_28841,N_28947);
nor U29151 (N_29151,N_29060,N_29020);
nor U29152 (N_29152,N_29064,N_28932);
or U29153 (N_29153,N_29079,N_28871);
nor U29154 (N_29154,N_28815,N_28961);
or U29155 (N_29155,N_29091,N_29003);
or U29156 (N_29156,N_28836,N_28828);
nor U29157 (N_29157,N_28930,N_28901);
nand U29158 (N_29158,N_28856,N_28959);
nand U29159 (N_29159,N_29000,N_28963);
nand U29160 (N_29160,N_28908,N_28968);
nor U29161 (N_29161,N_28940,N_28954);
or U29162 (N_29162,N_28918,N_29085);
and U29163 (N_29163,N_28862,N_28998);
and U29164 (N_29164,N_28885,N_28888);
xnor U29165 (N_29165,N_29053,N_28922);
nand U29166 (N_29166,N_28878,N_28889);
nor U29167 (N_29167,N_28910,N_29025);
xor U29168 (N_29168,N_29054,N_28863);
nand U29169 (N_29169,N_29037,N_28872);
and U29170 (N_29170,N_29042,N_28834);
or U29171 (N_29171,N_29050,N_28801);
nand U29172 (N_29172,N_29081,N_28883);
and U29173 (N_29173,N_29088,N_28906);
and U29174 (N_29174,N_28958,N_28988);
or U29175 (N_29175,N_28921,N_29008);
and U29176 (N_29176,N_28967,N_28924);
or U29177 (N_29177,N_29006,N_28832);
xnor U29178 (N_29178,N_28847,N_29082);
and U29179 (N_29179,N_28886,N_28807);
nor U29180 (N_29180,N_29063,N_28972);
xor U29181 (N_29181,N_28898,N_28950);
and U29182 (N_29182,N_28899,N_29013);
nor U29183 (N_29183,N_28966,N_28939);
xor U29184 (N_29184,N_29070,N_28937);
or U29185 (N_29185,N_29058,N_28960);
nor U29186 (N_29186,N_29068,N_28849);
and U29187 (N_29187,N_29077,N_28964);
nor U29188 (N_29188,N_28844,N_28843);
and U29189 (N_29189,N_28934,N_28833);
nand U29190 (N_29190,N_28880,N_28903);
nor U29191 (N_29191,N_28982,N_29044);
or U29192 (N_29192,N_28865,N_28993);
or U29193 (N_29193,N_29014,N_28949);
nor U29194 (N_29194,N_29078,N_28827);
nor U29195 (N_29195,N_28946,N_28826);
or U29196 (N_29196,N_28858,N_28948);
xnor U29197 (N_29197,N_29004,N_28990);
nand U29198 (N_29198,N_28879,N_29016);
or U29199 (N_29199,N_28971,N_28840);
or U29200 (N_29200,N_28819,N_28866);
and U29201 (N_29201,N_29075,N_29045);
or U29202 (N_29202,N_28848,N_28882);
or U29203 (N_29203,N_29049,N_28911);
and U29204 (N_29204,N_28936,N_29052);
nor U29205 (N_29205,N_29022,N_29033);
and U29206 (N_29206,N_29073,N_29057);
nand U29207 (N_29207,N_28929,N_28915);
or U29208 (N_29208,N_29015,N_29021);
or U29209 (N_29209,N_29018,N_29062);
nand U29210 (N_29210,N_28805,N_28875);
or U29211 (N_29211,N_28821,N_29093);
or U29212 (N_29212,N_28859,N_29001);
or U29213 (N_29213,N_29061,N_29087);
xor U29214 (N_29214,N_28851,N_28978);
xnor U29215 (N_29215,N_28808,N_29072);
or U29216 (N_29216,N_28867,N_28926);
xor U29217 (N_29217,N_29076,N_29096);
and U29218 (N_29218,N_28802,N_28887);
nor U29219 (N_29219,N_28980,N_29012);
or U29220 (N_29220,N_28902,N_28953);
and U29221 (N_29221,N_29036,N_29056);
and U29222 (N_29222,N_29009,N_28907);
nor U29223 (N_29223,N_28809,N_29019);
nor U29224 (N_29224,N_28838,N_29034);
nand U29225 (N_29225,N_29094,N_28857);
xnor U29226 (N_29226,N_28974,N_29040);
nand U29227 (N_29227,N_29017,N_28850);
xor U29228 (N_29228,N_29011,N_28837);
and U29229 (N_29229,N_28952,N_28904);
xor U29230 (N_29230,N_29027,N_29069);
or U29231 (N_29231,N_28962,N_28985);
and U29232 (N_29232,N_28829,N_28803);
xnor U29233 (N_29233,N_28842,N_29055);
nor U29234 (N_29234,N_28927,N_28925);
nand U29235 (N_29235,N_28981,N_28822);
or U29236 (N_29236,N_28951,N_28997);
xor U29237 (N_29237,N_28979,N_29038);
nand U29238 (N_29238,N_28855,N_28816);
xor U29239 (N_29239,N_29010,N_28999);
or U29240 (N_29240,N_28864,N_28943);
nand U29241 (N_29241,N_28893,N_28919);
nor U29242 (N_29242,N_29084,N_28909);
nand U29243 (N_29243,N_29031,N_28839);
and U29244 (N_29244,N_28992,N_28935);
nor U29245 (N_29245,N_28874,N_28965);
nand U29246 (N_29246,N_28976,N_28877);
nand U29247 (N_29247,N_28970,N_28931);
xor U29248 (N_29248,N_28853,N_28876);
nand U29249 (N_29249,N_28983,N_28881);
nand U29250 (N_29250,N_28854,N_28866);
nor U29251 (N_29251,N_29012,N_28969);
xnor U29252 (N_29252,N_28902,N_28806);
xnor U29253 (N_29253,N_28882,N_28883);
nand U29254 (N_29254,N_28965,N_28820);
xor U29255 (N_29255,N_29070,N_28802);
and U29256 (N_29256,N_28873,N_28953);
and U29257 (N_29257,N_28884,N_29028);
xor U29258 (N_29258,N_28909,N_28943);
xor U29259 (N_29259,N_29079,N_29073);
and U29260 (N_29260,N_29065,N_29026);
nor U29261 (N_29261,N_29082,N_28995);
nor U29262 (N_29262,N_29011,N_28839);
nor U29263 (N_29263,N_28836,N_28928);
and U29264 (N_29264,N_28956,N_29002);
xnor U29265 (N_29265,N_28944,N_28948);
xor U29266 (N_29266,N_28886,N_28922);
and U29267 (N_29267,N_28857,N_28921);
and U29268 (N_29268,N_28973,N_29034);
or U29269 (N_29269,N_28810,N_28981);
nand U29270 (N_29270,N_29003,N_28971);
nor U29271 (N_29271,N_29030,N_28931);
and U29272 (N_29272,N_28992,N_28993);
and U29273 (N_29273,N_28827,N_29093);
nor U29274 (N_29274,N_28896,N_28851);
and U29275 (N_29275,N_29061,N_29029);
nand U29276 (N_29276,N_28846,N_28955);
or U29277 (N_29277,N_28960,N_28911);
xnor U29278 (N_29278,N_29036,N_28960);
nand U29279 (N_29279,N_29010,N_28930);
xnor U29280 (N_29280,N_28993,N_28818);
xor U29281 (N_29281,N_28929,N_29051);
nand U29282 (N_29282,N_28872,N_29024);
and U29283 (N_29283,N_28916,N_28896);
nand U29284 (N_29284,N_28912,N_29072);
nand U29285 (N_29285,N_29006,N_28963);
or U29286 (N_29286,N_28887,N_29086);
and U29287 (N_29287,N_28906,N_28922);
nor U29288 (N_29288,N_29095,N_28877);
nor U29289 (N_29289,N_28837,N_28811);
nor U29290 (N_29290,N_28896,N_29077);
xor U29291 (N_29291,N_28846,N_28967);
and U29292 (N_29292,N_28922,N_28997);
nand U29293 (N_29293,N_28839,N_29033);
xor U29294 (N_29294,N_29018,N_28871);
xor U29295 (N_29295,N_28972,N_28979);
or U29296 (N_29296,N_28923,N_28918);
nand U29297 (N_29297,N_29017,N_29037);
nand U29298 (N_29298,N_28899,N_28904);
or U29299 (N_29299,N_28953,N_28977);
xor U29300 (N_29300,N_28827,N_28948);
nor U29301 (N_29301,N_28925,N_28864);
xor U29302 (N_29302,N_28915,N_28966);
xor U29303 (N_29303,N_28918,N_28812);
xnor U29304 (N_29304,N_29015,N_28818);
nor U29305 (N_29305,N_29081,N_28807);
xnor U29306 (N_29306,N_28922,N_28968);
nor U29307 (N_29307,N_28992,N_29020);
xor U29308 (N_29308,N_29021,N_28941);
xor U29309 (N_29309,N_28867,N_29054);
xnor U29310 (N_29310,N_29031,N_28873);
or U29311 (N_29311,N_28847,N_29062);
nand U29312 (N_29312,N_29020,N_28964);
nand U29313 (N_29313,N_29079,N_28926);
nand U29314 (N_29314,N_28956,N_28985);
nor U29315 (N_29315,N_28931,N_29026);
and U29316 (N_29316,N_28825,N_28905);
and U29317 (N_29317,N_28986,N_28927);
or U29318 (N_29318,N_28968,N_28986);
xnor U29319 (N_29319,N_28863,N_28972);
nor U29320 (N_29320,N_28874,N_28993);
nand U29321 (N_29321,N_29017,N_28960);
xnor U29322 (N_29322,N_29043,N_29096);
or U29323 (N_29323,N_28848,N_29073);
xnor U29324 (N_29324,N_28822,N_28813);
or U29325 (N_29325,N_29063,N_28854);
xor U29326 (N_29326,N_28950,N_28871);
and U29327 (N_29327,N_28855,N_29080);
xor U29328 (N_29328,N_28937,N_28996);
and U29329 (N_29329,N_28827,N_28864);
and U29330 (N_29330,N_28801,N_29001);
or U29331 (N_29331,N_29087,N_28999);
or U29332 (N_29332,N_29000,N_28973);
or U29333 (N_29333,N_28974,N_28847);
and U29334 (N_29334,N_29032,N_28880);
nor U29335 (N_29335,N_28806,N_29057);
or U29336 (N_29336,N_28964,N_29007);
nor U29337 (N_29337,N_28807,N_28814);
or U29338 (N_29338,N_28888,N_28900);
xor U29339 (N_29339,N_28965,N_28967);
and U29340 (N_29340,N_29091,N_28921);
nand U29341 (N_29341,N_28876,N_29005);
and U29342 (N_29342,N_28967,N_28857);
or U29343 (N_29343,N_28921,N_28987);
nor U29344 (N_29344,N_29028,N_28937);
nand U29345 (N_29345,N_28950,N_28899);
and U29346 (N_29346,N_29081,N_28952);
xnor U29347 (N_29347,N_29089,N_29062);
and U29348 (N_29348,N_29028,N_28959);
nor U29349 (N_29349,N_28913,N_29083);
nand U29350 (N_29350,N_29016,N_29093);
xor U29351 (N_29351,N_28929,N_28808);
or U29352 (N_29352,N_28862,N_28873);
nand U29353 (N_29353,N_28936,N_28958);
xnor U29354 (N_29354,N_29007,N_28913);
or U29355 (N_29355,N_29062,N_29039);
nand U29356 (N_29356,N_29040,N_29060);
and U29357 (N_29357,N_29089,N_28928);
nor U29358 (N_29358,N_29049,N_29056);
and U29359 (N_29359,N_29012,N_29001);
or U29360 (N_29360,N_28976,N_29092);
and U29361 (N_29361,N_29078,N_28832);
nand U29362 (N_29362,N_28951,N_29029);
or U29363 (N_29363,N_28884,N_29011);
nor U29364 (N_29364,N_28959,N_28931);
xor U29365 (N_29365,N_28957,N_28985);
and U29366 (N_29366,N_28924,N_28833);
nor U29367 (N_29367,N_29088,N_29016);
nand U29368 (N_29368,N_28803,N_28910);
xor U29369 (N_29369,N_29055,N_29066);
or U29370 (N_29370,N_28999,N_28997);
xor U29371 (N_29371,N_29069,N_28982);
xnor U29372 (N_29372,N_28955,N_28962);
nor U29373 (N_29373,N_28956,N_28994);
and U29374 (N_29374,N_28801,N_29008);
nand U29375 (N_29375,N_28936,N_29036);
or U29376 (N_29376,N_28835,N_28961);
xor U29377 (N_29377,N_28895,N_29040);
nand U29378 (N_29378,N_28983,N_28960);
and U29379 (N_29379,N_28906,N_28813);
nand U29380 (N_29380,N_29067,N_29030);
nor U29381 (N_29381,N_29081,N_28864);
and U29382 (N_29382,N_28879,N_28967);
xor U29383 (N_29383,N_28813,N_28826);
nor U29384 (N_29384,N_28823,N_28906);
xor U29385 (N_29385,N_28984,N_29096);
xnor U29386 (N_29386,N_28827,N_28973);
or U29387 (N_29387,N_28818,N_28814);
nor U29388 (N_29388,N_28849,N_28997);
or U29389 (N_29389,N_28877,N_29091);
and U29390 (N_29390,N_28943,N_28982);
nor U29391 (N_29391,N_29059,N_29006);
xor U29392 (N_29392,N_29055,N_29049);
nor U29393 (N_29393,N_28824,N_28811);
xnor U29394 (N_29394,N_29018,N_28998);
or U29395 (N_29395,N_29026,N_29080);
and U29396 (N_29396,N_28874,N_29070);
or U29397 (N_29397,N_28862,N_28955);
xnor U29398 (N_29398,N_29067,N_28934);
or U29399 (N_29399,N_28880,N_29072);
and U29400 (N_29400,N_29249,N_29103);
and U29401 (N_29401,N_29229,N_29284);
nand U29402 (N_29402,N_29164,N_29319);
nor U29403 (N_29403,N_29297,N_29379);
and U29404 (N_29404,N_29124,N_29341);
xnor U29405 (N_29405,N_29174,N_29367);
xnor U29406 (N_29406,N_29226,N_29377);
nor U29407 (N_29407,N_29157,N_29102);
nand U29408 (N_29408,N_29293,N_29294);
and U29409 (N_29409,N_29242,N_29209);
or U29410 (N_29410,N_29150,N_29220);
and U29411 (N_29411,N_29354,N_29146);
nand U29412 (N_29412,N_29210,N_29136);
xnor U29413 (N_29413,N_29222,N_29274);
xnor U29414 (N_29414,N_29173,N_29251);
nand U29415 (N_29415,N_29259,N_29148);
nor U29416 (N_29416,N_29121,N_29374);
and U29417 (N_29417,N_29171,N_29214);
nand U29418 (N_29418,N_29200,N_29307);
xnor U29419 (N_29419,N_29328,N_29218);
nor U29420 (N_29420,N_29140,N_29114);
nand U29421 (N_29421,N_29277,N_29276);
and U29422 (N_29422,N_29394,N_29355);
nor U29423 (N_29423,N_29370,N_29378);
or U29424 (N_29424,N_29193,N_29390);
and U29425 (N_29425,N_29356,N_29175);
or U29426 (N_29426,N_29368,N_29237);
nor U29427 (N_29427,N_29324,N_29330);
nor U29428 (N_29428,N_29278,N_29396);
and U29429 (N_29429,N_29326,N_29160);
nor U29430 (N_29430,N_29117,N_29199);
nand U29431 (N_29431,N_29194,N_29399);
and U29432 (N_29432,N_29298,N_29190);
nor U29433 (N_29433,N_29316,N_29185);
and U29434 (N_29434,N_29296,N_29305);
xnor U29435 (N_29435,N_29167,N_29187);
or U29436 (N_29436,N_29139,N_29219);
nor U29437 (N_29437,N_29228,N_29303);
or U29438 (N_29438,N_29299,N_29270);
xnor U29439 (N_29439,N_29147,N_29292);
xor U29440 (N_29440,N_29338,N_29262);
nand U29441 (N_29441,N_29142,N_29295);
nor U29442 (N_29442,N_29353,N_29323);
and U29443 (N_29443,N_29230,N_29216);
xnor U29444 (N_29444,N_29310,N_29149);
or U29445 (N_29445,N_29331,N_29119);
and U29446 (N_29446,N_29311,N_29345);
nand U29447 (N_29447,N_29232,N_29375);
or U29448 (N_29448,N_29246,N_29360);
xnor U29449 (N_29449,N_29285,N_29108);
nor U29450 (N_29450,N_29280,N_29327);
xor U29451 (N_29451,N_29332,N_29196);
nand U29452 (N_29452,N_29176,N_29234);
xor U29453 (N_29453,N_29395,N_29301);
and U29454 (N_29454,N_29155,N_29129);
nand U29455 (N_29455,N_29256,N_29227);
and U29456 (N_29456,N_29236,N_29380);
nor U29457 (N_29457,N_29239,N_29302);
and U29458 (N_29458,N_29221,N_29392);
xnor U29459 (N_29459,N_29289,N_29349);
nand U29460 (N_29460,N_29244,N_29267);
nand U29461 (N_29461,N_29318,N_29189);
xor U29462 (N_29462,N_29115,N_29342);
nand U29463 (N_29463,N_29208,N_29329);
and U29464 (N_29464,N_29233,N_29126);
and U29465 (N_29465,N_29195,N_29120);
nand U29466 (N_29466,N_29260,N_29335);
or U29467 (N_29467,N_29381,N_29321);
xnor U29468 (N_29468,N_29385,N_29373);
nand U29469 (N_29469,N_29104,N_29206);
nor U29470 (N_29470,N_29290,N_29144);
and U29471 (N_29471,N_29398,N_29231);
nor U29472 (N_29472,N_29275,N_29107);
nor U29473 (N_29473,N_29204,N_29281);
or U29474 (N_29474,N_29145,N_29106);
or U29475 (N_29475,N_29391,N_29192);
nand U29476 (N_29476,N_29158,N_29138);
nand U29477 (N_29477,N_29132,N_29170);
xnor U29478 (N_29478,N_29271,N_29197);
and U29479 (N_29479,N_29178,N_29263);
or U29480 (N_29480,N_29334,N_29201);
and U29481 (N_29481,N_29252,N_29151);
nor U29482 (N_29482,N_29291,N_29112);
nor U29483 (N_29483,N_29163,N_29363);
xnor U29484 (N_29484,N_29369,N_29172);
or U29485 (N_29485,N_29388,N_29122);
nand U29486 (N_29486,N_29168,N_29340);
and U29487 (N_29487,N_29205,N_29336);
nand U29488 (N_29488,N_29165,N_29133);
nand U29489 (N_29489,N_29339,N_29154);
and U29490 (N_29490,N_29109,N_29350);
nand U29491 (N_29491,N_29382,N_29179);
xor U29492 (N_29492,N_29287,N_29243);
or U29493 (N_29493,N_29347,N_29153);
nor U29494 (N_29494,N_29372,N_29143);
nor U29495 (N_29495,N_29105,N_29257);
and U29496 (N_29496,N_29288,N_29362);
xor U29497 (N_29497,N_29241,N_29300);
nor U29498 (N_29498,N_29180,N_29358);
and U29499 (N_29499,N_29183,N_29212);
nor U29500 (N_29500,N_29337,N_29266);
or U29501 (N_29501,N_29207,N_29203);
and U29502 (N_29502,N_29186,N_29286);
nor U29503 (N_29503,N_29134,N_29255);
nor U29504 (N_29504,N_29188,N_29113);
nand U29505 (N_29505,N_29211,N_29304);
xor U29506 (N_29506,N_29137,N_29156);
or U29507 (N_29507,N_29261,N_29346);
and U29508 (N_29508,N_29128,N_29215);
nand U29509 (N_29509,N_29343,N_29235);
nand U29510 (N_29510,N_29265,N_29269);
nand U29511 (N_29511,N_29127,N_29344);
and U29512 (N_29512,N_29159,N_29166);
xnor U29513 (N_29513,N_29125,N_29162);
nand U29514 (N_29514,N_29359,N_29313);
nor U29515 (N_29515,N_29245,N_29223);
nor U29516 (N_29516,N_29364,N_29169);
xor U29517 (N_29517,N_29312,N_29315);
nand U29518 (N_29518,N_29135,N_29238);
nor U29519 (N_29519,N_29308,N_29202);
nand U29520 (N_29520,N_29250,N_29365);
nor U29521 (N_29521,N_29309,N_29272);
nand U29522 (N_29522,N_29333,N_29282);
and U29523 (N_29523,N_29387,N_29352);
nor U29524 (N_29524,N_29264,N_29198);
and U29525 (N_29525,N_29357,N_29225);
nor U29526 (N_29526,N_29177,N_29123);
and U29527 (N_29527,N_29268,N_29181);
xor U29528 (N_29528,N_29376,N_29254);
and U29529 (N_29529,N_29116,N_29111);
xnor U29530 (N_29530,N_29306,N_29182);
and U29531 (N_29531,N_29389,N_29161);
or U29532 (N_29532,N_29118,N_29351);
and U29533 (N_29533,N_29283,N_29361);
or U29534 (N_29534,N_29253,N_29184);
nand U29535 (N_29535,N_29213,N_29371);
or U29536 (N_29536,N_29141,N_29397);
and U29537 (N_29537,N_29240,N_29322);
nand U29538 (N_29538,N_29131,N_29110);
nor U29539 (N_29539,N_29100,N_29224);
nand U29540 (N_29540,N_29386,N_29314);
or U29541 (N_29541,N_29101,N_29393);
xor U29542 (N_29542,N_29348,N_29130);
and U29543 (N_29543,N_29317,N_29384);
nor U29544 (N_29544,N_29383,N_29366);
nor U29545 (N_29545,N_29258,N_29248);
nand U29546 (N_29546,N_29325,N_29152);
nand U29547 (N_29547,N_29191,N_29320);
xor U29548 (N_29548,N_29217,N_29247);
nand U29549 (N_29549,N_29273,N_29279);
nor U29550 (N_29550,N_29384,N_29378);
and U29551 (N_29551,N_29280,N_29129);
or U29552 (N_29552,N_29332,N_29146);
xnor U29553 (N_29553,N_29262,N_29203);
nor U29554 (N_29554,N_29191,N_29354);
xnor U29555 (N_29555,N_29376,N_29366);
xor U29556 (N_29556,N_29130,N_29194);
and U29557 (N_29557,N_29271,N_29340);
xnor U29558 (N_29558,N_29295,N_29151);
and U29559 (N_29559,N_29142,N_29173);
nor U29560 (N_29560,N_29150,N_29107);
and U29561 (N_29561,N_29352,N_29310);
xnor U29562 (N_29562,N_29345,N_29117);
nor U29563 (N_29563,N_29370,N_29137);
nor U29564 (N_29564,N_29143,N_29398);
nand U29565 (N_29565,N_29282,N_29265);
nor U29566 (N_29566,N_29108,N_29364);
nor U29567 (N_29567,N_29114,N_29326);
or U29568 (N_29568,N_29191,N_29182);
or U29569 (N_29569,N_29210,N_29178);
xor U29570 (N_29570,N_29199,N_29193);
and U29571 (N_29571,N_29141,N_29235);
or U29572 (N_29572,N_29118,N_29183);
nor U29573 (N_29573,N_29229,N_29142);
xor U29574 (N_29574,N_29349,N_29303);
and U29575 (N_29575,N_29142,N_29393);
and U29576 (N_29576,N_29275,N_29349);
nor U29577 (N_29577,N_29216,N_29189);
or U29578 (N_29578,N_29284,N_29385);
nand U29579 (N_29579,N_29105,N_29129);
nand U29580 (N_29580,N_29119,N_29250);
nor U29581 (N_29581,N_29138,N_29317);
nand U29582 (N_29582,N_29344,N_29330);
nor U29583 (N_29583,N_29111,N_29160);
and U29584 (N_29584,N_29360,N_29318);
nand U29585 (N_29585,N_29283,N_29370);
and U29586 (N_29586,N_29165,N_29350);
nand U29587 (N_29587,N_29281,N_29380);
or U29588 (N_29588,N_29331,N_29343);
or U29589 (N_29589,N_29141,N_29132);
nand U29590 (N_29590,N_29283,N_29207);
or U29591 (N_29591,N_29184,N_29241);
or U29592 (N_29592,N_29321,N_29233);
nor U29593 (N_29593,N_29305,N_29192);
xnor U29594 (N_29594,N_29161,N_29125);
or U29595 (N_29595,N_29293,N_29103);
or U29596 (N_29596,N_29205,N_29373);
or U29597 (N_29597,N_29252,N_29270);
or U29598 (N_29598,N_29217,N_29198);
nand U29599 (N_29599,N_29340,N_29230);
xnor U29600 (N_29600,N_29187,N_29154);
xor U29601 (N_29601,N_29136,N_29327);
nand U29602 (N_29602,N_29314,N_29227);
nand U29603 (N_29603,N_29146,N_29288);
nor U29604 (N_29604,N_29379,N_29326);
nor U29605 (N_29605,N_29377,N_29358);
or U29606 (N_29606,N_29353,N_29225);
nor U29607 (N_29607,N_29320,N_29157);
and U29608 (N_29608,N_29270,N_29102);
or U29609 (N_29609,N_29369,N_29384);
nor U29610 (N_29610,N_29254,N_29272);
and U29611 (N_29611,N_29302,N_29147);
or U29612 (N_29612,N_29218,N_29371);
xor U29613 (N_29613,N_29244,N_29309);
xnor U29614 (N_29614,N_29243,N_29178);
nor U29615 (N_29615,N_29128,N_29380);
xor U29616 (N_29616,N_29386,N_29100);
nand U29617 (N_29617,N_29141,N_29319);
or U29618 (N_29618,N_29268,N_29240);
nand U29619 (N_29619,N_29156,N_29218);
and U29620 (N_29620,N_29269,N_29394);
xnor U29621 (N_29621,N_29304,N_29161);
nor U29622 (N_29622,N_29212,N_29364);
xor U29623 (N_29623,N_29310,N_29137);
nand U29624 (N_29624,N_29215,N_29220);
xnor U29625 (N_29625,N_29347,N_29157);
and U29626 (N_29626,N_29101,N_29371);
nor U29627 (N_29627,N_29105,N_29240);
xor U29628 (N_29628,N_29213,N_29211);
nand U29629 (N_29629,N_29330,N_29302);
and U29630 (N_29630,N_29293,N_29399);
nor U29631 (N_29631,N_29130,N_29260);
nor U29632 (N_29632,N_29237,N_29375);
nand U29633 (N_29633,N_29188,N_29232);
or U29634 (N_29634,N_29194,N_29157);
and U29635 (N_29635,N_29129,N_29206);
nand U29636 (N_29636,N_29379,N_29303);
nand U29637 (N_29637,N_29173,N_29383);
or U29638 (N_29638,N_29354,N_29147);
xnor U29639 (N_29639,N_29189,N_29304);
nand U29640 (N_29640,N_29136,N_29398);
nand U29641 (N_29641,N_29146,N_29106);
or U29642 (N_29642,N_29153,N_29156);
nand U29643 (N_29643,N_29206,N_29145);
and U29644 (N_29644,N_29329,N_29346);
nand U29645 (N_29645,N_29386,N_29211);
or U29646 (N_29646,N_29191,N_29390);
nor U29647 (N_29647,N_29275,N_29202);
xnor U29648 (N_29648,N_29314,N_29383);
nor U29649 (N_29649,N_29163,N_29196);
xnor U29650 (N_29650,N_29104,N_29145);
nor U29651 (N_29651,N_29125,N_29114);
or U29652 (N_29652,N_29208,N_29149);
or U29653 (N_29653,N_29320,N_29259);
xnor U29654 (N_29654,N_29391,N_29213);
and U29655 (N_29655,N_29201,N_29395);
nand U29656 (N_29656,N_29350,N_29219);
and U29657 (N_29657,N_29285,N_29231);
and U29658 (N_29658,N_29123,N_29200);
xor U29659 (N_29659,N_29323,N_29127);
xnor U29660 (N_29660,N_29364,N_29159);
or U29661 (N_29661,N_29175,N_29355);
or U29662 (N_29662,N_29208,N_29377);
or U29663 (N_29663,N_29271,N_29390);
and U29664 (N_29664,N_29322,N_29145);
nand U29665 (N_29665,N_29146,N_29230);
xor U29666 (N_29666,N_29332,N_29299);
and U29667 (N_29667,N_29313,N_29379);
and U29668 (N_29668,N_29122,N_29257);
nor U29669 (N_29669,N_29131,N_29359);
and U29670 (N_29670,N_29398,N_29317);
nor U29671 (N_29671,N_29203,N_29122);
xnor U29672 (N_29672,N_29285,N_29194);
nor U29673 (N_29673,N_29145,N_29164);
nand U29674 (N_29674,N_29244,N_29206);
nor U29675 (N_29675,N_29226,N_29341);
xor U29676 (N_29676,N_29316,N_29323);
xor U29677 (N_29677,N_29250,N_29381);
and U29678 (N_29678,N_29204,N_29383);
and U29679 (N_29679,N_29143,N_29278);
nand U29680 (N_29680,N_29170,N_29247);
xnor U29681 (N_29681,N_29166,N_29277);
or U29682 (N_29682,N_29272,N_29386);
nor U29683 (N_29683,N_29382,N_29210);
nand U29684 (N_29684,N_29329,N_29152);
or U29685 (N_29685,N_29126,N_29196);
or U29686 (N_29686,N_29285,N_29178);
nor U29687 (N_29687,N_29249,N_29204);
and U29688 (N_29688,N_29241,N_29219);
xnor U29689 (N_29689,N_29291,N_29368);
and U29690 (N_29690,N_29151,N_29190);
nor U29691 (N_29691,N_29283,N_29296);
or U29692 (N_29692,N_29153,N_29184);
nand U29693 (N_29693,N_29175,N_29196);
and U29694 (N_29694,N_29299,N_29346);
and U29695 (N_29695,N_29318,N_29215);
xor U29696 (N_29696,N_29139,N_29281);
and U29697 (N_29697,N_29174,N_29381);
xor U29698 (N_29698,N_29175,N_29242);
or U29699 (N_29699,N_29284,N_29371);
xnor U29700 (N_29700,N_29585,N_29582);
nand U29701 (N_29701,N_29698,N_29647);
nand U29702 (N_29702,N_29689,N_29683);
and U29703 (N_29703,N_29478,N_29475);
nand U29704 (N_29704,N_29401,N_29587);
or U29705 (N_29705,N_29521,N_29574);
nand U29706 (N_29706,N_29464,N_29442);
nor U29707 (N_29707,N_29668,N_29631);
nand U29708 (N_29708,N_29640,N_29550);
nor U29709 (N_29709,N_29461,N_29581);
nor U29710 (N_29710,N_29694,N_29412);
nand U29711 (N_29711,N_29637,N_29458);
nand U29712 (N_29712,N_29416,N_29513);
nand U29713 (N_29713,N_29607,N_29674);
nor U29714 (N_29714,N_29570,N_29455);
nor U29715 (N_29715,N_29596,N_29646);
xor U29716 (N_29716,N_29453,N_29598);
nand U29717 (N_29717,N_29542,N_29434);
nand U29718 (N_29718,N_29402,N_29452);
and U29719 (N_29719,N_29456,N_29414);
and U29720 (N_29720,N_29451,N_29400);
or U29721 (N_29721,N_29500,N_29468);
xor U29722 (N_29722,N_29490,N_29693);
xor U29723 (N_29723,N_29463,N_29555);
and U29724 (N_29724,N_29527,N_29422);
and U29725 (N_29725,N_29409,N_29566);
nand U29726 (N_29726,N_29484,N_29404);
or U29727 (N_29727,N_29438,N_29526);
or U29728 (N_29728,N_29488,N_29466);
nor U29729 (N_29729,N_29630,N_29440);
nand U29730 (N_29730,N_29415,N_29473);
nor U29731 (N_29731,N_29548,N_29428);
or U29732 (N_29732,N_29532,N_29430);
nor U29733 (N_29733,N_29540,N_29608);
xnor U29734 (N_29734,N_29545,N_29684);
nor U29735 (N_29735,N_29667,N_29489);
nor U29736 (N_29736,N_29651,N_29445);
xor U29737 (N_29737,N_29588,N_29600);
nand U29738 (N_29738,N_29676,N_29612);
and U29739 (N_29739,N_29411,N_29539);
nor U29740 (N_29740,N_29580,N_29433);
nand U29741 (N_29741,N_29556,N_29613);
and U29742 (N_29742,N_29685,N_29663);
nand U29743 (N_29743,N_29517,N_29690);
and U29744 (N_29744,N_29454,N_29688);
xor U29745 (N_29745,N_29501,N_29657);
nand U29746 (N_29746,N_29655,N_29408);
and U29747 (N_29747,N_29460,N_29618);
or U29748 (N_29748,N_29692,N_29572);
xor U29749 (N_29749,N_29533,N_29495);
and U29750 (N_29750,N_29699,N_29506);
or U29751 (N_29751,N_29603,N_29601);
nor U29752 (N_29752,N_29591,N_29405);
or U29753 (N_29753,N_29465,N_29469);
and U29754 (N_29754,N_29424,N_29658);
xor U29755 (N_29755,N_29649,N_29546);
xor U29756 (N_29756,N_29622,N_29474);
nand U29757 (N_29757,N_29523,N_29642);
nand U29758 (N_29758,N_29579,N_29487);
nor U29759 (N_29759,N_29577,N_29459);
nor U29760 (N_29760,N_29560,N_29565);
nand U29761 (N_29761,N_29514,N_29530);
nor U29762 (N_29762,N_29639,N_29571);
and U29763 (N_29763,N_29511,N_29602);
xnor U29764 (N_29764,N_29564,N_29609);
nand U29765 (N_29765,N_29606,N_29595);
nor U29766 (N_29766,N_29615,N_29496);
or U29767 (N_29767,N_29691,N_29502);
and U29768 (N_29768,N_29576,N_29629);
and U29769 (N_29769,N_29450,N_29671);
or U29770 (N_29770,N_29632,N_29610);
or U29771 (N_29771,N_29436,N_29472);
nor U29772 (N_29772,N_29648,N_29432);
or U29773 (N_29773,N_29679,N_29420);
nand U29774 (N_29774,N_29439,N_29441);
or U29775 (N_29775,N_29696,N_29573);
or U29776 (N_29776,N_29482,N_29672);
or U29777 (N_29777,N_29578,N_29659);
nor U29778 (N_29778,N_29470,N_29423);
and U29779 (N_29779,N_29537,N_29522);
and U29780 (N_29780,N_29462,N_29593);
nand U29781 (N_29781,N_29551,N_29483);
nor U29782 (N_29782,N_29525,N_29619);
xor U29783 (N_29783,N_29457,N_29636);
and U29784 (N_29784,N_29589,N_29583);
nor U29785 (N_29785,N_29599,N_29427);
and U29786 (N_29786,N_29562,N_29625);
xor U29787 (N_29787,N_29549,N_29561);
and U29788 (N_29788,N_29635,N_29605);
and U29789 (N_29789,N_29481,N_29510);
xnor U29790 (N_29790,N_29505,N_29643);
or U29791 (N_29791,N_29611,N_29673);
nand U29792 (N_29792,N_29425,N_29553);
nand U29793 (N_29793,N_29681,N_29678);
xnor U29794 (N_29794,N_29638,N_29467);
xor U29795 (N_29795,N_29435,N_29528);
xnor U29796 (N_29796,N_29641,N_29654);
xor U29797 (N_29797,N_29644,N_29535);
nand U29798 (N_29798,N_29682,N_29507);
nor U29799 (N_29799,N_29558,N_29534);
xnor U29800 (N_29800,N_29443,N_29695);
or U29801 (N_29801,N_29634,N_29544);
and U29802 (N_29802,N_29406,N_29519);
nand U29803 (N_29803,N_29493,N_29697);
xnor U29804 (N_29804,N_29626,N_29418);
xor U29805 (N_29805,N_29686,N_29567);
and U29806 (N_29806,N_29499,N_29543);
and U29807 (N_29807,N_29413,N_29665);
nand U29808 (N_29808,N_29621,N_29666);
xor U29809 (N_29809,N_29431,N_29446);
nand U29810 (N_29810,N_29617,N_29590);
and U29811 (N_29811,N_29503,N_29531);
and U29812 (N_29812,N_29687,N_29476);
nor U29813 (N_29813,N_29492,N_29497);
and U29814 (N_29814,N_29614,N_29633);
and U29815 (N_29815,N_29437,N_29645);
or U29816 (N_29816,N_29515,N_29650);
or U29817 (N_29817,N_29444,N_29664);
or U29818 (N_29818,N_29557,N_29520);
nor U29819 (N_29819,N_29627,N_29559);
or U29820 (N_29820,N_29592,N_29677);
and U29821 (N_29821,N_29477,N_29449);
xor U29822 (N_29822,N_29547,N_29653);
xor U29823 (N_29823,N_29662,N_29675);
and U29824 (N_29824,N_29568,N_29623);
or U29825 (N_29825,N_29421,N_29670);
or U29826 (N_29826,N_29504,N_29604);
nand U29827 (N_29827,N_29586,N_29624);
xnor U29828 (N_29828,N_29575,N_29508);
nor U29829 (N_29829,N_29494,N_29518);
nor U29830 (N_29830,N_29538,N_29447);
or U29831 (N_29831,N_29616,N_29448);
xor U29832 (N_29832,N_29516,N_29524);
or U29833 (N_29833,N_29552,N_29480);
or U29834 (N_29834,N_29529,N_29569);
xnor U29835 (N_29835,N_29410,N_29536);
and U29836 (N_29836,N_29479,N_29563);
and U29837 (N_29837,N_29429,N_29419);
nand U29838 (N_29838,N_29417,N_29597);
nand U29839 (N_29839,N_29485,N_29661);
xnor U29840 (N_29840,N_29486,N_29407);
nor U29841 (N_29841,N_29403,N_29471);
or U29842 (N_29842,N_29426,N_29512);
nand U29843 (N_29843,N_29584,N_29509);
or U29844 (N_29844,N_29594,N_29554);
nor U29845 (N_29845,N_29660,N_29628);
xor U29846 (N_29846,N_29652,N_29541);
nand U29847 (N_29847,N_29669,N_29620);
nor U29848 (N_29848,N_29498,N_29491);
or U29849 (N_29849,N_29680,N_29656);
or U29850 (N_29850,N_29498,N_29514);
and U29851 (N_29851,N_29439,N_29510);
or U29852 (N_29852,N_29466,N_29661);
xnor U29853 (N_29853,N_29483,N_29562);
or U29854 (N_29854,N_29539,N_29533);
xnor U29855 (N_29855,N_29604,N_29567);
nand U29856 (N_29856,N_29579,N_29454);
nor U29857 (N_29857,N_29494,N_29603);
or U29858 (N_29858,N_29562,N_29621);
and U29859 (N_29859,N_29466,N_29411);
or U29860 (N_29860,N_29430,N_29572);
and U29861 (N_29861,N_29405,N_29574);
xor U29862 (N_29862,N_29585,N_29698);
or U29863 (N_29863,N_29603,N_29683);
and U29864 (N_29864,N_29683,N_29622);
xnor U29865 (N_29865,N_29547,N_29657);
xnor U29866 (N_29866,N_29621,N_29699);
xor U29867 (N_29867,N_29679,N_29669);
xnor U29868 (N_29868,N_29435,N_29561);
nand U29869 (N_29869,N_29629,N_29556);
nor U29870 (N_29870,N_29465,N_29553);
nand U29871 (N_29871,N_29603,N_29682);
and U29872 (N_29872,N_29429,N_29534);
and U29873 (N_29873,N_29591,N_29586);
nand U29874 (N_29874,N_29485,N_29663);
or U29875 (N_29875,N_29457,N_29455);
xor U29876 (N_29876,N_29416,N_29451);
nand U29877 (N_29877,N_29491,N_29591);
or U29878 (N_29878,N_29566,N_29689);
nor U29879 (N_29879,N_29630,N_29634);
xor U29880 (N_29880,N_29405,N_29443);
nor U29881 (N_29881,N_29600,N_29623);
and U29882 (N_29882,N_29489,N_29512);
xnor U29883 (N_29883,N_29695,N_29460);
or U29884 (N_29884,N_29680,N_29555);
nand U29885 (N_29885,N_29560,N_29672);
or U29886 (N_29886,N_29579,N_29547);
nand U29887 (N_29887,N_29697,N_29687);
and U29888 (N_29888,N_29691,N_29512);
xnor U29889 (N_29889,N_29644,N_29622);
and U29890 (N_29890,N_29544,N_29590);
and U29891 (N_29891,N_29539,N_29635);
nand U29892 (N_29892,N_29550,N_29526);
and U29893 (N_29893,N_29486,N_29570);
nor U29894 (N_29894,N_29429,N_29485);
and U29895 (N_29895,N_29591,N_29628);
or U29896 (N_29896,N_29567,N_29524);
nand U29897 (N_29897,N_29643,N_29646);
and U29898 (N_29898,N_29490,N_29494);
or U29899 (N_29899,N_29538,N_29552);
nor U29900 (N_29900,N_29482,N_29488);
nor U29901 (N_29901,N_29562,N_29620);
nor U29902 (N_29902,N_29651,N_29467);
xnor U29903 (N_29903,N_29543,N_29538);
nand U29904 (N_29904,N_29482,N_29466);
nand U29905 (N_29905,N_29517,N_29639);
nand U29906 (N_29906,N_29662,N_29401);
nor U29907 (N_29907,N_29433,N_29601);
nand U29908 (N_29908,N_29569,N_29692);
xnor U29909 (N_29909,N_29584,N_29542);
nor U29910 (N_29910,N_29509,N_29480);
or U29911 (N_29911,N_29662,N_29644);
nor U29912 (N_29912,N_29524,N_29505);
xor U29913 (N_29913,N_29519,N_29539);
and U29914 (N_29914,N_29617,N_29480);
nor U29915 (N_29915,N_29477,N_29680);
or U29916 (N_29916,N_29691,N_29545);
or U29917 (N_29917,N_29580,N_29686);
xnor U29918 (N_29918,N_29613,N_29594);
and U29919 (N_29919,N_29571,N_29506);
or U29920 (N_29920,N_29615,N_29667);
nor U29921 (N_29921,N_29540,N_29411);
nand U29922 (N_29922,N_29493,N_29401);
nand U29923 (N_29923,N_29567,N_29677);
nor U29924 (N_29924,N_29429,N_29670);
xnor U29925 (N_29925,N_29420,N_29475);
and U29926 (N_29926,N_29494,N_29590);
nor U29927 (N_29927,N_29499,N_29584);
xor U29928 (N_29928,N_29425,N_29607);
nand U29929 (N_29929,N_29453,N_29487);
nor U29930 (N_29930,N_29662,N_29445);
xnor U29931 (N_29931,N_29660,N_29546);
nand U29932 (N_29932,N_29512,N_29682);
nor U29933 (N_29933,N_29433,N_29560);
xor U29934 (N_29934,N_29537,N_29551);
nand U29935 (N_29935,N_29654,N_29436);
xnor U29936 (N_29936,N_29684,N_29468);
xor U29937 (N_29937,N_29423,N_29696);
xor U29938 (N_29938,N_29494,N_29503);
and U29939 (N_29939,N_29446,N_29636);
and U29940 (N_29940,N_29684,N_29414);
or U29941 (N_29941,N_29659,N_29468);
and U29942 (N_29942,N_29621,N_29643);
and U29943 (N_29943,N_29420,N_29541);
and U29944 (N_29944,N_29636,N_29625);
nand U29945 (N_29945,N_29463,N_29676);
xnor U29946 (N_29946,N_29469,N_29562);
nand U29947 (N_29947,N_29565,N_29587);
nand U29948 (N_29948,N_29673,N_29693);
xnor U29949 (N_29949,N_29551,N_29504);
nor U29950 (N_29950,N_29561,N_29471);
or U29951 (N_29951,N_29405,N_29490);
and U29952 (N_29952,N_29600,N_29471);
nor U29953 (N_29953,N_29482,N_29599);
nor U29954 (N_29954,N_29679,N_29634);
or U29955 (N_29955,N_29661,N_29591);
and U29956 (N_29956,N_29658,N_29638);
xnor U29957 (N_29957,N_29617,N_29587);
xnor U29958 (N_29958,N_29463,N_29513);
xnor U29959 (N_29959,N_29562,N_29614);
and U29960 (N_29960,N_29573,N_29558);
and U29961 (N_29961,N_29460,N_29444);
xnor U29962 (N_29962,N_29633,N_29506);
or U29963 (N_29963,N_29469,N_29448);
or U29964 (N_29964,N_29543,N_29515);
xor U29965 (N_29965,N_29618,N_29537);
or U29966 (N_29966,N_29458,N_29522);
and U29967 (N_29967,N_29617,N_29544);
nand U29968 (N_29968,N_29648,N_29578);
nor U29969 (N_29969,N_29489,N_29675);
xnor U29970 (N_29970,N_29663,N_29672);
xor U29971 (N_29971,N_29640,N_29528);
and U29972 (N_29972,N_29688,N_29646);
and U29973 (N_29973,N_29517,N_29477);
and U29974 (N_29974,N_29664,N_29667);
nand U29975 (N_29975,N_29678,N_29445);
nand U29976 (N_29976,N_29592,N_29417);
xor U29977 (N_29977,N_29672,N_29653);
or U29978 (N_29978,N_29448,N_29523);
and U29979 (N_29979,N_29610,N_29640);
or U29980 (N_29980,N_29521,N_29402);
nor U29981 (N_29981,N_29524,N_29424);
nor U29982 (N_29982,N_29627,N_29576);
nand U29983 (N_29983,N_29597,N_29573);
or U29984 (N_29984,N_29539,N_29466);
or U29985 (N_29985,N_29618,N_29413);
nand U29986 (N_29986,N_29663,N_29428);
or U29987 (N_29987,N_29615,N_29644);
xnor U29988 (N_29988,N_29484,N_29692);
or U29989 (N_29989,N_29647,N_29567);
nand U29990 (N_29990,N_29617,N_29492);
xnor U29991 (N_29991,N_29411,N_29664);
and U29992 (N_29992,N_29670,N_29430);
nor U29993 (N_29993,N_29646,N_29556);
and U29994 (N_29994,N_29579,N_29449);
xnor U29995 (N_29995,N_29429,N_29464);
nand U29996 (N_29996,N_29668,N_29562);
nor U29997 (N_29997,N_29421,N_29684);
nand U29998 (N_29998,N_29541,N_29612);
nand U29999 (N_29999,N_29468,N_29403);
nor UO_0 (O_0,N_29945,N_29898);
nand UO_1 (O_1,N_29881,N_29882);
xnor UO_2 (O_2,N_29878,N_29923);
xor UO_3 (O_3,N_29744,N_29999);
nor UO_4 (O_4,N_29883,N_29937);
nor UO_5 (O_5,N_29803,N_29816);
or UO_6 (O_6,N_29818,N_29905);
nand UO_7 (O_7,N_29766,N_29833);
xor UO_8 (O_8,N_29787,N_29704);
or UO_9 (O_9,N_29954,N_29807);
xor UO_10 (O_10,N_29758,N_29895);
xnor UO_11 (O_11,N_29777,N_29864);
nand UO_12 (O_12,N_29773,N_29862);
or UO_13 (O_13,N_29910,N_29849);
nand UO_14 (O_14,N_29746,N_29956);
or UO_15 (O_15,N_29771,N_29997);
nand UO_16 (O_16,N_29958,N_29735);
nor UO_17 (O_17,N_29951,N_29934);
and UO_18 (O_18,N_29942,N_29713);
nor UO_19 (O_19,N_29795,N_29877);
xor UO_20 (O_20,N_29949,N_29812);
xnor UO_21 (O_21,N_29897,N_29835);
nor UO_22 (O_22,N_29706,N_29874);
and UO_23 (O_23,N_29707,N_29860);
nor UO_24 (O_24,N_29928,N_29995);
nor UO_25 (O_25,N_29834,N_29988);
nor UO_26 (O_26,N_29739,N_29723);
or UO_27 (O_27,N_29939,N_29983);
or UO_28 (O_28,N_29893,N_29770);
or UO_29 (O_29,N_29960,N_29798);
and UO_30 (O_30,N_29708,N_29901);
nor UO_31 (O_31,N_29973,N_29786);
or UO_32 (O_32,N_29852,N_29953);
xnor UO_33 (O_33,N_29915,N_29793);
or UO_34 (O_34,N_29848,N_29872);
and UO_35 (O_35,N_29709,N_29823);
nand UO_36 (O_36,N_29894,N_29809);
and UO_37 (O_37,N_29909,N_29902);
or UO_38 (O_38,N_29844,N_29733);
or UO_39 (O_39,N_29718,N_29725);
xor UO_40 (O_40,N_29900,N_29979);
and UO_41 (O_41,N_29879,N_29828);
and UO_42 (O_42,N_29841,N_29932);
xnor UO_43 (O_43,N_29734,N_29761);
and UO_44 (O_44,N_29726,N_29991);
and UO_45 (O_45,N_29782,N_29944);
nor UO_46 (O_46,N_29873,N_29821);
nor UO_47 (O_47,N_29822,N_29980);
xor UO_48 (O_48,N_29763,N_29985);
nor UO_49 (O_49,N_29742,N_29840);
and UO_50 (O_50,N_29913,N_29720);
or UO_51 (O_51,N_29886,N_29775);
nand UO_52 (O_52,N_29745,N_29867);
nand UO_53 (O_53,N_29941,N_29866);
nor UO_54 (O_54,N_29887,N_29748);
or UO_55 (O_55,N_29926,N_29827);
or UO_56 (O_56,N_29847,N_29754);
nor UO_57 (O_57,N_29992,N_29929);
xnor UO_58 (O_58,N_29851,N_29832);
nor UO_59 (O_59,N_29868,N_29890);
and UO_60 (O_60,N_29729,N_29751);
nand UO_61 (O_61,N_29857,N_29755);
nand UO_62 (O_62,N_29715,N_29931);
nand UO_63 (O_63,N_29994,N_29876);
xor UO_64 (O_64,N_29853,N_29955);
or UO_65 (O_65,N_29719,N_29998);
or UO_66 (O_66,N_29826,N_29837);
or UO_67 (O_67,N_29804,N_29981);
and UO_68 (O_68,N_29730,N_29982);
nor UO_69 (O_69,N_29987,N_29836);
nand UO_70 (O_70,N_29757,N_29785);
and UO_71 (O_71,N_29800,N_29788);
nand UO_72 (O_72,N_29781,N_29925);
or UO_73 (O_73,N_29967,N_29977);
xnor UO_74 (O_74,N_29768,N_29854);
and UO_75 (O_75,N_29968,N_29774);
nand UO_76 (O_76,N_29728,N_29825);
and UO_77 (O_77,N_29721,N_29701);
nand UO_78 (O_78,N_29984,N_29789);
or UO_79 (O_79,N_29914,N_29861);
nand UO_80 (O_80,N_29815,N_29888);
or UO_81 (O_81,N_29889,N_29790);
xor UO_82 (O_82,N_29884,N_29738);
nor UO_83 (O_83,N_29990,N_29700);
or UO_84 (O_84,N_29917,N_29957);
nor UO_85 (O_85,N_29924,N_29869);
and UO_86 (O_86,N_29904,N_29747);
xnor UO_87 (O_87,N_29920,N_29703);
nand UO_88 (O_88,N_29830,N_29717);
xnor UO_89 (O_89,N_29753,N_29989);
xor UO_90 (O_90,N_29710,N_29791);
or UO_91 (O_91,N_29845,N_29938);
xor UO_92 (O_92,N_29965,N_29930);
and UO_93 (O_93,N_29855,N_29737);
xnor UO_94 (O_94,N_29797,N_29767);
or UO_95 (O_95,N_29842,N_29727);
xnor UO_96 (O_96,N_29950,N_29760);
or UO_97 (O_97,N_29740,N_29711);
nand UO_98 (O_98,N_29962,N_29952);
nor UO_99 (O_99,N_29783,N_29974);
nor UO_100 (O_100,N_29899,N_29839);
and UO_101 (O_101,N_29824,N_29871);
xnor UO_102 (O_102,N_29750,N_29940);
nor UO_103 (O_103,N_29817,N_29922);
nor UO_104 (O_104,N_29801,N_29892);
or UO_105 (O_105,N_29732,N_29759);
nand UO_106 (O_106,N_29891,N_29880);
xnor UO_107 (O_107,N_29705,N_29858);
nand UO_108 (O_108,N_29769,N_29943);
and UO_109 (O_109,N_29896,N_29933);
nand UO_110 (O_110,N_29850,N_29903);
xor UO_111 (O_111,N_29838,N_29731);
nor UO_112 (O_112,N_29870,N_29946);
xnor UO_113 (O_113,N_29908,N_29947);
or UO_114 (O_114,N_29784,N_29918);
and UO_115 (O_115,N_29741,N_29978);
nand UO_116 (O_116,N_29752,N_29736);
and UO_117 (O_117,N_29846,N_29970);
and UO_118 (O_118,N_29813,N_29794);
xnor UO_119 (O_119,N_29843,N_29765);
xor UO_120 (O_120,N_29811,N_29756);
and UO_121 (O_121,N_29814,N_29819);
and UO_122 (O_122,N_29986,N_29961);
nand UO_123 (O_123,N_29875,N_29796);
nor UO_124 (O_124,N_29764,N_29863);
and UO_125 (O_125,N_29969,N_29959);
nand UO_126 (O_126,N_29993,N_29966);
and UO_127 (O_127,N_29964,N_29780);
nor UO_128 (O_128,N_29912,N_29805);
xnor UO_129 (O_129,N_29820,N_29919);
nor UO_130 (O_130,N_29972,N_29911);
or UO_131 (O_131,N_29963,N_29859);
and UO_132 (O_132,N_29935,N_29885);
and UO_133 (O_133,N_29916,N_29802);
nor UO_134 (O_134,N_29948,N_29778);
and UO_135 (O_135,N_29716,N_29856);
and UO_136 (O_136,N_29749,N_29971);
xnor UO_137 (O_137,N_29996,N_29762);
and UO_138 (O_138,N_29779,N_29975);
nand UO_139 (O_139,N_29906,N_29776);
nor UO_140 (O_140,N_29927,N_29702);
nand UO_141 (O_141,N_29714,N_29799);
xor UO_142 (O_142,N_29976,N_29806);
nand UO_143 (O_143,N_29936,N_29792);
and UO_144 (O_144,N_29772,N_29743);
or UO_145 (O_145,N_29808,N_29722);
nand UO_146 (O_146,N_29810,N_29921);
and UO_147 (O_147,N_29829,N_29712);
nand UO_148 (O_148,N_29865,N_29907);
and UO_149 (O_149,N_29724,N_29831);
xor UO_150 (O_150,N_29968,N_29864);
xnor UO_151 (O_151,N_29974,N_29782);
nor UO_152 (O_152,N_29944,N_29965);
and UO_153 (O_153,N_29822,N_29936);
or UO_154 (O_154,N_29799,N_29824);
xnor UO_155 (O_155,N_29946,N_29839);
nand UO_156 (O_156,N_29717,N_29885);
nand UO_157 (O_157,N_29799,N_29843);
and UO_158 (O_158,N_29891,N_29757);
or UO_159 (O_159,N_29969,N_29999);
xnor UO_160 (O_160,N_29719,N_29951);
nand UO_161 (O_161,N_29751,N_29884);
nor UO_162 (O_162,N_29791,N_29819);
xnor UO_163 (O_163,N_29961,N_29851);
and UO_164 (O_164,N_29710,N_29943);
and UO_165 (O_165,N_29882,N_29880);
nand UO_166 (O_166,N_29900,N_29962);
and UO_167 (O_167,N_29713,N_29723);
or UO_168 (O_168,N_29943,N_29878);
or UO_169 (O_169,N_29935,N_29806);
xnor UO_170 (O_170,N_29915,N_29923);
nand UO_171 (O_171,N_29768,N_29734);
nand UO_172 (O_172,N_29947,N_29826);
nor UO_173 (O_173,N_29815,N_29869);
nor UO_174 (O_174,N_29811,N_29746);
nor UO_175 (O_175,N_29912,N_29723);
xnor UO_176 (O_176,N_29894,N_29917);
and UO_177 (O_177,N_29701,N_29787);
and UO_178 (O_178,N_29829,N_29783);
nor UO_179 (O_179,N_29971,N_29801);
or UO_180 (O_180,N_29985,N_29943);
xnor UO_181 (O_181,N_29796,N_29743);
and UO_182 (O_182,N_29774,N_29830);
and UO_183 (O_183,N_29829,N_29906);
nand UO_184 (O_184,N_29801,N_29873);
xnor UO_185 (O_185,N_29863,N_29780);
xnor UO_186 (O_186,N_29840,N_29934);
xor UO_187 (O_187,N_29721,N_29962);
or UO_188 (O_188,N_29813,N_29821);
xnor UO_189 (O_189,N_29889,N_29920);
and UO_190 (O_190,N_29737,N_29760);
or UO_191 (O_191,N_29853,N_29913);
nor UO_192 (O_192,N_29799,N_29816);
and UO_193 (O_193,N_29825,N_29719);
and UO_194 (O_194,N_29784,N_29703);
nand UO_195 (O_195,N_29993,N_29723);
or UO_196 (O_196,N_29924,N_29830);
xnor UO_197 (O_197,N_29838,N_29804);
or UO_198 (O_198,N_29778,N_29878);
nand UO_199 (O_199,N_29911,N_29881);
nor UO_200 (O_200,N_29996,N_29708);
or UO_201 (O_201,N_29712,N_29791);
nor UO_202 (O_202,N_29715,N_29724);
nor UO_203 (O_203,N_29714,N_29858);
nand UO_204 (O_204,N_29869,N_29958);
or UO_205 (O_205,N_29796,N_29838);
nand UO_206 (O_206,N_29770,N_29941);
or UO_207 (O_207,N_29807,N_29969);
and UO_208 (O_208,N_29783,N_29935);
xor UO_209 (O_209,N_29748,N_29733);
and UO_210 (O_210,N_29819,N_29881);
and UO_211 (O_211,N_29832,N_29786);
or UO_212 (O_212,N_29978,N_29754);
xnor UO_213 (O_213,N_29801,N_29902);
or UO_214 (O_214,N_29794,N_29945);
nor UO_215 (O_215,N_29947,N_29722);
or UO_216 (O_216,N_29879,N_29837);
nor UO_217 (O_217,N_29898,N_29712);
nand UO_218 (O_218,N_29821,N_29843);
xnor UO_219 (O_219,N_29978,N_29716);
nand UO_220 (O_220,N_29941,N_29822);
or UO_221 (O_221,N_29784,N_29728);
xnor UO_222 (O_222,N_29969,N_29792);
or UO_223 (O_223,N_29737,N_29817);
and UO_224 (O_224,N_29854,N_29859);
or UO_225 (O_225,N_29957,N_29715);
and UO_226 (O_226,N_29808,N_29861);
xnor UO_227 (O_227,N_29834,N_29845);
nor UO_228 (O_228,N_29875,N_29838);
or UO_229 (O_229,N_29774,N_29948);
nand UO_230 (O_230,N_29741,N_29731);
or UO_231 (O_231,N_29815,N_29761);
and UO_232 (O_232,N_29848,N_29827);
xor UO_233 (O_233,N_29956,N_29969);
or UO_234 (O_234,N_29723,N_29792);
nor UO_235 (O_235,N_29913,N_29724);
nand UO_236 (O_236,N_29923,N_29876);
xor UO_237 (O_237,N_29780,N_29972);
and UO_238 (O_238,N_29713,N_29929);
xor UO_239 (O_239,N_29825,N_29704);
and UO_240 (O_240,N_29769,N_29862);
or UO_241 (O_241,N_29896,N_29907);
nor UO_242 (O_242,N_29732,N_29790);
or UO_243 (O_243,N_29853,N_29937);
or UO_244 (O_244,N_29843,N_29863);
xor UO_245 (O_245,N_29881,N_29995);
xor UO_246 (O_246,N_29869,N_29940);
or UO_247 (O_247,N_29977,N_29722);
and UO_248 (O_248,N_29850,N_29709);
nand UO_249 (O_249,N_29707,N_29951);
and UO_250 (O_250,N_29709,N_29854);
nand UO_251 (O_251,N_29966,N_29708);
or UO_252 (O_252,N_29952,N_29789);
nor UO_253 (O_253,N_29765,N_29745);
or UO_254 (O_254,N_29949,N_29817);
nand UO_255 (O_255,N_29890,N_29755);
or UO_256 (O_256,N_29817,N_29867);
and UO_257 (O_257,N_29947,N_29997);
nor UO_258 (O_258,N_29782,N_29769);
xnor UO_259 (O_259,N_29838,N_29819);
or UO_260 (O_260,N_29784,N_29740);
xnor UO_261 (O_261,N_29934,N_29853);
xor UO_262 (O_262,N_29813,N_29722);
nor UO_263 (O_263,N_29740,N_29975);
or UO_264 (O_264,N_29776,N_29980);
xnor UO_265 (O_265,N_29920,N_29925);
xnor UO_266 (O_266,N_29819,N_29786);
or UO_267 (O_267,N_29790,N_29774);
xor UO_268 (O_268,N_29889,N_29873);
and UO_269 (O_269,N_29922,N_29735);
nor UO_270 (O_270,N_29746,N_29933);
xor UO_271 (O_271,N_29959,N_29908);
and UO_272 (O_272,N_29914,N_29729);
xor UO_273 (O_273,N_29852,N_29840);
or UO_274 (O_274,N_29801,N_29738);
or UO_275 (O_275,N_29933,N_29909);
or UO_276 (O_276,N_29817,N_29805);
and UO_277 (O_277,N_29773,N_29821);
nor UO_278 (O_278,N_29975,N_29943);
or UO_279 (O_279,N_29838,N_29757);
or UO_280 (O_280,N_29939,N_29967);
xor UO_281 (O_281,N_29891,N_29747);
nor UO_282 (O_282,N_29774,N_29999);
or UO_283 (O_283,N_29977,N_29944);
nand UO_284 (O_284,N_29965,N_29990);
xnor UO_285 (O_285,N_29733,N_29932);
nor UO_286 (O_286,N_29711,N_29807);
nor UO_287 (O_287,N_29903,N_29986);
xnor UO_288 (O_288,N_29784,N_29849);
and UO_289 (O_289,N_29988,N_29860);
nand UO_290 (O_290,N_29700,N_29786);
nor UO_291 (O_291,N_29982,N_29718);
and UO_292 (O_292,N_29897,N_29740);
nor UO_293 (O_293,N_29892,N_29828);
or UO_294 (O_294,N_29775,N_29736);
or UO_295 (O_295,N_29995,N_29745);
and UO_296 (O_296,N_29831,N_29848);
nor UO_297 (O_297,N_29761,N_29800);
nor UO_298 (O_298,N_29908,N_29865);
nor UO_299 (O_299,N_29873,N_29905);
and UO_300 (O_300,N_29863,N_29809);
nor UO_301 (O_301,N_29974,N_29701);
nand UO_302 (O_302,N_29713,N_29760);
xnor UO_303 (O_303,N_29716,N_29984);
xor UO_304 (O_304,N_29763,N_29965);
xor UO_305 (O_305,N_29789,N_29909);
xor UO_306 (O_306,N_29811,N_29896);
and UO_307 (O_307,N_29878,N_29749);
and UO_308 (O_308,N_29834,N_29843);
xor UO_309 (O_309,N_29704,N_29842);
or UO_310 (O_310,N_29830,N_29716);
and UO_311 (O_311,N_29759,N_29853);
xnor UO_312 (O_312,N_29925,N_29706);
and UO_313 (O_313,N_29883,N_29840);
nor UO_314 (O_314,N_29884,N_29777);
or UO_315 (O_315,N_29793,N_29712);
nor UO_316 (O_316,N_29729,N_29860);
and UO_317 (O_317,N_29721,N_29933);
xor UO_318 (O_318,N_29754,N_29943);
or UO_319 (O_319,N_29974,N_29848);
nand UO_320 (O_320,N_29790,N_29915);
nand UO_321 (O_321,N_29777,N_29916);
xor UO_322 (O_322,N_29982,N_29925);
or UO_323 (O_323,N_29872,N_29748);
xor UO_324 (O_324,N_29812,N_29866);
nor UO_325 (O_325,N_29709,N_29814);
and UO_326 (O_326,N_29723,N_29988);
and UO_327 (O_327,N_29814,N_29825);
nand UO_328 (O_328,N_29793,N_29951);
xnor UO_329 (O_329,N_29723,N_29770);
and UO_330 (O_330,N_29719,N_29776);
or UO_331 (O_331,N_29736,N_29977);
xnor UO_332 (O_332,N_29878,N_29884);
and UO_333 (O_333,N_29785,N_29868);
nand UO_334 (O_334,N_29824,N_29942);
nor UO_335 (O_335,N_29990,N_29801);
xnor UO_336 (O_336,N_29764,N_29890);
nor UO_337 (O_337,N_29733,N_29754);
xnor UO_338 (O_338,N_29728,N_29869);
and UO_339 (O_339,N_29917,N_29967);
nand UO_340 (O_340,N_29968,N_29914);
nor UO_341 (O_341,N_29710,N_29842);
or UO_342 (O_342,N_29819,N_29912);
nand UO_343 (O_343,N_29773,N_29964);
nand UO_344 (O_344,N_29949,N_29885);
xnor UO_345 (O_345,N_29740,N_29846);
nor UO_346 (O_346,N_29801,N_29732);
or UO_347 (O_347,N_29774,N_29924);
and UO_348 (O_348,N_29929,N_29873);
xnor UO_349 (O_349,N_29949,N_29783);
and UO_350 (O_350,N_29754,N_29871);
nand UO_351 (O_351,N_29943,N_29851);
and UO_352 (O_352,N_29734,N_29889);
nor UO_353 (O_353,N_29782,N_29701);
nand UO_354 (O_354,N_29878,N_29900);
nand UO_355 (O_355,N_29966,N_29745);
or UO_356 (O_356,N_29919,N_29809);
nor UO_357 (O_357,N_29862,N_29897);
and UO_358 (O_358,N_29703,N_29807);
xnor UO_359 (O_359,N_29896,N_29732);
or UO_360 (O_360,N_29798,N_29817);
or UO_361 (O_361,N_29885,N_29915);
xor UO_362 (O_362,N_29923,N_29824);
nor UO_363 (O_363,N_29815,N_29727);
nand UO_364 (O_364,N_29746,N_29989);
nand UO_365 (O_365,N_29783,N_29870);
xor UO_366 (O_366,N_29936,N_29750);
or UO_367 (O_367,N_29762,N_29769);
and UO_368 (O_368,N_29741,N_29798);
and UO_369 (O_369,N_29946,N_29931);
or UO_370 (O_370,N_29957,N_29975);
and UO_371 (O_371,N_29880,N_29701);
xnor UO_372 (O_372,N_29896,N_29816);
nor UO_373 (O_373,N_29827,N_29735);
and UO_374 (O_374,N_29755,N_29853);
nand UO_375 (O_375,N_29832,N_29892);
nand UO_376 (O_376,N_29892,N_29739);
and UO_377 (O_377,N_29772,N_29704);
nand UO_378 (O_378,N_29784,N_29895);
and UO_379 (O_379,N_29902,N_29784);
or UO_380 (O_380,N_29777,N_29735);
nor UO_381 (O_381,N_29758,N_29770);
and UO_382 (O_382,N_29951,N_29746);
or UO_383 (O_383,N_29701,N_29870);
or UO_384 (O_384,N_29842,N_29998);
and UO_385 (O_385,N_29949,N_29702);
xor UO_386 (O_386,N_29882,N_29797);
xnor UO_387 (O_387,N_29902,N_29919);
xor UO_388 (O_388,N_29955,N_29808);
nor UO_389 (O_389,N_29772,N_29898);
nor UO_390 (O_390,N_29969,N_29914);
or UO_391 (O_391,N_29770,N_29899);
xor UO_392 (O_392,N_29910,N_29835);
nor UO_393 (O_393,N_29795,N_29723);
nor UO_394 (O_394,N_29811,N_29985);
or UO_395 (O_395,N_29946,N_29922);
or UO_396 (O_396,N_29842,N_29928);
nand UO_397 (O_397,N_29842,N_29730);
and UO_398 (O_398,N_29824,N_29785);
or UO_399 (O_399,N_29772,N_29782);
nand UO_400 (O_400,N_29831,N_29720);
nand UO_401 (O_401,N_29977,N_29938);
nor UO_402 (O_402,N_29959,N_29841);
nand UO_403 (O_403,N_29755,N_29707);
nand UO_404 (O_404,N_29939,N_29784);
and UO_405 (O_405,N_29950,N_29778);
or UO_406 (O_406,N_29701,N_29998);
nand UO_407 (O_407,N_29884,N_29705);
and UO_408 (O_408,N_29836,N_29728);
nor UO_409 (O_409,N_29943,N_29755);
and UO_410 (O_410,N_29733,N_29865);
nor UO_411 (O_411,N_29974,N_29875);
or UO_412 (O_412,N_29949,N_29863);
or UO_413 (O_413,N_29828,N_29803);
or UO_414 (O_414,N_29891,N_29812);
and UO_415 (O_415,N_29991,N_29946);
nand UO_416 (O_416,N_29738,N_29994);
or UO_417 (O_417,N_29793,N_29727);
nor UO_418 (O_418,N_29985,N_29968);
nand UO_419 (O_419,N_29870,N_29824);
xnor UO_420 (O_420,N_29833,N_29996);
or UO_421 (O_421,N_29857,N_29811);
nand UO_422 (O_422,N_29774,N_29702);
nor UO_423 (O_423,N_29931,N_29907);
or UO_424 (O_424,N_29947,N_29903);
nand UO_425 (O_425,N_29729,N_29874);
or UO_426 (O_426,N_29760,N_29968);
nor UO_427 (O_427,N_29713,N_29890);
xor UO_428 (O_428,N_29972,N_29773);
nor UO_429 (O_429,N_29836,N_29771);
and UO_430 (O_430,N_29830,N_29759);
nand UO_431 (O_431,N_29966,N_29702);
nand UO_432 (O_432,N_29801,N_29912);
nand UO_433 (O_433,N_29940,N_29703);
nand UO_434 (O_434,N_29987,N_29740);
nor UO_435 (O_435,N_29820,N_29717);
nor UO_436 (O_436,N_29891,N_29777);
nand UO_437 (O_437,N_29731,N_29903);
nor UO_438 (O_438,N_29804,N_29781);
xnor UO_439 (O_439,N_29779,N_29753);
and UO_440 (O_440,N_29984,N_29753);
nor UO_441 (O_441,N_29866,N_29888);
xnor UO_442 (O_442,N_29932,N_29850);
and UO_443 (O_443,N_29710,N_29756);
or UO_444 (O_444,N_29773,N_29746);
or UO_445 (O_445,N_29909,N_29801);
xnor UO_446 (O_446,N_29765,N_29828);
or UO_447 (O_447,N_29846,N_29825);
nand UO_448 (O_448,N_29887,N_29891);
nor UO_449 (O_449,N_29849,N_29776);
xnor UO_450 (O_450,N_29963,N_29824);
nor UO_451 (O_451,N_29790,N_29910);
and UO_452 (O_452,N_29809,N_29719);
nor UO_453 (O_453,N_29911,N_29764);
nor UO_454 (O_454,N_29927,N_29978);
or UO_455 (O_455,N_29705,N_29978);
and UO_456 (O_456,N_29820,N_29895);
xnor UO_457 (O_457,N_29974,N_29939);
xor UO_458 (O_458,N_29949,N_29880);
and UO_459 (O_459,N_29785,N_29780);
or UO_460 (O_460,N_29818,N_29796);
nor UO_461 (O_461,N_29918,N_29871);
nand UO_462 (O_462,N_29948,N_29738);
and UO_463 (O_463,N_29858,N_29845);
nor UO_464 (O_464,N_29828,N_29702);
xnor UO_465 (O_465,N_29821,N_29757);
or UO_466 (O_466,N_29756,N_29925);
nand UO_467 (O_467,N_29986,N_29742);
and UO_468 (O_468,N_29887,N_29792);
nand UO_469 (O_469,N_29741,N_29892);
and UO_470 (O_470,N_29840,N_29804);
and UO_471 (O_471,N_29797,N_29943);
and UO_472 (O_472,N_29967,N_29807);
nor UO_473 (O_473,N_29981,N_29950);
nand UO_474 (O_474,N_29863,N_29723);
xnor UO_475 (O_475,N_29910,N_29932);
and UO_476 (O_476,N_29744,N_29878);
xor UO_477 (O_477,N_29999,N_29807);
xnor UO_478 (O_478,N_29861,N_29926);
nand UO_479 (O_479,N_29908,N_29835);
xor UO_480 (O_480,N_29912,N_29980);
xor UO_481 (O_481,N_29881,N_29735);
xnor UO_482 (O_482,N_29941,N_29867);
and UO_483 (O_483,N_29813,N_29929);
or UO_484 (O_484,N_29703,N_29944);
nand UO_485 (O_485,N_29908,N_29741);
or UO_486 (O_486,N_29896,N_29850);
nand UO_487 (O_487,N_29888,N_29771);
and UO_488 (O_488,N_29744,N_29949);
nor UO_489 (O_489,N_29977,N_29936);
nor UO_490 (O_490,N_29738,N_29730);
and UO_491 (O_491,N_29768,N_29919);
nor UO_492 (O_492,N_29830,N_29907);
xnor UO_493 (O_493,N_29989,N_29972);
xor UO_494 (O_494,N_29997,N_29739);
xor UO_495 (O_495,N_29722,N_29927);
nor UO_496 (O_496,N_29733,N_29960);
and UO_497 (O_497,N_29727,N_29760);
nor UO_498 (O_498,N_29941,N_29719);
nor UO_499 (O_499,N_29995,N_29707);
and UO_500 (O_500,N_29957,N_29873);
xnor UO_501 (O_501,N_29796,N_29863);
nand UO_502 (O_502,N_29800,N_29845);
nor UO_503 (O_503,N_29757,N_29855);
nand UO_504 (O_504,N_29847,N_29828);
and UO_505 (O_505,N_29724,N_29884);
or UO_506 (O_506,N_29847,N_29982);
nor UO_507 (O_507,N_29862,N_29792);
nor UO_508 (O_508,N_29711,N_29943);
xor UO_509 (O_509,N_29805,N_29793);
nand UO_510 (O_510,N_29755,N_29848);
and UO_511 (O_511,N_29782,N_29805);
and UO_512 (O_512,N_29926,N_29891);
or UO_513 (O_513,N_29703,N_29732);
and UO_514 (O_514,N_29886,N_29840);
or UO_515 (O_515,N_29770,N_29838);
and UO_516 (O_516,N_29936,N_29985);
and UO_517 (O_517,N_29851,N_29781);
nor UO_518 (O_518,N_29776,N_29791);
nand UO_519 (O_519,N_29885,N_29819);
xor UO_520 (O_520,N_29818,N_29951);
and UO_521 (O_521,N_29999,N_29916);
xor UO_522 (O_522,N_29882,N_29929);
or UO_523 (O_523,N_29751,N_29835);
nand UO_524 (O_524,N_29736,N_29866);
and UO_525 (O_525,N_29710,N_29855);
and UO_526 (O_526,N_29865,N_29810);
nand UO_527 (O_527,N_29975,N_29728);
or UO_528 (O_528,N_29736,N_29926);
xnor UO_529 (O_529,N_29960,N_29833);
nor UO_530 (O_530,N_29879,N_29858);
and UO_531 (O_531,N_29811,N_29903);
or UO_532 (O_532,N_29724,N_29734);
xor UO_533 (O_533,N_29828,N_29994);
nand UO_534 (O_534,N_29818,N_29930);
and UO_535 (O_535,N_29817,N_29869);
nor UO_536 (O_536,N_29912,N_29709);
nand UO_537 (O_537,N_29856,N_29895);
or UO_538 (O_538,N_29824,N_29924);
and UO_539 (O_539,N_29702,N_29963);
nor UO_540 (O_540,N_29971,N_29942);
nor UO_541 (O_541,N_29902,N_29825);
xor UO_542 (O_542,N_29997,N_29819);
xor UO_543 (O_543,N_29875,N_29996);
or UO_544 (O_544,N_29804,N_29717);
or UO_545 (O_545,N_29876,N_29953);
nand UO_546 (O_546,N_29739,N_29864);
and UO_547 (O_547,N_29795,N_29944);
xnor UO_548 (O_548,N_29977,N_29984);
nor UO_549 (O_549,N_29935,N_29842);
xnor UO_550 (O_550,N_29867,N_29772);
or UO_551 (O_551,N_29955,N_29781);
xnor UO_552 (O_552,N_29871,N_29774);
or UO_553 (O_553,N_29875,N_29811);
nor UO_554 (O_554,N_29762,N_29913);
nor UO_555 (O_555,N_29823,N_29837);
or UO_556 (O_556,N_29880,N_29857);
xnor UO_557 (O_557,N_29700,N_29840);
or UO_558 (O_558,N_29832,N_29818);
and UO_559 (O_559,N_29922,N_29871);
nor UO_560 (O_560,N_29777,N_29756);
or UO_561 (O_561,N_29863,N_29890);
nand UO_562 (O_562,N_29709,N_29926);
or UO_563 (O_563,N_29938,N_29901);
nand UO_564 (O_564,N_29748,N_29835);
or UO_565 (O_565,N_29862,N_29974);
or UO_566 (O_566,N_29715,N_29987);
xnor UO_567 (O_567,N_29881,N_29723);
nor UO_568 (O_568,N_29904,N_29969);
or UO_569 (O_569,N_29939,N_29788);
xnor UO_570 (O_570,N_29787,N_29897);
or UO_571 (O_571,N_29728,N_29903);
nor UO_572 (O_572,N_29912,N_29764);
nand UO_573 (O_573,N_29761,N_29897);
and UO_574 (O_574,N_29924,N_29733);
xor UO_575 (O_575,N_29913,N_29800);
nor UO_576 (O_576,N_29722,N_29934);
xnor UO_577 (O_577,N_29705,N_29788);
and UO_578 (O_578,N_29834,N_29894);
nand UO_579 (O_579,N_29889,N_29908);
nor UO_580 (O_580,N_29963,N_29781);
xor UO_581 (O_581,N_29998,N_29982);
nand UO_582 (O_582,N_29983,N_29742);
and UO_583 (O_583,N_29720,N_29804);
and UO_584 (O_584,N_29803,N_29984);
and UO_585 (O_585,N_29766,N_29991);
or UO_586 (O_586,N_29943,N_29707);
xnor UO_587 (O_587,N_29711,N_29751);
nor UO_588 (O_588,N_29752,N_29982);
and UO_589 (O_589,N_29923,N_29919);
or UO_590 (O_590,N_29902,N_29920);
and UO_591 (O_591,N_29916,N_29795);
or UO_592 (O_592,N_29799,N_29913);
or UO_593 (O_593,N_29777,N_29788);
or UO_594 (O_594,N_29735,N_29778);
nor UO_595 (O_595,N_29810,N_29967);
nor UO_596 (O_596,N_29753,N_29789);
nor UO_597 (O_597,N_29888,N_29783);
nand UO_598 (O_598,N_29951,N_29871);
nand UO_599 (O_599,N_29960,N_29708);
or UO_600 (O_600,N_29737,N_29792);
xnor UO_601 (O_601,N_29807,N_29968);
nor UO_602 (O_602,N_29756,N_29896);
or UO_603 (O_603,N_29868,N_29941);
nand UO_604 (O_604,N_29831,N_29737);
nand UO_605 (O_605,N_29790,N_29865);
nor UO_606 (O_606,N_29950,N_29824);
nor UO_607 (O_607,N_29756,N_29922);
nand UO_608 (O_608,N_29999,N_29760);
and UO_609 (O_609,N_29965,N_29909);
xor UO_610 (O_610,N_29716,N_29745);
or UO_611 (O_611,N_29711,N_29884);
and UO_612 (O_612,N_29837,N_29943);
or UO_613 (O_613,N_29985,N_29933);
and UO_614 (O_614,N_29741,N_29939);
xnor UO_615 (O_615,N_29967,N_29842);
or UO_616 (O_616,N_29727,N_29861);
and UO_617 (O_617,N_29796,N_29997);
nand UO_618 (O_618,N_29967,N_29840);
xor UO_619 (O_619,N_29845,N_29896);
xnor UO_620 (O_620,N_29777,N_29936);
nand UO_621 (O_621,N_29809,N_29908);
xor UO_622 (O_622,N_29736,N_29961);
nand UO_623 (O_623,N_29848,N_29940);
and UO_624 (O_624,N_29723,N_29914);
nand UO_625 (O_625,N_29783,N_29779);
xor UO_626 (O_626,N_29958,N_29926);
nor UO_627 (O_627,N_29765,N_29983);
nor UO_628 (O_628,N_29832,N_29945);
xor UO_629 (O_629,N_29997,N_29792);
nand UO_630 (O_630,N_29704,N_29707);
or UO_631 (O_631,N_29841,N_29853);
xnor UO_632 (O_632,N_29704,N_29713);
xor UO_633 (O_633,N_29711,N_29918);
nor UO_634 (O_634,N_29965,N_29811);
nor UO_635 (O_635,N_29848,N_29771);
or UO_636 (O_636,N_29928,N_29827);
nor UO_637 (O_637,N_29938,N_29752);
nor UO_638 (O_638,N_29712,N_29874);
nor UO_639 (O_639,N_29902,N_29778);
or UO_640 (O_640,N_29999,N_29913);
nand UO_641 (O_641,N_29758,N_29808);
xnor UO_642 (O_642,N_29723,N_29728);
or UO_643 (O_643,N_29702,N_29852);
and UO_644 (O_644,N_29926,N_29920);
nor UO_645 (O_645,N_29967,N_29989);
xor UO_646 (O_646,N_29940,N_29983);
xor UO_647 (O_647,N_29828,N_29749);
and UO_648 (O_648,N_29879,N_29747);
and UO_649 (O_649,N_29860,N_29963);
or UO_650 (O_650,N_29734,N_29760);
xor UO_651 (O_651,N_29767,N_29729);
or UO_652 (O_652,N_29952,N_29911);
xnor UO_653 (O_653,N_29879,N_29731);
nand UO_654 (O_654,N_29727,N_29881);
xnor UO_655 (O_655,N_29950,N_29848);
xnor UO_656 (O_656,N_29739,N_29947);
nor UO_657 (O_657,N_29858,N_29824);
nor UO_658 (O_658,N_29866,N_29969);
or UO_659 (O_659,N_29709,N_29703);
or UO_660 (O_660,N_29922,N_29763);
nand UO_661 (O_661,N_29836,N_29738);
or UO_662 (O_662,N_29722,N_29915);
nand UO_663 (O_663,N_29791,N_29986);
nor UO_664 (O_664,N_29779,N_29872);
xnor UO_665 (O_665,N_29811,N_29921);
nand UO_666 (O_666,N_29740,N_29847);
nor UO_667 (O_667,N_29991,N_29741);
and UO_668 (O_668,N_29875,N_29742);
or UO_669 (O_669,N_29986,N_29829);
and UO_670 (O_670,N_29728,N_29764);
nor UO_671 (O_671,N_29711,N_29793);
or UO_672 (O_672,N_29774,N_29845);
or UO_673 (O_673,N_29840,N_29799);
nor UO_674 (O_674,N_29912,N_29717);
nand UO_675 (O_675,N_29843,N_29717);
or UO_676 (O_676,N_29891,N_29851);
nand UO_677 (O_677,N_29898,N_29991);
or UO_678 (O_678,N_29955,N_29798);
nor UO_679 (O_679,N_29974,N_29943);
nor UO_680 (O_680,N_29976,N_29825);
nand UO_681 (O_681,N_29820,N_29831);
and UO_682 (O_682,N_29867,N_29792);
nor UO_683 (O_683,N_29879,N_29965);
nand UO_684 (O_684,N_29765,N_29806);
and UO_685 (O_685,N_29759,N_29902);
and UO_686 (O_686,N_29840,N_29753);
and UO_687 (O_687,N_29950,N_29834);
or UO_688 (O_688,N_29846,N_29803);
xor UO_689 (O_689,N_29896,N_29838);
and UO_690 (O_690,N_29807,N_29702);
or UO_691 (O_691,N_29763,N_29717);
and UO_692 (O_692,N_29895,N_29806);
and UO_693 (O_693,N_29870,N_29880);
nor UO_694 (O_694,N_29860,N_29811);
or UO_695 (O_695,N_29892,N_29884);
or UO_696 (O_696,N_29988,N_29814);
nand UO_697 (O_697,N_29948,N_29848);
or UO_698 (O_698,N_29768,N_29863);
nor UO_699 (O_699,N_29975,N_29947);
nand UO_700 (O_700,N_29811,N_29871);
nand UO_701 (O_701,N_29713,N_29869);
xnor UO_702 (O_702,N_29974,N_29990);
xnor UO_703 (O_703,N_29810,N_29701);
nand UO_704 (O_704,N_29926,N_29797);
nor UO_705 (O_705,N_29949,N_29972);
or UO_706 (O_706,N_29882,N_29759);
xnor UO_707 (O_707,N_29894,N_29755);
nor UO_708 (O_708,N_29768,N_29872);
and UO_709 (O_709,N_29794,N_29835);
and UO_710 (O_710,N_29728,N_29805);
nor UO_711 (O_711,N_29944,N_29982);
nor UO_712 (O_712,N_29968,N_29779);
xnor UO_713 (O_713,N_29878,N_29718);
nand UO_714 (O_714,N_29712,N_29753);
or UO_715 (O_715,N_29877,N_29985);
xor UO_716 (O_716,N_29707,N_29765);
nand UO_717 (O_717,N_29796,N_29907);
and UO_718 (O_718,N_29798,N_29870);
nor UO_719 (O_719,N_29817,N_29848);
and UO_720 (O_720,N_29827,N_29972);
nor UO_721 (O_721,N_29857,N_29831);
and UO_722 (O_722,N_29707,N_29930);
nand UO_723 (O_723,N_29755,N_29948);
xnor UO_724 (O_724,N_29852,N_29929);
nor UO_725 (O_725,N_29977,N_29768);
nor UO_726 (O_726,N_29952,N_29910);
nor UO_727 (O_727,N_29818,N_29709);
nor UO_728 (O_728,N_29709,N_29928);
xnor UO_729 (O_729,N_29809,N_29932);
or UO_730 (O_730,N_29993,N_29744);
xor UO_731 (O_731,N_29707,N_29862);
or UO_732 (O_732,N_29955,N_29927);
or UO_733 (O_733,N_29801,N_29923);
nor UO_734 (O_734,N_29924,N_29741);
nor UO_735 (O_735,N_29719,N_29796);
or UO_736 (O_736,N_29829,N_29726);
or UO_737 (O_737,N_29767,N_29926);
xor UO_738 (O_738,N_29834,N_29797);
and UO_739 (O_739,N_29924,N_29765);
nand UO_740 (O_740,N_29985,N_29856);
and UO_741 (O_741,N_29852,N_29823);
nand UO_742 (O_742,N_29783,N_29971);
nor UO_743 (O_743,N_29742,N_29862);
nand UO_744 (O_744,N_29954,N_29718);
xor UO_745 (O_745,N_29753,N_29981);
nand UO_746 (O_746,N_29721,N_29838);
nand UO_747 (O_747,N_29879,N_29953);
nand UO_748 (O_748,N_29835,N_29796);
or UO_749 (O_749,N_29753,N_29922);
or UO_750 (O_750,N_29913,N_29889);
xor UO_751 (O_751,N_29944,N_29731);
or UO_752 (O_752,N_29741,N_29733);
nand UO_753 (O_753,N_29835,N_29872);
and UO_754 (O_754,N_29910,N_29853);
xor UO_755 (O_755,N_29704,N_29788);
xnor UO_756 (O_756,N_29887,N_29769);
and UO_757 (O_757,N_29736,N_29980);
xor UO_758 (O_758,N_29841,N_29872);
or UO_759 (O_759,N_29821,N_29886);
xor UO_760 (O_760,N_29865,N_29970);
nor UO_761 (O_761,N_29846,N_29933);
nand UO_762 (O_762,N_29900,N_29798);
xnor UO_763 (O_763,N_29738,N_29838);
xnor UO_764 (O_764,N_29760,N_29725);
nand UO_765 (O_765,N_29822,N_29958);
xnor UO_766 (O_766,N_29716,N_29726);
nand UO_767 (O_767,N_29796,N_29815);
xor UO_768 (O_768,N_29959,N_29779);
nor UO_769 (O_769,N_29807,N_29915);
and UO_770 (O_770,N_29919,N_29803);
or UO_771 (O_771,N_29857,N_29727);
or UO_772 (O_772,N_29988,N_29859);
and UO_773 (O_773,N_29945,N_29760);
xor UO_774 (O_774,N_29970,N_29736);
or UO_775 (O_775,N_29806,N_29990);
or UO_776 (O_776,N_29835,N_29847);
xor UO_777 (O_777,N_29719,N_29761);
nor UO_778 (O_778,N_29750,N_29714);
nor UO_779 (O_779,N_29914,N_29721);
xnor UO_780 (O_780,N_29791,N_29931);
nand UO_781 (O_781,N_29874,N_29838);
xor UO_782 (O_782,N_29722,N_29875);
nand UO_783 (O_783,N_29887,N_29849);
xor UO_784 (O_784,N_29882,N_29903);
or UO_785 (O_785,N_29885,N_29826);
nand UO_786 (O_786,N_29896,N_29765);
nor UO_787 (O_787,N_29939,N_29857);
or UO_788 (O_788,N_29821,N_29725);
nand UO_789 (O_789,N_29941,N_29840);
nand UO_790 (O_790,N_29706,N_29792);
xor UO_791 (O_791,N_29759,N_29757);
nand UO_792 (O_792,N_29701,N_29752);
or UO_793 (O_793,N_29960,N_29846);
xor UO_794 (O_794,N_29891,N_29845);
and UO_795 (O_795,N_29703,N_29992);
xnor UO_796 (O_796,N_29989,N_29727);
xor UO_797 (O_797,N_29981,N_29906);
nand UO_798 (O_798,N_29701,N_29852);
nand UO_799 (O_799,N_29719,N_29830);
xnor UO_800 (O_800,N_29858,N_29929);
and UO_801 (O_801,N_29792,N_29812);
or UO_802 (O_802,N_29968,N_29899);
or UO_803 (O_803,N_29909,N_29895);
and UO_804 (O_804,N_29810,N_29735);
xor UO_805 (O_805,N_29892,N_29886);
and UO_806 (O_806,N_29741,N_29703);
nor UO_807 (O_807,N_29816,N_29795);
xor UO_808 (O_808,N_29736,N_29720);
and UO_809 (O_809,N_29918,N_29844);
nor UO_810 (O_810,N_29845,N_29737);
or UO_811 (O_811,N_29724,N_29876);
or UO_812 (O_812,N_29766,N_29784);
nand UO_813 (O_813,N_29843,N_29716);
nor UO_814 (O_814,N_29920,N_29987);
and UO_815 (O_815,N_29718,N_29830);
or UO_816 (O_816,N_29857,N_29991);
nor UO_817 (O_817,N_29990,N_29729);
or UO_818 (O_818,N_29750,N_29989);
xnor UO_819 (O_819,N_29754,N_29782);
or UO_820 (O_820,N_29761,N_29781);
nand UO_821 (O_821,N_29878,N_29844);
nor UO_822 (O_822,N_29990,N_29777);
or UO_823 (O_823,N_29921,N_29766);
nor UO_824 (O_824,N_29798,N_29729);
or UO_825 (O_825,N_29715,N_29899);
nand UO_826 (O_826,N_29938,N_29906);
or UO_827 (O_827,N_29981,N_29776);
xnor UO_828 (O_828,N_29776,N_29767);
nand UO_829 (O_829,N_29822,N_29992);
xnor UO_830 (O_830,N_29759,N_29751);
and UO_831 (O_831,N_29798,N_29939);
nand UO_832 (O_832,N_29701,N_29707);
and UO_833 (O_833,N_29741,N_29783);
or UO_834 (O_834,N_29730,N_29723);
or UO_835 (O_835,N_29890,N_29792);
or UO_836 (O_836,N_29947,N_29901);
or UO_837 (O_837,N_29749,N_29786);
nor UO_838 (O_838,N_29764,N_29717);
nand UO_839 (O_839,N_29718,N_29859);
and UO_840 (O_840,N_29816,N_29856);
nand UO_841 (O_841,N_29954,N_29800);
nand UO_842 (O_842,N_29921,N_29738);
nor UO_843 (O_843,N_29728,N_29909);
nor UO_844 (O_844,N_29960,N_29790);
nor UO_845 (O_845,N_29760,N_29946);
and UO_846 (O_846,N_29933,N_29795);
nor UO_847 (O_847,N_29745,N_29971);
xor UO_848 (O_848,N_29727,N_29710);
xnor UO_849 (O_849,N_29756,N_29858);
and UO_850 (O_850,N_29923,N_29785);
xor UO_851 (O_851,N_29894,N_29821);
xor UO_852 (O_852,N_29867,N_29917);
nand UO_853 (O_853,N_29978,N_29961);
nand UO_854 (O_854,N_29830,N_29767);
nand UO_855 (O_855,N_29852,N_29821);
xor UO_856 (O_856,N_29867,N_29737);
nor UO_857 (O_857,N_29923,N_29928);
or UO_858 (O_858,N_29748,N_29886);
or UO_859 (O_859,N_29963,N_29747);
xnor UO_860 (O_860,N_29803,N_29836);
xor UO_861 (O_861,N_29924,N_29941);
xor UO_862 (O_862,N_29936,N_29901);
nor UO_863 (O_863,N_29966,N_29863);
and UO_864 (O_864,N_29818,N_29866);
nor UO_865 (O_865,N_29859,N_29840);
nand UO_866 (O_866,N_29731,N_29794);
nand UO_867 (O_867,N_29837,N_29971);
nand UO_868 (O_868,N_29861,N_29934);
nand UO_869 (O_869,N_29808,N_29866);
nor UO_870 (O_870,N_29993,N_29973);
and UO_871 (O_871,N_29769,N_29778);
xor UO_872 (O_872,N_29967,N_29713);
or UO_873 (O_873,N_29806,N_29924);
and UO_874 (O_874,N_29979,N_29929);
or UO_875 (O_875,N_29873,N_29902);
nor UO_876 (O_876,N_29928,N_29967);
nand UO_877 (O_877,N_29874,N_29802);
or UO_878 (O_878,N_29853,N_29743);
and UO_879 (O_879,N_29779,N_29895);
or UO_880 (O_880,N_29828,N_29843);
nand UO_881 (O_881,N_29726,N_29781);
nand UO_882 (O_882,N_29715,N_29905);
nor UO_883 (O_883,N_29811,N_29972);
nor UO_884 (O_884,N_29767,N_29700);
or UO_885 (O_885,N_29880,N_29877);
nand UO_886 (O_886,N_29721,N_29892);
and UO_887 (O_887,N_29976,N_29847);
nor UO_888 (O_888,N_29877,N_29909);
xnor UO_889 (O_889,N_29946,N_29909);
nand UO_890 (O_890,N_29887,N_29707);
or UO_891 (O_891,N_29902,N_29750);
xnor UO_892 (O_892,N_29873,N_29984);
xor UO_893 (O_893,N_29722,N_29898);
nor UO_894 (O_894,N_29846,N_29824);
xnor UO_895 (O_895,N_29860,N_29884);
and UO_896 (O_896,N_29769,N_29750);
xor UO_897 (O_897,N_29870,N_29763);
nor UO_898 (O_898,N_29870,N_29903);
nor UO_899 (O_899,N_29963,N_29841);
xnor UO_900 (O_900,N_29894,N_29745);
or UO_901 (O_901,N_29992,N_29937);
xor UO_902 (O_902,N_29759,N_29917);
nor UO_903 (O_903,N_29830,N_29985);
and UO_904 (O_904,N_29700,N_29892);
xnor UO_905 (O_905,N_29890,N_29773);
nor UO_906 (O_906,N_29837,N_29788);
nand UO_907 (O_907,N_29942,N_29947);
and UO_908 (O_908,N_29892,N_29820);
nand UO_909 (O_909,N_29931,N_29846);
nand UO_910 (O_910,N_29758,N_29941);
and UO_911 (O_911,N_29781,N_29993);
xor UO_912 (O_912,N_29974,N_29994);
nor UO_913 (O_913,N_29772,N_29960);
nand UO_914 (O_914,N_29953,N_29748);
xnor UO_915 (O_915,N_29799,N_29793);
or UO_916 (O_916,N_29756,N_29723);
and UO_917 (O_917,N_29905,N_29729);
or UO_918 (O_918,N_29769,N_29802);
or UO_919 (O_919,N_29985,N_29910);
nor UO_920 (O_920,N_29762,N_29721);
or UO_921 (O_921,N_29893,N_29883);
and UO_922 (O_922,N_29749,N_29787);
nand UO_923 (O_923,N_29720,N_29938);
nand UO_924 (O_924,N_29955,N_29832);
nor UO_925 (O_925,N_29796,N_29862);
xnor UO_926 (O_926,N_29844,N_29842);
xnor UO_927 (O_927,N_29781,N_29950);
xor UO_928 (O_928,N_29799,N_29865);
and UO_929 (O_929,N_29817,N_29806);
xor UO_930 (O_930,N_29847,N_29937);
or UO_931 (O_931,N_29924,N_29898);
nand UO_932 (O_932,N_29832,N_29847);
nor UO_933 (O_933,N_29777,N_29874);
nor UO_934 (O_934,N_29818,N_29968);
xnor UO_935 (O_935,N_29955,N_29771);
nand UO_936 (O_936,N_29814,N_29907);
xor UO_937 (O_937,N_29926,N_29852);
or UO_938 (O_938,N_29850,N_29785);
xor UO_939 (O_939,N_29842,N_29981);
nand UO_940 (O_940,N_29923,N_29752);
xor UO_941 (O_941,N_29787,N_29938);
nand UO_942 (O_942,N_29962,N_29926);
and UO_943 (O_943,N_29702,N_29740);
nor UO_944 (O_944,N_29799,N_29788);
or UO_945 (O_945,N_29926,N_29700);
xnor UO_946 (O_946,N_29712,N_29775);
and UO_947 (O_947,N_29969,N_29756);
nand UO_948 (O_948,N_29749,N_29907);
nor UO_949 (O_949,N_29780,N_29709);
nor UO_950 (O_950,N_29831,N_29983);
and UO_951 (O_951,N_29893,N_29867);
nor UO_952 (O_952,N_29841,N_29753);
nand UO_953 (O_953,N_29792,N_29848);
and UO_954 (O_954,N_29741,N_29868);
or UO_955 (O_955,N_29812,N_29867);
nand UO_956 (O_956,N_29780,N_29839);
xnor UO_957 (O_957,N_29828,N_29762);
nor UO_958 (O_958,N_29717,N_29882);
nor UO_959 (O_959,N_29753,N_29909);
and UO_960 (O_960,N_29874,N_29927);
or UO_961 (O_961,N_29871,N_29958);
xnor UO_962 (O_962,N_29852,N_29931);
and UO_963 (O_963,N_29840,N_29905);
nand UO_964 (O_964,N_29815,N_29819);
nand UO_965 (O_965,N_29765,N_29783);
or UO_966 (O_966,N_29706,N_29846);
or UO_967 (O_967,N_29755,N_29849);
nor UO_968 (O_968,N_29805,N_29763);
xor UO_969 (O_969,N_29901,N_29896);
and UO_970 (O_970,N_29813,N_29739);
and UO_971 (O_971,N_29898,N_29863);
nor UO_972 (O_972,N_29764,N_29807);
nor UO_973 (O_973,N_29814,N_29837);
and UO_974 (O_974,N_29934,N_29901);
nand UO_975 (O_975,N_29927,N_29711);
and UO_976 (O_976,N_29804,N_29825);
nor UO_977 (O_977,N_29915,N_29759);
xor UO_978 (O_978,N_29880,N_29759);
or UO_979 (O_979,N_29824,N_29843);
nand UO_980 (O_980,N_29947,N_29860);
nand UO_981 (O_981,N_29960,N_29880);
or UO_982 (O_982,N_29913,N_29918);
or UO_983 (O_983,N_29965,N_29841);
or UO_984 (O_984,N_29749,N_29998);
nand UO_985 (O_985,N_29868,N_29781);
nor UO_986 (O_986,N_29807,N_29821);
nand UO_987 (O_987,N_29984,N_29939);
or UO_988 (O_988,N_29866,N_29722);
and UO_989 (O_989,N_29780,N_29985);
or UO_990 (O_990,N_29785,N_29974);
or UO_991 (O_991,N_29722,N_29795);
or UO_992 (O_992,N_29861,N_29929);
or UO_993 (O_993,N_29981,N_29724);
nand UO_994 (O_994,N_29711,N_29764);
nand UO_995 (O_995,N_29820,N_29834);
nand UO_996 (O_996,N_29971,N_29926);
nand UO_997 (O_997,N_29717,N_29724);
or UO_998 (O_998,N_29761,N_29807);
and UO_999 (O_999,N_29867,N_29701);
or UO_1000 (O_1000,N_29851,N_29731);
or UO_1001 (O_1001,N_29947,N_29713);
and UO_1002 (O_1002,N_29732,N_29938);
or UO_1003 (O_1003,N_29812,N_29782);
nor UO_1004 (O_1004,N_29864,N_29946);
or UO_1005 (O_1005,N_29769,N_29996);
nand UO_1006 (O_1006,N_29891,N_29992);
and UO_1007 (O_1007,N_29731,N_29850);
and UO_1008 (O_1008,N_29798,N_29706);
nand UO_1009 (O_1009,N_29932,N_29725);
or UO_1010 (O_1010,N_29872,N_29700);
or UO_1011 (O_1011,N_29766,N_29930);
or UO_1012 (O_1012,N_29996,N_29790);
and UO_1013 (O_1013,N_29872,N_29756);
nand UO_1014 (O_1014,N_29790,N_29711);
xnor UO_1015 (O_1015,N_29715,N_29970);
or UO_1016 (O_1016,N_29726,N_29968);
and UO_1017 (O_1017,N_29828,N_29944);
or UO_1018 (O_1018,N_29713,N_29817);
xor UO_1019 (O_1019,N_29724,N_29927);
and UO_1020 (O_1020,N_29870,N_29854);
nand UO_1021 (O_1021,N_29765,N_29780);
nor UO_1022 (O_1022,N_29726,N_29793);
or UO_1023 (O_1023,N_29907,N_29768);
or UO_1024 (O_1024,N_29964,N_29864);
xor UO_1025 (O_1025,N_29916,N_29735);
or UO_1026 (O_1026,N_29934,N_29762);
or UO_1027 (O_1027,N_29846,N_29742);
and UO_1028 (O_1028,N_29750,N_29758);
or UO_1029 (O_1029,N_29718,N_29921);
nand UO_1030 (O_1030,N_29942,N_29937);
xnor UO_1031 (O_1031,N_29879,N_29952);
and UO_1032 (O_1032,N_29943,N_29938);
and UO_1033 (O_1033,N_29898,N_29926);
xor UO_1034 (O_1034,N_29706,N_29801);
or UO_1035 (O_1035,N_29785,N_29744);
and UO_1036 (O_1036,N_29963,N_29789);
and UO_1037 (O_1037,N_29923,N_29742);
nand UO_1038 (O_1038,N_29760,N_29929);
or UO_1039 (O_1039,N_29706,N_29932);
nand UO_1040 (O_1040,N_29729,N_29922);
nand UO_1041 (O_1041,N_29925,N_29835);
nor UO_1042 (O_1042,N_29974,N_29763);
or UO_1043 (O_1043,N_29843,N_29845);
nor UO_1044 (O_1044,N_29750,N_29751);
xnor UO_1045 (O_1045,N_29721,N_29999);
or UO_1046 (O_1046,N_29819,N_29934);
and UO_1047 (O_1047,N_29970,N_29794);
nand UO_1048 (O_1048,N_29700,N_29779);
or UO_1049 (O_1049,N_29721,N_29822);
xor UO_1050 (O_1050,N_29773,N_29795);
xor UO_1051 (O_1051,N_29850,N_29810);
xnor UO_1052 (O_1052,N_29981,N_29732);
and UO_1053 (O_1053,N_29932,N_29913);
and UO_1054 (O_1054,N_29893,N_29700);
xor UO_1055 (O_1055,N_29956,N_29967);
nor UO_1056 (O_1056,N_29893,N_29702);
nand UO_1057 (O_1057,N_29962,N_29717);
nor UO_1058 (O_1058,N_29921,N_29906);
or UO_1059 (O_1059,N_29834,N_29904);
nor UO_1060 (O_1060,N_29795,N_29985);
and UO_1061 (O_1061,N_29917,N_29840);
nor UO_1062 (O_1062,N_29784,N_29797);
xnor UO_1063 (O_1063,N_29968,N_29940);
and UO_1064 (O_1064,N_29906,N_29956);
nand UO_1065 (O_1065,N_29700,N_29930);
or UO_1066 (O_1066,N_29828,N_29750);
or UO_1067 (O_1067,N_29865,N_29793);
xnor UO_1068 (O_1068,N_29973,N_29755);
nor UO_1069 (O_1069,N_29792,N_29838);
and UO_1070 (O_1070,N_29731,N_29828);
nor UO_1071 (O_1071,N_29967,N_29973);
nor UO_1072 (O_1072,N_29970,N_29762);
xor UO_1073 (O_1073,N_29934,N_29764);
nor UO_1074 (O_1074,N_29855,N_29941);
nor UO_1075 (O_1075,N_29776,N_29916);
nor UO_1076 (O_1076,N_29813,N_29941);
or UO_1077 (O_1077,N_29939,N_29894);
nor UO_1078 (O_1078,N_29862,N_29783);
nor UO_1079 (O_1079,N_29721,N_29964);
xor UO_1080 (O_1080,N_29787,N_29862);
and UO_1081 (O_1081,N_29965,N_29907);
or UO_1082 (O_1082,N_29718,N_29775);
nor UO_1083 (O_1083,N_29719,N_29773);
and UO_1084 (O_1084,N_29960,N_29889);
nand UO_1085 (O_1085,N_29939,N_29993);
nor UO_1086 (O_1086,N_29939,N_29936);
and UO_1087 (O_1087,N_29902,N_29746);
xnor UO_1088 (O_1088,N_29785,N_29718);
xor UO_1089 (O_1089,N_29786,N_29704);
nand UO_1090 (O_1090,N_29893,N_29746);
and UO_1091 (O_1091,N_29910,N_29935);
xnor UO_1092 (O_1092,N_29930,N_29887);
or UO_1093 (O_1093,N_29816,N_29941);
nand UO_1094 (O_1094,N_29887,N_29823);
nor UO_1095 (O_1095,N_29827,N_29952);
nand UO_1096 (O_1096,N_29872,N_29844);
nand UO_1097 (O_1097,N_29860,N_29908);
nor UO_1098 (O_1098,N_29856,N_29952);
nand UO_1099 (O_1099,N_29883,N_29906);
and UO_1100 (O_1100,N_29989,N_29763);
and UO_1101 (O_1101,N_29708,N_29843);
nand UO_1102 (O_1102,N_29734,N_29819);
or UO_1103 (O_1103,N_29725,N_29883);
nand UO_1104 (O_1104,N_29919,N_29808);
and UO_1105 (O_1105,N_29772,N_29809);
and UO_1106 (O_1106,N_29763,N_29806);
and UO_1107 (O_1107,N_29775,N_29969);
or UO_1108 (O_1108,N_29884,N_29997);
or UO_1109 (O_1109,N_29738,N_29843);
or UO_1110 (O_1110,N_29993,N_29851);
xor UO_1111 (O_1111,N_29731,N_29736);
and UO_1112 (O_1112,N_29825,N_29904);
nor UO_1113 (O_1113,N_29918,N_29910);
xor UO_1114 (O_1114,N_29971,N_29832);
nand UO_1115 (O_1115,N_29977,N_29818);
and UO_1116 (O_1116,N_29955,N_29712);
xor UO_1117 (O_1117,N_29999,N_29892);
xnor UO_1118 (O_1118,N_29740,N_29948);
nand UO_1119 (O_1119,N_29964,N_29934);
xor UO_1120 (O_1120,N_29919,N_29814);
or UO_1121 (O_1121,N_29707,N_29749);
xor UO_1122 (O_1122,N_29965,N_29793);
nand UO_1123 (O_1123,N_29790,N_29776);
xor UO_1124 (O_1124,N_29899,N_29921);
and UO_1125 (O_1125,N_29781,N_29778);
nand UO_1126 (O_1126,N_29835,N_29918);
nor UO_1127 (O_1127,N_29995,N_29963);
xor UO_1128 (O_1128,N_29790,N_29821);
nor UO_1129 (O_1129,N_29787,N_29822);
nor UO_1130 (O_1130,N_29708,N_29806);
or UO_1131 (O_1131,N_29761,N_29768);
nand UO_1132 (O_1132,N_29709,N_29950);
nor UO_1133 (O_1133,N_29848,N_29999);
nor UO_1134 (O_1134,N_29805,N_29882);
nand UO_1135 (O_1135,N_29868,N_29723);
nor UO_1136 (O_1136,N_29788,N_29781);
and UO_1137 (O_1137,N_29881,N_29840);
xnor UO_1138 (O_1138,N_29964,N_29926);
nand UO_1139 (O_1139,N_29986,N_29847);
and UO_1140 (O_1140,N_29826,N_29737);
or UO_1141 (O_1141,N_29731,N_29976);
or UO_1142 (O_1142,N_29852,N_29930);
and UO_1143 (O_1143,N_29988,N_29737);
nand UO_1144 (O_1144,N_29814,N_29802);
and UO_1145 (O_1145,N_29974,N_29850);
nor UO_1146 (O_1146,N_29976,N_29728);
nor UO_1147 (O_1147,N_29764,N_29769);
nor UO_1148 (O_1148,N_29782,N_29716);
and UO_1149 (O_1149,N_29993,N_29810);
nor UO_1150 (O_1150,N_29838,N_29876);
nor UO_1151 (O_1151,N_29946,N_29869);
nand UO_1152 (O_1152,N_29883,N_29966);
xor UO_1153 (O_1153,N_29927,N_29823);
nor UO_1154 (O_1154,N_29991,N_29809);
nor UO_1155 (O_1155,N_29812,N_29791);
nand UO_1156 (O_1156,N_29783,N_29807);
nor UO_1157 (O_1157,N_29870,N_29853);
or UO_1158 (O_1158,N_29761,N_29737);
xnor UO_1159 (O_1159,N_29922,N_29973);
nor UO_1160 (O_1160,N_29975,N_29721);
xor UO_1161 (O_1161,N_29869,N_29888);
and UO_1162 (O_1162,N_29867,N_29836);
or UO_1163 (O_1163,N_29710,N_29732);
and UO_1164 (O_1164,N_29886,N_29995);
nor UO_1165 (O_1165,N_29817,N_29703);
nand UO_1166 (O_1166,N_29950,N_29762);
or UO_1167 (O_1167,N_29994,N_29741);
xor UO_1168 (O_1168,N_29929,N_29732);
nand UO_1169 (O_1169,N_29953,N_29738);
xnor UO_1170 (O_1170,N_29835,N_29744);
and UO_1171 (O_1171,N_29932,N_29921);
and UO_1172 (O_1172,N_29830,N_29991);
and UO_1173 (O_1173,N_29798,N_29938);
xor UO_1174 (O_1174,N_29732,N_29829);
xnor UO_1175 (O_1175,N_29787,N_29813);
or UO_1176 (O_1176,N_29802,N_29733);
and UO_1177 (O_1177,N_29803,N_29730);
and UO_1178 (O_1178,N_29862,N_29822);
xor UO_1179 (O_1179,N_29961,N_29751);
nand UO_1180 (O_1180,N_29736,N_29860);
nor UO_1181 (O_1181,N_29982,N_29995);
nor UO_1182 (O_1182,N_29858,N_29916);
or UO_1183 (O_1183,N_29997,N_29875);
nor UO_1184 (O_1184,N_29833,N_29997);
nor UO_1185 (O_1185,N_29894,N_29879);
nand UO_1186 (O_1186,N_29716,N_29986);
nand UO_1187 (O_1187,N_29730,N_29721);
nand UO_1188 (O_1188,N_29713,N_29893);
nor UO_1189 (O_1189,N_29950,N_29979);
or UO_1190 (O_1190,N_29723,N_29797);
xor UO_1191 (O_1191,N_29755,N_29877);
xnor UO_1192 (O_1192,N_29935,N_29709);
xor UO_1193 (O_1193,N_29915,N_29879);
xnor UO_1194 (O_1194,N_29731,N_29764);
and UO_1195 (O_1195,N_29997,N_29980);
or UO_1196 (O_1196,N_29802,N_29766);
nand UO_1197 (O_1197,N_29786,N_29964);
nand UO_1198 (O_1198,N_29981,N_29946);
nor UO_1199 (O_1199,N_29782,N_29829);
or UO_1200 (O_1200,N_29808,N_29959);
or UO_1201 (O_1201,N_29729,N_29852);
xor UO_1202 (O_1202,N_29796,N_29799);
xor UO_1203 (O_1203,N_29937,N_29901);
nand UO_1204 (O_1204,N_29799,N_29851);
nand UO_1205 (O_1205,N_29741,N_29811);
nand UO_1206 (O_1206,N_29755,N_29763);
nor UO_1207 (O_1207,N_29885,N_29737);
and UO_1208 (O_1208,N_29946,N_29865);
nor UO_1209 (O_1209,N_29731,N_29779);
nor UO_1210 (O_1210,N_29776,N_29938);
xnor UO_1211 (O_1211,N_29933,N_29826);
or UO_1212 (O_1212,N_29818,N_29853);
nor UO_1213 (O_1213,N_29807,N_29985);
and UO_1214 (O_1214,N_29783,N_29799);
nand UO_1215 (O_1215,N_29853,N_29729);
nor UO_1216 (O_1216,N_29836,N_29942);
or UO_1217 (O_1217,N_29872,N_29782);
nor UO_1218 (O_1218,N_29952,N_29853);
xor UO_1219 (O_1219,N_29807,N_29840);
nand UO_1220 (O_1220,N_29752,N_29964);
nor UO_1221 (O_1221,N_29758,N_29722);
or UO_1222 (O_1222,N_29803,N_29900);
xor UO_1223 (O_1223,N_29879,N_29785);
or UO_1224 (O_1224,N_29707,N_29708);
nand UO_1225 (O_1225,N_29827,N_29792);
xnor UO_1226 (O_1226,N_29918,N_29942);
or UO_1227 (O_1227,N_29996,N_29727);
nor UO_1228 (O_1228,N_29851,N_29787);
xor UO_1229 (O_1229,N_29843,N_29901);
nor UO_1230 (O_1230,N_29715,N_29727);
xor UO_1231 (O_1231,N_29800,N_29930);
xnor UO_1232 (O_1232,N_29957,N_29891);
and UO_1233 (O_1233,N_29761,N_29845);
nor UO_1234 (O_1234,N_29908,N_29932);
xor UO_1235 (O_1235,N_29778,N_29745);
xor UO_1236 (O_1236,N_29855,N_29972);
xnor UO_1237 (O_1237,N_29946,N_29806);
nand UO_1238 (O_1238,N_29760,N_29965);
xor UO_1239 (O_1239,N_29944,N_29878);
xor UO_1240 (O_1240,N_29811,N_29796);
xnor UO_1241 (O_1241,N_29730,N_29760);
nor UO_1242 (O_1242,N_29754,N_29981);
xnor UO_1243 (O_1243,N_29902,N_29831);
xnor UO_1244 (O_1244,N_29747,N_29850);
nand UO_1245 (O_1245,N_29739,N_29966);
and UO_1246 (O_1246,N_29741,N_29792);
xor UO_1247 (O_1247,N_29979,N_29957);
nor UO_1248 (O_1248,N_29998,N_29805);
or UO_1249 (O_1249,N_29828,N_29751);
nor UO_1250 (O_1250,N_29767,N_29845);
nand UO_1251 (O_1251,N_29815,N_29722);
nand UO_1252 (O_1252,N_29847,N_29714);
and UO_1253 (O_1253,N_29860,N_29936);
nand UO_1254 (O_1254,N_29730,N_29823);
nor UO_1255 (O_1255,N_29861,N_29806);
nor UO_1256 (O_1256,N_29784,N_29836);
nand UO_1257 (O_1257,N_29925,N_29883);
nor UO_1258 (O_1258,N_29877,N_29857);
nand UO_1259 (O_1259,N_29830,N_29989);
or UO_1260 (O_1260,N_29748,N_29992);
nor UO_1261 (O_1261,N_29843,N_29836);
or UO_1262 (O_1262,N_29741,N_29728);
xor UO_1263 (O_1263,N_29864,N_29831);
xor UO_1264 (O_1264,N_29752,N_29837);
and UO_1265 (O_1265,N_29804,N_29773);
xnor UO_1266 (O_1266,N_29822,N_29964);
and UO_1267 (O_1267,N_29878,N_29980);
nor UO_1268 (O_1268,N_29777,N_29957);
nand UO_1269 (O_1269,N_29902,N_29976);
xnor UO_1270 (O_1270,N_29915,N_29705);
nor UO_1271 (O_1271,N_29936,N_29745);
nand UO_1272 (O_1272,N_29747,N_29724);
and UO_1273 (O_1273,N_29940,N_29793);
and UO_1274 (O_1274,N_29857,N_29821);
and UO_1275 (O_1275,N_29891,N_29770);
nand UO_1276 (O_1276,N_29756,N_29850);
nand UO_1277 (O_1277,N_29735,N_29796);
nand UO_1278 (O_1278,N_29768,N_29829);
or UO_1279 (O_1279,N_29898,N_29812);
nor UO_1280 (O_1280,N_29817,N_29877);
or UO_1281 (O_1281,N_29889,N_29760);
xnor UO_1282 (O_1282,N_29846,N_29975);
or UO_1283 (O_1283,N_29922,N_29995);
nand UO_1284 (O_1284,N_29964,N_29826);
xnor UO_1285 (O_1285,N_29870,N_29791);
and UO_1286 (O_1286,N_29743,N_29979);
or UO_1287 (O_1287,N_29735,N_29882);
nor UO_1288 (O_1288,N_29960,N_29710);
nand UO_1289 (O_1289,N_29791,N_29744);
or UO_1290 (O_1290,N_29834,N_29781);
nand UO_1291 (O_1291,N_29949,N_29758);
and UO_1292 (O_1292,N_29977,N_29729);
or UO_1293 (O_1293,N_29739,N_29775);
nand UO_1294 (O_1294,N_29919,N_29925);
or UO_1295 (O_1295,N_29724,N_29946);
nor UO_1296 (O_1296,N_29817,N_29935);
xnor UO_1297 (O_1297,N_29994,N_29993);
nor UO_1298 (O_1298,N_29741,N_29854);
or UO_1299 (O_1299,N_29905,N_29767);
nor UO_1300 (O_1300,N_29707,N_29852);
xnor UO_1301 (O_1301,N_29785,N_29848);
xor UO_1302 (O_1302,N_29936,N_29970);
and UO_1303 (O_1303,N_29724,N_29805);
and UO_1304 (O_1304,N_29951,N_29956);
nand UO_1305 (O_1305,N_29758,N_29762);
xor UO_1306 (O_1306,N_29997,N_29773);
nand UO_1307 (O_1307,N_29716,N_29788);
or UO_1308 (O_1308,N_29935,N_29933);
nor UO_1309 (O_1309,N_29729,N_29704);
and UO_1310 (O_1310,N_29805,N_29925);
nor UO_1311 (O_1311,N_29766,N_29911);
or UO_1312 (O_1312,N_29868,N_29747);
nor UO_1313 (O_1313,N_29761,N_29922);
xor UO_1314 (O_1314,N_29982,N_29994);
xor UO_1315 (O_1315,N_29901,N_29836);
nor UO_1316 (O_1316,N_29833,N_29919);
or UO_1317 (O_1317,N_29861,N_29700);
nand UO_1318 (O_1318,N_29880,N_29971);
xnor UO_1319 (O_1319,N_29938,N_29850);
xnor UO_1320 (O_1320,N_29792,N_29715);
and UO_1321 (O_1321,N_29953,N_29888);
or UO_1322 (O_1322,N_29833,N_29810);
xor UO_1323 (O_1323,N_29736,N_29760);
nor UO_1324 (O_1324,N_29999,N_29937);
nand UO_1325 (O_1325,N_29952,N_29755);
nor UO_1326 (O_1326,N_29852,N_29999);
xnor UO_1327 (O_1327,N_29888,N_29719);
and UO_1328 (O_1328,N_29841,N_29887);
and UO_1329 (O_1329,N_29819,N_29925);
and UO_1330 (O_1330,N_29800,N_29776);
and UO_1331 (O_1331,N_29844,N_29781);
and UO_1332 (O_1332,N_29956,N_29710);
and UO_1333 (O_1333,N_29977,N_29777);
nor UO_1334 (O_1334,N_29817,N_29878);
and UO_1335 (O_1335,N_29985,N_29967);
nand UO_1336 (O_1336,N_29739,N_29714);
xor UO_1337 (O_1337,N_29825,N_29958);
nand UO_1338 (O_1338,N_29937,N_29990);
and UO_1339 (O_1339,N_29879,N_29853);
or UO_1340 (O_1340,N_29847,N_29912);
xnor UO_1341 (O_1341,N_29995,N_29728);
nor UO_1342 (O_1342,N_29727,N_29981);
or UO_1343 (O_1343,N_29963,N_29739);
nor UO_1344 (O_1344,N_29808,N_29981);
nand UO_1345 (O_1345,N_29948,N_29946);
nor UO_1346 (O_1346,N_29771,N_29743);
or UO_1347 (O_1347,N_29709,N_29715);
nand UO_1348 (O_1348,N_29925,N_29803);
and UO_1349 (O_1349,N_29961,N_29859);
nor UO_1350 (O_1350,N_29951,N_29800);
and UO_1351 (O_1351,N_29941,N_29913);
and UO_1352 (O_1352,N_29966,N_29816);
or UO_1353 (O_1353,N_29732,N_29890);
nor UO_1354 (O_1354,N_29868,N_29703);
xnor UO_1355 (O_1355,N_29812,N_29746);
nor UO_1356 (O_1356,N_29804,N_29878);
xor UO_1357 (O_1357,N_29932,N_29930);
xnor UO_1358 (O_1358,N_29735,N_29946);
and UO_1359 (O_1359,N_29706,N_29873);
xor UO_1360 (O_1360,N_29888,N_29838);
nor UO_1361 (O_1361,N_29973,N_29760);
nor UO_1362 (O_1362,N_29812,N_29999);
or UO_1363 (O_1363,N_29769,N_29746);
or UO_1364 (O_1364,N_29967,N_29853);
or UO_1365 (O_1365,N_29705,N_29850);
nor UO_1366 (O_1366,N_29827,N_29913);
nand UO_1367 (O_1367,N_29983,N_29786);
or UO_1368 (O_1368,N_29782,N_29821);
or UO_1369 (O_1369,N_29745,N_29815);
nand UO_1370 (O_1370,N_29794,N_29932);
nor UO_1371 (O_1371,N_29853,N_29830);
or UO_1372 (O_1372,N_29774,N_29752);
and UO_1373 (O_1373,N_29964,N_29987);
nor UO_1374 (O_1374,N_29930,N_29785);
nand UO_1375 (O_1375,N_29859,N_29951);
or UO_1376 (O_1376,N_29852,N_29879);
nor UO_1377 (O_1377,N_29800,N_29809);
nor UO_1378 (O_1378,N_29969,N_29934);
nand UO_1379 (O_1379,N_29757,N_29920);
nor UO_1380 (O_1380,N_29950,N_29891);
and UO_1381 (O_1381,N_29767,N_29896);
nor UO_1382 (O_1382,N_29770,N_29700);
or UO_1383 (O_1383,N_29804,N_29988);
nand UO_1384 (O_1384,N_29954,N_29774);
nor UO_1385 (O_1385,N_29876,N_29757);
and UO_1386 (O_1386,N_29703,N_29818);
nor UO_1387 (O_1387,N_29777,N_29998);
xnor UO_1388 (O_1388,N_29962,N_29932);
xnor UO_1389 (O_1389,N_29963,N_29724);
xnor UO_1390 (O_1390,N_29952,N_29818);
and UO_1391 (O_1391,N_29830,N_29860);
nand UO_1392 (O_1392,N_29754,N_29865);
nand UO_1393 (O_1393,N_29867,N_29899);
nor UO_1394 (O_1394,N_29829,N_29952);
nand UO_1395 (O_1395,N_29736,N_29807);
or UO_1396 (O_1396,N_29816,N_29894);
nand UO_1397 (O_1397,N_29724,N_29851);
xnor UO_1398 (O_1398,N_29994,N_29778);
xnor UO_1399 (O_1399,N_29878,N_29872);
nand UO_1400 (O_1400,N_29724,N_29881);
nor UO_1401 (O_1401,N_29711,N_29878);
nand UO_1402 (O_1402,N_29857,N_29976);
and UO_1403 (O_1403,N_29782,N_29892);
or UO_1404 (O_1404,N_29945,N_29989);
and UO_1405 (O_1405,N_29860,N_29713);
nor UO_1406 (O_1406,N_29801,N_29734);
and UO_1407 (O_1407,N_29862,N_29981);
nor UO_1408 (O_1408,N_29965,N_29947);
or UO_1409 (O_1409,N_29707,N_29962);
nand UO_1410 (O_1410,N_29818,N_29993);
xor UO_1411 (O_1411,N_29950,N_29922);
nor UO_1412 (O_1412,N_29929,N_29725);
nor UO_1413 (O_1413,N_29902,N_29703);
nor UO_1414 (O_1414,N_29767,N_29852);
xnor UO_1415 (O_1415,N_29771,N_29948);
and UO_1416 (O_1416,N_29918,N_29791);
and UO_1417 (O_1417,N_29872,N_29715);
or UO_1418 (O_1418,N_29784,N_29968);
and UO_1419 (O_1419,N_29717,N_29749);
xnor UO_1420 (O_1420,N_29726,N_29721);
nand UO_1421 (O_1421,N_29921,N_29767);
and UO_1422 (O_1422,N_29845,N_29728);
nor UO_1423 (O_1423,N_29801,N_29940);
nor UO_1424 (O_1424,N_29934,N_29739);
nand UO_1425 (O_1425,N_29707,N_29734);
or UO_1426 (O_1426,N_29766,N_29708);
and UO_1427 (O_1427,N_29808,N_29746);
xor UO_1428 (O_1428,N_29833,N_29883);
nand UO_1429 (O_1429,N_29733,N_29933);
and UO_1430 (O_1430,N_29782,N_29733);
or UO_1431 (O_1431,N_29768,N_29847);
nand UO_1432 (O_1432,N_29801,N_29807);
nor UO_1433 (O_1433,N_29956,N_29839);
nor UO_1434 (O_1434,N_29808,N_29862);
nor UO_1435 (O_1435,N_29883,N_29868);
and UO_1436 (O_1436,N_29734,N_29767);
and UO_1437 (O_1437,N_29979,N_29815);
nand UO_1438 (O_1438,N_29926,N_29855);
xnor UO_1439 (O_1439,N_29748,N_29750);
nor UO_1440 (O_1440,N_29820,N_29956);
nand UO_1441 (O_1441,N_29873,N_29965);
or UO_1442 (O_1442,N_29801,N_29929);
and UO_1443 (O_1443,N_29741,N_29938);
nor UO_1444 (O_1444,N_29819,N_29774);
xor UO_1445 (O_1445,N_29965,N_29816);
and UO_1446 (O_1446,N_29741,N_29791);
nor UO_1447 (O_1447,N_29990,N_29772);
xor UO_1448 (O_1448,N_29746,N_29977);
nand UO_1449 (O_1449,N_29805,N_29865);
xor UO_1450 (O_1450,N_29869,N_29853);
xnor UO_1451 (O_1451,N_29944,N_29759);
nand UO_1452 (O_1452,N_29701,N_29898);
xnor UO_1453 (O_1453,N_29935,N_29769);
xnor UO_1454 (O_1454,N_29935,N_29779);
xor UO_1455 (O_1455,N_29911,N_29912);
or UO_1456 (O_1456,N_29818,N_29708);
and UO_1457 (O_1457,N_29800,N_29860);
and UO_1458 (O_1458,N_29747,N_29964);
or UO_1459 (O_1459,N_29908,N_29977);
nor UO_1460 (O_1460,N_29719,N_29700);
nor UO_1461 (O_1461,N_29901,N_29729);
xor UO_1462 (O_1462,N_29869,N_29822);
nand UO_1463 (O_1463,N_29876,N_29779);
nor UO_1464 (O_1464,N_29754,N_29931);
or UO_1465 (O_1465,N_29725,N_29980);
xor UO_1466 (O_1466,N_29978,N_29747);
or UO_1467 (O_1467,N_29756,N_29736);
xnor UO_1468 (O_1468,N_29708,N_29877);
xor UO_1469 (O_1469,N_29953,N_29819);
nand UO_1470 (O_1470,N_29838,N_29710);
nand UO_1471 (O_1471,N_29741,N_29734);
xor UO_1472 (O_1472,N_29855,N_29907);
nor UO_1473 (O_1473,N_29978,N_29948);
and UO_1474 (O_1474,N_29857,N_29839);
or UO_1475 (O_1475,N_29934,N_29810);
nand UO_1476 (O_1476,N_29888,N_29770);
or UO_1477 (O_1477,N_29785,N_29749);
nor UO_1478 (O_1478,N_29757,N_29742);
or UO_1479 (O_1479,N_29737,N_29937);
xnor UO_1480 (O_1480,N_29996,N_29923);
or UO_1481 (O_1481,N_29991,N_29982);
and UO_1482 (O_1482,N_29835,N_29960);
xor UO_1483 (O_1483,N_29711,N_29802);
nand UO_1484 (O_1484,N_29792,N_29730);
and UO_1485 (O_1485,N_29747,N_29876);
and UO_1486 (O_1486,N_29836,N_29953);
or UO_1487 (O_1487,N_29905,N_29849);
nand UO_1488 (O_1488,N_29919,N_29805);
nand UO_1489 (O_1489,N_29736,N_29784);
nand UO_1490 (O_1490,N_29855,N_29858);
nor UO_1491 (O_1491,N_29839,N_29777);
nand UO_1492 (O_1492,N_29721,N_29960);
or UO_1493 (O_1493,N_29916,N_29737);
xnor UO_1494 (O_1494,N_29835,N_29756);
xor UO_1495 (O_1495,N_29779,N_29919);
xnor UO_1496 (O_1496,N_29798,N_29732);
or UO_1497 (O_1497,N_29859,N_29797);
nand UO_1498 (O_1498,N_29832,N_29770);
xor UO_1499 (O_1499,N_29991,N_29865);
or UO_1500 (O_1500,N_29735,N_29745);
nand UO_1501 (O_1501,N_29982,N_29939);
nor UO_1502 (O_1502,N_29983,N_29776);
nor UO_1503 (O_1503,N_29997,N_29720);
or UO_1504 (O_1504,N_29996,N_29735);
nand UO_1505 (O_1505,N_29778,N_29944);
and UO_1506 (O_1506,N_29893,N_29938);
nand UO_1507 (O_1507,N_29994,N_29767);
xor UO_1508 (O_1508,N_29834,N_29933);
or UO_1509 (O_1509,N_29973,N_29961);
xor UO_1510 (O_1510,N_29923,N_29993);
nand UO_1511 (O_1511,N_29715,N_29783);
and UO_1512 (O_1512,N_29959,N_29765);
nand UO_1513 (O_1513,N_29807,N_29905);
and UO_1514 (O_1514,N_29818,N_29816);
nand UO_1515 (O_1515,N_29812,N_29817);
and UO_1516 (O_1516,N_29904,N_29731);
nand UO_1517 (O_1517,N_29791,N_29827);
and UO_1518 (O_1518,N_29747,N_29996);
or UO_1519 (O_1519,N_29726,N_29720);
nor UO_1520 (O_1520,N_29788,N_29707);
nand UO_1521 (O_1521,N_29910,N_29854);
and UO_1522 (O_1522,N_29987,N_29750);
xor UO_1523 (O_1523,N_29762,N_29854);
or UO_1524 (O_1524,N_29810,N_29774);
nor UO_1525 (O_1525,N_29895,N_29728);
xnor UO_1526 (O_1526,N_29996,N_29851);
nor UO_1527 (O_1527,N_29721,N_29840);
nand UO_1528 (O_1528,N_29712,N_29990);
nor UO_1529 (O_1529,N_29719,N_29752);
or UO_1530 (O_1530,N_29752,N_29891);
or UO_1531 (O_1531,N_29716,N_29852);
xnor UO_1532 (O_1532,N_29928,N_29822);
nand UO_1533 (O_1533,N_29945,N_29897);
xnor UO_1534 (O_1534,N_29912,N_29815);
nor UO_1535 (O_1535,N_29945,N_29783);
and UO_1536 (O_1536,N_29719,N_29994);
or UO_1537 (O_1537,N_29973,N_29820);
and UO_1538 (O_1538,N_29881,N_29795);
and UO_1539 (O_1539,N_29737,N_29950);
or UO_1540 (O_1540,N_29739,N_29869);
nor UO_1541 (O_1541,N_29754,N_29870);
nand UO_1542 (O_1542,N_29735,N_29907);
and UO_1543 (O_1543,N_29805,N_29729);
nor UO_1544 (O_1544,N_29753,N_29760);
xnor UO_1545 (O_1545,N_29996,N_29870);
and UO_1546 (O_1546,N_29936,N_29905);
or UO_1547 (O_1547,N_29894,N_29707);
and UO_1548 (O_1548,N_29946,N_29786);
nand UO_1549 (O_1549,N_29763,N_29821);
or UO_1550 (O_1550,N_29989,N_29807);
or UO_1551 (O_1551,N_29962,N_29897);
xor UO_1552 (O_1552,N_29922,N_29706);
xor UO_1553 (O_1553,N_29854,N_29927);
xnor UO_1554 (O_1554,N_29869,N_29771);
or UO_1555 (O_1555,N_29783,N_29894);
nor UO_1556 (O_1556,N_29968,N_29804);
nand UO_1557 (O_1557,N_29751,N_29798);
nand UO_1558 (O_1558,N_29855,N_29800);
nand UO_1559 (O_1559,N_29941,N_29934);
xnor UO_1560 (O_1560,N_29870,N_29786);
nor UO_1561 (O_1561,N_29970,N_29973);
or UO_1562 (O_1562,N_29941,N_29976);
nand UO_1563 (O_1563,N_29937,N_29895);
and UO_1564 (O_1564,N_29859,N_29780);
nor UO_1565 (O_1565,N_29799,N_29880);
and UO_1566 (O_1566,N_29775,N_29836);
or UO_1567 (O_1567,N_29736,N_29855);
or UO_1568 (O_1568,N_29787,N_29716);
or UO_1569 (O_1569,N_29956,N_29908);
nand UO_1570 (O_1570,N_29729,N_29891);
or UO_1571 (O_1571,N_29920,N_29816);
nand UO_1572 (O_1572,N_29880,N_29793);
nand UO_1573 (O_1573,N_29771,N_29938);
or UO_1574 (O_1574,N_29997,N_29751);
and UO_1575 (O_1575,N_29939,N_29930);
or UO_1576 (O_1576,N_29778,N_29969);
and UO_1577 (O_1577,N_29738,N_29735);
nor UO_1578 (O_1578,N_29919,N_29796);
nand UO_1579 (O_1579,N_29878,N_29723);
and UO_1580 (O_1580,N_29936,N_29808);
and UO_1581 (O_1581,N_29760,N_29764);
or UO_1582 (O_1582,N_29870,N_29756);
or UO_1583 (O_1583,N_29868,N_29876);
and UO_1584 (O_1584,N_29956,N_29913);
nor UO_1585 (O_1585,N_29746,N_29775);
nand UO_1586 (O_1586,N_29973,N_29798);
nand UO_1587 (O_1587,N_29962,N_29705);
or UO_1588 (O_1588,N_29813,N_29911);
or UO_1589 (O_1589,N_29992,N_29935);
and UO_1590 (O_1590,N_29845,N_29890);
xnor UO_1591 (O_1591,N_29834,N_29794);
and UO_1592 (O_1592,N_29739,N_29746);
or UO_1593 (O_1593,N_29731,N_29810);
nand UO_1594 (O_1594,N_29801,N_29752);
nor UO_1595 (O_1595,N_29829,N_29773);
nand UO_1596 (O_1596,N_29867,N_29846);
nand UO_1597 (O_1597,N_29855,N_29945);
or UO_1598 (O_1598,N_29834,N_29837);
nand UO_1599 (O_1599,N_29987,N_29931);
and UO_1600 (O_1600,N_29938,N_29818);
xor UO_1601 (O_1601,N_29778,N_29808);
nand UO_1602 (O_1602,N_29968,N_29858);
nor UO_1603 (O_1603,N_29727,N_29999);
nor UO_1604 (O_1604,N_29757,N_29959);
and UO_1605 (O_1605,N_29833,N_29821);
nor UO_1606 (O_1606,N_29746,N_29872);
nand UO_1607 (O_1607,N_29797,N_29747);
xor UO_1608 (O_1608,N_29814,N_29924);
xor UO_1609 (O_1609,N_29959,N_29915);
or UO_1610 (O_1610,N_29719,N_29709);
nor UO_1611 (O_1611,N_29770,N_29865);
nor UO_1612 (O_1612,N_29952,N_29953);
xnor UO_1613 (O_1613,N_29834,N_29718);
nor UO_1614 (O_1614,N_29847,N_29851);
nand UO_1615 (O_1615,N_29803,N_29741);
nor UO_1616 (O_1616,N_29931,N_29790);
and UO_1617 (O_1617,N_29735,N_29948);
and UO_1618 (O_1618,N_29876,N_29920);
and UO_1619 (O_1619,N_29900,N_29862);
nor UO_1620 (O_1620,N_29949,N_29859);
nor UO_1621 (O_1621,N_29815,N_29998);
and UO_1622 (O_1622,N_29745,N_29989);
and UO_1623 (O_1623,N_29843,N_29785);
or UO_1624 (O_1624,N_29861,N_29859);
and UO_1625 (O_1625,N_29940,N_29907);
or UO_1626 (O_1626,N_29755,N_29788);
and UO_1627 (O_1627,N_29754,N_29730);
nand UO_1628 (O_1628,N_29741,N_29761);
nor UO_1629 (O_1629,N_29762,N_29779);
or UO_1630 (O_1630,N_29753,N_29759);
xor UO_1631 (O_1631,N_29961,N_29994);
or UO_1632 (O_1632,N_29860,N_29812);
nand UO_1633 (O_1633,N_29756,N_29718);
xnor UO_1634 (O_1634,N_29863,N_29738);
nand UO_1635 (O_1635,N_29861,N_29965);
nand UO_1636 (O_1636,N_29725,N_29747);
or UO_1637 (O_1637,N_29709,N_29867);
xnor UO_1638 (O_1638,N_29851,N_29974);
xor UO_1639 (O_1639,N_29929,N_29785);
or UO_1640 (O_1640,N_29838,N_29787);
and UO_1641 (O_1641,N_29892,N_29701);
xor UO_1642 (O_1642,N_29731,N_29784);
xor UO_1643 (O_1643,N_29856,N_29992);
xnor UO_1644 (O_1644,N_29706,N_29973);
nor UO_1645 (O_1645,N_29988,N_29947);
nand UO_1646 (O_1646,N_29855,N_29722);
xnor UO_1647 (O_1647,N_29824,N_29728);
or UO_1648 (O_1648,N_29855,N_29990);
nand UO_1649 (O_1649,N_29782,N_29900);
nand UO_1650 (O_1650,N_29752,N_29983);
or UO_1651 (O_1651,N_29840,N_29865);
nor UO_1652 (O_1652,N_29977,N_29912);
or UO_1653 (O_1653,N_29812,N_29967);
xnor UO_1654 (O_1654,N_29793,N_29730);
nand UO_1655 (O_1655,N_29920,N_29866);
xor UO_1656 (O_1656,N_29966,N_29700);
xor UO_1657 (O_1657,N_29851,N_29859);
nand UO_1658 (O_1658,N_29728,N_29942);
nand UO_1659 (O_1659,N_29795,N_29940);
nor UO_1660 (O_1660,N_29890,N_29834);
nor UO_1661 (O_1661,N_29707,N_29975);
and UO_1662 (O_1662,N_29926,N_29851);
xor UO_1663 (O_1663,N_29974,N_29822);
nand UO_1664 (O_1664,N_29913,N_29882);
and UO_1665 (O_1665,N_29975,N_29857);
nor UO_1666 (O_1666,N_29716,N_29790);
nand UO_1667 (O_1667,N_29853,N_29711);
xor UO_1668 (O_1668,N_29852,N_29995);
xor UO_1669 (O_1669,N_29901,N_29768);
nor UO_1670 (O_1670,N_29970,N_29748);
nor UO_1671 (O_1671,N_29783,N_29739);
and UO_1672 (O_1672,N_29871,N_29907);
nand UO_1673 (O_1673,N_29747,N_29842);
nand UO_1674 (O_1674,N_29858,N_29965);
or UO_1675 (O_1675,N_29983,N_29916);
xor UO_1676 (O_1676,N_29821,N_29806);
xnor UO_1677 (O_1677,N_29706,N_29755);
nand UO_1678 (O_1678,N_29828,N_29757);
nand UO_1679 (O_1679,N_29976,N_29974);
xnor UO_1680 (O_1680,N_29868,N_29725);
xor UO_1681 (O_1681,N_29916,N_29940);
nand UO_1682 (O_1682,N_29790,N_29956);
xnor UO_1683 (O_1683,N_29838,N_29981);
nor UO_1684 (O_1684,N_29807,N_29870);
and UO_1685 (O_1685,N_29713,N_29739);
and UO_1686 (O_1686,N_29831,N_29816);
xor UO_1687 (O_1687,N_29837,N_29989);
or UO_1688 (O_1688,N_29933,N_29750);
and UO_1689 (O_1689,N_29737,N_29842);
xnor UO_1690 (O_1690,N_29916,N_29944);
or UO_1691 (O_1691,N_29839,N_29869);
xnor UO_1692 (O_1692,N_29701,N_29891);
xnor UO_1693 (O_1693,N_29905,N_29738);
nor UO_1694 (O_1694,N_29889,N_29991);
xnor UO_1695 (O_1695,N_29925,N_29767);
or UO_1696 (O_1696,N_29725,N_29801);
xnor UO_1697 (O_1697,N_29876,N_29930);
xor UO_1698 (O_1698,N_29733,N_29895);
nor UO_1699 (O_1699,N_29738,N_29782);
xnor UO_1700 (O_1700,N_29927,N_29921);
or UO_1701 (O_1701,N_29717,N_29713);
nor UO_1702 (O_1702,N_29956,N_29829);
nand UO_1703 (O_1703,N_29911,N_29992);
and UO_1704 (O_1704,N_29708,N_29957);
xor UO_1705 (O_1705,N_29865,N_29727);
nand UO_1706 (O_1706,N_29898,N_29904);
nand UO_1707 (O_1707,N_29879,N_29923);
nand UO_1708 (O_1708,N_29753,N_29777);
and UO_1709 (O_1709,N_29836,N_29990);
and UO_1710 (O_1710,N_29787,N_29811);
xnor UO_1711 (O_1711,N_29737,N_29835);
and UO_1712 (O_1712,N_29949,N_29921);
and UO_1713 (O_1713,N_29724,N_29898);
nor UO_1714 (O_1714,N_29812,N_29804);
xnor UO_1715 (O_1715,N_29959,N_29798);
and UO_1716 (O_1716,N_29762,N_29705);
xnor UO_1717 (O_1717,N_29787,N_29782);
and UO_1718 (O_1718,N_29770,N_29740);
nor UO_1719 (O_1719,N_29944,N_29991);
or UO_1720 (O_1720,N_29753,N_29903);
nand UO_1721 (O_1721,N_29938,N_29749);
or UO_1722 (O_1722,N_29973,N_29876);
xnor UO_1723 (O_1723,N_29972,N_29726);
xnor UO_1724 (O_1724,N_29924,N_29906);
nor UO_1725 (O_1725,N_29844,N_29700);
xnor UO_1726 (O_1726,N_29821,N_29997);
or UO_1727 (O_1727,N_29709,N_29848);
nor UO_1728 (O_1728,N_29981,N_29766);
nand UO_1729 (O_1729,N_29864,N_29804);
xnor UO_1730 (O_1730,N_29715,N_29823);
nand UO_1731 (O_1731,N_29974,N_29852);
nor UO_1732 (O_1732,N_29792,N_29778);
or UO_1733 (O_1733,N_29756,N_29982);
or UO_1734 (O_1734,N_29710,N_29867);
nand UO_1735 (O_1735,N_29905,N_29900);
or UO_1736 (O_1736,N_29848,N_29788);
nor UO_1737 (O_1737,N_29778,N_29813);
or UO_1738 (O_1738,N_29976,N_29919);
or UO_1739 (O_1739,N_29711,N_29787);
or UO_1740 (O_1740,N_29741,N_29708);
or UO_1741 (O_1741,N_29882,N_29916);
xnor UO_1742 (O_1742,N_29731,N_29952);
nor UO_1743 (O_1743,N_29782,N_29912);
nor UO_1744 (O_1744,N_29713,N_29865);
nand UO_1745 (O_1745,N_29831,N_29735);
nor UO_1746 (O_1746,N_29837,N_29858);
nor UO_1747 (O_1747,N_29982,N_29774);
and UO_1748 (O_1748,N_29760,N_29744);
and UO_1749 (O_1749,N_29792,N_29727);
or UO_1750 (O_1750,N_29994,N_29858);
xnor UO_1751 (O_1751,N_29966,N_29918);
nand UO_1752 (O_1752,N_29773,N_29840);
or UO_1753 (O_1753,N_29896,N_29832);
nand UO_1754 (O_1754,N_29803,N_29743);
xor UO_1755 (O_1755,N_29927,N_29794);
or UO_1756 (O_1756,N_29745,N_29771);
or UO_1757 (O_1757,N_29912,N_29802);
nor UO_1758 (O_1758,N_29901,N_29860);
nor UO_1759 (O_1759,N_29930,N_29961);
nand UO_1760 (O_1760,N_29860,N_29738);
xor UO_1761 (O_1761,N_29977,N_29701);
and UO_1762 (O_1762,N_29966,N_29979);
and UO_1763 (O_1763,N_29911,N_29980);
xnor UO_1764 (O_1764,N_29786,N_29804);
or UO_1765 (O_1765,N_29889,N_29789);
xor UO_1766 (O_1766,N_29804,N_29963);
xor UO_1767 (O_1767,N_29700,N_29879);
nand UO_1768 (O_1768,N_29787,N_29707);
xor UO_1769 (O_1769,N_29873,N_29860);
xnor UO_1770 (O_1770,N_29719,N_29844);
and UO_1771 (O_1771,N_29778,N_29920);
xor UO_1772 (O_1772,N_29855,N_29786);
or UO_1773 (O_1773,N_29707,N_29784);
xor UO_1774 (O_1774,N_29932,N_29744);
nand UO_1775 (O_1775,N_29827,N_29946);
or UO_1776 (O_1776,N_29734,N_29826);
and UO_1777 (O_1777,N_29800,N_29911);
and UO_1778 (O_1778,N_29744,N_29751);
nand UO_1779 (O_1779,N_29798,N_29759);
and UO_1780 (O_1780,N_29868,N_29906);
or UO_1781 (O_1781,N_29836,N_29903);
or UO_1782 (O_1782,N_29911,N_29823);
and UO_1783 (O_1783,N_29824,N_29742);
xnor UO_1784 (O_1784,N_29974,N_29928);
nand UO_1785 (O_1785,N_29797,N_29709);
nor UO_1786 (O_1786,N_29751,N_29776);
nor UO_1787 (O_1787,N_29786,N_29857);
and UO_1788 (O_1788,N_29717,N_29902);
or UO_1789 (O_1789,N_29937,N_29759);
or UO_1790 (O_1790,N_29857,N_29863);
and UO_1791 (O_1791,N_29889,N_29990);
nand UO_1792 (O_1792,N_29903,N_29945);
or UO_1793 (O_1793,N_29849,N_29717);
nand UO_1794 (O_1794,N_29797,N_29925);
and UO_1795 (O_1795,N_29965,N_29786);
xor UO_1796 (O_1796,N_29852,N_29732);
nor UO_1797 (O_1797,N_29970,N_29961);
or UO_1798 (O_1798,N_29792,N_29990);
nor UO_1799 (O_1799,N_29779,N_29900);
and UO_1800 (O_1800,N_29923,N_29777);
and UO_1801 (O_1801,N_29736,N_29987);
nand UO_1802 (O_1802,N_29910,N_29908);
nand UO_1803 (O_1803,N_29934,N_29858);
or UO_1804 (O_1804,N_29891,N_29961);
xor UO_1805 (O_1805,N_29775,N_29802);
xnor UO_1806 (O_1806,N_29908,N_29995);
nor UO_1807 (O_1807,N_29750,N_29980);
xor UO_1808 (O_1808,N_29751,N_29975);
nor UO_1809 (O_1809,N_29774,N_29743);
nand UO_1810 (O_1810,N_29882,N_29984);
nand UO_1811 (O_1811,N_29907,N_29841);
or UO_1812 (O_1812,N_29758,N_29714);
nand UO_1813 (O_1813,N_29902,N_29844);
nand UO_1814 (O_1814,N_29787,N_29773);
nand UO_1815 (O_1815,N_29792,N_29799);
or UO_1816 (O_1816,N_29827,N_29951);
and UO_1817 (O_1817,N_29836,N_29817);
xnor UO_1818 (O_1818,N_29933,N_29992);
nor UO_1819 (O_1819,N_29889,N_29803);
or UO_1820 (O_1820,N_29900,N_29858);
or UO_1821 (O_1821,N_29772,N_29912);
nand UO_1822 (O_1822,N_29814,N_29845);
or UO_1823 (O_1823,N_29829,N_29724);
or UO_1824 (O_1824,N_29712,N_29993);
nor UO_1825 (O_1825,N_29712,N_29916);
and UO_1826 (O_1826,N_29889,N_29775);
and UO_1827 (O_1827,N_29728,N_29761);
nand UO_1828 (O_1828,N_29942,N_29958);
xnor UO_1829 (O_1829,N_29808,N_29787);
nor UO_1830 (O_1830,N_29804,N_29892);
or UO_1831 (O_1831,N_29718,N_29957);
xor UO_1832 (O_1832,N_29941,N_29706);
xor UO_1833 (O_1833,N_29866,N_29863);
xnor UO_1834 (O_1834,N_29757,N_29712);
xor UO_1835 (O_1835,N_29857,N_29954);
and UO_1836 (O_1836,N_29790,N_29813);
xnor UO_1837 (O_1837,N_29748,N_29948);
xnor UO_1838 (O_1838,N_29748,N_29997);
xor UO_1839 (O_1839,N_29809,N_29837);
xnor UO_1840 (O_1840,N_29768,N_29995);
or UO_1841 (O_1841,N_29791,N_29787);
xnor UO_1842 (O_1842,N_29809,N_29812);
or UO_1843 (O_1843,N_29952,N_29832);
nor UO_1844 (O_1844,N_29858,N_29820);
xor UO_1845 (O_1845,N_29951,N_29944);
nor UO_1846 (O_1846,N_29984,N_29712);
nor UO_1847 (O_1847,N_29772,N_29759);
nor UO_1848 (O_1848,N_29855,N_29716);
or UO_1849 (O_1849,N_29863,N_29952);
or UO_1850 (O_1850,N_29936,N_29845);
nand UO_1851 (O_1851,N_29989,N_29999);
nor UO_1852 (O_1852,N_29962,N_29993);
and UO_1853 (O_1853,N_29933,N_29895);
xor UO_1854 (O_1854,N_29999,N_29810);
nor UO_1855 (O_1855,N_29929,N_29730);
and UO_1856 (O_1856,N_29988,N_29773);
and UO_1857 (O_1857,N_29771,N_29788);
and UO_1858 (O_1858,N_29829,N_29797);
nand UO_1859 (O_1859,N_29916,N_29757);
or UO_1860 (O_1860,N_29834,N_29865);
nand UO_1861 (O_1861,N_29939,N_29810);
xor UO_1862 (O_1862,N_29716,N_29786);
nor UO_1863 (O_1863,N_29965,N_29707);
nand UO_1864 (O_1864,N_29948,N_29707);
or UO_1865 (O_1865,N_29815,N_29922);
nor UO_1866 (O_1866,N_29725,N_29768);
and UO_1867 (O_1867,N_29879,N_29906);
nor UO_1868 (O_1868,N_29700,N_29775);
nand UO_1869 (O_1869,N_29819,N_29914);
or UO_1870 (O_1870,N_29850,N_29948);
nor UO_1871 (O_1871,N_29806,N_29792);
xor UO_1872 (O_1872,N_29985,N_29855);
nand UO_1873 (O_1873,N_29754,N_29830);
and UO_1874 (O_1874,N_29930,N_29866);
and UO_1875 (O_1875,N_29877,N_29932);
nand UO_1876 (O_1876,N_29992,N_29837);
xor UO_1877 (O_1877,N_29890,N_29872);
xor UO_1878 (O_1878,N_29911,N_29959);
nor UO_1879 (O_1879,N_29779,N_29983);
nand UO_1880 (O_1880,N_29968,N_29741);
or UO_1881 (O_1881,N_29714,N_29979);
nor UO_1882 (O_1882,N_29810,N_29927);
xnor UO_1883 (O_1883,N_29856,N_29802);
nand UO_1884 (O_1884,N_29880,N_29924);
and UO_1885 (O_1885,N_29980,N_29829);
or UO_1886 (O_1886,N_29951,N_29905);
xor UO_1887 (O_1887,N_29703,N_29926);
or UO_1888 (O_1888,N_29882,N_29745);
xnor UO_1889 (O_1889,N_29983,N_29897);
xor UO_1890 (O_1890,N_29879,N_29839);
and UO_1891 (O_1891,N_29900,N_29985);
nor UO_1892 (O_1892,N_29885,N_29938);
xnor UO_1893 (O_1893,N_29937,N_29785);
xnor UO_1894 (O_1894,N_29759,N_29824);
or UO_1895 (O_1895,N_29887,N_29837);
nand UO_1896 (O_1896,N_29700,N_29783);
nor UO_1897 (O_1897,N_29798,N_29733);
nor UO_1898 (O_1898,N_29889,N_29766);
nor UO_1899 (O_1899,N_29986,N_29832);
nand UO_1900 (O_1900,N_29908,N_29895);
and UO_1901 (O_1901,N_29802,N_29922);
nand UO_1902 (O_1902,N_29747,N_29739);
and UO_1903 (O_1903,N_29971,N_29835);
nand UO_1904 (O_1904,N_29715,N_29829);
and UO_1905 (O_1905,N_29764,N_29849);
xnor UO_1906 (O_1906,N_29996,N_29906);
or UO_1907 (O_1907,N_29968,N_29707);
nand UO_1908 (O_1908,N_29933,N_29772);
or UO_1909 (O_1909,N_29875,N_29851);
nand UO_1910 (O_1910,N_29876,N_29938);
nand UO_1911 (O_1911,N_29946,N_29898);
xor UO_1912 (O_1912,N_29790,N_29730);
nand UO_1913 (O_1913,N_29860,N_29724);
xor UO_1914 (O_1914,N_29745,N_29755);
and UO_1915 (O_1915,N_29790,N_29738);
and UO_1916 (O_1916,N_29920,N_29872);
nor UO_1917 (O_1917,N_29750,N_29934);
nor UO_1918 (O_1918,N_29704,N_29768);
nor UO_1919 (O_1919,N_29843,N_29962);
nand UO_1920 (O_1920,N_29886,N_29991);
or UO_1921 (O_1921,N_29768,N_29923);
nand UO_1922 (O_1922,N_29833,N_29908);
or UO_1923 (O_1923,N_29860,N_29752);
xor UO_1924 (O_1924,N_29883,N_29713);
or UO_1925 (O_1925,N_29963,N_29970);
xor UO_1926 (O_1926,N_29819,N_29917);
xor UO_1927 (O_1927,N_29922,N_29795);
nor UO_1928 (O_1928,N_29781,N_29897);
nor UO_1929 (O_1929,N_29880,N_29767);
xnor UO_1930 (O_1930,N_29803,N_29753);
or UO_1931 (O_1931,N_29708,N_29884);
nor UO_1932 (O_1932,N_29756,N_29935);
or UO_1933 (O_1933,N_29916,N_29877);
xnor UO_1934 (O_1934,N_29838,N_29882);
and UO_1935 (O_1935,N_29849,N_29958);
xnor UO_1936 (O_1936,N_29768,N_29798);
xnor UO_1937 (O_1937,N_29704,N_29864);
or UO_1938 (O_1938,N_29716,N_29722);
nand UO_1939 (O_1939,N_29799,N_29983);
nor UO_1940 (O_1940,N_29901,N_29945);
xnor UO_1941 (O_1941,N_29894,N_29752);
nor UO_1942 (O_1942,N_29955,N_29936);
or UO_1943 (O_1943,N_29875,N_29746);
nand UO_1944 (O_1944,N_29968,N_29980);
or UO_1945 (O_1945,N_29783,N_29846);
nand UO_1946 (O_1946,N_29799,N_29794);
xnor UO_1947 (O_1947,N_29803,N_29815);
nand UO_1948 (O_1948,N_29823,N_29861);
nor UO_1949 (O_1949,N_29967,N_29855);
nand UO_1950 (O_1950,N_29812,N_29995);
or UO_1951 (O_1951,N_29789,N_29999);
and UO_1952 (O_1952,N_29855,N_29885);
or UO_1953 (O_1953,N_29978,N_29749);
and UO_1954 (O_1954,N_29881,N_29938);
nand UO_1955 (O_1955,N_29751,N_29801);
or UO_1956 (O_1956,N_29820,N_29879);
or UO_1957 (O_1957,N_29801,N_29964);
or UO_1958 (O_1958,N_29854,N_29748);
xor UO_1959 (O_1959,N_29813,N_29762);
and UO_1960 (O_1960,N_29861,N_29754);
and UO_1961 (O_1961,N_29904,N_29907);
and UO_1962 (O_1962,N_29766,N_29748);
nand UO_1963 (O_1963,N_29955,N_29760);
nor UO_1964 (O_1964,N_29740,N_29958);
xor UO_1965 (O_1965,N_29919,N_29772);
nand UO_1966 (O_1966,N_29840,N_29780);
xnor UO_1967 (O_1967,N_29750,N_29884);
and UO_1968 (O_1968,N_29766,N_29926);
nand UO_1969 (O_1969,N_29929,N_29878);
and UO_1970 (O_1970,N_29958,N_29808);
nor UO_1971 (O_1971,N_29715,N_29782);
nand UO_1972 (O_1972,N_29834,N_29772);
xnor UO_1973 (O_1973,N_29736,N_29835);
xor UO_1974 (O_1974,N_29714,N_29820);
or UO_1975 (O_1975,N_29822,N_29849);
nand UO_1976 (O_1976,N_29952,N_29938);
nor UO_1977 (O_1977,N_29887,N_29802);
and UO_1978 (O_1978,N_29798,N_29930);
nand UO_1979 (O_1979,N_29774,N_29748);
and UO_1980 (O_1980,N_29879,N_29993);
nor UO_1981 (O_1981,N_29857,N_29828);
xor UO_1982 (O_1982,N_29952,N_29770);
nand UO_1983 (O_1983,N_29765,N_29733);
and UO_1984 (O_1984,N_29716,N_29861);
and UO_1985 (O_1985,N_29833,N_29804);
nor UO_1986 (O_1986,N_29755,N_29968);
nor UO_1987 (O_1987,N_29960,N_29959);
xnor UO_1988 (O_1988,N_29726,N_29931);
or UO_1989 (O_1989,N_29907,N_29996);
nor UO_1990 (O_1990,N_29896,N_29846);
or UO_1991 (O_1991,N_29798,N_29904);
xor UO_1992 (O_1992,N_29906,N_29832);
nand UO_1993 (O_1993,N_29848,N_29978);
xor UO_1994 (O_1994,N_29923,N_29762);
and UO_1995 (O_1995,N_29910,N_29961);
xnor UO_1996 (O_1996,N_29706,N_29716);
nand UO_1997 (O_1997,N_29905,N_29941);
or UO_1998 (O_1998,N_29890,N_29821);
nand UO_1999 (O_1999,N_29716,N_29906);
or UO_2000 (O_2000,N_29907,N_29809);
and UO_2001 (O_2001,N_29745,N_29797);
nand UO_2002 (O_2002,N_29742,N_29750);
nand UO_2003 (O_2003,N_29823,N_29817);
nor UO_2004 (O_2004,N_29763,N_29822);
nor UO_2005 (O_2005,N_29820,N_29875);
and UO_2006 (O_2006,N_29717,N_29863);
xnor UO_2007 (O_2007,N_29730,N_29762);
xnor UO_2008 (O_2008,N_29978,N_29966);
and UO_2009 (O_2009,N_29776,N_29726);
nand UO_2010 (O_2010,N_29949,N_29973);
xnor UO_2011 (O_2011,N_29847,N_29922);
nand UO_2012 (O_2012,N_29844,N_29951);
xnor UO_2013 (O_2013,N_29878,N_29974);
and UO_2014 (O_2014,N_29750,N_29921);
and UO_2015 (O_2015,N_29715,N_29991);
xor UO_2016 (O_2016,N_29967,N_29781);
nor UO_2017 (O_2017,N_29795,N_29702);
nor UO_2018 (O_2018,N_29730,N_29984);
and UO_2019 (O_2019,N_29714,N_29985);
xor UO_2020 (O_2020,N_29780,N_29834);
nor UO_2021 (O_2021,N_29707,N_29976);
and UO_2022 (O_2022,N_29813,N_29761);
nand UO_2023 (O_2023,N_29860,N_29839);
xor UO_2024 (O_2024,N_29984,N_29724);
xnor UO_2025 (O_2025,N_29889,N_29850);
and UO_2026 (O_2026,N_29876,N_29847);
xnor UO_2027 (O_2027,N_29978,N_29939);
and UO_2028 (O_2028,N_29805,N_29894);
and UO_2029 (O_2029,N_29915,N_29957);
and UO_2030 (O_2030,N_29962,N_29846);
and UO_2031 (O_2031,N_29999,N_29971);
xnor UO_2032 (O_2032,N_29710,N_29721);
xnor UO_2033 (O_2033,N_29886,N_29889);
nand UO_2034 (O_2034,N_29987,N_29705);
xor UO_2035 (O_2035,N_29950,N_29759);
and UO_2036 (O_2036,N_29994,N_29878);
xnor UO_2037 (O_2037,N_29901,N_29797);
nor UO_2038 (O_2038,N_29961,N_29933);
nand UO_2039 (O_2039,N_29722,N_29830);
and UO_2040 (O_2040,N_29819,N_29913);
or UO_2041 (O_2041,N_29958,N_29748);
nor UO_2042 (O_2042,N_29757,N_29950);
and UO_2043 (O_2043,N_29880,N_29768);
or UO_2044 (O_2044,N_29967,N_29933);
xnor UO_2045 (O_2045,N_29895,N_29808);
or UO_2046 (O_2046,N_29983,N_29992);
or UO_2047 (O_2047,N_29985,N_29760);
or UO_2048 (O_2048,N_29785,N_29727);
xor UO_2049 (O_2049,N_29799,N_29768);
nand UO_2050 (O_2050,N_29711,N_29872);
nand UO_2051 (O_2051,N_29717,N_29911);
xor UO_2052 (O_2052,N_29973,N_29726);
nor UO_2053 (O_2053,N_29770,N_29902);
or UO_2054 (O_2054,N_29748,N_29730);
xor UO_2055 (O_2055,N_29919,N_29819);
and UO_2056 (O_2056,N_29896,N_29771);
nor UO_2057 (O_2057,N_29795,N_29959);
nand UO_2058 (O_2058,N_29900,N_29788);
xor UO_2059 (O_2059,N_29738,N_29746);
nand UO_2060 (O_2060,N_29808,N_29943);
nor UO_2061 (O_2061,N_29735,N_29950);
or UO_2062 (O_2062,N_29797,N_29997);
nand UO_2063 (O_2063,N_29972,N_29960);
nor UO_2064 (O_2064,N_29960,N_29711);
and UO_2065 (O_2065,N_29995,N_29700);
nor UO_2066 (O_2066,N_29806,N_29798);
nand UO_2067 (O_2067,N_29931,N_29809);
and UO_2068 (O_2068,N_29795,N_29943);
xnor UO_2069 (O_2069,N_29718,N_29770);
or UO_2070 (O_2070,N_29705,N_29936);
and UO_2071 (O_2071,N_29811,N_29996);
nor UO_2072 (O_2072,N_29776,N_29865);
xnor UO_2073 (O_2073,N_29906,N_29711);
nand UO_2074 (O_2074,N_29725,N_29873);
nand UO_2075 (O_2075,N_29871,N_29872);
and UO_2076 (O_2076,N_29850,N_29954);
or UO_2077 (O_2077,N_29725,N_29773);
and UO_2078 (O_2078,N_29828,N_29854);
xnor UO_2079 (O_2079,N_29994,N_29764);
and UO_2080 (O_2080,N_29921,N_29998);
or UO_2081 (O_2081,N_29994,N_29914);
nor UO_2082 (O_2082,N_29715,N_29762);
nor UO_2083 (O_2083,N_29746,N_29945);
or UO_2084 (O_2084,N_29958,N_29700);
or UO_2085 (O_2085,N_29905,N_29894);
or UO_2086 (O_2086,N_29867,N_29702);
nor UO_2087 (O_2087,N_29750,N_29861);
nand UO_2088 (O_2088,N_29952,N_29985);
or UO_2089 (O_2089,N_29883,N_29875);
xnor UO_2090 (O_2090,N_29839,N_29741);
xnor UO_2091 (O_2091,N_29773,N_29940);
and UO_2092 (O_2092,N_29903,N_29936);
nand UO_2093 (O_2093,N_29823,N_29758);
nand UO_2094 (O_2094,N_29941,N_29884);
nor UO_2095 (O_2095,N_29854,N_29993);
nor UO_2096 (O_2096,N_29855,N_29904);
or UO_2097 (O_2097,N_29752,N_29850);
nand UO_2098 (O_2098,N_29990,N_29979);
xor UO_2099 (O_2099,N_29745,N_29777);
nor UO_2100 (O_2100,N_29834,N_29908);
xnor UO_2101 (O_2101,N_29801,N_29927);
and UO_2102 (O_2102,N_29706,N_29900);
xor UO_2103 (O_2103,N_29732,N_29855);
nor UO_2104 (O_2104,N_29749,N_29790);
nand UO_2105 (O_2105,N_29975,N_29833);
nand UO_2106 (O_2106,N_29939,N_29768);
xor UO_2107 (O_2107,N_29964,N_29841);
nor UO_2108 (O_2108,N_29908,N_29864);
nand UO_2109 (O_2109,N_29733,N_29760);
and UO_2110 (O_2110,N_29714,N_29989);
nor UO_2111 (O_2111,N_29977,N_29709);
xor UO_2112 (O_2112,N_29901,N_29988);
or UO_2113 (O_2113,N_29884,N_29804);
nand UO_2114 (O_2114,N_29798,N_29703);
and UO_2115 (O_2115,N_29804,N_29908);
nand UO_2116 (O_2116,N_29825,N_29873);
or UO_2117 (O_2117,N_29817,N_29849);
nor UO_2118 (O_2118,N_29733,N_29925);
nor UO_2119 (O_2119,N_29877,N_29964);
nor UO_2120 (O_2120,N_29990,N_29839);
nand UO_2121 (O_2121,N_29958,N_29845);
nor UO_2122 (O_2122,N_29719,N_29723);
or UO_2123 (O_2123,N_29933,N_29841);
nand UO_2124 (O_2124,N_29965,N_29751);
or UO_2125 (O_2125,N_29734,N_29702);
and UO_2126 (O_2126,N_29869,N_29801);
nor UO_2127 (O_2127,N_29710,N_29968);
or UO_2128 (O_2128,N_29917,N_29741);
or UO_2129 (O_2129,N_29729,N_29801);
and UO_2130 (O_2130,N_29795,N_29942);
nand UO_2131 (O_2131,N_29959,N_29823);
nand UO_2132 (O_2132,N_29721,N_29827);
nor UO_2133 (O_2133,N_29747,N_29745);
or UO_2134 (O_2134,N_29803,N_29987);
nand UO_2135 (O_2135,N_29719,N_29840);
nand UO_2136 (O_2136,N_29879,N_29924);
xnor UO_2137 (O_2137,N_29811,N_29839);
nor UO_2138 (O_2138,N_29744,N_29701);
nor UO_2139 (O_2139,N_29775,N_29805);
or UO_2140 (O_2140,N_29964,N_29741);
nand UO_2141 (O_2141,N_29896,N_29888);
and UO_2142 (O_2142,N_29766,N_29726);
or UO_2143 (O_2143,N_29710,N_29834);
xor UO_2144 (O_2144,N_29727,N_29977);
or UO_2145 (O_2145,N_29834,N_29883);
nor UO_2146 (O_2146,N_29986,N_29826);
nor UO_2147 (O_2147,N_29711,N_29834);
xor UO_2148 (O_2148,N_29919,N_29816);
xnor UO_2149 (O_2149,N_29822,N_29801);
nor UO_2150 (O_2150,N_29820,N_29870);
nor UO_2151 (O_2151,N_29972,N_29764);
or UO_2152 (O_2152,N_29832,N_29740);
and UO_2153 (O_2153,N_29746,N_29728);
nand UO_2154 (O_2154,N_29990,N_29947);
and UO_2155 (O_2155,N_29901,N_29774);
or UO_2156 (O_2156,N_29974,N_29820);
xor UO_2157 (O_2157,N_29775,N_29767);
and UO_2158 (O_2158,N_29827,N_29909);
or UO_2159 (O_2159,N_29741,N_29789);
nand UO_2160 (O_2160,N_29974,N_29921);
nand UO_2161 (O_2161,N_29790,N_29936);
or UO_2162 (O_2162,N_29829,N_29843);
nand UO_2163 (O_2163,N_29828,N_29747);
and UO_2164 (O_2164,N_29770,N_29818);
or UO_2165 (O_2165,N_29859,N_29857);
and UO_2166 (O_2166,N_29850,N_29748);
nand UO_2167 (O_2167,N_29823,N_29886);
nor UO_2168 (O_2168,N_29945,N_29716);
and UO_2169 (O_2169,N_29902,N_29957);
xnor UO_2170 (O_2170,N_29796,N_29742);
and UO_2171 (O_2171,N_29893,N_29794);
nor UO_2172 (O_2172,N_29754,N_29840);
nand UO_2173 (O_2173,N_29822,N_29918);
or UO_2174 (O_2174,N_29830,N_29800);
and UO_2175 (O_2175,N_29943,N_29999);
xor UO_2176 (O_2176,N_29940,N_29958);
or UO_2177 (O_2177,N_29915,N_29968);
nor UO_2178 (O_2178,N_29783,N_29948);
xnor UO_2179 (O_2179,N_29955,N_29948);
nor UO_2180 (O_2180,N_29863,N_29720);
or UO_2181 (O_2181,N_29811,N_29993);
nor UO_2182 (O_2182,N_29963,N_29709);
nor UO_2183 (O_2183,N_29759,N_29961);
and UO_2184 (O_2184,N_29938,N_29785);
nand UO_2185 (O_2185,N_29838,N_29703);
xor UO_2186 (O_2186,N_29832,N_29836);
xnor UO_2187 (O_2187,N_29881,N_29799);
nand UO_2188 (O_2188,N_29943,N_29842);
or UO_2189 (O_2189,N_29702,N_29758);
nor UO_2190 (O_2190,N_29721,N_29749);
and UO_2191 (O_2191,N_29736,N_29791);
nor UO_2192 (O_2192,N_29746,N_29754);
nor UO_2193 (O_2193,N_29988,N_29975);
and UO_2194 (O_2194,N_29855,N_29902);
xnor UO_2195 (O_2195,N_29809,N_29843);
nor UO_2196 (O_2196,N_29793,N_29776);
nor UO_2197 (O_2197,N_29857,N_29904);
nand UO_2198 (O_2198,N_29869,N_29886);
nor UO_2199 (O_2199,N_29749,N_29973);
nand UO_2200 (O_2200,N_29888,N_29735);
nor UO_2201 (O_2201,N_29804,N_29801);
and UO_2202 (O_2202,N_29727,N_29824);
or UO_2203 (O_2203,N_29997,N_29756);
nor UO_2204 (O_2204,N_29750,N_29728);
or UO_2205 (O_2205,N_29882,N_29945);
and UO_2206 (O_2206,N_29735,N_29756);
nand UO_2207 (O_2207,N_29897,N_29805);
or UO_2208 (O_2208,N_29714,N_29783);
nand UO_2209 (O_2209,N_29715,N_29947);
or UO_2210 (O_2210,N_29894,N_29708);
or UO_2211 (O_2211,N_29712,N_29786);
or UO_2212 (O_2212,N_29878,N_29888);
nor UO_2213 (O_2213,N_29910,N_29808);
nand UO_2214 (O_2214,N_29851,N_29790);
and UO_2215 (O_2215,N_29729,N_29786);
and UO_2216 (O_2216,N_29752,N_29969);
nor UO_2217 (O_2217,N_29892,N_29996);
nand UO_2218 (O_2218,N_29785,N_29801);
nor UO_2219 (O_2219,N_29809,N_29708);
nor UO_2220 (O_2220,N_29840,N_29740);
or UO_2221 (O_2221,N_29784,N_29857);
nor UO_2222 (O_2222,N_29930,N_29954);
and UO_2223 (O_2223,N_29932,N_29833);
nor UO_2224 (O_2224,N_29810,N_29929);
or UO_2225 (O_2225,N_29919,N_29823);
xor UO_2226 (O_2226,N_29762,N_29858);
or UO_2227 (O_2227,N_29786,N_29767);
nand UO_2228 (O_2228,N_29751,N_29706);
or UO_2229 (O_2229,N_29811,N_29893);
xor UO_2230 (O_2230,N_29816,N_29737);
or UO_2231 (O_2231,N_29838,N_29719);
or UO_2232 (O_2232,N_29917,N_29914);
and UO_2233 (O_2233,N_29825,N_29851);
xnor UO_2234 (O_2234,N_29727,N_29751);
nand UO_2235 (O_2235,N_29719,N_29850);
or UO_2236 (O_2236,N_29728,N_29703);
nand UO_2237 (O_2237,N_29968,N_29929);
nor UO_2238 (O_2238,N_29829,N_29931);
nand UO_2239 (O_2239,N_29786,N_29966);
xor UO_2240 (O_2240,N_29892,N_29710);
nand UO_2241 (O_2241,N_29907,N_29898);
xor UO_2242 (O_2242,N_29709,N_29973);
or UO_2243 (O_2243,N_29906,N_29992);
and UO_2244 (O_2244,N_29904,N_29749);
nor UO_2245 (O_2245,N_29863,N_29941);
and UO_2246 (O_2246,N_29848,N_29875);
nand UO_2247 (O_2247,N_29731,N_29943);
or UO_2248 (O_2248,N_29747,N_29944);
or UO_2249 (O_2249,N_29986,N_29743);
xnor UO_2250 (O_2250,N_29977,N_29708);
nor UO_2251 (O_2251,N_29762,N_29812);
xnor UO_2252 (O_2252,N_29982,N_29776);
nor UO_2253 (O_2253,N_29957,N_29871);
nand UO_2254 (O_2254,N_29912,N_29886);
nor UO_2255 (O_2255,N_29774,N_29765);
nor UO_2256 (O_2256,N_29989,N_29943);
nor UO_2257 (O_2257,N_29938,N_29739);
or UO_2258 (O_2258,N_29859,N_29778);
nor UO_2259 (O_2259,N_29754,N_29937);
nand UO_2260 (O_2260,N_29941,N_29925);
or UO_2261 (O_2261,N_29767,N_29713);
nor UO_2262 (O_2262,N_29935,N_29891);
and UO_2263 (O_2263,N_29871,N_29974);
xnor UO_2264 (O_2264,N_29827,N_29769);
or UO_2265 (O_2265,N_29706,N_29899);
nand UO_2266 (O_2266,N_29970,N_29999);
or UO_2267 (O_2267,N_29844,N_29778);
xnor UO_2268 (O_2268,N_29876,N_29957);
xnor UO_2269 (O_2269,N_29715,N_29810);
nor UO_2270 (O_2270,N_29781,N_29978);
and UO_2271 (O_2271,N_29992,N_29708);
nor UO_2272 (O_2272,N_29836,N_29740);
and UO_2273 (O_2273,N_29737,N_29864);
nor UO_2274 (O_2274,N_29985,N_29845);
or UO_2275 (O_2275,N_29890,N_29885);
and UO_2276 (O_2276,N_29782,N_29758);
nor UO_2277 (O_2277,N_29746,N_29905);
and UO_2278 (O_2278,N_29929,N_29705);
and UO_2279 (O_2279,N_29925,N_29826);
nor UO_2280 (O_2280,N_29909,N_29791);
and UO_2281 (O_2281,N_29739,N_29909);
nand UO_2282 (O_2282,N_29806,N_29701);
and UO_2283 (O_2283,N_29877,N_29833);
nand UO_2284 (O_2284,N_29878,N_29762);
nor UO_2285 (O_2285,N_29759,N_29803);
and UO_2286 (O_2286,N_29720,N_29899);
xnor UO_2287 (O_2287,N_29860,N_29827);
xnor UO_2288 (O_2288,N_29788,N_29826);
nand UO_2289 (O_2289,N_29854,N_29773);
nor UO_2290 (O_2290,N_29831,N_29791);
nand UO_2291 (O_2291,N_29939,N_29823);
or UO_2292 (O_2292,N_29890,N_29947);
nand UO_2293 (O_2293,N_29866,N_29966);
nand UO_2294 (O_2294,N_29982,N_29987);
and UO_2295 (O_2295,N_29964,N_29885);
nor UO_2296 (O_2296,N_29796,N_29700);
xor UO_2297 (O_2297,N_29773,N_29990);
nor UO_2298 (O_2298,N_29756,N_29789);
nor UO_2299 (O_2299,N_29994,N_29978);
or UO_2300 (O_2300,N_29897,N_29750);
xor UO_2301 (O_2301,N_29869,N_29851);
nand UO_2302 (O_2302,N_29962,N_29783);
or UO_2303 (O_2303,N_29933,N_29794);
or UO_2304 (O_2304,N_29981,N_29745);
nand UO_2305 (O_2305,N_29762,N_29925);
xor UO_2306 (O_2306,N_29724,N_29810);
xnor UO_2307 (O_2307,N_29950,N_29926);
and UO_2308 (O_2308,N_29929,N_29798);
or UO_2309 (O_2309,N_29892,N_29905);
and UO_2310 (O_2310,N_29785,N_29993);
xor UO_2311 (O_2311,N_29999,N_29912);
and UO_2312 (O_2312,N_29711,N_29961);
and UO_2313 (O_2313,N_29710,N_29891);
nand UO_2314 (O_2314,N_29715,N_29854);
and UO_2315 (O_2315,N_29989,N_29944);
nand UO_2316 (O_2316,N_29997,N_29881);
and UO_2317 (O_2317,N_29770,N_29714);
nor UO_2318 (O_2318,N_29862,N_29804);
and UO_2319 (O_2319,N_29978,N_29867);
or UO_2320 (O_2320,N_29774,N_29793);
or UO_2321 (O_2321,N_29739,N_29726);
xor UO_2322 (O_2322,N_29941,N_29827);
nor UO_2323 (O_2323,N_29852,N_29898);
and UO_2324 (O_2324,N_29863,N_29744);
xor UO_2325 (O_2325,N_29807,N_29752);
or UO_2326 (O_2326,N_29928,N_29742);
and UO_2327 (O_2327,N_29702,N_29880);
nand UO_2328 (O_2328,N_29712,N_29718);
nand UO_2329 (O_2329,N_29930,N_29729);
and UO_2330 (O_2330,N_29725,N_29765);
nor UO_2331 (O_2331,N_29960,N_29968);
nand UO_2332 (O_2332,N_29826,N_29928);
nor UO_2333 (O_2333,N_29916,N_29862);
nand UO_2334 (O_2334,N_29780,N_29980);
or UO_2335 (O_2335,N_29968,N_29733);
and UO_2336 (O_2336,N_29805,N_29735);
or UO_2337 (O_2337,N_29863,N_29874);
nor UO_2338 (O_2338,N_29964,N_29811);
nand UO_2339 (O_2339,N_29752,N_29897);
nand UO_2340 (O_2340,N_29861,N_29709);
nor UO_2341 (O_2341,N_29941,N_29769);
and UO_2342 (O_2342,N_29776,N_29902);
and UO_2343 (O_2343,N_29956,N_29731);
or UO_2344 (O_2344,N_29824,N_29860);
xnor UO_2345 (O_2345,N_29729,N_29733);
or UO_2346 (O_2346,N_29968,N_29744);
xor UO_2347 (O_2347,N_29760,N_29801);
nand UO_2348 (O_2348,N_29749,N_29820);
nand UO_2349 (O_2349,N_29719,N_29853);
or UO_2350 (O_2350,N_29729,N_29899);
nor UO_2351 (O_2351,N_29917,N_29805);
nor UO_2352 (O_2352,N_29820,N_29757);
nor UO_2353 (O_2353,N_29831,N_29856);
nand UO_2354 (O_2354,N_29746,N_29881);
or UO_2355 (O_2355,N_29840,N_29995);
xor UO_2356 (O_2356,N_29835,N_29758);
xnor UO_2357 (O_2357,N_29844,N_29928);
nand UO_2358 (O_2358,N_29977,N_29851);
xor UO_2359 (O_2359,N_29995,N_29827);
nand UO_2360 (O_2360,N_29949,N_29860);
xnor UO_2361 (O_2361,N_29985,N_29955);
and UO_2362 (O_2362,N_29741,N_29913);
or UO_2363 (O_2363,N_29829,N_29755);
nor UO_2364 (O_2364,N_29956,N_29726);
or UO_2365 (O_2365,N_29818,N_29768);
or UO_2366 (O_2366,N_29858,N_29987);
or UO_2367 (O_2367,N_29972,N_29842);
or UO_2368 (O_2368,N_29860,N_29706);
nand UO_2369 (O_2369,N_29902,N_29897);
xor UO_2370 (O_2370,N_29989,N_29719);
and UO_2371 (O_2371,N_29839,N_29864);
or UO_2372 (O_2372,N_29950,N_29944);
or UO_2373 (O_2373,N_29706,N_29859);
xnor UO_2374 (O_2374,N_29777,N_29846);
nand UO_2375 (O_2375,N_29804,N_29916);
and UO_2376 (O_2376,N_29874,N_29954);
nor UO_2377 (O_2377,N_29706,N_29794);
xor UO_2378 (O_2378,N_29941,N_29789);
and UO_2379 (O_2379,N_29887,N_29787);
nand UO_2380 (O_2380,N_29775,N_29769);
xor UO_2381 (O_2381,N_29908,N_29872);
and UO_2382 (O_2382,N_29944,N_29820);
nand UO_2383 (O_2383,N_29859,N_29822);
nor UO_2384 (O_2384,N_29752,N_29775);
xor UO_2385 (O_2385,N_29773,N_29816);
or UO_2386 (O_2386,N_29742,N_29929);
or UO_2387 (O_2387,N_29780,N_29894);
or UO_2388 (O_2388,N_29945,N_29709);
nor UO_2389 (O_2389,N_29792,N_29772);
or UO_2390 (O_2390,N_29920,N_29901);
nor UO_2391 (O_2391,N_29941,N_29761);
and UO_2392 (O_2392,N_29948,N_29869);
nor UO_2393 (O_2393,N_29778,N_29891);
nor UO_2394 (O_2394,N_29945,N_29987);
and UO_2395 (O_2395,N_29898,N_29965);
and UO_2396 (O_2396,N_29835,N_29815);
and UO_2397 (O_2397,N_29700,N_29886);
nor UO_2398 (O_2398,N_29862,N_29725);
nor UO_2399 (O_2399,N_29814,N_29768);
nor UO_2400 (O_2400,N_29800,N_29810);
xnor UO_2401 (O_2401,N_29746,N_29943);
nand UO_2402 (O_2402,N_29805,N_29845);
or UO_2403 (O_2403,N_29930,N_29715);
and UO_2404 (O_2404,N_29846,N_29898);
nand UO_2405 (O_2405,N_29779,N_29867);
nand UO_2406 (O_2406,N_29821,N_29983);
and UO_2407 (O_2407,N_29978,N_29946);
nor UO_2408 (O_2408,N_29905,N_29785);
and UO_2409 (O_2409,N_29864,N_29942);
nor UO_2410 (O_2410,N_29961,N_29846);
or UO_2411 (O_2411,N_29961,N_29865);
or UO_2412 (O_2412,N_29728,N_29817);
xor UO_2413 (O_2413,N_29854,N_29875);
nor UO_2414 (O_2414,N_29950,N_29733);
xnor UO_2415 (O_2415,N_29753,N_29804);
xor UO_2416 (O_2416,N_29719,N_29977);
nand UO_2417 (O_2417,N_29702,N_29908);
xnor UO_2418 (O_2418,N_29920,N_29817);
xnor UO_2419 (O_2419,N_29837,N_29915);
xor UO_2420 (O_2420,N_29755,N_29945);
or UO_2421 (O_2421,N_29914,N_29715);
nand UO_2422 (O_2422,N_29779,N_29898);
nand UO_2423 (O_2423,N_29904,N_29803);
nand UO_2424 (O_2424,N_29914,N_29950);
and UO_2425 (O_2425,N_29707,N_29746);
and UO_2426 (O_2426,N_29792,N_29875);
nor UO_2427 (O_2427,N_29771,N_29755);
nor UO_2428 (O_2428,N_29877,N_29738);
or UO_2429 (O_2429,N_29940,N_29726);
and UO_2430 (O_2430,N_29832,N_29921);
xnor UO_2431 (O_2431,N_29919,N_29767);
xnor UO_2432 (O_2432,N_29961,N_29748);
or UO_2433 (O_2433,N_29976,N_29955);
or UO_2434 (O_2434,N_29912,N_29924);
or UO_2435 (O_2435,N_29810,N_29775);
or UO_2436 (O_2436,N_29825,N_29830);
nand UO_2437 (O_2437,N_29783,N_29960);
and UO_2438 (O_2438,N_29988,N_29747);
nand UO_2439 (O_2439,N_29770,N_29769);
xnor UO_2440 (O_2440,N_29905,N_29704);
nor UO_2441 (O_2441,N_29870,N_29869);
or UO_2442 (O_2442,N_29943,N_29825);
nand UO_2443 (O_2443,N_29952,N_29710);
nor UO_2444 (O_2444,N_29961,N_29796);
nor UO_2445 (O_2445,N_29815,N_29933);
nand UO_2446 (O_2446,N_29987,N_29900);
or UO_2447 (O_2447,N_29888,N_29779);
or UO_2448 (O_2448,N_29837,N_29719);
nor UO_2449 (O_2449,N_29820,N_29962);
and UO_2450 (O_2450,N_29770,N_29988);
xor UO_2451 (O_2451,N_29850,N_29745);
xnor UO_2452 (O_2452,N_29924,N_29896);
and UO_2453 (O_2453,N_29879,N_29936);
nand UO_2454 (O_2454,N_29857,N_29948);
or UO_2455 (O_2455,N_29813,N_29820);
nand UO_2456 (O_2456,N_29935,N_29977);
and UO_2457 (O_2457,N_29799,N_29904);
nor UO_2458 (O_2458,N_29787,N_29769);
and UO_2459 (O_2459,N_29793,N_29977);
and UO_2460 (O_2460,N_29914,N_29966);
and UO_2461 (O_2461,N_29726,N_29978);
or UO_2462 (O_2462,N_29868,N_29857);
nand UO_2463 (O_2463,N_29842,N_29899);
and UO_2464 (O_2464,N_29995,N_29753);
xnor UO_2465 (O_2465,N_29809,N_29723);
xnor UO_2466 (O_2466,N_29922,N_29700);
or UO_2467 (O_2467,N_29728,N_29843);
or UO_2468 (O_2468,N_29949,N_29980);
xor UO_2469 (O_2469,N_29782,N_29752);
or UO_2470 (O_2470,N_29989,N_29871);
and UO_2471 (O_2471,N_29967,N_29711);
nand UO_2472 (O_2472,N_29917,N_29966);
xor UO_2473 (O_2473,N_29918,N_29714);
xnor UO_2474 (O_2474,N_29944,N_29708);
or UO_2475 (O_2475,N_29747,N_29763);
or UO_2476 (O_2476,N_29924,N_29931);
and UO_2477 (O_2477,N_29954,N_29858);
or UO_2478 (O_2478,N_29983,N_29977);
nor UO_2479 (O_2479,N_29732,N_29850);
nand UO_2480 (O_2480,N_29967,N_29872);
and UO_2481 (O_2481,N_29812,N_29976);
and UO_2482 (O_2482,N_29740,N_29988);
xnor UO_2483 (O_2483,N_29716,N_29791);
and UO_2484 (O_2484,N_29967,N_29988);
nor UO_2485 (O_2485,N_29708,N_29790);
xor UO_2486 (O_2486,N_29719,N_29737);
nor UO_2487 (O_2487,N_29728,N_29853);
nor UO_2488 (O_2488,N_29960,N_29919);
nor UO_2489 (O_2489,N_29753,N_29736);
xnor UO_2490 (O_2490,N_29985,N_29737);
and UO_2491 (O_2491,N_29939,N_29702);
nand UO_2492 (O_2492,N_29788,N_29764);
xnor UO_2493 (O_2493,N_29922,N_29843);
xor UO_2494 (O_2494,N_29843,N_29803);
xnor UO_2495 (O_2495,N_29851,N_29853);
xnor UO_2496 (O_2496,N_29756,N_29737);
and UO_2497 (O_2497,N_29960,N_29719);
xnor UO_2498 (O_2498,N_29838,N_29997);
nor UO_2499 (O_2499,N_29903,N_29962);
nand UO_2500 (O_2500,N_29706,N_29741);
nand UO_2501 (O_2501,N_29703,N_29701);
nor UO_2502 (O_2502,N_29831,N_29893);
nand UO_2503 (O_2503,N_29985,N_29901);
nand UO_2504 (O_2504,N_29926,N_29798);
nor UO_2505 (O_2505,N_29976,N_29724);
nand UO_2506 (O_2506,N_29989,N_29735);
xor UO_2507 (O_2507,N_29985,N_29865);
nand UO_2508 (O_2508,N_29917,N_29980);
xor UO_2509 (O_2509,N_29827,N_29775);
and UO_2510 (O_2510,N_29941,N_29907);
or UO_2511 (O_2511,N_29710,N_29790);
nand UO_2512 (O_2512,N_29730,N_29829);
and UO_2513 (O_2513,N_29925,N_29954);
nor UO_2514 (O_2514,N_29867,N_29790);
nand UO_2515 (O_2515,N_29828,N_29867);
nand UO_2516 (O_2516,N_29825,N_29837);
nor UO_2517 (O_2517,N_29742,N_29955);
or UO_2518 (O_2518,N_29957,N_29908);
and UO_2519 (O_2519,N_29963,N_29706);
and UO_2520 (O_2520,N_29905,N_29932);
nand UO_2521 (O_2521,N_29751,N_29704);
nor UO_2522 (O_2522,N_29809,N_29761);
nand UO_2523 (O_2523,N_29969,N_29749);
nand UO_2524 (O_2524,N_29803,N_29869);
nand UO_2525 (O_2525,N_29856,N_29709);
nor UO_2526 (O_2526,N_29729,N_29759);
and UO_2527 (O_2527,N_29787,N_29839);
or UO_2528 (O_2528,N_29725,N_29962);
xnor UO_2529 (O_2529,N_29918,N_29908);
nor UO_2530 (O_2530,N_29807,N_29893);
nor UO_2531 (O_2531,N_29776,N_29924);
xor UO_2532 (O_2532,N_29858,N_29870);
xor UO_2533 (O_2533,N_29910,N_29912);
or UO_2534 (O_2534,N_29748,N_29867);
xor UO_2535 (O_2535,N_29905,N_29720);
or UO_2536 (O_2536,N_29733,N_29989);
or UO_2537 (O_2537,N_29954,N_29949);
nor UO_2538 (O_2538,N_29948,N_29958);
nand UO_2539 (O_2539,N_29883,N_29956);
nand UO_2540 (O_2540,N_29961,N_29787);
xnor UO_2541 (O_2541,N_29851,N_29777);
xnor UO_2542 (O_2542,N_29731,N_29941);
xor UO_2543 (O_2543,N_29855,N_29890);
nor UO_2544 (O_2544,N_29743,N_29775);
and UO_2545 (O_2545,N_29864,N_29885);
and UO_2546 (O_2546,N_29713,N_29800);
nor UO_2547 (O_2547,N_29859,N_29821);
nand UO_2548 (O_2548,N_29775,N_29761);
and UO_2549 (O_2549,N_29934,N_29922);
xor UO_2550 (O_2550,N_29707,N_29724);
nor UO_2551 (O_2551,N_29830,N_29813);
and UO_2552 (O_2552,N_29914,N_29883);
and UO_2553 (O_2553,N_29804,N_29737);
and UO_2554 (O_2554,N_29786,N_29747);
xor UO_2555 (O_2555,N_29893,N_29968);
nor UO_2556 (O_2556,N_29793,N_29861);
xor UO_2557 (O_2557,N_29721,N_29997);
xnor UO_2558 (O_2558,N_29896,N_29780);
or UO_2559 (O_2559,N_29975,N_29715);
or UO_2560 (O_2560,N_29790,N_29901);
nand UO_2561 (O_2561,N_29897,N_29913);
or UO_2562 (O_2562,N_29956,N_29964);
nand UO_2563 (O_2563,N_29950,N_29753);
or UO_2564 (O_2564,N_29758,N_29777);
nor UO_2565 (O_2565,N_29917,N_29969);
nor UO_2566 (O_2566,N_29885,N_29934);
or UO_2567 (O_2567,N_29990,N_29877);
xor UO_2568 (O_2568,N_29873,N_29960);
or UO_2569 (O_2569,N_29725,N_29919);
nor UO_2570 (O_2570,N_29874,N_29903);
or UO_2571 (O_2571,N_29895,N_29949);
and UO_2572 (O_2572,N_29853,N_29858);
or UO_2573 (O_2573,N_29793,N_29749);
and UO_2574 (O_2574,N_29849,N_29747);
and UO_2575 (O_2575,N_29989,N_29994);
nor UO_2576 (O_2576,N_29729,N_29724);
xnor UO_2577 (O_2577,N_29865,N_29960);
xor UO_2578 (O_2578,N_29949,N_29773);
nand UO_2579 (O_2579,N_29818,N_29785);
nor UO_2580 (O_2580,N_29955,N_29995);
or UO_2581 (O_2581,N_29958,N_29972);
or UO_2582 (O_2582,N_29703,N_29806);
nand UO_2583 (O_2583,N_29952,N_29845);
and UO_2584 (O_2584,N_29944,N_29876);
xnor UO_2585 (O_2585,N_29958,N_29757);
nand UO_2586 (O_2586,N_29912,N_29822);
or UO_2587 (O_2587,N_29759,N_29928);
nand UO_2588 (O_2588,N_29994,N_29891);
xor UO_2589 (O_2589,N_29871,N_29857);
nand UO_2590 (O_2590,N_29843,N_29784);
or UO_2591 (O_2591,N_29731,N_29792);
or UO_2592 (O_2592,N_29768,N_29841);
nor UO_2593 (O_2593,N_29870,N_29785);
or UO_2594 (O_2594,N_29710,N_29730);
and UO_2595 (O_2595,N_29842,N_29755);
or UO_2596 (O_2596,N_29929,N_29762);
or UO_2597 (O_2597,N_29797,N_29982);
and UO_2598 (O_2598,N_29748,N_29824);
and UO_2599 (O_2599,N_29884,N_29744);
nand UO_2600 (O_2600,N_29797,N_29824);
xnor UO_2601 (O_2601,N_29809,N_29913);
nor UO_2602 (O_2602,N_29824,N_29991);
nand UO_2603 (O_2603,N_29783,N_29744);
or UO_2604 (O_2604,N_29767,N_29968);
or UO_2605 (O_2605,N_29803,N_29965);
xor UO_2606 (O_2606,N_29860,N_29799);
or UO_2607 (O_2607,N_29855,N_29988);
and UO_2608 (O_2608,N_29948,N_29706);
or UO_2609 (O_2609,N_29812,N_29947);
xor UO_2610 (O_2610,N_29772,N_29793);
nor UO_2611 (O_2611,N_29796,N_29730);
nor UO_2612 (O_2612,N_29978,N_29970);
or UO_2613 (O_2613,N_29856,N_29707);
nor UO_2614 (O_2614,N_29850,N_29754);
and UO_2615 (O_2615,N_29813,N_29960);
and UO_2616 (O_2616,N_29856,N_29862);
or UO_2617 (O_2617,N_29884,N_29897);
or UO_2618 (O_2618,N_29764,N_29703);
and UO_2619 (O_2619,N_29923,N_29772);
nand UO_2620 (O_2620,N_29984,N_29852);
xor UO_2621 (O_2621,N_29930,N_29872);
nor UO_2622 (O_2622,N_29981,N_29963);
or UO_2623 (O_2623,N_29831,N_29963);
nand UO_2624 (O_2624,N_29806,N_29991);
xor UO_2625 (O_2625,N_29705,N_29995);
nor UO_2626 (O_2626,N_29935,N_29776);
xor UO_2627 (O_2627,N_29862,N_29748);
or UO_2628 (O_2628,N_29919,N_29812);
and UO_2629 (O_2629,N_29984,N_29793);
and UO_2630 (O_2630,N_29940,N_29815);
nor UO_2631 (O_2631,N_29793,N_29882);
nand UO_2632 (O_2632,N_29729,N_29768);
nand UO_2633 (O_2633,N_29892,N_29834);
nand UO_2634 (O_2634,N_29814,N_29931);
nor UO_2635 (O_2635,N_29718,N_29854);
nand UO_2636 (O_2636,N_29701,N_29812);
and UO_2637 (O_2637,N_29868,N_29796);
xnor UO_2638 (O_2638,N_29802,N_29815);
xor UO_2639 (O_2639,N_29913,N_29986);
xnor UO_2640 (O_2640,N_29836,N_29893);
nand UO_2641 (O_2641,N_29974,N_29713);
nand UO_2642 (O_2642,N_29945,N_29892);
xnor UO_2643 (O_2643,N_29740,N_29907);
nand UO_2644 (O_2644,N_29952,N_29787);
and UO_2645 (O_2645,N_29808,N_29830);
nor UO_2646 (O_2646,N_29763,N_29932);
or UO_2647 (O_2647,N_29726,N_29834);
and UO_2648 (O_2648,N_29820,N_29814);
and UO_2649 (O_2649,N_29795,N_29929);
xor UO_2650 (O_2650,N_29765,N_29861);
or UO_2651 (O_2651,N_29794,N_29961);
xor UO_2652 (O_2652,N_29995,N_29847);
or UO_2653 (O_2653,N_29980,N_29925);
and UO_2654 (O_2654,N_29815,N_29771);
nor UO_2655 (O_2655,N_29700,N_29849);
and UO_2656 (O_2656,N_29981,N_29935);
or UO_2657 (O_2657,N_29880,N_29965);
nor UO_2658 (O_2658,N_29839,N_29950);
xnor UO_2659 (O_2659,N_29727,N_29998);
nor UO_2660 (O_2660,N_29936,N_29945);
xor UO_2661 (O_2661,N_29934,N_29834);
nand UO_2662 (O_2662,N_29982,N_29786);
nor UO_2663 (O_2663,N_29722,N_29807);
or UO_2664 (O_2664,N_29911,N_29773);
xor UO_2665 (O_2665,N_29782,N_29827);
and UO_2666 (O_2666,N_29795,N_29827);
xor UO_2667 (O_2667,N_29767,N_29899);
nor UO_2668 (O_2668,N_29761,N_29866);
or UO_2669 (O_2669,N_29700,N_29928);
nor UO_2670 (O_2670,N_29976,N_29992);
xor UO_2671 (O_2671,N_29741,N_29815);
nand UO_2672 (O_2672,N_29792,N_29820);
nand UO_2673 (O_2673,N_29941,N_29900);
and UO_2674 (O_2674,N_29891,N_29980);
and UO_2675 (O_2675,N_29985,N_29805);
xnor UO_2676 (O_2676,N_29722,N_29924);
and UO_2677 (O_2677,N_29777,N_29953);
or UO_2678 (O_2678,N_29714,N_29942);
nor UO_2679 (O_2679,N_29878,N_29986);
and UO_2680 (O_2680,N_29969,N_29717);
nand UO_2681 (O_2681,N_29772,N_29843);
or UO_2682 (O_2682,N_29794,N_29978);
and UO_2683 (O_2683,N_29882,N_29990);
nor UO_2684 (O_2684,N_29757,N_29861);
or UO_2685 (O_2685,N_29924,N_29913);
and UO_2686 (O_2686,N_29848,N_29745);
or UO_2687 (O_2687,N_29960,N_29975);
xnor UO_2688 (O_2688,N_29820,N_29769);
and UO_2689 (O_2689,N_29944,N_29946);
and UO_2690 (O_2690,N_29750,N_29965);
xnor UO_2691 (O_2691,N_29815,N_29790);
xor UO_2692 (O_2692,N_29942,N_29710);
and UO_2693 (O_2693,N_29738,N_29929);
and UO_2694 (O_2694,N_29931,N_29703);
xnor UO_2695 (O_2695,N_29920,N_29879);
nor UO_2696 (O_2696,N_29973,N_29785);
xor UO_2697 (O_2697,N_29919,N_29744);
nand UO_2698 (O_2698,N_29902,N_29758);
or UO_2699 (O_2699,N_29731,N_29880);
nor UO_2700 (O_2700,N_29811,N_29777);
nor UO_2701 (O_2701,N_29878,N_29713);
nor UO_2702 (O_2702,N_29750,N_29789);
or UO_2703 (O_2703,N_29965,N_29837);
nand UO_2704 (O_2704,N_29983,N_29891);
and UO_2705 (O_2705,N_29723,N_29748);
or UO_2706 (O_2706,N_29991,N_29899);
or UO_2707 (O_2707,N_29768,N_29897);
and UO_2708 (O_2708,N_29836,N_29880);
xor UO_2709 (O_2709,N_29875,N_29710);
xnor UO_2710 (O_2710,N_29933,N_29893);
nand UO_2711 (O_2711,N_29712,N_29944);
nor UO_2712 (O_2712,N_29847,N_29898);
or UO_2713 (O_2713,N_29826,N_29725);
or UO_2714 (O_2714,N_29741,N_29990);
and UO_2715 (O_2715,N_29880,N_29722);
or UO_2716 (O_2716,N_29713,N_29897);
or UO_2717 (O_2717,N_29910,N_29834);
or UO_2718 (O_2718,N_29942,N_29924);
nand UO_2719 (O_2719,N_29997,N_29885);
and UO_2720 (O_2720,N_29870,N_29980);
or UO_2721 (O_2721,N_29813,N_29951);
nand UO_2722 (O_2722,N_29735,N_29820);
nand UO_2723 (O_2723,N_29916,N_29834);
or UO_2724 (O_2724,N_29973,N_29975);
nand UO_2725 (O_2725,N_29828,N_29711);
and UO_2726 (O_2726,N_29814,N_29788);
nor UO_2727 (O_2727,N_29728,N_29747);
xor UO_2728 (O_2728,N_29740,N_29939);
xnor UO_2729 (O_2729,N_29806,N_29926);
or UO_2730 (O_2730,N_29874,N_29722);
nor UO_2731 (O_2731,N_29789,N_29712);
xor UO_2732 (O_2732,N_29856,N_29776);
and UO_2733 (O_2733,N_29975,N_29768);
and UO_2734 (O_2734,N_29840,N_29997);
nand UO_2735 (O_2735,N_29886,N_29904);
nand UO_2736 (O_2736,N_29791,N_29878);
xor UO_2737 (O_2737,N_29855,N_29943);
or UO_2738 (O_2738,N_29931,N_29967);
xnor UO_2739 (O_2739,N_29767,N_29800);
or UO_2740 (O_2740,N_29757,N_29810);
nor UO_2741 (O_2741,N_29893,N_29996);
nor UO_2742 (O_2742,N_29993,N_29720);
nand UO_2743 (O_2743,N_29754,N_29936);
nand UO_2744 (O_2744,N_29738,N_29845);
nor UO_2745 (O_2745,N_29748,N_29911);
nor UO_2746 (O_2746,N_29835,N_29852);
xor UO_2747 (O_2747,N_29890,N_29842);
nor UO_2748 (O_2748,N_29916,N_29747);
xor UO_2749 (O_2749,N_29718,N_29811);
or UO_2750 (O_2750,N_29840,N_29750);
xnor UO_2751 (O_2751,N_29838,N_29963);
xnor UO_2752 (O_2752,N_29862,N_29957);
nand UO_2753 (O_2753,N_29721,N_29900);
nand UO_2754 (O_2754,N_29833,N_29962);
nand UO_2755 (O_2755,N_29892,N_29851);
nand UO_2756 (O_2756,N_29755,N_29850);
nand UO_2757 (O_2757,N_29908,N_29757);
nand UO_2758 (O_2758,N_29781,N_29903);
and UO_2759 (O_2759,N_29934,N_29775);
nand UO_2760 (O_2760,N_29853,N_29993);
nand UO_2761 (O_2761,N_29839,N_29880);
nand UO_2762 (O_2762,N_29713,N_29765);
xor UO_2763 (O_2763,N_29760,N_29740);
nor UO_2764 (O_2764,N_29958,N_29745);
or UO_2765 (O_2765,N_29707,N_29822);
nand UO_2766 (O_2766,N_29954,N_29809);
or UO_2767 (O_2767,N_29825,N_29792);
nand UO_2768 (O_2768,N_29779,N_29990);
nand UO_2769 (O_2769,N_29980,N_29741);
or UO_2770 (O_2770,N_29987,N_29814);
or UO_2771 (O_2771,N_29752,N_29995);
xor UO_2772 (O_2772,N_29802,N_29990);
xnor UO_2773 (O_2773,N_29837,N_29899);
nand UO_2774 (O_2774,N_29743,N_29740);
or UO_2775 (O_2775,N_29864,N_29953);
xnor UO_2776 (O_2776,N_29932,N_29895);
nor UO_2777 (O_2777,N_29868,N_29853);
nand UO_2778 (O_2778,N_29981,N_29958);
and UO_2779 (O_2779,N_29953,N_29784);
or UO_2780 (O_2780,N_29821,N_29818);
nand UO_2781 (O_2781,N_29837,N_29986);
or UO_2782 (O_2782,N_29818,N_29966);
xnor UO_2783 (O_2783,N_29740,N_29758);
nor UO_2784 (O_2784,N_29775,N_29903);
nor UO_2785 (O_2785,N_29804,N_29936);
or UO_2786 (O_2786,N_29779,N_29989);
nand UO_2787 (O_2787,N_29953,N_29971);
or UO_2788 (O_2788,N_29835,N_29944);
nand UO_2789 (O_2789,N_29744,N_29909);
nor UO_2790 (O_2790,N_29760,N_29891);
xnor UO_2791 (O_2791,N_29916,N_29856);
or UO_2792 (O_2792,N_29892,N_29902);
nand UO_2793 (O_2793,N_29861,N_29898);
nor UO_2794 (O_2794,N_29740,N_29938);
xnor UO_2795 (O_2795,N_29819,N_29884);
or UO_2796 (O_2796,N_29869,N_29911);
or UO_2797 (O_2797,N_29904,N_29879);
nand UO_2798 (O_2798,N_29798,N_29716);
nor UO_2799 (O_2799,N_29984,N_29970);
xor UO_2800 (O_2800,N_29792,N_29918);
and UO_2801 (O_2801,N_29786,N_29791);
and UO_2802 (O_2802,N_29730,N_29771);
xnor UO_2803 (O_2803,N_29831,N_29845);
or UO_2804 (O_2804,N_29808,N_29797);
and UO_2805 (O_2805,N_29812,N_29763);
and UO_2806 (O_2806,N_29876,N_29852);
nor UO_2807 (O_2807,N_29814,N_29913);
nor UO_2808 (O_2808,N_29991,N_29968);
and UO_2809 (O_2809,N_29802,N_29779);
xor UO_2810 (O_2810,N_29834,N_29899);
nor UO_2811 (O_2811,N_29847,N_29926);
nand UO_2812 (O_2812,N_29808,N_29834);
xor UO_2813 (O_2813,N_29790,N_29854);
and UO_2814 (O_2814,N_29736,N_29946);
or UO_2815 (O_2815,N_29892,N_29771);
and UO_2816 (O_2816,N_29896,N_29814);
and UO_2817 (O_2817,N_29980,N_29820);
and UO_2818 (O_2818,N_29783,N_29771);
and UO_2819 (O_2819,N_29991,N_29811);
nor UO_2820 (O_2820,N_29725,N_29894);
nor UO_2821 (O_2821,N_29923,N_29702);
or UO_2822 (O_2822,N_29869,N_29862);
xor UO_2823 (O_2823,N_29720,N_29853);
nor UO_2824 (O_2824,N_29878,N_29758);
nand UO_2825 (O_2825,N_29928,N_29892);
nand UO_2826 (O_2826,N_29721,N_29874);
nor UO_2827 (O_2827,N_29870,N_29825);
nor UO_2828 (O_2828,N_29940,N_29765);
or UO_2829 (O_2829,N_29826,N_29961);
xor UO_2830 (O_2830,N_29800,N_29958);
nor UO_2831 (O_2831,N_29791,N_29941);
nor UO_2832 (O_2832,N_29888,N_29786);
or UO_2833 (O_2833,N_29805,N_29766);
xor UO_2834 (O_2834,N_29873,N_29876);
nor UO_2835 (O_2835,N_29740,N_29943);
xnor UO_2836 (O_2836,N_29880,N_29884);
or UO_2837 (O_2837,N_29739,N_29976);
nor UO_2838 (O_2838,N_29943,N_29873);
xor UO_2839 (O_2839,N_29877,N_29730);
nand UO_2840 (O_2840,N_29887,N_29863);
nor UO_2841 (O_2841,N_29796,N_29712);
nand UO_2842 (O_2842,N_29741,N_29790);
or UO_2843 (O_2843,N_29756,N_29801);
nand UO_2844 (O_2844,N_29856,N_29964);
nand UO_2845 (O_2845,N_29848,N_29802);
and UO_2846 (O_2846,N_29785,N_29994);
or UO_2847 (O_2847,N_29837,N_29892);
nand UO_2848 (O_2848,N_29871,N_29955);
and UO_2849 (O_2849,N_29962,N_29821);
xor UO_2850 (O_2850,N_29754,N_29724);
and UO_2851 (O_2851,N_29814,N_29821);
nand UO_2852 (O_2852,N_29799,N_29884);
and UO_2853 (O_2853,N_29875,N_29928);
nand UO_2854 (O_2854,N_29863,N_29799);
nand UO_2855 (O_2855,N_29984,N_29871);
xnor UO_2856 (O_2856,N_29906,N_29931);
nor UO_2857 (O_2857,N_29771,N_29839);
and UO_2858 (O_2858,N_29759,N_29976);
xnor UO_2859 (O_2859,N_29935,N_29976);
xnor UO_2860 (O_2860,N_29924,N_29835);
nand UO_2861 (O_2861,N_29760,N_29960);
nand UO_2862 (O_2862,N_29954,N_29795);
or UO_2863 (O_2863,N_29753,N_29808);
nor UO_2864 (O_2864,N_29717,N_29791);
xor UO_2865 (O_2865,N_29886,N_29723);
or UO_2866 (O_2866,N_29835,N_29849);
nand UO_2867 (O_2867,N_29895,N_29970);
or UO_2868 (O_2868,N_29817,N_29965);
or UO_2869 (O_2869,N_29952,N_29877);
nand UO_2870 (O_2870,N_29724,N_29875);
xnor UO_2871 (O_2871,N_29962,N_29750);
nand UO_2872 (O_2872,N_29964,N_29787);
and UO_2873 (O_2873,N_29893,N_29859);
and UO_2874 (O_2874,N_29806,N_29897);
and UO_2875 (O_2875,N_29784,N_29865);
or UO_2876 (O_2876,N_29837,N_29828);
nand UO_2877 (O_2877,N_29961,N_29738);
nand UO_2878 (O_2878,N_29879,N_29959);
nor UO_2879 (O_2879,N_29790,N_29872);
nand UO_2880 (O_2880,N_29892,N_29826);
nor UO_2881 (O_2881,N_29711,N_29868);
or UO_2882 (O_2882,N_29853,N_29906);
xnor UO_2883 (O_2883,N_29779,N_29869);
and UO_2884 (O_2884,N_29993,N_29943);
xnor UO_2885 (O_2885,N_29933,N_29878);
or UO_2886 (O_2886,N_29932,N_29786);
nand UO_2887 (O_2887,N_29963,N_29765);
xor UO_2888 (O_2888,N_29813,N_29913);
and UO_2889 (O_2889,N_29872,N_29702);
xor UO_2890 (O_2890,N_29757,N_29987);
nand UO_2891 (O_2891,N_29962,N_29863);
and UO_2892 (O_2892,N_29767,N_29793);
xnor UO_2893 (O_2893,N_29980,N_29959);
or UO_2894 (O_2894,N_29954,N_29854);
or UO_2895 (O_2895,N_29975,N_29797);
nand UO_2896 (O_2896,N_29821,N_29781);
nand UO_2897 (O_2897,N_29759,N_29743);
nand UO_2898 (O_2898,N_29814,N_29973);
nor UO_2899 (O_2899,N_29785,N_29954);
nor UO_2900 (O_2900,N_29883,N_29979);
nor UO_2901 (O_2901,N_29998,N_29876);
or UO_2902 (O_2902,N_29988,N_29802);
xnor UO_2903 (O_2903,N_29813,N_29808);
nand UO_2904 (O_2904,N_29806,N_29851);
and UO_2905 (O_2905,N_29945,N_29943);
or UO_2906 (O_2906,N_29873,N_29980);
xor UO_2907 (O_2907,N_29920,N_29803);
or UO_2908 (O_2908,N_29945,N_29829);
nor UO_2909 (O_2909,N_29847,N_29749);
nor UO_2910 (O_2910,N_29971,N_29833);
nor UO_2911 (O_2911,N_29885,N_29768);
nand UO_2912 (O_2912,N_29714,N_29951);
and UO_2913 (O_2913,N_29767,N_29780);
and UO_2914 (O_2914,N_29736,N_29878);
xor UO_2915 (O_2915,N_29891,N_29714);
or UO_2916 (O_2916,N_29960,N_29984);
nand UO_2917 (O_2917,N_29719,N_29812);
nand UO_2918 (O_2918,N_29789,N_29724);
xor UO_2919 (O_2919,N_29715,N_29921);
nand UO_2920 (O_2920,N_29800,N_29747);
nand UO_2921 (O_2921,N_29852,N_29914);
xnor UO_2922 (O_2922,N_29827,N_29780);
or UO_2923 (O_2923,N_29827,N_29889);
nand UO_2924 (O_2924,N_29982,N_29788);
or UO_2925 (O_2925,N_29958,N_29824);
or UO_2926 (O_2926,N_29905,N_29891);
and UO_2927 (O_2927,N_29740,N_29838);
xor UO_2928 (O_2928,N_29794,N_29805);
or UO_2929 (O_2929,N_29715,N_29879);
nand UO_2930 (O_2930,N_29767,N_29801);
nor UO_2931 (O_2931,N_29858,N_29804);
or UO_2932 (O_2932,N_29784,N_29920);
and UO_2933 (O_2933,N_29874,N_29816);
nor UO_2934 (O_2934,N_29920,N_29832);
or UO_2935 (O_2935,N_29711,N_29888);
or UO_2936 (O_2936,N_29713,N_29790);
nand UO_2937 (O_2937,N_29757,N_29736);
nand UO_2938 (O_2938,N_29997,N_29726);
nor UO_2939 (O_2939,N_29957,N_29820);
or UO_2940 (O_2940,N_29815,N_29847);
xnor UO_2941 (O_2941,N_29809,N_29923);
and UO_2942 (O_2942,N_29952,N_29898);
and UO_2943 (O_2943,N_29937,N_29721);
and UO_2944 (O_2944,N_29940,N_29962);
nor UO_2945 (O_2945,N_29790,N_29873);
nor UO_2946 (O_2946,N_29855,N_29887);
nand UO_2947 (O_2947,N_29934,N_29768);
and UO_2948 (O_2948,N_29861,N_29880);
xor UO_2949 (O_2949,N_29952,N_29931);
nor UO_2950 (O_2950,N_29896,N_29946);
and UO_2951 (O_2951,N_29855,N_29982);
and UO_2952 (O_2952,N_29930,N_29907);
nor UO_2953 (O_2953,N_29745,N_29985);
and UO_2954 (O_2954,N_29955,N_29880);
xnor UO_2955 (O_2955,N_29740,N_29837);
or UO_2956 (O_2956,N_29839,N_29856);
xor UO_2957 (O_2957,N_29767,N_29731);
nand UO_2958 (O_2958,N_29910,N_29844);
nor UO_2959 (O_2959,N_29804,N_29887);
nor UO_2960 (O_2960,N_29818,N_29971);
nand UO_2961 (O_2961,N_29735,N_29729);
nor UO_2962 (O_2962,N_29983,N_29914);
nor UO_2963 (O_2963,N_29922,N_29957);
or UO_2964 (O_2964,N_29930,N_29891);
or UO_2965 (O_2965,N_29847,N_29807);
xnor UO_2966 (O_2966,N_29870,N_29886);
xnor UO_2967 (O_2967,N_29753,N_29978);
nand UO_2968 (O_2968,N_29962,N_29992);
and UO_2969 (O_2969,N_29776,N_29951);
and UO_2970 (O_2970,N_29989,N_29993);
nand UO_2971 (O_2971,N_29829,N_29927);
or UO_2972 (O_2972,N_29990,N_29747);
or UO_2973 (O_2973,N_29821,N_29769);
xor UO_2974 (O_2974,N_29744,N_29841);
nor UO_2975 (O_2975,N_29852,N_29976);
nor UO_2976 (O_2976,N_29991,N_29935);
and UO_2977 (O_2977,N_29972,N_29885);
nor UO_2978 (O_2978,N_29880,N_29829);
and UO_2979 (O_2979,N_29938,N_29862);
xnor UO_2980 (O_2980,N_29881,N_29848);
or UO_2981 (O_2981,N_29967,N_29908);
and UO_2982 (O_2982,N_29835,N_29839);
xnor UO_2983 (O_2983,N_29996,N_29844);
nor UO_2984 (O_2984,N_29789,N_29923);
and UO_2985 (O_2985,N_29968,N_29875);
and UO_2986 (O_2986,N_29826,N_29740);
nor UO_2987 (O_2987,N_29745,N_29707);
and UO_2988 (O_2988,N_29969,N_29732);
and UO_2989 (O_2989,N_29800,N_29804);
or UO_2990 (O_2990,N_29777,N_29850);
nor UO_2991 (O_2991,N_29819,N_29921);
and UO_2992 (O_2992,N_29882,N_29907);
and UO_2993 (O_2993,N_29985,N_29948);
and UO_2994 (O_2994,N_29787,N_29821);
nand UO_2995 (O_2995,N_29825,N_29925);
and UO_2996 (O_2996,N_29848,N_29809);
xor UO_2997 (O_2997,N_29950,N_29827);
or UO_2998 (O_2998,N_29778,N_29938);
nand UO_2999 (O_2999,N_29704,N_29994);
nand UO_3000 (O_3000,N_29754,N_29715);
or UO_3001 (O_3001,N_29766,N_29797);
nor UO_3002 (O_3002,N_29700,N_29833);
nor UO_3003 (O_3003,N_29984,N_29841);
nor UO_3004 (O_3004,N_29904,N_29779);
nand UO_3005 (O_3005,N_29942,N_29888);
nor UO_3006 (O_3006,N_29957,N_29733);
nand UO_3007 (O_3007,N_29967,N_29706);
xnor UO_3008 (O_3008,N_29749,N_29728);
or UO_3009 (O_3009,N_29767,N_29879);
and UO_3010 (O_3010,N_29716,N_29890);
and UO_3011 (O_3011,N_29945,N_29864);
xor UO_3012 (O_3012,N_29876,N_29895);
nor UO_3013 (O_3013,N_29715,N_29998);
nand UO_3014 (O_3014,N_29970,N_29997);
and UO_3015 (O_3015,N_29708,N_29768);
xnor UO_3016 (O_3016,N_29711,N_29999);
and UO_3017 (O_3017,N_29964,N_29955);
xor UO_3018 (O_3018,N_29853,N_29832);
nand UO_3019 (O_3019,N_29969,N_29902);
nor UO_3020 (O_3020,N_29794,N_29937);
nand UO_3021 (O_3021,N_29821,N_29847);
xor UO_3022 (O_3022,N_29750,N_29865);
nor UO_3023 (O_3023,N_29772,N_29877);
or UO_3024 (O_3024,N_29973,N_29863);
nor UO_3025 (O_3025,N_29925,N_29997);
nor UO_3026 (O_3026,N_29940,N_29718);
nand UO_3027 (O_3027,N_29734,N_29875);
nand UO_3028 (O_3028,N_29866,N_29764);
nor UO_3029 (O_3029,N_29838,N_29771);
and UO_3030 (O_3030,N_29973,N_29826);
nand UO_3031 (O_3031,N_29850,N_29712);
nor UO_3032 (O_3032,N_29914,N_29939);
xnor UO_3033 (O_3033,N_29934,N_29835);
or UO_3034 (O_3034,N_29837,N_29816);
xnor UO_3035 (O_3035,N_29775,N_29938);
and UO_3036 (O_3036,N_29932,N_29804);
and UO_3037 (O_3037,N_29972,N_29889);
nor UO_3038 (O_3038,N_29838,N_29988);
and UO_3039 (O_3039,N_29788,N_29844);
or UO_3040 (O_3040,N_29752,N_29831);
xor UO_3041 (O_3041,N_29955,N_29820);
nor UO_3042 (O_3042,N_29755,N_29938);
xor UO_3043 (O_3043,N_29851,N_29918);
nand UO_3044 (O_3044,N_29861,N_29922);
or UO_3045 (O_3045,N_29985,N_29731);
nand UO_3046 (O_3046,N_29729,N_29712);
nor UO_3047 (O_3047,N_29975,N_29881);
xor UO_3048 (O_3048,N_29880,N_29748);
nor UO_3049 (O_3049,N_29717,N_29836);
or UO_3050 (O_3050,N_29711,N_29778);
nor UO_3051 (O_3051,N_29951,N_29965);
nor UO_3052 (O_3052,N_29821,N_29950);
and UO_3053 (O_3053,N_29756,N_29936);
or UO_3054 (O_3054,N_29943,N_29821);
nor UO_3055 (O_3055,N_29742,N_29791);
or UO_3056 (O_3056,N_29919,N_29982);
and UO_3057 (O_3057,N_29894,N_29953);
xor UO_3058 (O_3058,N_29721,N_29768);
and UO_3059 (O_3059,N_29971,N_29828);
and UO_3060 (O_3060,N_29985,N_29809);
xnor UO_3061 (O_3061,N_29725,N_29780);
nand UO_3062 (O_3062,N_29900,N_29982);
and UO_3063 (O_3063,N_29718,N_29839);
xnor UO_3064 (O_3064,N_29738,N_29965);
nor UO_3065 (O_3065,N_29822,N_29896);
nand UO_3066 (O_3066,N_29913,N_29744);
nand UO_3067 (O_3067,N_29857,N_29898);
and UO_3068 (O_3068,N_29863,N_29824);
xnor UO_3069 (O_3069,N_29854,N_29822);
nor UO_3070 (O_3070,N_29720,N_29906);
nand UO_3071 (O_3071,N_29799,N_29967);
and UO_3072 (O_3072,N_29754,N_29954);
xor UO_3073 (O_3073,N_29906,N_29872);
nand UO_3074 (O_3074,N_29811,N_29713);
xor UO_3075 (O_3075,N_29892,N_29957);
nand UO_3076 (O_3076,N_29764,N_29925);
nor UO_3077 (O_3077,N_29784,N_29991);
xnor UO_3078 (O_3078,N_29944,N_29751);
nand UO_3079 (O_3079,N_29975,N_29934);
or UO_3080 (O_3080,N_29821,N_29740);
and UO_3081 (O_3081,N_29991,N_29949);
nor UO_3082 (O_3082,N_29705,N_29881);
or UO_3083 (O_3083,N_29840,N_29707);
xnor UO_3084 (O_3084,N_29939,N_29718);
and UO_3085 (O_3085,N_29787,N_29817);
nand UO_3086 (O_3086,N_29856,N_29743);
xnor UO_3087 (O_3087,N_29773,N_29711);
xor UO_3088 (O_3088,N_29959,N_29764);
xnor UO_3089 (O_3089,N_29836,N_29943);
and UO_3090 (O_3090,N_29721,N_29824);
nor UO_3091 (O_3091,N_29705,N_29824);
xnor UO_3092 (O_3092,N_29903,N_29933);
nor UO_3093 (O_3093,N_29875,N_29800);
or UO_3094 (O_3094,N_29754,N_29914);
and UO_3095 (O_3095,N_29997,N_29930);
and UO_3096 (O_3096,N_29896,N_29778);
nand UO_3097 (O_3097,N_29821,N_29748);
and UO_3098 (O_3098,N_29892,N_29794);
xnor UO_3099 (O_3099,N_29885,N_29905);
nor UO_3100 (O_3100,N_29820,N_29961);
nor UO_3101 (O_3101,N_29850,N_29815);
nor UO_3102 (O_3102,N_29973,N_29799);
or UO_3103 (O_3103,N_29803,N_29878);
xnor UO_3104 (O_3104,N_29808,N_29979);
nand UO_3105 (O_3105,N_29703,N_29864);
nand UO_3106 (O_3106,N_29875,N_29807);
or UO_3107 (O_3107,N_29883,N_29767);
nor UO_3108 (O_3108,N_29847,N_29865);
xnor UO_3109 (O_3109,N_29915,N_29938);
nand UO_3110 (O_3110,N_29871,N_29905);
xnor UO_3111 (O_3111,N_29710,N_29769);
or UO_3112 (O_3112,N_29915,N_29826);
xor UO_3113 (O_3113,N_29838,N_29833);
or UO_3114 (O_3114,N_29738,N_29930);
or UO_3115 (O_3115,N_29971,N_29800);
nand UO_3116 (O_3116,N_29796,N_29858);
nor UO_3117 (O_3117,N_29971,N_29997);
and UO_3118 (O_3118,N_29950,N_29880);
and UO_3119 (O_3119,N_29780,N_29885);
xor UO_3120 (O_3120,N_29974,N_29825);
nand UO_3121 (O_3121,N_29866,N_29842);
nand UO_3122 (O_3122,N_29804,N_29905);
and UO_3123 (O_3123,N_29786,N_29868);
xor UO_3124 (O_3124,N_29839,N_29785);
nand UO_3125 (O_3125,N_29993,N_29731);
xor UO_3126 (O_3126,N_29818,N_29990);
nand UO_3127 (O_3127,N_29720,N_29743);
and UO_3128 (O_3128,N_29801,N_29961);
or UO_3129 (O_3129,N_29946,N_29832);
nand UO_3130 (O_3130,N_29870,N_29942);
nand UO_3131 (O_3131,N_29929,N_29831);
and UO_3132 (O_3132,N_29820,N_29878);
or UO_3133 (O_3133,N_29883,N_29740);
or UO_3134 (O_3134,N_29915,N_29861);
or UO_3135 (O_3135,N_29893,N_29957);
and UO_3136 (O_3136,N_29809,N_29901);
nand UO_3137 (O_3137,N_29966,N_29884);
or UO_3138 (O_3138,N_29718,N_29794);
xor UO_3139 (O_3139,N_29935,N_29716);
xor UO_3140 (O_3140,N_29922,N_29989);
nor UO_3141 (O_3141,N_29911,N_29976);
nor UO_3142 (O_3142,N_29802,N_29927);
or UO_3143 (O_3143,N_29913,N_29888);
nand UO_3144 (O_3144,N_29701,N_29956);
xnor UO_3145 (O_3145,N_29779,N_29831);
nand UO_3146 (O_3146,N_29975,N_29984);
nand UO_3147 (O_3147,N_29702,N_29792);
nor UO_3148 (O_3148,N_29741,N_29833);
and UO_3149 (O_3149,N_29828,N_29957);
xnor UO_3150 (O_3150,N_29753,N_29799);
or UO_3151 (O_3151,N_29905,N_29881);
xor UO_3152 (O_3152,N_29731,N_29966);
or UO_3153 (O_3153,N_29704,N_29784);
and UO_3154 (O_3154,N_29792,N_29776);
or UO_3155 (O_3155,N_29731,N_29781);
nor UO_3156 (O_3156,N_29851,N_29944);
or UO_3157 (O_3157,N_29904,N_29944);
and UO_3158 (O_3158,N_29926,N_29823);
nor UO_3159 (O_3159,N_29970,N_29876);
and UO_3160 (O_3160,N_29882,N_29791);
and UO_3161 (O_3161,N_29820,N_29929);
nor UO_3162 (O_3162,N_29897,N_29934);
or UO_3163 (O_3163,N_29748,N_29841);
nand UO_3164 (O_3164,N_29788,N_29745);
nor UO_3165 (O_3165,N_29976,N_29722);
nand UO_3166 (O_3166,N_29779,N_29899);
and UO_3167 (O_3167,N_29903,N_29957);
nand UO_3168 (O_3168,N_29949,N_29844);
xor UO_3169 (O_3169,N_29895,N_29911);
or UO_3170 (O_3170,N_29896,N_29866);
nor UO_3171 (O_3171,N_29818,N_29914);
nand UO_3172 (O_3172,N_29884,N_29984);
or UO_3173 (O_3173,N_29896,N_29759);
xnor UO_3174 (O_3174,N_29896,N_29996);
nand UO_3175 (O_3175,N_29839,N_29999);
nand UO_3176 (O_3176,N_29857,N_29881);
nor UO_3177 (O_3177,N_29701,N_29781);
xnor UO_3178 (O_3178,N_29927,N_29804);
nor UO_3179 (O_3179,N_29818,N_29848);
or UO_3180 (O_3180,N_29889,N_29981);
or UO_3181 (O_3181,N_29766,N_29992);
nand UO_3182 (O_3182,N_29884,N_29836);
or UO_3183 (O_3183,N_29847,N_29709);
nand UO_3184 (O_3184,N_29851,N_29715);
nand UO_3185 (O_3185,N_29749,N_29975);
xnor UO_3186 (O_3186,N_29825,N_29808);
and UO_3187 (O_3187,N_29956,N_29949);
nand UO_3188 (O_3188,N_29929,N_29821);
nor UO_3189 (O_3189,N_29867,N_29734);
or UO_3190 (O_3190,N_29873,N_29802);
xnor UO_3191 (O_3191,N_29929,N_29824);
or UO_3192 (O_3192,N_29757,N_29947);
xor UO_3193 (O_3193,N_29934,N_29830);
xnor UO_3194 (O_3194,N_29773,N_29945);
nand UO_3195 (O_3195,N_29996,N_29856);
nor UO_3196 (O_3196,N_29991,N_29997);
nand UO_3197 (O_3197,N_29779,N_29896);
or UO_3198 (O_3198,N_29901,N_29795);
nor UO_3199 (O_3199,N_29909,N_29966);
or UO_3200 (O_3200,N_29879,N_29909);
or UO_3201 (O_3201,N_29864,N_29924);
xnor UO_3202 (O_3202,N_29781,N_29714);
xor UO_3203 (O_3203,N_29875,N_29840);
nor UO_3204 (O_3204,N_29779,N_29796);
nor UO_3205 (O_3205,N_29820,N_29724);
or UO_3206 (O_3206,N_29946,N_29950);
nor UO_3207 (O_3207,N_29955,N_29870);
nor UO_3208 (O_3208,N_29814,N_29917);
or UO_3209 (O_3209,N_29744,N_29854);
or UO_3210 (O_3210,N_29889,N_29892);
xnor UO_3211 (O_3211,N_29854,N_29815);
xor UO_3212 (O_3212,N_29983,N_29957);
nor UO_3213 (O_3213,N_29952,N_29852);
or UO_3214 (O_3214,N_29841,N_29976);
and UO_3215 (O_3215,N_29891,N_29803);
or UO_3216 (O_3216,N_29850,N_29912);
and UO_3217 (O_3217,N_29805,N_29938);
or UO_3218 (O_3218,N_29956,N_29901);
nand UO_3219 (O_3219,N_29804,N_29827);
and UO_3220 (O_3220,N_29862,N_29977);
nor UO_3221 (O_3221,N_29859,N_29906);
or UO_3222 (O_3222,N_29792,N_29815);
xor UO_3223 (O_3223,N_29998,N_29827);
and UO_3224 (O_3224,N_29895,N_29905);
nand UO_3225 (O_3225,N_29881,N_29987);
xor UO_3226 (O_3226,N_29813,N_29940);
and UO_3227 (O_3227,N_29806,N_29828);
and UO_3228 (O_3228,N_29901,N_29914);
and UO_3229 (O_3229,N_29874,N_29957);
xnor UO_3230 (O_3230,N_29764,N_29805);
xnor UO_3231 (O_3231,N_29908,N_29769);
xnor UO_3232 (O_3232,N_29726,N_29902);
or UO_3233 (O_3233,N_29813,N_29931);
nand UO_3234 (O_3234,N_29800,N_29846);
nor UO_3235 (O_3235,N_29770,N_29913);
nand UO_3236 (O_3236,N_29871,N_29940);
or UO_3237 (O_3237,N_29825,N_29782);
nand UO_3238 (O_3238,N_29781,N_29861);
and UO_3239 (O_3239,N_29854,N_29948);
nor UO_3240 (O_3240,N_29983,N_29773);
and UO_3241 (O_3241,N_29846,N_29772);
or UO_3242 (O_3242,N_29876,N_29807);
nor UO_3243 (O_3243,N_29763,N_29944);
nand UO_3244 (O_3244,N_29874,N_29934);
nand UO_3245 (O_3245,N_29782,N_29755);
or UO_3246 (O_3246,N_29900,N_29752);
and UO_3247 (O_3247,N_29790,N_29892);
or UO_3248 (O_3248,N_29740,N_29797);
and UO_3249 (O_3249,N_29820,N_29801);
nor UO_3250 (O_3250,N_29987,N_29802);
nor UO_3251 (O_3251,N_29755,N_29702);
nand UO_3252 (O_3252,N_29983,N_29710);
xnor UO_3253 (O_3253,N_29702,N_29815);
and UO_3254 (O_3254,N_29752,N_29840);
or UO_3255 (O_3255,N_29873,N_29752);
nor UO_3256 (O_3256,N_29762,N_29966);
and UO_3257 (O_3257,N_29869,N_29893);
nand UO_3258 (O_3258,N_29813,N_29858);
or UO_3259 (O_3259,N_29831,N_29972);
and UO_3260 (O_3260,N_29777,N_29742);
xnor UO_3261 (O_3261,N_29941,N_29701);
nand UO_3262 (O_3262,N_29876,N_29858);
and UO_3263 (O_3263,N_29710,N_29764);
and UO_3264 (O_3264,N_29884,N_29765);
or UO_3265 (O_3265,N_29722,N_29708);
nand UO_3266 (O_3266,N_29914,N_29903);
xnor UO_3267 (O_3267,N_29837,N_29869);
nand UO_3268 (O_3268,N_29762,N_29835);
and UO_3269 (O_3269,N_29922,N_29765);
xnor UO_3270 (O_3270,N_29997,N_29916);
nand UO_3271 (O_3271,N_29940,N_29911);
nor UO_3272 (O_3272,N_29931,N_29888);
xnor UO_3273 (O_3273,N_29851,N_29931);
or UO_3274 (O_3274,N_29758,N_29844);
xor UO_3275 (O_3275,N_29883,N_29820);
and UO_3276 (O_3276,N_29726,N_29724);
and UO_3277 (O_3277,N_29757,N_29934);
nand UO_3278 (O_3278,N_29786,N_29752);
or UO_3279 (O_3279,N_29902,N_29924);
nor UO_3280 (O_3280,N_29843,N_29883);
and UO_3281 (O_3281,N_29853,N_29809);
and UO_3282 (O_3282,N_29958,N_29832);
and UO_3283 (O_3283,N_29702,N_29929);
nor UO_3284 (O_3284,N_29949,N_29767);
xor UO_3285 (O_3285,N_29870,N_29718);
nor UO_3286 (O_3286,N_29965,N_29972);
or UO_3287 (O_3287,N_29785,N_29812);
or UO_3288 (O_3288,N_29808,N_29718);
nand UO_3289 (O_3289,N_29773,N_29815);
xor UO_3290 (O_3290,N_29849,N_29763);
nand UO_3291 (O_3291,N_29968,N_29717);
xor UO_3292 (O_3292,N_29891,N_29878);
xor UO_3293 (O_3293,N_29733,N_29812);
nor UO_3294 (O_3294,N_29952,N_29955);
or UO_3295 (O_3295,N_29947,N_29946);
nor UO_3296 (O_3296,N_29983,N_29833);
or UO_3297 (O_3297,N_29781,N_29968);
and UO_3298 (O_3298,N_29947,N_29815);
xnor UO_3299 (O_3299,N_29724,N_29880);
or UO_3300 (O_3300,N_29889,N_29808);
nand UO_3301 (O_3301,N_29882,N_29706);
and UO_3302 (O_3302,N_29970,N_29769);
or UO_3303 (O_3303,N_29906,N_29917);
nor UO_3304 (O_3304,N_29876,N_29821);
and UO_3305 (O_3305,N_29715,N_29807);
xnor UO_3306 (O_3306,N_29840,N_29893);
or UO_3307 (O_3307,N_29732,N_29859);
nand UO_3308 (O_3308,N_29762,N_29947);
nor UO_3309 (O_3309,N_29740,N_29913);
nor UO_3310 (O_3310,N_29952,N_29799);
nor UO_3311 (O_3311,N_29851,N_29829);
xor UO_3312 (O_3312,N_29802,N_29949);
xor UO_3313 (O_3313,N_29815,N_29735);
nand UO_3314 (O_3314,N_29942,N_29747);
or UO_3315 (O_3315,N_29859,N_29786);
nor UO_3316 (O_3316,N_29957,N_29951);
nor UO_3317 (O_3317,N_29758,N_29807);
nor UO_3318 (O_3318,N_29720,N_29953);
nor UO_3319 (O_3319,N_29954,N_29970);
nand UO_3320 (O_3320,N_29863,N_29751);
and UO_3321 (O_3321,N_29807,N_29808);
xnor UO_3322 (O_3322,N_29947,N_29937);
or UO_3323 (O_3323,N_29809,N_29721);
nand UO_3324 (O_3324,N_29909,N_29970);
nor UO_3325 (O_3325,N_29843,N_29779);
xnor UO_3326 (O_3326,N_29722,N_29776);
or UO_3327 (O_3327,N_29766,N_29816);
xnor UO_3328 (O_3328,N_29719,N_29759);
xor UO_3329 (O_3329,N_29940,N_29975);
or UO_3330 (O_3330,N_29739,N_29771);
nor UO_3331 (O_3331,N_29961,N_29735);
nor UO_3332 (O_3332,N_29784,N_29842);
and UO_3333 (O_3333,N_29908,N_29734);
nand UO_3334 (O_3334,N_29975,N_29978);
nor UO_3335 (O_3335,N_29706,N_29737);
xor UO_3336 (O_3336,N_29700,N_29828);
nor UO_3337 (O_3337,N_29994,N_29840);
xnor UO_3338 (O_3338,N_29715,N_29925);
and UO_3339 (O_3339,N_29745,N_29845);
nor UO_3340 (O_3340,N_29717,N_29771);
nor UO_3341 (O_3341,N_29757,N_29747);
xor UO_3342 (O_3342,N_29931,N_29903);
or UO_3343 (O_3343,N_29823,N_29779);
and UO_3344 (O_3344,N_29784,N_29743);
nor UO_3345 (O_3345,N_29703,N_29876);
or UO_3346 (O_3346,N_29849,N_29806);
and UO_3347 (O_3347,N_29828,N_29848);
or UO_3348 (O_3348,N_29711,N_29781);
nor UO_3349 (O_3349,N_29819,N_29861);
and UO_3350 (O_3350,N_29941,N_29917);
nor UO_3351 (O_3351,N_29902,N_29761);
xnor UO_3352 (O_3352,N_29958,N_29842);
nor UO_3353 (O_3353,N_29803,N_29827);
nand UO_3354 (O_3354,N_29985,N_29866);
xnor UO_3355 (O_3355,N_29992,N_29874);
xnor UO_3356 (O_3356,N_29929,N_29717);
xor UO_3357 (O_3357,N_29797,N_29802);
nand UO_3358 (O_3358,N_29867,N_29759);
and UO_3359 (O_3359,N_29841,N_29941);
or UO_3360 (O_3360,N_29941,N_29919);
xnor UO_3361 (O_3361,N_29734,N_29722);
or UO_3362 (O_3362,N_29882,N_29964);
nand UO_3363 (O_3363,N_29823,N_29874);
or UO_3364 (O_3364,N_29898,N_29733);
or UO_3365 (O_3365,N_29753,N_29716);
or UO_3366 (O_3366,N_29981,N_29864);
nor UO_3367 (O_3367,N_29753,N_29718);
xnor UO_3368 (O_3368,N_29937,N_29881);
nor UO_3369 (O_3369,N_29981,N_29988);
or UO_3370 (O_3370,N_29764,N_29716);
and UO_3371 (O_3371,N_29762,N_29822);
or UO_3372 (O_3372,N_29987,N_29941);
xnor UO_3373 (O_3373,N_29946,N_29807);
nand UO_3374 (O_3374,N_29822,N_29753);
and UO_3375 (O_3375,N_29811,N_29735);
xor UO_3376 (O_3376,N_29953,N_29903);
or UO_3377 (O_3377,N_29939,N_29767);
nor UO_3378 (O_3378,N_29711,N_29950);
nor UO_3379 (O_3379,N_29742,N_29850);
nor UO_3380 (O_3380,N_29826,N_29921);
nand UO_3381 (O_3381,N_29705,N_29772);
nand UO_3382 (O_3382,N_29735,N_29986);
nand UO_3383 (O_3383,N_29916,N_29978);
and UO_3384 (O_3384,N_29708,N_29952);
nor UO_3385 (O_3385,N_29877,N_29780);
xnor UO_3386 (O_3386,N_29840,N_29761);
nand UO_3387 (O_3387,N_29860,N_29951);
and UO_3388 (O_3388,N_29764,N_29823);
nor UO_3389 (O_3389,N_29888,N_29785);
nand UO_3390 (O_3390,N_29965,N_29883);
nand UO_3391 (O_3391,N_29976,N_29800);
or UO_3392 (O_3392,N_29754,N_29716);
and UO_3393 (O_3393,N_29876,N_29761);
xor UO_3394 (O_3394,N_29823,N_29722);
nand UO_3395 (O_3395,N_29758,N_29971);
nand UO_3396 (O_3396,N_29731,N_29720);
xnor UO_3397 (O_3397,N_29825,N_29705);
xnor UO_3398 (O_3398,N_29952,N_29903);
xnor UO_3399 (O_3399,N_29732,N_29714);
nor UO_3400 (O_3400,N_29958,N_29993);
nand UO_3401 (O_3401,N_29969,N_29706);
nand UO_3402 (O_3402,N_29789,N_29759);
or UO_3403 (O_3403,N_29861,N_29990);
and UO_3404 (O_3404,N_29844,N_29932);
or UO_3405 (O_3405,N_29970,N_29870);
and UO_3406 (O_3406,N_29952,N_29717);
or UO_3407 (O_3407,N_29914,N_29825);
nand UO_3408 (O_3408,N_29882,N_29731);
xor UO_3409 (O_3409,N_29957,N_29943);
xor UO_3410 (O_3410,N_29824,N_29734);
xnor UO_3411 (O_3411,N_29929,N_29857);
and UO_3412 (O_3412,N_29989,N_29744);
nor UO_3413 (O_3413,N_29875,N_29935);
and UO_3414 (O_3414,N_29987,N_29983);
nor UO_3415 (O_3415,N_29841,N_29783);
nor UO_3416 (O_3416,N_29746,N_29999);
and UO_3417 (O_3417,N_29712,N_29989);
and UO_3418 (O_3418,N_29716,N_29821);
xnor UO_3419 (O_3419,N_29804,N_29769);
nand UO_3420 (O_3420,N_29704,N_29769);
xnor UO_3421 (O_3421,N_29999,N_29964);
nand UO_3422 (O_3422,N_29714,N_29997);
and UO_3423 (O_3423,N_29722,N_29897);
or UO_3424 (O_3424,N_29776,N_29885);
nand UO_3425 (O_3425,N_29929,N_29851);
and UO_3426 (O_3426,N_29981,N_29978);
nand UO_3427 (O_3427,N_29989,N_29846);
nor UO_3428 (O_3428,N_29878,N_29834);
nor UO_3429 (O_3429,N_29903,N_29772);
or UO_3430 (O_3430,N_29787,N_29759);
xnor UO_3431 (O_3431,N_29834,N_29893);
and UO_3432 (O_3432,N_29957,N_29816);
xor UO_3433 (O_3433,N_29797,N_29887);
nor UO_3434 (O_3434,N_29962,N_29960);
or UO_3435 (O_3435,N_29753,N_29778);
nor UO_3436 (O_3436,N_29814,N_29727);
nand UO_3437 (O_3437,N_29982,N_29834);
xor UO_3438 (O_3438,N_29739,N_29870);
xor UO_3439 (O_3439,N_29769,N_29749);
xor UO_3440 (O_3440,N_29717,N_29828);
xor UO_3441 (O_3441,N_29857,N_29967);
or UO_3442 (O_3442,N_29783,N_29762);
nand UO_3443 (O_3443,N_29797,N_29858);
nor UO_3444 (O_3444,N_29767,N_29837);
nor UO_3445 (O_3445,N_29823,N_29993);
xnor UO_3446 (O_3446,N_29717,N_29918);
xnor UO_3447 (O_3447,N_29924,N_29850);
nor UO_3448 (O_3448,N_29761,N_29795);
xor UO_3449 (O_3449,N_29896,N_29898);
and UO_3450 (O_3450,N_29700,N_29896);
and UO_3451 (O_3451,N_29945,N_29881);
xnor UO_3452 (O_3452,N_29911,N_29962);
nor UO_3453 (O_3453,N_29948,N_29941);
nor UO_3454 (O_3454,N_29839,N_29981);
or UO_3455 (O_3455,N_29893,N_29952);
or UO_3456 (O_3456,N_29700,N_29851);
nand UO_3457 (O_3457,N_29733,N_29849);
xor UO_3458 (O_3458,N_29905,N_29870);
nor UO_3459 (O_3459,N_29905,N_29830);
nand UO_3460 (O_3460,N_29820,N_29876);
or UO_3461 (O_3461,N_29867,N_29994);
or UO_3462 (O_3462,N_29829,N_29863);
or UO_3463 (O_3463,N_29905,N_29835);
nand UO_3464 (O_3464,N_29855,N_29820);
nor UO_3465 (O_3465,N_29889,N_29963);
nor UO_3466 (O_3466,N_29823,N_29940);
nand UO_3467 (O_3467,N_29778,N_29827);
xor UO_3468 (O_3468,N_29749,N_29990);
or UO_3469 (O_3469,N_29856,N_29973);
nor UO_3470 (O_3470,N_29748,N_29902);
nand UO_3471 (O_3471,N_29879,N_29882);
xor UO_3472 (O_3472,N_29731,N_29819);
or UO_3473 (O_3473,N_29814,N_29826);
nor UO_3474 (O_3474,N_29769,N_29962);
and UO_3475 (O_3475,N_29953,N_29966);
and UO_3476 (O_3476,N_29996,N_29925);
nor UO_3477 (O_3477,N_29878,N_29876);
nor UO_3478 (O_3478,N_29893,N_29715);
or UO_3479 (O_3479,N_29877,N_29831);
nor UO_3480 (O_3480,N_29990,N_29832);
xnor UO_3481 (O_3481,N_29755,N_29729);
xor UO_3482 (O_3482,N_29842,N_29802);
nand UO_3483 (O_3483,N_29879,N_29788);
or UO_3484 (O_3484,N_29717,N_29727);
and UO_3485 (O_3485,N_29922,N_29862);
and UO_3486 (O_3486,N_29753,N_29731);
xnor UO_3487 (O_3487,N_29739,N_29831);
xor UO_3488 (O_3488,N_29769,N_29910);
and UO_3489 (O_3489,N_29880,N_29879);
xnor UO_3490 (O_3490,N_29885,N_29930);
and UO_3491 (O_3491,N_29915,N_29701);
and UO_3492 (O_3492,N_29967,N_29966);
or UO_3493 (O_3493,N_29781,N_29736);
or UO_3494 (O_3494,N_29992,N_29932);
and UO_3495 (O_3495,N_29913,N_29784);
and UO_3496 (O_3496,N_29967,N_29922);
or UO_3497 (O_3497,N_29725,N_29884);
nor UO_3498 (O_3498,N_29986,N_29894);
and UO_3499 (O_3499,N_29814,N_29838);
endmodule