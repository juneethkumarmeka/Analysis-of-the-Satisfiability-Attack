module basic_5000_50000_5000_10_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_303,In_2742);
or U1 (N_1,In_796,In_4900);
nor U2 (N_2,In_2523,In_2243);
and U3 (N_3,In_3568,In_378);
or U4 (N_4,In_310,In_3029);
xor U5 (N_5,In_1072,In_2750);
nand U6 (N_6,In_2337,In_4462);
nor U7 (N_7,In_4912,In_1316);
nor U8 (N_8,In_343,In_581);
nor U9 (N_9,In_3686,In_144);
xor U10 (N_10,In_3747,In_464);
nand U11 (N_11,In_4944,In_3595);
nor U12 (N_12,In_4114,In_4987);
nand U13 (N_13,In_547,In_119);
or U14 (N_14,In_4608,In_1881);
nor U15 (N_15,In_4202,In_2648);
nand U16 (N_16,In_2514,In_1825);
xnor U17 (N_17,In_4057,In_2776);
or U18 (N_18,In_1475,In_2618);
nor U19 (N_19,In_2864,In_1957);
nor U20 (N_20,In_3063,In_4730);
xor U21 (N_21,In_1396,In_1174);
or U22 (N_22,In_438,In_4668);
and U23 (N_23,In_1867,In_2660);
or U24 (N_24,In_103,In_4731);
xnor U25 (N_25,In_1462,In_4161);
nand U26 (N_26,In_593,In_64);
and U27 (N_27,In_4620,In_1077);
nor U28 (N_28,In_3275,In_2096);
or U29 (N_29,In_3477,In_430);
nand U30 (N_30,In_3114,In_3690);
nor U31 (N_31,In_4431,In_4934);
or U32 (N_32,In_1736,In_1169);
xor U33 (N_33,In_3535,In_1635);
and U34 (N_34,In_4818,In_2814);
and U35 (N_35,In_4226,In_4998);
and U36 (N_36,In_3195,In_314);
and U37 (N_37,In_1468,In_3427);
or U38 (N_38,In_758,In_8);
or U39 (N_39,In_1641,In_889);
or U40 (N_40,In_179,In_1719);
or U41 (N_41,In_465,In_3494);
nand U42 (N_42,In_3046,In_1677);
and U43 (N_43,In_1019,In_1424);
nor U44 (N_44,In_2909,In_995);
nand U45 (N_45,In_1243,In_4747);
nand U46 (N_46,In_2334,In_3077);
nor U47 (N_47,In_2710,In_281);
xor U48 (N_48,In_3881,In_4243);
nand U49 (N_49,In_2822,In_3167);
or U50 (N_50,In_4284,In_1097);
xor U51 (N_51,In_4170,In_1513);
or U52 (N_52,In_2242,In_4723);
xnor U53 (N_53,In_3099,In_866);
nand U54 (N_54,In_1387,In_2195);
or U55 (N_55,In_970,In_2778);
nand U56 (N_56,In_2331,In_2664);
and U57 (N_57,In_3390,In_3559);
nor U58 (N_58,In_3693,In_1416);
or U59 (N_59,In_3854,In_3829);
or U60 (N_60,In_655,In_3463);
and U61 (N_61,In_748,In_2262);
nor U62 (N_62,In_4376,In_1787);
xnor U63 (N_63,In_606,In_4205);
and U64 (N_64,In_2610,In_1645);
and U65 (N_65,In_4097,In_2715);
nand U66 (N_66,In_861,In_2511);
nand U67 (N_67,In_1070,In_1160);
nor U68 (N_68,In_4929,In_2852);
nor U69 (N_69,In_448,In_2916);
nand U70 (N_70,In_1355,In_2259);
or U71 (N_71,In_1841,In_2111);
or U72 (N_72,In_4615,In_4704);
nand U73 (N_73,In_3132,In_3300);
and U74 (N_74,In_4296,In_3953);
nor U75 (N_75,In_4952,In_2122);
nor U76 (N_76,In_791,In_2609);
nand U77 (N_77,In_466,In_4880);
or U78 (N_78,In_2194,In_597);
or U79 (N_79,In_4819,In_4549);
xnor U80 (N_80,In_2290,In_2665);
or U81 (N_81,In_35,In_4684);
nor U82 (N_82,In_4933,In_3957);
nor U83 (N_83,In_2491,In_3749);
nand U84 (N_84,In_420,In_2824);
nor U85 (N_85,In_185,In_4456);
and U86 (N_86,In_1898,In_28);
nor U87 (N_87,In_684,In_1571);
nor U88 (N_88,In_2878,In_749);
nor U89 (N_89,In_1220,In_4102);
nand U90 (N_90,In_164,In_4834);
nand U91 (N_91,In_1613,In_3960);
nand U92 (N_92,In_2135,In_1259);
xnor U93 (N_93,In_1235,In_1830);
nand U94 (N_94,In_541,In_4569);
and U95 (N_95,In_3079,In_719);
or U96 (N_96,In_138,In_1066);
and U97 (N_97,In_3653,In_1069);
nor U98 (N_98,In_910,In_3235);
nand U99 (N_99,In_1938,In_3567);
or U100 (N_100,In_1680,In_2938);
nand U101 (N_101,In_1073,In_4911);
xnor U102 (N_102,In_2058,In_3807);
nand U103 (N_103,In_4106,In_191);
and U104 (N_104,In_1793,In_817);
xnor U105 (N_105,In_3504,In_523);
or U106 (N_106,In_682,In_2036);
xnor U107 (N_107,In_1529,In_1615);
nor U108 (N_108,In_4306,In_1247);
and U109 (N_109,In_4414,In_352);
or U110 (N_110,In_3194,In_538);
and U111 (N_111,In_3355,In_3307);
or U112 (N_112,In_2284,In_1662);
and U113 (N_113,In_4075,In_694);
and U114 (N_114,In_605,In_4194);
xor U115 (N_115,In_4460,In_2448);
nand U116 (N_116,In_3705,In_2304);
and U117 (N_117,In_4318,In_683);
nand U118 (N_118,In_2318,In_3124);
xnor U119 (N_119,In_2042,In_4021);
and U120 (N_120,In_1435,In_1059);
and U121 (N_121,In_1765,In_2592);
nand U122 (N_122,In_1398,In_1415);
or U123 (N_123,In_356,In_1391);
and U124 (N_124,In_4491,In_3349);
nor U125 (N_125,In_2109,In_950);
nand U126 (N_126,In_4871,In_4344);
and U127 (N_127,In_4768,In_2282);
or U128 (N_128,In_3088,In_4196);
and U129 (N_129,In_884,In_2067);
or U130 (N_130,In_2309,In_1519);
and U131 (N_131,In_920,In_1277);
nor U132 (N_132,In_2395,In_3110);
nand U133 (N_133,In_4508,In_1324);
or U134 (N_134,In_453,In_1317);
nand U135 (N_135,In_1597,In_4369);
xor U136 (N_136,In_2552,In_2169);
and U137 (N_137,In_2171,In_4585);
xnor U138 (N_138,In_1692,In_4428);
and U139 (N_139,In_1623,In_2877);
xor U140 (N_140,In_668,In_1079);
nand U141 (N_141,In_3399,In_4770);
or U142 (N_142,In_1711,In_92);
and U143 (N_143,In_3579,In_4283);
xnor U144 (N_144,In_3263,In_2057);
xor U145 (N_145,In_3666,In_4693);
xnor U146 (N_146,In_4148,In_399);
xor U147 (N_147,In_3825,In_3987);
or U148 (N_148,In_2206,In_4332);
nor U149 (N_149,In_1983,In_4991);
xnor U150 (N_150,In_2876,In_4985);
and U151 (N_151,In_2208,In_2717);
nand U152 (N_152,In_1768,In_1928);
xnor U153 (N_153,In_3652,In_2120);
nand U154 (N_154,In_4586,In_3994);
or U155 (N_155,In_3419,In_2931);
xor U156 (N_156,In_4294,In_4697);
nand U157 (N_157,In_967,In_1804);
and U158 (N_158,In_4430,In_4004);
and U159 (N_159,In_4316,In_2933);
and U160 (N_160,In_2322,In_2566);
nor U161 (N_161,In_2930,In_2502);
or U162 (N_162,In_4212,In_1353);
or U163 (N_163,In_3348,In_3182);
nor U164 (N_164,In_251,In_37);
nand U165 (N_165,In_3270,In_4796);
nand U166 (N_166,In_1642,In_20);
and U167 (N_167,In_672,In_3415);
or U168 (N_168,In_1427,In_4429);
nand U169 (N_169,In_3345,In_4725);
and U170 (N_170,In_902,In_1944);
xor U171 (N_171,In_981,In_1155);
nor U172 (N_172,In_4099,In_3901);
nor U173 (N_173,In_2755,In_3185);
xor U174 (N_174,In_4341,In_4745);
nand U175 (N_175,In_3128,In_3658);
nand U176 (N_176,In_4994,In_2232);
xor U177 (N_177,In_4084,In_1278);
xor U178 (N_178,In_4143,In_2899);
xnor U179 (N_179,In_3847,In_3288);
nor U180 (N_180,In_1031,In_3269);
or U181 (N_181,In_1693,In_4046);
xor U182 (N_182,In_3860,In_4830);
or U183 (N_183,In_4901,In_4996);
or U184 (N_184,In_789,In_3186);
nor U185 (N_185,In_1028,In_3346);
nor U186 (N_186,In_4250,In_3111);
nand U187 (N_187,In_4217,In_3197);
nand U188 (N_188,In_1889,In_3143);
nor U189 (N_189,In_3622,In_1902);
nor U190 (N_190,In_4310,In_3880);
and U191 (N_191,In_1258,In_4338);
nand U192 (N_192,In_355,In_2073);
and U193 (N_193,In_2779,In_2244);
xor U194 (N_194,In_2917,In_4554);
or U195 (N_195,In_2270,In_26);
xnor U196 (N_196,In_1085,In_972);
or U197 (N_197,In_1647,In_2196);
and U198 (N_198,In_3806,In_4314);
or U199 (N_199,In_1150,In_2412);
xnor U200 (N_200,In_4023,In_864);
xnor U201 (N_201,In_1912,In_3213);
or U202 (N_202,In_562,In_460);
or U203 (N_203,In_1018,In_418);
or U204 (N_204,In_2557,In_3898);
nor U205 (N_205,In_70,In_67);
and U206 (N_206,In_1884,In_2786);
xor U207 (N_207,In_2966,In_2758);
nand U208 (N_208,In_1837,In_3924);
or U209 (N_209,In_3552,In_170);
and U210 (N_210,In_2355,In_3000);
xnor U211 (N_211,In_282,In_3203);
and U212 (N_212,In_3508,In_4577);
xnor U213 (N_213,In_1555,In_3907);
and U214 (N_214,In_245,In_763);
nand U215 (N_215,In_2039,In_3671);
xnor U216 (N_216,In_4187,In_4055);
nand U217 (N_217,In_2103,In_2882);
or U218 (N_218,In_4896,In_2614);
nand U219 (N_219,In_781,In_2080);
xnor U220 (N_220,In_3222,In_1113);
nor U221 (N_221,In_4018,In_1458);
nand U222 (N_222,In_3314,In_897);
or U223 (N_223,In_2836,In_4122);
nand U224 (N_224,In_3464,In_3104);
nand U225 (N_225,In_706,In_1893);
or U226 (N_226,In_1173,In_1817);
nor U227 (N_227,In_2869,In_4476);
nand U228 (N_228,In_3048,In_2847);
nor U229 (N_229,In_2908,In_1466);
or U230 (N_230,In_2469,In_360);
nand U231 (N_231,In_4446,In_1709);
or U232 (N_232,In_2394,In_3835);
nand U233 (N_233,In_4763,In_954);
or U234 (N_234,In_1949,In_2172);
nor U235 (N_235,In_3233,In_1095);
nor U236 (N_236,In_2349,In_3527);
nand U237 (N_237,In_1128,In_2512);
or U238 (N_238,In_2147,In_2524);
nor U239 (N_239,In_4445,In_2804);
xor U240 (N_240,In_34,In_3695);
nand U241 (N_241,In_3159,In_1646);
nor U242 (N_242,In_4164,In_4119);
and U243 (N_243,In_2799,In_3020);
xnor U244 (N_244,In_3443,In_1335);
xnor U245 (N_245,In_731,In_792);
nor U246 (N_246,In_582,In_3561);
or U247 (N_247,In_4596,In_3261);
or U248 (N_248,In_1992,In_4583);
nor U249 (N_249,In_4346,In_753);
nor U250 (N_250,In_2853,In_4881);
xnor U251 (N_251,In_1120,In_1661);
xor U252 (N_252,In_1565,In_4126);
nand U253 (N_253,In_4765,In_3905);
and U254 (N_254,In_2672,In_4893);
nand U255 (N_255,In_1005,In_560);
or U256 (N_256,In_2104,In_4947);
or U257 (N_257,In_1965,In_256);
xnor U258 (N_258,In_3726,In_4696);
and U259 (N_259,In_3207,In_528);
nand U260 (N_260,In_4755,In_3512);
and U261 (N_261,In_1552,In_2163);
xor U262 (N_262,In_3677,In_2955);
nor U263 (N_263,In_81,In_2994);
nand U264 (N_264,In_4022,In_2288);
xnor U265 (N_265,In_769,In_105);
xnor U266 (N_266,In_1907,In_490);
nor U267 (N_267,In_4829,In_760);
xnor U268 (N_268,In_4859,In_72);
or U269 (N_269,In_3578,In_3290);
nand U270 (N_270,In_501,In_3796);
nand U271 (N_271,In_4516,In_627);
nand U272 (N_272,In_4210,In_1051);
or U273 (N_273,In_3748,In_2019);
and U274 (N_274,In_4091,In_4375);
and U275 (N_275,In_3500,In_1913);
nor U276 (N_276,In_389,In_2500);
and U277 (N_277,In_422,In_3335);
xor U278 (N_278,In_1503,In_2953);
xnor U279 (N_279,In_3574,In_4120);
nand U280 (N_280,In_610,In_3189);
and U281 (N_281,In_2637,In_3838);
xor U282 (N_282,In_3721,In_3712);
or U283 (N_283,In_3416,In_2054);
or U284 (N_284,In_2276,In_2508);
or U285 (N_285,In_3632,In_31);
nor U286 (N_286,In_4070,In_4690);
nor U287 (N_287,In_90,In_3708);
or U288 (N_288,In_3562,In_236);
or U289 (N_289,In_18,In_2981);
nand U290 (N_290,In_533,In_4812);
or U291 (N_291,In_1242,In_3776);
xor U292 (N_292,In_386,In_1759);
or U293 (N_293,In_2956,In_4035);
xnor U294 (N_294,In_612,In_2835);
xnor U295 (N_295,In_4427,In_1358);
or U296 (N_296,In_1506,In_2445);
nand U297 (N_297,In_2993,In_730);
nor U298 (N_298,In_205,In_4221);
xor U299 (N_299,In_203,In_4042);
or U300 (N_300,In_4008,In_359);
or U301 (N_301,In_2001,In_4032);
xnor U302 (N_302,In_1831,In_845);
and U303 (N_303,In_140,In_306);
or U304 (N_304,In_2510,In_3981);
or U305 (N_305,In_805,In_1791);
nand U306 (N_306,In_4398,In_860);
nand U307 (N_307,In_3435,In_2941);
and U308 (N_308,In_3947,In_3147);
nand U309 (N_309,In_461,In_3809);
or U310 (N_310,In_1050,In_145);
nand U311 (N_311,In_3858,In_638);
or U312 (N_312,In_39,In_268);
and U313 (N_313,In_557,In_3986);
xnor U314 (N_314,In_3551,In_1764);
nand U315 (N_315,In_3886,In_2404);
xor U316 (N_316,In_4232,In_3141);
and U317 (N_317,In_894,In_291);
nor U318 (N_318,In_2181,In_1723);
xnor U319 (N_319,In_4926,In_4739);
nor U320 (N_320,In_1780,In_1578);
and U321 (N_321,In_955,In_1846);
nor U322 (N_322,In_292,In_4636);
and U323 (N_323,In_4865,In_1257);
and U324 (N_324,In_463,In_1172);
and U325 (N_325,In_1592,In_1682);
xor U326 (N_326,In_4879,In_2704);
nor U327 (N_327,In_576,In_3083);
or U328 (N_328,In_1722,In_3801);
xor U329 (N_329,In_1036,In_2924);
nor U330 (N_330,In_3526,In_3585);
and U331 (N_331,In_4658,In_3889);
nand U332 (N_332,In_4754,In_3340);
or U333 (N_333,In_870,In_1761);
nor U334 (N_334,In_1741,In_2185);
nand U335 (N_335,In_3215,In_2198);
or U336 (N_336,In_1266,In_2892);
nor U337 (N_337,In_1991,In_1164);
nor U338 (N_338,In_2601,In_1784);
nor U339 (N_339,In_3816,In_4289);
xor U340 (N_340,In_1946,In_1074);
xnor U341 (N_341,In_2652,In_3379);
nand U342 (N_342,In_1744,In_568);
xor U343 (N_343,In_928,In_1593);
nand U344 (N_344,In_4117,In_669);
and U345 (N_345,In_658,In_4822);
and U346 (N_346,In_4737,In_4335);
and U347 (N_347,In_3172,In_4707);
and U348 (N_348,In_519,In_1012);
or U349 (N_349,In_1269,In_2929);
nor U350 (N_350,In_656,In_4965);
nor U351 (N_351,In_2587,In_3092);
or U352 (N_352,In_226,In_1419);
and U353 (N_353,In_896,In_3109);
xnor U354 (N_354,In_3402,In_2435);
and U355 (N_355,In_1751,In_2602);
nor U356 (N_356,In_1168,In_235);
or U357 (N_357,In_2119,In_1094);
and U358 (N_358,In_4849,In_3962);
and U359 (N_359,In_1632,In_4744);
nand U360 (N_360,In_720,In_4719);
or U361 (N_361,In_3645,In_4802);
xor U362 (N_362,In_3298,In_1034);
nand U363 (N_363,In_521,In_1481);
or U364 (N_364,In_414,In_4557);
and U365 (N_365,In_3452,In_1332);
and U366 (N_366,In_3573,In_1049);
nand U367 (N_367,In_2999,In_1796);
nor U368 (N_368,In_2798,In_4756);
or U369 (N_369,In_4786,In_3468);
and U370 (N_370,In_3667,In_951);
xor U371 (N_371,In_3429,In_62);
nor U372 (N_372,In_278,In_471);
nand U373 (N_373,In_2562,In_1381);
and U374 (N_374,In_4823,In_3700);
xnor U375 (N_375,In_1700,In_696);
xor U376 (N_376,In_2371,In_3306);
nand U377 (N_377,In_108,In_4342);
nor U378 (N_378,In_4072,In_212);
nand U379 (N_379,In_3584,In_4534);
or U380 (N_380,In_3055,In_439);
xor U381 (N_381,In_3267,In_3187);
xnor U382 (N_382,In_4689,In_1039);
or U383 (N_383,In_1076,In_1895);
nand U384 (N_384,In_797,In_2539);
nand U385 (N_385,In_4125,In_4563);
and U386 (N_386,In_1188,In_2784);
xor U387 (N_387,In_623,In_2731);
or U388 (N_388,In_1286,In_2176);
nand U389 (N_389,In_2806,In_1507);
or U390 (N_390,In_3763,In_4374);
xnor U391 (N_391,In_1828,In_1017);
and U392 (N_392,In_3012,In_2537);
nor U393 (N_393,In_1718,In_1921);
nor U394 (N_394,In_36,In_755);
nand U395 (N_395,In_2811,In_1403);
or U396 (N_396,In_1640,In_2772);
nand U397 (N_397,In_3711,In_2497);
nand U398 (N_398,In_2534,In_1870);
nor U399 (N_399,In_3511,In_2273);
nor U400 (N_400,In_1591,In_2366);
and U401 (N_401,In_1222,In_4886);
and U402 (N_402,In_11,In_2974);
or U403 (N_403,In_3190,In_2378);
and U404 (N_404,In_2760,In_4477);
xnor U405 (N_405,In_3470,In_4144);
nor U406 (N_406,In_2662,In_1282);
xnor U407 (N_407,In_3210,In_4784);
nor U408 (N_408,In_2724,In_3674);
xnor U409 (N_409,In_4954,In_1575);
xor U410 (N_410,In_4264,In_2516);
or U411 (N_411,In_1371,In_4505);
or U412 (N_412,In_3474,In_590);
xor U413 (N_413,In_980,In_770);
or U414 (N_414,In_3204,In_1467);
nand U415 (N_415,In_3246,In_4809);
and U416 (N_416,In_3952,In_1892);
nor U417 (N_417,In_1852,In_553);
and U418 (N_418,In_4415,In_1924);
nand U419 (N_419,In_2671,In_2248);
or U420 (N_420,In_2018,In_1900);
nand U421 (N_421,In_487,In_2630);
nor U422 (N_422,In_4349,In_4942);
nor U423 (N_423,In_1140,In_738);
xor U424 (N_424,In_3804,In_1411);
nand U425 (N_425,In_4280,In_953);
nand U426 (N_426,In_2160,In_1811);
nor U427 (N_427,In_4957,In_299);
nand U428 (N_428,In_847,In_3506);
and U429 (N_429,In_221,In_509);
or U430 (N_430,In_1544,In_1600);
xor U431 (N_431,In_419,In_4927);
nand U432 (N_432,In_2984,In_3687);
or U433 (N_433,In_2440,In_2749);
and U434 (N_434,In_3027,In_611);
xor U435 (N_435,In_428,In_2686);
and U436 (N_436,In_2962,In_2744);
xor U437 (N_437,In_4172,In_4788);
or U438 (N_438,In_3615,In_3681);
nand U439 (N_439,In_252,In_741);
nor U440 (N_440,In_341,In_1872);
nand U441 (N_441,In_2850,In_1724);
or U442 (N_442,In_165,In_3098);
or U443 (N_443,In_2972,In_2659);
nor U444 (N_444,In_2029,In_1522);
or U445 (N_445,In_3780,In_1747);
nor U446 (N_446,In_587,In_3094);
xnor U447 (N_447,In_784,In_670);
and U448 (N_448,In_2090,In_3575);
or U449 (N_449,In_2875,In_2789);
nand U450 (N_450,In_503,In_549);
nand U451 (N_451,In_3179,In_4902);
nor U452 (N_452,In_2961,In_3397);
nand U453 (N_453,In_3163,In_187);
and U454 (N_454,In_4895,In_2775);
nor U455 (N_455,In_3741,In_1654);
nor U456 (N_456,In_4160,In_2912);
or U457 (N_457,In_2757,In_2900);
and U458 (N_458,In_3129,In_4391);
xor U459 (N_459,In_4108,In_4635);
or U460 (N_460,In_2204,In_1096);
or U461 (N_461,In_957,In_2024);
nand U462 (N_462,In_1136,In_2433);
xnor U463 (N_463,In_3643,In_3557);
xnor U464 (N_464,In_288,In_1910);
nor U465 (N_465,In_4846,In_3155);
and U466 (N_466,In_313,In_1885);
and U467 (N_467,In_2990,In_2560);
and U468 (N_468,In_1997,In_4095);
nand U469 (N_469,In_3078,In_4597);
and U470 (N_470,In_2680,In_134);
xor U471 (N_471,In_3217,In_1084);
nor U472 (N_472,In_827,In_883);
xnor U473 (N_473,In_2365,In_3059);
nor U474 (N_474,In_4654,In_3154);
nor U475 (N_475,In_2517,In_558);
or U476 (N_476,In_1275,In_3972);
and U477 (N_477,In_2780,In_1489);
xor U478 (N_478,In_4783,In_4634);
and U479 (N_479,In_302,In_4225);
nor U480 (N_480,In_410,In_1926);
and U481 (N_481,In_2110,In_952);
and U482 (N_482,In_1117,In_449);
xor U483 (N_483,In_4141,In_4197);
or U484 (N_484,In_3606,In_3438);
xnor U485 (N_485,In_956,In_4490);
or U486 (N_486,In_2342,In_2154);
xor U487 (N_487,In_1664,In_3792);
and U488 (N_488,In_1213,In_1303);
or U489 (N_489,In_4452,In_2808);
xnor U490 (N_490,In_3382,In_869);
nand U491 (N_491,In_1206,In_842);
xor U492 (N_492,In_2092,In_4357);
and U493 (N_493,In_2921,In_1280);
xor U494 (N_494,In_4053,In_1650);
nand U495 (N_495,In_2466,In_492);
or U496 (N_496,In_859,In_290);
nand U497 (N_497,In_2957,In_2874);
nor U498 (N_498,In_4595,In_1483);
or U499 (N_499,In_630,In_4740);
nand U500 (N_500,In_1875,In_392);
nand U501 (N_501,In_3710,In_765);
or U502 (N_502,In_795,In_3149);
nand U503 (N_503,In_445,In_697);
and U504 (N_504,In_4525,In_385);
nor U505 (N_505,In_3973,In_156);
nand U506 (N_506,In_4,In_402);
and U507 (N_507,In_2859,In_2487);
xnor U508 (N_508,In_485,In_4526);
and U509 (N_509,In_3242,In_2829);
xor U510 (N_510,In_1495,In_530);
xor U511 (N_511,In_1116,In_559);
xor U512 (N_512,In_1347,In_403);
nor U513 (N_513,In_580,In_3845);
xor U514 (N_514,In_371,In_575);
or U515 (N_515,In_493,In_1832);
or U516 (N_516,In_1879,In_4631);
nor U517 (N_517,In_4074,In_3505);
nor U518 (N_518,In_2881,In_878);
or U519 (N_519,In_284,In_150);
nor U520 (N_520,In_275,In_2509);
xor U521 (N_521,In_318,In_3798);
or U522 (N_522,In_2234,In_3948);
nand U523 (N_523,In_2589,In_4797);
nand U524 (N_524,In_4265,In_3752);
and U525 (N_525,In_916,In_2620);
or U526 (N_526,In_939,In_3214);
xnor U527 (N_527,In_4492,In_4111);
or U528 (N_528,In_2475,In_1834);
or U529 (N_529,In_4803,In_2422);
or U530 (N_530,In_4839,In_4598);
and U531 (N_531,In_3238,In_4573);
xnor U532 (N_532,In_243,In_1134);
nor U533 (N_533,In_1102,In_622);
or U534 (N_534,In_1839,In_634);
nand U535 (N_535,In_4591,In_429);
or U536 (N_536,In_1093,In_908);
xnor U537 (N_537,In_2237,In_227);
and U538 (N_538,In_1713,In_2649);
and U539 (N_539,In_2866,In_4662);
or U540 (N_540,In_2828,In_2893);
nor U541 (N_541,In_4025,In_3691);
nor U542 (N_542,In_2987,In_848);
nor U543 (N_543,In_4890,In_1224);
or U544 (N_544,In_396,In_4457);
xor U545 (N_545,In_3802,In_384);
nor U546 (N_546,In_2161,In_478);
and U547 (N_547,In_2666,In_3004);
nand U548 (N_548,In_2040,In_4641);
nor U549 (N_549,In_3684,In_4567);
nand U550 (N_550,In_3177,In_4527);
nor U551 (N_551,In_931,In_2207);
nand U552 (N_552,In_2805,In_2896);
nand U553 (N_553,In_2920,In_3656);
and U554 (N_554,In_937,In_2880);
nand U555 (N_555,In_3469,In_1183);
nor U556 (N_556,In_1379,In_4067);
and U557 (N_557,In_4007,In_3015);
or U558 (N_558,In_2505,In_3625);
nor U559 (N_559,In_4547,In_2411);
xor U560 (N_560,In_4961,In_3844);
or U561 (N_561,In_4995,In_716);
nor U562 (N_562,In_3761,In_4971);
nor U563 (N_563,In_3380,In_551);
or U564 (N_564,In_4633,In_4162);
or U565 (N_565,In_1402,In_189);
nand U566 (N_566,In_4211,In_4293);
and U567 (N_567,In_2464,In_3910);
or U568 (N_568,In_4899,In_1769);
nor U569 (N_569,In_2703,In_3897);
or U570 (N_570,In_3929,In_2354);
or U571 (N_571,In_4909,In_131);
nor U572 (N_572,In_527,In_19);
or U573 (N_573,In_4069,In_4485);
or U574 (N_574,In_1365,In_628);
nor U575 (N_575,In_4279,In_442);
nand U576 (N_576,In_4531,In_4907);
xor U577 (N_577,In_707,In_4750);
nor U578 (N_578,In_3302,In_3673);
or U579 (N_579,In_1145,In_3689);
nor U580 (N_580,In_477,In_2060);
nor U581 (N_581,In_4945,In_4079);
nand U582 (N_582,In_2837,In_564);
and U583 (N_583,In_3513,In_3425);
or U584 (N_584,In_374,In_890);
and U585 (N_585,In_4045,In_3198);
or U586 (N_586,In_2542,In_1690);
and U587 (N_587,In_2545,In_3982);
or U588 (N_588,In_88,In_2240);
and U589 (N_589,In_3707,In_473);
nor U590 (N_590,In_2532,In_229);
nand U591 (N_591,In_3030,In_1757);
nor U592 (N_592,In_4436,In_2834);
or U593 (N_593,In_2886,In_1630);
or U594 (N_594,In_1810,In_2613);
xnor U595 (N_595,In_3842,In_3950);
nand U596 (N_596,In_1166,In_3264);
nand U597 (N_597,In_280,In_3192);
or U598 (N_598,In_3954,In_3590);
and U599 (N_599,In_2567,In_2948);
nor U600 (N_600,In_1955,In_1378);
nand U601 (N_601,In_1638,In_3258);
and U602 (N_602,In_3492,In_4440);
or U603 (N_603,In_2481,In_2434);
xor U604 (N_604,In_1037,In_4278);
xor U605 (N_605,In_3401,In_821);
and U606 (N_606,In_4556,In_66);
or U607 (N_607,In_2173,In_3205);
xor U608 (N_608,In_2007,In_1651);
nand U609 (N_609,In_2151,In_3138);
nor U610 (N_610,In_2314,In_2627);
nand U611 (N_611,In_3945,In_1903);
and U612 (N_612,In_4983,In_1433);
nand U613 (N_613,In_4568,In_2551);
and U614 (N_614,In_3356,In_616);
xnor U615 (N_615,In_660,In_544);
nor U616 (N_616,In_1734,In_1437);
nand U617 (N_617,In_688,In_534);
xnor U618 (N_618,In_1459,In_76);
nor U619 (N_619,In_3158,In_1216);
or U620 (N_620,In_1288,In_416);
xor U621 (N_621,In_4326,In_4666);
nor U622 (N_622,In_1157,In_3032);
xor U623 (N_623,In_3593,In_4671);
and U624 (N_624,In_3661,In_2651);
or U625 (N_625,In_1801,In_846);
or U626 (N_626,In_2306,In_3529);
nand U627 (N_627,In_4432,In_3161);
and U628 (N_628,In_238,In_1314);
and U629 (N_629,In_1687,In_4758);
nand U630 (N_630,In_1492,In_3255);
xor U631 (N_631,In_2611,In_193);
nor U632 (N_632,In_3805,In_1141);
xor U633 (N_633,In_162,In_4820);
and U634 (N_634,In_1197,In_1816);
nand U635 (N_635,In_2606,In_787);
or U636 (N_636,In_3344,In_132);
nand U637 (N_637,In_68,In_2714);
nor U638 (N_638,In_537,In_2531);
or U639 (N_639,In_1,In_3028);
and U640 (N_640,In_824,In_2139);
xor U641 (N_641,In_3540,In_914);
or U642 (N_642,In_2530,In_4800);
nor U643 (N_643,In_3934,In_3280);
xnor U644 (N_644,In_2568,In_4129);
and U645 (N_645,In_3496,In_161);
nand U646 (N_646,In_4274,In_3966);
and U647 (N_647,In_3130,In_515);
nand U648 (N_648,In_714,In_3913);
xnor U649 (N_649,In_4914,In_4582);
nor U650 (N_650,In_1629,In_3228);
or U651 (N_651,In_1812,In_3760);
and U652 (N_652,In_269,In_3826);
xor U653 (N_653,In_3704,In_1573);
nand U654 (N_654,In_4098,In_3808);
nor U655 (N_655,In_4152,In_2344);
xnor U656 (N_656,In_3122,In_1679);
and U657 (N_657,In_1950,In_4151);
nor U658 (N_658,In_1289,In_4333);
and U659 (N_659,In_903,In_2155);
nor U660 (N_660,In_3025,In_4845);
nand U661 (N_661,In_918,In_4168);
or U662 (N_662,In_1177,In_2050);
xnor U663 (N_663,In_502,In_960);
nor U664 (N_664,In_764,In_4254);
xor U665 (N_665,In_4702,In_3361);
xor U666 (N_666,In_3084,In_3308);
or U667 (N_667,In_904,In_2529);
or U668 (N_668,In_1790,In_4063);
xnor U669 (N_669,In_2116,In_4300);
xor U670 (N_670,In_1425,In_2231);
xnor U671 (N_671,In_3788,In_1129);
nor U672 (N_672,In_3911,In_3767);
xnor U673 (N_673,In_3627,In_4267);
nor U674 (N_674,In_286,In_4115);
xor U675 (N_675,In_309,In_2034);
xnor U676 (N_676,In_3619,In_906);
xnor U677 (N_677,In_2549,In_4566);
or U678 (N_678,In_667,In_1673);
and U679 (N_679,In_1504,In_214);
xnor U680 (N_680,In_1773,In_4155);
and U681 (N_681,In_2197,In_4715);
xor U682 (N_682,In_3417,In_474);
nand U683 (N_683,In_4883,In_4963);
or U684 (N_684,In_77,In_3915);
or U685 (N_685,In_512,In_3811);
nor U686 (N_686,In_2547,In_3904);
and U687 (N_687,In_2410,In_3961);
nor U688 (N_688,In_3148,In_218);
or U689 (N_689,In_2889,In_32);
or U690 (N_690,In_4334,In_2949);
nor U691 (N_691,In_736,In_888);
or U692 (N_692,In_387,In_3594);
or U693 (N_693,In_3520,In_4459);
nor U694 (N_694,In_2037,In_4271);
or U695 (N_695,In_2011,In_2741);
or U696 (N_696,In_3362,In_3353);
and U697 (N_697,In_1753,In_1126);
or U698 (N_698,In_2450,In_2209);
or U699 (N_699,In_1236,In_2328);
nand U700 (N_700,In_3067,In_806);
xor U701 (N_701,In_1055,In_1523);
nand U702 (N_702,In_3317,In_4928);
nand U703 (N_703,In_421,In_4124);
nor U704 (N_704,In_3370,In_3279);
xnor U705 (N_705,In_520,In_2483);
nor U706 (N_706,In_271,In_44);
and U707 (N_707,In_1917,In_3550);
or U708 (N_708,In_86,In_2321);
xnor U709 (N_709,In_3329,In_1344);
and U710 (N_710,In_2088,In_3662);
or U711 (N_711,In_517,In_3241);
or U712 (N_712,In_932,In_3586);
nor U713 (N_713,In_1710,In_4672);
xor U714 (N_714,In_1244,In_4686);
or U715 (N_715,In_2260,In_4711);
nor U716 (N_716,In_1449,In_4365);
nor U717 (N_717,In_1271,In_2363);
and U718 (N_718,In_1535,In_3794);
or U719 (N_719,In_4331,In_912);
nor U720 (N_720,In_1302,In_2636);
or U721 (N_721,In_815,In_469);
xnor U722 (N_722,In_4564,In_1214);
nand U723 (N_723,In_369,In_3497);
nor U724 (N_724,In_2752,In_1189);
xnor U725 (N_725,In_577,In_2635);
nand U726 (N_726,In_2527,In_4565);
nand U727 (N_727,In_3284,In_2420);
and U728 (N_728,In_516,In_267);
and U729 (N_729,In_2105,In_3983);
xnor U730 (N_730,In_3388,In_740);
xnor U731 (N_731,In_3038,In_4924);
nor U732 (N_732,In_2312,In_1840);
and U733 (N_733,In_3820,In_617);
nor U734 (N_734,In_4135,In_1699);
nor U735 (N_735,In_4033,In_4777);
nand U736 (N_736,In_2661,In_4000);
xor U737 (N_737,In_2238,In_2826);
xor U738 (N_738,In_2657,In_1968);
or U739 (N_739,In_4680,In_4343);
and U740 (N_740,In_4051,In_3107);
or U741 (N_741,In_836,In_2584);
and U742 (N_742,In_1845,In_4691);
nand U743 (N_743,In_2967,In_2159);
xnor U744 (N_744,In_4204,In_963);
and U745 (N_745,In_1428,In_979);
nor U746 (N_746,In_532,In_186);
nand U747 (N_747,In_2436,In_4512);
or U748 (N_748,In_1669,In_607);
or U749 (N_749,In_3278,In_4513);
xor U750 (N_750,In_1041,In_3781);
nor U751 (N_751,In_3998,In_3657);
or U752 (N_752,In_4638,In_1372);
nor U753 (N_753,In_996,In_813);
nand U754 (N_754,In_1694,In_3990);
nand U755 (N_755,In_4260,In_2723);
or U756 (N_756,In_1981,In_1374);
xor U757 (N_757,In_4856,In_3180);
xnor U758 (N_758,In_771,In_1100);
xnor U759 (N_759,In_2867,In_983);
xnor U760 (N_760,In_892,In_2272);
nor U761 (N_761,In_4869,In_270);
nand U762 (N_762,In_63,In_871);
or U763 (N_763,In_4767,In_3162);
or U764 (N_764,In_2452,In_4515);
or U765 (N_765,In_3456,In_2573);
xnor U766 (N_766,In_1730,In_4397);
nor U767 (N_767,In_1715,In_4530);
nand U768 (N_768,In_3928,In_3243);
xor U769 (N_769,In_2214,In_3955);
xor U770 (N_770,In_1445,In_2323);
or U771 (N_771,In_799,In_4005);
and U772 (N_772,In_2998,In_244);
nand U773 (N_773,In_2117,In_4769);
nand U774 (N_774,In_366,In_1016);
xnor U775 (N_775,In_3085,In_1331);
xor U776 (N_776,In_3126,In_2683);
xor U777 (N_777,In_1375,In_4936);
and U778 (N_778,In_3378,In_1338);
nor U779 (N_779,In_4872,In_1482);
nand U780 (N_780,In_1937,In_98);
or U781 (N_781,In_4694,In_938);
xnor U782 (N_782,In_2146,In_1726);
xnor U783 (N_783,In_2470,In_12);
nor U784 (N_784,In_2447,In_793);
and U785 (N_785,In_4855,In_536);
and U786 (N_786,In_3864,In_3439);
xnor U787 (N_787,In_4675,In_768);
xor U788 (N_788,In_2794,In_4701);
nor U789 (N_789,In_2091,In_2303);
and U790 (N_790,In_3978,In_196);
xor U791 (N_791,In_4898,In_4612);
or U792 (N_792,In_4507,In_2935);
and U793 (N_793,In_653,In_4986);
nor U794 (N_794,In_3226,In_4760);
nor U795 (N_795,In_2415,In_3856);
xnor U796 (N_796,In_2203,In_315);
or U797 (N_797,In_1549,In_1742);
nand U798 (N_798,In_3450,In_1583);
nand U799 (N_799,In_1854,In_2414);
or U800 (N_800,In_4503,In_3001);
and U801 (N_801,In_4623,In_4759);
xor U802 (N_802,In_2125,In_4682);
xor U803 (N_803,In_1754,In_2078);
nor U804 (N_804,In_1478,In_3927);
and U805 (N_805,In_3,In_3894);
and U806 (N_806,In_3799,In_2764);
and U807 (N_807,In_1634,In_1191);
or U808 (N_808,In_4989,In_1982);
and U809 (N_809,In_3688,In_2417);
nor U810 (N_810,In_2390,In_840);
nor U811 (N_811,In_4736,In_58);
or U812 (N_812,In_3714,In_3610);
nand U813 (N_813,In_2076,In_2175);
or U814 (N_814,In_3582,In_2021);
nand U815 (N_815,In_4404,In_1024);
or U816 (N_816,In_1505,In_1139);
or U817 (N_817,In_4313,In_2766);
nor U818 (N_818,In_2771,In_3640);
or U819 (N_819,In_1211,In_3676);
nor U820 (N_820,In_973,In_2586);
xnor U821 (N_821,In_2519,In_169);
nand U822 (N_822,In_880,In_4572);
or U823 (N_823,In_3524,In_4030);
nand U824 (N_824,In_388,In_3768);
nand U825 (N_825,In_488,In_1948);
or U826 (N_826,In_1038,In_3735);
nand U827 (N_827,In_2245,In_60);
xor U828 (N_828,In_820,In_2484);
and U829 (N_829,In_3117,In_750);
and U830 (N_830,In_4257,In_1617);
and U831 (N_831,In_3589,In_4191);
nor U832 (N_832,In_2849,In_807);
or U833 (N_833,In_143,In_2376);
or U834 (N_834,In_1023,In_3765);
xnor U835 (N_835,In_4817,In_2184);
nand U836 (N_836,In_217,In_739);
nand U837 (N_837,In_2168,In_3785);
and U838 (N_838,In_879,In_637);
xnor U839 (N_839,In_1514,In_2157);
nand U840 (N_840,In_231,In_3738);
and U841 (N_841,In_1720,In_3895);
or U842 (N_842,In_2643,In_1137);
nor U843 (N_843,In_3626,In_4486);
nor U844 (N_844,In_2398,In_2301);
nor U845 (N_845,In_1748,In_1287);
nor U846 (N_846,In_1400,In_2668);
or U847 (N_847,In_2945,In_2918);
xnor U848 (N_848,In_3414,In_4661);
and U849 (N_849,In_1359,In_2988);
nor U850 (N_850,In_3404,In_2358);
nand U851 (N_851,In_565,In_4831);
or U852 (N_852,In_2253,In_3216);
nand U853 (N_853,In_4203,In_4287);
and U854 (N_854,In_276,In_3102);
nand U855 (N_855,In_907,In_4522);
nor U856 (N_856,In_1326,In_3156);
nor U857 (N_857,In_228,In_620);
xnor U858 (N_858,In_2619,In_1829);
nor U859 (N_859,In_1301,In_3153);
nor U860 (N_860,In_33,In_2631);
or U861 (N_861,In_4149,In_4145);
or U862 (N_862,In_3305,In_4717);
or U863 (N_863,In_2191,In_1382);
and U864 (N_864,In_3613,In_4977);
and U865 (N_865,In_4288,In_1688);
nand U866 (N_866,In_1473,In_3719);
xor U867 (N_867,In_320,In_3997);
nor U868 (N_868,In_1994,In_2641);
nor U869 (N_869,In_2293,In_1620);
or U870 (N_870,In_3750,In_1062);
nand U871 (N_871,In_2359,In_3906);
xnor U872 (N_872,In_3769,In_2138);
or U873 (N_873,In_2149,In_3672);
or U874 (N_874,In_182,In_1484);
and U875 (N_875,In_4622,In_895);
and U876 (N_876,In_3432,In_1605);
or U877 (N_877,In_2241,In_4487);
or U878 (N_878,In_1684,In_298);
or U879 (N_879,In_2997,In_2158);
and U880 (N_880,In_1826,In_1299);
and U881 (N_881,In_3993,In_3350);
and U882 (N_882,In_1607,In_74);
xor U883 (N_883,In_2838,In_1265);
or U884 (N_884,In_3131,In_4273);
xnor U885 (N_885,In_4495,In_596);
and U886 (N_886,In_722,In_427);
nand U887 (N_887,In_4499,In_2170);
nand U888 (N_888,In_3598,In_2426);
or U889 (N_889,In_437,In_2577);
nand U890 (N_890,In_4482,In_1476);
nor U891 (N_891,In_4798,In_1046);
nor U892 (N_892,In_2737,In_96);
or U893 (N_893,In_1930,In_393);
or U894 (N_894,In_1705,In_2051);
and U895 (N_895,In_1383,In_3006);
xor U896 (N_896,In_1132,In_4474);
or U897 (N_897,In_4781,In_3387);
nand U898 (N_898,In_1906,In_2843);
xnor U899 (N_899,In_881,In_555);
nor U900 (N_900,In_55,In_4669);
and U901 (N_901,In_451,In_2970);
nor U902 (N_902,In_3090,In_4811);
xor U903 (N_903,In_1625,In_2901);
nand U904 (N_904,In_1368,In_1670);
xnor U905 (N_905,In_332,In_1827);
xor U906 (N_906,In_3709,In_2885);
nand U907 (N_907,In_433,In_61);
nand U908 (N_908,In_4101,In_710);
nor U909 (N_909,In_4253,In_4105);
xnor U910 (N_910,In_3281,In_2368);
nand U911 (N_911,In_3428,In_4234);
and U912 (N_912,In_2427,In_2280);
nor U913 (N_913,In_3146,In_4003);
nor U914 (N_914,In_3940,In_223);
or U915 (N_915,In_113,In_1963);
or U916 (N_916,In_1609,In_80);
xor U917 (N_917,In_4175,In_1611);
xor U918 (N_918,In_4442,In_3398);
nand U919 (N_919,In_595,In_4877);
xnor U920 (N_920,In_136,In_930);
xnor U921 (N_921,In_614,In_4843);
nand U922 (N_922,In_3465,In_1252);
xnor U923 (N_923,In_921,In_1360);
or U924 (N_924,In_1914,In_197);
nand U925 (N_925,In_2563,In_3166);
xnor U926 (N_926,In_2707,In_2521);
and U927 (N_927,In_1561,In_1614);
and U928 (N_928,In_927,In_2969);
nand U929 (N_929,In_408,In_4870);
and U930 (N_930,In_4068,In_2725);
and U931 (N_931,In_4560,In_4728);
and U932 (N_932,In_4814,In_2095);
xnor U933 (N_933,In_1940,In_1871);
xor U934 (N_934,In_2989,In_3373);
xor U935 (N_935,In_602,In_915);
nor U936 (N_936,In_2727,In_4384);
xnor U937 (N_937,In_1295,In_3074);
nor U938 (N_938,In_644,In_3989);
or U939 (N_939,In_2106,In_2670);
or U940 (N_940,In_1758,In_3566);
or U941 (N_941,In_417,In_1752);
or U942 (N_942,In_258,In_1138);
nand U943 (N_943,In_2658,In_3392);
nand U944 (N_944,In_188,In_2596);
or U945 (N_945,In_3276,In_1836);
nand U946 (N_946,In_4347,In_2554);
nor U947 (N_947,In_4382,In_2431);
and U948 (N_948,In_599,In_3389);
or U949 (N_949,In_4087,In_1525);
xnor U950 (N_950,In_1007,In_934);
nand U951 (N_951,In_365,In_3611);
and U952 (N_952,In_1104,In_2082);
nor U953 (N_953,In_2851,In_2059);
and U954 (N_954,In_654,In_4588);
nand U955 (N_955,In_2144,In_3871);
and U956 (N_956,In_69,In_3791);
xor U957 (N_957,In_3023,In_16);
and U958 (N_958,In_3171,In_2216);
xor U959 (N_959,In_4721,In_3617);
and U960 (N_960,In_2468,In_4052);
xnor U961 (N_961,In_3930,In_3501);
and U962 (N_962,In_3777,In_3837);
xnor U963 (N_963,In_4953,In_4208);
and U964 (N_964,In_2129,In_3959);
or U965 (N_965,In_1749,In_3070);
and U966 (N_966,In_2819,In_3165);
or U967 (N_967,In_102,In_1200);
xnor U968 (N_968,In_625,In_2380);
nand U969 (N_969,In_4127,In_4174);
nor U970 (N_970,In_1953,In_3437);
xnor U971 (N_971,In_2733,In_380);
or U972 (N_972,In_3056,In_3925);
xor U973 (N_973,In_4408,In_1413);
and U974 (N_974,In_3274,In_1735);
and U975 (N_975,In_2709,In_693);
nor U976 (N_976,In_2030,In_1805);
and U977 (N_977,In_2022,In_2773);
xnor U978 (N_978,In_3876,In_3026);
xnor U979 (N_979,In_594,In_822);
xor U980 (N_980,In_261,In_3853);
nand U981 (N_981,In_1407,In_3252);
and U982 (N_982,In_2408,In_1212);
and U983 (N_983,In_1219,In_4041);
xnor U984 (N_984,In_4908,In_3720);
nor U985 (N_985,In_1978,In_2887);
or U986 (N_986,In_4107,In_4532);
nand U987 (N_987,In_4010,In_689);
nand U988 (N_988,In_2550,In_2165);
nand U989 (N_989,In_4673,In_675);
nor U990 (N_990,In_462,In_1847);
and U991 (N_991,In_123,In_4233);
or U992 (N_992,In_2490,In_4602);
xor U993 (N_993,In_4131,In_1541);
xnor U994 (N_994,In_1672,In_2821);
nand U995 (N_995,In_2113,In_2311);
nand U996 (N_996,In_4766,In_0);
nor U997 (N_997,In_1520,In_4688);
or U998 (N_998,In_2372,In_4077);
nor U999 (N_999,In_1436,In_1357);
nand U1000 (N_1000,In_1652,In_1621);
nor U1001 (N_1001,In_1112,In_4708);
nand U1002 (N_1002,In_2308,In_4443);
nand U1003 (N_1003,In_851,In_4461);
and U1004 (N_1004,In_89,In_1232);
xor U1005 (N_1005,In_3827,In_4301);
nand U1006 (N_1006,In_4975,In_2716);
or U1007 (N_1007,In_2236,In_4972);
xor U1008 (N_1008,In_4860,In_2279);
or U1009 (N_1009,In_2246,In_190);
nor U1010 (N_1010,In_3762,In_3532);
nand U1011 (N_1011,In_598,In_4537);
and U1012 (N_1012,In_2538,In_4874);
nor U1013 (N_1013,In_3412,In_3113);
and U1014 (N_1014,In_3440,In_3531);
xor U1015 (N_1015,In_2320,In_4433);
or U1016 (N_1016,In_1192,In_2910);
nor U1017 (N_1017,In_3988,In_3538);
nor U1018 (N_1018,In_3764,In_4286);
and U1019 (N_1019,In_316,In_1986);
nor U1020 (N_1020,In_3836,In_2356);
or U1021 (N_1021,In_2256,In_4088);
nor U1022 (N_1022,In_4764,In_3849);
or U1023 (N_1023,In_255,In_3075);
and U1024 (N_1024,In_4182,In_317);
or U1025 (N_1025,In_4677,In_2409);
and U1026 (N_1026,In_4940,In_1230);
xor U1027 (N_1027,In_3637,In_4026);
nor U1028 (N_1028,In_1323,In_1943);
and U1029 (N_1029,In_2504,In_4962);
xor U1030 (N_1030,In_909,In_45);
nor U1031 (N_1031,In_1103,In_1423);
xnor U1032 (N_1032,In_4450,In_116);
nand U1033 (N_1033,In_2350,In_2336);
nor U1034 (N_1034,In_563,In_2233);
nand U1035 (N_1035,In_4815,In_4552);
xor U1036 (N_1036,In_4360,In_3251);
nand U1037 (N_1037,In_4646,In_2283);
nor U1038 (N_1038,In_603,In_1869);
and U1039 (N_1039,In_2628,In_4096);
nor U1040 (N_1040,In_2438,In_363);
xor U1041 (N_1041,In_84,In_3271);
and U1042 (N_1042,In_2012,In_3819);
or U1043 (N_1043,In_2285,In_495);
nand U1044 (N_1044,In_3115,In_233);
xor U1045 (N_1045,In_2857,In_2654);
nor U1046 (N_1046,In_2518,In_621);
or U1047 (N_1047,In_2871,In_1606);
or U1048 (N_1048,In_3563,In_1493);
xnor U1049 (N_1049,In_3057,In_2897);
nor U1050 (N_1050,In_1686,In_3958);
nand U1051 (N_1051,In_3293,In_3301);
xnor U1052 (N_1052,In_4761,In_129);
nor U1053 (N_1053,In_917,In_1766);
or U1054 (N_1054,In_3660,In_4158);
nor U1055 (N_1055,In_4793,In_2818);
xor U1056 (N_1056,In_1306,In_3601);
xnor U1057 (N_1057,In_1421,In_3939);
or U1058 (N_1058,In_3377,In_3360);
nand U1059 (N_1059,In_3445,In_201);
nor U1060 (N_1060,In_2790,In_1328);
and U1061 (N_1061,In_253,In_3872);
xor U1062 (N_1062,In_2939,In_1849);
and U1063 (N_1063,In_1533,In_2360);
or U1064 (N_1064,In_571,In_2831);
xor U1065 (N_1065,In_4625,In_1628);
and U1066 (N_1066,In_2580,In_3202);
nor U1067 (N_1067,In_550,In_1494);
or U1068 (N_1068,In_17,In_4118);
nor U1069 (N_1069,In_3073,In_216);
and U1070 (N_1070,In_2848,In_4297);
xor U1071 (N_1071,In_4787,In_4150);
and U1072 (N_1072,In_4464,In_4875);
nor U1073 (N_1073,In_3441,In_2827);
nor U1074 (N_1074,In_3053,In_1985);
and U1075 (N_1075,In_4801,In_242);
nand U1076 (N_1076,In_4082,In_3703);
nand U1077 (N_1077,In_2754,In_2472);
and U1078 (N_1078,In_220,In_681);
and U1079 (N_1079,In_1860,In_285);
nor U1080 (N_1080,In_733,In_774);
xnor U1081 (N_1081,In_1274,In_900);
xnor U1082 (N_1082,In_2142,In_3678);
nand U1083 (N_1083,In_4029,In_2048);
nor U1084 (N_1084,In_2669,In_4206);
and U1085 (N_1085,In_2068,In_825);
xnor U1086 (N_1086,In_2603,In_159);
nor U1087 (N_1087,In_1498,In_3303);
nand U1088 (N_1088,In_2985,In_1431);
xor U1089 (N_1089,In_3442,In_4395);
and U1090 (N_1090,In_2753,In_671);
and U1091 (N_1091,In_2265,In_3120);
nor U1092 (N_1092,In_535,In_2003);
or U1093 (N_1093,In_773,In_1029);
or U1094 (N_1094,In_2501,In_2379);
nor U1095 (N_1095,In_1158,In_4795);
and U1096 (N_1096,In_857,In_494);
nand U1097 (N_1097,In_350,In_4290);
nand U1098 (N_1098,In_3320,In_1240);
nor U1099 (N_1099,In_4657,In_1843);
nand U1100 (N_1100,In_2081,In_1732);
or U1101 (N_1101,In_1880,In_1778);
and U1102 (N_1102,In_2094,In_4587);
nand U1103 (N_1103,In_1285,In_3514);
nor U1104 (N_1104,In_2923,In_171);
nor U1105 (N_1105,In_3995,In_2520);
nor U1106 (N_1106,In_1729,In_4782);
nor U1107 (N_1107,In_3754,In_368);
nor U1108 (N_1108,In_3604,In_2227);
xor U1109 (N_1109,In_112,In_2870);
and U1110 (N_1110,In_4437,In_2656);
nor U1111 (N_1111,In_225,In_14);
nor U1112 (N_1112,In_2595,In_4916);
nor U1113 (N_1113,In_1486,In_1185);
xor U1114 (N_1114,In_4494,In_3614);
nand U1115 (N_1115,In_181,In_459);
nor U1116 (N_1116,In_2213,In_3460);
nor U1117 (N_1117,In_4319,In_2927);
and U1118 (N_1118,In_4034,In_4799);
xor U1119 (N_1119,In_1131,In_2153);
nand U1120 (N_1120,In_2299,In_1420);
xnor U1121 (N_1121,In_4861,In_1022);
xor U1122 (N_1122,In_624,In_2053);
xor U1123 (N_1123,In_4590,In_4967);
nor U1124 (N_1124,In_1856,In_4309);
and U1125 (N_1125,In_2492,In_798);
nand U1126 (N_1126,In_3332,In_1215);
nand U1127 (N_1127,In_1065,In_1739);
and U1128 (N_1128,In_4364,In_2100);
or U1129 (N_1129,In_4727,In_3250);
nand U1130 (N_1130,In_2062,In_4742);
xnor U1131 (N_1131,In_3737,In_38);
or U1132 (N_1132,In_1585,In_4399);
xnor U1133 (N_1133,In_3668,In_2140);
nor U1134 (N_1134,In_646,In_1636);
xnor U1135 (N_1135,In_4687,In_4980);
or U1136 (N_1136,In_4643,In_48);
or U1137 (N_1137,In_2792,In_850);
and U1138 (N_1138,In_2330,In_542);
nand U1139 (N_1139,In_3724,In_457);
and U1140 (N_1140,In_1367,In_886);
nand U1141 (N_1141,In_126,In_3884);
nor U1142 (N_1142,In_1612,In_2788);
nand U1143 (N_1143,In_334,In_2623);
nor U1144 (N_1144,In_4060,In_2726);
nor U1145 (N_1145,In_3793,In_2269);
nand U1146 (N_1146,In_2928,In_3985);
or U1147 (N_1147,In_1975,In_767);
or U1148 (N_1148,In_4937,In_4520);
nor U1149 (N_1149,In_2644,In_3774);
nand U1150 (N_1150,In_3821,In_29);
nor U1151 (N_1151,In_312,In_412);
and U1152 (N_1152,In_2830,In_4850);
nor U1153 (N_1153,In_4593,In_778);
and U1154 (N_1154,In_3728,In_1461);
or U1155 (N_1155,In_3206,In_985);
nor U1156 (N_1156,In_3685,In_260);
nor U1157 (N_1157,In_4417,In_4483);
or U1158 (N_1158,In_1738,In_4824);
and U1159 (N_1159,In_2626,In_3385);
nand U1160 (N_1160,In_1604,In_1737);
nand U1161 (N_1161,In_3480,In_1866);
xnor U1162 (N_1162,In_325,In_1346);
xor U1163 (N_1163,In_1184,In_3034);
nand U1164 (N_1164,In_2982,In_818);
nor U1165 (N_1165,In_3339,In_54);
xor U1166 (N_1166,In_2730,In_1127);
and U1167 (N_1167,In_2065,In_4259);
xnor U1168 (N_1168,In_4639,In_1315);
nor U1169 (N_1169,In_4090,In_4992);
or U1170 (N_1170,In_1974,In_3286);
xor U1171 (N_1171,In_1590,In_2944);
xor U1172 (N_1172,In_398,In_552);
nor U1173 (N_1173,In_994,In_2721);
nand U1174 (N_1174,In_239,In_4842);
and U1175 (N_1175,In_3778,In_1887);
nor U1176 (N_1176,In_1237,In_4387);
nand U1177 (N_1177,In_911,In_120);
xnor U1178 (N_1178,In_2977,In_4044);
nor U1179 (N_1179,In_2883,In_3509);
nand U1180 (N_1180,In_3548,In_1818);
xnor U1181 (N_1181,In_2591,In_988);
and U1182 (N_1182,In_2399,In_2401);
or U1183 (N_1183,In_3650,In_1262);
or U1184 (N_1184,In_4218,In_3372);
nand U1185 (N_1185,In_3591,In_3534);
or U1186 (N_1186,In_569,In_3755);
nor U1187 (N_1187,In_3326,In_4002);
xnor U1188 (N_1188,In_4528,In_1822);
or U1189 (N_1189,In_2638,In_3581);
nor U1190 (N_1190,In_3336,In_4020);
or U1191 (N_1191,In_3739,In_1702);
and U1192 (N_1192,In_2257,In_4071);
nand U1193 (N_1193,In_2043,In_2218);
or U1194 (N_1194,In_357,In_4862);
and U1195 (N_1195,In_666,In_3478);
and U1196 (N_1196,In_2084,In_1815);
nand U1197 (N_1197,In_4167,In_1241);
nand U1198 (N_1198,In_1808,In_2854);
xor U1199 (N_1199,In_4237,In_1774);
xnor U1200 (N_1200,In_4720,In_2761);
and U1201 (N_1201,In_4943,In_711);
and U1202 (N_1202,In_2061,In_1666);
nand U1203 (N_1203,In_531,In_2687);
and U1204 (N_1204,In_2565,In_148);
nand U1205 (N_1205,In_4235,In_1438);
nand U1206 (N_1206,In_834,In_4919);
nand U1207 (N_1207,In_589,In_4076);
nor U1208 (N_1208,In_2148,In_943);
and U1209 (N_1209,In_540,In_4390);
or U1210 (N_1210,In_1179,In_1819);
or U1211 (N_1211,In_4810,In_3702);
and U1212 (N_1212,In_2370,In_1227);
nor U1213 (N_1213,In_1538,In_2423);
or U1214 (N_1214,In_2548,In_4379);
xor U1215 (N_1215,In_546,In_4510);
xor U1216 (N_1216,In_3571,In_674);
or U1217 (N_1217,In_3424,In_3868);
nand U1218 (N_1218,In_3444,In_2797);
xor U1219 (N_1219,In_936,In_4248);
or U1220 (N_1220,In_3779,In_2903);
nand U1221 (N_1221,In_608,In_2179);
or U1222 (N_1222,In_4231,In_382);
and U1223 (N_1223,In_3283,In_4305);
and U1224 (N_1224,In_435,In_3669);
nand U1225 (N_1225,In_2582,In_4959);
nand U1226 (N_1226,In_27,In_82);
or U1227 (N_1227,In_1993,In_1786);
nand U1228 (N_1228,In_4613,In_1644);
or U1229 (N_1229,In_97,In_4988);
xnor U1230 (N_1230,In_1310,In_1354);
xor U1231 (N_1231,In_2226,In_1643);
nand U1232 (N_1232,In_1532,In_4159);
nand U1233 (N_1233,In_2633,In_1497);
or U1234 (N_1234,In_1509,In_1337);
and U1235 (N_1235,In_308,In_2369);
xor U1236 (N_1236,In_3043,In_1385);
xnor U1237 (N_1237,In_326,In_2458);
nor U1238 (N_1238,In_1234,In_4841);
xor U1239 (N_1239,In_1649,In_3733);
and U1240 (N_1240,In_4277,In_4308);
nand U1241 (N_1241,In_811,In_2418);
and U1242 (N_1242,In_1610,In_353);
nand U1243 (N_1243,In_446,In_3376);
or U1244 (N_1244,In_756,In_3291);
nand U1245 (N_1245,In_4359,In_128);
nor U1246 (N_1246,In_2625,In_2667);
nor U1247 (N_1247,In_3522,In_2576);
or U1248 (N_1248,In_1064,In_484);
nand U1249 (N_1249,In_1369,In_3770);
nor U1250 (N_1250,In_2178,In_1995);
or U1251 (N_1251,In_3941,In_4239);
and U1252 (N_1252,In_2476,In_4276);
nand U1253 (N_1253,In_1665,In_1580);
and U1254 (N_1254,In_3782,In_3039);
or U1255 (N_1255,In_3393,In_514);
or U1256 (N_1256,In_591,In_73);
or U1257 (N_1257,In_65,In_898);
nand U1258 (N_1258,In_293,In_4645);
nor U1259 (N_1259,In_2345,In_1027);
and U1260 (N_1260,In_498,In_2579);
or U1261 (N_1261,In_456,In_263);
or U1262 (N_1262,In_4263,In_4036);
nor U1263 (N_1263,In_130,In_1901);
and U1264 (N_1264,In_826,In_3729);
nor U1265 (N_1265,In_10,In_3888);
xor U1266 (N_1266,In_100,In_1162);
or U1267 (N_1267,In_2964,In_3800);
nor U1268 (N_1268,In_2581,In_3965);
or U1269 (N_1269,In_111,In_1204);
and U1270 (N_1270,In_4738,In_759);
xor U1271 (N_1271,In_4816,In_1800);
nand U1272 (N_1272,In_3731,In_2449);
nor U1273 (N_1273,In_301,In_2740);
and U1274 (N_1274,In_2319,In_2463);
or U1275 (N_1275,In_4422,In_2934);
nor U1276 (N_1276,In_1659,In_2210);
and U1277 (N_1277,In_454,In_2166);
or U1278 (N_1278,In_3797,In_1977);
nand U1279 (N_1279,In_1261,In_250);
nand U1280 (N_1280,In_998,In_1560);
nand U1281 (N_1281,In_3565,In_949);
xnor U1282 (N_1282,In_2890,In_2066);
nor U1283 (N_1283,In_830,In_1181);
nor U1284 (N_1284,In_4882,In_2325);
nor U1285 (N_1285,In_3975,In_2277);
nor U1286 (N_1286,In_3946,In_3828);
nand U1287 (N_1287,In_4015,In_2570);
or U1288 (N_1288,In_945,In_1857);
xor U1289 (N_1289,In_1226,In_3257);
and U1290 (N_1290,In_1460,In_829);
nand U1291 (N_1291,In_1671,In_2617);
or U1292 (N_1292,In_3035,In_3221);
xnor U1293 (N_1293,In_2802,In_1010);
xor U1294 (N_1294,In_751,In_304);
nor U1295 (N_1295,In_4833,In_2796);
nand U1296 (N_1296,In_3670,In_3181);
xor U1297 (N_1297,In_3164,In_4303);
or U1298 (N_1298,In_1683,In_1297);
nor U1299 (N_1299,In_2787,In_4616);
nand U1300 (N_1300,In_1728,In_588);
nor U1301 (N_1301,In_394,In_307);
xnor U1302 (N_1302,In_4214,In_2598);
or U1303 (N_1303,In_4722,In_1021);
xnor U1304 (N_1304,In_2275,In_3051);
or U1305 (N_1305,In_3602,In_567);
or U1306 (N_1306,In_4383,In_1006);
nor U1307 (N_1307,In_4714,In_2339);
and U1308 (N_1308,In_3840,In_3256);
or U1309 (N_1309,In_3112,In_99);
xor U1310 (N_1310,In_3896,In_3231);
nand U1311 (N_1311,In_4594,In_2220);
nor U1312 (N_1312,In_4960,In_4207);
nand U1313 (N_1313,In_373,In_1551);
xor U1314 (N_1314,In_3639,In_3022);
and U1315 (N_1315,In_3846,In_3771);
nor U1316 (N_1316,In_2077,In_1443);
or U1317 (N_1317,In_1238,In_3125);
xnor U1318 (N_1318,In_1531,In_232);
or U1319 (N_1319,In_1362,In_701);
and U1320 (N_1320,In_3218,In_3682);
and U1321 (N_1321,In_2971,In_2333);
nor U1322 (N_1322,In_3980,In_4733);
xor U1323 (N_1323,In_1133,In_2465);
xor U1324 (N_1324,In_4465,In_3473);
xnor U1325 (N_1325,In_2942,In_3718);
or U1326 (N_1326,In_776,In_1970);
or U1327 (N_1327,In_2432,In_4039);
nand U1328 (N_1328,In_3903,In_833);
xnor U1329 (N_1329,In_990,In_192);
nand U1330 (N_1330,In_3583,In_3459);
nand U1331 (N_1331,In_3253,In_3142);
nand U1332 (N_1332,In_3715,In_3665);
nor U1333 (N_1333,In_4441,In_3471);
and U1334 (N_1334,In_1920,In_2706);
nor U1335 (N_1335,In_1434,In_2751);
nand U1336 (N_1336,In_4242,In_1848);
or U1337 (N_1337,In_1122,In_168);
or U1338 (N_1338,In_786,In_4367);
nand U1339 (N_1339,In_4178,In_3893);
or U1340 (N_1340,In_4540,In_3227);
nor U1341 (N_1341,In_381,In_2008);
or U1342 (N_1342,In_1685,In_1201);
xor U1343 (N_1343,In_865,In_3236);
and U1344 (N_1344,In_1756,In_702);
nor U1345 (N_1345,In_4922,In_1300);
nor U1346 (N_1346,In_4252,In_3101);
or U1347 (N_1347,In_4917,In_3830);
xor U1348 (N_1348,In_1294,In_1806);
xor U1349 (N_1349,In_1110,In_3265);
nor U1350 (N_1350,In_1099,In_1704);
or U1351 (N_1351,In_4753,In_1154);
nor U1352 (N_1352,In_4085,In_3347);
and U1353 (N_1353,In_1296,In_4789);
or U1354 (N_1354,In_4255,In_854);
nand U1355 (N_1355,In_925,In_1030);
xnor U1356 (N_1356,In_3211,In_1147);
xnor U1357 (N_1357,In_1176,In_1342);
xnor U1358 (N_1358,In_4027,In_1149);
and U1359 (N_1359,In_3621,In_2891);
nand U1360 (N_1360,In_984,In_4163);
and U1361 (N_1361,In_1198,In_1594);
or U1362 (N_1362,In_2774,In_3875);
nor U1363 (N_1363,In_4580,In_4848);
xnor U1364 (N_1364,In_1251,In_3413);
xor U1365 (N_1365,In_1063,In_3631);
nand U1366 (N_1366,In_3044,In_3753);
nand U1367 (N_1367,In_2085,In_3342);
nand U1368 (N_1368,In_142,In_1088);
nor U1369 (N_1369,In_1485,In_3899);
nand U1370 (N_1370,In_1698,In_819);
xor U1371 (N_1371,In_2035,In_1109);
nand U1372 (N_1372,In_3543,In_2713);
nand U1373 (N_1373,In_2353,In_2108);
nor U1374 (N_1374,In_4386,In_3521);
and U1375 (N_1375,In_4256,In_772);
xor U1376 (N_1376,In_4589,In_1414);
and U1377 (N_1377,In_3488,In_1056);
nor U1378 (N_1378,In_3259,In_2);
nand U1379 (N_1379,In_4539,In_3991);
and U1380 (N_1380,In_3587,In_704);
xor U1381 (N_1381,In_3815,In_3033);
nand U1382 (N_1382,In_4592,In_3483);
xnor U1383 (N_1383,In_1626,In_3654);
and U1384 (N_1384,In_788,In_1456);
nor U1385 (N_1385,In_4920,In_1973);
or U1386 (N_1386,In_2748,In_1508);
and U1387 (N_1387,In_4223,In_4718);
nor U1388 (N_1388,In_1121,In_2768);
xnor U1389 (N_1389,In_3968,In_3176);
and U1390 (N_1390,In_1890,In_977);
nor U1391 (N_1391,In_4930,In_3951);
and U1392 (N_1392,In_1569,In_2083);
or U1393 (N_1393,In_274,In_401);
nor U1394 (N_1394,In_1393,In_1417);
xor U1395 (N_1395,In_924,In_1622);
nand U1396 (N_1396,In_2137,In_1624);
xnor U1397 (N_1397,In_4400,In_1952);
or U1398 (N_1398,In_440,In_1171);
xor U1399 (N_1399,In_4559,In_3150);
nand U1400 (N_1400,In_4128,In_4016);
nor U1401 (N_1401,In_4642,In_1935);
and U1402 (N_1402,In_4352,In_3394);
xnor U1403 (N_1403,In_1004,In_3923);
nor U1404 (N_1404,In_41,In_1186);
nand U1405 (N_1405,In_3783,In_247);
or U1406 (N_1406,In_4837,In_2846);
xnor U1407 (N_1407,In_4863,In_1599);
xor U1408 (N_1408,In_1542,In_362);
nand U1409 (N_1409,In_2684,In_3628);
or U1410 (N_1410,In_1320,In_4544);
and U1411 (N_1411,In_4416,In_4268);
or U1412 (N_1412,In_3938,In_3013);
or U1413 (N_1413,In_210,In_1334);
nand U1414 (N_1414,In_2522,In_2597);
and U1415 (N_1415,In_2599,In_887);
xnor U1416 (N_1416,In_1054,In_2406);
nand U1417 (N_1417,In_3659,In_2052);
nand U1418 (N_1418,In_1092,In_4017);
nor U1419 (N_1419,In_2047,In_2904);
nor U1420 (N_1420,In_4181,In_1564);
xor U1421 (N_1421,In_1518,In_415);
and U1422 (N_1422,In_3727,In_1725);
xor U1423 (N_1423,In_3890,In_698);
nor U1424 (N_1424,In_1559,In_3834);
nor U1425 (N_1425,In_4609,In_311);
or U1426 (N_1426,In_2499,In_1763);
nor U1427 (N_1427,In_2201,In_1472);
nor U1428 (N_1428,In_2868,In_1304);
and U1429 (N_1429,In_1562,In_324);
xnor U1430 (N_1430,In_2402,In_2453);
xor U1431 (N_1431,In_4050,In_1487);
xnor U1432 (N_1432,In_1733,In_2027);
and U1433 (N_1433,In_2820,In_195);
nand U1434 (N_1434,In_106,In_2583);
nand U1435 (N_1435,In_4652,In_444);
and U1436 (N_1436,In_2604,In_110);
nand U1437 (N_1437,In_3510,In_346);
or U1438 (N_1438,In_4377,In_141);
nor U1439 (N_1439,In_1003,In_329);
nand U1440 (N_1440,In_1678,In_4463);
and U1441 (N_1441,In_876,In_1695);
nand U1442 (N_1442,In_1067,In_2397);
nor U1443 (N_1443,In_615,In_1637);
nor U1444 (N_1444,In_647,In_1245);
nor U1445 (N_1445,In_2712,In_4112);
nand U1446 (N_1446,In_1052,In_2503);
nor U1447 (N_1447,In_2951,In_3430);
and U1448 (N_1448,In_3174,In_2860);
or U1449 (N_1449,In_636,In_3588);
xnor U1450 (N_1450,In_3359,In_2813);
nor U1451 (N_1451,In_4199,In_4317);
or U1452 (N_1452,In_3082,In_1470);
and U1453 (N_1453,In_3268,In_686);
or U1454 (N_1454,In_3648,In_4419);
nand U1455 (N_1455,In_2678,In_2264);
nor U1456 (N_1456,In_1151,In_2952);
nor U1457 (N_1457,In_3224,In_2292);
nor U1458 (N_1458,In_4009,In_4241);
and U1459 (N_1459,In_3299,In_57);
or U1460 (N_1460,In_2295,In_3212);
or U1461 (N_1461,In_1574,In_643);
xor U1462 (N_1462,In_2327,In_4887);
xnor U1463 (N_1463,In_3698,In_4078);
and U1464 (N_1464,In_816,In_295);
nand U1465 (N_1465,In_208,In_1703);
nor U1466 (N_1466,In_3479,In_1979);
nand U1467 (N_1467,In_4330,In_511);
nand U1468 (N_1468,In_4180,In_2528);
xnor U1469 (N_1469,In_4847,In_744);
nand U1470 (N_1470,In_1035,In_1660);
and U1471 (N_1471,In_679,In_1448);
and U1472 (N_1472,In_296,In_3140);
or U1473 (N_1473,In_1905,In_651);
or U1474 (N_1474,In_4219,In_4712);
xor U1475 (N_1475,In_1190,In_823);
nand U1476 (N_1476,In_4147,In_2605);
nand U1477 (N_1477,In_1229,In_4650);
nand U1478 (N_1478,In_4906,In_1964);
and U1479 (N_1479,In_1667,In_875);
nor U1480 (N_1480,In_4866,In_2688);
or U1481 (N_1481,In_2767,In_4550);
nor U1482 (N_1482,In_1776,In_391);
nand U1483 (N_1483,In_4956,In_104);
xor U1484 (N_1484,In_3248,In_342);
or U1485 (N_1485,In_499,In_3515);
or U1486 (N_1486,In_2009,In_3843);
nand U1487 (N_1487,In_198,In_1515);
xor U1488 (N_1488,In_1000,In_3338);
nand U1489 (N_1489,In_1833,In_2873);
xnor U1490 (N_1490,In_663,In_3133);
and U1491 (N_1491,In_3937,In_1961);
nor U1492 (N_1492,In_779,In_3309);
nor U1493 (N_1493,In_2222,In_2629);
nor U1494 (N_1494,In_862,In_4200);
xor U1495 (N_1495,In_518,In_2590);
nor U1496 (N_1496,In_4405,In_2249);
nor U1497 (N_1497,In_1962,In_3549);
and U1498 (N_1498,In_1479,In_4621);
nor U1499 (N_1499,In_1550,In_3651);
or U1500 (N_1500,In_1312,In_206);
nand U1501 (N_1501,In_3254,In_2493);
nor U1502 (N_1502,In_4337,In_4394);
and U1503 (N_1503,In_1707,In_987);
or U1504 (N_1504,In_1588,In_3106);
and U1505 (N_1505,In_2347,In_4435);
xor U1506 (N_1506,In_2128,In_3734);
and U1507 (N_1507,In_1558,In_2496);
or U1508 (N_1508,In_680,In_958);
nand U1509 (N_1509,In_723,In_4024);
xnor U1510 (N_1510,In_1389,In_3436);
nor U1511 (N_1511,In_700,In_4904);
nand U1512 (N_1512,In_479,In_3240);
and U1513 (N_1513,In_1689,In_4692);
nand U1514 (N_1514,In_2442,In_4037);
nand U1515 (N_1515,In_3949,In_1386);
nand U1516 (N_1516,In_1330,In_1014);
nand U1517 (N_1517,In_4227,In_1570);
and U1518 (N_1518,In_4562,In_713);
and U1519 (N_1519,In_2702,In_1942);
or U1520 (N_1520,In_2541,In_1098);
and U1521 (N_1521,In_2718,In_4851);
or U1522 (N_1522,In_481,In_1851);
xnor U1523 (N_1523,In_2561,In_5);
nand U1524 (N_1524,In_2803,In_4518);
nor U1525 (N_1525,In_1557,In_3775);
and U1526 (N_1526,In_2430,In_3354);
and U1527 (N_1527,In_1178,In_3482);
nor U1528 (N_1528,In_2247,In_968);
xnor U1529 (N_1529,In_3694,In_404);
xnor U1530 (N_1530,In_330,In_2126);
nand U1531 (N_1531,In_3865,In_2677);
or U1532 (N_1532,In_1798,In_1044);
nor U1533 (N_1533,In_1307,In_4600);
xor U1534 (N_1534,In_2855,In_158);
or U1535 (N_1535,In_3969,In_3009);
or U1536 (N_1536,In_1380,In_3086);
xor U1537 (N_1537,In_1799,In_2186);
nor U1538 (N_1538,In_3503,In_3121);
nor U1539 (N_1539,In_3325,In_172);
nand U1540 (N_1540,In_3007,In_3080);
or U1541 (N_1541,In_2268,In_1584);
nand U1542 (N_1542,In_2141,In_2719);
and U1543 (N_1543,In_139,In_4056);
or U1544 (N_1544,In_3200,In_2689);
xnor U1545 (N_1545,In_539,In_1293);
nand U1546 (N_1546,In_3011,In_2071);
nor U1547 (N_1547,In_1813,In_1352);
and U1548 (N_1548,In_3134,In_2063);
nor U1549 (N_1549,In_976,In_1537);
and U1550 (N_1550,In_1745,In_4511);
nand U1551 (N_1551,In_4137,In_4649);
nor U1552 (N_1552,In_4327,In_1858);
or U1553 (N_1553,In_2235,In_1450);
or U1554 (N_1554,In_3105,In_335);
and U1555 (N_1555,In_4134,In_4772);
xor U1556 (N_1556,In_677,In_2405);
xor U1557 (N_1557,In_3597,In_2482);
nand U1558 (N_1558,In_975,In_1270);
xnor U1559 (N_1559,In_2400,In_3996);
and U1560 (N_1560,In_3453,In_2428);
nor U1561 (N_1561,In_734,In_579);
or U1562 (N_1562,In_3209,In_2615);
and U1563 (N_1563,In_3486,In_4894);
or U1564 (N_1564,In_1457,In_2199);
and U1565 (N_1565,In_1341,In_1205);
nor U1566 (N_1566,In_1406,In_3857);
and U1567 (N_1567,In_3123,In_585);
nor U1568 (N_1568,In_2546,In_2558);
and U1569 (N_1569,In_2697,In_690);
nand U1570 (N_1570,In_273,In_3877);
xor U1571 (N_1571,In_114,In_4136);
or U1572 (N_1572,In_999,In_3411);
nand U1573 (N_1573,In_4121,In_3406);
nand U1574 (N_1574,In_3855,In_1455);
xnor U1575 (N_1575,In_2745,In_2823);
xor U1576 (N_1576,In_1268,In_3433);
nand U1577 (N_1577,In_3902,In_4361);
xor U1578 (N_1578,In_2594,In_3331);
nand U1579 (N_1579,In_709,In_1080);
and U1580 (N_1580,In_522,In_2894);
xnor U1581 (N_1581,In_4142,In_3498);
nor U1582 (N_1582,In_3408,In_3572);
xor U1583 (N_1583,In_3546,In_4950);
and U1584 (N_1584,In_1988,In_4897);
nor U1585 (N_1585,In_2274,In_4328);
and U1586 (N_1586,In_3912,In_2229);
nor U1587 (N_1587,In_2305,In_53);
and U1588 (N_1588,In_42,In_1135);
nor U1589 (N_1589,In_645,In_3069);
nand U1590 (N_1590,In_1496,In_4049);
nor U1591 (N_1591,In_3603,In_1356);
nand U1592 (N_1592,In_584,In_4285);
or U1593 (N_1593,In_1231,In_2025);
xor U1594 (N_1594,In_3706,In_4109);
or U1595 (N_1595,In_1013,In_673);
nor U1596 (N_1596,In_4100,In_3921);
xor U1597 (N_1597,In_2732,In_3455);
xor U1598 (N_1598,In_1002,In_3740);
and U1599 (N_1599,In_3065,In_2212);
nand U1600 (N_1600,In_3979,In_1311);
and U1601 (N_1601,In_2180,In_2392);
and U1602 (N_1602,In_2759,In_4420);
nor U1603 (N_1603,In_1105,In_3333);
nor U1604 (N_1604,In_3087,In_4603);
and U1605 (N_1605,In_855,In_639);
nand U1606 (N_1606,In_724,In_2267);
nor U1607 (N_1607,In_4553,In_1480);
nand U1608 (N_1608,In_1361,In_4558);
and U1609 (N_1609,In_4868,In_1043);
or U1610 (N_1610,In_147,In_4905);
nand U1611 (N_1611,In_4371,In_4089);
and U1612 (N_1612,In_2000,In_3635);
or U1613 (N_1613,In_483,In_3679);
and U1614 (N_1614,In_1256,In_2473);
nand U1615 (N_1615,In_1091,In_4910);
nor U1616 (N_1616,In_3692,In_3487);
nor U1617 (N_1617,In_2271,In_3005);
or U1618 (N_1618,In_676,In_1217);
nor U1619 (N_1619,In_1408,In_3530);
or U1620 (N_1620,In_2800,In_2074);
nand U1621 (N_1621,In_1908,In_2569);
nand U1622 (N_1622,In_1899,In_91);
xnor U1623 (N_1623,In_166,In_1491);
and U1624 (N_1624,In_794,In_1086);
and U1625 (N_1625,In_1390,In_3461);
nand U1626 (N_1626,In_3368,In_4864);
xnor U1627 (N_1627,In_4570,In_661);
or U1628 (N_1628,In_1228,In_202);
nand U1629 (N_1629,In_2825,In_3813);
xnor U1630 (N_1630,In_1255,In_4627);
nand U1631 (N_1631,In_3421,In_2460);
nor U1632 (N_1632,In_4312,In_455);
nand U1633 (N_1633,In_1081,In_194);
and U1634 (N_1634,In_1877,In_1325);
and U1635 (N_1635,In_2571,In_489);
nor U1636 (N_1636,In_933,In_1298);
nand U1637 (N_1637,In_1376,In_4488);
and U1638 (N_1638,In_844,In_3047);
and U1639 (N_1639,In_3384,In_2016);
and U1640 (N_1640,In_777,In_4421);
nand U1641 (N_1641,In_2294,In_25);
nand U1642 (N_1642,In_1708,In_2477);
nor U1643 (N_1643,In_4351,In_4103);
nor U1644 (N_1644,In_9,In_882);
nor U1645 (N_1645,In_3570,In_678);
and U1646 (N_1646,In_4130,In_3169);
and U1647 (N_1647,In_2215,In_3014);
or U1648 (N_1648,In_4605,In_425);
xor U1649 (N_1649,In_2842,In_3766);
nand U1650 (N_1650,In_2101,In_237);
xnor U1651 (N_1651,In_1292,In_1934);
xor U1652 (N_1652,In_3891,In_837);
and U1653 (N_1653,In_3634,In_2374);
nand U1654 (N_1654,In_3773,In_3605);
or U1655 (N_1655,In_4038,In_3144);
nor U1656 (N_1656,In_4425,In_747);
nand U1657 (N_1657,In_1971,In_1061);
xor U1658 (N_1658,In_4183,In_4455);
nor U1659 (N_1659,In_2884,In_370);
nand U1660 (N_1660,In_1984,In_4471);
xor U1661 (N_1661,In_3675,In_1276);
or U1662 (N_1662,In_2785,In_3151);
nand U1663 (N_1663,In_4805,In_4941);
xor U1664 (N_1664,In_3541,In_1931);
and U1665 (N_1665,In_1273,In_3919);
nand U1666 (N_1666,In_4195,In_4424);
or U1667 (N_1667,In_4320,In_1394);
and U1668 (N_1668,In_2056,In_4407);
or U1669 (N_1669,In_397,In_1633);
or U1670 (N_1670,In_4156,In_2416);
xor U1671 (N_1671,In_726,In_2291);
nand U1672 (N_1672,In_4062,In_4852);
xor U1673 (N_1673,In_4601,In_1263);
xor U1674 (N_1674,In_2377,In_4216);
and U1675 (N_1675,In_3664,In_1999);
nor U1676 (N_1676,In_727,In_3553);
nand U1677 (N_1677,In_1040,In_4339);
and U1678 (N_1678,In_3272,In_2136);
or U1679 (N_1679,In_1453,In_3042);
or U1680 (N_1680,In_3199,In_327);
or U1681 (N_1681,In_566,In_959);
and U1682 (N_1682,In_989,In_3191);
nand U1683 (N_1683,In_2783,In_1797);
and U1684 (N_1684,In_3316,In_500);
and U1685 (N_1685,In_2364,In_2494);
xnor U1686 (N_1686,In_3485,In_1465);
nor U1687 (N_1687,In_944,In_4667);
xor U1688 (N_1688,In_3920,In_1143);
and U1689 (N_1689,In_4110,In_2384);
nor U1690 (N_1690,In_2017,In_4470);
or U1691 (N_1691,In_1947,In_3262);
or U1692 (N_1692,In_4475,In_4773);
xor U1693 (N_1693,In_2192,In_4579);
or U1694 (N_1694,In_1681,In_1321);
nand U1695 (N_1695,In_328,In_1918);
or U1696 (N_1696,In_3239,In_4844);
nand U1697 (N_1697,In_2419,In_3725);
nor U1698 (N_1698,In_785,In_4629);
and U1699 (N_1699,In_835,In_619);
and U1700 (N_1700,In_115,In_4350);
nand U1701 (N_1701,In_2004,In_3914);
xor U1702 (N_1702,In_2743,In_4885);
nand U1703 (N_1703,In_2769,In_4171);
and U1704 (N_1704,In_4249,In_3742);
and U1705 (N_1705,In_3184,In_4706);
nor U1706 (N_1706,In_1412,In_1546);
xnor U1707 (N_1707,In_3984,In_721);
and U1708 (N_1708,In_1500,In_578);
nand U1709 (N_1709,In_4447,In_2979);
nor U1710 (N_1710,In_3178,In_4599);
nor U1711 (N_1711,In_4955,In_687);
nor U1712 (N_1712,In_3789,In_2278);
nand U1713 (N_1713,In_3119,In_87);
or U1714 (N_1714,In_4523,In_1272);
nor U1715 (N_1715,In_234,In_941);
nand U1716 (N_1716,In_3374,In_472);
nor U1717 (N_1717,In_4660,In_376);
xor U1718 (N_1718,In_545,In_4481);
nand U1719 (N_1719,In_3859,In_2396);
and U1720 (N_1720,In_3744,In_4438);
or U1721 (N_1721,In_2239,In_2642);
xnor U1722 (N_1722,In_2121,In_1283);
nor U1723 (N_1723,In_1329,In_4774);
or U1724 (N_1724,In_4978,In_125);
or U1725 (N_1725,In_1802,In_2572);
nand U1726 (N_1726,In_2457,In_2720);
xor U1727 (N_1727,In_3851,In_1418);
nor U1728 (N_1728,In_4093,In_961);
xnor U1729 (N_1729,In_4363,In_2795);
nor U1730 (N_1730,In_3304,In_2674);
or U1731 (N_1731,In_1156,In_4244);
xor U1732 (N_1732,In_4663,In_1501);
and U1733 (N_1733,In_3232,In_762);
xnor U1734 (N_1734,In_4734,In_79);
and U1735 (N_1735,In_601,In_3758);
or U1736 (N_1736,In_2840,In_180);
nand U1737 (N_1737,In_2044,In_3970);
nand U1738 (N_1738,In_1032,In_4385);
nand U1739 (N_1739,In_4184,In_2107);
nor U1740 (N_1740,In_1835,In_810);
xnor U1741 (N_1741,In_3716,In_4705);
and U1742 (N_1742,In_3964,In_2578);
xnor U1743 (N_1743,In_2258,In_4981);
or U1744 (N_1744,In_4778,In_1540);
or U1745 (N_1745,In_1587,In_1207);
xor U1746 (N_1746,In_1553,In_1058);
and U1747 (N_1747,In_3375,In_2673);
xor U1748 (N_1748,In_3396,In_513);
xor U1749 (N_1749,In_265,In_452);
nand U1750 (N_1750,In_3713,In_3873);
nand U1751 (N_1751,In_2205,In_1124);
xnor U1752 (N_1752,In_199,In_852);
and U1753 (N_1753,In_4999,In_441);
nor U1754 (N_1754,In_4061,In_375);
nor U1755 (N_1755,In_3451,In_3861);
nor U1756 (N_1756,In_2991,In_71);
xor U1757 (N_1757,In_1119,In_4230);
or U1758 (N_1758,In_2425,In_4574);
nand U1759 (N_1759,In_3076,In_1026);
or U1760 (N_1760,In_3992,In_3431);
or U1761 (N_1761,In_3363,In_2167);
xnor U1762 (N_1762,In_177,In_1868);
and U1763 (N_1763,In_3052,In_4700);
and U1764 (N_1764,In_4504,In_2075);
xor U1765 (N_1765,In_4853,In_592);
xor U1766 (N_1766,In_1426,In_3607);
nand U1767 (N_1767,In_717,In_2041);
and U1768 (N_1768,In_4270,In_2289);
or U1769 (N_1769,In_1430,In_4665);
and U1770 (N_1770,In_4921,In_1608);
and U1771 (N_1771,In_83,In_1108);
or U1772 (N_1772,In_1960,In_157);
and U1773 (N_1773,In_3234,In_1842);
xnor U1774 (N_1774,In_2816,In_691);
nand U1775 (N_1775,In_4710,In_1363);
nor U1776 (N_1776,In_2098,In_1008);
nor U1777 (N_1777,In_4974,In_657);
and U1778 (N_1778,In_1399,In_4185);
nor U1779 (N_1779,In_1060,In_3528);
and U1780 (N_1780,In_926,In_3277);
and U1781 (N_1781,In_3817,In_708);
or U1782 (N_1782,In_3462,In_1193);
nor U1783 (N_1783,In_858,In_548);
xor U1784 (N_1784,In_4355,In_841);
xor U1785 (N_1785,In_1696,In_2872);
xor U1786 (N_1786,In_3089,In_4472);
or U1787 (N_1787,In_219,In_3933);
or U1788 (N_1788,In_1308,In_1788);
and U1789 (N_1789,In_200,In_3874);
xnor U1790 (N_1790,In_2588,In_22);
and U1791 (N_1791,In_1248,In_2281);
or U1792 (N_1792,In_2115,In_812);
xnor U1793 (N_1793,In_1336,In_1998);
and U1794 (N_1794,In_174,In_3323);
nor U1795 (N_1795,In_2118,In_3371);
nor U1796 (N_1796,In_4083,In_685);
xor U1797 (N_1797,In_4388,In_1279);
and U1798 (N_1798,In_1929,In_2489);
xor U1799 (N_1799,In_2089,In_1554);
xnor U1800 (N_1800,In_3287,In_3193);
nand U1801 (N_1801,In_4838,In_4664);
or U1802 (N_1802,In_2162,In_732);
nor U1803 (N_1803,In_2189,In_2650);
xnor U1804 (N_1804,In_424,In_1291);
nand U1805 (N_1805,In_3366,In_3599);
xnor U1806 (N_1806,In_4743,In_1530);
xor U1807 (N_1807,In_814,In_2747);
nand U1808 (N_1808,In_289,In_336);
nand U1809 (N_1809,In_3100,In_4261);
nor U1810 (N_1810,In_283,In_1697);
nor U1811 (N_1811,In_1327,In_3420);
nand U1812 (N_1812,In_2087,In_2986);
nor U1813 (N_1813,In_2403,In_2515);
nand U1814 (N_1814,In_176,In_3862);
nand U1815 (N_1815,In_4891,In_705);
or U1816 (N_1816,In_377,In_4323);
and U1817 (N_1817,In_4165,In_4238);
nand U1818 (N_1818,In_109,In_839);
or U1819 (N_1819,In_4451,In_2632);
nand U1820 (N_1820,In_1850,In_4548);
nor U1821 (N_1821,In_93,In_4418);
nor U1822 (N_1822,In_2559,In_2302);
nor U1823 (N_1823,In_3467,In_4201);
nor U1824 (N_1824,In_1653,In_3556);
and U1825 (N_1825,In_2600,In_2152);
nand U1826 (N_1826,In_2188,In_1223);
or U1827 (N_1827,In_4683,In_2607);
or U1828 (N_1828,In_3743,In_662);
nand U1829 (N_1829,In_3021,In_3493);
or U1830 (N_1830,In_1712,In_3786);
xor U1831 (N_1831,In_2841,In_2393);
nand U1832 (N_1832,In_1349,In_4188);
xor U1833 (N_1833,In_1404,In_3018);
and U1834 (N_1834,In_178,In_1528);
or U1835 (N_1835,In_1894,In_2488);
nand U1836 (N_1836,In_3852,In_2387);
nand U1837 (N_1837,In_2069,In_2738);
and U1838 (N_1838,In_986,In_3313);
and U1839 (N_1839,In_4617,In_1442);
nand U1840 (N_1840,In_3315,In_3917);
nand U1841 (N_1841,In_151,In_2200);
xnor U1842 (N_1842,In_728,In_4054);
nor U1843 (N_1843,In_4964,In_4509);
xnor U1844 (N_1844,In_3697,In_3024);
and U1845 (N_1845,In_2187,In_4307);
nor U1846 (N_1846,In_4236,In_1996);
nor U1847 (N_1847,In_1377,In_2462);
and U1848 (N_1848,In_1392,In_1524);
nor U1849 (N_1849,In_1152,In_4966);
or U1850 (N_1850,In_3041,In_1163);
nor U1851 (N_1851,In_2777,In_3863);
and U1852 (N_1852,In_3641,In_3145);
nor U1853 (N_1853,In_1792,In_3405);
and U1854 (N_1854,In_2467,In_618);
nand U1855 (N_1855,In_1452,In_2936);
nand U1856 (N_1856,In_4132,In_4368);
xor U1857 (N_1857,In_3294,In_2391);
nand U1858 (N_1858,In_4345,In_3810);
nor U1859 (N_1859,In_3576,In_1844);
and U1860 (N_1860,In_650,In_2992);
nor U1861 (N_1861,In_2691,In_443);
or U1862 (N_1862,In_458,In_167);
and U1863 (N_1863,In_4519,In_982);
nand U1864 (N_1864,In_2407,In_2862);
nand U1865 (N_1865,In_1366,In_2833);
or U1866 (N_1866,In_2701,In_2296);
nand U1867 (N_1867,In_347,In_4467);
nand U1868 (N_1868,In_1691,In_856);
xor U1869 (N_1869,In_2112,In_1896);
or U1870 (N_1870,In_1203,In_405);
nor U1871 (N_1871,In_2544,In_4892);
nor U1872 (N_1872,In_3127,In_294);
or U1873 (N_1873,In_248,In_338);
nor U1874 (N_1874,In_529,In_3642);
xor U1875 (N_1875,In_3410,In_117);
and U1876 (N_1876,In_1967,In_2914);
or U1877 (N_1877,In_524,In_2217);
xnor U1878 (N_1878,In_222,In_3696);
or U1879 (N_1879,In_1577,In_4502);
or U1880 (N_1880,In_4246,In_809);
or U1881 (N_1881,In_3137,In_3045);
xnor U1882 (N_1882,In_3545,In_4606);
nor U1883 (N_1883,In_2454,In_2536);
and U1884 (N_1884,In_3971,In_3449);
nand U1885 (N_1885,In_1932,In_2177);
nand U1886 (N_1886,In_2915,In_2809);
nor U1887 (N_1887,In_3832,In_574);
or U1888 (N_1888,In_2287,In_4716);
and U1889 (N_1889,In_1488,In_1675);
and U1890 (N_1890,In_3448,In_2049);
nand U1891 (N_1891,In_3173,In_3008);
nor U1892 (N_1892,In_1107,In_1083);
nand U1893 (N_1893,In_230,In_3418);
xnor U1894 (N_1894,In_4048,In_2895);
xnor U1895 (N_1895,In_4113,In_2711);
nand U1896 (N_1896,In_3093,In_2708);
and U1897 (N_1897,In_1595,In_3916);
nand U1898 (N_1898,In_2316,In_3183);
nand U1899 (N_1899,In_2926,In_319);
and U1900 (N_1900,In_2367,In_4401);
xor U1901 (N_1901,In_407,In_2793);
nor U1902 (N_1902,In_2352,In_703);
nor U1903 (N_1903,In_4222,In_3839);
nand U1904 (N_1904,In_3963,In_4969);
or U1905 (N_1905,In_1009,In_2286);
or U1906 (N_1906,In_348,In_4498);
xor U1907 (N_1907,In_3017,In_808);
and U1908 (N_1908,In_1777,In_2616);
or U1909 (N_1909,In_4888,In_1838);
or U1910 (N_1910,In_3942,In_361);
nor U1911 (N_1911,In_4637,In_3790);
nor U1912 (N_1912,In_149,In_1490);
nor U1913 (N_1913,In_4807,In_2996);
nor U1914 (N_1914,In_1536,In_1125);
nand U1915 (N_1915,In_966,In_4576);
or U1916 (N_1916,In_4381,In_3831);
nand U1917 (N_1917,In_2429,In_2362);
nor U1918 (N_1918,In_525,In_664);
nand U1919 (N_1919,In_1410,In_3967);
or U1920 (N_1920,In_1429,In_2608);
nor U1921 (N_1921,In_2739,In_3787);
xor U1922 (N_1922,In_4990,In_2221);
nand U1923 (N_1923,In_2968,In_372);
nand U1924 (N_1924,In_4220,In_4047);
nor U1925 (N_1925,In_2647,In_1075);
or U1926 (N_1926,In_4951,In_4469);
nand U1927 (N_1927,In_1318,In_4179);
xor U1928 (N_1928,In_2919,In_4014);
or U1929 (N_1929,In_3491,In_3663);
and U1930 (N_1930,In_1210,In_2346);
nand U1931 (N_1931,In_2131,In_3369);
nor U1932 (N_1932,In_85,In_2026);
and U1933 (N_1933,In_2485,In_4299);
xor U1934 (N_1934,In_3502,In_322);
xor U1935 (N_1935,In_2343,In_4611);
nand U1936 (N_1936,In_1260,In_3608);
xnor U1937 (N_1937,In_1397,In_1958);
xnor U1938 (N_1938,In_297,In_4524);
and U1939 (N_1939,In_4884,In_801);
xnor U1940 (N_1940,In_4791,In_838);
xor U1941 (N_1941,In_467,In_3908);
nor U1942 (N_1942,In_2762,In_1239);
xnor U1943 (N_1943,In_3999,In_743);
and U1944 (N_1944,In_1783,In_4932);
nor U1945 (N_1945,In_2791,In_849);
nand U1946 (N_1946,In_4154,In_2134);
nand U1947 (N_1947,In_4011,In_279);
nand U1948 (N_1948,In_4939,In_3935);
xor U1949 (N_1949,In_3245,In_241);
nor U1950 (N_1950,In_1904,In_4771);
and U1951 (N_1951,In_124,In_4348);
and U1952 (N_1952,In_3701,In_586);
nand U1953 (N_1953,In_2746,In_556);
nor U1954 (N_1954,In_1161,In_215);
or U1955 (N_1955,In_423,In_3623);
nand U1956 (N_1956,In_4209,In_4703);
nor U1957 (N_1957,In_1820,In_648);
nand U1958 (N_1958,In_4292,In_1598);
nand U1959 (N_1959,In_1794,In_331);
xnor U1960 (N_1960,In_1727,In_2211);
nand U1961 (N_1961,In_4448,In_4123);
nor U1962 (N_1962,In_2263,In_3956);
and U1963 (N_1963,In_3118,In_432);
and U1964 (N_1964,In_1548,In_4735);
nand U1965 (N_1965,In_4444,In_2543);
xnor U1966 (N_1966,In_1454,In_259);
nand U1967 (N_1967,In_1253,In_1862);
xnor U1968 (N_1968,In_2735,In_3324);
nand U1969 (N_1969,In_2906,In_4031);
xor U1970 (N_1970,In_1087,In_1743);
xor U1971 (N_1971,In_1987,In_3386);
xor U1972 (N_1972,In_4012,In_1888);
nand U1973 (N_1973,In_3616,In_1517);
nor U1974 (N_1974,In_1941,In_4857);
and U1975 (N_1975,In_2564,In_4094);
and U1976 (N_1976,In_604,In_974);
xor U1977 (N_1977,In_2332,In_652);
and U1978 (N_1978,In_344,In_3516);
xnor U1979 (N_1979,In_3638,In_2261);
and U1980 (N_1980,In_1576,In_2655);
and U1981 (N_1981,In_1539,In_2031);
nand U1982 (N_1982,In_358,In_4790);
nand U1983 (N_1983,In_3848,In_4578);
nand U1984 (N_1984,In_4913,In_1405);
xor U1985 (N_1985,In_790,In_507);
xnor U1986 (N_1986,In_4648,In_2114);
and U1987 (N_1987,In_2361,In_4709);
and U1988 (N_1988,In_3974,In_1563);
or U1989 (N_1989,In_4543,In_47);
and U1990 (N_1990,In_4019,In_3883);
or U1991 (N_1991,In_506,In_3644);
xnor U1992 (N_1992,In_526,In_1469);
nor U1993 (N_1993,In_277,In_46);
nor U1994 (N_1994,In_3139,In_1463);
and U1995 (N_1995,In_1803,In_94);
and U1996 (N_1996,In_4541,In_3081);
nor U1997 (N_1997,In_3577,In_3878);
xor U1998 (N_1998,In_1772,In_4059);
and U1999 (N_1999,In_3475,In_1115);
nor U2000 (N_2000,In_287,In_1911);
and U2001 (N_2001,In_4434,In_367);
xor U2002 (N_2002,In_155,In_2143);
nand U2003 (N_2003,In_3814,In_1989);
and U2004 (N_2004,In_3977,In_4938);
or U2005 (N_2005,In_4517,In_1976);
and U2006 (N_2006,In_2765,In_2251);
or U2007 (N_2007,In_4804,In_1855);
nand U2008 (N_2008,In_783,In_3327);
and U2009 (N_2009,In_3533,In_4291);
or U2010 (N_2010,In_913,In_4925);
nand U2011 (N_2011,In_1586,In_3882);
and U2012 (N_2012,In_735,In_1809);
nor U2013 (N_2013,In_3031,In_2038);
and U2014 (N_2014,In_3357,In_1319);
xor U2015 (N_2015,In_3135,In_4656);
xor U2016 (N_2016,In_4412,In_572);
and U2017 (N_2017,In_175,In_447);
nor U2018 (N_2018,In_1814,In_4275);
nand U2019 (N_2019,In_4086,In_1471);
nor U2020 (N_2020,In_3655,In_2498);
and U2021 (N_2021,In_2696,In_4311);
xor U2022 (N_2022,In_3003,In_4653);
or U2023 (N_2023,In_1782,In_2911);
or U2024 (N_2024,In_1208,In_832);
or U2025 (N_2025,In_3612,In_413);
nand U2026 (N_2026,In_4116,In_2351);
or U2027 (N_2027,In_1706,In_3343);
xnor U2028 (N_2028,In_561,In_3580);
and U2029 (N_2029,In_1589,In_4192);
or U2030 (N_2030,In_4058,In_4500);
or U2031 (N_2031,In_3803,In_4262);
xnor U2032 (N_2032,In_1422,In_4040);
nor U2033 (N_2033,In_4189,In_4193);
and U2034 (N_2034,In_2341,In_2297);
nand U2035 (N_2035,In_333,In_2940);
xnor U2036 (N_2036,In_804,In_4946);
or U2037 (N_2037,In_3866,In_2734);
nor U2038 (N_2038,In_853,In_1451);
xor U2039 (N_2039,In_2946,In_613);
xor U2040 (N_2040,In_699,In_4984);
nand U2041 (N_2041,In_3600,In_2698);
nand U2042 (N_2042,In_1951,In_3296);
xnor U2043 (N_2043,In_997,In_1864);
or U2044 (N_2044,In_1339,In_1925);
nand U2045 (N_2045,In_3457,In_3943);
nand U2046 (N_2046,In_3680,In_3759);
and U2047 (N_2047,In_4258,In_2123);
nand U2048 (N_2048,In_1601,In_2728);
or U2049 (N_2049,In_2676,In_1144);
and U2050 (N_2050,In_504,In_2373);
nand U2051 (N_2051,In_4449,In_4322);
nor U2052 (N_2052,In_4402,In_1082);
nor U2053 (N_2053,In_583,In_922);
and U2054 (N_2054,In_52,In_1511);
and U2055 (N_2055,In_4632,In_1111);
nand U2056 (N_2056,In_153,In_1936);
xnor U2057 (N_2057,In_1618,In_3337);
and U2058 (N_2058,In_1863,In_4266);
nor U2059 (N_2059,In_3160,In_3544);
or U2060 (N_2060,In_1534,In_4535);
nand U2061 (N_2061,In_4315,In_2383);
or U2062 (N_2062,In_3096,In_4968);
xor U2063 (N_2063,In_1432,In_2815);
or U2064 (N_2064,In_3220,In_7);
or U2065 (N_2065,In_2250,In_1446);
and U2066 (N_2066,In_3539,In_4628);
or U2067 (N_2067,In_2817,In_2002);
and U2068 (N_2068,In_4514,In_3932);
or U2069 (N_2069,In_4794,In_2879);
xor U2070 (N_2070,In_15,In_1025);
and U2071 (N_2071,In_2032,In_2937);
and U2072 (N_2072,In_4324,In_1527);
nor U2073 (N_2073,In_1821,In_1333);
or U2074 (N_2074,In_3542,In_867);
and U2075 (N_2075,In_2646,In_4775);
xnor U2076 (N_2076,In_1130,In_2266);
and U2077 (N_2077,In_4659,In_4484);
xnor U2078 (N_2078,In_2471,In_3310);
nor U2079 (N_2079,In_2663,In_4479);
and U2080 (N_2080,In_2905,In_2132);
nand U2081 (N_2081,In_3736,In_1464);
and U2082 (N_2082,In_4948,In_4493);
nor U2083 (N_2083,In_4354,In_4403);
xnor U2084 (N_2084,In_4732,In_3466);
xnor U2085 (N_2085,In_3517,In_4674);
and U2086 (N_2086,In_2844,In_1089);
and U2087 (N_2087,In_4655,In_2553);
nor U2088 (N_2088,In_2888,In_3537);
nor U2089 (N_2089,In_4302,In_3841);
xor U2090 (N_2090,In_2907,In_742);
nand U2091 (N_2091,In_3352,In_4393);
xnor U2092 (N_2092,In_2097,In_2225);
or U2093 (N_2093,In_75,In_3407);
and U2094 (N_2094,In_1233,In_4679);
xor U2095 (N_2095,In_3292,In_508);
and U2096 (N_2096,In_4624,In_3620);
and U2097 (N_2097,In_3900,In_828);
or U2098 (N_2098,In_1909,In_3746);
nand U2099 (N_2099,In_2593,In_2093);
nand U2100 (N_2100,In_4757,In_2801);
xnor U2101 (N_2101,In_2863,In_3058);
or U2102 (N_2102,In_1566,In_4224);
nand U2103 (N_2103,In_339,In_2832);
and U2104 (N_2104,In_137,In_2086);
or U2105 (N_2105,In_3064,In_3812);
nor U2106 (N_2106,In_4729,In_4752);
and U2107 (N_2107,In_3097,In_2480);
nand U2108 (N_2108,In_4358,In_2540);
nand U2109 (N_2109,In_4836,In_2164);
or U2110 (N_2110,In_411,In_3699);
nand U2111 (N_2111,In_4006,In_2478);
xnor U2112 (N_2112,In_4931,In_3116);
nand U2113 (N_2113,In_1114,In_2913);
nand U2114 (N_2114,In_4478,In_2444);
nor U2115 (N_2115,In_1348,In_4949);
xor U2116 (N_2116,In_2150,In_4779);
nor U2117 (N_2117,In_4619,In_4506);
or U2118 (N_2118,In_497,In_40);
and U2119 (N_2119,In_570,In_1199);
or U2120 (N_2120,In_3383,In_2947);
xor U2121 (N_2121,In_3909,In_3321);
nand U2122 (N_2122,In_1033,In_3596);
and U2123 (N_2123,In_1581,In_1543);
nor U2124 (N_2124,In_1305,In_1655);
xor U2125 (N_2125,In_4298,In_3297);
nor U2126 (N_2126,In_2252,In_2228);
and U2127 (N_2127,In_4854,In_2446);
xnor U2128 (N_2128,In_3757,In_782);
and U2129 (N_2129,In_2055,In_4373);
xnor U2130 (N_2130,In_1209,In_1153);
xnor U2131 (N_2131,In_426,In_4013);
xor U2132 (N_2132,In_1165,In_3334);
xnor U2133 (N_2133,In_4751,In_752);
nand U2134 (N_2134,In_3730,In_3472);
and U2135 (N_2135,In_4190,In_3476);
xor U2136 (N_2136,In_872,In_3446);
nand U2137 (N_2137,In_901,In_2932);
or U2138 (N_2138,In_725,In_3554);
nor U2139 (N_2139,In_1221,In_154);
and U2140 (N_2140,In_2190,In_4378);
xnor U2141 (N_2141,In_1159,In_3870);
nand U2142 (N_2142,In_554,In_340);
or U2143 (N_2143,In_3403,In_885);
and U2144 (N_2144,In_2382,In_4466);
or U2145 (N_2145,In_2621,In_1502);
nor U2146 (N_2146,In_3273,In_2653);
nor U2147 (N_2147,In_4533,In_3484);
and U2148 (N_2148,In_3330,In_3784);
nor U2149 (N_2149,In_2507,In_2474);
or U2150 (N_2150,In_2839,In_4982);
xor U2151 (N_2151,In_2013,In_1182);
or U2152 (N_2152,In_4153,In_4080);
nor U2153 (N_2153,In_1582,In_321);
and U2154 (N_2154,In_757,In_3061);
nor U2155 (N_2155,In_434,In_2130);
xnor U2156 (N_2156,In_3060,In_4104);
and U2157 (N_2157,In_4698,In_3646);
nor U2158 (N_2158,In_935,In_2902);
or U2159 (N_2159,In_3887,In_1322);
nor U2160 (N_2160,In_4614,In_1020);
xor U2161 (N_2161,In_2963,In_1567);
nand U2162 (N_2162,In_2845,In_4295);
nor U2163 (N_2163,In_3391,In_2357);
nand U2164 (N_2164,In_4028,In_4228);
and U2165 (N_2165,In_4282,In_475);
nand U2166 (N_2166,In_4423,In_633);
and U2167 (N_2167,In_3152,In_2925);
or U2168 (N_2168,In_1547,In_345);
or U2169 (N_2169,In_4454,In_1966);
nor U2170 (N_2170,In_1923,In_1290);
nor U2171 (N_2171,In_3592,In_4724);
or U2172 (N_2172,In_803,In_3002);
nand U2173 (N_2173,In_3499,In_4555);
and U2174 (N_2174,In_491,In_4876);
nand U2175 (N_2175,In_2763,In_163);
nand U2176 (N_2176,In_1142,In_891);
nand U2177 (N_2177,In_1350,In_4092);
and U2178 (N_2178,In_1619,In_3507);
nor U2179 (N_2179,In_1441,In_224);
and U2180 (N_2180,In_2980,In_436);
and U2181 (N_2181,In_877,In_1874);
nand U2182 (N_2182,In_400,In_2315);
and U2183 (N_2183,In_3244,In_4832);
nor U2184 (N_2184,In_4245,In_4389);
or U2185 (N_2185,In_4630,In_1657);
nor U2186 (N_2186,In_4340,In_409);
or U2187 (N_2187,In_2729,In_2694);
nand U2188 (N_2188,In_3285,In_3722);
xor U2189 (N_2189,In_3318,In_1048);
or U2190 (N_2190,In_1556,In_2461);
nor U2191 (N_2191,In_2861,In_2102);
nor U2192 (N_2192,In_2424,In_4828);
or U2193 (N_2193,In_4043,In_4695);
xnor U2194 (N_2194,In_4269,In_3423);
and U2195 (N_2195,In_2479,In_1011);
nor U2196 (N_2196,In_56,In_3647);
or U2197 (N_2197,In_1731,In_3618);
xor U2198 (N_2198,In_249,In_1779);
nand U2199 (N_2199,In_1602,In_3201);
nand U2200 (N_2200,In_450,In_3936);
nor U2201 (N_2201,In_609,In_4699);
nand U2202 (N_2202,In_1676,In_3636);
or U2203 (N_2203,In_3040,In_6);
nand U2204 (N_2204,In_2219,In_4858);
or U2205 (N_2205,In_2014,In_4501);
xor U2206 (N_2206,In_4997,In_4138);
and U2207 (N_2207,In_2692,In_4915);
nor U2208 (N_2208,In_635,In_4979);
or U2209 (N_2209,In_3519,In_305);
nand U2210 (N_2210,In_3458,In_3208);
xnor U2211 (N_2211,In_3683,In_2456);
nor U2212 (N_2212,In_3931,In_2183);
or U2213 (N_2213,In_2230,In_213);
nor U2214 (N_2214,In_4644,In_2389);
nor U2215 (N_2215,In_4808,In_2348);
nand U2216 (N_2216,In_23,In_4581);
and U2217 (N_2217,In_480,In_4551);
or U2218 (N_2218,In_2812,In_4336);
and U2219 (N_2219,In_1196,In_4521);
and U2220 (N_2220,In_1499,In_2335);
or U2221 (N_2221,In_1639,In_1785);
and U2222 (N_2222,In_354,In_629);
xor U2223 (N_2223,In_4670,In_4785);
nand U2224 (N_2224,In_1656,In_665);
nand U2225 (N_2225,In_183,In_2513);
or U2226 (N_2226,In_754,In_1364);
and U2227 (N_2227,In_874,In_2995);
xnor U2228 (N_2228,In_1795,In_940);
and U2229 (N_2229,In_729,In_1886);
and U2230 (N_2230,In_95,In_969);
nor U2231 (N_2231,In_3103,In_649);
xor U2232 (N_2232,In_3772,In_2950);
nand U2233 (N_2233,In_2156,In_1572);
nor U2234 (N_2234,In_1477,In_3495);
and U2235 (N_2235,In_1250,In_3188);
xor U2236 (N_2236,In_3885,In_1118);
and U2237 (N_2237,In_2960,In_2028);
or U2238 (N_2238,In_3049,In_3136);
nor U2239 (N_2239,In_4610,In_3196);
and U2240 (N_2240,In_2555,In_2386);
and U2241 (N_2241,In_2682,In_1340);
nand U2242 (N_2242,In_3518,In_510);
xor U2243 (N_2243,In_254,In_1603);
and U2244 (N_2244,In_3037,In_2679);
nand U2245 (N_2245,In_4409,In_2255);
nor U2246 (N_2246,In_919,In_1170);
xnor U2247 (N_2247,In_1521,In_1068);
nor U2248 (N_2248,In_3157,In_2223);
nand U2249 (N_2249,In_1370,In_2020);
xor U2250 (N_2250,In_50,In_3976);
or U2251 (N_2251,In_3630,In_4993);
or U2252 (N_2252,In_843,In_3745);
xor U2253 (N_2253,In_337,In_4889);
nor U2254 (N_2254,In_3490,In_1401);
and U2255 (N_2255,In_470,In_1373);
nor U2256 (N_2256,In_4177,In_4157);
xor U2257 (N_2257,In_3072,In_3223);
nor U2258 (N_2258,In_3536,In_3564);
xnor U2259 (N_2259,In_640,In_4426);
xor U2260 (N_2260,In_2338,In_3649);
nand U2261 (N_2261,In_4066,In_2807);
or U2262 (N_2262,In_1919,In_3569);
nor U2263 (N_2263,In_1701,In_3230);
or U2264 (N_2264,In_3633,In_632);
nand U2265 (N_2265,In_4406,In_2965);
or U2266 (N_2266,In_2858,In_3168);
and U2267 (N_2267,In_1281,In_1516);
and U2268 (N_2268,In_1015,In_3818);
nor U2269 (N_2269,In_2685,In_2298);
and U2270 (N_2270,In_3560,In_2639);
xnor U2271 (N_2271,In_4356,In_1180);
nand U2272 (N_2272,In_1927,In_3833);
or U2273 (N_2273,In_1762,In_1047);
nand U2274 (N_2274,In_2388,In_978);
nor U2275 (N_2275,In_3447,In_4362);
xor U2276 (N_2276,In_1447,In_4413);
and U2277 (N_2277,In_1284,In_4272);
and U2278 (N_2278,In_1246,In_1264);
and U2279 (N_2279,In_947,In_4545);
or U2280 (N_2280,In_692,In_946);
nand U2281 (N_2281,In_948,In_2385);
and U2282 (N_2282,In_1716,In_476);
nand U2283 (N_2283,In_1939,In_3260);
xnor U2284 (N_2284,In_3609,In_2645);
nand U2285 (N_2285,In_3892,In_2533);
xor U2286 (N_2286,In_4607,In_746);
and U2287 (N_2287,In_2634,In_1249);
or U2288 (N_2288,In_2313,In_3869);
and U2289 (N_2289,In_4713,In_383);
xnor U2290 (N_2290,In_4776,In_2983);
nand U2291 (N_2291,In_1746,In_4678);
xor U2292 (N_2292,In_4923,In_160);
and U2293 (N_2293,In_2705,In_1202);
and U2294 (N_2294,In_3054,In_1760);
or U2295 (N_2295,In_3381,In_1865);
xor U2296 (N_2296,In_406,In_2046);
or U2297 (N_2297,In_4321,In_1990);
xnor U2298 (N_2298,In_4903,In_1648);
nor U2299 (N_2299,In_3341,In_1313);
nor U2300 (N_2300,In_4213,In_2193);
and U2301 (N_2301,In_257,In_1781);
and U2302 (N_2302,In_3175,In_2973);
or U2303 (N_2303,In_831,In_3237);
xnor U2304 (N_2304,In_4561,In_1254);
nor U2305 (N_2305,In_4325,In_173);
xnor U2306 (N_2306,In_4813,In_3010);
xor U2307 (N_2307,In_4762,In_3351);
and U2308 (N_2308,In_30,In_1440);
or U2309 (N_2309,In_2064,In_3364);
and U2310 (N_2310,In_3879,In_482);
nand U2311 (N_2311,In_4867,In_4651);
nor U2312 (N_2312,In_1915,In_873);
nor U2313 (N_2313,In_107,In_2326);
or U2314 (N_2314,In_3944,In_2124);
or U2315 (N_2315,In_146,In_1876);
nand U2316 (N_2316,In_3922,In_2556);
nand U2317 (N_2317,In_1658,In_3850);
nand U2318 (N_2318,In_2976,In_2310);
nor U2319 (N_2319,In_3409,In_1309);
xnor U2320 (N_2320,In_4480,In_3229);
nor U2321 (N_2321,In_3225,In_3547);
or U2322 (N_2322,In_4439,In_2455);
and U2323 (N_2323,In_4173,In_4835);
and U2324 (N_2324,In_3555,In_3629);
nor U2325 (N_2325,In_1045,In_1474);
xnor U2326 (N_2326,In_2865,In_993);
or U2327 (N_2327,In_1225,In_4186);
nand U2328 (N_2328,In_1384,In_4281);
xnor U2329 (N_2329,In_3723,In_4497);
or U2330 (N_2330,In_1194,In_2535);
nand U2331 (N_2331,In_3822,In_2700);
nand U2332 (N_2332,In_2421,In_4529);
xor U2333 (N_2333,In_1740,In_1674);
nand U2334 (N_2334,In_2307,In_3170);
nand U2335 (N_2335,In_3108,In_991);
or U2336 (N_2336,In_3071,In_964);
nand U2337 (N_2337,In_2324,In_431);
or U2338 (N_2338,In_4353,In_2898);
xor U2339 (N_2339,In_184,In_4411);
xnor U2340 (N_2340,In_364,In_4746);
or U2341 (N_2341,In_4918,In_4396);
and U2342 (N_2342,In_4748,In_4726);
nor U2343 (N_2343,In_4468,In_4827);
and U2344 (N_2344,In_3824,In_4685);
nand U2345 (N_2345,In_642,In_3365);
xnor U2346 (N_2346,In_1167,In_2675);
or U2347 (N_2347,In_4496,In_3249);
nor U2348 (N_2348,In_4780,In_3823);
xor U2349 (N_2349,In_761,In_4198);
or U2350 (N_2350,In_2690,In_2622);
or U2351 (N_2351,In_4251,In_863);
xnor U2352 (N_2352,In_1824,In_3400);
xnor U2353 (N_2353,In_1616,In_4792);
nand U2354 (N_2354,In_272,In_4410);
nand U2355 (N_2355,In_899,In_573);
or U2356 (N_2356,In_4542,In_4473);
and U2357 (N_2357,In_1579,In_4840);
and U2358 (N_2358,In_4604,In_3091);
nand U2359 (N_2359,In_1770,In_929);
nand U2360 (N_2360,In_262,In_4538);
nand U2361 (N_2361,In_3525,In_3016);
or U2362 (N_2362,In_122,In_2681);
nor U2363 (N_2363,In_2699,In_211);
xnor U2364 (N_2364,In_2612,In_3328);
or U2365 (N_2365,In_4618,In_1767);
or U2366 (N_2366,In_240,In_1388);
and U2367 (N_2367,In_2810,In_1807);
and U2368 (N_2368,In_2381,In_1882);
nor U2369 (N_2369,In_2224,In_2526);
xor U2370 (N_2370,In_4935,In_1959);
nor U2371 (N_2371,In_641,In_1545);
and U2372 (N_2372,In_2145,In_1631);
nor U2373 (N_2373,In_4229,In_3756);
or U2374 (N_2374,In_264,In_505);
nor U2375 (N_2375,In_1956,In_2441);
or U2376 (N_2376,In_1873,In_2693);
nand U2377 (N_2377,In_775,In_600);
or U2378 (N_2378,In_3319,In_1922);
and U2379 (N_2379,In_715,In_390);
or U2380 (N_2380,In_1789,In_1444);
nand U2381 (N_2381,In_13,In_1954);
xnor U2382 (N_2382,In_21,In_2978);
nor U2383 (N_2383,In_4453,In_1395);
nor U2384 (N_2384,In_4536,In_4826);
nor U2385 (N_2385,In_4065,In_3454);
nor U2386 (N_2386,In_4372,In_2525);
xor U2387 (N_2387,In_4873,In_24);
nand U2388 (N_2388,In_718,In_1933);
xor U2389 (N_2389,In_1668,In_135);
or U2390 (N_2390,In_3717,In_1512);
and U2391 (N_2391,In_1053,In_3322);
nor U2392 (N_2392,In_4546,In_1123);
nand U2393 (N_2393,In_152,In_2495);
nor U2394 (N_2394,In_1916,In_4073);
nand U2395 (N_2395,In_4647,In_2072);
nor U2396 (N_2396,In_1078,In_323);
nand U2397 (N_2397,In_4806,In_1627);
nand U2398 (N_2398,In_2756,In_2254);
nor U2399 (N_2399,In_1771,In_992);
nand U2400 (N_2400,In_2856,In_2695);
nor U2401 (N_2401,In_1663,In_3751);
nor U2402 (N_2402,In_4640,In_1218);
nor U2403 (N_2403,In_2437,In_659);
or U2404 (N_2404,In_2954,In_3434);
xor U2405 (N_2405,In_4370,In_3422);
nand U2406 (N_2406,In_3926,In_543);
nand U2407 (N_2407,In_3395,In_1891);
nor U2408 (N_2408,In_1859,In_2959);
xor U2409 (N_2409,In_3426,In_4571);
xnor U2410 (N_2410,In_3367,In_2413);
nor U2411 (N_2411,In_4749,In_4878);
and U2412 (N_2412,In_4825,In_1090);
xor U2413 (N_2413,In_3036,In_2340);
nand U2414 (N_2414,In_3247,In_127);
or U2415 (N_2415,In_209,In_2015);
nor U2416 (N_2416,In_3358,In_712);
and U2417 (N_2417,In_1969,In_1717);
and U2418 (N_2418,In_766,In_1861);
xor U2419 (N_2419,In_2010,In_266);
or U2420 (N_2420,In_1439,In_3311);
nand U2421 (N_2421,In_2439,In_1071);
and U2422 (N_2422,In_4081,In_4166);
nor U2423 (N_2423,In_1596,In_1823);
xor U2424 (N_2424,In_121,In_2736);
nand U2425 (N_2425,In_351,In_2459);
xnor U2426 (N_2426,In_3068,In_2640);
nand U2427 (N_2427,In_1101,In_1897);
nand U2428 (N_2428,In_1775,In_2023);
xnor U2429 (N_2429,In_1343,In_43);
nand U2430 (N_2430,In_4958,In_204);
nand U2431 (N_2431,In_3523,In_4973);
or U2432 (N_2432,In_1351,In_2005);
nand U2433 (N_2433,In_1878,In_737);
nand U2434 (N_2434,In_1568,In_2375);
or U2435 (N_2435,In_3558,In_4380);
nor U2436 (N_2436,In_4741,In_2506);
nand U2437 (N_2437,In_971,In_300);
and U2438 (N_2438,In_3481,In_923);
and U2439 (N_2439,In_3489,In_101);
nand U2440 (N_2440,In_3219,In_1042);
and U2441 (N_2441,In_4140,In_4976);
or U2442 (N_2442,In_1195,In_2575);
xor U2443 (N_2443,In_2585,In_2045);
nor U2444 (N_2444,In_395,In_2033);
nor U2445 (N_2445,In_3732,In_3062);
nor U2446 (N_2446,In_3282,In_1001);
nor U2447 (N_2447,In_1187,In_2486);
nand U2448 (N_2448,In_3918,In_118);
nand U2449 (N_2449,In_468,In_2722);
and U2450 (N_2450,In_1750,In_49);
xnor U2451 (N_2451,In_2781,In_4146);
or U2452 (N_2452,In_4575,In_4676);
nand U2453 (N_2453,In_2174,In_4489);
and U2454 (N_2454,In_2770,In_3867);
nor U2455 (N_2455,In_59,In_3266);
nor U2456 (N_2456,In_1853,In_1057);
xor U2457 (N_2457,In_2133,In_1106);
or U2458 (N_2458,In_2317,In_349);
nor U2459 (N_2459,In_2182,In_4064);
nand U2460 (N_2460,In_1714,In_962);
xor U2461 (N_2461,In_4329,In_868);
and U2462 (N_2462,In_631,In_4304);
nor U2463 (N_2463,In_2443,In_2079);
and U2464 (N_2464,In_2329,In_486);
nand U2465 (N_2465,In_1526,In_133);
nor U2466 (N_2466,In_2782,In_893);
nand U2467 (N_2467,In_965,In_802);
xor U2468 (N_2468,In_2574,In_3066);
or U2469 (N_2469,In_3312,In_4681);
and U2470 (N_2470,In_1755,In_2127);
nand U2471 (N_2471,In_4970,In_1267);
and U2472 (N_2472,In_2451,In_3624);
nor U2473 (N_2473,In_2300,In_3295);
nand U2474 (N_2474,In_246,In_2975);
or U2475 (N_2475,In_2099,In_4626);
nand U2476 (N_2476,In_1175,In_1148);
nor U2477 (N_2477,In_4169,In_4366);
and U2478 (N_2478,In_905,In_4176);
nor U2479 (N_2479,In_1409,In_2202);
and U2480 (N_2480,In_1980,In_3095);
xor U2481 (N_2481,In_695,In_800);
or U2482 (N_2482,In_4821,In_1345);
and U2483 (N_2483,In_78,In_1146);
xnor U2484 (N_2484,In_496,In_4247);
nor U2485 (N_2485,In_1721,In_1883);
xnor U2486 (N_2486,In_207,In_4240);
and U2487 (N_2487,In_3050,In_4001);
nor U2488 (N_2488,In_4139,In_626);
or U2489 (N_2489,In_2006,In_1945);
and U2490 (N_2490,In_2922,In_2958);
and U2491 (N_2491,In_1972,In_1510);
nor U2492 (N_2492,In_2943,In_942);
and U2493 (N_2493,In_2070,In_780);
nand U2494 (N_2494,In_4392,In_2624);
nand U2495 (N_2495,In_745,In_4584);
xor U2496 (N_2496,In_51,In_3289);
or U2497 (N_2497,In_4133,In_379);
nor U2498 (N_2498,In_3019,In_4215);
nor U2499 (N_2499,In_4458,In_3795);
nor U2500 (N_2500,In_2704,In_3214);
and U2501 (N_2501,In_2048,In_1819);
nand U2502 (N_2502,In_2899,In_2786);
or U2503 (N_2503,In_2849,In_4865);
and U2504 (N_2504,In_4342,In_2567);
xor U2505 (N_2505,In_1021,In_3008);
or U2506 (N_2506,In_2163,In_4410);
or U2507 (N_2507,In_4169,In_2302);
or U2508 (N_2508,In_3780,In_4646);
and U2509 (N_2509,In_2341,In_4879);
or U2510 (N_2510,In_2449,In_2330);
xnor U2511 (N_2511,In_3339,In_4204);
nand U2512 (N_2512,In_3343,In_973);
nor U2513 (N_2513,In_1642,In_2605);
xor U2514 (N_2514,In_3615,In_4541);
or U2515 (N_2515,In_877,In_1983);
nand U2516 (N_2516,In_3891,In_1688);
nand U2517 (N_2517,In_3037,In_4978);
and U2518 (N_2518,In_2653,In_44);
xor U2519 (N_2519,In_561,In_2081);
nor U2520 (N_2520,In_681,In_3941);
and U2521 (N_2521,In_4982,In_4261);
nand U2522 (N_2522,In_4528,In_3234);
xnor U2523 (N_2523,In_1273,In_309);
or U2524 (N_2524,In_2183,In_422);
nand U2525 (N_2525,In_4608,In_3449);
and U2526 (N_2526,In_4436,In_4602);
nand U2527 (N_2527,In_4481,In_2324);
nand U2528 (N_2528,In_2322,In_3767);
nand U2529 (N_2529,In_340,In_2825);
nand U2530 (N_2530,In_4622,In_2123);
nand U2531 (N_2531,In_478,In_3099);
and U2532 (N_2532,In_4677,In_1652);
nor U2533 (N_2533,In_4721,In_4743);
nor U2534 (N_2534,In_2919,In_2621);
or U2535 (N_2535,In_1230,In_4528);
nand U2536 (N_2536,In_4208,In_2799);
or U2537 (N_2537,In_2248,In_255);
or U2538 (N_2538,In_3442,In_3066);
or U2539 (N_2539,In_1773,In_4881);
xor U2540 (N_2540,In_155,In_4550);
or U2541 (N_2541,In_4980,In_4002);
or U2542 (N_2542,In_4441,In_4569);
nor U2543 (N_2543,In_1478,In_2684);
nand U2544 (N_2544,In_1383,In_3575);
xnor U2545 (N_2545,In_4454,In_3606);
xnor U2546 (N_2546,In_2064,In_3529);
and U2547 (N_2547,In_3216,In_209);
nor U2548 (N_2548,In_1420,In_307);
or U2549 (N_2549,In_1867,In_4764);
nor U2550 (N_2550,In_575,In_1136);
nand U2551 (N_2551,In_2954,In_1795);
or U2552 (N_2552,In_3064,In_4339);
nand U2553 (N_2553,In_4732,In_3951);
and U2554 (N_2554,In_2866,In_2209);
or U2555 (N_2555,In_2167,In_2156);
nand U2556 (N_2556,In_174,In_703);
xnor U2557 (N_2557,In_4607,In_4308);
nand U2558 (N_2558,In_3473,In_4163);
nor U2559 (N_2559,In_3078,In_2686);
or U2560 (N_2560,In_4295,In_3424);
xor U2561 (N_2561,In_819,In_1107);
xor U2562 (N_2562,In_1341,In_4565);
xor U2563 (N_2563,In_2364,In_1704);
xnor U2564 (N_2564,In_2083,In_1657);
xor U2565 (N_2565,In_4837,In_4478);
xor U2566 (N_2566,In_1592,In_2739);
or U2567 (N_2567,In_1269,In_2950);
and U2568 (N_2568,In_2257,In_2573);
nor U2569 (N_2569,In_2801,In_244);
or U2570 (N_2570,In_2654,In_1443);
nor U2571 (N_2571,In_784,In_4774);
xor U2572 (N_2572,In_2639,In_4911);
xor U2573 (N_2573,In_2200,In_1918);
and U2574 (N_2574,In_4818,In_1521);
nand U2575 (N_2575,In_1597,In_3276);
xor U2576 (N_2576,In_4048,In_219);
xnor U2577 (N_2577,In_3840,In_4177);
nor U2578 (N_2578,In_604,In_1769);
and U2579 (N_2579,In_4259,In_792);
nor U2580 (N_2580,In_3604,In_1578);
or U2581 (N_2581,In_2968,In_4604);
or U2582 (N_2582,In_2495,In_1270);
and U2583 (N_2583,In_4641,In_3469);
nand U2584 (N_2584,In_1080,In_2705);
nand U2585 (N_2585,In_3923,In_4755);
nor U2586 (N_2586,In_276,In_26);
xnor U2587 (N_2587,In_523,In_4820);
and U2588 (N_2588,In_4703,In_3251);
or U2589 (N_2589,In_3288,In_1248);
nand U2590 (N_2590,In_4007,In_1772);
nand U2591 (N_2591,In_1946,In_353);
and U2592 (N_2592,In_4020,In_3466);
xnor U2593 (N_2593,In_3839,In_2952);
and U2594 (N_2594,In_4005,In_1538);
nor U2595 (N_2595,In_3333,In_4741);
nand U2596 (N_2596,In_2081,In_3082);
nor U2597 (N_2597,In_198,In_1088);
or U2598 (N_2598,In_3973,In_371);
and U2599 (N_2599,In_4060,In_987);
or U2600 (N_2600,In_1462,In_4273);
and U2601 (N_2601,In_3169,In_4370);
nand U2602 (N_2602,In_3825,In_3426);
xor U2603 (N_2603,In_1586,In_2756);
nand U2604 (N_2604,In_301,In_3694);
nand U2605 (N_2605,In_289,In_3958);
nand U2606 (N_2606,In_3172,In_197);
or U2607 (N_2607,In_627,In_1507);
nor U2608 (N_2608,In_3467,In_3035);
or U2609 (N_2609,In_623,In_3085);
and U2610 (N_2610,In_2758,In_4966);
xnor U2611 (N_2611,In_4468,In_2139);
nor U2612 (N_2612,In_2585,In_2909);
nor U2613 (N_2613,In_3299,In_1054);
and U2614 (N_2614,In_4637,In_3719);
and U2615 (N_2615,In_3641,In_1654);
or U2616 (N_2616,In_2127,In_1378);
xor U2617 (N_2617,In_2750,In_3471);
or U2618 (N_2618,In_2653,In_640);
nand U2619 (N_2619,In_4239,In_164);
nand U2620 (N_2620,In_2248,In_3547);
xor U2621 (N_2621,In_3430,In_2044);
or U2622 (N_2622,In_4640,In_2013);
xnor U2623 (N_2623,In_1222,In_4508);
and U2624 (N_2624,In_2769,In_2827);
or U2625 (N_2625,In_1725,In_2582);
nand U2626 (N_2626,In_2571,In_1605);
nor U2627 (N_2627,In_4717,In_246);
xor U2628 (N_2628,In_1624,In_809);
nand U2629 (N_2629,In_3698,In_1897);
nor U2630 (N_2630,In_4908,In_210);
xnor U2631 (N_2631,In_4670,In_3197);
nor U2632 (N_2632,In_2346,In_3097);
nor U2633 (N_2633,In_1900,In_3760);
nand U2634 (N_2634,In_233,In_601);
and U2635 (N_2635,In_4796,In_1804);
xnor U2636 (N_2636,In_4222,In_1104);
xnor U2637 (N_2637,In_2662,In_646);
and U2638 (N_2638,In_1817,In_1886);
and U2639 (N_2639,In_2436,In_4338);
and U2640 (N_2640,In_2058,In_2349);
xor U2641 (N_2641,In_2399,In_4851);
or U2642 (N_2642,In_4983,In_1945);
and U2643 (N_2643,In_1760,In_1797);
or U2644 (N_2644,In_4508,In_2860);
nand U2645 (N_2645,In_3395,In_3342);
xnor U2646 (N_2646,In_3601,In_1710);
or U2647 (N_2647,In_4805,In_2366);
or U2648 (N_2648,In_2365,In_2802);
nor U2649 (N_2649,In_2218,In_3651);
nor U2650 (N_2650,In_2223,In_3131);
and U2651 (N_2651,In_1916,In_3590);
and U2652 (N_2652,In_3239,In_780);
xnor U2653 (N_2653,In_692,In_235);
nor U2654 (N_2654,In_4415,In_4197);
xor U2655 (N_2655,In_3239,In_613);
nand U2656 (N_2656,In_96,In_1859);
and U2657 (N_2657,In_3414,In_2858);
and U2658 (N_2658,In_3060,In_1468);
nor U2659 (N_2659,In_2048,In_143);
and U2660 (N_2660,In_282,In_3718);
xor U2661 (N_2661,In_2389,In_1673);
or U2662 (N_2662,In_2690,In_2332);
or U2663 (N_2663,In_2104,In_4261);
and U2664 (N_2664,In_4328,In_281);
nand U2665 (N_2665,In_2704,In_3655);
or U2666 (N_2666,In_1274,In_3452);
and U2667 (N_2667,In_596,In_4456);
xnor U2668 (N_2668,In_3088,In_1417);
xor U2669 (N_2669,In_912,In_4017);
nand U2670 (N_2670,In_3420,In_8);
xor U2671 (N_2671,In_3301,In_2678);
nor U2672 (N_2672,In_281,In_2729);
nor U2673 (N_2673,In_525,In_1796);
or U2674 (N_2674,In_2304,In_3953);
and U2675 (N_2675,In_4274,In_22);
or U2676 (N_2676,In_1936,In_989);
nand U2677 (N_2677,In_97,In_3855);
and U2678 (N_2678,In_1369,In_3149);
nor U2679 (N_2679,In_3585,In_3670);
and U2680 (N_2680,In_221,In_2823);
or U2681 (N_2681,In_4412,In_3114);
nor U2682 (N_2682,In_3208,In_1160);
and U2683 (N_2683,In_512,In_748);
and U2684 (N_2684,In_2680,In_777);
and U2685 (N_2685,In_1789,In_310);
and U2686 (N_2686,In_883,In_4203);
nor U2687 (N_2687,In_2066,In_3157);
nand U2688 (N_2688,In_1189,In_1038);
nand U2689 (N_2689,In_2520,In_793);
and U2690 (N_2690,In_4578,In_4079);
nand U2691 (N_2691,In_1472,In_2748);
nand U2692 (N_2692,In_3684,In_3711);
or U2693 (N_2693,In_4725,In_1424);
or U2694 (N_2694,In_4118,In_582);
nand U2695 (N_2695,In_3041,In_3605);
or U2696 (N_2696,In_1270,In_2352);
nand U2697 (N_2697,In_143,In_835);
xor U2698 (N_2698,In_1628,In_2972);
nor U2699 (N_2699,In_2272,In_1574);
nand U2700 (N_2700,In_3788,In_1148);
xor U2701 (N_2701,In_3213,In_3628);
and U2702 (N_2702,In_4912,In_888);
xor U2703 (N_2703,In_3607,In_242);
nor U2704 (N_2704,In_1459,In_3455);
nand U2705 (N_2705,In_1314,In_980);
or U2706 (N_2706,In_3523,In_4240);
or U2707 (N_2707,In_3718,In_3113);
xnor U2708 (N_2708,In_1768,In_1718);
nand U2709 (N_2709,In_4884,In_4940);
xnor U2710 (N_2710,In_3177,In_1153);
nor U2711 (N_2711,In_2805,In_2727);
nor U2712 (N_2712,In_3383,In_2839);
nor U2713 (N_2713,In_2898,In_4513);
xor U2714 (N_2714,In_695,In_776);
nor U2715 (N_2715,In_3851,In_3980);
or U2716 (N_2716,In_2949,In_38);
xor U2717 (N_2717,In_3025,In_565);
nor U2718 (N_2718,In_4595,In_287);
nand U2719 (N_2719,In_4096,In_2370);
or U2720 (N_2720,In_4816,In_539);
and U2721 (N_2721,In_693,In_684);
and U2722 (N_2722,In_823,In_136);
or U2723 (N_2723,In_4717,In_126);
nand U2724 (N_2724,In_1399,In_1355);
nand U2725 (N_2725,In_878,In_4187);
xnor U2726 (N_2726,In_1551,In_893);
nor U2727 (N_2727,In_4863,In_3021);
and U2728 (N_2728,In_2225,In_2231);
nor U2729 (N_2729,In_2513,In_1732);
nor U2730 (N_2730,In_1989,In_4637);
nand U2731 (N_2731,In_3555,In_848);
xnor U2732 (N_2732,In_3118,In_4794);
nand U2733 (N_2733,In_4432,In_1479);
nand U2734 (N_2734,In_2930,In_2233);
xnor U2735 (N_2735,In_3881,In_3669);
or U2736 (N_2736,In_2066,In_1867);
nor U2737 (N_2737,In_1989,In_3611);
nor U2738 (N_2738,In_4217,In_2543);
and U2739 (N_2739,In_374,In_1844);
nor U2740 (N_2740,In_2910,In_1182);
nor U2741 (N_2741,In_2180,In_814);
or U2742 (N_2742,In_4344,In_188);
nand U2743 (N_2743,In_2185,In_1989);
nor U2744 (N_2744,In_4625,In_1123);
nor U2745 (N_2745,In_4963,In_887);
nor U2746 (N_2746,In_1918,In_4210);
nor U2747 (N_2747,In_4409,In_2559);
nand U2748 (N_2748,In_848,In_2237);
nor U2749 (N_2749,In_2642,In_4218);
nor U2750 (N_2750,In_4322,In_1708);
nand U2751 (N_2751,In_2905,In_4618);
nand U2752 (N_2752,In_95,In_4881);
nor U2753 (N_2753,In_2639,In_3666);
xor U2754 (N_2754,In_2357,In_514);
xor U2755 (N_2755,In_4001,In_2584);
nor U2756 (N_2756,In_431,In_3756);
and U2757 (N_2757,In_4719,In_1433);
or U2758 (N_2758,In_524,In_573);
nor U2759 (N_2759,In_4154,In_3105);
nor U2760 (N_2760,In_600,In_3252);
or U2761 (N_2761,In_2732,In_900);
nor U2762 (N_2762,In_1229,In_3602);
xnor U2763 (N_2763,In_3425,In_2333);
and U2764 (N_2764,In_2971,In_464);
nand U2765 (N_2765,In_1679,In_4809);
nand U2766 (N_2766,In_2310,In_1105);
xnor U2767 (N_2767,In_1537,In_2985);
and U2768 (N_2768,In_4255,In_1105);
and U2769 (N_2769,In_307,In_1135);
or U2770 (N_2770,In_2011,In_538);
or U2771 (N_2771,In_2480,In_4619);
or U2772 (N_2772,In_1623,In_1884);
or U2773 (N_2773,In_4607,In_944);
nand U2774 (N_2774,In_2902,In_3156);
nand U2775 (N_2775,In_1127,In_803);
and U2776 (N_2776,In_243,In_3110);
and U2777 (N_2777,In_4551,In_1091);
xor U2778 (N_2778,In_2782,In_4958);
or U2779 (N_2779,In_3625,In_2309);
and U2780 (N_2780,In_4718,In_1759);
nor U2781 (N_2781,In_2328,In_4295);
and U2782 (N_2782,In_2623,In_782);
xor U2783 (N_2783,In_1988,In_2487);
nor U2784 (N_2784,In_2418,In_4791);
or U2785 (N_2785,In_4522,In_641);
nor U2786 (N_2786,In_1293,In_3659);
and U2787 (N_2787,In_2591,In_1231);
nand U2788 (N_2788,In_781,In_339);
nor U2789 (N_2789,In_1560,In_3721);
nand U2790 (N_2790,In_3645,In_2686);
and U2791 (N_2791,In_490,In_115);
and U2792 (N_2792,In_2816,In_4911);
or U2793 (N_2793,In_2959,In_2111);
nor U2794 (N_2794,In_3759,In_4131);
and U2795 (N_2795,In_2989,In_3892);
xnor U2796 (N_2796,In_73,In_4146);
nor U2797 (N_2797,In_490,In_587);
nand U2798 (N_2798,In_2628,In_2113);
or U2799 (N_2799,In_2113,In_3141);
nand U2800 (N_2800,In_4083,In_2529);
nor U2801 (N_2801,In_1466,In_1670);
or U2802 (N_2802,In_2309,In_2311);
nand U2803 (N_2803,In_4524,In_4650);
xnor U2804 (N_2804,In_838,In_351);
nand U2805 (N_2805,In_4953,In_3947);
or U2806 (N_2806,In_4117,In_77);
xnor U2807 (N_2807,In_1159,In_602);
or U2808 (N_2808,In_518,In_683);
nor U2809 (N_2809,In_349,In_887);
and U2810 (N_2810,In_4432,In_2803);
xor U2811 (N_2811,In_1383,In_2906);
or U2812 (N_2812,In_2165,In_93);
or U2813 (N_2813,In_966,In_4265);
or U2814 (N_2814,In_333,In_4693);
or U2815 (N_2815,In_2709,In_3529);
nor U2816 (N_2816,In_2523,In_2706);
xor U2817 (N_2817,In_3825,In_1349);
or U2818 (N_2818,In_3944,In_1677);
or U2819 (N_2819,In_825,In_51);
and U2820 (N_2820,In_618,In_1176);
xor U2821 (N_2821,In_4335,In_4647);
xnor U2822 (N_2822,In_2903,In_3977);
nor U2823 (N_2823,In_1807,In_2730);
xnor U2824 (N_2824,In_3434,In_2116);
nor U2825 (N_2825,In_2543,In_3056);
xor U2826 (N_2826,In_2851,In_766);
or U2827 (N_2827,In_2905,In_3754);
xor U2828 (N_2828,In_3186,In_1729);
and U2829 (N_2829,In_1856,In_4875);
nor U2830 (N_2830,In_406,In_1694);
xor U2831 (N_2831,In_2338,In_965);
nand U2832 (N_2832,In_4390,In_191);
nand U2833 (N_2833,In_836,In_1813);
nor U2834 (N_2834,In_877,In_837);
nand U2835 (N_2835,In_4519,In_858);
xnor U2836 (N_2836,In_3709,In_623);
and U2837 (N_2837,In_3230,In_2518);
nand U2838 (N_2838,In_1269,In_3458);
and U2839 (N_2839,In_3987,In_4048);
xnor U2840 (N_2840,In_3960,In_2888);
or U2841 (N_2841,In_130,In_1926);
xor U2842 (N_2842,In_3263,In_2986);
nand U2843 (N_2843,In_811,In_1177);
or U2844 (N_2844,In_3674,In_709);
nor U2845 (N_2845,In_2644,In_3478);
xnor U2846 (N_2846,In_3163,In_4177);
nor U2847 (N_2847,In_3386,In_819);
or U2848 (N_2848,In_4595,In_638);
nand U2849 (N_2849,In_80,In_3768);
and U2850 (N_2850,In_4766,In_1104);
or U2851 (N_2851,In_2815,In_3942);
nand U2852 (N_2852,In_2099,In_4844);
nor U2853 (N_2853,In_3799,In_4858);
or U2854 (N_2854,In_2557,In_111);
nor U2855 (N_2855,In_22,In_2320);
xnor U2856 (N_2856,In_1345,In_3024);
nor U2857 (N_2857,In_507,In_2161);
or U2858 (N_2858,In_802,In_3391);
and U2859 (N_2859,In_972,In_3034);
xnor U2860 (N_2860,In_4817,In_3605);
xor U2861 (N_2861,In_564,In_4336);
nor U2862 (N_2862,In_3530,In_392);
and U2863 (N_2863,In_343,In_3976);
nand U2864 (N_2864,In_2958,In_4640);
nand U2865 (N_2865,In_984,In_2192);
or U2866 (N_2866,In_837,In_3524);
or U2867 (N_2867,In_1678,In_2190);
nor U2868 (N_2868,In_431,In_2915);
nor U2869 (N_2869,In_3820,In_3210);
xnor U2870 (N_2870,In_2201,In_838);
nand U2871 (N_2871,In_258,In_779);
and U2872 (N_2872,In_4103,In_4313);
nand U2873 (N_2873,In_2058,In_2296);
nor U2874 (N_2874,In_4973,In_2430);
or U2875 (N_2875,In_1410,In_1218);
nor U2876 (N_2876,In_568,In_2675);
or U2877 (N_2877,In_4992,In_4732);
nand U2878 (N_2878,In_1279,In_4086);
and U2879 (N_2879,In_3341,In_1918);
and U2880 (N_2880,In_983,In_2374);
xor U2881 (N_2881,In_1736,In_2335);
nor U2882 (N_2882,In_4276,In_2451);
xor U2883 (N_2883,In_970,In_2185);
xor U2884 (N_2884,In_4635,In_4931);
or U2885 (N_2885,In_3442,In_835);
or U2886 (N_2886,In_2598,In_407);
and U2887 (N_2887,In_1813,In_912);
nand U2888 (N_2888,In_14,In_672);
and U2889 (N_2889,In_2831,In_3947);
xnor U2890 (N_2890,In_3225,In_316);
nor U2891 (N_2891,In_3404,In_2120);
nand U2892 (N_2892,In_2069,In_4189);
or U2893 (N_2893,In_468,In_56);
nor U2894 (N_2894,In_342,In_2537);
nor U2895 (N_2895,In_774,In_701);
and U2896 (N_2896,In_4755,In_3925);
or U2897 (N_2897,In_4698,In_4082);
xor U2898 (N_2898,In_2771,In_4180);
nand U2899 (N_2899,In_2642,In_2280);
or U2900 (N_2900,In_2568,In_2248);
and U2901 (N_2901,In_1804,In_152);
nand U2902 (N_2902,In_352,In_386);
and U2903 (N_2903,In_3740,In_4069);
or U2904 (N_2904,In_4472,In_1771);
nor U2905 (N_2905,In_2540,In_30);
nand U2906 (N_2906,In_2155,In_775);
and U2907 (N_2907,In_1308,In_2525);
and U2908 (N_2908,In_817,In_4893);
or U2909 (N_2909,In_3033,In_2059);
nor U2910 (N_2910,In_4414,In_273);
or U2911 (N_2911,In_4934,In_3466);
nand U2912 (N_2912,In_4080,In_4273);
and U2913 (N_2913,In_4213,In_1689);
or U2914 (N_2914,In_4818,In_2115);
or U2915 (N_2915,In_4581,In_3033);
nor U2916 (N_2916,In_4384,In_3298);
xnor U2917 (N_2917,In_1003,In_3122);
nor U2918 (N_2918,In_2822,In_4845);
or U2919 (N_2919,In_57,In_4657);
xor U2920 (N_2920,In_2790,In_4386);
nand U2921 (N_2921,In_3302,In_857);
and U2922 (N_2922,In_2177,In_4006);
nand U2923 (N_2923,In_2968,In_1211);
and U2924 (N_2924,In_23,In_652);
and U2925 (N_2925,In_2801,In_1797);
nor U2926 (N_2926,In_2180,In_186);
and U2927 (N_2927,In_4484,In_3430);
or U2928 (N_2928,In_2934,In_1117);
nand U2929 (N_2929,In_4867,In_3790);
xnor U2930 (N_2930,In_2689,In_4307);
and U2931 (N_2931,In_791,In_4448);
nor U2932 (N_2932,In_2281,In_696);
xnor U2933 (N_2933,In_1792,In_427);
and U2934 (N_2934,In_3862,In_1527);
xor U2935 (N_2935,In_527,In_2806);
or U2936 (N_2936,In_2914,In_1792);
nor U2937 (N_2937,In_2033,In_4669);
nor U2938 (N_2938,In_1020,In_63);
or U2939 (N_2939,In_2077,In_2167);
xor U2940 (N_2940,In_1399,In_3178);
nand U2941 (N_2941,In_1946,In_2456);
nand U2942 (N_2942,In_2710,In_1288);
xor U2943 (N_2943,In_509,In_494);
nor U2944 (N_2944,In_1962,In_4431);
nor U2945 (N_2945,In_1549,In_4516);
nand U2946 (N_2946,In_846,In_830);
nor U2947 (N_2947,In_4886,In_1453);
nand U2948 (N_2948,In_704,In_4603);
nand U2949 (N_2949,In_4880,In_4610);
and U2950 (N_2950,In_4131,In_2008);
and U2951 (N_2951,In_3221,In_1462);
and U2952 (N_2952,In_2721,In_1490);
nor U2953 (N_2953,In_100,In_2817);
nor U2954 (N_2954,In_3660,In_1546);
nand U2955 (N_2955,In_4573,In_494);
xnor U2956 (N_2956,In_4983,In_3906);
xor U2957 (N_2957,In_964,In_2421);
or U2958 (N_2958,In_627,In_3485);
nor U2959 (N_2959,In_3097,In_2757);
xnor U2960 (N_2960,In_4343,In_1382);
nor U2961 (N_2961,In_246,In_1395);
nand U2962 (N_2962,In_3802,In_4057);
and U2963 (N_2963,In_1544,In_2395);
xnor U2964 (N_2964,In_938,In_2383);
or U2965 (N_2965,In_2525,In_2093);
or U2966 (N_2966,In_678,In_4422);
nand U2967 (N_2967,In_1812,In_1296);
nor U2968 (N_2968,In_4253,In_2086);
and U2969 (N_2969,In_4258,In_1682);
or U2970 (N_2970,In_941,In_671);
nand U2971 (N_2971,In_2146,In_4904);
nor U2972 (N_2972,In_3496,In_4770);
nand U2973 (N_2973,In_2483,In_3286);
nor U2974 (N_2974,In_237,In_3889);
nand U2975 (N_2975,In_3156,In_2590);
nand U2976 (N_2976,In_1613,In_3456);
nand U2977 (N_2977,In_2117,In_4190);
and U2978 (N_2978,In_2895,In_4242);
and U2979 (N_2979,In_3956,In_1225);
and U2980 (N_2980,In_598,In_1368);
xor U2981 (N_2981,In_3119,In_2554);
or U2982 (N_2982,In_3753,In_2706);
nor U2983 (N_2983,In_2828,In_3133);
xnor U2984 (N_2984,In_838,In_3817);
nand U2985 (N_2985,In_3838,In_291);
or U2986 (N_2986,In_195,In_1102);
xnor U2987 (N_2987,In_267,In_4943);
xnor U2988 (N_2988,In_3842,In_2939);
and U2989 (N_2989,In_343,In_3427);
nor U2990 (N_2990,In_3059,In_153);
or U2991 (N_2991,In_412,In_1579);
nand U2992 (N_2992,In_4846,In_1482);
and U2993 (N_2993,In_2100,In_2414);
xor U2994 (N_2994,In_299,In_2755);
nor U2995 (N_2995,In_531,In_4795);
or U2996 (N_2996,In_4301,In_4673);
xnor U2997 (N_2997,In_80,In_3323);
or U2998 (N_2998,In_3220,In_4379);
or U2999 (N_2999,In_3152,In_4408);
nand U3000 (N_3000,In_1885,In_3011);
and U3001 (N_3001,In_4331,In_2317);
xor U3002 (N_3002,In_1259,In_3620);
and U3003 (N_3003,In_2308,In_2806);
nor U3004 (N_3004,In_4969,In_1432);
and U3005 (N_3005,In_4368,In_290);
nand U3006 (N_3006,In_3718,In_2431);
xor U3007 (N_3007,In_4188,In_2876);
xor U3008 (N_3008,In_831,In_3222);
nand U3009 (N_3009,In_2168,In_1264);
xor U3010 (N_3010,In_3321,In_4476);
and U3011 (N_3011,In_4269,In_4328);
or U3012 (N_3012,In_61,In_4978);
and U3013 (N_3013,In_1965,In_110);
nor U3014 (N_3014,In_4502,In_2408);
xor U3015 (N_3015,In_668,In_4295);
and U3016 (N_3016,In_3025,In_3886);
nor U3017 (N_3017,In_1420,In_3882);
and U3018 (N_3018,In_4874,In_1668);
nor U3019 (N_3019,In_4332,In_2187);
xor U3020 (N_3020,In_4289,In_61);
or U3021 (N_3021,In_1416,In_262);
nand U3022 (N_3022,In_847,In_4503);
or U3023 (N_3023,In_2905,In_1993);
nand U3024 (N_3024,In_1677,In_3913);
and U3025 (N_3025,In_4102,In_4248);
or U3026 (N_3026,In_1948,In_4489);
or U3027 (N_3027,In_614,In_581);
nor U3028 (N_3028,In_3132,In_472);
xnor U3029 (N_3029,In_2573,In_4531);
nand U3030 (N_3030,In_335,In_3471);
xor U3031 (N_3031,In_1578,In_2814);
and U3032 (N_3032,In_571,In_3006);
xor U3033 (N_3033,In_220,In_2704);
nand U3034 (N_3034,In_4250,In_2606);
or U3035 (N_3035,In_1096,In_3986);
and U3036 (N_3036,In_3948,In_1202);
nand U3037 (N_3037,In_673,In_1308);
xnor U3038 (N_3038,In_2708,In_2838);
nand U3039 (N_3039,In_2479,In_1565);
nand U3040 (N_3040,In_948,In_1424);
or U3041 (N_3041,In_146,In_3888);
nand U3042 (N_3042,In_3241,In_2431);
nand U3043 (N_3043,In_1395,In_2016);
and U3044 (N_3044,In_3126,In_2024);
nor U3045 (N_3045,In_3853,In_1133);
xnor U3046 (N_3046,In_3637,In_2986);
xnor U3047 (N_3047,In_593,In_3259);
nand U3048 (N_3048,In_710,In_2389);
nand U3049 (N_3049,In_86,In_314);
and U3050 (N_3050,In_781,In_3816);
xor U3051 (N_3051,In_4148,In_3235);
nand U3052 (N_3052,In_3399,In_2865);
nor U3053 (N_3053,In_3816,In_3370);
nand U3054 (N_3054,In_3807,In_3578);
or U3055 (N_3055,In_4148,In_3487);
nand U3056 (N_3056,In_1186,In_2875);
or U3057 (N_3057,In_2459,In_1662);
nor U3058 (N_3058,In_3088,In_424);
nand U3059 (N_3059,In_170,In_1851);
nor U3060 (N_3060,In_4214,In_826);
xor U3061 (N_3061,In_4841,In_2258);
or U3062 (N_3062,In_3302,In_2793);
and U3063 (N_3063,In_405,In_4815);
xnor U3064 (N_3064,In_1161,In_4571);
nand U3065 (N_3065,In_4725,In_2622);
or U3066 (N_3066,In_3620,In_3808);
or U3067 (N_3067,In_4559,In_188);
xnor U3068 (N_3068,In_2305,In_732);
or U3069 (N_3069,In_3613,In_2798);
and U3070 (N_3070,In_1022,In_4654);
or U3071 (N_3071,In_3722,In_36);
xnor U3072 (N_3072,In_2925,In_592);
and U3073 (N_3073,In_133,In_2657);
nand U3074 (N_3074,In_2423,In_1220);
nor U3075 (N_3075,In_1816,In_3943);
nand U3076 (N_3076,In_76,In_1033);
xor U3077 (N_3077,In_1402,In_3957);
or U3078 (N_3078,In_4475,In_3923);
or U3079 (N_3079,In_153,In_2142);
and U3080 (N_3080,In_3337,In_16);
and U3081 (N_3081,In_169,In_4262);
nor U3082 (N_3082,In_4223,In_2944);
xnor U3083 (N_3083,In_1724,In_4522);
and U3084 (N_3084,In_1333,In_534);
and U3085 (N_3085,In_3059,In_1511);
and U3086 (N_3086,In_2043,In_2559);
nor U3087 (N_3087,In_210,In_19);
nand U3088 (N_3088,In_2265,In_408);
xor U3089 (N_3089,In_291,In_2107);
and U3090 (N_3090,In_3550,In_285);
and U3091 (N_3091,In_2566,In_2530);
or U3092 (N_3092,In_3000,In_212);
nor U3093 (N_3093,In_1108,In_2655);
xnor U3094 (N_3094,In_4186,In_4302);
or U3095 (N_3095,In_811,In_1494);
and U3096 (N_3096,In_3126,In_865);
nor U3097 (N_3097,In_3135,In_470);
or U3098 (N_3098,In_671,In_9);
nand U3099 (N_3099,In_4858,In_620);
nor U3100 (N_3100,In_2963,In_3977);
nor U3101 (N_3101,In_1428,In_137);
xnor U3102 (N_3102,In_2246,In_3224);
nor U3103 (N_3103,In_1616,In_483);
xor U3104 (N_3104,In_1810,In_411);
and U3105 (N_3105,In_1395,In_904);
nand U3106 (N_3106,In_1061,In_2658);
or U3107 (N_3107,In_694,In_3926);
nor U3108 (N_3108,In_4922,In_1512);
nand U3109 (N_3109,In_996,In_2064);
nor U3110 (N_3110,In_2964,In_1065);
and U3111 (N_3111,In_2467,In_2305);
and U3112 (N_3112,In_3733,In_3602);
nor U3113 (N_3113,In_2858,In_2001);
and U3114 (N_3114,In_889,In_3034);
or U3115 (N_3115,In_4949,In_4783);
and U3116 (N_3116,In_3505,In_4868);
nand U3117 (N_3117,In_4140,In_4736);
nand U3118 (N_3118,In_1687,In_4449);
or U3119 (N_3119,In_647,In_3324);
nor U3120 (N_3120,In_1275,In_394);
nand U3121 (N_3121,In_1831,In_902);
and U3122 (N_3122,In_1864,In_486);
xnor U3123 (N_3123,In_2572,In_1736);
nor U3124 (N_3124,In_2573,In_2311);
nor U3125 (N_3125,In_1524,In_4488);
and U3126 (N_3126,In_1963,In_569);
nand U3127 (N_3127,In_4701,In_3312);
or U3128 (N_3128,In_390,In_1977);
and U3129 (N_3129,In_771,In_3175);
xnor U3130 (N_3130,In_232,In_2949);
nand U3131 (N_3131,In_4183,In_4492);
nand U3132 (N_3132,In_2372,In_109);
xor U3133 (N_3133,In_685,In_4341);
and U3134 (N_3134,In_4623,In_1482);
and U3135 (N_3135,In_3803,In_438);
or U3136 (N_3136,In_2802,In_1830);
nor U3137 (N_3137,In_4494,In_1893);
nor U3138 (N_3138,In_3208,In_137);
nand U3139 (N_3139,In_217,In_1416);
nor U3140 (N_3140,In_360,In_2974);
or U3141 (N_3141,In_2581,In_2821);
xor U3142 (N_3142,In_3823,In_1555);
xor U3143 (N_3143,In_3501,In_227);
xor U3144 (N_3144,In_1126,In_3984);
xor U3145 (N_3145,In_2926,In_1054);
and U3146 (N_3146,In_2562,In_4854);
or U3147 (N_3147,In_4689,In_4065);
or U3148 (N_3148,In_2944,In_4807);
or U3149 (N_3149,In_4865,In_2631);
and U3150 (N_3150,In_3433,In_2349);
nor U3151 (N_3151,In_864,In_583);
nand U3152 (N_3152,In_4649,In_3517);
xnor U3153 (N_3153,In_222,In_3459);
nor U3154 (N_3154,In_1298,In_3559);
nor U3155 (N_3155,In_1218,In_3474);
xor U3156 (N_3156,In_4945,In_1742);
xnor U3157 (N_3157,In_4233,In_3735);
nor U3158 (N_3158,In_2721,In_1221);
and U3159 (N_3159,In_868,In_1958);
and U3160 (N_3160,In_4046,In_4779);
nor U3161 (N_3161,In_3258,In_4574);
xnor U3162 (N_3162,In_2400,In_512);
and U3163 (N_3163,In_1211,In_4050);
and U3164 (N_3164,In_1916,In_3789);
nor U3165 (N_3165,In_1381,In_867);
nor U3166 (N_3166,In_2961,In_2765);
nor U3167 (N_3167,In_1913,In_668);
or U3168 (N_3168,In_4393,In_583);
nor U3169 (N_3169,In_101,In_3623);
xor U3170 (N_3170,In_2690,In_2012);
xnor U3171 (N_3171,In_1985,In_491);
xnor U3172 (N_3172,In_2839,In_3054);
nor U3173 (N_3173,In_2533,In_3403);
and U3174 (N_3174,In_2857,In_3481);
and U3175 (N_3175,In_3661,In_1060);
and U3176 (N_3176,In_2927,In_1678);
xor U3177 (N_3177,In_2584,In_4186);
xor U3178 (N_3178,In_3715,In_4224);
xnor U3179 (N_3179,In_1517,In_2867);
or U3180 (N_3180,In_317,In_2500);
nor U3181 (N_3181,In_3838,In_3689);
or U3182 (N_3182,In_1167,In_3829);
xor U3183 (N_3183,In_2370,In_3544);
nor U3184 (N_3184,In_4283,In_3120);
or U3185 (N_3185,In_917,In_2800);
and U3186 (N_3186,In_460,In_3008);
xor U3187 (N_3187,In_4896,In_3682);
and U3188 (N_3188,In_2039,In_3218);
xor U3189 (N_3189,In_1966,In_3366);
and U3190 (N_3190,In_2785,In_828);
xor U3191 (N_3191,In_812,In_4519);
or U3192 (N_3192,In_2227,In_3849);
and U3193 (N_3193,In_3080,In_4510);
nand U3194 (N_3194,In_1014,In_450);
or U3195 (N_3195,In_1529,In_1090);
nor U3196 (N_3196,In_2858,In_413);
xor U3197 (N_3197,In_3428,In_3181);
and U3198 (N_3198,In_759,In_4333);
xnor U3199 (N_3199,In_101,In_1595);
xor U3200 (N_3200,In_2315,In_490);
or U3201 (N_3201,In_3256,In_830);
nor U3202 (N_3202,In_694,In_1877);
nand U3203 (N_3203,In_805,In_2193);
nand U3204 (N_3204,In_2651,In_538);
nand U3205 (N_3205,In_3723,In_3001);
nand U3206 (N_3206,In_3747,In_102);
nand U3207 (N_3207,In_4111,In_4254);
nor U3208 (N_3208,In_1172,In_3420);
xor U3209 (N_3209,In_2042,In_1300);
nand U3210 (N_3210,In_3355,In_2157);
and U3211 (N_3211,In_3416,In_2275);
nor U3212 (N_3212,In_4077,In_3576);
and U3213 (N_3213,In_4595,In_291);
or U3214 (N_3214,In_4718,In_2829);
xor U3215 (N_3215,In_318,In_4115);
nor U3216 (N_3216,In_3953,In_1375);
and U3217 (N_3217,In_3278,In_448);
nor U3218 (N_3218,In_725,In_1715);
nor U3219 (N_3219,In_23,In_4576);
or U3220 (N_3220,In_4407,In_1170);
and U3221 (N_3221,In_4075,In_4254);
xor U3222 (N_3222,In_1653,In_1238);
or U3223 (N_3223,In_2655,In_929);
xor U3224 (N_3224,In_4695,In_4674);
and U3225 (N_3225,In_3747,In_3082);
and U3226 (N_3226,In_84,In_708);
or U3227 (N_3227,In_672,In_1246);
or U3228 (N_3228,In_835,In_3447);
xnor U3229 (N_3229,In_1899,In_4691);
nand U3230 (N_3230,In_4141,In_2625);
and U3231 (N_3231,In_4285,In_2514);
or U3232 (N_3232,In_2091,In_3805);
xor U3233 (N_3233,In_4449,In_806);
or U3234 (N_3234,In_4886,In_298);
or U3235 (N_3235,In_1911,In_36);
nor U3236 (N_3236,In_137,In_749);
nor U3237 (N_3237,In_4222,In_183);
or U3238 (N_3238,In_4963,In_4374);
or U3239 (N_3239,In_1910,In_909);
xnor U3240 (N_3240,In_3769,In_2387);
or U3241 (N_3241,In_727,In_2125);
or U3242 (N_3242,In_564,In_1838);
nand U3243 (N_3243,In_4783,In_333);
nand U3244 (N_3244,In_672,In_3046);
and U3245 (N_3245,In_219,In_2074);
and U3246 (N_3246,In_2592,In_70);
xor U3247 (N_3247,In_3088,In_2470);
nor U3248 (N_3248,In_4803,In_1247);
nand U3249 (N_3249,In_1602,In_3980);
nand U3250 (N_3250,In_2726,In_3959);
xor U3251 (N_3251,In_1858,In_3646);
and U3252 (N_3252,In_3621,In_354);
nor U3253 (N_3253,In_129,In_254);
or U3254 (N_3254,In_2419,In_4404);
nand U3255 (N_3255,In_1127,In_2102);
and U3256 (N_3256,In_2154,In_3022);
and U3257 (N_3257,In_4601,In_4974);
nor U3258 (N_3258,In_3798,In_2104);
nand U3259 (N_3259,In_2703,In_292);
and U3260 (N_3260,In_2754,In_3554);
xor U3261 (N_3261,In_4176,In_1280);
nor U3262 (N_3262,In_4760,In_4639);
xor U3263 (N_3263,In_1383,In_4071);
or U3264 (N_3264,In_183,In_3);
xor U3265 (N_3265,In_4299,In_403);
and U3266 (N_3266,In_4081,In_1820);
or U3267 (N_3267,In_958,In_3479);
nor U3268 (N_3268,In_1479,In_2946);
or U3269 (N_3269,In_2294,In_4103);
nor U3270 (N_3270,In_1529,In_2371);
and U3271 (N_3271,In_3369,In_1813);
nand U3272 (N_3272,In_445,In_1027);
nor U3273 (N_3273,In_962,In_4296);
or U3274 (N_3274,In_1213,In_3651);
or U3275 (N_3275,In_3517,In_984);
and U3276 (N_3276,In_3625,In_2777);
nor U3277 (N_3277,In_904,In_2167);
nand U3278 (N_3278,In_1814,In_3210);
or U3279 (N_3279,In_2604,In_2368);
and U3280 (N_3280,In_23,In_1463);
nor U3281 (N_3281,In_2512,In_2050);
or U3282 (N_3282,In_1991,In_369);
or U3283 (N_3283,In_1584,In_1696);
nand U3284 (N_3284,In_4808,In_4442);
and U3285 (N_3285,In_2544,In_4697);
nand U3286 (N_3286,In_1422,In_1544);
nand U3287 (N_3287,In_1610,In_3324);
or U3288 (N_3288,In_234,In_2349);
xnor U3289 (N_3289,In_1611,In_754);
or U3290 (N_3290,In_2967,In_2495);
xnor U3291 (N_3291,In_952,In_110);
nor U3292 (N_3292,In_3648,In_3239);
nand U3293 (N_3293,In_20,In_4025);
nand U3294 (N_3294,In_3351,In_2807);
or U3295 (N_3295,In_1944,In_4581);
and U3296 (N_3296,In_2790,In_899);
xnor U3297 (N_3297,In_4277,In_1557);
nor U3298 (N_3298,In_4290,In_3038);
xnor U3299 (N_3299,In_2275,In_1734);
nand U3300 (N_3300,In_2710,In_284);
nand U3301 (N_3301,In_2005,In_3019);
and U3302 (N_3302,In_450,In_4618);
nand U3303 (N_3303,In_12,In_3406);
nand U3304 (N_3304,In_3478,In_764);
xnor U3305 (N_3305,In_1259,In_469);
and U3306 (N_3306,In_2872,In_2934);
nor U3307 (N_3307,In_4150,In_3786);
nor U3308 (N_3308,In_1082,In_1354);
xnor U3309 (N_3309,In_3751,In_2675);
xor U3310 (N_3310,In_2282,In_3326);
xor U3311 (N_3311,In_1972,In_341);
or U3312 (N_3312,In_3416,In_3887);
and U3313 (N_3313,In_780,In_4427);
xnor U3314 (N_3314,In_3577,In_4532);
and U3315 (N_3315,In_891,In_1154);
or U3316 (N_3316,In_1663,In_127);
and U3317 (N_3317,In_2126,In_576);
or U3318 (N_3318,In_4522,In_304);
nand U3319 (N_3319,In_282,In_2652);
nor U3320 (N_3320,In_4268,In_4324);
xor U3321 (N_3321,In_4414,In_2711);
xor U3322 (N_3322,In_653,In_1032);
nor U3323 (N_3323,In_3640,In_2781);
nor U3324 (N_3324,In_424,In_2182);
nand U3325 (N_3325,In_880,In_4356);
nand U3326 (N_3326,In_3654,In_3331);
nor U3327 (N_3327,In_2652,In_4258);
nor U3328 (N_3328,In_2374,In_1241);
nand U3329 (N_3329,In_2934,In_1838);
and U3330 (N_3330,In_975,In_4713);
nor U3331 (N_3331,In_3796,In_3760);
and U3332 (N_3332,In_2325,In_2171);
xnor U3333 (N_3333,In_647,In_4844);
nand U3334 (N_3334,In_3366,In_1778);
and U3335 (N_3335,In_298,In_1544);
nor U3336 (N_3336,In_3318,In_4963);
and U3337 (N_3337,In_1587,In_150);
and U3338 (N_3338,In_296,In_3373);
and U3339 (N_3339,In_320,In_1171);
xor U3340 (N_3340,In_4672,In_4147);
or U3341 (N_3341,In_448,In_1718);
nand U3342 (N_3342,In_3926,In_3440);
nand U3343 (N_3343,In_3406,In_4581);
nor U3344 (N_3344,In_2678,In_1573);
nand U3345 (N_3345,In_103,In_316);
nor U3346 (N_3346,In_1462,In_829);
nand U3347 (N_3347,In_1792,In_1192);
and U3348 (N_3348,In_1724,In_4827);
or U3349 (N_3349,In_640,In_2612);
nand U3350 (N_3350,In_82,In_1297);
xnor U3351 (N_3351,In_4229,In_106);
xor U3352 (N_3352,In_2854,In_4559);
nand U3353 (N_3353,In_3634,In_4944);
and U3354 (N_3354,In_2410,In_2014);
or U3355 (N_3355,In_4389,In_226);
xnor U3356 (N_3356,In_214,In_583);
nand U3357 (N_3357,In_4307,In_724);
nand U3358 (N_3358,In_595,In_2310);
nor U3359 (N_3359,In_3158,In_1124);
xnor U3360 (N_3360,In_1907,In_4520);
or U3361 (N_3361,In_4497,In_1055);
nand U3362 (N_3362,In_2806,In_3344);
xnor U3363 (N_3363,In_1537,In_1165);
and U3364 (N_3364,In_1714,In_953);
nand U3365 (N_3365,In_2068,In_622);
nor U3366 (N_3366,In_4733,In_3620);
nor U3367 (N_3367,In_1909,In_900);
nand U3368 (N_3368,In_2307,In_429);
or U3369 (N_3369,In_747,In_1700);
and U3370 (N_3370,In_3041,In_3557);
or U3371 (N_3371,In_3926,In_2036);
or U3372 (N_3372,In_483,In_1640);
or U3373 (N_3373,In_1622,In_4736);
or U3374 (N_3374,In_423,In_4794);
or U3375 (N_3375,In_612,In_3872);
xor U3376 (N_3376,In_2959,In_1720);
and U3377 (N_3377,In_3435,In_3869);
xnor U3378 (N_3378,In_4365,In_3576);
xor U3379 (N_3379,In_2389,In_3907);
nand U3380 (N_3380,In_1424,In_4153);
or U3381 (N_3381,In_2254,In_2600);
nor U3382 (N_3382,In_1142,In_354);
and U3383 (N_3383,In_2814,In_2626);
nand U3384 (N_3384,In_1443,In_3515);
or U3385 (N_3385,In_3299,In_1079);
or U3386 (N_3386,In_237,In_4564);
nand U3387 (N_3387,In_3508,In_2304);
nand U3388 (N_3388,In_690,In_4248);
nor U3389 (N_3389,In_2227,In_935);
xnor U3390 (N_3390,In_1691,In_1443);
xnor U3391 (N_3391,In_3758,In_79);
nor U3392 (N_3392,In_1133,In_2796);
nor U3393 (N_3393,In_1238,In_2585);
xnor U3394 (N_3394,In_3084,In_3236);
and U3395 (N_3395,In_1489,In_1512);
xnor U3396 (N_3396,In_1508,In_3688);
nor U3397 (N_3397,In_3668,In_4511);
nor U3398 (N_3398,In_4035,In_1407);
nor U3399 (N_3399,In_4397,In_4345);
nor U3400 (N_3400,In_1897,In_663);
xnor U3401 (N_3401,In_3035,In_718);
nand U3402 (N_3402,In_2388,In_996);
and U3403 (N_3403,In_895,In_254);
xnor U3404 (N_3404,In_261,In_2356);
or U3405 (N_3405,In_489,In_544);
nor U3406 (N_3406,In_425,In_4248);
nor U3407 (N_3407,In_762,In_721);
nor U3408 (N_3408,In_2741,In_2540);
xnor U3409 (N_3409,In_601,In_1169);
and U3410 (N_3410,In_2942,In_4390);
nor U3411 (N_3411,In_2608,In_3636);
or U3412 (N_3412,In_1370,In_4989);
nand U3413 (N_3413,In_4973,In_4962);
or U3414 (N_3414,In_4615,In_2260);
and U3415 (N_3415,In_1551,In_1541);
and U3416 (N_3416,In_2099,In_844);
nor U3417 (N_3417,In_4686,In_4812);
xor U3418 (N_3418,In_1858,In_1477);
xnor U3419 (N_3419,In_1174,In_2360);
and U3420 (N_3420,In_769,In_846);
or U3421 (N_3421,In_4307,In_3491);
and U3422 (N_3422,In_2002,In_1171);
xnor U3423 (N_3423,In_3774,In_76);
and U3424 (N_3424,In_4425,In_837);
xor U3425 (N_3425,In_2004,In_2003);
or U3426 (N_3426,In_4534,In_192);
and U3427 (N_3427,In_881,In_2715);
and U3428 (N_3428,In_1126,In_1345);
xor U3429 (N_3429,In_1282,In_2032);
nand U3430 (N_3430,In_1266,In_3150);
and U3431 (N_3431,In_1275,In_479);
and U3432 (N_3432,In_1820,In_2980);
nor U3433 (N_3433,In_2849,In_2054);
and U3434 (N_3434,In_2299,In_4766);
and U3435 (N_3435,In_597,In_3486);
nand U3436 (N_3436,In_1209,In_1400);
and U3437 (N_3437,In_2898,In_846);
nor U3438 (N_3438,In_2809,In_1538);
xnor U3439 (N_3439,In_667,In_2636);
xnor U3440 (N_3440,In_3987,In_4542);
nand U3441 (N_3441,In_4867,In_1213);
xor U3442 (N_3442,In_699,In_4248);
nand U3443 (N_3443,In_1151,In_2978);
or U3444 (N_3444,In_4829,In_2275);
or U3445 (N_3445,In_2285,In_1277);
and U3446 (N_3446,In_365,In_2334);
and U3447 (N_3447,In_1231,In_3873);
xor U3448 (N_3448,In_1291,In_752);
xor U3449 (N_3449,In_2163,In_54);
nor U3450 (N_3450,In_2747,In_869);
xnor U3451 (N_3451,In_4056,In_3633);
and U3452 (N_3452,In_172,In_2440);
or U3453 (N_3453,In_1864,In_3380);
or U3454 (N_3454,In_1637,In_270);
nand U3455 (N_3455,In_3278,In_635);
and U3456 (N_3456,In_1451,In_3846);
xnor U3457 (N_3457,In_3241,In_4663);
nand U3458 (N_3458,In_1183,In_3079);
nor U3459 (N_3459,In_1068,In_213);
and U3460 (N_3460,In_4461,In_2440);
and U3461 (N_3461,In_2336,In_431);
nand U3462 (N_3462,In_2642,In_2614);
or U3463 (N_3463,In_1279,In_2902);
xnor U3464 (N_3464,In_4479,In_1219);
nand U3465 (N_3465,In_2364,In_4979);
and U3466 (N_3466,In_296,In_4236);
or U3467 (N_3467,In_2946,In_1168);
nand U3468 (N_3468,In_1287,In_2635);
nand U3469 (N_3469,In_1327,In_4837);
or U3470 (N_3470,In_3512,In_2658);
nor U3471 (N_3471,In_1502,In_1665);
xor U3472 (N_3472,In_1708,In_4581);
nor U3473 (N_3473,In_1230,In_4275);
and U3474 (N_3474,In_4444,In_852);
and U3475 (N_3475,In_167,In_1541);
xor U3476 (N_3476,In_4872,In_2942);
xnor U3477 (N_3477,In_1798,In_3542);
or U3478 (N_3478,In_2978,In_1234);
xnor U3479 (N_3479,In_1301,In_732);
xnor U3480 (N_3480,In_447,In_3366);
nand U3481 (N_3481,In_4421,In_3402);
nor U3482 (N_3482,In_3368,In_3726);
and U3483 (N_3483,In_3704,In_292);
nand U3484 (N_3484,In_165,In_3517);
or U3485 (N_3485,In_3073,In_1960);
and U3486 (N_3486,In_4951,In_241);
nand U3487 (N_3487,In_3629,In_2450);
nand U3488 (N_3488,In_4307,In_355);
xnor U3489 (N_3489,In_2627,In_1409);
or U3490 (N_3490,In_330,In_1553);
or U3491 (N_3491,In_790,In_1949);
nor U3492 (N_3492,In_3450,In_3004);
xor U3493 (N_3493,In_479,In_3109);
nor U3494 (N_3494,In_1447,In_4725);
nor U3495 (N_3495,In_4873,In_1141);
nand U3496 (N_3496,In_4874,In_2332);
nand U3497 (N_3497,In_1473,In_1971);
xor U3498 (N_3498,In_3571,In_913);
xnor U3499 (N_3499,In_4503,In_718);
nand U3500 (N_3500,In_629,In_3674);
nor U3501 (N_3501,In_2738,In_836);
nor U3502 (N_3502,In_401,In_2793);
or U3503 (N_3503,In_1163,In_679);
or U3504 (N_3504,In_2235,In_1844);
xnor U3505 (N_3505,In_3003,In_4394);
xnor U3506 (N_3506,In_4624,In_1644);
xor U3507 (N_3507,In_4766,In_1691);
nand U3508 (N_3508,In_333,In_3791);
and U3509 (N_3509,In_842,In_4738);
xor U3510 (N_3510,In_4886,In_471);
xnor U3511 (N_3511,In_2426,In_4850);
nand U3512 (N_3512,In_3114,In_4830);
and U3513 (N_3513,In_4672,In_4462);
nand U3514 (N_3514,In_2232,In_3518);
and U3515 (N_3515,In_3476,In_4488);
xnor U3516 (N_3516,In_4931,In_1518);
nor U3517 (N_3517,In_3965,In_2187);
xnor U3518 (N_3518,In_4677,In_3066);
nor U3519 (N_3519,In_412,In_2385);
or U3520 (N_3520,In_2007,In_4280);
and U3521 (N_3521,In_1988,In_2184);
and U3522 (N_3522,In_1299,In_1666);
nand U3523 (N_3523,In_1369,In_3935);
nor U3524 (N_3524,In_4250,In_4786);
nor U3525 (N_3525,In_2193,In_3303);
and U3526 (N_3526,In_3044,In_1464);
nand U3527 (N_3527,In_2871,In_1141);
nand U3528 (N_3528,In_140,In_3851);
nor U3529 (N_3529,In_2489,In_2784);
xnor U3530 (N_3530,In_4549,In_32);
or U3531 (N_3531,In_2163,In_4997);
xor U3532 (N_3532,In_1087,In_3520);
xor U3533 (N_3533,In_2813,In_1023);
or U3534 (N_3534,In_2320,In_469);
nand U3535 (N_3535,In_285,In_2496);
xor U3536 (N_3536,In_319,In_2536);
nand U3537 (N_3537,In_2145,In_3643);
nand U3538 (N_3538,In_52,In_2061);
or U3539 (N_3539,In_2139,In_54);
nor U3540 (N_3540,In_4341,In_4787);
or U3541 (N_3541,In_749,In_1453);
nand U3542 (N_3542,In_4615,In_1813);
xor U3543 (N_3543,In_4390,In_2854);
and U3544 (N_3544,In_1279,In_3721);
nor U3545 (N_3545,In_735,In_4728);
nor U3546 (N_3546,In_518,In_1183);
or U3547 (N_3547,In_2316,In_1438);
nor U3548 (N_3548,In_3593,In_3607);
xnor U3549 (N_3549,In_559,In_4875);
xor U3550 (N_3550,In_3163,In_884);
nand U3551 (N_3551,In_428,In_4150);
or U3552 (N_3552,In_2954,In_1025);
nor U3553 (N_3553,In_3325,In_2402);
xnor U3554 (N_3554,In_3779,In_2788);
nand U3555 (N_3555,In_1319,In_198);
or U3556 (N_3556,In_55,In_4268);
nor U3557 (N_3557,In_152,In_3776);
nor U3558 (N_3558,In_157,In_4586);
nand U3559 (N_3559,In_2533,In_2760);
and U3560 (N_3560,In_1775,In_4122);
and U3561 (N_3561,In_634,In_2256);
xor U3562 (N_3562,In_1154,In_2907);
or U3563 (N_3563,In_1460,In_430);
xnor U3564 (N_3564,In_4850,In_1474);
or U3565 (N_3565,In_1789,In_3377);
nand U3566 (N_3566,In_1932,In_1740);
or U3567 (N_3567,In_2466,In_1660);
or U3568 (N_3568,In_4080,In_548);
nand U3569 (N_3569,In_2015,In_2399);
or U3570 (N_3570,In_774,In_3740);
nand U3571 (N_3571,In_2958,In_883);
or U3572 (N_3572,In_1089,In_1583);
and U3573 (N_3573,In_4530,In_1045);
or U3574 (N_3574,In_2348,In_827);
and U3575 (N_3575,In_4656,In_3500);
nor U3576 (N_3576,In_461,In_4550);
nor U3577 (N_3577,In_3287,In_1960);
nor U3578 (N_3578,In_3061,In_3198);
and U3579 (N_3579,In_2337,In_1313);
and U3580 (N_3580,In_2870,In_4362);
and U3581 (N_3581,In_1304,In_1573);
nor U3582 (N_3582,In_250,In_3154);
xor U3583 (N_3583,In_3498,In_2821);
nand U3584 (N_3584,In_1191,In_4861);
nor U3585 (N_3585,In_849,In_3746);
nand U3586 (N_3586,In_3527,In_1508);
and U3587 (N_3587,In_3528,In_4889);
and U3588 (N_3588,In_2885,In_409);
xor U3589 (N_3589,In_750,In_2002);
xnor U3590 (N_3590,In_4526,In_3125);
and U3591 (N_3591,In_3246,In_2914);
nand U3592 (N_3592,In_4677,In_4645);
and U3593 (N_3593,In_2567,In_2756);
nor U3594 (N_3594,In_3966,In_4790);
nand U3595 (N_3595,In_689,In_2855);
xor U3596 (N_3596,In_318,In_358);
nand U3597 (N_3597,In_2669,In_4973);
xor U3598 (N_3598,In_4386,In_1742);
xnor U3599 (N_3599,In_2893,In_1654);
nand U3600 (N_3600,In_1533,In_4503);
nor U3601 (N_3601,In_465,In_1601);
nand U3602 (N_3602,In_266,In_4001);
nand U3603 (N_3603,In_4626,In_2614);
nand U3604 (N_3604,In_609,In_3910);
nor U3605 (N_3605,In_1637,In_766);
xnor U3606 (N_3606,In_4257,In_1601);
and U3607 (N_3607,In_289,In_4910);
and U3608 (N_3608,In_2812,In_384);
xor U3609 (N_3609,In_792,In_4650);
and U3610 (N_3610,In_2205,In_563);
xnor U3611 (N_3611,In_4442,In_1951);
and U3612 (N_3612,In_2608,In_2881);
nor U3613 (N_3613,In_3154,In_424);
nand U3614 (N_3614,In_1413,In_3073);
or U3615 (N_3615,In_2135,In_525);
and U3616 (N_3616,In_514,In_4850);
xnor U3617 (N_3617,In_3764,In_2175);
xnor U3618 (N_3618,In_606,In_732);
xnor U3619 (N_3619,In_1360,In_3765);
xor U3620 (N_3620,In_1325,In_1808);
nand U3621 (N_3621,In_387,In_2312);
nand U3622 (N_3622,In_4341,In_3287);
xnor U3623 (N_3623,In_2170,In_4251);
xor U3624 (N_3624,In_3825,In_1300);
or U3625 (N_3625,In_3362,In_4990);
and U3626 (N_3626,In_1934,In_2919);
nand U3627 (N_3627,In_3353,In_1348);
xnor U3628 (N_3628,In_1505,In_783);
nand U3629 (N_3629,In_4561,In_2538);
nor U3630 (N_3630,In_2921,In_3248);
xor U3631 (N_3631,In_2864,In_1863);
and U3632 (N_3632,In_10,In_2224);
or U3633 (N_3633,In_3711,In_6);
or U3634 (N_3634,In_996,In_2358);
or U3635 (N_3635,In_4532,In_3840);
nor U3636 (N_3636,In_2618,In_2926);
xnor U3637 (N_3637,In_1537,In_4547);
or U3638 (N_3638,In_2489,In_4666);
and U3639 (N_3639,In_3891,In_3647);
nand U3640 (N_3640,In_2404,In_1805);
or U3641 (N_3641,In_892,In_1634);
nand U3642 (N_3642,In_1789,In_277);
nand U3643 (N_3643,In_2866,In_1710);
xnor U3644 (N_3644,In_3093,In_733);
and U3645 (N_3645,In_2752,In_1773);
xor U3646 (N_3646,In_3287,In_3765);
and U3647 (N_3647,In_1733,In_3503);
or U3648 (N_3648,In_1008,In_4814);
and U3649 (N_3649,In_3069,In_3370);
nand U3650 (N_3650,In_4821,In_4887);
or U3651 (N_3651,In_955,In_1460);
xor U3652 (N_3652,In_334,In_353);
xnor U3653 (N_3653,In_2629,In_1608);
and U3654 (N_3654,In_1249,In_2262);
nand U3655 (N_3655,In_4831,In_589);
nor U3656 (N_3656,In_442,In_1963);
nand U3657 (N_3657,In_4853,In_3687);
nand U3658 (N_3658,In_3098,In_1205);
or U3659 (N_3659,In_2386,In_2019);
nor U3660 (N_3660,In_2548,In_3875);
and U3661 (N_3661,In_4900,In_1465);
and U3662 (N_3662,In_4857,In_1768);
nand U3663 (N_3663,In_1686,In_4863);
xor U3664 (N_3664,In_3164,In_4155);
nor U3665 (N_3665,In_2891,In_402);
nor U3666 (N_3666,In_2836,In_2369);
xor U3667 (N_3667,In_1814,In_2280);
nand U3668 (N_3668,In_240,In_3242);
xor U3669 (N_3669,In_3944,In_3381);
nor U3670 (N_3670,In_250,In_2661);
or U3671 (N_3671,In_4577,In_2132);
nand U3672 (N_3672,In_4620,In_400);
or U3673 (N_3673,In_441,In_731);
or U3674 (N_3674,In_357,In_2362);
xor U3675 (N_3675,In_981,In_3913);
xnor U3676 (N_3676,In_23,In_57);
xor U3677 (N_3677,In_1692,In_1921);
and U3678 (N_3678,In_4837,In_4074);
nor U3679 (N_3679,In_4379,In_4426);
xor U3680 (N_3680,In_1353,In_577);
xor U3681 (N_3681,In_853,In_233);
or U3682 (N_3682,In_4699,In_3951);
nor U3683 (N_3683,In_453,In_3816);
nor U3684 (N_3684,In_2751,In_2095);
nand U3685 (N_3685,In_3146,In_1343);
and U3686 (N_3686,In_1820,In_3787);
xnor U3687 (N_3687,In_1906,In_4191);
nand U3688 (N_3688,In_1918,In_1887);
or U3689 (N_3689,In_4782,In_3689);
and U3690 (N_3690,In_155,In_4167);
xor U3691 (N_3691,In_4668,In_778);
nor U3692 (N_3692,In_296,In_2549);
and U3693 (N_3693,In_4375,In_2704);
or U3694 (N_3694,In_2581,In_2089);
nor U3695 (N_3695,In_2057,In_4415);
or U3696 (N_3696,In_4328,In_3507);
nand U3697 (N_3697,In_599,In_2892);
and U3698 (N_3698,In_829,In_1677);
xnor U3699 (N_3699,In_2565,In_432);
xor U3700 (N_3700,In_4265,In_1843);
nor U3701 (N_3701,In_3638,In_579);
nand U3702 (N_3702,In_4730,In_2209);
nor U3703 (N_3703,In_2660,In_3005);
and U3704 (N_3704,In_2856,In_2543);
nor U3705 (N_3705,In_2653,In_666);
nor U3706 (N_3706,In_998,In_4381);
nor U3707 (N_3707,In_1504,In_1397);
nand U3708 (N_3708,In_1557,In_1357);
and U3709 (N_3709,In_3889,In_1283);
or U3710 (N_3710,In_4671,In_2382);
and U3711 (N_3711,In_805,In_352);
and U3712 (N_3712,In_2199,In_4497);
nor U3713 (N_3713,In_1954,In_4574);
xor U3714 (N_3714,In_582,In_3419);
or U3715 (N_3715,In_3551,In_3630);
xnor U3716 (N_3716,In_4577,In_2087);
nand U3717 (N_3717,In_586,In_3978);
nor U3718 (N_3718,In_3697,In_3213);
and U3719 (N_3719,In_2685,In_2116);
xnor U3720 (N_3720,In_3402,In_2071);
xor U3721 (N_3721,In_2119,In_2952);
or U3722 (N_3722,In_3792,In_2467);
xor U3723 (N_3723,In_4031,In_71);
and U3724 (N_3724,In_3697,In_4327);
nor U3725 (N_3725,In_2967,In_3302);
nand U3726 (N_3726,In_1867,In_1692);
and U3727 (N_3727,In_4986,In_4195);
nor U3728 (N_3728,In_2253,In_2818);
xor U3729 (N_3729,In_1503,In_3097);
nand U3730 (N_3730,In_3577,In_2380);
and U3731 (N_3731,In_1980,In_1554);
xnor U3732 (N_3732,In_2770,In_1459);
or U3733 (N_3733,In_1102,In_2590);
nand U3734 (N_3734,In_1275,In_136);
nand U3735 (N_3735,In_81,In_3602);
or U3736 (N_3736,In_2738,In_2285);
nor U3737 (N_3737,In_3302,In_2964);
or U3738 (N_3738,In_4326,In_4463);
nor U3739 (N_3739,In_2819,In_2671);
nand U3740 (N_3740,In_2451,In_1052);
nand U3741 (N_3741,In_2843,In_4981);
or U3742 (N_3742,In_631,In_188);
nand U3743 (N_3743,In_3106,In_1534);
nor U3744 (N_3744,In_744,In_4963);
and U3745 (N_3745,In_782,In_3384);
or U3746 (N_3746,In_3151,In_3839);
xor U3747 (N_3747,In_3046,In_3662);
xor U3748 (N_3748,In_1752,In_3378);
or U3749 (N_3749,In_4193,In_883);
and U3750 (N_3750,In_4268,In_2901);
nand U3751 (N_3751,In_544,In_1483);
nand U3752 (N_3752,In_1229,In_3317);
or U3753 (N_3753,In_4671,In_901);
xor U3754 (N_3754,In_755,In_1844);
nor U3755 (N_3755,In_483,In_1770);
nand U3756 (N_3756,In_1999,In_4361);
and U3757 (N_3757,In_4348,In_3851);
nor U3758 (N_3758,In_3340,In_3264);
xnor U3759 (N_3759,In_4747,In_179);
nand U3760 (N_3760,In_3461,In_4513);
xnor U3761 (N_3761,In_4378,In_3264);
xor U3762 (N_3762,In_115,In_1719);
nand U3763 (N_3763,In_1977,In_2237);
xnor U3764 (N_3764,In_328,In_3070);
nand U3765 (N_3765,In_4371,In_3358);
or U3766 (N_3766,In_1693,In_2403);
or U3767 (N_3767,In_3272,In_1193);
nand U3768 (N_3768,In_33,In_2335);
xnor U3769 (N_3769,In_2907,In_3608);
nand U3770 (N_3770,In_674,In_4056);
xnor U3771 (N_3771,In_4744,In_434);
nor U3772 (N_3772,In_2851,In_2971);
nand U3773 (N_3773,In_955,In_4122);
nor U3774 (N_3774,In_3670,In_469);
xnor U3775 (N_3775,In_1353,In_3796);
nor U3776 (N_3776,In_1950,In_2996);
nand U3777 (N_3777,In_3310,In_4960);
and U3778 (N_3778,In_2576,In_2614);
nor U3779 (N_3779,In_3637,In_2883);
or U3780 (N_3780,In_2360,In_3933);
nor U3781 (N_3781,In_13,In_635);
nor U3782 (N_3782,In_396,In_4753);
xor U3783 (N_3783,In_77,In_3571);
nor U3784 (N_3784,In_3595,In_1495);
or U3785 (N_3785,In_272,In_3363);
nor U3786 (N_3786,In_303,In_564);
nor U3787 (N_3787,In_1765,In_4465);
nand U3788 (N_3788,In_2976,In_2476);
or U3789 (N_3789,In_1465,In_27);
and U3790 (N_3790,In_4560,In_2940);
xor U3791 (N_3791,In_415,In_912);
nand U3792 (N_3792,In_765,In_4236);
or U3793 (N_3793,In_3738,In_4610);
xor U3794 (N_3794,In_3640,In_45);
and U3795 (N_3795,In_3735,In_1005);
nand U3796 (N_3796,In_3501,In_140);
xor U3797 (N_3797,In_1955,In_2524);
nand U3798 (N_3798,In_3236,In_4887);
or U3799 (N_3799,In_2616,In_546);
nand U3800 (N_3800,In_1780,In_216);
xor U3801 (N_3801,In_2163,In_4372);
xor U3802 (N_3802,In_3646,In_435);
xor U3803 (N_3803,In_1704,In_3521);
nand U3804 (N_3804,In_365,In_3989);
and U3805 (N_3805,In_2336,In_2086);
and U3806 (N_3806,In_2431,In_363);
or U3807 (N_3807,In_4045,In_1001);
and U3808 (N_3808,In_2672,In_3122);
or U3809 (N_3809,In_3407,In_3231);
xor U3810 (N_3810,In_4013,In_1129);
or U3811 (N_3811,In_4053,In_4404);
or U3812 (N_3812,In_1086,In_825);
nand U3813 (N_3813,In_4659,In_2004);
nand U3814 (N_3814,In_2206,In_4400);
nor U3815 (N_3815,In_3828,In_393);
nor U3816 (N_3816,In_2404,In_4906);
nand U3817 (N_3817,In_1411,In_2447);
nand U3818 (N_3818,In_456,In_3198);
nor U3819 (N_3819,In_1658,In_2257);
xnor U3820 (N_3820,In_1300,In_386);
nand U3821 (N_3821,In_935,In_3285);
and U3822 (N_3822,In_2852,In_3958);
and U3823 (N_3823,In_1149,In_46);
or U3824 (N_3824,In_3916,In_4307);
and U3825 (N_3825,In_2655,In_1503);
and U3826 (N_3826,In_4627,In_3999);
and U3827 (N_3827,In_4129,In_2810);
xor U3828 (N_3828,In_323,In_1608);
xor U3829 (N_3829,In_345,In_3669);
and U3830 (N_3830,In_678,In_3922);
and U3831 (N_3831,In_4396,In_4386);
or U3832 (N_3832,In_2203,In_1749);
or U3833 (N_3833,In_958,In_1568);
and U3834 (N_3834,In_613,In_3585);
and U3835 (N_3835,In_4761,In_1963);
xor U3836 (N_3836,In_1777,In_4764);
xor U3837 (N_3837,In_4559,In_2361);
and U3838 (N_3838,In_841,In_4385);
or U3839 (N_3839,In_4006,In_2822);
nor U3840 (N_3840,In_527,In_624);
and U3841 (N_3841,In_1197,In_1115);
nand U3842 (N_3842,In_2220,In_2028);
and U3843 (N_3843,In_2986,In_23);
xnor U3844 (N_3844,In_1776,In_1545);
xnor U3845 (N_3845,In_4609,In_746);
or U3846 (N_3846,In_315,In_404);
nand U3847 (N_3847,In_872,In_2030);
or U3848 (N_3848,In_2146,In_441);
nand U3849 (N_3849,In_4338,In_2712);
and U3850 (N_3850,In_96,In_4048);
xor U3851 (N_3851,In_3051,In_4711);
nand U3852 (N_3852,In_1327,In_4397);
xor U3853 (N_3853,In_1819,In_2709);
or U3854 (N_3854,In_3264,In_3784);
or U3855 (N_3855,In_1535,In_106);
nand U3856 (N_3856,In_1431,In_4559);
or U3857 (N_3857,In_65,In_2213);
nor U3858 (N_3858,In_2077,In_4704);
or U3859 (N_3859,In_1398,In_854);
or U3860 (N_3860,In_2190,In_1495);
and U3861 (N_3861,In_2997,In_1);
or U3862 (N_3862,In_4403,In_2816);
and U3863 (N_3863,In_3840,In_2594);
nor U3864 (N_3864,In_4015,In_3403);
xor U3865 (N_3865,In_3372,In_2866);
xnor U3866 (N_3866,In_4507,In_2586);
and U3867 (N_3867,In_240,In_1304);
and U3868 (N_3868,In_3533,In_1330);
or U3869 (N_3869,In_3940,In_3601);
and U3870 (N_3870,In_3386,In_220);
nor U3871 (N_3871,In_2089,In_641);
nand U3872 (N_3872,In_3546,In_2750);
nor U3873 (N_3873,In_2212,In_3882);
xor U3874 (N_3874,In_4936,In_4841);
and U3875 (N_3875,In_3899,In_2471);
xor U3876 (N_3876,In_2856,In_2414);
nand U3877 (N_3877,In_3754,In_2854);
xnor U3878 (N_3878,In_3806,In_2506);
nand U3879 (N_3879,In_2659,In_2349);
nor U3880 (N_3880,In_2985,In_2759);
xor U3881 (N_3881,In_4181,In_1665);
nor U3882 (N_3882,In_3332,In_4909);
or U3883 (N_3883,In_1735,In_4144);
nor U3884 (N_3884,In_1935,In_655);
nand U3885 (N_3885,In_2222,In_630);
nand U3886 (N_3886,In_1130,In_184);
nor U3887 (N_3887,In_4001,In_519);
nor U3888 (N_3888,In_3503,In_4940);
or U3889 (N_3889,In_3602,In_3902);
nor U3890 (N_3890,In_2958,In_3453);
nand U3891 (N_3891,In_2995,In_1384);
or U3892 (N_3892,In_1411,In_587);
and U3893 (N_3893,In_1146,In_2499);
nor U3894 (N_3894,In_4417,In_2499);
nand U3895 (N_3895,In_1505,In_2641);
nor U3896 (N_3896,In_2008,In_2293);
or U3897 (N_3897,In_2972,In_3074);
or U3898 (N_3898,In_3578,In_196);
nand U3899 (N_3899,In_4142,In_89);
nand U3900 (N_3900,In_2008,In_1047);
xor U3901 (N_3901,In_3085,In_2943);
and U3902 (N_3902,In_223,In_3107);
xnor U3903 (N_3903,In_2387,In_2433);
and U3904 (N_3904,In_712,In_1727);
nand U3905 (N_3905,In_4453,In_229);
and U3906 (N_3906,In_1987,In_4911);
and U3907 (N_3907,In_383,In_2016);
xor U3908 (N_3908,In_3626,In_1737);
xor U3909 (N_3909,In_2792,In_3015);
xnor U3910 (N_3910,In_731,In_2031);
nor U3911 (N_3911,In_4323,In_147);
and U3912 (N_3912,In_1004,In_2397);
or U3913 (N_3913,In_4776,In_1325);
xor U3914 (N_3914,In_1144,In_3089);
and U3915 (N_3915,In_4578,In_1183);
xor U3916 (N_3916,In_1085,In_3543);
or U3917 (N_3917,In_4411,In_2560);
nand U3918 (N_3918,In_3768,In_3032);
nor U3919 (N_3919,In_9,In_762);
xnor U3920 (N_3920,In_4081,In_4812);
nor U3921 (N_3921,In_3249,In_1672);
xnor U3922 (N_3922,In_327,In_3997);
and U3923 (N_3923,In_1044,In_2113);
nor U3924 (N_3924,In_993,In_842);
and U3925 (N_3925,In_2587,In_1144);
nor U3926 (N_3926,In_845,In_3615);
or U3927 (N_3927,In_3009,In_4866);
and U3928 (N_3928,In_3372,In_1183);
xnor U3929 (N_3929,In_818,In_98);
nor U3930 (N_3930,In_4356,In_2897);
xnor U3931 (N_3931,In_914,In_790);
xnor U3932 (N_3932,In_3386,In_194);
xor U3933 (N_3933,In_1277,In_2526);
nand U3934 (N_3934,In_3962,In_1052);
xor U3935 (N_3935,In_1921,In_2111);
or U3936 (N_3936,In_2845,In_1994);
or U3937 (N_3937,In_3548,In_2472);
nand U3938 (N_3938,In_4034,In_861);
nor U3939 (N_3939,In_4538,In_4470);
or U3940 (N_3940,In_4259,In_294);
xnor U3941 (N_3941,In_3101,In_3051);
xor U3942 (N_3942,In_1599,In_2590);
xor U3943 (N_3943,In_2899,In_3647);
nor U3944 (N_3944,In_4247,In_4225);
nor U3945 (N_3945,In_1853,In_3905);
xor U3946 (N_3946,In_1269,In_3009);
nand U3947 (N_3947,In_4405,In_4878);
xnor U3948 (N_3948,In_3881,In_713);
nand U3949 (N_3949,In_1417,In_1355);
xor U3950 (N_3950,In_4425,In_2134);
or U3951 (N_3951,In_4886,In_2529);
and U3952 (N_3952,In_764,In_2874);
and U3953 (N_3953,In_2419,In_3288);
or U3954 (N_3954,In_607,In_2641);
xor U3955 (N_3955,In_4737,In_3660);
nand U3956 (N_3956,In_4697,In_2279);
and U3957 (N_3957,In_3575,In_1734);
nor U3958 (N_3958,In_3548,In_2774);
nor U3959 (N_3959,In_1377,In_3763);
or U3960 (N_3960,In_4633,In_3430);
and U3961 (N_3961,In_4984,In_3150);
or U3962 (N_3962,In_4979,In_676);
xnor U3963 (N_3963,In_1151,In_3076);
and U3964 (N_3964,In_626,In_1144);
xor U3965 (N_3965,In_3764,In_1454);
nand U3966 (N_3966,In_4604,In_1680);
nor U3967 (N_3967,In_1210,In_4720);
nand U3968 (N_3968,In_281,In_2025);
and U3969 (N_3969,In_73,In_4209);
xor U3970 (N_3970,In_508,In_3946);
xor U3971 (N_3971,In_3920,In_118);
nor U3972 (N_3972,In_4986,In_1626);
nor U3973 (N_3973,In_347,In_201);
nor U3974 (N_3974,In_4291,In_23);
and U3975 (N_3975,In_2103,In_3060);
xor U3976 (N_3976,In_4954,In_177);
or U3977 (N_3977,In_1052,In_2263);
or U3978 (N_3978,In_3287,In_4462);
nor U3979 (N_3979,In_243,In_2249);
xnor U3980 (N_3980,In_2887,In_1337);
xnor U3981 (N_3981,In_2948,In_4717);
xnor U3982 (N_3982,In_40,In_4773);
or U3983 (N_3983,In_4070,In_870);
xor U3984 (N_3984,In_518,In_50);
xor U3985 (N_3985,In_2416,In_78);
xor U3986 (N_3986,In_2714,In_1363);
nand U3987 (N_3987,In_1168,In_4329);
nor U3988 (N_3988,In_3060,In_1059);
or U3989 (N_3989,In_1537,In_3007);
and U3990 (N_3990,In_1200,In_2176);
or U3991 (N_3991,In_1453,In_4190);
and U3992 (N_3992,In_1317,In_2255);
nor U3993 (N_3993,In_3982,In_2987);
xnor U3994 (N_3994,In_3214,In_141);
nor U3995 (N_3995,In_3717,In_975);
nor U3996 (N_3996,In_2551,In_2267);
nand U3997 (N_3997,In_2164,In_2296);
nand U3998 (N_3998,In_2439,In_1573);
nor U3999 (N_3999,In_4003,In_2623);
or U4000 (N_4000,In_2992,In_4266);
and U4001 (N_4001,In_3995,In_1234);
or U4002 (N_4002,In_3230,In_1738);
nand U4003 (N_4003,In_1743,In_3588);
xor U4004 (N_4004,In_4968,In_3413);
nand U4005 (N_4005,In_3311,In_1073);
or U4006 (N_4006,In_2125,In_827);
nor U4007 (N_4007,In_4863,In_3029);
nor U4008 (N_4008,In_234,In_3963);
nor U4009 (N_4009,In_4238,In_4139);
nor U4010 (N_4010,In_4070,In_1913);
and U4011 (N_4011,In_3185,In_2395);
nand U4012 (N_4012,In_1473,In_4669);
xor U4013 (N_4013,In_3037,In_3758);
or U4014 (N_4014,In_2223,In_1306);
or U4015 (N_4015,In_1497,In_565);
and U4016 (N_4016,In_258,In_2823);
or U4017 (N_4017,In_2183,In_2833);
or U4018 (N_4018,In_778,In_726);
nand U4019 (N_4019,In_2922,In_4579);
nand U4020 (N_4020,In_4091,In_4090);
or U4021 (N_4021,In_2351,In_3234);
and U4022 (N_4022,In_4843,In_4333);
and U4023 (N_4023,In_1757,In_863);
or U4024 (N_4024,In_2864,In_904);
nor U4025 (N_4025,In_4002,In_3820);
xor U4026 (N_4026,In_2440,In_3810);
nor U4027 (N_4027,In_4451,In_3731);
nor U4028 (N_4028,In_2104,In_976);
or U4029 (N_4029,In_964,In_2833);
or U4030 (N_4030,In_3919,In_1320);
nor U4031 (N_4031,In_2842,In_1725);
or U4032 (N_4032,In_1209,In_2670);
and U4033 (N_4033,In_2924,In_4696);
xor U4034 (N_4034,In_1541,In_1930);
xnor U4035 (N_4035,In_4057,In_4861);
nor U4036 (N_4036,In_1024,In_3475);
nand U4037 (N_4037,In_877,In_886);
xnor U4038 (N_4038,In_3827,In_2726);
nor U4039 (N_4039,In_2167,In_3427);
nand U4040 (N_4040,In_5,In_3514);
nor U4041 (N_4041,In_1509,In_3442);
nor U4042 (N_4042,In_2929,In_2337);
nor U4043 (N_4043,In_1919,In_2708);
nand U4044 (N_4044,In_259,In_4862);
or U4045 (N_4045,In_2227,In_4230);
nor U4046 (N_4046,In_2047,In_1515);
xnor U4047 (N_4047,In_1451,In_4263);
nor U4048 (N_4048,In_1807,In_3136);
and U4049 (N_4049,In_801,In_2395);
xor U4050 (N_4050,In_878,In_4848);
nand U4051 (N_4051,In_1668,In_3321);
nand U4052 (N_4052,In_760,In_1066);
and U4053 (N_4053,In_1122,In_1448);
nand U4054 (N_4054,In_2505,In_3658);
and U4055 (N_4055,In_497,In_516);
or U4056 (N_4056,In_964,In_2193);
nor U4057 (N_4057,In_442,In_631);
or U4058 (N_4058,In_1321,In_2810);
nand U4059 (N_4059,In_689,In_4596);
or U4060 (N_4060,In_4098,In_201);
or U4061 (N_4061,In_1549,In_494);
and U4062 (N_4062,In_4858,In_1431);
and U4063 (N_4063,In_2879,In_4085);
or U4064 (N_4064,In_3853,In_3955);
xnor U4065 (N_4065,In_312,In_4399);
nand U4066 (N_4066,In_1100,In_663);
xnor U4067 (N_4067,In_3829,In_3049);
xor U4068 (N_4068,In_3902,In_1294);
or U4069 (N_4069,In_2028,In_4326);
and U4070 (N_4070,In_3299,In_708);
or U4071 (N_4071,In_921,In_653);
nand U4072 (N_4072,In_677,In_503);
and U4073 (N_4073,In_1764,In_4343);
or U4074 (N_4074,In_3754,In_352);
and U4075 (N_4075,In_118,In_4414);
or U4076 (N_4076,In_686,In_4654);
or U4077 (N_4077,In_1394,In_3234);
xor U4078 (N_4078,In_2905,In_4592);
xnor U4079 (N_4079,In_1337,In_4918);
nor U4080 (N_4080,In_2691,In_2777);
and U4081 (N_4081,In_3825,In_885);
or U4082 (N_4082,In_2427,In_3318);
or U4083 (N_4083,In_4855,In_1546);
nor U4084 (N_4084,In_3931,In_864);
nand U4085 (N_4085,In_1339,In_1364);
xnor U4086 (N_4086,In_2723,In_3597);
or U4087 (N_4087,In_1492,In_3441);
and U4088 (N_4088,In_1670,In_840);
nor U4089 (N_4089,In_1119,In_1055);
nand U4090 (N_4090,In_812,In_346);
nand U4091 (N_4091,In_3526,In_453);
nand U4092 (N_4092,In_998,In_1862);
or U4093 (N_4093,In_4782,In_412);
xor U4094 (N_4094,In_3005,In_1053);
xnor U4095 (N_4095,In_2828,In_2426);
nand U4096 (N_4096,In_3417,In_1008);
nand U4097 (N_4097,In_2424,In_1383);
nor U4098 (N_4098,In_1477,In_3787);
or U4099 (N_4099,In_3347,In_4863);
and U4100 (N_4100,In_4170,In_3644);
nor U4101 (N_4101,In_3846,In_3258);
xor U4102 (N_4102,In_163,In_292);
and U4103 (N_4103,In_588,In_2356);
or U4104 (N_4104,In_426,In_625);
and U4105 (N_4105,In_3413,In_4785);
or U4106 (N_4106,In_568,In_3465);
or U4107 (N_4107,In_4191,In_4773);
xor U4108 (N_4108,In_775,In_2168);
nand U4109 (N_4109,In_1021,In_2285);
and U4110 (N_4110,In_2692,In_4079);
nor U4111 (N_4111,In_1701,In_3788);
and U4112 (N_4112,In_680,In_3585);
and U4113 (N_4113,In_3873,In_4616);
and U4114 (N_4114,In_2838,In_997);
xnor U4115 (N_4115,In_60,In_1464);
and U4116 (N_4116,In_4096,In_895);
and U4117 (N_4117,In_1919,In_311);
and U4118 (N_4118,In_116,In_184);
or U4119 (N_4119,In_1404,In_2633);
nand U4120 (N_4120,In_4502,In_4852);
nor U4121 (N_4121,In_1143,In_2816);
and U4122 (N_4122,In_4028,In_4233);
or U4123 (N_4123,In_1160,In_2289);
or U4124 (N_4124,In_4306,In_3741);
and U4125 (N_4125,In_3267,In_2480);
xnor U4126 (N_4126,In_3748,In_780);
and U4127 (N_4127,In_1747,In_3799);
nor U4128 (N_4128,In_862,In_1873);
nor U4129 (N_4129,In_51,In_2851);
xnor U4130 (N_4130,In_2331,In_138);
nor U4131 (N_4131,In_2240,In_2951);
nand U4132 (N_4132,In_855,In_4136);
or U4133 (N_4133,In_3357,In_1232);
nand U4134 (N_4134,In_2564,In_1474);
or U4135 (N_4135,In_1004,In_3207);
xnor U4136 (N_4136,In_1323,In_1856);
or U4137 (N_4137,In_3799,In_2231);
xor U4138 (N_4138,In_3261,In_1476);
nand U4139 (N_4139,In_1558,In_482);
nand U4140 (N_4140,In_3217,In_3206);
nand U4141 (N_4141,In_3744,In_4497);
xnor U4142 (N_4142,In_4704,In_3149);
or U4143 (N_4143,In_1727,In_3066);
nand U4144 (N_4144,In_2776,In_3519);
or U4145 (N_4145,In_2246,In_1825);
nand U4146 (N_4146,In_469,In_4962);
nor U4147 (N_4147,In_873,In_2407);
and U4148 (N_4148,In_3305,In_1710);
or U4149 (N_4149,In_1014,In_3312);
xor U4150 (N_4150,In_98,In_3908);
xor U4151 (N_4151,In_1610,In_324);
and U4152 (N_4152,In_139,In_448);
or U4153 (N_4153,In_240,In_574);
nor U4154 (N_4154,In_2902,In_4575);
nor U4155 (N_4155,In_371,In_1339);
xor U4156 (N_4156,In_4463,In_3275);
nand U4157 (N_4157,In_3961,In_3184);
or U4158 (N_4158,In_3605,In_3146);
nor U4159 (N_4159,In_3423,In_2153);
nand U4160 (N_4160,In_439,In_3264);
or U4161 (N_4161,In_4007,In_256);
nor U4162 (N_4162,In_1770,In_493);
nor U4163 (N_4163,In_2554,In_2065);
nor U4164 (N_4164,In_1044,In_2578);
nor U4165 (N_4165,In_2736,In_3489);
xor U4166 (N_4166,In_2988,In_206);
or U4167 (N_4167,In_1487,In_3285);
or U4168 (N_4168,In_182,In_669);
or U4169 (N_4169,In_3634,In_1796);
nor U4170 (N_4170,In_1155,In_4735);
nand U4171 (N_4171,In_3061,In_1553);
xnor U4172 (N_4172,In_2594,In_1679);
nand U4173 (N_4173,In_4650,In_4085);
nand U4174 (N_4174,In_2111,In_1498);
nand U4175 (N_4175,In_3898,In_4415);
and U4176 (N_4176,In_2711,In_4893);
nor U4177 (N_4177,In_4431,In_1898);
nand U4178 (N_4178,In_3997,In_216);
nor U4179 (N_4179,In_2567,In_4221);
and U4180 (N_4180,In_876,In_1474);
and U4181 (N_4181,In_1208,In_15);
and U4182 (N_4182,In_369,In_4780);
nand U4183 (N_4183,In_388,In_1974);
xnor U4184 (N_4184,In_2108,In_243);
and U4185 (N_4185,In_133,In_1932);
and U4186 (N_4186,In_2350,In_3252);
and U4187 (N_4187,In_4888,In_2391);
xor U4188 (N_4188,In_3300,In_2033);
and U4189 (N_4189,In_3779,In_4006);
nor U4190 (N_4190,In_3060,In_3412);
and U4191 (N_4191,In_1589,In_4224);
nand U4192 (N_4192,In_3049,In_1937);
nor U4193 (N_4193,In_3522,In_2494);
or U4194 (N_4194,In_2897,In_4081);
or U4195 (N_4195,In_2610,In_2268);
xor U4196 (N_4196,In_1817,In_4462);
nand U4197 (N_4197,In_1702,In_1075);
xor U4198 (N_4198,In_2176,In_3091);
nor U4199 (N_4199,In_2059,In_4023);
or U4200 (N_4200,In_1753,In_3104);
or U4201 (N_4201,In_4590,In_4390);
and U4202 (N_4202,In_1997,In_3935);
and U4203 (N_4203,In_3284,In_2684);
nand U4204 (N_4204,In_408,In_2039);
or U4205 (N_4205,In_2768,In_32);
nor U4206 (N_4206,In_2308,In_4140);
xor U4207 (N_4207,In_2020,In_3127);
or U4208 (N_4208,In_3762,In_1295);
and U4209 (N_4209,In_4601,In_1779);
nand U4210 (N_4210,In_2982,In_2668);
nand U4211 (N_4211,In_3580,In_2342);
nand U4212 (N_4212,In_1876,In_4986);
and U4213 (N_4213,In_2097,In_1186);
and U4214 (N_4214,In_1747,In_3486);
nor U4215 (N_4215,In_1565,In_4437);
and U4216 (N_4216,In_820,In_3063);
xor U4217 (N_4217,In_3759,In_1030);
or U4218 (N_4218,In_2371,In_3311);
and U4219 (N_4219,In_4956,In_3929);
or U4220 (N_4220,In_4638,In_4428);
or U4221 (N_4221,In_4128,In_4510);
nand U4222 (N_4222,In_139,In_4836);
xnor U4223 (N_4223,In_4354,In_510);
xnor U4224 (N_4224,In_2320,In_3528);
and U4225 (N_4225,In_2511,In_2842);
nor U4226 (N_4226,In_4001,In_494);
nor U4227 (N_4227,In_730,In_4204);
nand U4228 (N_4228,In_1582,In_2418);
nor U4229 (N_4229,In_4820,In_2461);
nand U4230 (N_4230,In_1585,In_4221);
nand U4231 (N_4231,In_813,In_3740);
or U4232 (N_4232,In_3458,In_3344);
xor U4233 (N_4233,In_1153,In_676);
or U4234 (N_4234,In_4504,In_917);
nand U4235 (N_4235,In_4357,In_3033);
or U4236 (N_4236,In_2247,In_387);
nand U4237 (N_4237,In_2397,In_4546);
nor U4238 (N_4238,In_4017,In_1706);
or U4239 (N_4239,In_2363,In_3253);
nor U4240 (N_4240,In_1793,In_2447);
and U4241 (N_4241,In_539,In_3869);
or U4242 (N_4242,In_4835,In_2768);
nand U4243 (N_4243,In_574,In_2219);
nor U4244 (N_4244,In_4755,In_4644);
or U4245 (N_4245,In_3991,In_4293);
xor U4246 (N_4246,In_3273,In_2890);
and U4247 (N_4247,In_4959,In_403);
or U4248 (N_4248,In_4701,In_3379);
or U4249 (N_4249,In_3280,In_1981);
nor U4250 (N_4250,In_964,In_923);
xnor U4251 (N_4251,In_4254,In_2493);
nor U4252 (N_4252,In_2518,In_3406);
or U4253 (N_4253,In_3567,In_2238);
nor U4254 (N_4254,In_2922,In_5);
or U4255 (N_4255,In_1967,In_1938);
and U4256 (N_4256,In_3706,In_2184);
and U4257 (N_4257,In_3364,In_1536);
nand U4258 (N_4258,In_1445,In_1863);
xor U4259 (N_4259,In_3163,In_4629);
nor U4260 (N_4260,In_3034,In_3026);
or U4261 (N_4261,In_1858,In_1981);
and U4262 (N_4262,In_2612,In_2846);
nor U4263 (N_4263,In_4613,In_1639);
or U4264 (N_4264,In_4292,In_2503);
and U4265 (N_4265,In_1827,In_240);
xnor U4266 (N_4266,In_862,In_1217);
nor U4267 (N_4267,In_3867,In_628);
nand U4268 (N_4268,In_1461,In_2402);
nand U4269 (N_4269,In_1044,In_956);
nor U4270 (N_4270,In_3476,In_4022);
or U4271 (N_4271,In_629,In_2562);
nand U4272 (N_4272,In_4204,In_2739);
and U4273 (N_4273,In_2087,In_697);
nand U4274 (N_4274,In_4588,In_1363);
xor U4275 (N_4275,In_2604,In_555);
or U4276 (N_4276,In_3836,In_3457);
and U4277 (N_4277,In_2489,In_2630);
and U4278 (N_4278,In_4758,In_3929);
xnor U4279 (N_4279,In_865,In_4923);
and U4280 (N_4280,In_1379,In_3421);
and U4281 (N_4281,In_3818,In_3412);
xor U4282 (N_4282,In_616,In_3828);
nor U4283 (N_4283,In_4450,In_4405);
or U4284 (N_4284,In_2967,In_2404);
nor U4285 (N_4285,In_3802,In_101);
nand U4286 (N_4286,In_4559,In_1406);
and U4287 (N_4287,In_3458,In_180);
nand U4288 (N_4288,In_165,In_614);
nand U4289 (N_4289,In_548,In_379);
xor U4290 (N_4290,In_3373,In_2224);
nand U4291 (N_4291,In_2625,In_1637);
xor U4292 (N_4292,In_2524,In_60);
xor U4293 (N_4293,In_3554,In_3024);
nand U4294 (N_4294,In_4903,In_3021);
and U4295 (N_4295,In_4418,In_22);
nor U4296 (N_4296,In_272,In_1457);
nor U4297 (N_4297,In_3387,In_3327);
nand U4298 (N_4298,In_2774,In_929);
xnor U4299 (N_4299,In_3168,In_1041);
xor U4300 (N_4300,In_1469,In_2503);
nor U4301 (N_4301,In_1940,In_4455);
nand U4302 (N_4302,In_3368,In_4481);
or U4303 (N_4303,In_3998,In_3642);
and U4304 (N_4304,In_2485,In_526);
xor U4305 (N_4305,In_2265,In_3578);
nor U4306 (N_4306,In_1538,In_2266);
and U4307 (N_4307,In_1038,In_1772);
nand U4308 (N_4308,In_2995,In_3575);
xnor U4309 (N_4309,In_2814,In_372);
and U4310 (N_4310,In_3148,In_4398);
xnor U4311 (N_4311,In_4715,In_3733);
or U4312 (N_4312,In_3209,In_2510);
nor U4313 (N_4313,In_2224,In_4252);
or U4314 (N_4314,In_3476,In_1632);
xnor U4315 (N_4315,In_4491,In_3761);
nor U4316 (N_4316,In_832,In_224);
or U4317 (N_4317,In_1322,In_1214);
nor U4318 (N_4318,In_819,In_3664);
xnor U4319 (N_4319,In_3786,In_302);
and U4320 (N_4320,In_173,In_3246);
nand U4321 (N_4321,In_1196,In_4480);
nand U4322 (N_4322,In_344,In_4818);
nand U4323 (N_4323,In_4019,In_1313);
nand U4324 (N_4324,In_1387,In_3522);
nand U4325 (N_4325,In_3223,In_480);
nand U4326 (N_4326,In_1913,In_963);
xor U4327 (N_4327,In_3637,In_4985);
xor U4328 (N_4328,In_2425,In_4501);
or U4329 (N_4329,In_2071,In_1362);
and U4330 (N_4330,In_1686,In_1354);
nand U4331 (N_4331,In_3192,In_2030);
and U4332 (N_4332,In_3430,In_3130);
nor U4333 (N_4333,In_2177,In_4474);
xnor U4334 (N_4334,In_959,In_3940);
nor U4335 (N_4335,In_406,In_1442);
or U4336 (N_4336,In_4973,In_3685);
nor U4337 (N_4337,In_2824,In_4806);
nand U4338 (N_4338,In_4264,In_3990);
or U4339 (N_4339,In_2941,In_2455);
and U4340 (N_4340,In_1745,In_4644);
or U4341 (N_4341,In_4733,In_1033);
xor U4342 (N_4342,In_112,In_2406);
or U4343 (N_4343,In_3970,In_4108);
xnor U4344 (N_4344,In_4559,In_3205);
xnor U4345 (N_4345,In_4269,In_3929);
xnor U4346 (N_4346,In_3452,In_2761);
or U4347 (N_4347,In_4718,In_4885);
nand U4348 (N_4348,In_2478,In_1959);
or U4349 (N_4349,In_3413,In_1358);
nor U4350 (N_4350,In_2142,In_2766);
xor U4351 (N_4351,In_709,In_1581);
and U4352 (N_4352,In_1947,In_1698);
nor U4353 (N_4353,In_2857,In_1648);
nor U4354 (N_4354,In_561,In_4668);
nand U4355 (N_4355,In_2502,In_4401);
nand U4356 (N_4356,In_4297,In_3934);
or U4357 (N_4357,In_4682,In_661);
and U4358 (N_4358,In_4345,In_712);
nor U4359 (N_4359,In_561,In_1563);
nand U4360 (N_4360,In_507,In_280);
or U4361 (N_4361,In_3192,In_788);
nand U4362 (N_4362,In_1554,In_3247);
nor U4363 (N_4363,In_4369,In_4236);
nor U4364 (N_4364,In_3537,In_4208);
nor U4365 (N_4365,In_2991,In_696);
nand U4366 (N_4366,In_563,In_4996);
nor U4367 (N_4367,In_2451,In_1359);
and U4368 (N_4368,In_1664,In_292);
or U4369 (N_4369,In_2251,In_4120);
xnor U4370 (N_4370,In_4160,In_244);
nand U4371 (N_4371,In_4931,In_3357);
xnor U4372 (N_4372,In_4895,In_4324);
and U4373 (N_4373,In_2247,In_2489);
xor U4374 (N_4374,In_1232,In_3921);
or U4375 (N_4375,In_3381,In_3779);
or U4376 (N_4376,In_2437,In_2608);
xnor U4377 (N_4377,In_4729,In_1837);
xor U4378 (N_4378,In_3447,In_1319);
nor U4379 (N_4379,In_1570,In_3263);
or U4380 (N_4380,In_1668,In_1280);
nand U4381 (N_4381,In_336,In_1600);
xor U4382 (N_4382,In_4611,In_129);
nor U4383 (N_4383,In_4741,In_407);
and U4384 (N_4384,In_53,In_2134);
or U4385 (N_4385,In_4784,In_2409);
nand U4386 (N_4386,In_2934,In_1762);
xor U4387 (N_4387,In_3378,In_485);
nor U4388 (N_4388,In_3643,In_1974);
and U4389 (N_4389,In_3282,In_2549);
and U4390 (N_4390,In_1865,In_3750);
or U4391 (N_4391,In_2107,In_4000);
xnor U4392 (N_4392,In_1705,In_4725);
xnor U4393 (N_4393,In_3389,In_2713);
nor U4394 (N_4394,In_887,In_3936);
nand U4395 (N_4395,In_3944,In_3826);
or U4396 (N_4396,In_631,In_2697);
nand U4397 (N_4397,In_3016,In_445);
or U4398 (N_4398,In_3529,In_2238);
nand U4399 (N_4399,In_3710,In_3220);
nand U4400 (N_4400,In_4407,In_1221);
or U4401 (N_4401,In_3646,In_4755);
and U4402 (N_4402,In_211,In_1384);
nand U4403 (N_4403,In_1063,In_380);
xor U4404 (N_4404,In_2485,In_4088);
xnor U4405 (N_4405,In_1465,In_3499);
nand U4406 (N_4406,In_4344,In_509);
and U4407 (N_4407,In_206,In_4589);
nand U4408 (N_4408,In_1974,In_4278);
nand U4409 (N_4409,In_4989,In_446);
xnor U4410 (N_4410,In_2841,In_1241);
or U4411 (N_4411,In_3539,In_2920);
and U4412 (N_4412,In_804,In_956);
nand U4413 (N_4413,In_3931,In_4641);
or U4414 (N_4414,In_4944,In_367);
xnor U4415 (N_4415,In_3966,In_4276);
xnor U4416 (N_4416,In_3214,In_513);
nor U4417 (N_4417,In_4354,In_4878);
nor U4418 (N_4418,In_2451,In_2340);
nand U4419 (N_4419,In_3680,In_3489);
xnor U4420 (N_4420,In_3571,In_774);
nor U4421 (N_4421,In_2191,In_2716);
xnor U4422 (N_4422,In_1447,In_4186);
nand U4423 (N_4423,In_809,In_3049);
xnor U4424 (N_4424,In_1457,In_2491);
xor U4425 (N_4425,In_2359,In_2973);
nand U4426 (N_4426,In_4000,In_3692);
nor U4427 (N_4427,In_3133,In_2962);
and U4428 (N_4428,In_4144,In_1757);
nand U4429 (N_4429,In_3672,In_2182);
and U4430 (N_4430,In_970,In_1746);
and U4431 (N_4431,In_673,In_3766);
and U4432 (N_4432,In_1372,In_2773);
nor U4433 (N_4433,In_1482,In_1965);
xnor U4434 (N_4434,In_1179,In_3535);
xor U4435 (N_4435,In_4334,In_347);
or U4436 (N_4436,In_262,In_1043);
xor U4437 (N_4437,In_3323,In_3202);
xnor U4438 (N_4438,In_1062,In_4446);
xnor U4439 (N_4439,In_26,In_2847);
xnor U4440 (N_4440,In_259,In_471);
or U4441 (N_4441,In_2212,In_4651);
and U4442 (N_4442,In_4076,In_1473);
and U4443 (N_4443,In_676,In_1219);
xnor U4444 (N_4444,In_2763,In_2499);
and U4445 (N_4445,In_4119,In_135);
or U4446 (N_4446,In_4160,In_3783);
nor U4447 (N_4447,In_292,In_67);
nor U4448 (N_4448,In_817,In_189);
xor U4449 (N_4449,In_1741,In_1789);
or U4450 (N_4450,In_4854,In_1623);
and U4451 (N_4451,In_3384,In_2163);
or U4452 (N_4452,In_842,In_790);
nand U4453 (N_4453,In_2676,In_4561);
nand U4454 (N_4454,In_3448,In_1201);
nor U4455 (N_4455,In_2490,In_342);
xnor U4456 (N_4456,In_3642,In_182);
nand U4457 (N_4457,In_3091,In_3232);
xor U4458 (N_4458,In_1404,In_259);
or U4459 (N_4459,In_1839,In_1797);
nor U4460 (N_4460,In_2410,In_2576);
nor U4461 (N_4461,In_1203,In_1435);
or U4462 (N_4462,In_2441,In_2393);
and U4463 (N_4463,In_1146,In_2668);
nor U4464 (N_4464,In_365,In_335);
nor U4465 (N_4465,In_140,In_1893);
xor U4466 (N_4466,In_418,In_268);
or U4467 (N_4467,In_1985,In_3408);
xor U4468 (N_4468,In_3860,In_685);
nor U4469 (N_4469,In_516,In_1481);
and U4470 (N_4470,In_16,In_978);
or U4471 (N_4471,In_2904,In_1571);
and U4472 (N_4472,In_2912,In_4332);
nor U4473 (N_4473,In_2696,In_3183);
or U4474 (N_4474,In_2143,In_72);
and U4475 (N_4475,In_461,In_818);
nand U4476 (N_4476,In_2212,In_851);
or U4477 (N_4477,In_3614,In_2113);
nor U4478 (N_4478,In_2625,In_1865);
nor U4479 (N_4479,In_4280,In_2657);
xnor U4480 (N_4480,In_4198,In_2662);
or U4481 (N_4481,In_4759,In_2985);
or U4482 (N_4482,In_4411,In_1535);
and U4483 (N_4483,In_4798,In_1717);
nand U4484 (N_4484,In_1912,In_440);
nor U4485 (N_4485,In_2936,In_1225);
or U4486 (N_4486,In_2274,In_2063);
and U4487 (N_4487,In_3439,In_4301);
nand U4488 (N_4488,In_2205,In_3114);
nand U4489 (N_4489,In_2018,In_2037);
nor U4490 (N_4490,In_3681,In_260);
nor U4491 (N_4491,In_4973,In_932);
xnor U4492 (N_4492,In_3476,In_4905);
or U4493 (N_4493,In_2989,In_4525);
or U4494 (N_4494,In_300,In_2541);
or U4495 (N_4495,In_452,In_2410);
xnor U4496 (N_4496,In_3240,In_1097);
or U4497 (N_4497,In_4228,In_3616);
or U4498 (N_4498,In_982,In_1418);
nor U4499 (N_4499,In_4068,In_3306);
or U4500 (N_4500,In_136,In_415);
and U4501 (N_4501,In_974,In_99);
xnor U4502 (N_4502,In_769,In_109);
or U4503 (N_4503,In_3595,In_1996);
xnor U4504 (N_4504,In_4409,In_3516);
nand U4505 (N_4505,In_4951,In_2427);
nor U4506 (N_4506,In_2727,In_2680);
xnor U4507 (N_4507,In_3224,In_3063);
and U4508 (N_4508,In_2736,In_4485);
nand U4509 (N_4509,In_4815,In_3107);
or U4510 (N_4510,In_3526,In_2998);
xnor U4511 (N_4511,In_4579,In_493);
xnor U4512 (N_4512,In_2449,In_1174);
xor U4513 (N_4513,In_1490,In_293);
nand U4514 (N_4514,In_4531,In_3596);
and U4515 (N_4515,In_631,In_2530);
and U4516 (N_4516,In_4760,In_1548);
xor U4517 (N_4517,In_963,In_3064);
xnor U4518 (N_4518,In_2493,In_3228);
nor U4519 (N_4519,In_3924,In_3016);
and U4520 (N_4520,In_4676,In_1327);
nand U4521 (N_4521,In_2696,In_1339);
xnor U4522 (N_4522,In_3014,In_3294);
nor U4523 (N_4523,In_3006,In_4461);
xnor U4524 (N_4524,In_1828,In_22);
nand U4525 (N_4525,In_1954,In_2855);
or U4526 (N_4526,In_4633,In_45);
xnor U4527 (N_4527,In_4704,In_1716);
or U4528 (N_4528,In_818,In_2615);
nand U4529 (N_4529,In_1480,In_2679);
xnor U4530 (N_4530,In_3884,In_2097);
or U4531 (N_4531,In_792,In_4463);
xnor U4532 (N_4532,In_4722,In_3619);
nor U4533 (N_4533,In_4422,In_4919);
or U4534 (N_4534,In_1240,In_502);
xor U4535 (N_4535,In_3356,In_3873);
xnor U4536 (N_4536,In_1137,In_1540);
nand U4537 (N_4537,In_3691,In_2708);
xor U4538 (N_4538,In_224,In_2650);
xor U4539 (N_4539,In_4373,In_4568);
or U4540 (N_4540,In_1770,In_4885);
xnor U4541 (N_4541,In_4256,In_273);
and U4542 (N_4542,In_3506,In_3067);
nand U4543 (N_4543,In_3611,In_4076);
and U4544 (N_4544,In_4595,In_3639);
nor U4545 (N_4545,In_804,In_2286);
or U4546 (N_4546,In_3412,In_4877);
or U4547 (N_4547,In_1300,In_1402);
nor U4548 (N_4548,In_328,In_1778);
nor U4549 (N_4549,In_4592,In_2840);
nand U4550 (N_4550,In_2178,In_3804);
and U4551 (N_4551,In_4647,In_4318);
and U4552 (N_4552,In_3632,In_2384);
nor U4553 (N_4553,In_4037,In_1734);
xnor U4554 (N_4554,In_2935,In_39);
xnor U4555 (N_4555,In_937,In_1883);
xor U4556 (N_4556,In_4820,In_4478);
nand U4557 (N_4557,In_1279,In_12);
nor U4558 (N_4558,In_2794,In_1713);
or U4559 (N_4559,In_3766,In_465);
and U4560 (N_4560,In_1732,In_426);
nor U4561 (N_4561,In_565,In_2645);
nor U4562 (N_4562,In_2102,In_781);
and U4563 (N_4563,In_474,In_2379);
xor U4564 (N_4564,In_68,In_4204);
nand U4565 (N_4565,In_2399,In_2667);
or U4566 (N_4566,In_991,In_1675);
xor U4567 (N_4567,In_622,In_2211);
and U4568 (N_4568,In_2786,In_3924);
and U4569 (N_4569,In_1958,In_2536);
nor U4570 (N_4570,In_4858,In_2116);
and U4571 (N_4571,In_692,In_2773);
or U4572 (N_4572,In_3594,In_2391);
xor U4573 (N_4573,In_4596,In_4272);
nand U4574 (N_4574,In_2463,In_760);
and U4575 (N_4575,In_122,In_2149);
or U4576 (N_4576,In_2916,In_3757);
xnor U4577 (N_4577,In_1088,In_4342);
nor U4578 (N_4578,In_789,In_2540);
xor U4579 (N_4579,In_1997,In_147);
and U4580 (N_4580,In_44,In_387);
nor U4581 (N_4581,In_2072,In_3391);
xor U4582 (N_4582,In_2798,In_2247);
or U4583 (N_4583,In_500,In_3473);
and U4584 (N_4584,In_4233,In_2387);
or U4585 (N_4585,In_10,In_438);
xor U4586 (N_4586,In_1292,In_3752);
or U4587 (N_4587,In_2262,In_3464);
and U4588 (N_4588,In_865,In_1919);
and U4589 (N_4589,In_4489,In_3534);
nand U4590 (N_4590,In_4989,In_1208);
or U4591 (N_4591,In_3728,In_1603);
and U4592 (N_4592,In_114,In_2146);
and U4593 (N_4593,In_1221,In_3448);
and U4594 (N_4594,In_4847,In_27);
xnor U4595 (N_4595,In_976,In_2324);
xor U4596 (N_4596,In_2993,In_3990);
nor U4597 (N_4597,In_3550,In_3176);
nand U4598 (N_4598,In_4733,In_2886);
xor U4599 (N_4599,In_2782,In_1573);
nand U4600 (N_4600,In_1811,In_628);
or U4601 (N_4601,In_4584,In_2471);
nor U4602 (N_4602,In_3972,In_3958);
and U4603 (N_4603,In_24,In_3697);
nand U4604 (N_4604,In_1243,In_2795);
nand U4605 (N_4605,In_4067,In_3751);
or U4606 (N_4606,In_2758,In_1436);
nand U4607 (N_4607,In_2827,In_3321);
and U4608 (N_4608,In_2431,In_2715);
xnor U4609 (N_4609,In_2597,In_1832);
nand U4610 (N_4610,In_16,In_1156);
xor U4611 (N_4611,In_2750,In_4756);
nand U4612 (N_4612,In_2954,In_100);
and U4613 (N_4613,In_4395,In_3395);
or U4614 (N_4614,In_3829,In_1518);
nand U4615 (N_4615,In_3978,In_2498);
nand U4616 (N_4616,In_377,In_3948);
nor U4617 (N_4617,In_2891,In_1185);
and U4618 (N_4618,In_1989,In_728);
and U4619 (N_4619,In_3682,In_571);
nor U4620 (N_4620,In_1816,In_1315);
or U4621 (N_4621,In_2103,In_4772);
and U4622 (N_4622,In_4440,In_3797);
xor U4623 (N_4623,In_1204,In_4418);
xnor U4624 (N_4624,In_1261,In_399);
nor U4625 (N_4625,In_155,In_174);
and U4626 (N_4626,In_1610,In_227);
and U4627 (N_4627,In_1406,In_3429);
or U4628 (N_4628,In_286,In_4129);
xor U4629 (N_4629,In_3168,In_3809);
and U4630 (N_4630,In_4010,In_4234);
nand U4631 (N_4631,In_190,In_3275);
nor U4632 (N_4632,In_2848,In_4049);
or U4633 (N_4633,In_4074,In_1580);
xor U4634 (N_4634,In_3245,In_2159);
or U4635 (N_4635,In_4447,In_4771);
xor U4636 (N_4636,In_2804,In_3431);
nand U4637 (N_4637,In_974,In_4097);
and U4638 (N_4638,In_3229,In_3726);
xor U4639 (N_4639,In_3172,In_633);
nor U4640 (N_4640,In_25,In_4978);
xor U4641 (N_4641,In_1489,In_3209);
and U4642 (N_4642,In_1117,In_4660);
or U4643 (N_4643,In_2650,In_3330);
and U4644 (N_4644,In_2289,In_2401);
or U4645 (N_4645,In_2624,In_3541);
or U4646 (N_4646,In_4478,In_4341);
nor U4647 (N_4647,In_4206,In_3085);
nand U4648 (N_4648,In_3785,In_2288);
and U4649 (N_4649,In_112,In_3191);
and U4650 (N_4650,In_3520,In_783);
xor U4651 (N_4651,In_0,In_4177);
or U4652 (N_4652,In_63,In_4272);
or U4653 (N_4653,In_4996,In_4277);
nand U4654 (N_4654,In_3177,In_4971);
or U4655 (N_4655,In_192,In_40);
xnor U4656 (N_4656,In_3746,In_2723);
xor U4657 (N_4657,In_2614,In_639);
and U4658 (N_4658,In_1577,In_3754);
nand U4659 (N_4659,In_4847,In_244);
nor U4660 (N_4660,In_1597,In_2072);
nand U4661 (N_4661,In_3629,In_3118);
or U4662 (N_4662,In_1653,In_4987);
and U4663 (N_4663,In_2509,In_4296);
and U4664 (N_4664,In_2273,In_4377);
and U4665 (N_4665,In_2996,In_501);
xnor U4666 (N_4666,In_1910,In_605);
and U4667 (N_4667,In_2432,In_430);
nor U4668 (N_4668,In_2436,In_4129);
and U4669 (N_4669,In_3013,In_4542);
xor U4670 (N_4670,In_4994,In_3331);
or U4671 (N_4671,In_4001,In_3981);
xor U4672 (N_4672,In_3040,In_4669);
or U4673 (N_4673,In_3354,In_349);
and U4674 (N_4674,In_3107,In_1255);
or U4675 (N_4675,In_1568,In_3408);
or U4676 (N_4676,In_2785,In_995);
nor U4677 (N_4677,In_4725,In_78);
nor U4678 (N_4678,In_333,In_3299);
or U4679 (N_4679,In_2802,In_4941);
nand U4680 (N_4680,In_745,In_3646);
nor U4681 (N_4681,In_2429,In_1058);
xnor U4682 (N_4682,In_884,In_4833);
or U4683 (N_4683,In_4972,In_4607);
xnor U4684 (N_4684,In_2818,In_3434);
and U4685 (N_4685,In_884,In_2487);
nor U4686 (N_4686,In_1519,In_2589);
xor U4687 (N_4687,In_3000,In_3818);
and U4688 (N_4688,In_771,In_2098);
xnor U4689 (N_4689,In_1071,In_2450);
nand U4690 (N_4690,In_3260,In_4123);
nand U4691 (N_4691,In_2800,In_1991);
nand U4692 (N_4692,In_4539,In_2248);
nor U4693 (N_4693,In_2423,In_3898);
and U4694 (N_4694,In_4604,In_670);
nand U4695 (N_4695,In_3215,In_906);
and U4696 (N_4696,In_4376,In_4334);
xnor U4697 (N_4697,In_2270,In_4885);
nor U4698 (N_4698,In_4616,In_256);
or U4699 (N_4699,In_73,In_4120);
nand U4700 (N_4700,In_466,In_1804);
nor U4701 (N_4701,In_1953,In_379);
and U4702 (N_4702,In_330,In_1302);
or U4703 (N_4703,In_2874,In_2746);
nor U4704 (N_4704,In_3767,In_250);
xor U4705 (N_4705,In_2625,In_2916);
and U4706 (N_4706,In_3032,In_2405);
and U4707 (N_4707,In_4575,In_1977);
nor U4708 (N_4708,In_3465,In_2124);
nand U4709 (N_4709,In_4473,In_2087);
nand U4710 (N_4710,In_4123,In_4353);
or U4711 (N_4711,In_232,In_1692);
xnor U4712 (N_4712,In_174,In_3992);
and U4713 (N_4713,In_2985,In_1073);
xor U4714 (N_4714,In_3298,In_4912);
xor U4715 (N_4715,In_755,In_174);
nand U4716 (N_4716,In_2434,In_4993);
nor U4717 (N_4717,In_2870,In_965);
nor U4718 (N_4718,In_2688,In_4708);
or U4719 (N_4719,In_4635,In_1835);
nor U4720 (N_4720,In_2234,In_4631);
xnor U4721 (N_4721,In_1764,In_3545);
nor U4722 (N_4722,In_2310,In_3733);
nand U4723 (N_4723,In_538,In_1926);
nor U4724 (N_4724,In_4033,In_504);
nand U4725 (N_4725,In_4986,In_4218);
and U4726 (N_4726,In_1730,In_1227);
or U4727 (N_4727,In_2760,In_4729);
or U4728 (N_4728,In_7,In_2620);
and U4729 (N_4729,In_3584,In_3657);
nor U4730 (N_4730,In_2495,In_3032);
nor U4731 (N_4731,In_2292,In_1902);
nand U4732 (N_4732,In_1313,In_2014);
or U4733 (N_4733,In_1243,In_3492);
nand U4734 (N_4734,In_2865,In_552);
nor U4735 (N_4735,In_1456,In_2415);
or U4736 (N_4736,In_1837,In_2718);
and U4737 (N_4737,In_734,In_702);
nand U4738 (N_4738,In_4632,In_4008);
nand U4739 (N_4739,In_1196,In_1337);
nand U4740 (N_4740,In_1023,In_1707);
nand U4741 (N_4741,In_2600,In_4621);
nand U4742 (N_4742,In_2619,In_2632);
or U4743 (N_4743,In_1648,In_1799);
nand U4744 (N_4744,In_2308,In_4612);
nand U4745 (N_4745,In_4020,In_3424);
nand U4746 (N_4746,In_1959,In_4238);
nand U4747 (N_4747,In_169,In_842);
xnor U4748 (N_4748,In_3740,In_3361);
xor U4749 (N_4749,In_4255,In_4091);
xnor U4750 (N_4750,In_545,In_900);
nand U4751 (N_4751,In_1793,In_4837);
nand U4752 (N_4752,In_1923,In_2796);
xnor U4753 (N_4753,In_3257,In_1885);
or U4754 (N_4754,In_2109,In_581);
xnor U4755 (N_4755,In_450,In_39);
xnor U4756 (N_4756,In_1685,In_19);
or U4757 (N_4757,In_1879,In_2771);
nand U4758 (N_4758,In_2820,In_668);
xor U4759 (N_4759,In_1602,In_148);
or U4760 (N_4760,In_264,In_995);
and U4761 (N_4761,In_248,In_4756);
xor U4762 (N_4762,In_278,In_3073);
nand U4763 (N_4763,In_2580,In_722);
or U4764 (N_4764,In_3069,In_2332);
and U4765 (N_4765,In_3249,In_3539);
nand U4766 (N_4766,In_2905,In_2050);
or U4767 (N_4767,In_1876,In_2646);
or U4768 (N_4768,In_2536,In_3220);
or U4769 (N_4769,In_4129,In_4506);
or U4770 (N_4770,In_362,In_3924);
or U4771 (N_4771,In_2639,In_1929);
nor U4772 (N_4772,In_3738,In_4799);
nor U4773 (N_4773,In_3483,In_3338);
nor U4774 (N_4774,In_2456,In_1140);
xnor U4775 (N_4775,In_2798,In_4952);
or U4776 (N_4776,In_1958,In_487);
or U4777 (N_4777,In_3248,In_4446);
or U4778 (N_4778,In_3596,In_2892);
or U4779 (N_4779,In_74,In_212);
or U4780 (N_4780,In_969,In_4188);
or U4781 (N_4781,In_4885,In_2955);
nor U4782 (N_4782,In_2290,In_1327);
nor U4783 (N_4783,In_4202,In_1997);
nand U4784 (N_4784,In_954,In_2509);
nor U4785 (N_4785,In_3570,In_3664);
or U4786 (N_4786,In_4039,In_1236);
xor U4787 (N_4787,In_1131,In_3296);
or U4788 (N_4788,In_4522,In_902);
nand U4789 (N_4789,In_1239,In_1331);
xnor U4790 (N_4790,In_2781,In_4093);
nor U4791 (N_4791,In_4475,In_1088);
nor U4792 (N_4792,In_4391,In_3014);
and U4793 (N_4793,In_4279,In_1881);
xnor U4794 (N_4794,In_464,In_4225);
xnor U4795 (N_4795,In_626,In_2605);
nand U4796 (N_4796,In_1563,In_1168);
nor U4797 (N_4797,In_1921,In_2725);
nand U4798 (N_4798,In_2386,In_612);
nand U4799 (N_4799,In_181,In_2958);
xor U4800 (N_4800,In_1676,In_4290);
xnor U4801 (N_4801,In_3877,In_2918);
xnor U4802 (N_4802,In_3067,In_2654);
and U4803 (N_4803,In_685,In_3946);
nor U4804 (N_4804,In_2654,In_2325);
xnor U4805 (N_4805,In_2445,In_296);
nand U4806 (N_4806,In_1112,In_797);
and U4807 (N_4807,In_936,In_4444);
nor U4808 (N_4808,In_2687,In_67);
nor U4809 (N_4809,In_2792,In_4668);
xor U4810 (N_4810,In_2518,In_2394);
xor U4811 (N_4811,In_3928,In_1557);
and U4812 (N_4812,In_4492,In_1210);
and U4813 (N_4813,In_1879,In_3306);
or U4814 (N_4814,In_4751,In_801);
or U4815 (N_4815,In_1245,In_4678);
nand U4816 (N_4816,In_4110,In_2057);
nor U4817 (N_4817,In_1293,In_1830);
and U4818 (N_4818,In_3520,In_642);
nand U4819 (N_4819,In_1301,In_4245);
nand U4820 (N_4820,In_764,In_74);
and U4821 (N_4821,In_3958,In_2877);
or U4822 (N_4822,In_2013,In_3574);
nor U4823 (N_4823,In_1599,In_2802);
or U4824 (N_4824,In_1950,In_2324);
and U4825 (N_4825,In_2729,In_85);
xor U4826 (N_4826,In_1704,In_181);
xnor U4827 (N_4827,In_4073,In_4107);
nand U4828 (N_4828,In_3463,In_2895);
xnor U4829 (N_4829,In_4300,In_3092);
nand U4830 (N_4830,In_1750,In_876);
nor U4831 (N_4831,In_1255,In_3048);
or U4832 (N_4832,In_1016,In_516);
nand U4833 (N_4833,In_247,In_4500);
and U4834 (N_4834,In_3290,In_1279);
nand U4835 (N_4835,In_1956,In_4525);
nor U4836 (N_4836,In_4056,In_1855);
and U4837 (N_4837,In_3510,In_4308);
xor U4838 (N_4838,In_810,In_4560);
xor U4839 (N_4839,In_4113,In_4597);
xor U4840 (N_4840,In_2743,In_1670);
nor U4841 (N_4841,In_4635,In_1852);
xor U4842 (N_4842,In_262,In_3422);
nand U4843 (N_4843,In_1541,In_4096);
or U4844 (N_4844,In_3341,In_1216);
or U4845 (N_4845,In_399,In_2120);
or U4846 (N_4846,In_755,In_4679);
nor U4847 (N_4847,In_1562,In_3354);
and U4848 (N_4848,In_2431,In_3975);
and U4849 (N_4849,In_2846,In_605);
nor U4850 (N_4850,In_1336,In_16);
nand U4851 (N_4851,In_1130,In_2851);
nand U4852 (N_4852,In_4307,In_2834);
nand U4853 (N_4853,In_3322,In_3443);
and U4854 (N_4854,In_4831,In_184);
nand U4855 (N_4855,In_3039,In_1558);
and U4856 (N_4856,In_4506,In_4011);
nor U4857 (N_4857,In_4279,In_4729);
or U4858 (N_4858,In_366,In_546);
nor U4859 (N_4859,In_3718,In_4891);
xnor U4860 (N_4860,In_2154,In_1773);
nand U4861 (N_4861,In_170,In_2104);
and U4862 (N_4862,In_3584,In_4798);
and U4863 (N_4863,In_1950,In_2377);
and U4864 (N_4864,In_84,In_4704);
and U4865 (N_4865,In_1439,In_3317);
and U4866 (N_4866,In_1681,In_4909);
or U4867 (N_4867,In_3847,In_1530);
nor U4868 (N_4868,In_2756,In_669);
nand U4869 (N_4869,In_3920,In_1959);
xor U4870 (N_4870,In_279,In_3810);
or U4871 (N_4871,In_869,In_4972);
or U4872 (N_4872,In_4590,In_3118);
and U4873 (N_4873,In_1406,In_1113);
nor U4874 (N_4874,In_1607,In_732);
or U4875 (N_4875,In_3237,In_174);
or U4876 (N_4876,In_3267,In_4273);
or U4877 (N_4877,In_1842,In_2972);
nor U4878 (N_4878,In_915,In_1395);
nor U4879 (N_4879,In_494,In_611);
and U4880 (N_4880,In_3507,In_2450);
xor U4881 (N_4881,In_4846,In_2837);
and U4882 (N_4882,In_1044,In_2640);
nor U4883 (N_4883,In_1560,In_4615);
nand U4884 (N_4884,In_3695,In_1045);
xor U4885 (N_4885,In_1501,In_4005);
nand U4886 (N_4886,In_895,In_496);
or U4887 (N_4887,In_3974,In_3761);
xor U4888 (N_4888,In_2232,In_750);
nor U4889 (N_4889,In_194,In_1523);
and U4890 (N_4890,In_3265,In_4042);
or U4891 (N_4891,In_2837,In_1961);
xnor U4892 (N_4892,In_4750,In_4457);
nor U4893 (N_4893,In_3329,In_24);
xor U4894 (N_4894,In_93,In_1805);
and U4895 (N_4895,In_3773,In_4622);
or U4896 (N_4896,In_2741,In_973);
nand U4897 (N_4897,In_1767,In_4139);
and U4898 (N_4898,In_4654,In_4445);
xnor U4899 (N_4899,In_2633,In_662);
xor U4900 (N_4900,In_840,In_2272);
and U4901 (N_4901,In_4266,In_1987);
or U4902 (N_4902,In_3244,In_1019);
nor U4903 (N_4903,In_2771,In_1373);
or U4904 (N_4904,In_838,In_3478);
nor U4905 (N_4905,In_4436,In_2374);
nand U4906 (N_4906,In_4615,In_3508);
and U4907 (N_4907,In_4472,In_216);
and U4908 (N_4908,In_3053,In_480);
xor U4909 (N_4909,In_1194,In_2477);
or U4910 (N_4910,In_649,In_4915);
nor U4911 (N_4911,In_4408,In_1662);
xor U4912 (N_4912,In_4941,In_3570);
nor U4913 (N_4913,In_747,In_1908);
or U4914 (N_4914,In_3959,In_3344);
nand U4915 (N_4915,In_1775,In_3783);
and U4916 (N_4916,In_4964,In_3536);
or U4917 (N_4917,In_4418,In_4070);
nor U4918 (N_4918,In_1436,In_950);
or U4919 (N_4919,In_265,In_1652);
or U4920 (N_4920,In_1218,In_1606);
xnor U4921 (N_4921,In_2753,In_4065);
nor U4922 (N_4922,In_1132,In_324);
nor U4923 (N_4923,In_3582,In_4387);
and U4924 (N_4924,In_2704,In_601);
nand U4925 (N_4925,In_4176,In_2482);
nand U4926 (N_4926,In_3497,In_4658);
xor U4927 (N_4927,In_4105,In_3147);
and U4928 (N_4928,In_3756,In_3623);
nand U4929 (N_4929,In_2736,In_3399);
or U4930 (N_4930,In_4009,In_1808);
and U4931 (N_4931,In_2839,In_499);
nor U4932 (N_4932,In_900,In_1467);
nand U4933 (N_4933,In_3932,In_1775);
nand U4934 (N_4934,In_3630,In_3304);
or U4935 (N_4935,In_4262,In_48);
and U4936 (N_4936,In_1293,In_2016);
xor U4937 (N_4937,In_3512,In_4485);
or U4938 (N_4938,In_3503,In_371);
or U4939 (N_4939,In_3697,In_2411);
or U4940 (N_4940,In_3942,In_3068);
nand U4941 (N_4941,In_1498,In_1480);
xnor U4942 (N_4942,In_519,In_1353);
nor U4943 (N_4943,In_3720,In_3568);
xor U4944 (N_4944,In_1974,In_2537);
or U4945 (N_4945,In_2852,In_4413);
or U4946 (N_4946,In_3293,In_527);
xnor U4947 (N_4947,In_3025,In_977);
nand U4948 (N_4948,In_2373,In_2193);
and U4949 (N_4949,In_342,In_1584);
nor U4950 (N_4950,In_3310,In_2231);
nand U4951 (N_4951,In_2759,In_3831);
xnor U4952 (N_4952,In_4047,In_2376);
xor U4953 (N_4953,In_1407,In_4907);
and U4954 (N_4954,In_3849,In_274);
xnor U4955 (N_4955,In_1428,In_4463);
or U4956 (N_4956,In_793,In_3086);
xor U4957 (N_4957,In_688,In_474);
or U4958 (N_4958,In_2342,In_959);
xnor U4959 (N_4959,In_1447,In_291);
and U4960 (N_4960,In_4122,In_1161);
xnor U4961 (N_4961,In_242,In_1751);
or U4962 (N_4962,In_2185,In_1794);
xnor U4963 (N_4963,In_4278,In_3705);
nand U4964 (N_4964,In_4177,In_293);
or U4965 (N_4965,In_4819,In_2389);
nor U4966 (N_4966,In_3805,In_417);
or U4967 (N_4967,In_1523,In_4606);
nand U4968 (N_4968,In_4024,In_1752);
or U4969 (N_4969,In_849,In_4013);
and U4970 (N_4970,In_2557,In_897);
and U4971 (N_4971,In_2480,In_2970);
xor U4972 (N_4972,In_3418,In_1312);
xnor U4973 (N_4973,In_4856,In_2962);
nand U4974 (N_4974,In_807,In_65);
xnor U4975 (N_4975,In_1801,In_540);
or U4976 (N_4976,In_2747,In_3672);
nand U4977 (N_4977,In_4982,In_3747);
nand U4978 (N_4978,In_3223,In_2339);
and U4979 (N_4979,In_364,In_4519);
xor U4980 (N_4980,In_3973,In_1400);
nor U4981 (N_4981,In_1238,In_2850);
or U4982 (N_4982,In_3084,In_1641);
and U4983 (N_4983,In_2890,In_2653);
and U4984 (N_4984,In_1840,In_974);
xnor U4985 (N_4985,In_4526,In_2461);
and U4986 (N_4986,In_2043,In_4680);
nor U4987 (N_4987,In_1901,In_1023);
and U4988 (N_4988,In_4966,In_3007);
nor U4989 (N_4989,In_2009,In_4466);
nor U4990 (N_4990,In_1097,In_3271);
nand U4991 (N_4991,In_2612,In_3234);
nand U4992 (N_4992,In_125,In_1708);
or U4993 (N_4993,In_3586,In_4613);
xor U4994 (N_4994,In_739,In_3438);
nand U4995 (N_4995,In_3134,In_372);
nand U4996 (N_4996,In_1489,In_590);
nor U4997 (N_4997,In_2552,In_51);
nor U4998 (N_4998,In_3100,In_4437);
nand U4999 (N_4999,In_1459,In_1627);
nand U5000 (N_5000,N_3076,N_3250);
nand U5001 (N_5001,N_2063,N_4522);
or U5002 (N_5002,N_1142,N_4838);
nor U5003 (N_5003,N_2448,N_3095);
or U5004 (N_5004,N_3072,N_4451);
nor U5005 (N_5005,N_3451,N_111);
and U5006 (N_5006,N_3321,N_4835);
and U5007 (N_5007,N_1849,N_134);
nor U5008 (N_5008,N_1132,N_1586);
and U5009 (N_5009,N_4825,N_2379);
and U5010 (N_5010,N_1382,N_3780);
and U5011 (N_5011,N_2928,N_759);
or U5012 (N_5012,N_1572,N_1841);
nor U5013 (N_5013,N_1332,N_179);
nand U5014 (N_5014,N_1263,N_3981);
and U5015 (N_5015,N_4015,N_2055);
or U5016 (N_5016,N_927,N_1922);
and U5017 (N_5017,N_3911,N_903);
xor U5018 (N_5018,N_4534,N_1595);
xnor U5019 (N_5019,N_803,N_949);
nand U5020 (N_5020,N_2827,N_4448);
or U5021 (N_5021,N_2706,N_4227);
and U5022 (N_5022,N_517,N_2870);
or U5023 (N_5023,N_4546,N_3417);
nand U5024 (N_5024,N_324,N_4122);
nand U5025 (N_5025,N_4925,N_1186);
or U5026 (N_5026,N_1214,N_1759);
or U5027 (N_5027,N_1268,N_2629);
nand U5028 (N_5028,N_3591,N_1091);
xnor U5029 (N_5029,N_172,N_1642);
and U5030 (N_5030,N_4132,N_2623);
and U5031 (N_5031,N_3037,N_1035);
and U5032 (N_5032,N_608,N_943);
xor U5033 (N_5033,N_3217,N_4208);
xor U5034 (N_5034,N_2573,N_3577);
nor U5035 (N_5035,N_2540,N_381);
nand U5036 (N_5036,N_1191,N_3529);
nor U5037 (N_5037,N_984,N_2054);
nor U5038 (N_5038,N_3562,N_1236);
or U5039 (N_5039,N_1245,N_4332);
and U5040 (N_5040,N_2316,N_1411);
nor U5041 (N_5041,N_2489,N_2222);
nand U5042 (N_5042,N_643,N_1379);
and U5043 (N_5043,N_3506,N_557);
nor U5044 (N_5044,N_1936,N_1068);
nor U5045 (N_5045,N_359,N_726);
or U5046 (N_5046,N_3766,N_4251);
and U5047 (N_5047,N_1896,N_2499);
nand U5048 (N_5048,N_3488,N_4259);
and U5049 (N_5049,N_2701,N_2925);
or U5050 (N_5050,N_4974,N_3950);
and U5051 (N_5051,N_1394,N_3336);
nor U5052 (N_5052,N_1745,N_4301);
xor U5053 (N_5053,N_2861,N_495);
or U5054 (N_5054,N_1094,N_2694);
nor U5055 (N_5055,N_4314,N_1565);
xnor U5056 (N_5056,N_245,N_142);
nor U5057 (N_5057,N_455,N_1979);
nor U5058 (N_5058,N_1467,N_3782);
xnor U5059 (N_5059,N_336,N_454);
xor U5060 (N_5060,N_2172,N_1291);
and U5061 (N_5061,N_3604,N_3288);
nor U5062 (N_5062,N_4071,N_4004);
nand U5063 (N_5063,N_1518,N_100);
and U5064 (N_5064,N_1788,N_4640);
nand U5065 (N_5065,N_4253,N_2116);
xor U5066 (N_5066,N_1978,N_57);
and U5067 (N_5067,N_3497,N_1898);
nor U5068 (N_5068,N_3500,N_4036);
nand U5069 (N_5069,N_1993,N_699);
and U5070 (N_5070,N_4630,N_267);
xnor U5071 (N_5071,N_3333,N_2248);
and U5072 (N_5072,N_3007,N_3086);
nand U5073 (N_5073,N_2099,N_4211);
or U5074 (N_5074,N_4169,N_4257);
and U5075 (N_5075,N_897,N_1597);
nor U5076 (N_5076,N_4535,N_4544);
and U5077 (N_5077,N_2105,N_2654);
or U5078 (N_5078,N_528,N_3262);
nor U5079 (N_5079,N_1298,N_4912);
nand U5080 (N_5080,N_964,N_2256);
and U5081 (N_5081,N_560,N_820);
nor U5082 (N_5082,N_4929,N_1342);
nor U5083 (N_5083,N_3310,N_4757);
or U5084 (N_5084,N_1280,N_4217);
nor U5085 (N_5085,N_3832,N_1847);
and U5086 (N_5086,N_911,N_2850);
or U5087 (N_5087,N_2298,N_4698);
nor U5088 (N_5088,N_3842,N_4962);
nand U5089 (N_5089,N_3283,N_593);
nand U5090 (N_5090,N_471,N_2755);
nand U5091 (N_5091,N_4039,N_3306);
nand U5092 (N_5092,N_854,N_1466);
nor U5093 (N_5093,N_635,N_259);
nor U5094 (N_5094,N_4858,N_1431);
xnor U5095 (N_5095,N_4876,N_2401);
xnor U5096 (N_5096,N_3660,N_4877);
and U5097 (N_5097,N_914,N_2957);
nor U5098 (N_5098,N_1010,N_816);
or U5099 (N_5099,N_4862,N_1807);
xor U5100 (N_5100,N_4268,N_3944);
xnor U5101 (N_5101,N_3522,N_1450);
xnor U5102 (N_5102,N_3483,N_4599);
xnor U5103 (N_5103,N_2249,N_915);
or U5104 (N_5104,N_286,N_2264);
and U5105 (N_5105,N_4981,N_1677);
xnor U5106 (N_5106,N_4933,N_4135);
nand U5107 (N_5107,N_2851,N_4394);
or U5108 (N_5108,N_930,N_2735);
and U5109 (N_5109,N_1724,N_1520);
nor U5110 (N_5110,N_4754,N_1140);
and U5111 (N_5111,N_4337,N_2787);
nor U5112 (N_5112,N_158,N_1353);
nor U5113 (N_5113,N_656,N_487);
nor U5114 (N_5114,N_3729,N_1076);
nor U5115 (N_5115,N_1503,N_2125);
xor U5116 (N_5116,N_1130,N_3212);
xnor U5117 (N_5117,N_1653,N_4238);
or U5118 (N_5118,N_2718,N_2660);
or U5119 (N_5119,N_379,N_107);
and U5120 (N_5120,N_4644,N_3247);
nand U5121 (N_5121,N_2395,N_3495);
xor U5122 (N_5122,N_2671,N_503);
xnor U5123 (N_5123,N_1723,N_2916);
or U5124 (N_5124,N_249,N_1716);
or U5125 (N_5125,N_1324,N_2644);
nand U5126 (N_5126,N_880,N_861);
and U5127 (N_5127,N_3746,N_2219);
xnor U5128 (N_5128,N_806,N_3230);
and U5129 (N_5129,N_1425,N_3942);
and U5130 (N_5130,N_2896,N_676);
nor U5131 (N_5131,N_3162,N_4673);
and U5132 (N_5132,N_909,N_60);
nor U5133 (N_5133,N_10,N_4119);
and U5134 (N_5134,N_266,N_2602);
or U5135 (N_5135,N_2495,N_1780);
nor U5136 (N_5136,N_867,N_4);
and U5137 (N_5137,N_3605,N_2323);
xnor U5138 (N_5138,N_2142,N_3665);
xor U5139 (N_5139,N_1292,N_646);
or U5140 (N_5140,N_3024,N_3438);
nor U5141 (N_5141,N_410,N_2403);
nor U5142 (N_5142,N_4773,N_3082);
nand U5143 (N_5143,N_4676,N_2051);
nand U5144 (N_5144,N_4367,N_4847);
or U5145 (N_5145,N_1444,N_125);
and U5146 (N_5146,N_1546,N_4559);
xor U5147 (N_5147,N_341,N_801);
xnor U5148 (N_5148,N_4371,N_1135);
and U5149 (N_5149,N_4146,N_2983);
and U5150 (N_5150,N_3485,N_2299);
nor U5151 (N_5151,N_4218,N_4973);
or U5152 (N_5152,N_2552,N_1602);
or U5153 (N_5153,N_3365,N_735);
xor U5154 (N_5154,N_4324,N_182);
xnor U5155 (N_5155,N_3923,N_1080);
nand U5156 (N_5156,N_4882,N_4789);
nand U5157 (N_5157,N_1088,N_288);
nor U5158 (N_5158,N_2458,N_4734);
or U5159 (N_5159,N_4903,N_1933);
or U5160 (N_5160,N_3499,N_4396);
nand U5161 (N_5161,N_1590,N_1935);
or U5162 (N_5162,N_3091,N_2663);
nand U5163 (N_5163,N_9,N_4984);
nand U5164 (N_5164,N_3254,N_3195);
nand U5165 (N_5165,N_4033,N_4315);
xor U5166 (N_5166,N_814,N_3236);
and U5167 (N_5167,N_4832,N_2149);
nand U5168 (N_5168,N_2881,N_2025);
xnor U5169 (N_5169,N_2453,N_4172);
nor U5170 (N_5170,N_4302,N_1853);
nor U5171 (N_5171,N_946,N_1383);
nand U5172 (N_5172,N_1900,N_4439);
xor U5173 (N_5173,N_1260,N_87);
xor U5174 (N_5174,N_2723,N_1034);
xnor U5175 (N_5175,N_4181,N_4814);
nand U5176 (N_5176,N_4088,N_3853);
or U5177 (N_5177,N_3512,N_1108);
nand U5178 (N_5178,N_4417,N_4867);
xor U5179 (N_5179,N_374,N_4567);
or U5180 (N_5180,N_2441,N_3213);
or U5181 (N_5181,N_4810,N_4025);
nor U5182 (N_5182,N_3996,N_4745);
xnor U5183 (N_5183,N_4796,N_2724);
and U5184 (N_5184,N_3580,N_745);
nand U5185 (N_5185,N_4688,N_2865);
and U5186 (N_5186,N_3801,N_3927);
or U5187 (N_5187,N_1127,N_2271);
and U5188 (N_5188,N_108,N_3104);
or U5189 (N_5189,N_2824,N_3433);
xnor U5190 (N_5190,N_68,N_1947);
or U5191 (N_5191,N_4478,N_678);
and U5192 (N_5192,N_4602,N_4591);
nor U5193 (N_5193,N_979,N_361);
and U5194 (N_5194,N_1064,N_3208);
nor U5195 (N_5195,N_4896,N_4628);
and U5196 (N_5196,N_4017,N_500);
or U5197 (N_5197,N_1888,N_1030);
and U5198 (N_5198,N_494,N_1687);
and U5199 (N_5199,N_2003,N_1011);
or U5200 (N_5200,N_3307,N_522);
nand U5201 (N_5201,N_2768,N_3342);
nor U5202 (N_5202,N_2417,N_21);
nor U5203 (N_5203,N_2531,N_3294);
or U5204 (N_5204,N_3285,N_1928);
xor U5205 (N_5205,N_1481,N_1469);
and U5206 (N_5206,N_3172,N_2998);
xnor U5207 (N_5207,N_3077,N_1519);
nor U5208 (N_5208,N_681,N_2347);
or U5209 (N_5209,N_3825,N_2225);
or U5210 (N_5210,N_4442,N_4714);
nand U5211 (N_5211,N_2900,N_169);
nand U5212 (N_5212,N_4505,N_2362);
xnor U5213 (N_5213,N_2775,N_2825);
nand U5214 (N_5214,N_3754,N_3376);
xor U5215 (N_5215,N_4086,N_2094);
or U5216 (N_5216,N_20,N_1406);
nand U5217 (N_5217,N_1567,N_3144);
xor U5218 (N_5218,N_3219,N_3034);
or U5219 (N_5219,N_3795,N_2652);
nor U5220 (N_5220,N_1905,N_1373);
nor U5221 (N_5221,N_3673,N_83);
nand U5222 (N_5222,N_393,N_2399);
nand U5223 (N_5223,N_1463,N_1131);
and U5224 (N_5224,N_67,N_862);
nand U5225 (N_5225,N_4307,N_4826);
and U5226 (N_5226,N_1402,N_287);
or U5227 (N_5227,N_874,N_2632);
and U5228 (N_5228,N_2292,N_4897);
xnor U5229 (N_5229,N_3183,N_250);
xnor U5230 (N_5230,N_4645,N_1533);
xor U5231 (N_5231,N_236,N_2965);
nand U5232 (N_5232,N_2402,N_542);
and U5233 (N_5233,N_4166,N_674);
nor U5234 (N_5234,N_123,N_2221);
nand U5235 (N_5235,N_2188,N_912);
and U5236 (N_5236,N_2015,N_918);
nand U5237 (N_5237,N_3636,N_4972);
nand U5238 (N_5238,N_1734,N_3722);
nor U5239 (N_5239,N_4006,N_1190);
or U5240 (N_5240,N_423,N_4229);
xor U5241 (N_5241,N_3860,N_4099);
and U5242 (N_5242,N_2022,N_4162);
and U5243 (N_5243,N_1470,N_1040);
or U5244 (N_5244,N_1483,N_4596);
or U5245 (N_5245,N_2630,N_1018);
nor U5246 (N_5246,N_1987,N_2875);
nor U5247 (N_5247,N_838,N_4340);
nand U5248 (N_5248,N_2554,N_1109);
and U5249 (N_5249,N_4914,N_3056);
xnor U5250 (N_5250,N_407,N_2367);
and U5251 (N_5251,N_599,N_3229);
or U5252 (N_5252,N_1920,N_1418);
nand U5253 (N_5253,N_3627,N_3468);
and U5254 (N_5254,N_4403,N_2129);
nor U5255 (N_5255,N_1377,N_4993);
or U5256 (N_5256,N_439,N_2559);
or U5257 (N_5257,N_2866,N_1715);
nor U5258 (N_5258,N_1072,N_3057);
nand U5259 (N_5259,N_334,N_181);
or U5260 (N_5260,N_665,N_3013);
xor U5261 (N_5261,N_2252,N_690);
nand U5262 (N_5262,N_2037,N_61);
xnor U5263 (N_5263,N_162,N_1721);
nor U5264 (N_5264,N_4863,N_1981);
and U5265 (N_5265,N_1711,N_269);
nand U5266 (N_5266,N_4750,N_680);
or U5267 (N_5267,N_103,N_2297);
or U5268 (N_5268,N_4120,N_8);
nor U5269 (N_5269,N_4298,N_1618);
and U5270 (N_5270,N_2538,N_1569);
and U5271 (N_5271,N_3119,N_2296);
and U5272 (N_5272,N_4947,N_4737);
nor U5273 (N_5273,N_2542,N_3012);
or U5274 (N_5274,N_1443,N_3735);
or U5275 (N_5275,N_4326,N_3620);
and U5276 (N_5276,N_4457,N_2800);
xor U5277 (N_5277,N_1587,N_2942);
nor U5278 (N_5278,N_1525,N_4999);
or U5279 (N_5279,N_1316,N_4627);
and U5280 (N_5280,N_62,N_1848);
xor U5281 (N_5281,N_2502,N_424);
nand U5282 (N_5282,N_1852,N_4704);
and U5283 (N_5283,N_1166,N_2912);
or U5284 (N_5284,N_3480,N_1966);
or U5285 (N_5285,N_2715,N_1516);
nor U5286 (N_5286,N_961,N_175);
nor U5287 (N_5287,N_1070,N_632);
and U5288 (N_5288,N_1434,N_3520);
and U5289 (N_5289,N_371,N_2636);
nand U5290 (N_5290,N_4322,N_2622);
and U5291 (N_5291,N_3980,N_2203);
or U5292 (N_5292,N_4222,N_4389);
and U5293 (N_5293,N_1955,N_318);
nand U5294 (N_5294,N_1649,N_161);
nand U5295 (N_5295,N_3978,N_3032);
and U5296 (N_5296,N_3784,N_2053);
and U5297 (N_5297,N_784,N_116);
xnor U5298 (N_5298,N_1453,N_4680);
or U5299 (N_5299,N_1976,N_2887);
or U5300 (N_5300,N_877,N_793);
xor U5301 (N_5301,N_4793,N_2781);
nor U5302 (N_5302,N_4202,N_4007);
or U5303 (N_5303,N_2158,N_2670);
and U5304 (N_5304,N_2693,N_3234);
nor U5305 (N_5305,N_4992,N_2014);
nand U5306 (N_5306,N_3994,N_1170);
xnor U5307 (N_5307,N_2430,N_240);
xor U5308 (N_5308,N_3816,N_4874);
nor U5309 (N_5309,N_569,N_4785);
or U5310 (N_5310,N_2832,N_4117);
and U5311 (N_5311,N_4312,N_1855);
and U5312 (N_5312,N_292,N_4192);
and U5313 (N_5313,N_2805,N_136);
nand U5314 (N_5314,N_3101,N_3679);
or U5315 (N_5315,N_4769,N_1247);
nor U5316 (N_5316,N_4583,N_4020);
xnor U5317 (N_5317,N_2212,N_3109);
or U5318 (N_5318,N_4566,N_247);
or U5319 (N_5319,N_2049,N_2553);
and U5320 (N_5320,N_1584,N_3384);
or U5321 (N_5321,N_37,N_316);
nand U5322 (N_5322,N_4724,N_3293);
xor U5323 (N_5323,N_4995,N_1760);
or U5324 (N_5324,N_4074,N_4141);
or U5325 (N_5325,N_3658,N_3667);
xor U5326 (N_5326,N_4030,N_514);
nor U5327 (N_5327,N_1158,N_2304);
and U5328 (N_5328,N_4647,N_2950);
nor U5329 (N_5329,N_1305,N_4184);
nor U5330 (N_5330,N_2589,N_4240);
and U5331 (N_5331,N_1959,N_2784);
and U5332 (N_5332,N_4341,N_4779);
nand U5333 (N_5333,N_3719,N_2618);
nor U5334 (N_5334,N_3,N_1908);
xor U5335 (N_5335,N_4935,N_2208);
nand U5336 (N_5336,N_3493,N_2904);
nor U5337 (N_5337,N_4594,N_2944);
nor U5338 (N_5338,N_2712,N_3023);
or U5339 (N_5339,N_3837,N_3706);
nand U5340 (N_5340,N_3134,N_293);
nand U5341 (N_5341,N_1143,N_2451);
nor U5342 (N_5342,N_3955,N_3595);
and U5343 (N_5343,N_3596,N_1562);
or U5344 (N_5344,N_660,N_769);
or U5345 (N_5345,N_426,N_1722);
xor U5346 (N_5346,N_3439,N_99);
nor U5347 (N_5347,N_1173,N_1782);
and U5348 (N_5348,N_2523,N_2348);
nor U5349 (N_5349,N_2518,N_2862);
nand U5350 (N_5350,N_1179,N_3871);
or U5351 (N_5351,N_4436,N_1641);
nand U5352 (N_5352,N_2019,N_513);
nor U5353 (N_5353,N_4890,N_4082);
xor U5354 (N_5354,N_4456,N_3872);
and U5355 (N_5355,N_4717,N_3074);
xnor U5356 (N_5356,N_4455,N_1574);
or U5357 (N_5357,N_3118,N_4305);
xnor U5358 (N_5358,N_2678,N_4803);
and U5359 (N_5359,N_4529,N_3299);
or U5360 (N_5360,N_412,N_3295);
and U5361 (N_5361,N_1363,N_3351);
or U5362 (N_5362,N_378,N_2634);
nand U5363 (N_5363,N_3277,N_2217);
and U5364 (N_5364,N_795,N_4770);
xor U5365 (N_5365,N_863,N_649);
xor U5366 (N_5366,N_2325,N_4986);
and U5367 (N_5367,N_1155,N_4143);
and U5368 (N_5368,N_3202,N_89);
nand U5369 (N_5369,N_655,N_997);
nand U5370 (N_5370,N_3715,N_1599);
or U5371 (N_5371,N_1776,N_1257);
nand U5372 (N_5372,N_4956,N_2387);
nand U5373 (N_5373,N_2835,N_2171);
xor U5374 (N_5374,N_804,N_1028);
xor U5375 (N_5375,N_1666,N_845);
nor U5376 (N_5376,N_1084,N_3607);
xor U5377 (N_5377,N_2426,N_2570);
xor U5378 (N_5378,N_1521,N_4351);
nand U5379 (N_5379,N_2389,N_3160);
xor U5380 (N_5380,N_591,N_567);
or U5381 (N_5381,N_1779,N_155);
xor U5382 (N_5382,N_4741,N_2072);
xnor U5383 (N_5383,N_2609,N_192);
nor U5384 (N_5384,N_3946,N_2673);
nor U5385 (N_5385,N_2988,N_3028);
nand U5386 (N_5386,N_2742,N_2612);
xnor U5387 (N_5387,N_2102,N_3696);
nor U5388 (N_5388,N_1426,N_3915);
or U5389 (N_5389,N_506,N_1032);
nand U5390 (N_5390,N_3089,N_2119);
and U5391 (N_5391,N_2516,N_4279);
or U5392 (N_5392,N_2211,N_4512);
nor U5393 (N_5393,N_3400,N_2720);
or U5394 (N_5394,N_3820,N_1523);
or U5395 (N_5395,N_3427,N_3773);
nor U5396 (N_5396,N_4648,N_581);
or U5397 (N_5397,N_4157,N_3800);
nand U5398 (N_5398,N_1542,N_2356);
nand U5399 (N_5399,N_1067,N_347);
xor U5400 (N_5400,N_1720,N_1694);
or U5401 (N_5401,N_3537,N_109);
nor U5402 (N_5402,N_686,N_2743);
or U5403 (N_5403,N_4092,N_3455);
or U5404 (N_5404,N_4811,N_3831);
nand U5405 (N_5405,N_2408,N_2065);
and U5406 (N_5406,N_4809,N_59);
nand U5407 (N_5407,N_3041,N_211);
or U5408 (N_5408,N_4880,N_572);
xnor U5409 (N_5409,N_2621,N_2600);
nor U5410 (N_5410,N_480,N_3066);
or U5411 (N_5411,N_2750,N_2093);
nand U5412 (N_5412,N_2889,N_4400);
nand U5413 (N_5413,N_2452,N_71);
nor U5414 (N_5414,N_1014,N_3446);
nand U5415 (N_5415,N_2884,N_4922);
nor U5416 (N_5416,N_3105,N_114);
and U5417 (N_5417,N_4023,N_32);
nand U5418 (N_5418,N_4467,N_3033);
nand U5419 (N_5419,N_4133,N_1029);
nand U5420 (N_5420,N_4778,N_3245);
and U5421 (N_5421,N_2682,N_3344);
and U5422 (N_5422,N_1526,N_2420);
and U5423 (N_5423,N_4420,N_153);
or U5424 (N_5424,N_2771,N_1207);
and U5425 (N_5425,N_1793,N_2593);
nor U5426 (N_5426,N_3249,N_648);
nor U5427 (N_5427,N_2463,N_4245);
xor U5428 (N_5428,N_2153,N_417);
xor U5429 (N_5429,N_3813,N_3507);
and U5430 (N_5430,N_3354,N_2938);
nand U5431 (N_5431,N_3828,N_2932);
and U5432 (N_5432,N_4252,N_2326);
xnor U5433 (N_5433,N_4387,N_3976);
nand U5434 (N_5434,N_3760,N_546);
xnor U5435 (N_5435,N_2337,N_3140);
xnor U5436 (N_5436,N_1013,N_4495);
nand U5437 (N_5437,N_1341,N_3919);
xnor U5438 (N_5438,N_762,N_4272);
or U5439 (N_5439,N_3243,N_4009);
xor U5440 (N_5440,N_1006,N_712);
nor U5441 (N_5441,N_3067,N_1834);
nor U5442 (N_5442,N_2295,N_609);
nand U5443 (N_5443,N_340,N_152);
and U5444 (N_5444,N_3962,N_3752);
or U5445 (N_5445,N_121,N_4357);
and U5446 (N_5446,N_976,N_2982);
or U5447 (N_5447,N_2036,N_4424);
nor U5448 (N_5448,N_3450,N_1772);
xnor U5449 (N_5449,N_3961,N_4255);
xor U5450 (N_5450,N_3684,N_3622);
nor U5451 (N_5451,N_958,N_4083);
and U5452 (N_5452,N_682,N_4979);
and U5453 (N_5453,N_4294,N_4637);
and U5454 (N_5454,N_3611,N_96);
or U5455 (N_5455,N_129,N_2493);
nand U5456 (N_5456,N_1369,N_4308);
nand U5457 (N_5457,N_688,N_3014);
nor U5458 (N_5458,N_1505,N_780);
nor U5459 (N_5459,N_75,N_117);
or U5460 (N_5460,N_3639,N_4376);
or U5461 (N_5461,N_945,N_4547);
and U5462 (N_5462,N_2159,N_4435);
or U5463 (N_5463,N_3064,N_538);
nand U5464 (N_5464,N_4418,N_1970);
or U5465 (N_5465,N_1536,N_4998);
and U5466 (N_5466,N_1648,N_3350);
or U5467 (N_5467,N_3535,N_388);
xor U5468 (N_5468,N_2937,N_4468);
and U5469 (N_5469,N_4213,N_437);
or U5470 (N_5470,N_4354,N_4244);
and U5471 (N_5471,N_550,N_4067);
or U5472 (N_5472,N_1455,N_1460);
and U5473 (N_5473,N_4289,N_3052);
or U5474 (N_5474,N_4454,N_855);
and U5475 (N_5475,N_3395,N_3316);
and U5476 (N_5476,N_3670,N_4554);
nand U5477 (N_5477,N_1038,N_1294);
or U5478 (N_5478,N_1507,N_1082);
or U5479 (N_5479,N_703,N_4084);
or U5480 (N_5480,N_1036,N_433);
xnor U5481 (N_5481,N_4089,N_4997);
nor U5482 (N_5482,N_4399,N_493);
xor U5483 (N_5483,N_3573,N_2915);
or U5484 (N_5484,N_2274,N_702);
and U5485 (N_5485,N_2869,N_3418);
nand U5486 (N_5486,N_625,N_3778);
nor U5487 (N_5487,N_3610,N_3758);
and U5488 (N_5488,N_4195,N_1833);
nor U5489 (N_5489,N_4790,N_3073);
nand U5490 (N_5490,N_2539,N_2422);
and U5491 (N_5491,N_305,N_1478);
or U5492 (N_5492,N_399,N_2338);
xnor U5493 (N_5493,N_4759,N_1001);
or U5494 (N_5494,N_2327,N_1891);
nor U5495 (N_5495,N_4118,N_4003);
and U5496 (N_5496,N_3601,N_3868);
and U5497 (N_5497,N_2684,N_131);
nand U5498 (N_5498,N_127,N_1151);
nor U5499 (N_5499,N_1835,N_2058);
xnor U5500 (N_5500,N_4585,N_427);
or U5501 (N_5501,N_2253,N_4582);
xnor U5502 (N_5502,N_3690,N_3796);
nand U5503 (N_5503,N_2744,N_3811);
xor U5504 (N_5504,N_4419,N_2178);
and U5505 (N_5505,N_418,N_4710);
and U5506 (N_5506,N_3000,N_3367);
xor U5507 (N_5507,N_1864,N_832);
nor U5508 (N_5508,N_1317,N_4210);
or U5509 (N_5509,N_2088,N_28);
nor U5510 (N_5510,N_4685,N_2586);
nand U5511 (N_5511,N_829,N_1413);
xnor U5512 (N_5512,N_3656,N_2601);
nor U5513 (N_5513,N_3258,N_3298);
nand U5514 (N_5514,N_113,N_3286);
nor U5515 (N_5515,N_3779,N_4675);
and U5516 (N_5516,N_2459,N_1424);
or U5517 (N_5517,N_2814,N_2527);
nor U5518 (N_5518,N_3492,N_2650);
xor U5519 (N_5519,N_952,N_4319);
xnor U5520 (N_5520,N_4760,N_3792);
nand U5521 (N_5521,N_3844,N_4488);
nor U5522 (N_5522,N_2890,N_2007);
xor U5523 (N_5523,N_2580,N_4140);
xnor U5524 (N_5524,N_4219,N_2310);
and U5525 (N_5525,N_1510,N_3867);
xor U5526 (N_5526,N_3705,N_4952);
nand U5527 (N_5527,N_636,N_26);
or U5528 (N_5528,N_1200,N_4413);
and U5529 (N_5529,N_4114,N_196);
and U5530 (N_5530,N_2797,N_2255);
nand U5531 (N_5531,N_130,N_3322);
nand U5532 (N_5532,N_1804,N_4855);
xnor U5533 (N_5533,N_3847,N_2853);
xor U5534 (N_5534,N_1764,N_2613);
xnor U5535 (N_5535,N_4048,N_856);
or U5536 (N_5536,N_1231,N_3121);
and U5537 (N_5537,N_326,N_3353);
or U5538 (N_5538,N_2440,N_2547);
and U5539 (N_5539,N_4701,N_3998);
or U5540 (N_5540,N_3478,N_405);
and U5541 (N_5541,N_344,N_4104);
nor U5542 (N_5542,N_4481,N_386);
nand U5543 (N_5543,N_449,N_694);
or U5544 (N_5544,N_978,N_1386);
nor U5545 (N_5545,N_3192,N_333);
xnor U5546 (N_5546,N_4946,N_1787);
or U5547 (N_5547,N_2237,N_1251);
xor U5548 (N_5548,N_2599,N_4438);
nand U5549 (N_5549,N_4500,N_3724);
and U5550 (N_5550,N_3125,N_4277);
or U5551 (N_5551,N_4957,N_264);
and U5552 (N_5552,N_3175,N_1675);
and U5553 (N_5553,N_2439,N_2154);
nand U5554 (N_5554,N_2184,N_791);
or U5555 (N_5555,N_4306,N_3514);
nor U5556 (N_5556,N_4005,N_1457);
or U5557 (N_5557,N_992,N_2511);
xnor U5558 (N_5558,N_1205,N_3669);
nand U5559 (N_5559,N_753,N_4123);
nor U5560 (N_5560,N_3435,N_3338);
nand U5561 (N_5561,N_2813,N_837);
xor U5562 (N_5562,N_3198,N_1558);
and U5563 (N_5563,N_508,N_637);
and U5564 (N_5564,N_4476,N_382);
nand U5565 (N_5565,N_3516,N_1707);
xnor U5566 (N_5566,N_3574,N_2729);
and U5567 (N_5567,N_2557,N_778);
nand U5568 (N_5568,N_4802,N_2012);
and U5569 (N_5569,N_4728,N_4942);
and U5570 (N_5570,N_422,N_2366);
xnor U5571 (N_5571,N_2114,N_2638);
xnor U5572 (N_5572,N_206,N_170);
and U5573 (N_5573,N_277,N_4856);
xor U5574 (N_5574,N_2226,N_2848);
xor U5575 (N_5575,N_4292,N_1632);
nor U5576 (N_5576,N_2961,N_1056);
and U5577 (N_5577,N_3572,N_1148);
xor U5578 (N_5578,N_2429,N_383);
nand U5579 (N_5579,N_4385,N_3829);
xnor U5580 (N_5580,N_605,N_545);
or U5581 (N_5581,N_1230,N_499);
and U5582 (N_5582,N_4483,N_3017);
xor U5583 (N_5583,N_4806,N_2675);
and U5584 (N_5584,N_835,N_434);
or U5585 (N_5585,N_3889,N_908);
nor U5586 (N_5586,N_3846,N_2123);
or U5587 (N_5587,N_2639,N_456);
nand U5588 (N_5588,N_3408,N_1459);
nor U5589 (N_5589,N_3268,N_432);
or U5590 (N_5590,N_1880,N_2436);
or U5591 (N_5591,N_4256,N_4393);
nor U5592 (N_5592,N_1279,N_731);
or U5593 (N_5593,N_4098,N_4702);
xor U5594 (N_5594,N_4026,N_607);
nor U5595 (N_5595,N_4697,N_2550);
nand U5596 (N_5596,N_3649,N_201);
and U5597 (N_5597,N_4684,N_327);
nand U5598 (N_5598,N_4926,N_2407);
xnor U5599 (N_5599,N_2576,N_1479);
xnor U5600 (N_5600,N_3775,N_2301);
xnor U5601 (N_5601,N_2287,N_2156);
nand U5602 (N_5602,N_3710,N_3371);
or U5603 (N_5603,N_1061,N_1354);
xor U5604 (N_5604,N_2239,N_1821);
or U5605 (N_5605,N_3939,N_2400);
xnor U5606 (N_5606,N_2421,N_4328);
nor U5607 (N_5607,N_623,N_1913);
or U5608 (N_5608,N_4771,N_3672);
or U5609 (N_5609,N_4248,N_1344);
nand U5610 (N_5610,N_2293,N_2761);
xor U5611 (N_5611,N_1529,N_1216);
xnor U5612 (N_5612,N_2331,N_3035);
nand U5613 (N_5613,N_317,N_1071);
xor U5614 (N_5614,N_1730,N_4706);
or U5615 (N_5615,N_4053,N_4853);
and U5616 (N_5616,N_4032,N_2628);
and U5617 (N_5617,N_4868,N_3080);
or U5618 (N_5618,N_4047,N_4681);
nor U5619 (N_5619,N_2981,N_4449);
or U5620 (N_5620,N_4885,N_4930);
nor U5621 (N_5621,N_813,N_1563);
nand U5622 (N_5622,N_3477,N_3732);
xnor U5623 (N_5623,N_2190,N_4078);
and U5624 (N_5624,N_2275,N_3539);
nor U5625 (N_5625,N_4907,N_4845);
nand U5626 (N_5626,N_3324,N_933);
and U5627 (N_5627,N_3659,N_1678);
nor U5628 (N_5628,N_3726,N_3986);
and U5629 (N_5629,N_1240,N_4545);
nor U5630 (N_5630,N_1327,N_4515);
and U5631 (N_5631,N_296,N_1199);
xnor U5632 (N_5632,N_617,N_3548);
nand U5633 (N_5633,N_1408,N_751);
nor U5634 (N_5634,N_1695,N_1578);
and U5635 (N_5635,N_925,N_3635);
and U5636 (N_5636,N_973,N_3644);
nor U5637 (N_5637,N_180,N_4911);
nand U5638 (N_5638,N_1926,N_3525);
and U5639 (N_5639,N_4107,N_2692);
and U5640 (N_5640,N_442,N_1492);
xnor U5641 (N_5641,N_3533,N_4953);
nor U5642 (N_5642,N_3135,N_2468);
or U5643 (N_5643,N_1708,N_4940);
nor U5644 (N_5644,N_670,N_3764);
nand U5645 (N_5645,N_3005,N_3972);
nor U5646 (N_5646,N_4295,N_1404);
or U5647 (N_5647,N_1893,N_2717);
or U5648 (N_5648,N_474,N_1322);
and U5649 (N_5649,N_4924,N_708);
or U5650 (N_5650,N_1917,N_3275);
and U5651 (N_5651,N_2060,N_802);
nor U5652 (N_5652,N_1557,N_3751);
and U5653 (N_5653,N_1881,N_88);
nor U5654 (N_5654,N_1644,N_586);
nand U5655 (N_5655,N_3407,N_337);
or U5656 (N_5656,N_4891,N_2457);
or U5657 (N_5657,N_4234,N_4423);
nand U5658 (N_5658,N_732,N_967);
nor U5659 (N_5659,N_4652,N_698);
and U5660 (N_5660,N_1664,N_2946);
nand U5661 (N_5661,N_705,N_2508);
nor U5662 (N_5662,N_2996,N_4461);
nor U5663 (N_5663,N_2033,N_2194);
nand U5664 (N_5664,N_1903,N_4689);
and U5665 (N_5665,N_1836,N_3030);
nand U5666 (N_5666,N_3975,N_3930);
nor U5667 (N_5667,N_2596,N_4008);
nand U5668 (N_5668,N_166,N_3389);
nand U5669 (N_5669,N_4818,N_2454);
and U5670 (N_5670,N_3940,N_3692);
or U5671 (N_5671,N_202,N_3788);
nand U5672 (N_5672,N_4293,N_3233);
or U5673 (N_5673,N_1911,N_1973);
xor U5674 (N_5674,N_1725,N_273);
nand U5675 (N_5675,N_507,N_783);
and U5676 (N_5676,N_1306,N_4404);
nand U5677 (N_5677,N_2042,N_4638);
nor U5678 (N_5678,N_4441,N_2767);
nand U5679 (N_5679,N_2524,N_4738);
xor U5680 (N_5680,N_302,N_53);
nand U5681 (N_5681,N_3585,N_425);
nand U5682 (N_5682,N_3209,N_3893);
nor U5683 (N_5683,N_2286,N_516);
or U5684 (N_5684,N_164,N_4193);
or U5685 (N_5685,N_3456,N_1269);
nor U5686 (N_5686,N_2284,N_2394);
and U5687 (N_5687,N_3097,N_1271);
and U5688 (N_5688,N_132,N_4991);
or U5689 (N_5689,N_631,N_4579);
nor U5690 (N_5690,N_1113,N_821);
nand U5691 (N_5691,N_2038,N_4543);
or U5692 (N_5692,N_2135,N_673);
or U5693 (N_5693,N_1549,N_3805);
nand U5694 (N_5694,N_2397,N_3567);
nor U5695 (N_5695,N_934,N_35);
nand U5696 (N_5696,N_4105,N_2278);
xor U5697 (N_5697,N_2734,N_1600);
nand U5698 (N_5698,N_176,N_2574);
nor U5699 (N_5699,N_1159,N_4669);
or U5700 (N_5700,N_1929,N_2103);
nor U5701 (N_5701,N_2005,N_3127);
xnor U5702 (N_5702,N_2235,N_342);
and U5703 (N_5703,N_1866,N_452);
nand U5704 (N_5704,N_1116,N_1514);
xnor U5705 (N_5705,N_895,N_4465);
or U5706 (N_5706,N_1609,N_3416);
and U5707 (N_5707,N_1568,N_2918);
xor U5708 (N_5708,N_4887,N_2204);
and U5709 (N_5709,N_1957,N_4270);
xor U5710 (N_5710,N_2335,N_4384);
nor U5711 (N_5711,N_3334,N_4024);
xnor U5712 (N_5712,N_2704,N_3689);
xnor U5713 (N_5713,N_482,N_2886);
xor U5714 (N_5714,N_4031,N_2611);
and U5715 (N_5715,N_810,N_4881);
or U5716 (N_5716,N_1551,N_1615);
nand U5717 (N_5717,N_3252,N_465);
nor U5718 (N_5718,N_1669,N_3568);
nor U5719 (N_5719,N_1177,N_3606);
xor U5720 (N_5720,N_840,N_3569);
xor U5721 (N_5721,N_1690,N_1005);
or U5722 (N_5722,N_2736,N_4733);
xor U5723 (N_5723,N_207,N_4052);
xnor U5724 (N_5724,N_2450,N_3861);
nand U5725 (N_5725,N_4223,N_736);
or U5726 (N_5726,N_2091,N_3903);
and U5727 (N_5727,N_4538,N_2345);
nor U5728 (N_5728,N_208,N_1497);
nand U5729 (N_5729,N_2776,N_4615);
or U5730 (N_5730,N_3267,N_1771);
and U5731 (N_5731,N_679,N_4447);
and U5732 (N_5732,N_4578,N_1472);
nand U5733 (N_5733,N_3637,N_1761);
nand U5734 (N_5734,N_1663,N_1717);
or U5735 (N_5735,N_2043,N_2066);
or U5736 (N_5736,N_4060,N_4236);
nand U5737 (N_5737,N_3841,N_3083);
nand U5738 (N_5738,N_2386,N_3008);
nand U5739 (N_5739,N_2838,N_4695);
and U5740 (N_5740,N_721,N_2230);
xor U5741 (N_5741,N_124,N_3711);
nor U5742 (N_5742,N_4840,N_2772);
or U5743 (N_5743,N_2849,N_147);
and U5744 (N_5744,N_1233,N_4022);
nand U5745 (N_5745,N_4791,N_3390);
or U5746 (N_5746,N_1938,N_3616);
xor U5747 (N_5747,N_4094,N_4233);
nor U5748 (N_5748,N_1953,N_2871);
or U5749 (N_5749,N_1685,N_2332);
xor U5750 (N_5750,N_4608,N_1218);
or U5751 (N_5751,N_3925,N_4869);
and U5752 (N_5752,N_3510,N_2197);
or U5753 (N_5753,N_246,N_790);
and U5754 (N_5754,N_3768,N_2138);
nand U5755 (N_5755,N_2118,N_4336);
and U5756 (N_5756,N_4327,N_476);
and U5757 (N_5757,N_1468,N_3892);
nand U5758 (N_5758,N_4125,N_2193);
nand U5759 (N_5759,N_988,N_1571);
and U5760 (N_5760,N_4524,N_42);
and U5761 (N_5761,N_4558,N_268);
nor U5762 (N_5762,N_2177,N_4601);
or U5763 (N_5763,N_1487,N_230);
nor U5764 (N_5764,N_1193,N_47);
nor U5765 (N_5765,N_160,N_2571);
xor U5766 (N_5766,N_511,N_3629);
xnor U5767 (N_5767,N_2196,N_400);
nand U5768 (N_5768,N_3597,N_2344);
and U5769 (N_5769,N_4109,N_2011);
and U5770 (N_5770,N_3436,N_3375);
or U5771 (N_5771,N_2201,N_4044);
nand U5772 (N_5772,N_2669,N_1352);
xnor U5773 (N_5773,N_1360,N_1357);
or U5774 (N_5774,N_2021,N_4246);
xnor U5775 (N_5775,N_1817,N_3878);
or U5776 (N_5776,N_3652,N_2668);
xnor U5777 (N_5777,N_2079,N_4168);
and U5778 (N_5778,N_3332,N_2096);
nand U5779 (N_5779,N_4232,N_537);
xor U5780 (N_5780,N_2350,N_1101);
xor U5781 (N_5781,N_4364,N_1700);
nor U5782 (N_5782,N_3501,N_1103);
or U5783 (N_5783,N_3460,N_4747);
nor U5784 (N_5784,N_616,N_1698);
and U5785 (N_5785,N_4372,N_2721);
and U5786 (N_5786,N_1650,N_1242);
nand U5787 (N_5787,N_1482,N_4459);
nor U5788 (N_5788,N_3887,N_4303);
nand U5789 (N_5789,N_1766,N_3683);
and U5790 (N_5790,N_4748,N_1594);
or U5791 (N_5791,N_1137,N_4365);
and U5792 (N_5792,N_3347,N_1697);
or U5793 (N_5793,N_647,N_2467);
and U5794 (N_5794,N_198,N_3458);
or U5795 (N_5795,N_276,N_3186);
nor U5796 (N_5796,N_574,N_2667);
nand U5797 (N_5797,N_2464,N_4446);
or U5798 (N_5798,N_2259,N_2311);
or U5799 (N_5799,N_1092,N_1133);
or U5800 (N_5800,N_3769,N_2223);
nand U5801 (N_5801,N_204,N_4658);
or U5802 (N_5802,N_3827,N_1640);
nand U5803 (N_5803,N_3146,N_847);
nand U5804 (N_5804,N_2919,N_3043);
and U5805 (N_5805,N_3021,N_329);
or U5806 (N_5806,N_3214,N_3188);
xnor U5807 (N_5807,N_1703,N_1634);
and U5808 (N_5808,N_2927,N_3269);
xor U5809 (N_5809,N_3228,N_571);
nor U5810 (N_5810,N_3092,N_1872);
nor U5811 (N_5811,N_44,N_1346);
or U5812 (N_5812,N_1286,N_2590);
or U5813 (N_5813,N_3244,N_1299);
xnor U5814 (N_5814,N_2864,N_242);
nor U5815 (N_5815,N_369,N_126);
and U5816 (N_5816,N_3624,N_2428);
xnor U5817 (N_5817,N_3169,N_4920);
or U5818 (N_5818,N_4249,N_1904);
or U5819 (N_5819,N_376,N_1112);
nand U5820 (N_5820,N_4100,N_4443);
or U5821 (N_5821,N_3157,N_4492);
xnor U5822 (N_5822,N_258,N_4831);
xnor U5823 (N_5823,N_3555,N_2725);
nor U5824 (N_5824,N_1656,N_1359);
nor U5825 (N_5825,N_2995,N_2307);
nor U5826 (N_5826,N_3425,N_2562);
nand U5827 (N_5827,N_2409,N_2308);
xor U5828 (N_5828,N_3810,N_4829);
xnor U5829 (N_5829,N_2097,N_956);
nor U5830 (N_5830,N_4572,N_2922);
or U5831 (N_5831,N_2645,N_2841);
or U5832 (N_5832,N_3329,N_1705);
and U5833 (N_5833,N_2819,N_3093);
nand U5834 (N_5834,N_1796,N_1621);
and U5835 (N_5835,N_3070,N_3809);
and U5836 (N_5836,N_770,N_4873);
or U5837 (N_5837,N_189,N_1392);
xor U5838 (N_5838,N_1427,N_4160);
nand U5839 (N_5839,N_4034,N_2716);
nand U5840 (N_5840,N_4923,N_3153);
nor U5841 (N_5841,N_3184,N_3708);
xor U5842 (N_5842,N_2526,N_2381);
nor U5843 (N_5843,N_515,N_4813);
or U5844 (N_5844,N_4426,N_3772);
nand U5845 (N_5845,N_661,N_521);
xnor U5846 (N_5846,N_566,N_1461);
or U5847 (N_5847,N_4339,N_1837);
or U5848 (N_5848,N_222,N_1845);
nor U5849 (N_5849,N_4703,N_6);
nor U5850 (N_5850,N_603,N_2823);
xor U5851 (N_5851,N_2305,N_1187);
nand U5852 (N_5852,N_3570,N_1337);
or U5853 (N_5853,N_3396,N_2705);
nand U5854 (N_5854,N_2954,N_3098);
and U5855 (N_5855,N_2830,N_720);
or U5856 (N_5856,N_2860,N_722);
nor U5857 (N_5857,N_78,N_3819);
or U5858 (N_5858,N_1120,N_95);
or U5859 (N_5859,N_1504,N_2795);
or U5860 (N_5860,N_3143,N_3527);
or U5861 (N_5861,N_2565,N_3123);
xor U5862 (N_5862,N_1289,N_401);
or U5863 (N_5863,N_4916,N_941);
nor U5864 (N_5864,N_3534,N_2352);
xor U5865 (N_5865,N_3936,N_1480);
nand U5866 (N_5866,N_2677,N_2018);
nor U5867 (N_5867,N_3279,N_4029);
or U5868 (N_5868,N_1613,N_4690);
and U5869 (N_5869,N_4110,N_3079);
xnor U5870 (N_5870,N_4080,N_1958);
nand U5871 (N_5871,N_1319,N_1867);
nor U5872 (N_5872,N_3099,N_2161);
and U5873 (N_5873,N_764,N_3688);
nand U5874 (N_5874,N_4893,N_3282);
xor U5875 (N_5875,N_1100,N_1388);
and U5876 (N_5876,N_4046,N_2418);
or U5877 (N_5877,N_54,N_3431);
and U5878 (N_5878,N_2713,N_666);
xnor U5879 (N_5879,N_2990,N_390);
nor U5880 (N_5880,N_4464,N_3265);
or U5881 (N_5881,N_3163,N_1395);
nand U5882 (N_5882,N_2266,N_4850);
and U5883 (N_5883,N_3716,N_2131);
and U5884 (N_5884,N_556,N_1676);
and U5885 (N_5885,N_191,N_4595);
nor U5886 (N_5886,N_2758,N_3524);
nor U5887 (N_5887,N_2515,N_1370);
nor U5888 (N_5888,N_380,N_1879);
xnor U5889 (N_5889,N_932,N_4370);
nor U5890 (N_5890,N_4756,N_2543);
and U5891 (N_5891,N_3638,N_612);
or U5892 (N_5892,N_1345,N_3276);
nor U5893 (N_5893,N_1688,N_3424);
nor U5894 (N_5894,N_1041,N_2578);
and U5895 (N_5895,N_1877,N_2891);
xor U5896 (N_5896,N_2688,N_1767);
or U5897 (N_5897,N_2500,N_3133);
nand U5898 (N_5898,N_2976,N_524);
xor U5899 (N_5899,N_689,N_592);
nand U5900 (N_5900,N_2505,N_4523);
and U5901 (N_5901,N_4621,N_727);
or U5902 (N_5902,N_763,N_1213);
and U5903 (N_5903,N_4470,N_2277);
nor U5904 (N_5904,N_3556,N_4865);
nand U5905 (N_5905,N_1522,N_186);
nor U5906 (N_5906,N_1050,N_2817);
nand U5907 (N_5907,N_1509,N_1844);
or U5908 (N_5908,N_601,N_1428);
or U5909 (N_5909,N_484,N_3977);
or U5910 (N_5910,N_4452,N_2828);
xnor U5911 (N_5911,N_1161,N_445);
nor U5912 (N_5912,N_459,N_595);
nor U5913 (N_5913,N_3156,N_1991);
or U5914 (N_5914,N_3774,N_2798);
nand U5915 (N_5915,N_227,N_3755);
and U5916 (N_5916,N_1785,N_972);
nand U5917 (N_5917,N_3129,N_4622);
or U5918 (N_5918,N_3896,N_3967);
and U5919 (N_5919,N_779,N_974);
or U5920 (N_5920,N_2000,N_926);
nor U5921 (N_5921,N_2240,N_4980);
or U5922 (N_5922,N_2039,N_1843);
xor U5923 (N_5923,N_910,N_1224);
xor U5924 (N_5924,N_4310,N_1384);
nand U5925 (N_5925,N_4383,N_1252);
and U5926 (N_5926,N_3062,N_3419);
xor U5927 (N_5927,N_734,N_416);
nand U5928 (N_5928,N_2947,N_281);
nand U5929 (N_5929,N_1696,N_102);
nand U5930 (N_5930,N_1626,N_3317);
nand U5931 (N_5931,N_216,N_3148);
xor U5932 (N_5932,N_4577,N_3890);
nor U5933 (N_5933,N_3714,N_4961);
or U5934 (N_5934,N_1596,N_4421);
nand U5935 (N_5935,N_4380,N_1899);
and U5936 (N_5936,N_2246,N_3479);
or U5937 (N_5937,N_4041,N_2077);
nor U5938 (N_5938,N_957,N_4216);
nand U5939 (N_5939,N_3327,N_3593);
xnor U5940 (N_5940,N_2176,N_4215);
xnor U5941 (N_5941,N_3260,N_4381);
or U5942 (N_5942,N_3740,N_1209);
nor U5943 (N_5943,N_1566,N_4902);
nand U5944 (N_5944,N_435,N_1797);
nand U5945 (N_5945,N_4768,N_4333);
and U5946 (N_5946,N_3155,N_4450);
nand U5947 (N_5947,N_1423,N_2175);
or U5948 (N_5948,N_3442,N_2955);
nand U5949 (N_5949,N_929,N_2522);
nor U5950 (N_5950,N_2808,N_231);
nand U5951 (N_5951,N_2269,N_3728);
and U5952 (N_5952,N_4230,N_561);
or U5953 (N_5953,N_1153,N_3901);
nand U5954 (N_5954,N_2858,N_4521);
and U5955 (N_5955,N_3979,N_2933);
nand U5956 (N_5956,N_29,N_4794);
and U5957 (N_5957,N_2561,N_4194);
nor U5958 (N_5958,N_1387,N_3687);
and U5959 (N_5959,N_1315,N_4898);
nor U5960 (N_5960,N_2358,N_3434);
or U5961 (N_5961,N_1749,N_1314);
and U5962 (N_5962,N_3747,N_3197);
or U5963 (N_5963,N_4050,N_4801);
nand U5964 (N_5964,N_3466,N_156);
nand U5965 (N_5965,N_4954,N_232);
nand U5966 (N_5966,N_1339,N_4927);
xor U5967 (N_5967,N_3532,N_45);
or U5968 (N_5968,N_3409,N_4715);
nand U5969 (N_5969,N_183,N_1994);
nand U5970 (N_5970,N_839,N_3657);
nand U5971 (N_5971,N_3363,N_385);
nand U5972 (N_5972,N_3059,N_3058);
and U5973 (N_5973,N_935,N_2703);
and U5974 (N_5974,N_3203,N_1051);
nor U5975 (N_5975,N_743,N_3564);
or U5976 (N_5976,N_1008,N_782);
or U5977 (N_5977,N_2363,N_966);
and U5978 (N_5978,N_373,N_4390);
xor U5979 (N_5979,N_2433,N_3029);
or U5980 (N_5980,N_1719,N_4755);
or U5981 (N_5981,N_3366,N_4069);
nor U5982 (N_5982,N_351,N_3985);
and U5983 (N_5983,N_2770,N_2566);
or U5984 (N_5984,N_3757,N_742);
xnor U5985 (N_5985,N_1090,N_3830);
and U5986 (N_5986,N_3136,N_2181);
nand U5987 (N_5987,N_1924,N_3223);
and U5988 (N_5988,N_1232,N_1683);
or U5989 (N_5989,N_260,N_4555);
xnor U5990 (N_5990,N_3122,N_2962);
nand U5991 (N_5991,N_2872,N_4479);
nor U5992 (N_5992,N_370,N_3655);
or U5993 (N_5993,N_2687,N_1410);
or U5994 (N_5994,N_4097,N_2369);
and U5995 (N_5995,N_3312,N_4260);
xnor U5996 (N_5996,N_4670,N_2993);
nand U5997 (N_5997,N_2969,N_4605);
or U5998 (N_5998,N_4359,N_3224);
or U5999 (N_5999,N_3949,N_2481);
nand U6000 (N_6000,N_4474,N_470);
or U6001 (N_6001,N_990,N_1617);
xnor U6002 (N_6002,N_4674,N_3463);
nor U6003 (N_6003,N_4556,N_598);
nor U6004 (N_6004,N_576,N_1865);
xor U6005 (N_6005,N_138,N_2728);
nor U6006 (N_6006,N_1927,N_1902);
nor U6007 (N_6007,N_3902,N_1939);
nand U6008 (N_6008,N_1165,N_33);
nor U6009 (N_6009,N_3001,N_3730);
xnor U6010 (N_6010,N_626,N_2110);
or U6011 (N_6011,N_257,N_1069);
xnor U6012 (N_6012,N_2773,N_940);
xor U6013 (N_6013,N_729,N_4580);
xnor U6014 (N_6014,N_785,N_2258);
nor U6015 (N_6015,N_677,N_4130);
xor U6016 (N_6016,N_2503,N_2588);
or U6017 (N_6017,N_3849,N_4154);
nor U6018 (N_6018,N_4343,N_1284);
or U6019 (N_6019,N_217,N_4996);
xnor U6020 (N_6020,N_2101,N_4782);
or U6021 (N_6021,N_1225,N_3540);
nand U6022 (N_6022,N_4884,N_2086);
nand U6023 (N_6023,N_1201,N_4068);
and U6024 (N_6024,N_2646,N_1275);
and U6025 (N_6025,N_2806,N_843);
nor U6026 (N_6026,N_4561,N_4788);
and U6027 (N_6027,N_2321,N_1405);
nor U6028 (N_6028,N_4723,N_3437);
and U6029 (N_6029,N_2711,N_3009);
and U6030 (N_6030,N_2191,N_3482);
nand U6031 (N_6031,N_3523,N_3221);
nand U6032 (N_6032,N_4368,N_1429);
and U6033 (N_6033,N_2432,N_3180);
xor U6034 (N_6034,N_2710,N_122);
nor U6035 (N_6035,N_1323,N_3877);
or U6036 (N_6036,N_159,N_3378);
xor U6037 (N_6037,N_315,N_3218);
nor U6038 (N_6038,N_890,N_1025);
or U6039 (N_6039,N_391,N_510);
and U6040 (N_6040,N_3246,N_4115);
xor U6041 (N_6041,N_3599,N_2232);
or U6042 (N_6042,N_483,N_2631);
and U6043 (N_6043,N_2229,N_989);
nor U6044 (N_6044,N_4860,N_1975);
nor U6045 (N_6045,N_3812,N_2551);
nor U6046 (N_6046,N_4525,N_387);
and U6047 (N_6047,N_1874,N_1238);
nand U6048 (N_6048,N_4254,N_39);
and U6049 (N_6049,N_356,N_429);
nor U6050 (N_6050,N_4042,N_1791);
xnor U6051 (N_6051,N_2616,N_3698);
and U6052 (N_6052,N_4490,N_3036);
xor U6053 (N_6053,N_2137,N_2651);
xnor U6054 (N_6054,N_4699,N_360);
xnor U6055 (N_6055,N_1407,N_2002);
or U6056 (N_6056,N_986,N_3614);
xnor U6057 (N_6057,N_1419,N_368);
xor U6058 (N_6058,N_2434,N_1645);
and U6059 (N_6059,N_4892,N_2406);
and U6060 (N_6060,N_3646,N_4792);
nor U6061 (N_6061,N_963,N_468);
xnor U6062 (N_6062,N_2740,N_4837);
nor U6063 (N_6063,N_4905,N_716);
and U6064 (N_6064,N_3770,N_1850);
xnor U6065 (N_6065,N_4550,N_4743);
xnor U6066 (N_6066,N_218,N_633);
and U6067 (N_6067,N_4584,N_2569);
nand U6068 (N_6068,N_3999,N_531);
nand U6069 (N_6069,N_4348,N_219);
xnor U6070 (N_6070,N_1906,N_4214);
and U6071 (N_6071,N_2517,N_1631);
nand U6072 (N_6072,N_1021,N_3633);
nand U6073 (N_6073,N_1185,N_406);
and U6074 (N_6074,N_4040,N_2473);
nor U6075 (N_6075,N_568,N_3387);
and U6076 (N_6076,N_1303,N_2377);
nand U6077 (N_6077,N_706,N_4719);
and U6078 (N_6078,N_3886,N_4967);
and U6079 (N_6079,N_3891,N_1901);
nor U6080 (N_6080,N_3797,N_1136);
or U6081 (N_6081,N_2455,N_2339);
and U6082 (N_6082,N_3255,N_2236);
nor U6083 (N_6083,N_1731,N_4427);
nor U6084 (N_6084,N_1355,N_1605);
xnor U6085 (N_6085,N_49,N_2456);
nor U6086 (N_6086,N_50,N_325);
nor U6087 (N_6087,N_3205,N_1282);
nand U6088 (N_6088,N_313,N_3948);
or U6089 (N_6089,N_3918,N_1119);
or U6090 (N_6090,N_685,N_866);
and U6091 (N_6091,N_262,N_403);
or U6092 (N_6092,N_4410,N_2372);
nor U6093 (N_6093,N_590,N_2730);
xor U6094 (N_6094,N_2419,N_3664);
and U6095 (N_6095,N_710,N_1986);
or U6096 (N_6096,N_4666,N_2791);
xnor U6097 (N_6097,N_2082,N_2680);
or U6098 (N_6098,N_1318,N_4919);
or U6099 (N_6099,N_875,N_1174);
nand U6100 (N_6100,N_901,N_2536);
xor U6101 (N_6101,N_3489,N_3717);
nor U6102 (N_6102,N_23,N_2164);
or U6103 (N_6103,N_4804,N_256);
xor U6104 (N_6104,N_2120,N_475);
nor U6105 (N_6105,N_3908,N_3454);
nand U6106 (N_6106,N_4764,N_2672);
and U6107 (N_6107,N_2685,N_2050);
or U6108 (N_6108,N_667,N_3702);
and U6109 (N_6109,N_2747,N_865);
and U6110 (N_6110,N_4895,N_3113);
xnor U6111 (N_6111,N_3839,N_1869);
nand U6112 (N_6112,N_4102,N_2525);
or U6113 (N_6113,N_1884,N_1538);
or U6114 (N_6114,N_2763,N_4226);
nor U6115 (N_6115,N_1104,N_4736);
and U6116 (N_6116,N_1589,N_3152);
xor U6117 (N_6117,N_4304,N_3632);
xnor U6118 (N_6118,N_4411,N_1585);
and U6119 (N_6119,N_831,N_3421);
and U6120 (N_6120,N_868,N_3798);
or U6121 (N_6121,N_3859,N_1087);
xor U6122 (N_6122,N_937,N_3020);
xnor U6123 (N_6123,N_4458,N_4313);
and U6124 (N_6124,N_3590,N_2139);
nor U6125 (N_6125,N_3045,N_4552);
and U6126 (N_6126,N_622,N_451);
nor U6127 (N_6127,N_1774,N_3467);
and U6128 (N_6128,N_4776,N_1249);
or U6129 (N_6129,N_2146,N_2936);
nand U6130 (N_6130,N_3368,N_3881);
xor U6131 (N_6131,N_1932,N_3137);
and U6132 (N_6132,N_1736,N_629);
or U6133 (N_6133,N_2575,N_3090);
nor U6134 (N_6134,N_453,N_3584);
or U6135 (N_6135,N_3284,N_1861);
or U6136 (N_6136,N_1513,N_2262);
and U6137 (N_6137,N_4573,N_3210);
or U6138 (N_6138,N_4338,N_58);
nand U6139 (N_6139,N_2626,N_18);
or U6140 (N_6140,N_2444,N_1351);
nand U6141 (N_6141,N_1556,N_1805);
and U6142 (N_6142,N_290,N_4281);
nand U6143 (N_6143,N_2941,N_133);
nor U6144 (N_6144,N_195,N_1181);
and U6145 (N_6145,N_3240,N_4147);
xnor U6146 (N_6146,N_4401,N_2247);
xnor U6147 (N_6147,N_3713,N_2816);
nor U6148 (N_6148,N_3040,N_4943);
or U6149 (N_6149,N_1326,N_4429);
or U6150 (N_6150,N_4823,N_1106);
or U6151 (N_6151,N_3834,N_714);
nand U6152 (N_6152,N_4043,N_4309);
nand U6153 (N_6153,N_749,N_104);
and U6154 (N_6154,N_2905,N_3309);
nand U6155 (N_6155,N_3589,N_3168);
or U6156 (N_6156,N_3793,N_3016);
nand U6157 (N_6157,N_3928,N_2257);
or U6158 (N_6158,N_2845,N_588);
nor U6159 (N_6159,N_409,N_3235);
or U6160 (N_6160,N_3449,N_168);
or U6161 (N_6161,N_2878,N_3653);
and U6162 (N_6162,N_981,N_1002);
xor U6163 (N_6163,N_4751,N_3791);
xor U6164 (N_6164,N_4795,N_2166);
nand U6165 (N_6165,N_3617,N_4526);
nor U6166 (N_6166,N_3685,N_4718);
and U6167 (N_6167,N_3691,N_2909);
nand U6168 (N_6168,N_184,N_2494);
and U6169 (N_6169,N_462,N_1829);
nor U6170 (N_6170,N_4581,N_4812);
xor U6171 (N_6171,N_1742,N_1347);
nor U6172 (N_6172,N_275,N_3642);
nand U6173 (N_6173,N_1699,N_1228);
nand U6174 (N_6174,N_1311,N_3050);
nor U6175 (N_6175,N_3377,N_4686);
nand U6176 (N_6176,N_2585,N_4405);
or U6177 (N_6177,N_4066,N_2371);
xor U6178 (N_6178,N_2376,N_4560);
nand U6179 (N_6179,N_1757,N_2897);
and U6180 (N_6180,N_3484,N_188);
and U6181 (N_6181,N_2846,N_2198);
nand U6182 (N_6182,N_2004,N_2793);
and U6183 (N_6183,N_489,N_594);
and U6184 (N_6184,N_4870,N_525);
xnor U6185 (N_6185,N_3835,N_2696);
or U6186 (N_6186,N_3031,N_4571);
and U6187 (N_6187,N_1422,N_748);
nand U6188 (N_6188,N_3364,N_2857);
nor U6189 (N_6189,N_4112,N_752);
xor U6190 (N_6190,N_1371,N_530);
nor U6191 (N_6191,N_3821,N_1343);
and U6192 (N_6192,N_1581,N_505);
nor U6193 (N_6193,N_4134,N_2971);
or U6194 (N_6194,N_808,N_4668);
nand U6195 (N_6195,N_238,N_527);
xor U6196 (N_6196,N_563,N_1389);
nand U6197 (N_6197,N_1952,N_2501);
nand U6198 (N_6198,N_3814,N_3700);
nor U6199 (N_6199,N_2210,N_2291);
xor U6200 (N_6200,N_4035,N_4633);
xnor U6201 (N_6201,N_859,N_69);
nor U6202 (N_6202,N_4378,N_4936);
and U6203 (N_6203,N_3508,N_1668);
nand U6204 (N_6204,N_4064,N_2794);
and U6205 (N_6205,N_2080,N_652);
nand U6206 (N_6206,N_3173,N_3579);
or U6207 (N_6207,N_2931,N_700);
nor U6208 (N_6208,N_719,N_805);
nor U6209 (N_6209,N_4126,N_2117);
nor U6210 (N_6210,N_1365,N_2867);
nand U6211 (N_6211,N_2564,N_3410);
and U6212 (N_6212,N_3879,N_1961);
and U6213 (N_6213,N_2949,N_4696);
nor U6214 (N_6214,N_43,N_31);
nand U6215 (N_6215,N_917,N_1024);
or U6216 (N_6216,N_4496,N_14);
nor U6217 (N_6217,N_2405,N_1129);
nor U6218 (N_6218,N_3278,N_1553);
nor U6219 (N_6219,N_2104,N_1770);
xor U6220 (N_6220,N_2023,N_332);
and U6221 (N_6221,N_1951,N_2924);
xor U6222 (N_6222,N_2985,N_534);
nor U6223 (N_6223,N_1203,N_4664);
or U6224 (N_6224,N_4908,N_2280);
or U6225 (N_6225,N_444,N_4278);
and U6226 (N_6226,N_701,N_675);
nor U6227 (N_6227,N_3496,N_4311);
or U6228 (N_6228,N_1000,N_4539);
xnor U6229 (N_6229,N_2147,N_3094);
nand U6230 (N_6230,N_1999,N_4434);
nand U6231 (N_6231,N_2953,N_1740);
nor U6232 (N_6232,N_2028,N_1147);
nand U6233 (N_6233,N_2342,N_2691);
and U6234 (N_6234,N_562,N_4271);
xor U6235 (N_6235,N_4342,N_2737);
or U6236 (N_6236,N_4124,N_2303);
or U6237 (N_6237,N_4611,N_3725);
or U6238 (N_6238,N_1543,N_2485);
and U6239 (N_6239,N_715,N_1693);
and U6240 (N_6240,N_1863,N_2057);
xnor U6241 (N_6241,N_4397,N_2958);
or U6242 (N_6242,N_1662,N_4656);
nor U6243 (N_6243,N_2207,N_3895);
nand U6244 (N_6244,N_2390,N_4489);
and U6245 (N_6245,N_397,N_312);
nand U6246 (N_6246,N_2582,N_3625);
and U6247 (N_6247,N_2577,N_3643);
nand U6248 (N_6248,N_955,N_1334);
and U6249 (N_6249,N_2991,N_2521);
nor U6250 (N_6250,N_1123,N_4329);
nor U6251 (N_6251,N_1267,N_4353);
and U6252 (N_6252,N_1755,N_4774);
or U6253 (N_6253,N_3357,N_4528);
or U6254 (N_6254,N_2479,N_4167);
nor U6255 (N_6255,N_4693,N_3423);
and U6256 (N_6256,N_3158,N_4173);
or U6257 (N_6257,N_3546,N_1498);
xnor U6258 (N_6258,N_1118,N_2324);
or U6259 (N_6259,N_1570,N_1117);
xor U6260 (N_6260,N_1102,N_3932);
xor U6261 (N_6261,N_4096,N_1714);
or U6262 (N_6262,N_3743,N_415);
and U6263 (N_6263,N_1246,N_1164);
or U6264 (N_6264,N_4516,N_3149);
xor U6265 (N_6265,N_3292,N_4846);
or U6266 (N_6266,N_1800,N_2276);
or U6267 (N_6267,N_1449,N_2469);
nand U6268 (N_6268,N_4727,N_4742);
and U6269 (N_6269,N_2731,N_4655);
nor U6270 (N_6270,N_589,N_1560);
and U6271 (N_6271,N_4273,N_2200);
and U6272 (N_6272,N_3211,N_4116);
nand U6273 (N_6273,N_2250,N_3164);
and U6274 (N_6274,N_953,N_2840);
and U6275 (N_6275,N_2385,N_695);
nor U6276 (N_6276,N_2843,N_331);
and U6277 (N_6277,N_1058,N_105);
nand U6278 (N_6278,N_2446,N_2424);
or U6279 (N_6279,N_2987,N_2608);
nand U6280 (N_6280,N_3969,N_1085);
nand U6281 (N_6281,N_1769,N_3621);
or U6282 (N_6282,N_684,N_398);
nor U6283 (N_6283,N_1042,N_4587);
xnor U6284 (N_6284,N_2655,N_1783);
xnor U6285 (N_6285,N_969,N_1733);
and U6286 (N_6286,N_1167,N_3862);
nand U6287 (N_6287,N_3349,N_3675);
and U6288 (N_6288,N_1673,N_1448);
xnor U6289 (N_6289,N_4913,N_3441);
or U6290 (N_6290,N_395,N_4720);
or U6291 (N_6291,N_3790,N_1398);
and U6292 (N_6292,N_1471,N_570);
and U6293 (N_6293,N_3968,N_2359);
nor U6294 (N_6294,N_558,N_284);
nand U6295 (N_6295,N_4276,N_776);
or U6296 (N_6296,N_2251,N_3362);
and U6297 (N_6297,N_1964,N_842);
or U6298 (N_6298,N_4513,N_2306);
and U6299 (N_6299,N_2242,N_4242);
xor U6300 (N_6300,N_4237,N_4985);
nor U6301 (N_6301,N_518,N_709);
nor U6302 (N_6302,N_3189,N_4355);
nand U6303 (N_6303,N_1825,N_2788);
or U6304 (N_6304,N_1329,N_3739);
nand U6305 (N_6305,N_2279,N_3626);
nand U6306 (N_6306,N_491,N_1530);
xnor U6307 (N_6307,N_4532,N_2071);
nor U6308 (N_6308,N_4527,N_3414);
and U6309 (N_6309,N_754,N_1432);
and U6310 (N_6310,N_3661,N_3531);
or U6311 (N_6311,N_939,N_3042);
and U6312 (N_6312,N_2910,N_887);
nand U6313 (N_6313,N_4155,N_3166);
or U6314 (N_6314,N_851,N_1397);
or U6315 (N_6315,N_244,N_2837);
xor U6316 (N_6316,N_4453,N_210);
or U6317 (N_6317,N_998,N_2766);
and U6318 (N_6318,N_4486,N_765);
or U6319 (N_6319,N_2112,N_2045);
or U6320 (N_6320,N_2027,N_4934);
and U6321 (N_6321,N_4212,N_1638);
xnor U6322 (N_6322,N_4531,N_761);
xor U6323 (N_6323,N_2069,N_881);
or U6324 (N_6324,N_2084,N_4989);
and U6325 (N_6325,N_1954,N_4735);
and U6326 (N_6326,N_3355,N_4864);
nor U6327 (N_6327,N_4906,N_3256);
nand U6328 (N_6328,N_1399,N_4473);
or U6329 (N_6329,N_2876,N_3051);
nor U6330 (N_6330,N_4749,N_4753);
and U6331 (N_6331,N_4152,N_2978);
and U6332 (N_6332,N_3019,N_2863);
and U6333 (N_6333,N_519,N_4190);
xor U6334 (N_6334,N_1963,N_1532);
and U6335 (N_6335,N_920,N_1099);
nand U6336 (N_6336,N_110,N_4659);
or U6337 (N_6337,N_2752,N_975);
or U6338 (N_6338,N_3933,N_2592);
nor U6339 (N_6339,N_3966,N_564);
nor U6340 (N_6340,N_2243,N_4484);
or U6341 (N_6341,N_739,N_2329);
and U6342 (N_6342,N_2765,N_1627);
nor U6343 (N_6343,N_4499,N_3461);
xnor U6344 (N_6344,N_2935,N_1);
xor U6345 (N_6345,N_642,N_1646);
nand U6346 (N_6346,N_2999,N_4191);
and U6347 (N_6347,N_2901,N_575);
or U6348 (N_6348,N_4179,N_2205);
or U6349 (N_6349,N_3145,N_1619);
xor U6350 (N_6350,N_1870,N_1266);
xor U6351 (N_6351,N_3103,N_19);
or U6352 (N_6352,N_2506,N_1003);
and U6353 (N_6353,N_3888,N_4013);
and U6354 (N_6354,N_252,N_4683);
nand U6355 (N_6355,N_1302,N_4266);
nand U6356 (N_6356,N_2528,N_335);
nor U6357 (N_6357,N_3022,N_4889);
nor U6358 (N_6358,N_4177,N_4288);
or U6359 (N_6359,N_4379,N_573);
nor U6360 (N_6360,N_3039,N_4878);
or U6361 (N_6361,N_1667,N_4350);
and U6362 (N_6362,N_3843,N_3193);
and U6363 (N_6363,N_4711,N_1960);
and U6364 (N_6364,N_323,N_638);
and U6365 (N_6365,N_4170,N_1670);
or U6366 (N_6366,N_3541,N_1689);
nand U6367 (N_6367,N_4682,N_1168);
nor U6368 (N_6368,N_3575,N_921);
xnor U6369 (N_6369,N_924,N_4207);
or U6370 (N_6370,N_3678,N_1561);
or U6371 (N_6371,N_3393,N_4344);
nand U6372 (N_6372,N_3487,N_760);
nand U6373 (N_6373,N_1489,N_767);
xnor U6374 (N_6374,N_2674,N_1494);
nand U6375 (N_6375,N_73,N_2973);
or U6376 (N_6376,N_2529,N_582);
nor U6377 (N_6377,N_1992,N_1486);
and U6378 (N_6378,N_1274,N_3995);
nor U6379 (N_6379,N_15,N_3503);
nor U6380 (N_6380,N_1206,N_3207);
or U6381 (N_6381,N_1944,N_2544);
or U6382 (N_6382,N_3141,N_4430);
or U6383 (N_6383,N_3231,N_3388);
xnor U6384 (N_6384,N_4510,N_4563);
xor U6385 (N_6385,N_443,N_4395);
nor U6386 (N_6386,N_2064,N_3297);
xnor U6387 (N_6387,N_4014,N_1819);
xor U6388 (N_6388,N_2764,N_4662);
nand U6389 (N_6389,N_4600,N_1496);
and U6390 (N_6390,N_3538,N_3065);
xor U6391 (N_6391,N_3951,N_1548);
and U6392 (N_6392,N_4672,N_3300);
xor U6393 (N_6393,N_1381,N_419);
xnor U6394 (N_6394,N_4150,N_2635);
nor U6395 (N_6395,N_4180,N_2604);
xor U6396 (N_6396,N_2960,N_555);
and U6397 (N_6397,N_3504,N_1235);
xnor U6398 (N_6398,N_3096,N_872);
nor U6399 (N_6399,N_1982,N_215);
xor U6400 (N_6400,N_4055,N_2227);
nand U6401 (N_6401,N_1033,N_1464);
nand U6402 (N_6402,N_1115,N_1718);
and U6403 (N_6403,N_4783,N_3826);
xor U6404 (N_6404,N_707,N_3974);
xnor U6405 (N_6405,N_1592,N_4205);
nor U6406 (N_6406,N_2756,N_4635);
xor U6407 (N_6407,N_2707,N_4287);
and U6408 (N_6408,N_1601,N_11);
and U6409 (N_6409,N_314,N_4772);
xor U6410 (N_6410,N_3666,N_3926);
nor U6411 (N_6411,N_2490,N_1276);
or U6412 (N_6412,N_4626,N_3379);
xor U6413 (N_6413,N_420,N_2108);
and U6414 (N_6414,N_826,N_3560);
or U6415 (N_6415,N_4949,N_1086);
and U6416 (N_6416,N_4121,N_2533);
xor U6417 (N_6417,N_209,N_38);
and U6418 (N_6418,N_3628,N_1790);
and U6419 (N_6419,N_41,N_2216);
xnor U6420 (N_6420,N_1204,N_497);
nand U6421 (N_6421,N_4729,N_4928);
nand U6422 (N_6422,N_4606,N_2388);
nand U6423 (N_6423,N_1923,N_2202);
and U6424 (N_6424,N_4915,N_4590);
xnor U6425 (N_6425,N_4021,N_2411);
nand U6426 (N_6426,N_1081,N_3993);
nor U6427 (N_6427,N_76,N_438);
nand U6428 (N_6428,N_4990,N_139);
xnor U6429 (N_6429,N_4093,N_4366);
or U6430 (N_6430,N_1273,N_1882);
nand U6431 (N_6431,N_2852,N_4262);
and U6432 (N_6432,N_962,N_2233);
nor U6433 (N_6433,N_4352,N_279);
nand U6434 (N_6434,N_144,N_2548);
or U6435 (N_6435,N_1059,N_3631);
xor U6436 (N_6436,N_3929,N_747);
nor U6437 (N_6437,N_3320,N_3938);
xnor U6438 (N_6438,N_3302,N_2885);
and U6439 (N_6439,N_339,N_1336);
xor U6440 (N_6440,N_1396,N_3750);
nand U6441 (N_6441,N_2537,N_830);
nand U6442 (N_6442,N_4691,N_1838);
nor U6443 (N_6443,N_1222,N_3745);
or U6444 (N_6444,N_3815,N_3151);
and U6445 (N_6445,N_604,N_1995);
xor U6446 (N_6446,N_3876,N_4937);
and U6447 (N_6447,N_3873,N_3906);
nand U6448 (N_6448,N_4542,N_1860);
nor U6449 (N_6449,N_1798,N_4038);
nor U6450 (N_6450,N_1873,N_2001);
nor U6451 (N_6451,N_2980,N_3291);
xnor U6452 (N_6452,N_3588,N_4849);
or U6453 (N_6453,N_4740,N_3997);
and U6454 (N_6454,N_3723,N_3864);
and U6455 (N_6455,N_1066,N_3581);
nor U6456 (N_6456,N_2322,N_4612);
xor U6457 (N_6457,N_4844,N_3271);
xnor U6458 (N_6458,N_3694,N_1026);
or U6459 (N_6459,N_3111,N_3361);
or U6460 (N_6460,N_4224,N_2375);
nor U6461 (N_6461,N_346,N_1074);
nor U6462 (N_6462,N_4839,N_1709);
and U6463 (N_6463,N_2106,N_1162);
nor U6464 (N_6464,N_213,N_4261);
xor U6465 (N_6465,N_4815,N_697);
and U6466 (N_6466,N_4073,N_4883);
xor U6467 (N_6467,N_4011,N_2751);
or U6468 (N_6468,N_3225,N_4178);
or U6469 (N_6469,N_4286,N_4472);
nand U6470 (N_6470,N_1756,N_2180);
nand U6471 (N_6471,N_1831,N_533);
xnor U6472 (N_6472,N_2396,N_536);
nor U6473 (N_6473,N_2496,N_852);
xor U6474 (N_6474,N_3547,N_3476);
or U6475 (N_6475,N_4206,N_1655);
nor U6476 (N_6476,N_261,N_3709);
or U6477 (N_6477,N_1534,N_2085);
xnor U6478 (N_6478,N_2633,N_1141);
or U6479 (N_6479,N_1184,N_2579);
nand U6480 (N_6480,N_2425,N_3738);
nor U6481 (N_6481,N_639,N_1416);
and U6482 (N_6482,N_4349,N_280);
nand U6483 (N_6483,N_774,N_2111);
nor U6484 (N_6484,N_3359,N_1178);
xor U6485 (N_6485,N_1244,N_3818);
nor U6486 (N_6486,N_3422,N_3179);
or U6487 (N_6487,N_4065,N_2334);
and U6488 (N_6488,N_501,N_2029);
nor U6489 (N_6489,N_2272,N_150);
xnor U6490 (N_6490,N_2136,N_4917);
nand U6491 (N_6491,N_3348,N_190);
xor U6492 (N_6492,N_367,N_2263);
nand U6493 (N_6493,N_3220,N_1259);
or U6494 (N_6494,N_2288,N_2760);
xor U6495 (N_6495,N_4412,N_3444);
or U6496 (N_6496,N_4901,N_4164);
and U6497 (N_6497,N_2967,N_3618);
and U6498 (N_6498,N_4113,N_4565);
nand U6499 (N_6499,N_4533,N_2510);
xor U6500 (N_6500,N_3515,N_2739);
xor U6501 (N_6501,N_4377,N_2130);
nand U6502 (N_6502,N_3274,N_46);
xnor U6503 (N_6503,N_2182,N_725);
and U6504 (N_6504,N_2234,N_1659);
or U6505 (N_6505,N_295,N_4994);
xnor U6506 (N_6506,N_3391,N_3600);
xnor U6507 (N_6507,N_2809,N_1762);
or U6508 (N_6508,N_1576,N_2929);
and U6509 (N_6509,N_3015,N_894);
xor U6510 (N_6510,N_2488,N_1192);
xor U6511 (N_6511,N_3078,N_3921);
nand U6512 (N_6512,N_1810,N_4576);
nand U6513 (N_6513,N_1799,N_4335);
nand U6514 (N_6514,N_2873,N_4541);
or U6515 (N_6515,N_4798,N_1763);
nand U6516 (N_6516,N_4564,N_4076);
or U6517 (N_6517,N_2460,N_48);
xnor U6518 (N_6518,N_2584,N_3046);
nor U6519 (N_6519,N_3619,N_640);
or U6520 (N_6520,N_1215,N_792);
and U6521 (N_6521,N_90,N_0);
nand U6522 (N_6522,N_3147,N_2662);
xnor U6523 (N_6523,N_1983,N_3177);
nand U6524 (N_6524,N_931,N_1728);
xnor U6525 (N_6525,N_1288,N_4145);
nand U6526 (N_6526,N_2319,N_1894);
nor U6527 (N_6527,N_4183,N_3490);
nor U6528 (N_6528,N_1729,N_3851);
nor U6529 (N_6529,N_4517,N_2241);
and U6530 (N_6530,N_4471,N_1393);
xor U6531 (N_6531,N_1604,N_3311);
xnor U6532 (N_6532,N_2059,N_1822);
xor U6533 (N_6533,N_4939,N_146);
nor U6534 (N_6534,N_2966,N_724);
and U6535 (N_6535,N_1814,N_307);
and U6536 (N_6536,N_1775,N_3464);
or U6537 (N_6537,N_2374,N_2519);
and U6538 (N_6538,N_741,N_928);
and U6539 (N_6539,N_1063,N_458);
xor U6540 (N_6540,N_239,N_662);
or U6541 (N_6541,N_2665,N_2783);
or U6542 (N_6542,N_3697,N_4888);
xor U6543 (N_6543,N_2360,N_786);
nor U6544 (N_6544,N_3856,N_2357);
or U6545 (N_6545,N_1364,N_4498);
xnor U6546 (N_6546,N_3301,N_1830);
or U6547 (N_6547,N_4297,N_4199);
nor U6548 (N_6548,N_4087,N_1515);
nor U6549 (N_6549,N_2888,N_2192);
and U6550 (N_6550,N_1474,N_559);
and U6551 (N_6551,N_4504,N_2940);
nor U6552 (N_6552,N_2462,N_265);
and U6553 (N_6553,N_4131,N_4692);
nand U6554 (N_6554,N_907,N_1043);
nand U6555 (N_6555,N_2062,N_2679);
xor U6556 (N_6556,N_1883,N_3561);
and U6557 (N_6557,N_1564,N_2774);
or U6558 (N_6558,N_3836,N_2921);
nand U6559 (N_6559,N_4221,N_4201);
xnor U6560 (N_6560,N_2555,N_4854);
nor U6561 (N_6561,N_4761,N_3405);
nand U6562 (N_6562,N_4274,N_413);
and U6563 (N_6563,N_3680,N_2512);
or U6564 (N_6564,N_1172,N_2498);
or U6565 (N_6565,N_3958,N_3550);
and U6566 (N_6566,N_1658,N_485);
or U6567 (N_6567,N_4174,N_2040);
nand U6568 (N_6568,N_1163,N_51);
or U6569 (N_6569,N_2351,N_2620);
nand U6570 (N_6570,N_2648,N_2480);
nand U6571 (N_6571,N_1320,N_4382);
or U6572 (N_6572,N_683,N_1628);
and U6573 (N_6573,N_2914,N_3742);
xor U6574 (N_6574,N_2148,N_3038);
or U6575 (N_6575,N_2656,N_4614);
nor U6576 (N_6576,N_1277,N_2056);
or U6577 (N_6577,N_2689,N_473);
or U6578 (N_6578,N_4619,N_2218);
or U6579 (N_6579,N_1629,N_744);
and U6580 (N_6580,N_3897,N_1527);
nand U6581 (N_6581,N_226,N_2282);
xnor U6582 (N_6582,N_509,N_597);
or U6583 (N_6583,N_809,N_350);
and U6584 (N_6584,N_187,N_3335);
xor U6585 (N_6585,N_1417,N_4586);
nor U6586 (N_6586,N_3727,N_4334);
nand U6587 (N_6587,N_1295,N_1611);
or U6588 (N_6588,N_253,N_4059);
nand U6589 (N_6589,N_3402,N_772);
and U6590 (N_6590,N_1897,N_120);
and U6591 (N_6591,N_4641,N_2934);
nor U6592 (N_6592,N_781,N_5);
nor U6593 (N_6593,N_1499,N_4731);
and U6594 (N_6594,N_659,N_3328);
and U6595 (N_6595,N_4469,N_4636);
nor U6596 (N_6596,N_1826,N_4373);
or U6597 (N_6597,N_1524,N_3662);
and U6598 (N_6598,N_4402,N_145);
xor U6599 (N_6599,N_1842,N_1660);
xor U6600 (N_6600,N_3115,N_540);
xor U6601 (N_6601,N_2068,N_3511);
xnor U6602 (N_6602,N_1652,N_2647);
nor U6603 (N_6603,N_3132,N_1647);
nor U6604 (N_6604,N_1442,N_3960);
nand U6605 (N_6605,N_1593,N_3475);
or U6606 (N_6606,N_2034,N_2133);
nand U6607 (N_6607,N_4800,N_4821);
or U6608 (N_6608,N_3822,N_876);
nor U6609 (N_6609,N_271,N_430);
or U6610 (N_6610,N_1027,N_4781);
or U6611 (N_6611,N_1555,N_4156);
and U6612 (N_6612,N_3767,N_4070);
nand U6613 (N_6613,N_4646,N_3686);
and U6614 (N_6614,N_3943,N_1748);
xor U6615 (N_6615,N_3957,N_532);
or U6616 (N_6616,N_2046,N_2483);
nand U6617 (N_6617,N_2844,N_4569);
xnor U6618 (N_6618,N_2478,N_4475);
and U6619 (N_6619,N_4976,N_2796);
and U6620 (N_6620,N_900,N_1758);
nand U6621 (N_6621,N_1015,N_2963);
or U6622 (N_6622,N_1813,N_3762);
nand U6623 (N_6623,N_3025,N_4824);
nor U6624 (N_6624,N_254,N_477);
nand U6625 (N_6625,N_3060,N_3296);
nor U6626 (N_6626,N_1608,N_3934);
and U6627 (N_6627,N_4062,N_4536);
and U6628 (N_6628,N_971,N_3069);
nor U6629 (N_6629,N_1490,N_1412);
xnor U6630 (N_6630,N_93,N_3894);
nor U6631 (N_6631,N_1331,N_3413);
or U6632 (N_6632,N_3273,N_2414);
and U6633 (N_6633,N_1330,N_3226);
nand U6634 (N_6634,N_3448,N_3912);
xnor U6635 (N_6635,N_663,N_2545);
or U6636 (N_6636,N_3107,N_4165);
or U6637 (N_6637,N_4651,N_4056);
nor U6638 (N_6638,N_2507,N_541);
xnor U6639 (N_6639,N_3916,N_2486);
nor U6640 (N_6640,N_2047,N_611);
nor U6641 (N_6641,N_902,N_3088);
xnor U6642 (N_6642,N_4258,N_1456);
nand U6643 (N_6643,N_1895,N_2826);
or U6644 (N_6644,N_1684,N_2615);
and U6645 (N_6645,N_3701,N_82);
xnor U6646 (N_6646,N_1942,N_2341);
and U6647 (N_6647,N_1134,N_2974);
xnor U6648 (N_6648,N_3552,N_1415);
or U6649 (N_6649,N_319,N_2477);
and U6650 (N_6650,N_310,N_1801);
or U6651 (N_6651,N_4016,N_3430);
or U6652 (N_6652,N_3634,N_2595);
xnor U6653 (N_6653,N_3521,N_1803);
nor U6654 (N_6654,N_2320,N_4431);
nand U6655 (N_6655,N_3406,N_2267);
nor U6656 (N_6656,N_2186,N_658);
nand U6657 (N_6657,N_3196,N_4460);
nand U6658 (N_6658,N_1447,N_807);
and U6659 (N_6659,N_857,N_2470);
xor U6660 (N_6660,N_1989,N_627);
nand U6661 (N_6661,N_4247,N_70);
nor U6662 (N_6662,N_580,N_1743);
nor U6663 (N_6663,N_4136,N_1815);
or U6664 (N_6664,N_1052,N_3248);
nor U6665 (N_6665,N_942,N_4285);
and U6666 (N_6666,N_4955,N_1500);
nor U6667 (N_6667,N_2330,N_1746);
xnor U6668 (N_6668,N_2879,N_3215);
or U6669 (N_6669,N_644,N_2898);
and U6670 (N_6670,N_693,N_1614);
nand U6671 (N_6671,N_2563,N_3330);
xnor U6672 (N_6672,N_467,N_2895);
nand U6673 (N_6673,N_1073,N_905);
xor U6674 (N_6674,N_3380,N_3304);
xor U6675 (N_6675,N_2779,N_3965);
xnor U6676 (N_6676,N_583,N_3850);
or U6677 (N_6677,N_547,N_1540);
or U6678 (N_6678,N_1636,N_321);
nor U6679 (N_6679,N_1237,N_228);
xnor U6680 (N_6680,N_650,N_4634);
nand U6681 (N_6681,N_4763,N_947);
and U6682 (N_6682,N_4416,N_92);
nor U6683 (N_6683,N_1726,N_624);
nor U6684 (N_6684,N_3287,N_1738);
or U6685 (N_6685,N_4497,N_1019);
or U6686 (N_6686,N_2132,N_4151);
xnor U6687 (N_6687,N_758,N_3671);
xor U6688 (N_6688,N_619,N_197);
nor U6689 (N_6689,N_52,N_3602);
or U6690 (N_6690,N_1828,N_2215);
nand U6691 (N_6691,N_2812,N_2410);
xor U6692 (N_6692,N_2074,N_3154);
xnor U6693 (N_6693,N_440,N_2746);
or U6694 (N_6694,N_1171,N_1692);
xnor U6695 (N_6695,N_1253,N_3120);
and U6696 (N_6696,N_819,N_3026);
xor U6697 (N_6697,N_2911,N_2260);
xnor U6698 (N_6698,N_504,N_4045);
nor U6699 (N_6699,N_3027,N_3018);
nor U6700 (N_6700,N_4414,N_3654);
nand U6701 (N_6701,N_1376,N_1878);
and U6702 (N_6702,N_4987,N_3703);
nor U6703 (N_6703,N_960,N_2702);
and U6704 (N_6704,N_585,N_1272);
nand U6705 (N_6705,N_106,N_1910);
xnor U6706 (N_6706,N_2709,N_2664);
nand U6707 (N_6707,N_1980,N_3470);
nand U6708 (N_6708,N_2970,N_3935);
xor U6709 (N_6709,N_3720,N_3447);
nand U6710 (N_6710,N_983,N_2048);
nor U6711 (N_6711,N_97,N_4204);
xor U6712 (N_6712,N_1682,N_2349);
nor U6713 (N_6713,N_3576,N_3913);
nand U6714 (N_6714,N_512,N_4398);
or U6715 (N_6715,N_2173,N_3914);
or U6716 (N_6716,N_2487,N_402);
xor U6717 (N_6717,N_651,N_1009);
nor U6718 (N_6718,N_4616,N_3117);
nor U6719 (N_6719,N_1654,N_1077);
xor U6720 (N_6720,N_4970,N_118);
nor U6721 (N_6721,N_2098,N_2785);
nor U6722 (N_6722,N_4593,N_1794);
and U6723 (N_6723,N_4091,N_3445);
or U6724 (N_6724,N_4631,N_4861);
or U6725 (N_6725,N_1777,N_309);
or U6726 (N_6726,N_906,N_3781);
nor U6727 (N_6727,N_4267,N_3150);
xnor U6728 (N_6728,N_3677,N_1887);
xnor U6729 (N_6729,N_2213,N_4746);
or U6730 (N_6730,N_3452,N_1264);
or U6731 (N_6731,N_539,N_3744);
nor U6732 (N_6732,N_579,N_4502);
or U6733 (N_6733,N_303,N_2189);
nor U6734 (N_6734,N_3068,N_1454);
xnor U6735 (N_6735,N_1475,N_4938);
xnor U6736 (N_6736,N_2209,N_4407);
and U6737 (N_6737,N_3748,N_2073);
xnor U6738 (N_6738,N_2591,N_4189);
and U6739 (N_6739,N_1915,N_1909);
and U6740 (N_6740,N_1022,N_4320);
xor U6741 (N_6741,N_2546,N_3242);
nand U6742 (N_6742,N_4239,N_112);
nor U6743 (N_6743,N_3991,N_3394);
and U6744 (N_6744,N_2474,N_1229);
nand U6745 (N_6745,N_1921,N_3398);
or U6746 (N_6746,N_2657,N_1435);
and U6747 (N_6747,N_4909,N_3854);
nand U6748 (N_6748,N_3874,N_3110);
and U6749 (N_6749,N_2619,N_2822);
nor U6750 (N_6750,N_3833,N_3206);
nor U6751 (N_6751,N_1512,N_3704);
xor U6752 (N_6752,N_3358,N_1686);
nand U6753 (N_6753,N_1977,N_22);
or U6754 (N_6754,N_2370,N_2700);
and U6755 (N_6755,N_4709,N_466);
or U6756 (N_6756,N_2035,N_4501);
xor U6757 (N_6757,N_3061,N_1004);
nor U6758 (N_6758,N_1573,N_140);
nor U6759 (N_6759,N_1495,N_1255);
nor U6760 (N_6760,N_3165,N_668);
nor U6761 (N_6761,N_4386,N_308);
xnor U6762 (N_6762,N_320,N_860);
nor U6763 (N_6763,N_1554,N_1517);
nor U6764 (N_6764,N_3954,N_4775);
nand U6765 (N_6765,N_1996,N_3200);
nor U6766 (N_6766,N_2642,N_2317);
or U6767 (N_6767,N_3536,N_4649);
xor U6768 (N_6768,N_154,N_3608);
nand U6769 (N_6769,N_2926,N_1075);
and U6770 (N_6770,N_968,N_3392);
xor U6771 (N_6771,N_2089,N_1598);
nor U6772 (N_6772,N_1079,N_3264);
xnor U6773 (N_6773,N_3270,N_488);
nand U6774 (N_6774,N_372,N_3904);
nand U6775 (N_6775,N_4409,N_618);
nand U6776 (N_6776,N_1811,N_1361);
and U6777 (N_6777,N_2353,N_2820);
nand U6778 (N_6778,N_2504,N_4807);
or U6779 (N_6779,N_544,N_1856);
or U6780 (N_6780,N_2894,N_1559);
nor U6781 (N_6781,N_3420,N_2155);
nor U6782 (N_6782,N_3823,N_4228);
xor U6783 (N_6783,N_520,N_1333);
nand U6784 (N_6784,N_3289,N_1967);
nand U6785 (N_6785,N_4487,N_4716);
or U6786 (N_6786,N_1293,N_849);
xnor U6787 (N_6787,N_285,N_3863);
or U6788 (N_6788,N_1545,N_3578);
xor U6789 (N_6789,N_2076,N_2614);
nand U6790 (N_6790,N_2560,N_1739);
nand U6791 (N_6791,N_2384,N_833);
or U6792 (N_6792,N_1868,N_55);
xor U6793 (N_6793,N_304,N_4072);
and U6794 (N_6794,N_1098,N_1285);
nand U6795 (N_6795,N_1476,N_3987);
xor U6796 (N_6796,N_994,N_3922);
or U6797 (N_6797,N_2572,N_2986);
xor U6798 (N_6798,N_4553,N_4819);
nor U6799 (N_6799,N_3992,N_3765);
xnor U6800 (N_6800,N_2466,N_996);
or U6801 (N_6801,N_3370,N_2789);
or U6802 (N_6802,N_551,N_811);
nand U6803 (N_6803,N_3759,N_3699);
or U6804 (N_6804,N_1107,N_2141);
nor U6805 (N_6805,N_4700,N_3803);
or U6806 (N_6806,N_1307,N_836);
or U6807 (N_6807,N_766,N_1338);
nor U6808 (N_6808,N_1735,N_1633);
nand U6809 (N_6809,N_4712,N_2690);
or U6810 (N_6810,N_436,N_2183);
and U6811 (N_6811,N_408,N_4941);
nand U6812 (N_6812,N_2610,N_185);
and U6813 (N_6813,N_3799,N_446);
nand U6814 (N_6814,N_1702,N_4265);
nor U6815 (N_6815,N_1639,N_1241);
nand U6816 (N_6816,N_2393,N_1195);
nor U6817 (N_6817,N_1580,N_3139);
or U6818 (N_6818,N_799,N_1437);
nor U6819 (N_6819,N_2008,N_463);
and U6820 (N_6820,N_4375,N_4331);
and U6821 (N_6821,N_789,N_457);
and U6822 (N_6822,N_4817,N_4678);
xor U6823 (N_6823,N_3313,N_2975);
nor U6824 (N_6824,N_12,N_2265);
nor U6825 (N_6825,N_606,N_3011);
and U6826 (N_6826,N_1606,N_4106);
xnor U6827 (N_6827,N_1057,N_4598);
or U6828 (N_6828,N_4613,N_3426);
nand U6829 (N_6829,N_1930,N_2100);
xor U6830 (N_6830,N_1890,N_3623);
nor U6831 (N_6831,N_822,N_815);
or U6832 (N_6832,N_1854,N_1300);
nand U6833 (N_6833,N_4463,N_3399);
and U6834 (N_6834,N_3191,N_1239);
and U6835 (N_6835,N_1680,N_4188);
xor U6836 (N_6836,N_389,N_3615);
or U6837 (N_6837,N_354,N_3990);
nand U6838 (N_6838,N_3481,N_2032);
nand U6839 (N_6839,N_1248,N_602);
nand U6840 (N_6840,N_3963,N_2052);
nor U6841 (N_6841,N_2447,N_3190);
nor U6842 (N_6842,N_4127,N_2443);
or U6843 (N_6843,N_220,N_1781);
nor U6844 (N_6844,N_2380,N_1366);
xnor U6845 (N_6845,N_846,N_664);
nor U6846 (N_6846,N_733,N_3824);
and U6847 (N_6847,N_3318,N_63);
and U6848 (N_6848,N_4280,N_2930);
nor U6849 (N_6849,N_4391,N_4028);
nand U6850 (N_6850,N_4406,N_4816);
and U6851 (N_6851,N_2244,N_4158);
nand U6852 (N_6852,N_653,N_212);
and U6853 (N_6853,N_3116,N_357);
nand U6854 (N_6854,N_923,N_4944);
xor U6855 (N_6855,N_1674,N_1859);
nor U6856 (N_6856,N_2782,N_4966);
xnor U6857 (N_6857,N_1706,N_535);
and U6858 (N_6858,N_4361,N_704);
nor U6859 (N_6859,N_1808,N_2603);
nor U6860 (N_6860,N_999,N_4568);
nand U6861 (N_6861,N_3869,N_263);
or U6862 (N_6862,N_291,N_824);
or U6863 (N_6863,N_1577,N_1007);
and U6864 (N_6864,N_3551,N_4153);
nand U6865 (N_6865,N_3518,N_2020);
nand U6866 (N_6866,N_775,N_1210);
nor U6867 (N_6867,N_1885,N_4570);
nor U6868 (N_6868,N_1062,N_1511);
nor U6869 (N_6869,N_4503,N_987);
and U6870 (N_6870,N_757,N_278);
nand U6871 (N_6871,N_2224,N_1948);
nand U6872 (N_6872,N_948,N_4765);
or U6873 (N_6873,N_1016,N_2030);
nor U6874 (N_6874,N_1892,N_1607);
nand U6875 (N_6875,N_718,N_2906);
xnor U6876 (N_6876,N_3486,N_282);
and U6877 (N_6877,N_2044,N_2643);
xnor U6878 (N_6878,N_3650,N_2977);
nand U6879 (N_6879,N_2637,N_4820);
and U6880 (N_6880,N_3613,N_2309);
or U6881 (N_6881,N_2497,N_4643);
xnor U6882 (N_6882,N_3440,N_1737);
or U6883 (N_6883,N_3411,N_1358);
nand U6884 (N_6884,N_4054,N_3305);
xnor U6885 (N_6885,N_2070,N_620);
nand U6886 (N_6886,N_4730,N_1778);
and U6887 (N_6887,N_3131,N_2520);
xnor U6888 (N_6888,N_2290,N_404);
nand U6889 (N_6889,N_2513,N_1312);
nor U6890 (N_6890,N_584,N_3263);
and U6891 (N_6891,N_4557,N_4960);
or U6892 (N_6892,N_3542,N_2134);
and U6893 (N_6893,N_4175,N_2627);
nor U6894 (N_6894,N_3161,N_919);
and U6895 (N_6895,N_2328,N_4623);
and U6896 (N_6896,N_2361,N_1672);
xnor U6897 (N_6897,N_223,N_2268);
nor U6898 (N_6898,N_274,N_3047);
or U6899 (N_6899,N_3494,N_4852);
nand U6900 (N_6900,N_3718,N_3044);
or U6901 (N_6901,N_1823,N_3866);
nand U6902 (N_6902,N_4142,N_1124);
nor U6903 (N_6903,N_4677,N_891);
xnor U6904 (N_6904,N_2167,N_1212);
xor U6905 (N_6905,N_1839,N_3403);
and U6906 (N_6906,N_3381,N_4642);
or U6907 (N_6907,N_3199,N_2315);
nor U6908 (N_6908,N_4665,N_3281);
nand U6909 (N_6909,N_1945,N_441);
or U6910 (N_6910,N_2992,N_3884);
and U6911 (N_6911,N_904,N_3290);
xnor U6912 (N_6912,N_2281,N_3373);
or U6913 (N_6913,N_3882,N_4241);
nor U6914 (N_6914,N_737,N_687);
and U6915 (N_6915,N_3266,N_34);
nand U6916 (N_6916,N_2391,N_1665);
and U6917 (N_6917,N_641,N_3314);
xnor U6918 (N_6918,N_3905,N_2318);
and U6919 (N_6919,N_4833,N_1941);
nor U6920 (N_6920,N_3505,N_1914);
or U6921 (N_6921,N_4290,N_4931);
xor U6922 (N_6922,N_827,N_3959);
or U6923 (N_6923,N_4362,N_2676);
xnor U6924 (N_6924,N_1250,N_2786);
nand U6925 (N_6925,N_2187,N_2968);
xor U6926 (N_6926,N_98,N_4061);
xor U6927 (N_6927,N_366,N_3794);
xor U6928 (N_6928,N_985,N_289);
nor U6929 (N_6929,N_1643,N_2514);
and U6930 (N_6930,N_4969,N_1283);
or U6931 (N_6931,N_2273,N_4766);
and U6932 (N_6932,N_3947,N_2471);
xnor U6933 (N_6933,N_338,N_3883);
or U6934 (N_6934,N_2732,N_823);
and U6935 (N_6935,N_1037,N_2294);
nor U6936 (N_6936,N_2491,N_251);
and U6937 (N_6937,N_3785,N_1055);
and U6938 (N_6938,N_4904,N_4951);
nand U6939 (N_6939,N_4317,N_3970);
xor U6940 (N_6940,N_4139,N_3100);
nand U6941 (N_6941,N_850,N_4425);
nor U6942 (N_6942,N_4462,N_2951);
nor U6943 (N_6943,N_2807,N_951);
xor U6944 (N_6944,N_1741,N_2174);
or U6945 (N_6945,N_898,N_2231);
or U6946 (N_6946,N_1219,N_1806);
or U6947 (N_6947,N_2606,N_2666);
and U6948 (N_6948,N_1765,N_4604);
or U6949 (N_6949,N_2802,N_4660);
nor U6950 (N_6950,N_692,N_3114);
and U6951 (N_6951,N_3128,N_755);
nand U6952 (N_6952,N_1840,N_2214);
or U6953 (N_6953,N_4597,N_4176);
nor U6954 (N_6954,N_1128,N_2831);
and U6955 (N_6955,N_2151,N_2);
and U6956 (N_6956,N_4300,N_1886);
xnor U6957 (N_6957,N_3612,N_1701);
and U6958 (N_6958,N_4744,N_355);
or U6959 (N_6959,N_1122,N_4687);
or U6960 (N_6960,N_1988,N_717);
nand U6961 (N_6961,N_94,N_1296);
xor U6962 (N_6962,N_1773,N_1160);
xor U6963 (N_6963,N_1356,N_4291);
xnor U6964 (N_6964,N_853,N_3383);
or U6965 (N_6965,N_878,N_554);
and U6966 (N_6966,N_798,N_4269);
nand U6967 (N_6967,N_4415,N_1335);
xor U6968 (N_6968,N_788,N_1552);
xnor U6969 (N_6969,N_1183,N_2300);
nor U6970 (N_6970,N_377,N_3526);
nand U6971 (N_6971,N_2140,N_965);
xnor U6972 (N_6972,N_3337,N_2880);
or U6973 (N_6973,N_2745,N_3472);
or U6974 (N_6974,N_3731,N_3553);
nand U6975 (N_6975,N_1971,N_1937);
xnor U6976 (N_6976,N_2641,N_3603);
nor U6977 (N_6977,N_2313,N_4589);
or U6978 (N_6978,N_4494,N_4968);
and U6979 (N_6979,N_1308,N_1045);
and U6980 (N_6980,N_3369,N_81);
nand U6981 (N_6981,N_1287,N_959);
nor U6982 (N_6982,N_3845,N_214);
nor U6983 (N_6983,N_24,N_1156);
or U6984 (N_6984,N_812,N_2535);
nand U6985 (N_6985,N_3323,N_56);
and U6986 (N_6986,N_4950,N_3647);
nand U6987 (N_6987,N_411,N_299);
or U6988 (N_6988,N_2583,N_1017);
or U6989 (N_6989,N_1196,N_3216);
or U6990 (N_6990,N_3204,N_3185);
or U6991 (N_6991,N_3582,N_1786);
and U6992 (N_6992,N_1946,N_1968);
and U6993 (N_6993,N_4530,N_4620);
nor U6994 (N_6994,N_173,N_2568);
and U6995 (N_6995,N_2165,N_1506);
xnor U6996 (N_6996,N_1421,N_4299);
nor U6997 (N_6997,N_36,N_229);
nand U6998 (N_6998,N_3372,N_4509);
xor U6999 (N_6999,N_2092,N_3973);
nor U7000 (N_7000,N_3241,N_2492);
xnor U7001 (N_7001,N_1194,N_1023);
nor U7002 (N_7002,N_1998,N_233);
nand U7003 (N_7003,N_3804,N_2727);
and U7004 (N_7004,N_1198,N_64);
or U7005 (N_7005,N_2556,N_4574);
or U7006 (N_7006,N_4705,N_2834);
or U7007 (N_7007,N_970,N_4879);
xor U7008 (N_7008,N_74,N_4857);
and U7009 (N_7009,N_771,N_4859);
nand U7010 (N_7010,N_1916,N_3112);
and U7011 (N_7011,N_529,N_1997);
or U7012 (N_7012,N_1328,N_4250);
xnor U7013 (N_7013,N_4607,N_4159);
or U7014 (N_7014,N_2150,N_1234);
nand U7015 (N_7015,N_3063,N_1325);
xnor U7016 (N_7016,N_301,N_2581);
nand U7017 (N_7017,N_2109,N_3102);
xnor U7018 (N_7018,N_298,N_1934);
nand U7019 (N_7019,N_3566,N_3707);
xor U7020 (N_7020,N_1501,N_2168);
nand U7021 (N_7021,N_2617,N_888);
or U7022 (N_7022,N_135,N_4485);
xnor U7023 (N_7023,N_4948,N_66);
xnor U7024 (N_7024,N_2597,N_2283);
nor U7025 (N_7025,N_3583,N_4762);
nand U7026 (N_7026,N_2972,N_365);
xor U7027 (N_7027,N_4721,N_4843);
xnor U7028 (N_7028,N_4899,N_4540);
nand U7029 (N_7029,N_3326,N_864);
or U7030 (N_7030,N_549,N_1065);
or U7031 (N_7031,N_352,N_2026);
nand U7032 (N_7032,N_3840,N_787);
xnor U7033 (N_7033,N_2364,N_3663);
and U7034 (N_7034,N_3917,N_3858);
or U7035 (N_7035,N_3645,N_1440);
or U7036 (N_7036,N_4296,N_3674);
and U7037 (N_7037,N_4667,N_2719);
nor U7038 (N_7038,N_713,N_1368);
nor U7039 (N_7039,N_84,N_1223);
xor U7040 (N_7040,N_3238,N_1096);
nand U7041 (N_7041,N_3130,N_1907);
and U7042 (N_7042,N_1832,N_1403);
nor U7043 (N_7043,N_2811,N_1258);
and U7044 (N_7044,N_328,N_1414);
nor U7045 (N_7045,N_4090,N_2778);
or U7046 (N_7046,N_2829,N_481);
nand U7047 (N_7047,N_1152,N_3385);
nand U7048 (N_7048,N_1012,N_3651);
or U7049 (N_7049,N_4363,N_3428);
or U7050 (N_7050,N_1372,N_4392);
nor U7051 (N_7051,N_2382,N_4519);
or U7052 (N_7052,N_954,N_128);
and U7053 (N_7053,N_3937,N_3941);
and U7054 (N_7054,N_553,N_1211);
nand U7055 (N_7055,N_1095,N_2398);
nor U7056 (N_7056,N_2126,N_1789);
nand U7057 (N_7057,N_3559,N_2877);
or U7058 (N_7058,N_1138,N_4679);
and U7059 (N_7059,N_174,N_991);
xnor U7060 (N_7060,N_4010,N_4632);
or U7061 (N_7061,N_543,N_2605);
and U7062 (N_7062,N_4975,N_794);
nor U7063 (N_7063,N_2899,N_3676);
or U7064 (N_7064,N_486,N_3356);
nor U7065 (N_7065,N_672,N_4629);
nand U7066 (N_7066,N_1436,N_2449);
and U7067 (N_7067,N_1451,N_2762);
nand U7068 (N_7068,N_4137,N_1493);
nand U7069 (N_7069,N_1261,N_2530);
or U7070 (N_7070,N_4650,N_4797);
nand U7071 (N_7071,N_4830,N_4722);
nor U7072 (N_7072,N_2127,N_2145);
xor U7073 (N_7073,N_2475,N_2285);
nand U7074 (N_7074,N_3084,N_1202);
nor U7075 (N_7075,N_384,N_2847);
nand U7076 (N_7076,N_2821,N_4012);
nor U7077 (N_7077,N_1795,N_91);
nand U7078 (N_7078,N_3360,N_1176);
nand U7079 (N_7079,N_1477,N_3343);
nand U7080 (N_7080,N_2302,N_255);
nor U7081 (N_7081,N_3201,N_2699);
nand U7082 (N_7082,N_163,N_205);
nor U7083 (N_7083,N_2959,N_1625);
and U7084 (N_7084,N_3598,N_944);
and U7085 (N_7085,N_3777,N_3469);
or U7086 (N_7086,N_4018,N_2818);
and U7087 (N_7087,N_25,N_1208);
xnor U7088 (N_7088,N_3753,N_1197);
xnor U7089 (N_7089,N_2121,N_2534);
and U7090 (N_7090,N_4654,N_696);
nor U7091 (N_7091,N_600,N_4963);
nor U7092 (N_7092,N_2245,N_738);
nand U7093 (N_7093,N_2649,N_1089);
nor U7094 (N_7094,N_2289,N_2698);
or U7095 (N_7095,N_4520,N_1620);
and U7096 (N_7096,N_4610,N_1943);
xnor U7097 (N_7097,N_3771,N_472);
nand U7098 (N_7098,N_889,N_4433);
nor U7099 (N_7099,N_3953,N_2162);
nand U7100 (N_7100,N_4592,N_4671);
xor U7101 (N_7101,N_2061,N_2333);
xor U7102 (N_7102,N_2431,N_1768);
xor U7103 (N_7103,N_2681,N_65);
xnor U7104 (N_7104,N_4445,N_3457);
or U7105 (N_7105,N_1679,N_178);
xor U7106 (N_7106,N_886,N_4713);
nand U7107 (N_7107,N_1623,N_913);
and U7108 (N_7108,N_1049,N_294);
nor U7109 (N_7109,N_502,N_1965);
xnor U7110 (N_7110,N_768,N_199);
or U7111 (N_7111,N_396,N_3586);
and U7112 (N_7112,N_1226,N_85);
or U7113 (N_7113,N_2859,N_3261);
nor U7114 (N_7114,N_1919,N_1637);
xor U7115 (N_7115,N_1262,N_1146);
nand U7116 (N_7116,N_4101,N_2016);
and U7117 (N_7117,N_2031,N_1657);
xor U7118 (N_7118,N_4848,N_353);
and U7119 (N_7119,N_283,N_2893);
nor U7120 (N_7120,N_137,N_3756);
nand U7121 (N_7121,N_4977,N_4514);
and U7122 (N_7122,N_363,N_1078);
nor U7123 (N_7123,N_243,N_2383);
and U7124 (N_7124,N_3346,N_634);
or U7125 (N_7125,N_4842,N_2994);
nand U7126 (N_7126,N_2254,N_1340);
and U7127 (N_7127,N_3253,N_330);
nand U7128 (N_7128,N_1876,N_3374);
or U7129 (N_7129,N_3880,N_2435);
and U7130 (N_7130,N_2083,N_4128);
nor U7131 (N_7131,N_3187,N_2509);
nor U7132 (N_7132,N_669,N_414);
nor U7133 (N_7133,N_4197,N_1732);
nor U7134 (N_7134,N_4493,N_3257);
or U7135 (N_7135,N_1114,N_3630);
xor U7136 (N_7136,N_3920,N_3401);
and U7137 (N_7137,N_1401,N_825);
and U7138 (N_7138,N_2378,N_1974);
and U7139 (N_7139,N_2270,N_2790);
or U7140 (N_7140,N_2476,N_4323);
or U7141 (N_7141,N_490,N_2754);
xnor U7142 (N_7142,N_3761,N_1265);
nor U7143 (N_7143,N_3227,N_728);
xnor U7144 (N_7144,N_4103,N_1985);
or U7145 (N_7145,N_17,N_3528);
nor U7146 (N_7146,N_1972,N_2757);
xnor U7147 (N_7147,N_614,N_2157);
nand U7148 (N_7148,N_1754,N_1409);
or U7149 (N_7149,N_740,N_4480);
xnor U7150 (N_7150,N_4921,N_4144);
and U7151 (N_7151,N_2923,N_235);
xnor U7152 (N_7152,N_1583,N_4808);
or U7153 (N_7153,N_2902,N_3259);
and U7154 (N_7154,N_3509,N_2013);
nor U7155 (N_7155,N_1420,N_4841);
nand U7156 (N_7156,N_4282,N_149);
xnor U7157 (N_7157,N_2107,N_2759);
or U7158 (N_7158,N_4432,N_885);
or U7159 (N_7159,N_358,N_4851);
nor U7160 (N_7160,N_2113,N_4283);
and U7161 (N_7161,N_2804,N_2952);
xor U7162 (N_7162,N_4786,N_464);
nand U7163 (N_7163,N_1144,N_2708);
nor U7164 (N_7164,N_1093,N_3171);
or U7165 (N_7165,N_3806,N_1931);
xor U7166 (N_7166,N_3749,N_2143);
xor U7167 (N_7167,N_3108,N_30);
or U7168 (N_7168,N_2979,N_2346);
and U7169 (N_7169,N_3737,N_980);
nand U7170 (N_7170,N_4422,N_1812);
or U7171 (N_7171,N_1105,N_2989);
nand U7172 (N_7172,N_1484,N_3006);
xor U7173 (N_7173,N_3004,N_4639);
nand U7174 (N_7174,N_3852,N_2437);
xor U7175 (N_7175,N_2009,N_1889);
or U7176 (N_7176,N_2484,N_3194);
and U7177 (N_7177,N_3855,N_977);
or U7178 (N_7178,N_1375,N_2695);
nor U7179 (N_7179,N_2368,N_4325);
and U7180 (N_7180,N_3545,N_4200);
nand U7181 (N_7181,N_3251,N_1281);
xnor U7182 (N_7182,N_1681,N_3106);
and U7183 (N_7183,N_3126,N_1465);
nor U7184 (N_7184,N_750,N_2541);
xor U7185 (N_7185,N_3432,N_4945);
or U7186 (N_7186,N_3075,N_3783);
nor U7187 (N_7187,N_4549,N_4149);
xor U7188 (N_7188,N_2741,N_1579);
or U7189 (N_7189,N_3982,N_3571);
and U7190 (N_7190,N_3341,N_86);
nor U7191 (N_7191,N_1550,N_428);
xnor U7192 (N_7192,N_2024,N_2354);
nand U7193 (N_7193,N_119,N_4225);
or U7194 (N_7194,N_3763,N_1508);
nand U7195 (N_7195,N_241,N_4624);
and U7196 (N_7196,N_171,N_1083);
nand U7197 (N_7197,N_2228,N_300);
or U7198 (N_7198,N_3989,N_893);
nor U7199 (N_7199,N_4971,N_773);
nor U7200 (N_7200,N_3308,N_151);
xnor U7201 (N_7201,N_4346,N_4027);
or U7202 (N_7202,N_1846,N_1488);
and U7203 (N_7203,N_2438,N_3924);
or U7204 (N_7204,N_3462,N_2948);
nand U7205 (N_7205,N_2803,N_1060);
and U7206 (N_7206,N_610,N_552);
nand U7207 (N_7207,N_3857,N_1984);
or U7208 (N_7208,N_3808,N_1254);
nor U7209 (N_7209,N_1150,N_1918);
or U7210 (N_7210,N_756,N_1278);
nor U7211 (N_7211,N_270,N_3802);
xor U7212 (N_7212,N_3415,N_4886);
nand U7213 (N_7213,N_348,N_3885);
nand U7214 (N_7214,N_141,N_4983);
or U7215 (N_7215,N_2472,N_1350);
and U7216 (N_7216,N_2075,N_4243);
nand U7217 (N_7217,N_4834,N_896);
xnor U7218 (N_7218,N_4111,N_3898);
nor U7219 (N_7219,N_3178,N_1582);
nor U7220 (N_7220,N_2624,N_2939);
and U7221 (N_7221,N_1169,N_1537);
xnor U7222 (N_7222,N_3239,N_1020);
nor U7223 (N_7223,N_4203,N_4518);
nand U7224 (N_7224,N_4732,N_3870);
or U7225 (N_7225,N_1189,N_818);
xnor U7226 (N_7226,N_1301,N_2152);
nand U7227 (N_7227,N_1588,N_3530);
xnor U7228 (N_7228,N_3695,N_3910);
or U7229 (N_7229,N_1802,N_1857);
or U7230 (N_7230,N_1541,N_2006);
nand U7231 (N_7231,N_4959,N_4657);
and U7232 (N_7232,N_1446,N_4694);
or U7233 (N_7233,N_4758,N_447);
xnor U7234 (N_7234,N_3340,N_1575);
or U7235 (N_7235,N_3789,N_4002);
xnor U7236 (N_7236,N_1031,N_1054);
or U7237 (N_7237,N_2917,N_1438);
xor U7238 (N_7238,N_2907,N_3182);
nor U7239 (N_7239,N_1962,N_3339);
nor U7240 (N_7240,N_4894,N_596);
xor U7241 (N_7241,N_3085,N_1297);
and U7242 (N_7242,N_3648,N_3352);
and U7243 (N_7243,N_3964,N_938);
or U7244 (N_7244,N_4625,N_1180);
nor U7245 (N_7245,N_2199,N_995);
nor U7246 (N_7246,N_2839,N_3693);
and U7247 (N_7247,N_4437,N_1630);
and U7248 (N_7248,N_2195,N_4739);
nor U7249 (N_7249,N_2726,N_2956);
or U7250 (N_7250,N_1270,N_3502);
nor U7251 (N_7251,N_1452,N_3549);
xor U7252 (N_7252,N_870,N_3776);
and U7253 (N_7253,N_461,N_2658);
xor U7254 (N_7254,N_2661,N_1391);
xor U7255 (N_7255,N_1616,N_498);
nand U7256 (N_7256,N_3404,N_548);
nand U7257 (N_7257,N_1290,N_3382);
nand U7258 (N_7258,N_1661,N_4872);
nor U7259 (N_7259,N_362,N_2427);
nand U7260 (N_7260,N_4063,N_2095);
and U7261 (N_7261,N_4161,N_297);
and U7262 (N_7262,N_1348,N_4982);
or U7263 (N_7263,N_630,N_1612);
xnor U7264 (N_7264,N_2733,N_4360);
and U7265 (N_7265,N_4408,N_4148);
nor U7266 (N_7266,N_1820,N_800);
and U7267 (N_7267,N_1349,N_3519);
or U7268 (N_7268,N_2738,N_1121);
nor U7269 (N_7269,N_3682,N_841);
xnor U7270 (N_7270,N_492,N_4784);
nand U7271 (N_7271,N_621,N_884);
xnor U7272 (N_7272,N_4900,N_2607);
nand U7273 (N_7273,N_2238,N_469);
or U7274 (N_7274,N_3087,N_3397);
or U7275 (N_7275,N_2442,N_115);
or U7276 (N_7276,N_40,N_3491);
nor U7277 (N_7277,N_3609,N_2081);
and U7278 (N_7278,N_3181,N_3345);
or U7279 (N_7279,N_3592,N_2842);
or U7280 (N_7280,N_143,N_4000);
xor U7281 (N_7281,N_3554,N_2815);
xnor U7282 (N_7282,N_1544,N_4618);
or U7283 (N_7283,N_2170,N_4081);
or U7284 (N_7284,N_2343,N_3587);
nor U7285 (N_7285,N_2067,N_479);
nand U7286 (N_7286,N_1374,N_2653);
xnor U7287 (N_7287,N_1310,N_3429);
or U7288 (N_7288,N_4866,N_3900);
and U7289 (N_7289,N_3170,N_3733);
and U7290 (N_7290,N_3712,N_4129);
xor U7291 (N_7291,N_873,N_4330);
nand U7292 (N_7292,N_2090,N_1473);
nand U7293 (N_7293,N_4777,N_248);
nand U7294 (N_7294,N_3594,N_711);
or U7295 (N_7295,N_2964,N_1956);
or U7296 (N_7296,N_3543,N_3848);
and U7297 (N_7297,N_421,N_4186);
and U7298 (N_7298,N_3280,N_2413);
nand U7299 (N_7299,N_200,N_4198);
nor U7300 (N_7300,N_4871,N_1990);
or U7301 (N_7301,N_1220,N_3563);
and U7302 (N_7302,N_1539,N_165);
nand U7303 (N_7303,N_234,N_922);
or U7304 (N_7304,N_730,N_3668);
nor U7305 (N_7305,N_4752,N_578);
nor U7306 (N_7306,N_1784,N_2640);
nand U7307 (N_7307,N_4537,N_1458);
nor U7308 (N_7308,N_3817,N_3081);
or U7309 (N_7309,N_3303,N_1610);
nand U7310 (N_7310,N_2686,N_1531);
nand U7311 (N_7311,N_4910,N_1969);
and U7312 (N_7312,N_1154,N_2404);
or U7313 (N_7313,N_4321,N_3071);
or U7314 (N_7314,N_1309,N_1430);
nor U7315 (N_7315,N_4508,N_194);
xnor U7316 (N_7316,N_3787,N_193);
or U7317 (N_7317,N_4828,N_817);
and U7318 (N_7318,N_691,N_1321);
and U7319 (N_7319,N_2769,N_1046);
nor U7320 (N_7320,N_892,N_4345);
nor U7321 (N_7321,N_177,N_1304);
and U7322 (N_7322,N_4428,N_3315);
xor U7323 (N_7323,N_2392,N_2780);
xor U7324 (N_7324,N_3049,N_4171);
nor U7325 (N_7325,N_3010,N_4506);
xnor U7326 (N_7326,N_167,N_3736);
nor U7327 (N_7327,N_2833,N_3875);
xor U7328 (N_7328,N_2913,N_2445);
xor U7329 (N_7329,N_478,N_2416);
nor U7330 (N_7330,N_1182,N_2206);
and U7331 (N_7331,N_3945,N_4477);
or U7332 (N_7332,N_3681,N_2412);
and U7333 (N_7333,N_4235,N_1111);
nor U7334 (N_7334,N_2945,N_2365);
or U7335 (N_7335,N_306,N_2722);
xor U7336 (N_7336,N_526,N_4019);
and U7337 (N_7337,N_871,N_3983);
nand U7338 (N_7338,N_4918,N_1385);
or U7339 (N_7339,N_1753,N_1949);
and U7340 (N_7340,N_3124,N_2017);
xor U7341 (N_7341,N_2160,N_2801);
and U7342 (N_7342,N_4263,N_2683);
and U7343 (N_7343,N_4707,N_1149);
nor U7344 (N_7344,N_3176,N_224);
nand U7345 (N_7345,N_4780,N_3053);
nor U7346 (N_7346,N_2792,N_1390);
or U7347 (N_7347,N_657,N_343);
nand U7348 (N_7348,N_1485,N_3474);
xnor U7349 (N_7349,N_615,N_1097);
xnor U7350 (N_7350,N_1712,N_2124);
and U7351 (N_7351,N_1751,N_4049);
or U7352 (N_7352,N_4805,N_3412);
nor U7353 (N_7353,N_4799,N_982);
or U7354 (N_7354,N_3807,N_3952);
and U7355 (N_7355,N_4726,N_4085);
nand U7356 (N_7356,N_4163,N_148);
xnor U7357 (N_7357,N_4482,N_2482);
or U7358 (N_7358,N_4187,N_1110);
nand U7359 (N_7359,N_496,N_2261);
nor U7360 (N_7360,N_936,N_3232);
xor U7361 (N_7361,N_3142,N_364);
xnor U7362 (N_7362,N_431,N_2336);
xor U7363 (N_7363,N_4562,N_1441);
nor U7364 (N_7364,N_3641,N_450);
nor U7365 (N_7365,N_2855,N_993);
and U7366 (N_7366,N_3325,N_4209);
nor U7367 (N_7367,N_3517,N_2874);
nor U7368 (N_7368,N_3721,N_4725);
nand U7369 (N_7369,N_3002,N_3984);
and U7370 (N_7370,N_2169,N_2753);
nand U7371 (N_7371,N_1750,N_1243);
or U7372 (N_7372,N_2836,N_628);
and U7373 (N_7373,N_2920,N_4358);
nor U7374 (N_7374,N_3899,N_3865);
and U7375 (N_7375,N_3167,N_834);
nor U7376 (N_7376,N_4095,N_2984);
nand U7377 (N_7377,N_1491,N_3544);
or U7378 (N_7378,N_1367,N_1139);
nor U7379 (N_7379,N_577,N_1313);
xnor U7380 (N_7380,N_225,N_1871);
xor U7381 (N_7381,N_899,N_4958);
xor U7382 (N_7382,N_1710,N_4057);
xor U7383 (N_7383,N_4708,N_3558);
and U7384 (N_7384,N_1752,N_1792);
nor U7385 (N_7385,N_2314,N_2355);
nor U7386 (N_7386,N_3907,N_2594);
nor U7387 (N_7387,N_613,N_4575);
and U7388 (N_7388,N_3174,N_4787);
and U7389 (N_7389,N_844,N_1809);
and U7390 (N_7390,N_797,N_777);
xor U7391 (N_7391,N_4964,N_1217);
nor U7392 (N_7392,N_3003,N_2312);
xnor U7393 (N_7393,N_448,N_4988);
and U7394 (N_7394,N_587,N_4079);
nand U7395 (N_7395,N_3471,N_1851);
or U7396 (N_7396,N_1378,N_4978);
and U7397 (N_7397,N_1380,N_1502);
nor U7398 (N_7398,N_101,N_2558);
nand U7399 (N_7399,N_1875,N_4511);
nand U7400 (N_7400,N_4374,N_2908);
and U7401 (N_7401,N_3055,N_1816);
and U7402 (N_7402,N_3838,N_4827);
and U7403 (N_7403,N_4182,N_883);
nand U7404 (N_7404,N_2163,N_4507);
and U7405 (N_7405,N_345,N_2465);
and U7406 (N_7406,N_4220,N_2883);
xnor U7407 (N_7407,N_4548,N_848);
or U7408 (N_7408,N_3453,N_3741);
or U7409 (N_7409,N_2373,N_1744);
nor U7410 (N_7410,N_375,N_4663);
xor U7411 (N_7411,N_394,N_2461);
or U7412 (N_7412,N_2903,N_796);
and U7413 (N_7413,N_2128,N_4037);
nand U7414 (N_7414,N_645,N_2340);
nor U7415 (N_7415,N_311,N_4617);
xnor U7416 (N_7416,N_1039,N_77);
xor U7417 (N_7417,N_2549,N_1950);
nand U7418 (N_7418,N_1862,N_3054);
nand U7419 (N_7419,N_1624,N_3272);
or U7420 (N_7420,N_1858,N_1547);
and U7421 (N_7421,N_4001,N_828);
nand U7422 (N_7422,N_2625,N_3331);
or U7423 (N_7423,N_2892,N_4275);
xor U7424 (N_7424,N_16,N_2423);
and U7425 (N_7425,N_13,N_4051);
or U7426 (N_7426,N_565,N_1433);
nand U7427 (N_7427,N_1691,N_3222);
or U7428 (N_7428,N_4822,N_723);
and U7429 (N_7429,N_4609,N_3473);
or U7430 (N_7430,N_1603,N_237);
nor U7431 (N_7431,N_2882,N_2041);
xor U7432 (N_7432,N_4318,N_4369);
xor U7433 (N_7433,N_80,N_4965);
or U7434 (N_7434,N_3048,N_3565);
nand U7435 (N_7435,N_1227,N_1824);
nand U7436 (N_7436,N_3909,N_2810);
and U7437 (N_7437,N_4440,N_523);
xnor U7438 (N_7438,N_1125,N_2854);
nand U7439 (N_7439,N_916,N_460);
and U7440 (N_7440,N_1145,N_1940);
nand U7441 (N_7441,N_1462,N_322);
or U7442 (N_7442,N_869,N_3786);
xnor U7443 (N_7443,N_1651,N_1221);
nor U7444 (N_7444,N_4767,N_3319);
nor U7445 (N_7445,N_4875,N_3237);
and U7446 (N_7446,N_2598,N_4058);
nand U7447 (N_7447,N_2185,N_671);
or U7448 (N_7448,N_1047,N_1747);
and U7449 (N_7449,N_4284,N_3971);
nor U7450 (N_7450,N_3386,N_4491);
and U7451 (N_7451,N_2749,N_1044);
or U7452 (N_7452,N_2078,N_746);
nor U7453 (N_7453,N_4388,N_1439);
nand U7454 (N_7454,N_4138,N_3988);
nand U7455 (N_7455,N_4551,N_3931);
nor U7456 (N_7456,N_3138,N_4356);
nor U7457 (N_7457,N_4075,N_1704);
xnor U7458 (N_7458,N_4196,N_2856);
and U7459 (N_7459,N_1818,N_2587);
or U7460 (N_7460,N_2144,N_3159);
or U7461 (N_7461,N_3734,N_221);
nor U7462 (N_7462,N_950,N_4316);
or U7463 (N_7463,N_2415,N_2943);
nor U7464 (N_7464,N_3443,N_1727);
nor U7465 (N_7465,N_858,N_1912);
xor U7466 (N_7466,N_1827,N_1053);
nor U7467 (N_7467,N_1126,N_3498);
and U7468 (N_7468,N_1535,N_2567);
nand U7469 (N_7469,N_4264,N_4444);
nor U7470 (N_7470,N_1157,N_2748);
nand U7471 (N_7471,N_654,N_2010);
nor U7472 (N_7472,N_3640,N_1622);
or U7473 (N_7473,N_4932,N_203);
nor U7474 (N_7474,N_392,N_4603);
and U7475 (N_7475,N_2087,N_1175);
or U7476 (N_7476,N_3956,N_1445);
nand U7477 (N_7477,N_7,N_3465);
or U7478 (N_7478,N_2777,N_2799);
and U7479 (N_7479,N_2997,N_2868);
nor U7480 (N_7480,N_272,N_1362);
xor U7481 (N_7481,N_1635,N_4466);
nor U7482 (N_7482,N_2115,N_1671);
nand U7483 (N_7483,N_2220,N_1400);
xnor U7484 (N_7484,N_27,N_4588);
nor U7485 (N_7485,N_1256,N_1713);
nand U7486 (N_7486,N_4661,N_72);
nand U7487 (N_7487,N_1048,N_1188);
nor U7488 (N_7488,N_1528,N_157);
nand U7489 (N_7489,N_4108,N_2179);
and U7490 (N_7490,N_4653,N_3557);
or U7491 (N_7491,N_2714,N_3513);
nand U7492 (N_7492,N_4231,N_2659);
xnor U7493 (N_7493,N_879,N_2532);
and U7494 (N_7494,N_1591,N_1925);
and U7495 (N_7495,N_4077,N_349);
nor U7496 (N_7496,N_2697,N_3459);
nor U7497 (N_7497,N_4347,N_79);
xnor U7498 (N_7498,N_2122,N_882);
nor U7499 (N_7499,N_4185,N_4836);
and U7500 (N_7500,N_261,N_3389);
nor U7501 (N_7501,N_3989,N_1913);
xor U7502 (N_7502,N_2053,N_2922);
or U7503 (N_7503,N_4002,N_2032);
nor U7504 (N_7504,N_4802,N_117);
nand U7505 (N_7505,N_1579,N_371);
or U7506 (N_7506,N_106,N_4845);
and U7507 (N_7507,N_3590,N_2093);
and U7508 (N_7508,N_7,N_1466);
nor U7509 (N_7509,N_776,N_3258);
or U7510 (N_7510,N_2859,N_1127);
or U7511 (N_7511,N_1446,N_1856);
xor U7512 (N_7512,N_424,N_2838);
xor U7513 (N_7513,N_817,N_4813);
nand U7514 (N_7514,N_1161,N_1547);
and U7515 (N_7515,N_397,N_1117);
xnor U7516 (N_7516,N_1433,N_4817);
xnor U7517 (N_7517,N_3459,N_574);
xnor U7518 (N_7518,N_2241,N_3220);
nor U7519 (N_7519,N_2764,N_3190);
nor U7520 (N_7520,N_948,N_1890);
or U7521 (N_7521,N_169,N_3937);
or U7522 (N_7522,N_4837,N_445);
xnor U7523 (N_7523,N_3739,N_1527);
or U7524 (N_7524,N_2744,N_1564);
or U7525 (N_7525,N_704,N_2658);
nand U7526 (N_7526,N_472,N_4631);
nand U7527 (N_7527,N_4289,N_1430);
nor U7528 (N_7528,N_2191,N_4590);
or U7529 (N_7529,N_216,N_4290);
nand U7530 (N_7530,N_760,N_4448);
nor U7531 (N_7531,N_3651,N_584);
xor U7532 (N_7532,N_1229,N_1561);
and U7533 (N_7533,N_2010,N_3534);
nor U7534 (N_7534,N_376,N_2140);
xnor U7535 (N_7535,N_4613,N_3723);
nor U7536 (N_7536,N_3912,N_1819);
or U7537 (N_7537,N_3635,N_4256);
or U7538 (N_7538,N_3628,N_3927);
xnor U7539 (N_7539,N_4261,N_3118);
nor U7540 (N_7540,N_1266,N_4778);
nand U7541 (N_7541,N_3201,N_2045);
nor U7542 (N_7542,N_67,N_4917);
nor U7543 (N_7543,N_3453,N_3143);
or U7544 (N_7544,N_3668,N_3300);
and U7545 (N_7545,N_526,N_1495);
nor U7546 (N_7546,N_2398,N_837);
nand U7547 (N_7547,N_565,N_1608);
xnor U7548 (N_7548,N_3246,N_1248);
nor U7549 (N_7549,N_718,N_2502);
or U7550 (N_7550,N_482,N_2996);
nand U7551 (N_7551,N_4332,N_2950);
nand U7552 (N_7552,N_3816,N_2116);
and U7553 (N_7553,N_3855,N_4898);
or U7554 (N_7554,N_2010,N_4874);
xor U7555 (N_7555,N_1901,N_14);
and U7556 (N_7556,N_2799,N_3620);
or U7557 (N_7557,N_983,N_2041);
xnor U7558 (N_7558,N_1229,N_1984);
or U7559 (N_7559,N_2517,N_3871);
xor U7560 (N_7560,N_4458,N_1868);
and U7561 (N_7561,N_3118,N_3064);
nor U7562 (N_7562,N_2785,N_261);
nor U7563 (N_7563,N_4809,N_2772);
nor U7564 (N_7564,N_4098,N_892);
nor U7565 (N_7565,N_4895,N_730);
xor U7566 (N_7566,N_1046,N_2377);
nand U7567 (N_7567,N_3111,N_1295);
nand U7568 (N_7568,N_3050,N_4847);
or U7569 (N_7569,N_3751,N_3920);
nor U7570 (N_7570,N_135,N_1836);
xor U7571 (N_7571,N_4671,N_4563);
and U7572 (N_7572,N_651,N_2544);
and U7573 (N_7573,N_576,N_2258);
and U7574 (N_7574,N_3918,N_3707);
and U7575 (N_7575,N_3780,N_803);
nand U7576 (N_7576,N_407,N_573);
and U7577 (N_7577,N_1072,N_981);
nor U7578 (N_7578,N_627,N_4354);
and U7579 (N_7579,N_337,N_3304);
nand U7580 (N_7580,N_1050,N_919);
xor U7581 (N_7581,N_2259,N_1298);
or U7582 (N_7582,N_2741,N_2259);
xor U7583 (N_7583,N_2161,N_796);
nand U7584 (N_7584,N_4906,N_560);
or U7585 (N_7585,N_2728,N_945);
nor U7586 (N_7586,N_4707,N_2802);
nor U7587 (N_7587,N_2982,N_1289);
nor U7588 (N_7588,N_3460,N_4902);
and U7589 (N_7589,N_3542,N_2655);
nand U7590 (N_7590,N_815,N_1949);
xor U7591 (N_7591,N_4288,N_821);
and U7592 (N_7592,N_4131,N_2437);
xor U7593 (N_7593,N_719,N_1696);
and U7594 (N_7594,N_1659,N_569);
xnor U7595 (N_7595,N_3017,N_2134);
nor U7596 (N_7596,N_1394,N_3339);
nand U7597 (N_7597,N_1993,N_716);
and U7598 (N_7598,N_752,N_459);
nor U7599 (N_7599,N_4700,N_927);
nor U7600 (N_7600,N_1240,N_3284);
and U7601 (N_7601,N_1959,N_3974);
and U7602 (N_7602,N_2084,N_3335);
nand U7603 (N_7603,N_2171,N_2551);
nor U7604 (N_7604,N_2953,N_1866);
or U7605 (N_7605,N_2866,N_1660);
nor U7606 (N_7606,N_4120,N_3800);
xnor U7607 (N_7607,N_4777,N_2703);
and U7608 (N_7608,N_2693,N_673);
nand U7609 (N_7609,N_552,N_1304);
nor U7610 (N_7610,N_4006,N_2171);
xnor U7611 (N_7611,N_2770,N_645);
and U7612 (N_7612,N_3841,N_1705);
or U7613 (N_7613,N_4515,N_1875);
and U7614 (N_7614,N_1433,N_257);
xor U7615 (N_7615,N_4085,N_4363);
nor U7616 (N_7616,N_1130,N_4619);
or U7617 (N_7617,N_124,N_1152);
nor U7618 (N_7618,N_4267,N_91);
and U7619 (N_7619,N_712,N_2851);
nor U7620 (N_7620,N_3387,N_2002);
or U7621 (N_7621,N_564,N_3193);
or U7622 (N_7622,N_4937,N_1347);
nor U7623 (N_7623,N_1757,N_4363);
xor U7624 (N_7624,N_3583,N_3443);
or U7625 (N_7625,N_2490,N_4435);
and U7626 (N_7626,N_1840,N_1076);
xor U7627 (N_7627,N_4726,N_3693);
nor U7628 (N_7628,N_3152,N_2981);
xnor U7629 (N_7629,N_4951,N_1929);
nor U7630 (N_7630,N_41,N_642);
xnor U7631 (N_7631,N_2671,N_2523);
or U7632 (N_7632,N_2627,N_929);
and U7633 (N_7633,N_2595,N_1544);
or U7634 (N_7634,N_4823,N_4896);
nand U7635 (N_7635,N_711,N_3149);
nand U7636 (N_7636,N_4173,N_4778);
xor U7637 (N_7637,N_3044,N_2900);
or U7638 (N_7638,N_4692,N_2684);
nand U7639 (N_7639,N_1252,N_3163);
or U7640 (N_7640,N_3118,N_1925);
or U7641 (N_7641,N_4080,N_320);
nand U7642 (N_7642,N_3220,N_4793);
xnor U7643 (N_7643,N_3692,N_4578);
or U7644 (N_7644,N_244,N_2718);
xor U7645 (N_7645,N_454,N_4518);
or U7646 (N_7646,N_476,N_4911);
nand U7647 (N_7647,N_3914,N_1920);
and U7648 (N_7648,N_18,N_3754);
nand U7649 (N_7649,N_3432,N_1076);
xnor U7650 (N_7650,N_4193,N_1538);
or U7651 (N_7651,N_4509,N_1358);
or U7652 (N_7652,N_2544,N_4755);
xor U7653 (N_7653,N_234,N_973);
or U7654 (N_7654,N_2268,N_776);
or U7655 (N_7655,N_3835,N_492);
nor U7656 (N_7656,N_1976,N_2527);
nor U7657 (N_7657,N_2300,N_1056);
xor U7658 (N_7658,N_378,N_913);
nor U7659 (N_7659,N_651,N_490);
nand U7660 (N_7660,N_2709,N_3622);
or U7661 (N_7661,N_4950,N_639);
nand U7662 (N_7662,N_4062,N_671);
nand U7663 (N_7663,N_3306,N_1844);
nand U7664 (N_7664,N_3935,N_850);
or U7665 (N_7665,N_144,N_1397);
nand U7666 (N_7666,N_4283,N_2054);
nand U7667 (N_7667,N_650,N_401);
or U7668 (N_7668,N_1464,N_4681);
xnor U7669 (N_7669,N_1785,N_1188);
nand U7670 (N_7670,N_1591,N_4803);
nor U7671 (N_7671,N_1169,N_3525);
nand U7672 (N_7672,N_1891,N_1048);
and U7673 (N_7673,N_2830,N_1073);
xor U7674 (N_7674,N_2785,N_2595);
nand U7675 (N_7675,N_3217,N_4985);
or U7676 (N_7676,N_3600,N_3346);
xor U7677 (N_7677,N_1909,N_42);
nor U7678 (N_7678,N_475,N_2204);
xor U7679 (N_7679,N_4959,N_4225);
nor U7680 (N_7680,N_3034,N_3374);
xor U7681 (N_7681,N_2150,N_443);
or U7682 (N_7682,N_1298,N_1048);
nand U7683 (N_7683,N_2131,N_2211);
or U7684 (N_7684,N_0,N_3625);
nand U7685 (N_7685,N_4858,N_710);
nor U7686 (N_7686,N_1870,N_2321);
and U7687 (N_7687,N_670,N_4519);
and U7688 (N_7688,N_2233,N_345);
nand U7689 (N_7689,N_2352,N_102);
nand U7690 (N_7690,N_462,N_1017);
xnor U7691 (N_7691,N_2561,N_51);
nor U7692 (N_7692,N_2294,N_2620);
nor U7693 (N_7693,N_4976,N_1644);
and U7694 (N_7694,N_4932,N_3524);
and U7695 (N_7695,N_1532,N_580);
xor U7696 (N_7696,N_4663,N_1857);
xnor U7697 (N_7697,N_3515,N_1323);
nor U7698 (N_7698,N_4223,N_3459);
or U7699 (N_7699,N_3285,N_3945);
or U7700 (N_7700,N_371,N_1564);
or U7701 (N_7701,N_63,N_2902);
nand U7702 (N_7702,N_228,N_3256);
or U7703 (N_7703,N_1574,N_226);
nor U7704 (N_7704,N_2740,N_1933);
nor U7705 (N_7705,N_2795,N_4456);
or U7706 (N_7706,N_995,N_49);
and U7707 (N_7707,N_4158,N_536);
and U7708 (N_7708,N_3111,N_1913);
and U7709 (N_7709,N_4010,N_2500);
or U7710 (N_7710,N_623,N_3140);
nor U7711 (N_7711,N_2706,N_3336);
nand U7712 (N_7712,N_4947,N_1904);
nor U7713 (N_7713,N_4153,N_1547);
nand U7714 (N_7714,N_1050,N_1727);
and U7715 (N_7715,N_4110,N_3652);
or U7716 (N_7716,N_2159,N_3686);
xnor U7717 (N_7717,N_4983,N_2043);
and U7718 (N_7718,N_1681,N_4862);
nand U7719 (N_7719,N_2346,N_4128);
and U7720 (N_7720,N_362,N_1827);
xnor U7721 (N_7721,N_3915,N_1471);
nor U7722 (N_7722,N_3377,N_2524);
nor U7723 (N_7723,N_395,N_841);
nand U7724 (N_7724,N_3125,N_4857);
or U7725 (N_7725,N_3925,N_2589);
nor U7726 (N_7726,N_605,N_160);
nand U7727 (N_7727,N_496,N_1734);
nor U7728 (N_7728,N_3269,N_2563);
nor U7729 (N_7729,N_2815,N_828);
and U7730 (N_7730,N_872,N_111);
and U7731 (N_7731,N_978,N_1174);
nand U7732 (N_7732,N_940,N_4307);
xnor U7733 (N_7733,N_4155,N_2758);
xor U7734 (N_7734,N_1885,N_4618);
or U7735 (N_7735,N_2133,N_1033);
or U7736 (N_7736,N_2854,N_1573);
xor U7737 (N_7737,N_962,N_2817);
nor U7738 (N_7738,N_4505,N_4496);
and U7739 (N_7739,N_4744,N_1442);
xor U7740 (N_7740,N_872,N_1980);
xor U7741 (N_7741,N_2279,N_2049);
nand U7742 (N_7742,N_4188,N_2657);
nand U7743 (N_7743,N_3209,N_2053);
nor U7744 (N_7744,N_271,N_4590);
nor U7745 (N_7745,N_1357,N_1741);
nand U7746 (N_7746,N_3858,N_3195);
or U7747 (N_7747,N_4333,N_4982);
and U7748 (N_7748,N_3972,N_2451);
or U7749 (N_7749,N_2484,N_4732);
nand U7750 (N_7750,N_2291,N_1274);
nand U7751 (N_7751,N_2164,N_1494);
nor U7752 (N_7752,N_3599,N_4236);
nand U7753 (N_7753,N_2694,N_710);
nand U7754 (N_7754,N_3613,N_1888);
and U7755 (N_7755,N_4251,N_4130);
nor U7756 (N_7756,N_2423,N_3338);
nand U7757 (N_7757,N_2691,N_3291);
and U7758 (N_7758,N_2172,N_2856);
nand U7759 (N_7759,N_3095,N_2871);
xor U7760 (N_7760,N_2717,N_3439);
and U7761 (N_7761,N_3267,N_3320);
xnor U7762 (N_7762,N_4350,N_731);
and U7763 (N_7763,N_4304,N_1686);
or U7764 (N_7764,N_2212,N_3618);
and U7765 (N_7765,N_2984,N_4496);
nor U7766 (N_7766,N_188,N_1667);
or U7767 (N_7767,N_1106,N_2194);
nor U7768 (N_7768,N_1938,N_2369);
and U7769 (N_7769,N_1932,N_3643);
and U7770 (N_7770,N_4593,N_411);
nor U7771 (N_7771,N_4771,N_3884);
xor U7772 (N_7772,N_429,N_170);
nand U7773 (N_7773,N_1119,N_4001);
nor U7774 (N_7774,N_1866,N_1670);
or U7775 (N_7775,N_3639,N_3042);
xor U7776 (N_7776,N_1356,N_1070);
and U7777 (N_7777,N_31,N_2204);
nand U7778 (N_7778,N_3474,N_2593);
and U7779 (N_7779,N_751,N_3200);
xnor U7780 (N_7780,N_1440,N_584);
xor U7781 (N_7781,N_3558,N_4953);
or U7782 (N_7782,N_4289,N_1336);
nor U7783 (N_7783,N_4556,N_865);
xor U7784 (N_7784,N_4308,N_3087);
or U7785 (N_7785,N_3185,N_3056);
nor U7786 (N_7786,N_4340,N_2983);
xnor U7787 (N_7787,N_3857,N_435);
and U7788 (N_7788,N_1323,N_2078);
nand U7789 (N_7789,N_2250,N_3850);
xor U7790 (N_7790,N_4398,N_2468);
nor U7791 (N_7791,N_164,N_1868);
xor U7792 (N_7792,N_1782,N_4200);
or U7793 (N_7793,N_3774,N_1539);
xnor U7794 (N_7794,N_4027,N_303);
and U7795 (N_7795,N_3233,N_3374);
or U7796 (N_7796,N_4309,N_1493);
or U7797 (N_7797,N_4918,N_3031);
and U7798 (N_7798,N_6,N_4491);
xnor U7799 (N_7799,N_1713,N_2410);
or U7800 (N_7800,N_306,N_2157);
nand U7801 (N_7801,N_1855,N_770);
nand U7802 (N_7802,N_3260,N_3686);
nor U7803 (N_7803,N_784,N_2708);
or U7804 (N_7804,N_1928,N_141);
xor U7805 (N_7805,N_722,N_312);
xor U7806 (N_7806,N_4066,N_4180);
nor U7807 (N_7807,N_3525,N_126);
or U7808 (N_7808,N_1147,N_2363);
and U7809 (N_7809,N_1013,N_1057);
or U7810 (N_7810,N_3706,N_4343);
nor U7811 (N_7811,N_2593,N_2787);
xor U7812 (N_7812,N_1497,N_2665);
and U7813 (N_7813,N_2525,N_1955);
nand U7814 (N_7814,N_1199,N_1985);
nand U7815 (N_7815,N_1914,N_4117);
xor U7816 (N_7816,N_373,N_3137);
xor U7817 (N_7817,N_743,N_1053);
and U7818 (N_7818,N_4056,N_4682);
and U7819 (N_7819,N_289,N_1346);
nor U7820 (N_7820,N_2792,N_3803);
nor U7821 (N_7821,N_2857,N_3132);
nor U7822 (N_7822,N_275,N_2952);
nor U7823 (N_7823,N_1695,N_2032);
nor U7824 (N_7824,N_1699,N_4479);
nor U7825 (N_7825,N_1074,N_4105);
or U7826 (N_7826,N_380,N_489);
and U7827 (N_7827,N_3005,N_2317);
nor U7828 (N_7828,N_4615,N_361);
xnor U7829 (N_7829,N_1829,N_937);
xnor U7830 (N_7830,N_4519,N_1607);
and U7831 (N_7831,N_3922,N_4512);
and U7832 (N_7832,N_1775,N_3079);
or U7833 (N_7833,N_4810,N_2425);
nor U7834 (N_7834,N_3489,N_193);
xor U7835 (N_7835,N_1392,N_1657);
and U7836 (N_7836,N_4875,N_444);
or U7837 (N_7837,N_621,N_3760);
xor U7838 (N_7838,N_2141,N_2109);
or U7839 (N_7839,N_3362,N_2220);
nor U7840 (N_7840,N_927,N_150);
nor U7841 (N_7841,N_4610,N_3238);
xor U7842 (N_7842,N_849,N_4235);
nand U7843 (N_7843,N_2364,N_4105);
or U7844 (N_7844,N_3219,N_3388);
nor U7845 (N_7845,N_3386,N_3719);
nand U7846 (N_7846,N_2722,N_4318);
and U7847 (N_7847,N_3546,N_691);
xnor U7848 (N_7848,N_3026,N_3588);
or U7849 (N_7849,N_49,N_3898);
or U7850 (N_7850,N_4453,N_965);
nand U7851 (N_7851,N_3431,N_2046);
xnor U7852 (N_7852,N_1217,N_3094);
xnor U7853 (N_7853,N_3679,N_2058);
xor U7854 (N_7854,N_1841,N_4133);
and U7855 (N_7855,N_1547,N_563);
and U7856 (N_7856,N_4185,N_4182);
or U7857 (N_7857,N_4270,N_4652);
and U7858 (N_7858,N_2942,N_167);
or U7859 (N_7859,N_4305,N_2666);
nor U7860 (N_7860,N_831,N_3004);
xor U7861 (N_7861,N_4808,N_4477);
or U7862 (N_7862,N_45,N_3720);
and U7863 (N_7863,N_3631,N_1640);
nor U7864 (N_7864,N_3036,N_3470);
nand U7865 (N_7865,N_4054,N_2758);
or U7866 (N_7866,N_2027,N_2711);
xnor U7867 (N_7867,N_4248,N_1327);
and U7868 (N_7868,N_2307,N_2981);
xor U7869 (N_7869,N_836,N_4895);
or U7870 (N_7870,N_3262,N_2582);
nand U7871 (N_7871,N_3534,N_3367);
and U7872 (N_7872,N_2920,N_3506);
or U7873 (N_7873,N_3009,N_3771);
or U7874 (N_7874,N_3495,N_543);
xor U7875 (N_7875,N_3503,N_3133);
and U7876 (N_7876,N_4383,N_4568);
nand U7877 (N_7877,N_4126,N_2352);
nor U7878 (N_7878,N_3000,N_1322);
xor U7879 (N_7879,N_3650,N_1339);
nand U7880 (N_7880,N_567,N_178);
or U7881 (N_7881,N_2313,N_4390);
or U7882 (N_7882,N_3618,N_17);
nor U7883 (N_7883,N_2632,N_2880);
nor U7884 (N_7884,N_4506,N_2966);
nor U7885 (N_7885,N_3012,N_4255);
nor U7886 (N_7886,N_1116,N_1435);
or U7887 (N_7887,N_3284,N_877);
or U7888 (N_7888,N_182,N_3236);
xnor U7889 (N_7889,N_700,N_829);
xnor U7890 (N_7890,N_3996,N_1489);
or U7891 (N_7891,N_4270,N_790);
nand U7892 (N_7892,N_274,N_2118);
or U7893 (N_7893,N_4869,N_3137);
nor U7894 (N_7894,N_4839,N_4867);
xor U7895 (N_7895,N_595,N_4395);
and U7896 (N_7896,N_4311,N_2526);
or U7897 (N_7897,N_4110,N_2368);
nand U7898 (N_7898,N_3707,N_303);
or U7899 (N_7899,N_158,N_695);
nand U7900 (N_7900,N_3282,N_4516);
xnor U7901 (N_7901,N_1403,N_328);
nand U7902 (N_7902,N_4384,N_3267);
nand U7903 (N_7903,N_1071,N_4042);
or U7904 (N_7904,N_4855,N_4308);
or U7905 (N_7905,N_3103,N_1373);
nand U7906 (N_7906,N_4453,N_2343);
xor U7907 (N_7907,N_2668,N_146);
nand U7908 (N_7908,N_4919,N_4788);
or U7909 (N_7909,N_1990,N_1);
nand U7910 (N_7910,N_170,N_4437);
and U7911 (N_7911,N_3924,N_2905);
or U7912 (N_7912,N_4337,N_3261);
nor U7913 (N_7913,N_3024,N_3365);
nand U7914 (N_7914,N_3810,N_721);
nand U7915 (N_7915,N_4857,N_1029);
and U7916 (N_7916,N_4453,N_2233);
nor U7917 (N_7917,N_1357,N_1774);
xor U7918 (N_7918,N_3931,N_1353);
and U7919 (N_7919,N_1825,N_2215);
nor U7920 (N_7920,N_870,N_1314);
or U7921 (N_7921,N_2591,N_2723);
nor U7922 (N_7922,N_2808,N_975);
nand U7923 (N_7923,N_38,N_1114);
nand U7924 (N_7924,N_3251,N_348);
xnor U7925 (N_7925,N_1673,N_2940);
nor U7926 (N_7926,N_1704,N_2802);
or U7927 (N_7927,N_3497,N_2905);
and U7928 (N_7928,N_4844,N_2261);
nor U7929 (N_7929,N_2413,N_387);
xnor U7930 (N_7930,N_3657,N_1174);
xnor U7931 (N_7931,N_4945,N_4900);
or U7932 (N_7932,N_1421,N_832);
nand U7933 (N_7933,N_1333,N_4568);
and U7934 (N_7934,N_1078,N_2729);
nand U7935 (N_7935,N_1601,N_4715);
nor U7936 (N_7936,N_1982,N_1521);
nor U7937 (N_7937,N_788,N_3174);
and U7938 (N_7938,N_1535,N_540);
nor U7939 (N_7939,N_1005,N_4256);
nand U7940 (N_7940,N_86,N_1837);
nor U7941 (N_7941,N_1409,N_857);
or U7942 (N_7942,N_3920,N_18);
nand U7943 (N_7943,N_3194,N_1005);
nor U7944 (N_7944,N_4362,N_3274);
xor U7945 (N_7945,N_3811,N_3533);
nand U7946 (N_7946,N_3297,N_987);
and U7947 (N_7947,N_4771,N_1070);
nand U7948 (N_7948,N_461,N_1744);
or U7949 (N_7949,N_4125,N_3362);
nand U7950 (N_7950,N_1651,N_221);
nand U7951 (N_7951,N_3369,N_3623);
or U7952 (N_7952,N_1484,N_3633);
xnor U7953 (N_7953,N_1732,N_3481);
or U7954 (N_7954,N_2065,N_1446);
nand U7955 (N_7955,N_369,N_3596);
and U7956 (N_7956,N_2383,N_700);
or U7957 (N_7957,N_1251,N_4401);
or U7958 (N_7958,N_2180,N_1190);
and U7959 (N_7959,N_2326,N_3695);
nor U7960 (N_7960,N_4749,N_1541);
nand U7961 (N_7961,N_3261,N_4776);
and U7962 (N_7962,N_4806,N_3165);
xor U7963 (N_7963,N_758,N_1591);
nor U7964 (N_7964,N_3156,N_1150);
nor U7965 (N_7965,N_4787,N_4019);
or U7966 (N_7966,N_3681,N_3030);
or U7967 (N_7967,N_1487,N_637);
or U7968 (N_7968,N_2359,N_3016);
nand U7969 (N_7969,N_1528,N_4418);
and U7970 (N_7970,N_925,N_4874);
xor U7971 (N_7971,N_4813,N_316);
nor U7972 (N_7972,N_1632,N_1316);
and U7973 (N_7973,N_2244,N_3821);
and U7974 (N_7974,N_1184,N_3689);
nand U7975 (N_7975,N_3241,N_2929);
nor U7976 (N_7976,N_4334,N_2408);
nand U7977 (N_7977,N_2208,N_265);
and U7978 (N_7978,N_1347,N_4752);
and U7979 (N_7979,N_2341,N_1279);
nor U7980 (N_7980,N_1220,N_2630);
xor U7981 (N_7981,N_2300,N_4582);
xnor U7982 (N_7982,N_1229,N_4981);
nand U7983 (N_7983,N_2700,N_2516);
nand U7984 (N_7984,N_3753,N_1918);
xnor U7985 (N_7985,N_2385,N_2260);
or U7986 (N_7986,N_1092,N_1979);
xor U7987 (N_7987,N_2237,N_396);
xor U7988 (N_7988,N_4769,N_986);
nor U7989 (N_7989,N_4937,N_1030);
nand U7990 (N_7990,N_3956,N_4924);
nor U7991 (N_7991,N_130,N_3794);
nor U7992 (N_7992,N_3381,N_1820);
nand U7993 (N_7993,N_2043,N_2820);
nor U7994 (N_7994,N_4923,N_3555);
nand U7995 (N_7995,N_2404,N_1935);
nand U7996 (N_7996,N_2470,N_1417);
nand U7997 (N_7997,N_1310,N_463);
nor U7998 (N_7998,N_1414,N_416);
and U7999 (N_7999,N_3579,N_2450);
or U8000 (N_8000,N_3991,N_3589);
or U8001 (N_8001,N_3396,N_4276);
nor U8002 (N_8002,N_2745,N_4495);
xor U8003 (N_8003,N_2087,N_4144);
or U8004 (N_8004,N_3165,N_2605);
nand U8005 (N_8005,N_1127,N_231);
nand U8006 (N_8006,N_918,N_2088);
and U8007 (N_8007,N_2273,N_3239);
nor U8008 (N_8008,N_577,N_4887);
nand U8009 (N_8009,N_3927,N_3449);
nor U8010 (N_8010,N_4768,N_1279);
xor U8011 (N_8011,N_2103,N_2489);
nor U8012 (N_8012,N_840,N_1130);
and U8013 (N_8013,N_2440,N_3887);
and U8014 (N_8014,N_4128,N_3249);
xor U8015 (N_8015,N_3456,N_1125);
nand U8016 (N_8016,N_802,N_3064);
and U8017 (N_8017,N_4329,N_4629);
nand U8018 (N_8018,N_4532,N_1908);
and U8019 (N_8019,N_368,N_2176);
or U8020 (N_8020,N_1742,N_2916);
and U8021 (N_8021,N_3242,N_1055);
nor U8022 (N_8022,N_155,N_4899);
or U8023 (N_8023,N_1036,N_3239);
nand U8024 (N_8024,N_3118,N_1918);
or U8025 (N_8025,N_924,N_4614);
nor U8026 (N_8026,N_3253,N_1292);
and U8027 (N_8027,N_3462,N_4788);
and U8028 (N_8028,N_4033,N_4979);
or U8029 (N_8029,N_4051,N_12);
or U8030 (N_8030,N_1544,N_2528);
xor U8031 (N_8031,N_4834,N_3689);
xnor U8032 (N_8032,N_3641,N_2200);
and U8033 (N_8033,N_4265,N_2255);
xnor U8034 (N_8034,N_4273,N_1561);
xnor U8035 (N_8035,N_3555,N_2388);
or U8036 (N_8036,N_4329,N_3203);
or U8037 (N_8037,N_3428,N_4066);
nand U8038 (N_8038,N_727,N_3123);
xor U8039 (N_8039,N_773,N_4907);
or U8040 (N_8040,N_3324,N_479);
nor U8041 (N_8041,N_2836,N_3271);
and U8042 (N_8042,N_3634,N_3628);
nand U8043 (N_8043,N_3183,N_3976);
xor U8044 (N_8044,N_1625,N_208);
nor U8045 (N_8045,N_3836,N_839);
xnor U8046 (N_8046,N_3607,N_631);
nand U8047 (N_8047,N_59,N_2059);
and U8048 (N_8048,N_3997,N_439);
or U8049 (N_8049,N_3907,N_3714);
xor U8050 (N_8050,N_2743,N_2096);
nor U8051 (N_8051,N_3012,N_3507);
nor U8052 (N_8052,N_4040,N_1347);
nor U8053 (N_8053,N_4736,N_4623);
nor U8054 (N_8054,N_4235,N_1950);
nand U8055 (N_8055,N_1867,N_3433);
nand U8056 (N_8056,N_337,N_1842);
xor U8057 (N_8057,N_4503,N_777);
and U8058 (N_8058,N_1147,N_593);
and U8059 (N_8059,N_4430,N_1833);
nand U8060 (N_8060,N_4703,N_2999);
and U8061 (N_8061,N_2814,N_473);
xor U8062 (N_8062,N_371,N_4316);
xnor U8063 (N_8063,N_2161,N_2441);
nand U8064 (N_8064,N_3350,N_4633);
or U8065 (N_8065,N_3727,N_3444);
and U8066 (N_8066,N_3309,N_3760);
nor U8067 (N_8067,N_354,N_3811);
and U8068 (N_8068,N_1395,N_371);
xor U8069 (N_8069,N_2494,N_4848);
nand U8070 (N_8070,N_707,N_2672);
or U8071 (N_8071,N_2635,N_3883);
or U8072 (N_8072,N_1854,N_647);
or U8073 (N_8073,N_1550,N_1144);
nand U8074 (N_8074,N_1371,N_4927);
or U8075 (N_8075,N_4255,N_1071);
or U8076 (N_8076,N_361,N_326);
xor U8077 (N_8077,N_2518,N_3403);
or U8078 (N_8078,N_431,N_2151);
nor U8079 (N_8079,N_3179,N_1664);
or U8080 (N_8080,N_2663,N_4145);
nand U8081 (N_8081,N_3217,N_4132);
and U8082 (N_8082,N_4788,N_4170);
or U8083 (N_8083,N_4367,N_3541);
xor U8084 (N_8084,N_1244,N_1524);
nor U8085 (N_8085,N_3395,N_675);
nand U8086 (N_8086,N_1589,N_1129);
nor U8087 (N_8087,N_534,N_3527);
or U8088 (N_8088,N_4446,N_1593);
nor U8089 (N_8089,N_1161,N_1180);
or U8090 (N_8090,N_1587,N_2803);
nand U8091 (N_8091,N_4418,N_213);
or U8092 (N_8092,N_970,N_4779);
nand U8093 (N_8093,N_1548,N_604);
nor U8094 (N_8094,N_527,N_4376);
nand U8095 (N_8095,N_2783,N_926);
xnor U8096 (N_8096,N_4779,N_4186);
nor U8097 (N_8097,N_1734,N_4169);
and U8098 (N_8098,N_552,N_4999);
or U8099 (N_8099,N_2817,N_2641);
or U8100 (N_8100,N_4141,N_2005);
nand U8101 (N_8101,N_2809,N_3170);
and U8102 (N_8102,N_3375,N_106);
nor U8103 (N_8103,N_3179,N_1866);
and U8104 (N_8104,N_2492,N_2370);
or U8105 (N_8105,N_4869,N_4395);
xnor U8106 (N_8106,N_1786,N_2879);
or U8107 (N_8107,N_3212,N_1561);
xnor U8108 (N_8108,N_3550,N_4199);
nor U8109 (N_8109,N_48,N_3366);
or U8110 (N_8110,N_1064,N_1160);
xnor U8111 (N_8111,N_1236,N_4474);
nor U8112 (N_8112,N_65,N_2534);
and U8113 (N_8113,N_2319,N_1406);
nand U8114 (N_8114,N_4188,N_20);
nor U8115 (N_8115,N_2312,N_1817);
nand U8116 (N_8116,N_4028,N_4610);
and U8117 (N_8117,N_2403,N_2346);
xor U8118 (N_8118,N_3119,N_4150);
nand U8119 (N_8119,N_3747,N_4753);
or U8120 (N_8120,N_2181,N_508);
or U8121 (N_8121,N_2273,N_4061);
xor U8122 (N_8122,N_1163,N_309);
nand U8123 (N_8123,N_3711,N_3743);
or U8124 (N_8124,N_2697,N_2829);
or U8125 (N_8125,N_1293,N_2603);
nand U8126 (N_8126,N_1048,N_3709);
xnor U8127 (N_8127,N_2612,N_152);
xnor U8128 (N_8128,N_3131,N_688);
nand U8129 (N_8129,N_3297,N_854);
or U8130 (N_8130,N_3889,N_4888);
xnor U8131 (N_8131,N_3296,N_4810);
and U8132 (N_8132,N_3096,N_3709);
xnor U8133 (N_8133,N_240,N_2700);
xor U8134 (N_8134,N_1192,N_4138);
xor U8135 (N_8135,N_421,N_1935);
nand U8136 (N_8136,N_3837,N_1574);
nor U8137 (N_8137,N_3192,N_558);
or U8138 (N_8138,N_2153,N_3700);
nand U8139 (N_8139,N_4030,N_237);
xor U8140 (N_8140,N_1574,N_3230);
nor U8141 (N_8141,N_4980,N_887);
nand U8142 (N_8142,N_2812,N_3555);
or U8143 (N_8143,N_1648,N_3978);
xor U8144 (N_8144,N_1076,N_2419);
xnor U8145 (N_8145,N_4916,N_4071);
and U8146 (N_8146,N_240,N_3310);
nand U8147 (N_8147,N_2606,N_4512);
and U8148 (N_8148,N_43,N_1547);
and U8149 (N_8149,N_1477,N_3022);
and U8150 (N_8150,N_1176,N_1242);
nand U8151 (N_8151,N_4370,N_149);
nor U8152 (N_8152,N_468,N_4488);
nand U8153 (N_8153,N_3533,N_1964);
nor U8154 (N_8154,N_1071,N_1934);
or U8155 (N_8155,N_1091,N_2734);
nand U8156 (N_8156,N_1842,N_4570);
nor U8157 (N_8157,N_4694,N_1770);
and U8158 (N_8158,N_2447,N_4247);
and U8159 (N_8159,N_4801,N_3006);
or U8160 (N_8160,N_3272,N_1333);
nor U8161 (N_8161,N_1116,N_167);
xnor U8162 (N_8162,N_4517,N_1517);
and U8163 (N_8163,N_2889,N_3118);
nor U8164 (N_8164,N_2198,N_3938);
nor U8165 (N_8165,N_745,N_4982);
and U8166 (N_8166,N_3143,N_3420);
and U8167 (N_8167,N_2447,N_679);
or U8168 (N_8168,N_4385,N_4303);
nand U8169 (N_8169,N_4911,N_2854);
and U8170 (N_8170,N_2534,N_1606);
and U8171 (N_8171,N_4463,N_1909);
or U8172 (N_8172,N_1880,N_2933);
or U8173 (N_8173,N_3714,N_1065);
nor U8174 (N_8174,N_4625,N_1885);
or U8175 (N_8175,N_3945,N_2515);
nor U8176 (N_8176,N_4224,N_3042);
nand U8177 (N_8177,N_3594,N_2124);
nand U8178 (N_8178,N_835,N_3744);
xnor U8179 (N_8179,N_2812,N_3034);
xnor U8180 (N_8180,N_624,N_1809);
xnor U8181 (N_8181,N_60,N_3176);
nor U8182 (N_8182,N_982,N_291);
nor U8183 (N_8183,N_3316,N_780);
nor U8184 (N_8184,N_2772,N_3411);
nand U8185 (N_8185,N_4329,N_1586);
and U8186 (N_8186,N_592,N_333);
nand U8187 (N_8187,N_1278,N_2952);
nand U8188 (N_8188,N_22,N_3127);
or U8189 (N_8189,N_2540,N_2220);
nand U8190 (N_8190,N_965,N_1488);
and U8191 (N_8191,N_3519,N_4367);
xnor U8192 (N_8192,N_4958,N_3926);
nand U8193 (N_8193,N_1720,N_138);
and U8194 (N_8194,N_565,N_3524);
nor U8195 (N_8195,N_4346,N_4622);
xnor U8196 (N_8196,N_4383,N_1477);
nor U8197 (N_8197,N_4145,N_4590);
and U8198 (N_8198,N_4428,N_1695);
xor U8199 (N_8199,N_3983,N_760);
xor U8200 (N_8200,N_2460,N_1068);
and U8201 (N_8201,N_2617,N_3179);
nor U8202 (N_8202,N_4472,N_3271);
nor U8203 (N_8203,N_2337,N_4959);
and U8204 (N_8204,N_1578,N_2428);
xnor U8205 (N_8205,N_2369,N_3935);
nand U8206 (N_8206,N_3400,N_2950);
and U8207 (N_8207,N_350,N_872);
or U8208 (N_8208,N_3509,N_4779);
nand U8209 (N_8209,N_133,N_207);
and U8210 (N_8210,N_4728,N_2918);
xor U8211 (N_8211,N_1015,N_1183);
or U8212 (N_8212,N_4079,N_3356);
xor U8213 (N_8213,N_451,N_3909);
xor U8214 (N_8214,N_583,N_4888);
nand U8215 (N_8215,N_2537,N_4593);
or U8216 (N_8216,N_2555,N_301);
xor U8217 (N_8217,N_805,N_450);
or U8218 (N_8218,N_2632,N_40);
and U8219 (N_8219,N_2954,N_2376);
xor U8220 (N_8220,N_4169,N_4952);
or U8221 (N_8221,N_4664,N_3145);
or U8222 (N_8222,N_3129,N_4496);
and U8223 (N_8223,N_3374,N_1803);
and U8224 (N_8224,N_4463,N_2137);
or U8225 (N_8225,N_1801,N_3188);
nor U8226 (N_8226,N_1071,N_885);
or U8227 (N_8227,N_4397,N_2692);
nand U8228 (N_8228,N_4868,N_61);
and U8229 (N_8229,N_3273,N_2503);
and U8230 (N_8230,N_840,N_2786);
xnor U8231 (N_8231,N_4569,N_4265);
nor U8232 (N_8232,N_4585,N_4014);
and U8233 (N_8233,N_1532,N_885);
nand U8234 (N_8234,N_1461,N_356);
nand U8235 (N_8235,N_3952,N_990);
and U8236 (N_8236,N_4736,N_4556);
and U8237 (N_8237,N_2371,N_2610);
nor U8238 (N_8238,N_3468,N_4797);
nor U8239 (N_8239,N_4555,N_4478);
xor U8240 (N_8240,N_3242,N_1071);
or U8241 (N_8241,N_2126,N_477);
or U8242 (N_8242,N_586,N_1845);
and U8243 (N_8243,N_1165,N_1612);
xnor U8244 (N_8244,N_4882,N_171);
nand U8245 (N_8245,N_4682,N_2103);
xor U8246 (N_8246,N_692,N_3032);
nor U8247 (N_8247,N_4641,N_950);
and U8248 (N_8248,N_2177,N_3899);
nor U8249 (N_8249,N_3625,N_4205);
and U8250 (N_8250,N_4930,N_754);
nor U8251 (N_8251,N_487,N_2110);
nand U8252 (N_8252,N_3508,N_364);
and U8253 (N_8253,N_175,N_966);
or U8254 (N_8254,N_3068,N_2591);
xnor U8255 (N_8255,N_1146,N_172);
xnor U8256 (N_8256,N_4346,N_1394);
nor U8257 (N_8257,N_3895,N_3187);
or U8258 (N_8258,N_4073,N_2326);
xnor U8259 (N_8259,N_3441,N_4269);
nand U8260 (N_8260,N_3301,N_423);
nand U8261 (N_8261,N_1388,N_1201);
and U8262 (N_8262,N_1091,N_1903);
nand U8263 (N_8263,N_2277,N_4637);
xnor U8264 (N_8264,N_1708,N_3107);
and U8265 (N_8265,N_2245,N_3295);
xnor U8266 (N_8266,N_821,N_1563);
or U8267 (N_8267,N_1449,N_4448);
nor U8268 (N_8268,N_3301,N_4664);
or U8269 (N_8269,N_3635,N_2742);
nand U8270 (N_8270,N_4717,N_4894);
nand U8271 (N_8271,N_2985,N_4763);
nand U8272 (N_8272,N_3084,N_517);
xor U8273 (N_8273,N_4113,N_2417);
xor U8274 (N_8274,N_2803,N_3993);
nor U8275 (N_8275,N_2489,N_896);
and U8276 (N_8276,N_3824,N_3910);
xnor U8277 (N_8277,N_4078,N_350);
nand U8278 (N_8278,N_3807,N_4991);
or U8279 (N_8279,N_1605,N_3186);
nor U8280 (N_8280,N_1808,N_2401);
and U8281 (N_8281,N_4668,N_3433);
xor U8282 (N_8282,N_2116,N_631);
and U8283 (N_8283,N_1692,N_1912);
nor U8284 (N_8284,N_1138,N_2238);
nand U8285 (N_8285,N_953,N_3439);
nand U8286 (N_8286,N_538,N_1552);
nor U8287 (N_8287,N_3395,N_225);
nor U8288 (N_8288,N_3728,N_910);
or U8289 (N_8289,N_4869,N_251);
nor U8290 (N_8290,N_834,N_3021);
and U8291 (N_8291,N_3185,N_1493);
nor U8292 (N_8292,N_1732,N_591);
and U8293 (N_8293,N_3023,N_2466);
nand U8294 (N_8294,N_4582,N_1788);
nand U8295 (N_8295,N_2940,N_1641);
or U8296 (N_8296,N_108,N_2641);
nand U8297 (N_8297,N_3687,N_4191);
and U8298 (N_8298,N_1382,N_2755);
and U8299 (N_8299,N_2272,N_3327);
nand U8300 (N_8300,N_1347,N_2672);
nor U8301 (N_8301,N_801,N_1852);
and U8302 (N_8302,N_896,N_4102);
and U8303 (N_8303,N_4984,N_4309);
nand U8304 (N_8304,N_292,N_2274);
or U8305 (N_8305,N_2572,N_3503);
and U8306 (N_8306,N_4170,N_4110);
nand U8307 (N_8307,N_4278,N_2909);
nor U8308 (N_8308,N_4125,N_1588);
xor U8309 (N_8309,N_3370,N_1730);
nor U8310 (N_8310,N_946,N_4537);
or U8311 (N_8311,N_3523,N_1881);
and U8312 (N_8312,N_4836,N_4873);
nand U8313 (N_8313,N_25,N_1090);
or U8314 (N_8314,N_98,N_3996);
nand U8315 (N_8315,N_1265,N_4872);
or U8316 (N_8316,N_317,N_4456);
nand U8317 (N_8317,N_1947,N_4492);
or U8318 (N_8318,N_1468,N_4137);
and U8319 (N_8319,N_431,N_3947);
xor U8320 (N_8320,N_4254,N_4477);
xnor U8321 (N_8321,N_76,N_504);
and U8322 (N_8322,N_2011,N_1580);
and U8323 (N_8323,N_3037,N_3434);
nand U8324 (N_8324,N_2137,N_2775);
nand U8325 (N_8325,N_4569,N_4934);
nor U8326 (N_8326,N_3340,N_3563);
and U8327 (N_8327,N_3816,N_123);
or U8328 (N_8328,N_239,N_3431);
xnor U8329 (N_8329,N_214,N_699);
xnor U8330 (N_8330,N_2993,N_1170);
nand U8331 (N_8331,N_4767,N_887);
nand U8332 (N_8332,N_3654,N_2330);
and U8333 (N_8333,N_2809,N_1101);
nor U8334 (N_8334,N_3596,N_4120);
nand U8335 (N_8335,N_2805,N_608);
nand U8336 (N_8336,N_3647,N_3127);
xor U8337 (N_8337,N_3377,N_3258);
or U8338 (N_8338,N_401,N_1347);
nor U8339 (N_8339,N_3012,N_3055);
or U8340 (N_8340,N_70,N_4507);
and U8341 (N_8341,N_2429,N_973);
or U8342 (N_8342,N_2322,N_2804);
nor U8343 (N_8343,N_2296,N_2731);
or U8344 (N_8344,N_4643,N_3228);
nor U8345 (N_8345,N_3061,N_4048);
and U8346 (N_8346,N_4795,N_4706);
or U8347 (N_8347,N_3650,N_1749);
xnor U8348 (N_8348,N_4842,N_4007);
and U8349 (N_8349,N_961,N_589);
or U8350 (N_8350,N_4532,N_2681);
xor U8351 (N_8351,N_1972,N_255);
or U8352 (N_8352,N_4385,N_345);
nand U8353 (N_8353,N_990,N_1830);
nand U8354 (N_8354,N_767,N_3178);
nand U8355 (N_8355,N_1601,N_717);
or U8356 (N_8356,N_3415,N_4233);
and U8357 (N_8357,N_148,N_2466);
or U8358 (N_8358,N_3382,N_2831);
and U8359 (N_8359,N_2580,N_1848);
and U8360 (N_8360,N_2271,N_4457);
or U8361 (N_8361,N_1916,N_2308);
xor U8362 (N_8362,N_4675,N_4817);
nand U8363 (N_8363,N_799,N_4136);
or U8364 (N_8364,N_4715,N_1558);
nor U8365 (N_8365,N_2442,N_4032);
and U8366 (N_8366,N_1798,N_4550);
xnor U8367 (N_8367,N_3224,N_4144);
and U8368 (N_8368,N_2401,N_3945);
nor U8369 (N_8369,N_1352,N_1147);
and U8370 (N_8370,N_3228,N_4143);
and U8371 (N_8371,N_177,N_521);
nor U8372 (N_8372,N_2993,N_1898);
xnor U8373 (N_8373,N_2864,N_3270);
and U8374 (N_8374,N_2707,N_27);
and U8375 (N_8375,N_1544,N_746);
and U8376 (N_8376,N_3761,N_1825);
and U8377 (N_8377,N_2659,N_1704);
xnor U8378 (N_8378,N_2236,N_126);
xnor U8379 (N_8379,N_3592,N_3974);
xor U8380 (N_8380,N_2694,N_4292);
and U8381 (N_8381,N_2725,N_4628);
or U8382 (N_8382,N_2214,N_947);
and U8383 (N_8383,N_3638,N_4999);
or U8384 (N_8384,N_3923,N_4254);
xor U8385 (N_8385,N_3598,N_4202);
and U8386 (N_8386,N_339,N_256);
or U8387 (N_8387,N_2014,N_2395);
nor U8388 (N_8388,N_2753,N_1209);
nand U8389 (N_8389,N_2221,N_3768);
or U8390 (N_8390,N_626,N_1181);
and U8391 (N_8391,N_1416,N_3908);
xnor U8392 (N_8392,N_1977,N_4097);
or U8393 (N_8393,N_3145,N_3039);
and U8394 (N_8394,N_4569,N_1949);
xor U8395 (N_8395,N_1294,N_832);
xnor U8396 (N_8396,N_3798,N_407);
nor U8397 (N_8397,N_2141,N_4949);
nand U8398 (N_8398,N_3570,N_1380);
or U8399 (N_8399,N_3557,N_2842);
and U8400 (N_8400,N_3944,N_2);
and U8401 (N_8401,N_2536,N_746);
or U8402 (N_8402,N_1020,N_4455);
or U8403 (N_8403,N_693,N_3108);
and U8404 (N_8404,N_113,N_2724);
nand U8405 (N_8405,N_2050,N_1258);
xor U8406 (N_8406,N_1052,N_1215);
or U8407 (N_8407,N_1348,N_4607);
xor U8408 (N_8408,N_4162,N_1193);
xnor U8409 (N_8409,N_423,N_4092);
nand U8410 (N_8410,N_3362,N_2092);
or U8411 (N_8411,N_2249,N_4817);
xor U8412 (N_8412,N_1683,N_1007);
nor U8413 (N_8413,N_1715,N_693);
nand U8414 (N_8414,N_989,N_595);
nor U8415 (N_8415,N_4989,N_3303);
nor U8416 (N_8416,N_4562,N_2066);
nor U8417 (N_8417,N_1381,N_2817);
or U8418 (N_8418,N_4594,N_1725);
or U8419 (N_8419,N_4992,N_2250);
nor U8420 (N_8420,N_4173,N_1623);
and U8421 (N_8421,N_4027,N_3784);
nor U8422 (N_8422,N_1042,N_3875);
or U8423 (N_8423,N_1719,N_3071);
or U8424 (N_8424,N_3184,N_3113);
nand U8425 (N_8425,N_3062,N_2918);
or U8426 (N_8426,N_184,N_392);
and U8427 (N_8427,N_1921,N_2207);
or U8428 (N_8428,N_1001,N_2542);
or U8429 (N_8429,N_1048,N_3718);
or U8430 (N_8430,N_886,N_436);
nor U8431 (N_8431,N_3192,N_2162);
xnor U8432 (N_8432,N_2454,N_4974);
or U8433 (N_8433,N_1239,N_2103);
nand U8434 (N_8434,N_660,N_4199);
nor U8435 (N_8435,N_55,N_2240);
or U8436 (N_8436,N_3641,N_4125);
and U8437 (N_8437,N_3095,N_2659);
nand U8438 (N_8438,N_4974,N_2967);
nor U8439 (N_8439,N_3771,N_3000);
and U8440 (N_8440,N_1727,N_3513);
or U8441 (N_8441,N_1605,N_2761);
or U8442 (N_8442,N_1044,N_2732);
xnor U8443 (N_8443,N_2824,N_1748);
nor U8444 (N_8444,N_4091,N_2965);
nand U8445 (N_8445,N_4225,N_463);
nand U8446 (N_8446,N_559,N_4082);
xor U8447 (N_8447,N_2065,N_2525);
and U8448 (N_8448,N_2887,N_3702);
or U8449 (N_8449,N_316,N_626);
nand U8450 (N_8450,N_697,N_3812);
nand U8451 (N_8451,N_3081,N_1318);
nand U8452 (N_8452,N_948,N_2367);
and U8453 (N_8453,N_383,N_3034);
xor U8454 (N_8454,N_1810,N_2150);
nor U8455 (N_8455,N_840,N_385);
or U8456 (N_8456,N_783,N_3978);
xor U8457 (N_8457,N_4672,N_4470);
xnor U8458 (N_8458,N_4745,N_3056);
nor U8459 (N_8459,N_2421,N_3651);
and U8460 (N_8460,N_3216,N_1502);
or U8461 (N_8461,N_1597,N_1951);
and U8462 (N_8462,N_2265,N_3117);
or U8463 (N_8463,N_4043,N_1719);
or U8464 (N_8464,N_3802,N_4684);
or U8465 (N_8465,N_1302,N_1828);
xnor U8466 (N_8466,N_1605,N_3009);
and U8467 (N_8467,N_4967,N_3666);
nand U8468 (N_8468,N_403,N_3905);
nand U8469 (N_8469,N_1259,N_1822);
or U8470 (N_8470,N_1726,N_541);
or U8471 (N_8471,N_1795,N_4173);
xnor U8472 (N_8472,N_208,N_4957);
or U8473 (N_8473,N_2793,N_4303);
nand U8474 (N_8474,N_1552,N_4052);
nor U8475 (N_8475,N_4812,N_2639);
and U8476 (N_8476,N_1033,N_2436);
xor U8477 (N_8477,N_138,N_2378);
nor U8478 (N_8478,N_4950,N_921);
or U8479 (N_8479,N_3551,N_4372);
nor U8480 (N_8480,N_1662,N_2519);
nor U8481 (N_8481,N_330,N_3033);
or U8482 (N_8482,N_4273,N_3292);
and U8483 (N_8483,N_2100,N_2070);
nor U8484 (N_8484,N_999,N_1219);
and U8485 (N_8485,N_2995,N_2702);
or U8486 (N_8486,N_1649,N_76);
nor U8487 (N_8487,N_3475,N_4048);
or U8488 (N_8488,N_1244,N_2666);
nor U8489 (N_8489,N_1973,N_3555);
nand U8490 (N_8490,N_3025,N_2752);
nand U8491 (N_8491,N_2649,N_2569);
and U8492 (N_8492,N_1296,N_3182);
and U8493 (N_8493,N_3374,N_2342);
nand U8494 (N_8494,N_1763,N_1636);
and U8495 (N_8495,N_4193,N_1721);
xnor U8496 (N_8496,N_4833,N_840);
xnor U8497 (N_8497,N_2298,N_4511);
nor U8498 (N_8498,N_1188,N_2039);
xor U8499 (N_8499,N_3622,N_1026);
and U8500 (N_8500,N_4874,N_1820);
or U8501 (N_8501,N_265,N_161);
and U8502 (N_8502,N_2320,N_1729);
nand U8503 (N_8503,N_551,N_3087);
or U8504 (N_8504,N_2089,N_202);
nor U8505 (N_8505,N_3074,N_2797);
xor U8506 (N_8506,N_4866,N_2618);
or U8507 (N_8507,N_1001,N_4568);
nor U8508 (N_8508,N_801,N_3680);
xor U8509 (N_8509,N_2845,N_4550);
and U8510 (N_8510,N_1926,N_2469);
and U8511 (N_8511,N_1899,N_886);
or U8512 (N_8512,N_106,N_3129);
nor U8513 (N_8513,N_4393,N_3045);
xor U8514 (N_8514,N_297,N_649);
and U8515 (N_8515,N_2420,N_4278);
nand U8516 (N_8516,N_3904,N_1805);
and U8517 (N_8517,N_4673,N_3295);
xnor U8518 (N_8518,N_4585,N_4124);
xnor U8519 (N_8519,N_1002,N_460);
nor U8520 (N_8520,N_4408,N_4493);
and U8521 (N_8521,N_70,N_3625);
nand U8522 (N_8522,N_2329,N_1576);
and U8523 (N_8523,N_3055,N_3163);
xor U8524 (N_8524,N_4300,N_1123);
nand U8525 (N_8525,N_3912,N_2918);
nand U8526 (N_8526,N_439,N_2499);
nor U8527 (N_8527,N_4719,N_2551);
and U8528 (N_8528,N_1937,N_3101);
and U8529 (N_8529,N_19,N_2079);
xor U8530 (N_8530,N_264,N_2664);
and U8531 (N_8531,N_227,N_4645);
xor U8532 (N_8532,N_1136,N_2887);
or U8533 (N_8533,N_1147,N_1995);
xor U8534 (N_8534,N_2633,N_1015);
xor U8535 (N_8535,N_1926,N_828);
or U8536 (N_8536,N_3435,N_2976);
xnor U8537 (N_8537,N_247,N_3471);
or U8538 (N_8538,N_1985,N_1454);
nor U8539 (N_8539,N_2883,N_3334);
and U8540 (N_8540,N_3393,N_1357);
xnor U8541 (N_8541,N_219,N_4384);
xnor U8542 (N_8542,N_3074,N_721);
nor U8543 (N_8543,N_3377,N_466);
nor U8544 (N_8544,N_1007,N_438);
xor U8545 (N_8545,N_77,N_4636);
and U8546 (N_8546,N_2989,N_1413);
xnor U8547 (N_8547,N_2895,N_1001);
xnor U8548 (N_8548,N_3914,N_2394);
and U8549 (N_8549,N_2488,N_74);
or U8550 (N_8550,N_1217,N_1502);
and U8551 (N_8551,N_4842,N_2246);
or U8552 (N_8552,N_4317,N_681);
xnor U8553 (N_8553,N_4974,N_3821);
or U8554 (N_8554,N_4496,N_3020);
or U8555 (N_8555,N_4990,N_4521);
or U8556 (N_8556,N_1881,N_2496);
and U8557 (N_8557,N_462,N_3870);
xor U8558 (N_8558,N_1642,N_1862);
nand U8559 (N_8559,N_674,N_1397);
nand U8560 (N_8560,N_526,N_2262);
nor U8561 (N_8561,N_4539,N_1469);
and U8562 (N_8562,N_1150,N_2602);
nand U8563 (N_8563,N_4077,N_3575);
or U8564 (N_8564,N_2636,N_1130);
xor U8565 (N_8565,N_247,N_3363);
or U8566 (N_8566,N_812,N_690);
xnor U8567 (N_8567,N_4229,N_1903);
or U8568 (N_8568,N_2316,N_2712);
or U8569 (N_8569,N_3867,N_2308);
and U8570 (N_8570,N_737,N_4334);
nand U8571 (N_8571,N_3196,N_2561);
xor U8572 (N_8572,N_4596,N_1776);
xor U8573 (N_8573,N_3559,N_1771);
and U8574 (N_8574,N_1146,N_1630);
xnor U8575 (N_8575,N_2891,N_2111);
nand U8576 (N_8576,N_471,N_3429);
or U8577 (N_8577,N_1614,N_712);
nand U8578 (N_8578,N_3869,N_2036);
nor U8579 (N_8579,N_3964,N_1587);
nor U8580 (N_8580,N_2963,N_3839);
or U8581 (N_8581,N_3715,N_1593);
nand U8582 (N_8582,N_606,N_1083);
and U8583 (N_8583,N_345,N_119);
xnor U8584 (N_8584,N_4169,N_4638);
xnor U8585 (N_8585,N_3722,N_3260);
xor U8586 (N_8586,N_807,N_814);
nand U8587 (N_8587,N_2263,N_3566);
or U8588 (N_8588,N_4915,N_3353);
or U8589 (N_8589,N_2509,N_3383);
nor U8590 (N_8590,N_3191,N_2972);
xnor U8591 (N_8591,N_642,N_2569);
or U8592 (N_8592,N_4143,N_248);
nand U8593 (N_8593,N_3154,N_2817);
nor U8594 (N_8594,N_653,N_3104);
nor U8595 (N_8595,N_4174,N_4138);
or U8596 (N_8596,N_2965,N_1161);
or U8597 (N_8597,N_1234,N_3513);
nand U8598 (N_8598,N_4711,N_2161);
and U8599 (N_8599,N_1544,N_1653);
xor U8600 (N_8600,N_1601,N_395);
xor U8601 (N_8601,N_1169,N_865);
xnor U8602 (N_8602,N_2551,N_1076);
nand U8603 (N_8603,N_1817,N_765);
nor U8604 (N_8604,N_363,N_3455);
or U8605 (N_8605,N_4024,N_2995);
and U8606 (N_8606,N_3383,N_1376);
nor U8607 (N_8607,N_1664,N_3281);
nand U8608 (N_8608,N_1687,N_4318);
and U8609 (N_8609,N_2132,N_4017);
and U8610 (N_8610,N_1802,N_3658);
xnor U8611 (N_8611,N_2982,N_1013);
and U8612 (N_8612,N_2867,N_1266);
or U8613 (N_8613,N_2490,N_471);
and U8614 (N_8614,N_2741,N_1504);
nand U8615 (N_8615,N_4307,N_1900);
and U8616 (N_8616,N_1401,N_4693);
nand U8617 (N_8617,N_547,N_1272);
or U8618 (N_8618,N_1497,N_869);
xnor U8619 (N_8619,N_1929,N_1540);
nor U8620 (N_8620,N_3420,N_4029);
and U8621 (N_8621,N_2413,N_4211);
xor U8622 (N_8622,N_3001,N_4825);
xor U8623 (N_8623,N_641,N_1614);
and U8624 (N_8624,N_4271,N_3618);
nor U8625 (N_8625,N_2494,N_4612);
nor U8626 (N_8626,N_3913,N_4363);
or U8627 (N_8627,N_2485,N_1977);
and U8628 (N_8628,N_3566,N_985);
nand U8629 (N_8629,N_3960,N_3140);
nor U8630 (N_8630,N_160,N_596);
nand U8631 (N_8631,N_4952,N_544);
or U8632 (N_8632,N_1613,N_2329);
xnor U8633 (N_8633,N_1789,N_4987);
or U8634 (N_8634,N_1412,N_1966);
xnor U8635 (N_8635,N_2308,N_1336);
xor U8636 (N_8636,N_3199,N_4714);
and U8637 (N_8637,N_3172,N_594);
or U8638 (N_8638,N_3466,N_3862);
and U8639 (N_8639,N_2715,N_384);
nor U8640 (N_8640,N_4457,N_1502);
nor U8641 (N_8641,N_3764,N_2300);
nor U8642 (N_8642,N_1289,N_2739);
nor U8643 (N_8643,N_233,N_3801);
nand U8644 (N_8644,N_1358,N_3571);
or U8645 (N_8645,N_1793,N_4521);
nand U8646 (N_8646,N_4321,N_3831);
xor U8647 (N_8647,N_2962,N_4591);
and U8648 (N_8648,N_1085,N_4088);
nor U8649 (N_8649,N_3048,N_3296);
xnor U8650 (N_8650,N_4014,N_1757);
nand U8651 (N_8651,N_1253,N_4785);
and U8652 (N_8652,N_813,N_4785);
nor U8653 (N_8653,N_2843,N_1338);
xor U8654 (N_8654,N_4433,N_3563);
nor U8655 (N_8655,N_4924,N_822);
nand U8656 (N_8656,N_3876,N_3310);
and U8657 (N_8657,N_370,N_2402);
nand U8658 (N_8658,N_3973,N_4089);
xor U8659 (N_8659,N_4351,N_3753);
nand U8660 (N_8660,N_1565,N_3047);
or U8661 (N_8661,N_1404,N_136);
nor U8662 (N_8662,N_3661,N_2352);
and U8663 (N_8663,N_207,N_1136);
nor U8664 (N_8664,N_4668,N_3118);
and U8665 (N_8665,N_459,N_931);
or U8666 (N_8666,N_3052,N_3351);
or U8667 (N_8667,N_751,N_4436);
xor U8668 (N_8668,N_1478,N_6);
nor U8669 (N_8669,N_2387,N_4920);
xor U8670 (N_8670,N_316,N_3499);
and U8671 (N_8671,N_86,N_880);
or U8672 (N_8672,N_1622,N_4295);
or U8673 (N_8673,N_4273,N_4297);
xor U8674 (N_8674,N_3077,N_3135);
nand U8675 (N_8675,N_1761,N_2082);
nand U8676 (N_8676,N_864,N_1641);
nor U8677 (N_8677,N_4904,N_4605);
and U8678 (N_8678,N_1954,N_4797);
nand U8679 (N_8679,N_4908,N_2238);
or U8680 (N_8680,N_440,N_4147);
or U8681 (N_8681,N_3101,N_4546);
nor U8682 (N_8682,N_4861,N_2253);
xor U8683 (N_8683,N_2553,N_1009);
or U8684 (N_8684,N_1817,N_1902);
nor U8685 (N_8685,N_1994,N_2350);
and U8686 (N_8686,N_4756,N_186);
nor U8687 (N_8687,N_404,N_681);
or U8688 (N_8688,N_2363,N_3028);
or U8689 (N_8689,N_3734,N_2805);
xnor U8690 (N_8690,N_1506,N_1689);
nor U8691 (N_8691,N_2791,N_449);
and U8692 (N_8692,N_906,N_588);
nand U8693 (N_8693,N_72,N_199);
or U8694 (N_8694,N_3277,N_2606);
and U8695 (N_8695,N_1774,N_3752);
nor U8696 (N_8696,N_1927,N_2357);
or U8697 (N_8697,N_3481,N_3496);
xor U8698 (N_8698,N_4920,N_3396);
and U8699 (N_8699,N_4761,N_3838);
nand U8700 (N_8700,N_3246,N_2849);
nand U8701 (N_8701,N_1814,N_4901);
nand U8702 (N_8702,N_4137,N_3619);
and U8703 (N_8703,N_2654,N_3136);
nand U8704 (N_8704,N_3798,N_3849);
nand U8705 (N_8705,N_580,N_1053);
nand U8706 (N_8706,N_3212,N_557);
nor U8707 (N_8707,N_2790,N_2616);
and U8708 (N_8708,N_1207,N_3262);
and U8709 (N_8709,N_87,N_585);
or U8710 (N_8710,N_270,N_131);
nor U8711 (N_8711,N_226,N_2196);
or U8712 (N_8712,N_522,N_1885);
nand U8713 (N_8713,N_2343,N_793);
or U8714 (N_8714,N_722,N_2799);
and U8715 (N_8715,N_3364,N_523);
or U8716 (N_8716,N_4825,N_1209);
nand U8717 (N_8717,N_1051,N_480);
or U8718 (N_8718,N_3950,N_4154);
and U8719 (N_8719,N_2454,N_4472);
nor U8720 (N_8720,N_422,N_3935);
xor U8721 (N_8721,N_2126,N_3249);
xor U8722 (N_8722,N_3696,N_2166);
nor U8723 (N_8723,N_726,N_857);
nor U8724 (N_8724,N_4369,N_3309);
xor U8725 (N_8725,N_2141,N_2682);
and U8726 (N_8726,N_4986,N_2903);
nor U8727 (N_8727,N_1871,N_1509);
nand U8728 (N_8728,N_3787,N_4656);
nor U8729 (N_8729,N_1287,N_317);
xor U8730 (N_8730,N_3646,N_3632);
or U8731 (N_8731,N_2223,N_2422);
nor U8732 (N_8732,N_3172,N_3944);
and U8733 (N_8733,N_1147,N_3284);
and U8734 (N_8734,N_4961,N_4);
or U8735 (N_8735,N_750,N_1037);
and U8736 (N_8736,N_4042,N_2370);
xnor U8737 (N_8737,N_1712,N_2232);
nand U8738 (N_8738,N_3127,N_126);
nor U8739 (N_8739,N_4371,N_4437);
or U8740 (N_8740,N_1959,N_4086);
nor U8741 (N_8741,N_634,N_3227);
or U8742 (N_8742,N_1237,N_2329);
nor U8743 (N_8743,N_3270,N_3358);
xor U8744 (N_8744,N_1980,N_2379);
xnor U8745 (N_8745,N_4847,N_2219);
or U8746 (N_8746,N_3587,N_1663);
nor U8747 (N_8747,N_215,N_3522);
nor U8748 (N_8748,N_1000,N_3175);
and U8749 (N_8749,N_2446,N_822);
and U8750 (N_8750,N_2330,N_3892);
nand U8751 (N_8751,N_61,N_723);
nor U8752 (N_8752,N_3931,N_424);
or U8753 (N_8753,N_1315,N_3747);
nor U8754 (N_8754,N_2616,N_2158);
nor U8755 (N_8755,N_2903,N_3200);
xor U8756 (N_8756,N_4408,N_1996);
nor U8757 (N_8757,N_1180,N_2685);
or U8758 (N_8758,N_4900,N_4527);
xnor U8759 (N_8759,N_2966,N_460);
nor U8760 (N_8760,N_1507,N_3342);
and U8761 (N_8761,N_2206,N_2326);
nor U8762 (N_8762,N_4036,N_757);
nand U8763 (N_8763,N_826,N_3824);
nand U8764 (N_8764,N_3396,N_26);
and U8765 (N_8765,N_243,N_4976);
or U8766 (N_8766,N_717,N_3910);
or U8767 (N_8767,N_473,N_2081);
and U8768 (N_8768,N_19,N_4869);
nand U8769 (N_8769,N_200,N_1429);
and U8770 (N_8770,N_391,N_4657);
or U8771 (N_8771,N_3517,N_3294);
nor U8772 (N_8772,N_4148,N_3192);
nor U8773 (N_8773,N_4037,N_2994);
xnor U8774 (N_8774,N_395,N_2522);
and U8775 (N_8775,N_941,N_885);
or U8776 (N_8776,N_4435,N_35);
nor U8777 (N_8777,N_1452,N_3596);
xor U8778 (N_8778,N_367,N_2490);
xor U8779 (N_8779,N_155,N_3217);
xnor U8780 (N_8780,N_3125,N_1273);
or U8781 (N_8781,N_2215,N_2437);
nand U8782 (N_8782,N_959,N_3089);
or U8783 (N_8783,N_4094,N_2790);
or U8784 (N_8784,N_3166,N_134);
nand U8785 (N_8785,N_4855,N_4538);
nor U8786 (N_8786,N_3669,N_2527);
and U8787 (N_8787,N_183,N_882);
or U8788 (N_8788,N_4888,N_2009);
and U8789 (N_8789,N_2543,N_4495);
or U8790 (N_8790,N_1880,N_4829);
and U8791 (N_8791,N_3284,N_3292);
nor U8792 (N_8792,N_2000,N_3174);
nor U8793 (N_8793,N_2776,N_1264);
nand U8794 (N_8794,N_2067,N_3907);
nor U8795 (N_8795,N_3380,N_4686);
nor U8796 (N_8796,N_2846,N_2697);
nand U8797 (N_8797,N_3398,N_4642);
nor U8798 (N_8798,N_3770,N_4494);
and U8799 (N_8799,N_3479,N_2521);
and U8800 (N_8800,N_1722,N_790);
nor U8801 (N_8801,N_3616,N_155);
and U8802 (N_8802,N_1541,N_4839);
xor U8803 (N_8803,N_1859,N_4291);
or U8804 (N_8804,N_2706,N_4374);
or U8805 (N_8805,N_163,N_4443);
and U8806 (N_8806,N_373,N_3766);
and U8807 (N_8807,N_3300,N_1596);
xnor U8808 (N_8808,N_3407,N_2931);
and U8809 (N_8809,N_1065,N_2159);
or U8810 (N_8810,N_358,N_2837);
or U8811 (N_8811,N_2944,N_1561);
nand U8812 (N_8812,N_4627,N_2670);
nor U8813 (N_8813,N_146,N_81);
and U8814 (N_8814,N_4533,N_2880);
or U8815 (N_8815,N_895,N_4177);
xor U8816 (N_8816,N_4180,N_2730);
and U8817 (N_8817,N_819,N_1234);
and U8818 (N_8818,N_2892,N_3900);
and U8819 (N_8819,N_3947,N_4928);
and U8820 (N_8820,N_3690,N_2825);
and U8821 (N_8821,N_2549,N_1073);
nand U8822 (N_8822,N_4316,N_4870);
or U8823 (N_8823,N_1235,N_2966);
and U8824 (N_8824,N_1500,N_1073);
nor U8825 (N_8825,N_3188,N_1800);
and U8826 (N_8826,N_1411,N_3276);
xnor U8827 (N_8827,N_4562,N_4457);
or U8828 (N_8828,N_3228,N_1737);
xnor U8829 (N_8829,N_122,N_3830);
nand U8830 (N_8830,N_453,N_3119);
nor U8831 (N_8831,N_1609,N_4732);
or U8832 (N_8832,N_4414,N_2916);
and U8833 (N_8833,N_2466,N_2356);
and U8834 (N_8834,N_4597,N_436);
xor U8835 (N_8835,N_364,N_4752);
nand U8836 (N_8836,N_2609,N_2104);
or U8837 (N_8837,N_1971,N_2815);
nand U8838 (N_8838,N_4133,N_964);
xor U8839 (N_8839,N_3975,N_4813);
or U8840 (N_8840,N_575,N_1284);
and U8841 (N_8841,N_512,N_899);
xnor U8842 (N_8842,N_3898,N_4896);
nand U8843 (N_8843,N_2669,N_3579);
nor U8844 (N_8844,N_4010,N_3762);
xor U8845 (N_8845,N_2787,N_1691);
or U8846 (N_8846,N_2279,N_4204);
or U8847 (N_8847,N_2035,N_2314);
nor U8848 (N_8848,N_2968,N_349);
and U8849 (N_8849,N_4820,N_3623);
xnor U8850 (N_8850,N_1248,N_2547);
nor U8851 (N_8851,N_41,N_2807);
xnor U8852 (N_8852,N_3037,N_30);
xor U8853 (N_8853,N_3666,N_1121);
nor U8854 (N_8854,N_2256,N_4279);
or U8855 (N_8855,N_515,N_3014);
nor U8856 (N_8856,N_139,N_1170);
or U8857 (N_8857,N_3133,N_4810);
nand U8858 (N_8858,N_3081,N_3617);
or U8859 (N_8859,N_1529,N_2259);
nand U8860 (N_8860,N_4524,N_2069);
nand U8861 (N_8861,N_2085,N_2399);
or U8862 (N_8862,N_1073,N_1498);
nand U8863 (N_8863,N_3753,N_61);
xnor U8864 (N_8864,N_2516,N_562);
nor U8865 (N_8865,N_4344,N_157);
and U8866 (N_8866,N_869,N_4974);
and U8867 (N_8867,N_1409,N_2854);
xnor U8868 (N_8868,N_157,N_856);
nor U8869 (N_8869,N_3715,N_116);
nor U8870 (N_8870,N_4654,N_186);
and U8871 (N_8871,N_1100,N_2255);
or U8872 (N_8872,N_467,N_2808);
and U8873 (N_8873,N_4806,N_4608);
nor U8874 (N_8874,N_2527,N_4105);
xnor U8875 (N_8875,N_4734,N_2478);
xnor U8876 (N_8876,N_2602,N_1516);
xnor U8877 (N_8877,N_109,N_2775);
and U8878 (N_8878,N_3680,N_3560);
nor U8879 (N_8879,N_1048,N_1501);
and U8880 (N_8880,N_1107,N_4948);
nor U8881 (N_8881,N_3476,N_1984);
nand U8882 (N_8882,N_686,N_940);
xnor U8883 (N_8883,N_2217,N_4249);
nand U8884 (N_8884,N_3574,N_4436);
and U8885 (N_8885,N_1674,N_3245);
nand U8886 (N_8886,N_1734,N_2584);
nand U8887 (N_8887,N_1888,N_4350);
and U8888 (N_8888,N_4341,N_4543);
and U8889 (N_8889,N_4624,N_4077);
or U8890 (N_8890,N_2009,N_3022);
nand U8891 (N_8891,N_2420,N_505);
and U8892 (N_8892,N_2117,N_614);
xor U8893 (N_8893,N_4742,N_1320);
or U8894 (N_8894,N_2348,N_2685);
nand U8895 (N_8895,N_111,N_1838);
or U8896 (N_8896,N_4398,N_4561);
nand U8897 (N_8897,N_3946,N_2690);
nand U8898 (N_8898,N_3863,N_2772);
nand U8899 (N_8899,N_3953,N_152);
or U8900 (N_8900,N_1538,N_2006);
xnor U8901 (N_8901,N_383,N_843);
nand U8902 (N_8902,N_3304,N_2743);
nand U8903 (N_8903,N_3971,N_4904);
and U8904 (N_8904,N_1710,N_1307);
or U8905 (N_8905,N_4175,N_3630);
or U8906 (N_8906,N_4124,N_4076);
nor U8907 (N_8907,N_3588,N_1505);
nor U8908 (N_8908,N_2238,N_33);
or U8909 (N_8909,N_4694,N_1554);
nor U8910 (N_8910,N_4809,N_4377);
xor U8911 (N_8911,N_115,N_844);
nor U8912 (N_8912,N_245,N_129);
or U8913 (N_8913,N_516,N_393);
nor U8914 (N_8914,N_990,N_1756);
and U8915 (N_8915,N_2927,N_1762);
or U8916 (N_8916,N_401,N_4483);
and U8917 (N_8917,N_3429,N_2001);
xor U8918 (N_8918,N_3465,N_4094);
or U8919 (N_8919,N_248,N_3322);
nand U8920 (N_8920,N_833,N_1378);
nand U8921 (N_8921,N_4506,N_3494);
nand U8922 (N_8922,N_1025,N_2629);
nor U8923 (N_8923,N_3492,N_3723);
or U8924 (N_8924,N_4207,N_3782);
nor U8925 (N_8925,N_4562,N_4887);
or U8926 (N_8926,N_3097,N_73);
nand U8927 (N_8927,N_1073,N_2901);
nor U8928 (N_8928,N_4972,N_2431);
nand U8929 (N_8929,N_3492,N_120);
or U8930 (N_8930,N_1063,N_4953);
nor U8931 (N_8931,N_1146,N_785);
xnor U8932 (N_8932,N_2592,N_645);
nor U8933 (N_8933,N_411,N_1856);
nor U8934 (N_8934,N_3956,N_3253);
or U8935 (N_8935,N_1286,N_2951);
or U8936 (N_8936,N_956,N_4569);
or U8937 (N_8937,N_314,N_2428);
nand U8938 (N_8938,N_1492,N_35);
nand U8939 (N_8939,N_2291,N_4322);
nand U8940 (N_8940,N_1721,N_4763);
xnor U8941 (N_8941,N_3110,N_1894);
and U8942 (N_8942,N_1872,N_2931);
and U8943 (N_8943,N_2966,N_2909);
xor U8944 (N_8944,N_1425,N_4788);
or U8945 (N_8945,N_2671,N_4520);
xor U8946 (N_8946,N_129,N_804);
xor U8947 (N_8947,N_611,N_1350);
and U8948 (N_8948,N_698,N_2663);
nor U8949 (N_8949,N_210,N_2759);
nor U8950 (N_8950,N_1081,N_899);
xor U8951 (N_8951,N_4867,N_1910);
xor U8952 (N_8952,N_4558,N_2677);
or U8953 (N_8953,N_2338,N_4317);
xor U8954 (N_8954,N_582,N_1782);
nor U8955 (N_8955,N_4441,N_3260);
or U8956 (N_8956,N_869,N_132);
nand U8957 (N_8957,N_2540,N_4690);
nor U8958 (N_8958,N_4739,N_810);
nor U8959 (N_8959,N_1338,N_83);
nor U8960 (N_8960,N_1476,N_4987);
nand U8961 (N_8961,N_4924,N_4437);
nand U8962 (N_8962,N_720,N_186);
and U8963 (N_8963,N_2339,N_3125);
or U8964 (N_8964,N_4796,N_387);
and U8965 (N_8965,N_1940,N_3119);
nor U8966 (N_8966,N_4995,N_3337);
and U8967 (N_8967,N_4935,N_337);
and U8968 (N_8968,N_753,N_4377);
and U8969 (N_8969,N_4924,N_3683);
or U8970 (N_8970,N_4777,N_974);
xor U8971 (N_8971,N_3591,N_4206);
or U8972 (N_8972,N_3597,N_4711);
xnor U8973 (N_8973,N_4632,N_2081);
or U8974 (N_8974,N_1836,N_1408);
nor U8975 (N_8975,N_3709,N_2130);
nand U8976 (N_8976,N_2404,N_4973);
or U8977 (N_8977,N_1700,N_3091);
nor U8978 (N_8978,N_4505,N_3531);
nand U8979 (N_8979,N_4068,N_2344);
and U8980 (N_8980,N_2124,N_1457);
or U8981 (N_8981,N_352,N_3819);
nand U8982 (N_8982,N_968,N_3016);
nor U8983 (N_8983,N_48,N_208);
and U8984 (N_8984,N_2267,N_2386);
xnor U8985 (N_8985,N_4979,N_1935);
or U8986 (N_8986,N_3001,N_4706);
nand U8987 (N_8987,N_1696,N_3122);
xnor U8988 (N_8988,N_2516,N_2466);
or U8989 (N_8989,N_1500,N_4222);
and U8990 (N_8990,N_2608,N_3852);
nor U8991 (N_8991,N_2852,N_4955);
and U8992 (N_8992,N_4148,N_1476);
nand U8993 (N_8993,N_3172,N_2938);
xor U8994 (N_8994,N_4040,N_3612);
and U8995 (N_8995,N_923,N_4317);
or U8996 (N_8996,N_1356,N_3781);
nor U8997 (N_8997,N_1304,N_2006);
or U8998 (N_8998,N_4864,N_1184);
nor U8999 (N_8999,N_1815,N_3484);
nor U9000 (N_9000,N_3990,N_4508);
and U9001 (N_9001,N_1483,N_1727);
nand U9002 (N_9002,N_2326,N_2933);
and U9003 (N_9003,N_3401,N_2825);
nand U9004 (N_9004,N_1445,N_2094);
nor U9005 (N_9005,N_3593,N_1274);
or U9006 (N_9006,N_3018,N_3016);
xor U9007 (N_9007,N_649,N_2005);
nor U9008 (N_9008,N_2906,N_2586);
nand U9009 (N_9009,N_1365,N_4881);
and U9010 (N_9010,N_2769,N_403);
nand U9011 (N_9011,N_1292,N_4089);
nand U9012 (N_9012,N_4,N_2498);
and U9013 (N_9013,N_2988,N_2144);
or U9014 (N_9014,N_861,N_2529);
nor U9015 (N_9015,N_1833,N_3332);
or U9016 (N_9016,N_1714,N_785);
and U9017 (N_9017,N_3987,N_3439);
or U9018 (N_9018,N_2148,N_3104);
and U9019 (N_9019,N_4355,N_77);
or U9020 (N_9020,N_3580,N_3980);
nor U9021 (N_9021,N_302,N_78);
xnor U9022 (N_9022,N_3566,N_3323);
or U9023 (N_9023,N_643,N_868);
nor U9024 (N_9024,N_1949,N_121);
xor U9025 (N_9025,N_2173,N_4304);
xor U9026 (N_9026,N_203,N_1450);
nand U9027 (N_9027,N_4118,N_1897);
xor U9028 (N_9028,N_2192,N_4532);
nor U9029 (N_9029,N_4983,N_1942);
and U9030 (N_9030,N_2069,N_3795);
and U9031 (N_9031,N_4374,N_1496);
nor U9032 (N_9032,N_1576,N_535);
xor U9033 (N_9033,N_3507,N_1742);
nor U9034 (N_9034,N_2177,N_2929);
nor U9035 (N_9035,N_4801,N_2607);
nand U9036 (N_9036,N_3784,N_2861);
xor U9037 (N_9037,N_2884,N_811);
and U9038 (N_9038,N_1769,N_1705);
xor U9039 (N_9039,N_663,N_1670);
nor U9040 (N_9040,N_4548,N_2388);
xnor U9041 (N_9041,N_4744,N_2247);
nand U9042 (N_9042,N_2603,N_3352);
nand U9043 (N_9043,N_4851,N_4057);
or U9044 (N_9044,N_782,N_3310);
and U9045 (N_9045,N_2366,N_1181);
or U9046 (N_9046,N_1268,N_2778);
nand U9047 (N_9047,N_4389,N_4511);
nand U9048 (N_9048,N_4839,N_690);
xnor U9049 (N_9049,N_1452,N_1752);
and U9050 (N_9050,N_4687,N_2611);
or U9051 (N_9051,N_4135,N_2144);
xnor U9052 (N_9052,N_1427,N_2313);
xor U9053 (N_9053,N_2634,N_521);
xor U9054 (N_9054,N_3781,N_2928);
xnor U9055 (N_9055,N_4828,N_4666);
nor U9056 (N_9056,N_1967,N_176);
nor U9057 (N_9057,N_589,N_4133);
and U9058 (N_9058,N_2815,N_3898);
nor U9059 (N_9059,N_1657,N_2565);
and U9060 (N_9060,N_916,N_1244);
nor U9061 (N_9061,N_4811,N_2127);
nand U9062 (N_9062,N_316,N_4408);
nand U9063 (N_9063,N_3363,N_3043);
nor U9064 (N_9064,N_3704,N_3341);
nand U9065 (N_9065,N_3463,N_1232);
or U9066 (N_9066,N_3433,N_1523);
xor U9067 (N_9067,N_3461,N_1662);
nand U9068 (N_9068,N_3177,N_3599);
nand U9069 (N_9069,N_2034,N_3506);
xnor U9070 (N_9070,N_305,N_120);
and U9071 (N_9071,N_892,N_231);
or U9072 (N_9072,N_2688,N_562);
or U9073 (N_9073,N_2318,N_404);
nand U9074 (N_9074,N_4023,N_3984);
and U9075 (N_9075,N_1647,N_2277);
xnor U9076 (N_9076,N_3713,N_3581);
or U9077 (N_9077,N_2546,N_1789);
nor U9078 (N_9078,N_2875,N_395);
nand U9079 (N_9079,N_389,N_2713);
xnor U9080 (N_9080,N_1451,N_1289);
nand U9081 (N_9081,N_3516,N_1040);
and U9082 (N_9082,N_944,N_347);
xnor U9083 (N_9083,N_3364,N_2645);
xor U9084 (N_9084,N_104,N_737);
and U9085 (N_9085,N_2065,N_2155);
nand U9086 (N_9086,N_3015,N_1875);
or U9087 (N_9087,N_4411,N_3385);
or U9088 (N_9088,N_463,N_3146);
nand U9089 (N_9089,N_2282,N_937);
xnor U9090 (N_9090,N_3209,N_4028);
nand U9091 (N_9091,N_2277,N_3338);
nor U9092 (N_9092,N_2442,N_3695);
xnor U9093 (N_9093,N_3193,N_577);
nor U9094 (N_9094,N_4914,N_1751);
or U9095 (N_9095,N_1161,N_2052);
and U9096 (N_9096,N_1833,N_926);
nor U9097 (N_9097,N_858,N_4008);
or U9098 (N_9098,N_1164,N_4494);
and U9099 (N_9099,N_2665,N_743);
or U9100 (N_9100,N_2269,N_431);
nand U9101 (N_9101,N_2278,N_2901);
and U9102 (N_9102,N_2037,N_552);
xor U9103 (N_9103,N_1478,N_4563);
nand U9104 (N_9104,N_3556,N_1322);
or U9105 (N_9105,N_2651,N_4656);
and U9106 (N_9106,N_1563,N_185);
and U9107 (N_9107,N_679,N_322);
xnor U9108 (N_9108,N_1858,N_3078);
and U9109 (N_9109,N_1817,N_1389);
xnor U9110 (N_9110,N_1429,N_3195);
nand U9111 (N_9111,N_4726,N_1312);
nor U9112 (N_9112,N_438,N_1278);
and U9113 (N_9113,N_1067,N_25);
and U9114 (N_9114,N_3697,N_4310);
or U9115 (N_9115,N_46,N_2068);
and U9116 (N_9116,N_412,N_2956);
or U9117 (N_9117,N_582,N_2354);
or U9118 (N_9118,N_4,N_3387);
nand U9119 (N_9119,N_4273,N_3787);
and U9120 (N_9120,N_2061,N_4164);
nand U9121 (N_9121,N_2384,N_2490);
nor U9122 (N_9122,N_1844,N_4400);
nor U9123 (N_9123,N_4236,N_3143);
nand U9124 (N_9124,N_4360,N_2506);
or U9125 (N_9125,N_2148,N_4960);
nor U9126 (N_9126,N_4649,N_3516);
nand U9127 (N_9127,N_3549,N_3317);
or U9128 (N_9128,N_4018,N_789);
nand U9129 (N_9129,N_2897,N_519);
nand U9130 (N_9130,N_2555,N_1699);
and U9131 (N_9131,N_3250,N_3078);
xnor U9132 (N_9132,N_3225,N_2711);
xor U9133 (N_9133,N_3365,N_11);
or U9134 (N_9134,N_1415,N_3126);
xnor U9135 (N_9135,N_3358,N_4320);
nor U9136 (N_9136,N_2632,N_1252);
or U9137 (N_9137,N_703,N_509);
or U9138 (N_9138,N_4617,N_56);
and U9139 (N_9139,N_3687,N_1909);
and U9140 (N_9140,N_1067,N_3450);
and U9141 (N_9141,N_4608,N_2323);
nand U9142 (N_9142,N_2967,N_2308);
nor U9143 (N_9143,N_2953,N_2393);
xor U9144 (N_9144,N_1066,N_4837);
and U9145 (N_9145,N_3726,N_3898);
or U9146 (N_9146,N_4435,N_3164);
and U9147 (N_9147,N_726,N_447);
nor U9148 (N_9148,N_429,N_1811);
and U9149 (N_9149,N_1349,N_3401);
or U9150 (N_9150,N_2292,N_3186);
nand U9151 (N_9151,N_710,N_3809);
and U9152 (N_9152,N_1972,N_2090);
xor U9153 (N_9153,N_4997,N_452);
and U9154 (N_9154,N_3437,N_2442);
nor U9155 (N_9155,N_1330,N_2127);
nor U9156 (N_9156,N_59,N_1792);
or U9157 (N_9157,N_4406,N_1735);
or U9158 (N_9158,N_2412,N_4682);
and U9159 (N_9159,N_4513,N_4300);
and U9160 (N_9160,N_2767,N_1135);
xnor U9161 (N_9161,N_4926,N_2570);
and U9162 (N_9162,N_1055,N_3729);
and U9163 (N_9163,N_402,N_737);
xor U9164 (N_9164,N_2840,N_3725);
xor U9165 (N_9165,N_1233,N_3723);
xor U9166 (N_9166,N_632,N_857);
nor U9167 (N_9167,N_1980,N_1454);
nor U9168 (N_9168,N_671,N_8);
and U9169 (N_9169,N_4759,N_354);
nand U9170 (N_9170,N_3839,N_901);
nand U9171 (N_9171,N_1451,N_1395);
xnor U9172 (N_9172,N_4829,N_64);
xor U9173 (N_9173,N_443,N_3040);
or U9174 (N_9174,N_4046,N_2783);
nor U9175 (N_9175,N_946,N_3730);
or U9176 (N_9176,N_3918,N_2644);
or U9177 (N_9177,N_3249,N_776);
nand U9178 (N_9178,N_47,N_4553);
xor U9179 (N_9179,N_1919,N_3811);
nand U9180 (N_9180,N_1037,N_1687);
nor U9181 (N_9181,N_4176,N_669);
or U9182 (N_9182,N_3038,N_941);
xor U9183 (N_9183,N_1345,N_254);
nor U9184 (N_9184,N_1487,N_4794);
nand U9185 (N_9185,N_2523,N_2602);
or U9186 (N_9186,N_46,N_649);
and U9187 (N_9187,N_4051,N_2175);
or U9188 (N_9188,N_4730,N_2726);
nand U9189 (N_9189,N_158,N_4286);
nor U9190 (N_9190,N_4741,N_1291);
xor U9191 (N_9191,N_2542,N_2830);
nor U9192 (N_9192,N_1122,N_2081);
or U9193 (N_9193,N_4215,N_3081);
nand U9194 (N_9194,N_4408,N_3441);
xnor U9195 (N_9195,N_1718,N_889);
nand U9196 (N_9196,N_4089,N_4420);
and U9197 (N_9197,N_521,N_3467);
nand U9198 (N_9198,N_4865,N_1797);
or U9199 (N_9199,N_690,N_2250);
nor U9200 (N_9200,N_4529,N_4018);
nor U9201 (N_9201,N_4482,N_1124);
and U9202 (N_9202,N_57,N_4287);
or U9203 (N_9203,N_3420,N_271);
nor U9204 (N_9204,N_14,N_1704);
nand U9205 (N_9205,N_2745,N_4217);
or U9206 (N_9206,N_2266,N_2534);
or U9207 (N_9207,N_1392,N_1641);
and U9208 (N_9208,N_320,N_4192);
or U9209 (N_9209,N_1419,N_793);
nor U9210 (N_9210,N_3420,N_3037);
nand U9211 (N_9211,N_2072,N_2192);
nand U9212 (N_9212,N_927,N_1820);
and U9213 (N_9213,N_2182,N_3304);
and U9214 (N_9214,N_1396,N_4659);
nor U9215 (N_9215,N_2161,N_2348);
or U9216 (N_9216,N_405,N_2370);
and U9217 (N_9217,N_2163,N_355);
nand U9218 (N_9218,N_1625,N_1782);
or U9219 (N_9219,N_72,N_3039);
xnor U9220 (N_9220,N_4728,N_637);
xor U9221 (N_9221,N_3674,N_1603);
nor U9222 (N_9222,N_3508,N_1473);
nand U9223 (N_9223,N_4885,N_2533);
xnor U9224 (N_9224,N_2844,N_2242);
or U9225 (N_9225,N_2703,N_120);
or U9226 (N_9226,N_1578,N_56);
nand U9227 (N_9227,N_565,N_1565);
or U9228 (N_9228,N_3900,N_3293);
xor U9229 (N_9229,N_355,N_4409);
xnor U9230 (N_9230,N_1904,N_4466);
xor U9231 (N_9231,N_3989,N_3229);
or U9232 (N_9232,N_1159,N_3902);
xor U9233 (N_9233,N_1770,N_550);
xor U9234 (N_9234,N_2925,N_4490);
nor U9235 (N_9235,N_2167,N_4692);
xnor U9236 (N_9236,N_2811,N_4078);
xor U9237 (N_9237,N_4610,N_2514);
or U9238 (N_9238,N_1144,N_1427);
xnor U9239 (N_9239,N_3938,N_2674);
nand U9240 (N_9240,N_2817,N_2480);
and U9241 (N_9241,N_2252,N_4222);
and U9242 (N_9242,N_2688,N_4564);
xor U9243 (N_9243,N_3404,N_3059);
nand U9244 (N_9244,N_489,N_4399);
nor U9245 (N_9245,N_3065,N_1888);
xnor U9246 (N_9246,N_3031,N_4171);
nand U9247 (N_9247,N_1662,N_1370);
nand U9248 (N_9248,N_4062,N_4085);
nor U9249 (N_9249,N_3928,N_4069);
xor U9250 (N_9250,N_4264,N_2753);
or U9251 (N_9251,N_741,N_4694);
xnor U9252 (N_9252,N_1332,N_3618);
nand U9253 (N_9253,N_3129,N_1550);
or U9254 (N_9254,N_64,N_2676);
nor U9255 (N_9255,N_3060,N_4274);
or U9256 (N_9256,N_3209,N_3411);
nand U9257 (N_9257,N_846,N_2678);
and U9258 (N_9258,N_960,N_4212);
nand U9259 (N_9259,N_4900,N_2853);
or U9260 (N_9260,N_2000,N_2475);
or U9261 (N_9261,N_2761,N_3606);
nand U9262 (N_9262,N_2484,N_4077);
nand U9263 (N_9263,N_4658,N_2814);
or U9264 (N_9264,N_3658,N_189);
or U9265 (N_9265,N_2493,N_4276);
xor U9266 (N_9266,N_660,N_4622);
nor U9267 (N_9267,N_4405,N_1077);
or U9268 (N_9268,N_4613,N_4001);
and U9269 (N_9269,N_2802,N_922);
nor U9270 (N_9270,N_2463,N_3239);
nand U9271 (N_9271,N_3688,N_2017);
xor U9272 (N_9272,N_3101,N_2736);
or U9273 (N_9273,N_1394,N_2943);
xor U9274 (N_9274,N_2120,N_4448);
and U9275 (N_9275,N_4187,N_1959);
xor U9276 (N_9276,N_2950,N_4940);
or U9277 (N_9277,N_2342,N_4865);
nand U9278 (N_9278,N_4836,N_3107);
xnor U9279 (N_9279,N_1695,N_2333);
nor U9280 (N_9280,N_308,N_2759);
and U9281 (N_9281,N_3594,N_4145);
nor U9282 (N_9282,N_4359,N_1600);
nand U9283 (N_9283,N_4464,N_1139);
or U9284 (N_9284,N_2435,N_4223);
or U9285 (N_9285,N_2606,N_4476);
nand U9286 (N_9286,N_4847,N_2741);
xnor U9287 (N_9287,N_2994,N_581);
nand U9288 (N_9288,N_3796,N_2622);
and U9289 (N_9289,N_707,N_2731);
xor U9290 (N_9290,N_3175,N_1217);
xor U9291 (N_9291,N_4071,N_2317);
or U9292 (N_9292,N_4840,N_2109);
nand U9293 (N_9293,N_4015,N_4179);
or U9294 (N_9294,N_131,N_940);
xnor U9295 (N_9295,N_815,N_3577);
nor U9296 (N_9296,N_3801,N_1896);
or U9297 (N_9297,N_3574,N_636);
nor U9298 (N_9298,N_4078,N_2459);
xor U9299 (N_9299,N_1310,N_195);
or U9300 (N_9300,N_370,N_1847);
xor U9301 (N_9301,N_3650,N_646);
xor U9302 (N_9302,N_2326,N_2892);
nand U9303 (N_9303,N_4711,N_4181);
or U9304 (N_9304,N_1314,N_785);
xnor U9305 (N_9305,N_1935,N_3272);
or U9306 (N_9306,N_448,N_3578);
nor U9307 (N_9307,N_1044,N_4525);
and U9308 (N_9308,N_1126,N_4894);
nor U9309 (N_9309,N_4810,N_3945);
xnor U9310 (N_9310,N_2314,N_2780);
nor U9311 (N_9311,N_1394,N_1250);
xor U9312 (N_9312,N_2741,N_1110);
and U9313 (N_9313,N_4464,N_3131);
or U9314 (N_9314,N_1823,N_4835);
nand U9315 (N_9315,N_460,N_3842);
or U9316 (N_9316,N_629,N_2447);
nor U9317 (N_9317,N_3625,N_934);
xnor U9318 (N_9318,N_1441,N_2215);
nand U9319 (N_9319,N_4795,N_1820);
and U9320 (N_9320,N_192,N_2622);
and U9321 (N_9321,N_1883,N_1779);
nor U9322 (N_9322,N_2696,N_1342);
nor U9323 (N_9323,N_3690,N_4468);
nor U9324 (N_9324,N_1366,N_4846);
nand U9325 (N_9325,N_4316,N_3348);
nand U9326 (N_9326,N_1365,N_2301);
nand U9327 (N_9327,N_3658,N_4333);
nor U9328 (N_9328,N_4135,N_1202);
xnor U9329 (N_9329,N_1623,N_1139);
nand U9330 (N_9330,N_4196,N_4780);
xnor U9331 (N_9331,N_551,N_2521);
and U9332 (N_9332,N_1058,N_3990);
and U9333 (N_9333,N_4308,N_1605);
and U9334 (N_9334,N_3190,N_3530);
nor U9335 (N_9335,N_2795,N_685);
nand U9336 (N_9336,N_4493,N_2900);
nand U9337 (N_9337,N_2528,N_2639);
nor U9338 (N_9338,N_3315,N_3312);
xor U9339 (N_9339,N_3626,N_2708);
or U9340 (N_9340,N_1388,N_3638);
or U9341 (N_9341,N_4940,N_2315);
and U9342 (N_9342,N_3714,N_2231);
and U9343 (N_9343,N_789,N_3166);
xnor U9344 (N_9344,N_279,N_908);
nand U9345 (N_9345,N_4135,N_3160);
nand U9346 (N_9346,N_3038,N_4891);
and U9347 (N_9347,N_1142,N_1557);
or U9348 (N_9348,N_3879,N_4431);
xnor U9349 (N_9349,N_1153,N_2198);
and U9350 (N_9350,N_2266,N_4786);
xnor U9351 (N_9351,N_1673,N_1802);
and U9352 (N_9352,N_3943,N_739);
and U9353 (N_9353,N_4287,N_2403);
xor U9354 (N_9354,N_202,N_3899);
nand U9355 (N_9355,N_4940,N_2379);
or U9356 (N_9356,N_3623,N_2481);
xnor U9357 (N_9357,N_3603,N_628);
xor U9358 (N_9358,N_1533,N_3830);
nor U9359 (N_9359,N_887,N_4140);
or U9360 (N_9360,N_4248,N_1681);
xor U9361 (N_9361,N_2145,N_4628);
nor U9362 (N_9362,N_3759,N_2347);
xor U9363 (N_9363,N_812,N_10);
xor U9364 (N_9364,N_4812,N_1916);
nand U9365 (N_9365,N_1491,N_2563);
xor U9366 (N_9366,N_4392,N_2975);
xnor U9367 (N_9367,N_3065,N_4335);
xor U9368 (N_9368,N_3239,N_2780);
or U9369 (N_9369,N_1567,N_3947);
nor U9370 (N_9370,N_2422,N_1866);
and U9371 (N_9371,N_3525,N_45);
nor U9372 (N_9372,N_4629,N_1034);
nand U9373 (N_9373,N_504,N_3057);
and U9374 (N_9374,N_3918,N_4965);
or U9375 (N_9375,N_462,N_3285);
xor U9376 (N_9376,N_3654,N_369);
nand U9377 (N_9377,N_1376,N_4553);
nand U9378 (N_9378,N_4615,N_2326);
xnor U9379 (N_9379,N_2553,N_2228);
nand U9380 (N_9380,N_2590,N_3912);
xor U9381 (N_9381,N_18,N_4838);
and U9382 (N_9382,N_3673,N_3200);
nor U9383 (N_9383,N_490,N_4836);
or U9384 (N_9384,N_2149,N_4624);
and U9385 (N_9385,N_779,N_3734);
and U9386 (N_9386,N_4461,N_1305);
nand U9387 (N_9387,N_3065,N_1134);
and U9388 (N_9388,N_1517,N_100);
or U9389 (N_9389,N_2294,N_3343);
nand U9390 (N_9390,N_262,N_2016);
and U9391 (N_9391,N_844,N_4674);
nand U9392 (N_9392,N_3775,N_4198);
nand U9393 (N_9393,N_1231,N_623);
xor U9394 (N_9394,N_2136,N_3113);
and U9395 (N_9395,N_519,N_2325);
xor U9396 (N_9396,N_3668,N_3111);
or U9397 (N_9397,N_1971,N_1236);
xnor U9398 (N_9398,N_2473,N_1968);
or U9399 (N_9399,N_2665,N_1606);
or U9400 (N_9400,N_3155,N_1236);
and U9401 (N_9401,N_3778,N_1142);
and U9402 (N_9402,N_1883,N_4539);
or U9403 (N_9403,N_3490,N_4446);
xnor U9404 (N_9404,N_1269,N_4803);
and U9405 (N_9405,N_3216,N_4848);
or U9406 (N_9406,N_1418,N_1512);
or U9407 (N_9407,N_3496,N_2213);
or U9408 (N_9408,N_2519,N_1242);
and U9409 (N_9409,N_75,N_2275);
xnor U9410 (N_9410,N_4040,N_1807);
or U9411 (N_9411,N_3298,N_3427);
xnor U9412 (N_9412,N_926,N_2719);
xor U9413 (N_9413,N_3163,N_3776);
nand U9414 (N_9414,N_782,N_3112);
xnor U9415 (N_9415,N_2519,N_3473);
and U9416 (N_9416,N_3720,N_665);
nor U9417 (N_9417,N_603,N_363);
xor U9418 (N_9418,N_3060,N_1743);
nor U9419 (N_9419,N_4612,N_578);
nand U9420 (N_9420,N_2146,N_383);
nand U9421 (N_9421,N_1806,N_2365);
xor U9422 (N_9422,N_3155,N_3044);
or U9423 (N_9423,N_3213,N_4125);
nand U9424 (N_9424,N_2118,N_3078);
nor U9425 (N_9425,N_273,N_2907);
or U9426 (N_9426,N_2868,N_1839);
and U9427 (N_9427,N_4305,N_2920);
and U9428 (N_9428,N_1948,N_4279);
or U9429 (N_9429,N_1985,N_1051);
xor U9430 (N_9430,N_899,N_3727);
nor U9431 (N_9431,N_2285,N_771);
and U9432 (N_9432,N_2319,N_4899);
nand U9433 (N_9433,N_166,N_2236);
nand U9434 (N_9434,N_741,N_1735);
nand U9435 (N_9435,N_3690,N_3054);
nor U9436 (N_9436,N_2079,N_3172);
nor U9437 (N_9437,N_3999,N_1842);
and U9438 (N_9438,N_4349,N_3329);
or U9439 (N_9439,N_4228,N_2842);
and U9440 (N_9440,N_314,N_3768);
nor U9441 (N_9441,N_2524,N_2311);
and U9442 (N_9442,N_1430,N_3209);
nand U9443 (N_9443,N_1147,N_3087);
nor U9444 (N_9444,N_2269,N_236);
nor U9445 (N_9445,N_1332,N_3636);
or U9446 (N_9446,N_2245,N_1312);
xor U9447 (N_9447,N_4320,N_3539);
nor U9448 (N_9448,N_3807,N_4138);
and U9449 (N_9449,N_293,N_1086);
xor U9450 (N_9450,N_2659,N_1232);
and U9451 (N_9451,N_70,N_2981);
and U9452 (N_9452,N_4663,N_2459);
xnor U9453 (N_9453,N_1120,N_803);
and U9454 (N_9454,N_2285,N_3190);
nor U9455 (N_9455,N_2816,N_2252);
or U9456 (N_9456,N_1951,N_830);
xnor U9457 (N_9457,N_3775,N_3106);
nor U9458 (N_9458,N_1035,N_1730);
nand U9459 (N_9459,N_2343,N_1970);
xnor U9460 (N_9460,N_3992,N_404);
nand U9461 (N_9461,N_1049,N_393);
nand U9462 (N_9462,N_1633,N_4389);
and U9463 (N_9463,N_1208,N_26);
xnor U9464 (N_9464,N_3882,N_4253);
nor U9465 (N_9465,N_1305,N_4394);
nor U9466 (N_9466,N_2637,N_370);
nor U9467 (N_9467,N_3572,N_2850);
nand U9468 (N_9468,N_1137,N_3784);
and U9469 (N_9469,N_2268,N_2830);
nor U9470 (N_9470,N_1467,N_1062);
and U9471 (N_9471,N_2944,N_3921);
xor U9472 (N_9472,N_2447,N_2426);
nand U9473 (N_9473,N_3309,N_733);
nor U9474 (N_9474,N_4374,N_1434);
and U9475 (N_9475,N_1821,N_981);
and U9476 (N_9476,N_3650,N_3011);
nor U9477 (N_9477,N_596,N_3473);
nand U9478 (N_9478,N_740,N_4218);
nor U9479 (N_9479,N_243,N_3822);
and U9480 (N_9480,N_63,N_4660);
and U9481 (N_9481,N_589,N_3453);
xnor U9482 (N_9482,N_1898,N_519);
nand U9483 (N_9483,N_3878,N_2598);
nand U9484 (N_9484,N_3260,N_1656);
nor U9485 (N_9485,N_2206,N_4039);
and U9486 (N_9486,N_331,N_2841);
or U9487 (N_9487,N_4746,N_1939);
xnor U9488 (N_9488,N_575,N_4997);
nand U9489 (N_9489,N_1851,N_4440);
xor U9490 (N_9490,N_3280,N_1761);
or U9491 (N_9491,N_2865,N_1147);
or U9492 (N_9492,N_4790,N_4634);
or U9493 (N_9493,N_4199,N_2114);
nor U9494 (N_9494,N_763,N_4434);
nand U9495 (N_9495,N_2008,N_4569);
nor U9496 (N_9496,N_2905,N_888);
nand U9497 (N_9497,N_3149,N_343);
or U9498 (N_9498,N_2305,N_3651);
or U9499 (N_9499,N_3054,N_4502);
or U9500 (N_9500,N_1634,N_3838);
xnor U9501 (N_9501,N_1995,N_3726);
nor U9502 (N_9502,N_3792,N_2580);
or U9503 (N_9503,N_3908,N_3895);
nand U9504 (N_9504,N_3685,N_2992);
nor U9505 (N_9505,N_3302,N_1702);
nand U9506 (N_9506,N_1872,N_1526);
and U9507 (N_9507,N_1707,N_329);
or U9508 (N_9508,N_366,N_3070);
or U9509 (N_9509,N_2353,N_864);
nor U9510 (N_9510,N_3985,N_2687);
or U9511 (N_9511,N_1983,N_1869);
xnor U9512 (N_9512,N_1823,N_1252);
nor U9513 (N_9513,N_225,N_2099);
or U9514 (N_9514,N_1698,N_1633);
or U9515 (N_9515,N_177,N_4444);
xnor U9516 (N_9516,N_2917,N_513);
xnor U9517 (N_9517,N_694,N_382);
or U9518 (N_9518,N_3806,N_3727);
or U9519 (N_9519,N_278,N_3710);
nor U9520 (N_9520,N_3315,N_3150);
xor U9521 (N_9521,N_2828,N_3847);
nor U9522 (N_9522,N_602,N_3309);
and U9523 (N_9523,N_3886,N_867);
nor U9524 (N_9524,N_3748,N_3917);
or U9525 (N_9525,N_3037,N_2543);
or U9526 (N_9526,N_3580,N_3746);
nand U9527 (N_9527,N_403,N_959);
or U9528 (N_9528,N_4801,N_1827);
nand U9529 (N_9529,N_2226,N_1655);
nor U9530 (N_9530,N_3004,N_3521);
nand U9531 (N_9531,N_1957,N_1512);
and U9532 (N_9532,N_4146,N_949);
and U9533 (N_9533,N_2037,N_3265);
xnor U9534 (N_9534,N_1254,N_3153);
nand U9535 (N_9535,N_4361,N_1720);
nand U9536 (N_9536,N_809,N_3666);
xnor U9537 (N_9537,N_2166,N_2515);
and U9538 (N_9538,N_3102,N_1953);
nor U9539 (N_9539,N_2960,N_2151);
and U9540 (N_9540,N_3375,N_1679);
and U9541 (N_9541,N_1656,N_4806);
nor U9542 (N_9542,N_3717,N_1495);
and U9543 (N_9543,N_3019,N_1382);
or U9544 (N_9544,N_1457,N_4153);
and U9545 (N_9545,N_3676,N_3888);
nand U9546 (N_9546,N_2076,N_4557);
nor U9547 (N_9547,N_4493,N_4348);
or U9548 (N_9548,N_3152,N_3127);
xor U9549 (N_9549,N_2373,N_2218);
or U9550 (N_9550,N_3877,N_1020);
nand U9551 (N_9551,N_1237,N_2079);
nor U9552 (N_9552,N_1401,N_64);
or U9553 (N_9553,N_3651,N_227);
nand U9554 (N_9554,N_3295,N_1582);
or U9555 (N_9555,N_4612,N_4468);
or U9556 (N_9556,N_3660,N_2101);
nor U9557 (N_9557,N_4765,N_318);
or U9558 (N_9558,N_2207,N_1617);
nor U9559 (N_9559,N_4272,N_4685);
and U9560 (N_9560,N_1654,N_4849);
nand U9561 (N_9561,N_3216,N_1217);
nand U9562 (N_9562,N_1813,N_1377);
xor U9563 (N_9563,N_584,N_4766);
nand U9564 (N_9564,N_2148,N_2327);
nand U9565 (N_9565,N_1238,N_4260);
nand U9566 (N_9566,N_437,N_4778);
and U9567 (N_9567,N_163,N_3410);
and U9568 (N_9568,N_2471,N_1900);
nor U9569 (N_9569,N_879,N_4108);
nand U9570 (N_9570,N_688,N_2152);
xor U9571 (N_9571,N_62,N_3902);
xnor U9572 (N_9572,N_3229,N_1809);
or U9573 (N_9573,N_1960,N_2642);
xnor U9574 (N_9574,N_4159,N_305);
nand U9575 (N_9575,N_4109,N_1515);
or U9576 (N_9576,N_3629,N_1527);
nand U9577 (N_9577,N_1490,N_3785);
nor U9578 (N_9578,N_2672,N_3429);
nor U9579 (N_9579,N_1664,N_3524);
and U9580 (N_9580,N_4169,N_2101);
or U9581 (N_9581,N_3378,N_534);
or U9582 (N_9582,N_4939,N_1088);
or U9583 (N_9583,N_336,N_2700);
xor U9584 (N_9584,N_4244,N_4550);
nand U9585 (N_9585,N_4680,N_2977);
and U9586 (N_9586,N_333,N_3910);
xor U9587 (N_9587,N_2463,N_4906);
and U9588 (N_9588,N_465,N_3271);
or U9589 (N_9589,N_1214,N_4581);
and U9590 (N_9590,N_4881,N_4425);
nand U9591 (N_9591,N_3937,N_1491);
and U9592 (N_9592,N_1381,N_1779);
and U9593 (N_9593,N_1237,N_1225);
nand U9594 (N_9594,N_2819,N_3846);
xor U9595 (N_9595,N_3269,N_2866);
and U9596 (N_9596,N_3596,N_4935);
nand U9597 (N_9597,N_2897,N_3831);
or U9598 (N_9598,N_3307,N_3084);
nand U9599 (N_9599,N_1330,N_2788);
nor U9600 (N_9600,N_1268,N_3170);
nand U9601 (N_9601,N_4795,N_4525);
or U9602 (N_9602,N_3027,N_2798);
nor U9603 (N_9603,N_252,N_1355);
or U9604 (N_9604,N_880,N_1497);
or U9605 (N_9605,N_1242,N_1501);
and U9606 (N_9606,N_4461,N_3785);
and U9607 (N_9607,N_1332,N_2822);
nand U9608 (N_9608,N_3185,N_2462);
nor U9609 (N_9609,N_4215,N_2463);
nor U9610 (N_9610,N_3398,N_2058);
and U9611 (N_9611,N_3984,N_3295);
xor U9612 (N_9612,N_4507,N_2377);
nor U9613 (N_9613,N_2018,N_2403);
xnor U9614 (N_9614,N_1297,N_395);
xnor U9615 (N_9615,N_3023,N_1202);
and U9616 (N_9616,N_1341,N_3594);
nor U9617 (N_9617,N_2929,N_4687);
and U9618 (N_9618,N_3173,N_1935);
nand U9619 (N_9619,N_1318,N_2713);
and U9620 (N_9620,N_3915,N_2199);
nor U9621 (N_9621,N_4081,N_2653);
nand U9622 (N_9622,N_3111,N_2665);
and U9623 (N_9623,N_4184,N_3308);
nor U9624 (N_9624,N_3863,N_4910);
xnor U9625 (N_9625,N_4980,N_4082);
and U9626 (N_9626,N_1663,N_2885);
nand U9627 (N_9627,N_3869,N_403);
nor U9628 (N_9628,N_629,N_2397);
nor U9629 (N_9629,N_4337,N_2370);
or U9630 (N_9630,N_4255,N_2550);
nand U9631 (N_9631,N_106,N_1028);
nand U9632 (N_9632,N_3988,N_3485);
and U9633 (N_9633,N_4637,N_626);
nand U9634 (N_9634,N_2273,N_1965);
nand U9635 (N_9635,N_3971,N_4493);
nor U9636 (N_9636,N_1661,N_4939);
xor U9637 (N_9637,N_2464,N_3908);
nand U9638 (N_9638,N_40,N_1268);
nand U9639 (N_9639,N_2890,N_1991);
or U9640 (N_9640,N_942,N_4409);
and U9641 (N_9641,N_3755,N_2689);
xnor U9642 (N_9642,N_801,N_4387);
nor U9643 (N_9643,N_4380,N_1066);
nand U9644 (N_9644,N_1738,N_4483);
and U9645 (N_9645,N_723,N_3575);
xor U9646 (N_9646,N_1258,N_3735);
nor U9647 (N_9647,N_3737,N_3571);
nand U9648 (N_9648,N_4413,N_3322);
xnor U9649 (N_9649,N_1244,N_2047);
nand U9650 (N_9650,N_3515,N_1218);
nor U9651 (N_9651,N_2276,N_4945);
nor U9652 (N_9652,N_3650,N_3725);
nor U9653 (N_9653,N_1391,N_1937);
or U9654 (N_9654,N_2813,N_1330);
nor U9655 (N_9655,N_2088,N_4914);
xor U9656 (N_9656,N_2439,N_1386);
and U9657 (N_9657,N_2473,N_3198);
nor U9658 (N_9658,N_4464,N_2719);
nand U9659 (N_9659,N_1275,N_203);
and U9660 (N_9660,N_4816,N_2079);
xnor U9661 (N_9661,N_160,N_4319);
and U9662 (N_9662,N_2547,N_3608);
or U9663 (N_9663,N_2506,N_2438);
nor U9664 (N_9664,N_1413,N_715);
or U9665 (N_9665,N_3916,N_2043);
and U9666 (N_9666,N_590,N_2865);
nand U9667 (N_9667,N_1658,N_1564);
and U9668 (N_9668,N_3919,N_4967);
or U9669 (N_9669,N_52,N_956);
xor U9670 (N_9670,N_764,N_2548);
nand U9671 (N_9671,N_1610,N_2135);
xnor U9672 (N_9672,N_2366,N_1352);
and U9673 (N_9673,N_1114,N_2890);
or U9674 (N_9674,N_1426,N_3592);
nand U9675 (N_9675,N_154,N_3320);
or U9676 (N_9676,N_1383,N_3058);
nor U9677 (N_9677,N_960,N_779);
and U9678 (N_9678,N_3770,N_2068);
nand U9679 (N_9679,N_2263,N_345);
and U9680 (N_9680,N_1255,N_820);
and U9681 (N_9681,N_2260,N_2379);
nor U9682 (N_9682,N_3913,N_4545);
or U9683 (N_9683,N_3846,N_828);
xnor U9684 (N_9684,N_261,N_2953);
and U9685 (N_9685,N_3178,N_4518);
and U9686 (N_9686,N_3328,N_4019);
nor U9687 (N_9687,N_1802,N_3760);
and U9688 (N_9688,N_2851,N_3169);
or U9689 (N_9689,N_3393,N_2787);
xnor U9690 (N_9690,N_1861,N_2600);
xnor U9691 (N_9691,N_3697,N_2597);
or U9692 (N_9692,N_279,N_2008);
nor U9693 (N_9693,N_848,N_856);
xor U9694 (N_9694,N_1435,N_4533);
xor U9695 (N_9695,N_2200,N_3843);
xnor U9696 (N_9696,N_701,N_3274);
nand U9697 (N_9697,N_4681,N_1155);
nand U9698 (N_9698,N_2542,N_224);
nor U9699 (N_9699,N_3050,N_3536);
and U9700 (N_9700,N_4458,N_2889);
or U9701 (N_9701,N_516,N_1000);
or U9702 (N_9702,N_4326,N_2919);
or U9703 (N_9703,N_4095,N_4404);
xnor U9704 (N_9704,N_3098,N_3265);
nor U9705 (N_9705,N_185,N_1146);
or U9706 (N_9706,N_3238,N_4803);
nand U9707 (N_9707,N_4952,N_1134);
nor U9708 (N_9708,N_3182,N_1349);
xnor U9709 (N_9709,N_3999,N_2033);
xor U9710 (N_9710,N_4553,N_1915);
or U9711 (N_9711,N_122,N_1302);
nand U9712 (N_9712,N_1885,N_2016);
nor U9713 (N_9713,N_752,N_1629);
and U9714 (N_9714,N_4342,N_3594);
or U9715 (N_9715,N_2944,N_4458);
xnor U9716 (N_9716,N_4928,N_732);
or U9717 (N_9717,N_516,N_731);
and U9718 (N_9718,N_1440,N_3572);
xor U9719 (N_9719,N_3396,N_3902);
or U9720 (N_9720,N_1249,N_4096);
xor U9721 (N_9721,N_1653,N_4556);
or U9722 (N_9722,N_3155,N_1735);
nor U9723 (N_9723,N_127,N_3266);
and U9724 (N_9724,N_2718,N_4191);
xnor U9725 (N_9725,N_988,N_1446);
xnor U9726 (N_9726,N_809,N_1755);
xor U9727 (N_9727,N_2289,N_387);
nor U9728 (N_9728,N_4345,N_298);
or U9729 (N_9729,N_231,N_1820);
xnor U9730 (N_9730,N_3180,N_2342);
or U9731 (N_9731,N_1503,N_107);
nand U9732 (N_9732,N_2160,N_1918);
and U9733 (N_9733,N_3841,N_4043);
xnor U9734 (N_9734,N_1871,N_4611);
xnor U9735 (N_9735,N_2724,N_4533);
and U9736 (N_9736,N_245,N_4278);
or U9737 (N_9737,N_692,N_1245);
xnor U9738 (N_9738,N_2805,N_155);
or U9739 (N_9739,N_1241,N_4714);
nor U9740 (N_9740,N_3380,N_176);
nand U9741 (N_9741,N_2592,N_2687);
nand U9742 (N_9742,N_1050,N_4939);
nand U9743 (N_9743,N_4686,N_4360);
and U9744 (N_9744,N_4100,N_1312);
xnor U9745 (N_9745,N_1834,N_1556);
nand U9746 (N_9746,N_987,N_4205);
nor U9747 (N_9747,N_1343,N_4501);
nand U9748 (N_9748,N_4992,N_3160);
and U9749 (N_9749,N_4670,N_958);
xor U9750 (N_9750,N_3427,N_3462);
nand U9751 (N_9751,N_665,N_3248);
nor U9752 (N_9752,N_3305,N_4055);
nand U9753 (N_9753,N_1246,N_121);
xnor U9754 (N_9754,N_288,N_3115);
or U9755 (N_9755,N_2191,N_3591);
nor U9756 (N_9756,N_4481,N_2576);
or U9757 (N_9757,N_3600,N_3324);
nor U9758 (N_9758,N_4198,N_2894);
or U9759 (N_9759,N_62,N_2233);
nand U9760 (N_9760,N_3197,N_717);
nand U9761 (N_9761,N_1770,N_2816);
nand U9762 (N_9762,N_4953,N_2837);
or U9763 (N_9763,N_4414,N_330);
or U9764 (N_9764,N_4698,N_3156);
and U9765 (N_9765,N_2749,N_3698);
nor U9766 (N_9766,N_3096,N_3434);
xor U9767 (N_9767,N_4810,N_818);
or U9768 (N_9768,N_3081,N_1188);
xnor U9769 (N_9769,N_4001,N_2283);
xnor U9770 (N_9770,N_3816,N_157);
or U9771 (N_9771,N_1061,N_2351);
xnor U9772 (N_9772,N_1428,N_1336);
and U9773 (N_9773,N_3653,N_3496);
xnor U9774 (N_9774,N_3807,N_2851);
nand U9775 (N_9775,N_4826,N_285);
or U9776 (N_9776,N_4694,N_4282);
xor U9777 (N_9777,N_3615,N_325);
nor U9778 (N_9778,N_315,N_110);
or U9779 (N_9779,N_379,N_2301);
nor U9780 (N_9780,N_2884,N_1756);
nand U9781 (N_9781,N_2083,N_1347);
or U9782 (N_9782,N_4925,N_2916);
nor U9783 (N_9783,N_4820,N_4924);
nor U9784 (N_9784,N_2175,N_4023);
nor U9785 (N_9785,N_2496,N_2877);
nand U9786 (N_9786,N_3110,N_2778);
nand U9787 (N_9787,N_1833,N_3065);
or U9788 (N_9788,N_1690,N_2026);
and U9789 (N_9789,N_413,N_4996);
nor U9790 (N_9790,N_2047,N_1233);
nand U9791 (N_9791,N_279,N_4163);
nor U9792 (N_9792,N_3143,N_1935);
xnor U9793 (N_9793,N_1625,N_4469);
xnor U9794 (N_9794,N_683,N_3268);
nor U9795 (N_9795,N_1414,N_3386);
or U9796 (N_9796,N_83,N_4311);
nand U9797 (N_9797,N_160,N_4110);
xnor U9798 (N_9798,N_1908,N_2047);
nand U9799 (N_9799,N_2382,N_2586);
nand U9800 (N_9800,N_229,N_3542);
and U9801 (N_9801,N_2048,N_3056);
xor U9802 (N_9802,N_2792,N_2320);
or U9803 (N_9803,N_872,N_1282);
or U9804 (N_9804,N_3119,N_354);
or U9805 (N_9805,N_2814,N_4292);
nand U9806 (N_9806,N_900,N_4169);
or U9807 (N_9807,N_4103,N_4079);
or U9808 (N_9808,N_1608,N_4716);
or U9809 (N_9809,N_3276,N_599);
or U9810 (N_9810,N_1268,N_1355);
xnor U9811 (N_9811,N_4376,N_4677);
nand U9812 (N_9812,N_3170,N_4201);
nor U9813 (N_9813,N_3319,N_1984);
nand U9814 (N_9814,N_3867,N_2066);
xnor U9815 (N_9815,N_2068,N_24);
xnor U9816 (N_9816,N_143,N_1006);
or U9817 (N_9817,N_4631,N_1590);
and U9818 (N_9818,N_1049,N_2925);
and U9819 (N_9819,N_4239,N_1717);
xor U9820 (N_9820,N_4186,N_2699);
or U9821 (N_9821,N_2659,N_2434);
nor U9822 (N_9822,N_4525,N_4908);
or U9823 (N_9823,N_3435,N_4599);
and U9824 (N_9824,N_4418,N_4281);
or U9825 (N_9825,N_1053,N_2083);
xnor U9826 (N_9826,N_2153,N_488);
nand U9827 (N_9827,N_1659,N_1479);
or U9828 (N_9828,N_4740,N_362);
or U9829 (N_9829,N_1139,N_2939);
or U9830 (N_9830,N_3964,N_1118);
and U9831 (N_9831,N_4045,N_2242);
nor U9832 (N_9832,N_3847,N_1534);
and U9833 (N_9833,N_1041,N_3305);
xor U9834 (N_9834,N_4858,N_4020);
or U9835 (N_9835,N_3138,N_1867);
or U9836 (N_9836,N_2098,N_4621);
or U9837 (N_9837,N_1764,N_1839);
and U9838 (N_9838,N_3719,N_4792);
nand U9839 (N_9839,N_3910,N_3709);
nor U9840 (N_9840,N_864,N_2929);
or U9841 (N_9841,N_3834,N_4611);
and U9842 (N_9842,N_2142,N_4762);
nor U9843 (N_9843,N_2685,N_1696);
and U9844 (N_9844,N_3256,N_4703);
nor U9845 (N_9845,N_1726,N_3502);
nand U9846 (N_9846,N_244,N_2544);
nand U9847 (N_9847,N_366,N_1557);
nor U9848 (N_9848,N_210,N_1292);
and U9849 (N_9849,N_3427,N_4964);
or U9850 (N_9850,N_4716,N_483);
or U9851 (N_9851,N_1520,N_3011);
or U9852 (N_9852,N_775,N_1461);
or U9853 (N_9853,N_4211,N_91);
xnor U9854 (N_9854,N_554,N_4851);
nand U9855 (N_9855,N_1911,N_313);
nand U9856 (N_9856,N_2689,N_1694);
or U9857 (N_9857,N_4144,N_2048);
nor U9858 (N_9858,N_3164,N_416);
nor U9859 (N_9859,N_1560,N_754);
or U9860 (N_9860,N_1006,N_4280);
xor U9861 (N_9861,N_2199,N_2714);
xnor U9862 (N_9862,N_1254,N_2003);
nand U9863 (N_9863,N_2195,N_4366);
or U9864 (N_9864,N_4746,N_626);
or U9865 (N_9865,N_1192,N_3748);
nor U9866 (N_9866,N_3573,N_998);
nor U9867 (N_9867,N_373,N_4554);
xor U9868 (N_9868,N_4010,N_640);
nor U9869 (N_9869,N_4655,N_962);
nor U9870 (N_9870,N_3223,N_2297);
nand U9871 (N_9871,N_3718,N_1044);
nand U9872 (N_9872,N_3581,N_3118);
nor U9873 (N_9873,N_1365,N_2523);
and U9874 (N_9874,N_4706,N_2301);
nor U9875 (N_9875,N_3543,N_386);
xnor U9876 (N_9876,N_473,N_2648);
nor U9877 (N_9877,N_3077,N_1231);
and U9878 (N_9878,N_4121,N_3146);
and U9879 (N_9879,N_1160,N_4757);
nor U9880 (N_9880,N_4740,N_3273);
xnor U9881 (N_9881,N_1662,N_3210);
nor U9882 (N_9882,N_4503,N_1316);
nand U9883 (N_9883,N_280,N_2393);
or U9884 (N_9884,N_4374,N_2697);
xor U9885 (N_9885,N_4568,N_828);
nand U9886 (N_9886,N_3194,N_2525);
or U9887 (N_9887,N_528,N_2088);
nor U9888 (N_9888,N_2485,N_2003);
xnor U9889 (N_9889,N_1060,N_4617);
xnor U9890 (N_9890,N_2704,N_4619);
nand U9891 (N_9891,N_4624,N_2192);
nand U9892 (N_9892,N_702,N_1127);
or U9893 (N_9893,N_3117,N_477);
or U9894 (N_9894,N_1389,N_4212);
and U9895 (N_9895,N_954,N_3326);
xor U9896 (N_9896,N_182,N_2150);
xor U9897 (N_9897,N_4536,N_878);
nor U9898 (N_9898,N_1490,N_4661);
nor U9899 (N_9899,N_858,N_1154);
and U9900 (N_9900,N_1502,N_363);
and U9901 (N_9901,N_1976,N_3078);
nor U9902 (N_9902,N_1555,N_989);
or U9903 (N_9903,N_4255,N_635);
xnor U9904 (N_9904,N_1002,N_3133);
xor U9905 (N_9905,N_2729,N_2774);
and U9906 (N_9906,N_3536,N_1378);
xnor U9907 (N_9907,N_4365,N_2876);
nor U9908 (N_9908,N_1519,N_242);
nand U9909 (N_9909,N_1171,N_3844);
or U9910 (N_9910,N_950,N_4669);
nand U9911 (N_9911,N_2870,N_3200);
nand U9912 (N_9912,N_3874,N_4951);
nand U9913 (N_9913,N_2117,N_2966);
nand U9914 (N_9914,N_3525,N_3497);
nor U9915 (N_9915,N_3180,N_3278);
or U9916 (N_9916,N_3255,N_480);
or U9917 (N_9917,N_3017,N_1518);
nor U9918 (N_9918,N_4040,N_1647);
xnor U9919 (N_9919,N_99,N_82);
and U9920 (N_9920,N_2394,N_3163);
nor U9921 (N_9921,N_2482,N_2536);
and U9922 (N_9922,N_1985,N_26);
xnor U9923 (N_9923,N_4545,N_987);
nand U9924 (N_9924,N_689,N_3832);
or U9925 (N_9925,N_4282,N_803);
nand U9926 (N_9926,N_2791,N_3753);
nor U9927 (N_9927,N_360,N_3444);
xor U9928 (N_9928,N_4635,N_1736);
nand U9929 (N_9929,N_4861,N_2911);
nand U9930 (N_9930,N_2715,N_3576);
and U9931 (N_9931,N_4546,N_2192);
nand U9932 (N_9932,N_2899,N_2920);
or U9933 (N_9933,N_694,N_1620);
or U9934 (N_9934,N_885,N_1135);
nand U9935 (N_9935,N_2733,N_4723);
xnor U9936 (N_9936,N_1569,N_3720);
nor U9937 (N_9937,N_1762,N_4988);
nand U9938 (N_9938,N_2876,N_17);
nand U9939 (N_9939,N_423,N_988);
nand U9940 (N_9940,N_3137,N_1406);
nor U9941 (N_9941,N_2459,N_1295);
nand U9942 (N_9942,N_4406,N_553);
and U9943 (N_9943,N_4174,N_4371);
xnor U9944 (N_9944,N_4151,N_2097);
nor U9945 (N_9945,N_3775,N_2811);
nor U9946 (N_9946,N_169,N_1993);
nor U9947 (N_9947,N_4583,N_1849);
or U9948 (N_9948,N_3421,N_1988);
nand U9949 (N_9949,N_469,N_2155);
and U9950 (N_9950,N_555,N_2532);
nor U9951 (N_9951,N_866,N_4741);
and U9952 (N_9952,N_286,N_2070);
or U9953 (N_9953,N_2936,N_4768);
and U9954 (N_9954,N_259,N_1171);
xor U9955 (N_9955,N_2131,N_2319);
xor U9956 (N_9956,N_2327,N_4576);
or U9957 (N_9957,N_824,N_4017);
or U9958 (N_9958,N_44,N_4686);
nand U9959 (N_9959,N_1459,N_4568);
nand U9960 (N_9960,N_116,N_204);
xor U9961 (N_9961,N_2488,N_1694);
and U9962 (N_9962,N_2197,N_4710);
and U9963 (N_9963,N_1594,N_353);
nor U9964 (N_9964,N_2302,N_4082);
and U9965 (N_9965,N_4556,N_4816);
nand U9966 (N_9966,N_1609,N_3635);
nor U9967 (N_9967,N_4843,N_4286);
nand U9968 (N_9968,N_2914,N_2769);
xnor U9969 (N_9969,N_688,N_3033);
or U9970 (N_9970,N_4168,N_1261);
or U9971 (N_9971,N_423,N_4980);
xor U9972 (N_9972,N_4053,N_1984);
nand U9973 (N_9973,N_4571,N_2945);
and U9974 (N_9974,N_3956,N_3023);
xor U9975 (N_9975,N_3427,N_348);
and U9976 (N_9976,N_165,N_96);
nand U9977 (N_9977,N_3032,N_2128);
xnor U9978 (N_9978,N_3349,N_1535);
nor U9979 (N_9979,N_1657,N_3544);
nor U9980 (N_9980,N_776,N_1292);
or U9981 (N_9981,N_2795,N_1996);
and U9982 (N_9982,N_2615,N_1993);
xor U9983 (N_9983,N_881,N_123);
xnor U9984 (N_9984,N_2334,N_3518);
nand U9985 (N_9985,N_1785,N_4284);
and U9986 (N_9986,N_3889,N_4950);
xnor U9987 (N_9987,N_4112,N_3581);
nand U9988 (N_9988,N_1551,N_4631);
nor U9989 (N_9989,N_4721,N_3008);
and U9990 (N_9990,N_1215,N_1258);
and U9991 (N_9991,N_362,N_4700);
nand U9992 (N_9992,N_3073,N_1761);
or U9993 (N_9993,N_4531,N_3106);
xnor U9994 (N_9994,N_209,N_2793);
or U9995 (N_9995,N_1743,N_4079);
xnor U9996 (N_9996,N_3942,N_355);
xor U9997 (N_9997,N_4700,N_3475);
nand U9998 (N_9998,N_3897,N_4907);
nand U9999 (N_9999,N_3256,N_221);
nor U10000 (N_10000,N_8068,N_7756);
xnor U10001 (N_10001,N_6373,N_9793);
or U10002 (N_10002,N_7956,N_7507);
and U10003 (N_10003,N_7683,N_7424);
xnor U10004 (N_10004,N_7573,N_5511);
and U10005 (N_10005,N_5136,N_7843);
or U10006 (N_10006,N_9447,N_6455);
or U10007 (N_10007,N_6606,N_5345);
and U10008 (N_10008,N_6332,N_8346);
or U10009 (N_10009,N_6170,N_5851);
nand U10010 (N_10010,N_9971,N_8999);
and U10011 (N_10011,N_5602,N_7081);
nand U10012 (N_10012,N_6178,N_9074);
nand U10013 (N_10013,N_6861,N_6388);
and U10014 (N_10014,N_7677,N_5570);
or U10015 (N_10015,N_8252,N_6234);
xor U10016 (N_10016,N_8279,N_9945);
nor U10017 (N_10017,N_8630,N_8738);
or U10018 (N_10018,N_8929,N_7347);
xor U10019 (N_10019,N_8997,N_7164);
or U10020 (N_10020,N_6534,N_6143);
nand U10021 (N_10021,N_8249,N_5043);
and U10022 (N_10022,N_9803,N_8573);
or U10023 (N_10023,N_6079,N_7777);
xor U10024 (N_10024,N_5133,N_8967);
and U10025 (N_10025,N_8169,N_8422);
and U10026 (N_10026,N_7189,N_6897);
nand U10027 (N_10027,N_7701,N_9530);
nor U10028 (N_10028,N_9229,N_8050);
nor U10029 (N_10029,N_5660,N_5295);
and U10030 (N_10030,N_6272,N_8183);
nor U10031 (N_10031,N_8828,N_6017);
nand U10032 (N_10032,N_7393,N_5535);
xnor U10033 (N_10033,N_8497,N_9920);
nor U10034 (N_10034,N_8141,N_6638);
nor U10035 (N_10035,N_5257,N_6696);
nand U10036 (N_10036,N_6258,N_8676);
nand U10037 (N_10037,N_9354,N_5126);
and U10038 (N_10038,N_9116,N_8774);
xor U10039 (N_10039,N_6888,N_8088);
nand U10040 (N_10040,N_5467,N_8148);
nor U10041 (N_10041,N_5614,N_5209);
or U10042 (N_10042,N_7784,N_5857);
nor U10043 (N_10043,N_8465,N_9451);
nor U10044 (N_10044,N_6653,N_6123);
and U10045 (N_10045,N_5744,N_7828);
or U10046 (N_10046,N_9919,N_5707);
xnor U10047 (N_10047,N_8485,N_7718);
nand U10048 (N_10048,N_5586,N_9981);
and U10049 (N_10049,N_8910,N_8221);
xnor U10050 (N_10050,N_8859,N_5530);
and U10051 (N_10051,N_9661,N_9257);
and U10052 (N_10052,N_8555,N_8207);
nor U10053 (N_10053,N_7229,N_9804);
or U10054 (N_10054,N_8103,N_9862);
or U10055 (N_10055,N_8082,N_7592);
xnor U10056 (N_10056,N_8768,N_7146);
nor U10057 (N_10057,N_7338,N_5553);
and U10058 (N_10058,N_7295,N_9228);
or U10059 (N_10059,N_6228,N_9104);
or U10060 (N_10060,N_5419,N_8228);
nand U10061 (N_10061,N_7589,N_8425);
xnor U10062 (N_10062,N_7243,N_5940);
nand U10063 (N_10063,N_6297,N_6049);
or U10064 (N_10064,N_5245,N_7052);
nor U10065 (N_10065,N_9321,N_8789);
nand U10066 (N_10066,N_6905,N_6129);
nand U10067 (N_10067,N_9733,N_9472);
xor U10068 (N_10068,N_9991,N_9882);
or U10069 (N_10069,N_9018,N_6563);
nand U10070 (N_10070,N_5066,N_6195);
xor U10071 (N_10071,N_7217,N_7272);
xnor U10072 (N_10072,N_9858,N_9526);
nor U10073 (N_10073,N_5781,N_8323);
or U10074 (N_10074,N_9111,N_7053);
and U10075 (N_10075,N_6276,N_8355);
nor U10076 (N_10076,N_9891,N_8753);
and U10077 (N_10077,N_6995,N_9412);
and U10078 (N_10078,N_5955,N_8351);
and U10079 (N_10079,N_7524,N_6298);
or U10080 (N_10080,N_8823,N_8212);
nand U10081 (N_10081,N_9968,N_9106);
nand U10082 (N_10082,N_7055,N_8939);
xor U10083 (N_10083,N_5791,N_5118);
or U10084 (N_10084,N_5160,N_5300);
or U10085 (N_10085,N_8627,N_6350);
xor U10086 (N_10086,N_6240,N_7208);
nand U10087 (N_10087,N_6421,N_6912);
or U10088 (N_10088,N_7618,N_7902);
xnor U10089 (N_10089,N_9827,N_7231);
and U10090 (N_10090,N_6061,N_8655);
or U10091 (N_10091,N_5391,N_9190);
and U10092 (N_10092,N_8399,N_6865);
or U10093 (N_10093,N_6620,N_6539);
xor U10094 (N_10094,N_9033,N_9698);
and U10095 (N_10095,N_6103,N_8136);
xnor U10096 (N_10096,N_7318,N_9380);
or U10097 (N_10097,N_5143,N_9892);
nand U10098 (N_10098,N_8913,N_9810);
and U10099 (N_10099,N_5090,N_5083);
and U10100 (N_10100,N_5282,N_8908);
and U10101 (N_10101,N_8161,N_5740);
nand U10102 (N_10102,N_8712,N_6891);
xnor U10103 (N_10103,N_9368,N_6952);
nand U10104 (N_10104,N_5218,N_9180);
and U10105 (N_10105,N_6675,N_9298);
nand U10106 (N_10106,N_9596,N_9914);
xor U10107 (N_10107,N_6244,N_6593);
or U10108 (N_10108,N_5520,N_8515);
and U10109 (N_10109,N_6855,N_7090);
nor U10110 (N_10110,N_6480,N_9520);
and U10111 (N_10111,N_6256,N_9478);
or U10112 (N_10112,N_5464,N_9797);
nand U10113 (N_10113,N_7493,N_5932);
xor U10114 (N_10114,N_8451,N_8966);
xor U10115 (N_10115,N_5790,N_6774);
and U10116 (N_10116,N_7102,N_9805);
nor U10117 (N_10117,N_9148,N_9603);
and U10118 (N_10118,N_5566,N_5347);
or U10119 (N_10119,N_9517,N_6836);
nand U10120 (N_10120,N_5946,N_5555);
xnor U10121 (N_10121,N_8875,N_5326);
xnor U10122 (N_10122,N_7521,N_7283);
or U10123 (N_10123,N_6608,N_5279);
nand U10124 (N_10124,N_8374,N_6441);
nor U10125 (N_10125,N_8771,N_5098);
and U10126 (N_10126,N_5310,N_7653);
or U10127 (N_10127,N_6409,N_5481);
nand U10128 (N_10128,N_7759,N_5825);
nor U10129 (N_10129,N_8609,N_5177);
xor U10130 (N_10130,N_7630,N_5531);
nor U10131 (N_10131,N_9786,N_9933);
xnor U10132 (N_10132,N_7781,N_9740);
and U10133 (N_10133,N_8008,N_7172);
nand U10134 (N_10134,N_9818,N_6470);
nand U10135 (N_10135,N_6317,N_6219);
and U10136 (N_10136,N_6138,N_7845);
nor U10137 (N_10137,N_8981,N_7080);
xnor U10138 (N_10138,N_9539,N_6878);
nand U10139 (N_10139,N_7133,N_5484);
or U10140 (N_10140,N_7232,N_5580);
and U10141 (N_10141,N_9364,N_7946);
xnor U10142 (N_10142,N_9582,N_5668);
and U10143 (N_10143,N_8414,N_9133);
or U10144 (N_10144,N_9170,N_6011);
nor U10145 (N_10145,N_6783,N_7517);
nor U10146 (N_10146,N_8651,N_6288);
nor U10147 (N_10147,N_6003,N_9140);
nor U10148 (N_10148,N_9842,N_8368);
or U10149 (N_10149,N_7026,N_9068);
and U10150 (N_10150,N_6943,N_5549);
nand U10151 (N_10151,N_6420,N_9870);
or U10152 (N_10152,N_5917,N_6902);
nand U10153 (N_10153,N_8385,N_5096);
xor U10154 (N_10154,N_8091,N_8752);
nor U10155 (N_10155,N_8253,N_6838);
nand U10156 (N_10156,N_6813,N_6767);
or U10157 (N_10157,N_8772,N_7639);
xnor U10158 (N_10158,N_5341,N_6166);
nand U10159 (N_10159,N_8729,N_7577);
and U10160 (N_10160,N_5967,N_7988);
nand U10161 (N_10161,N_8064,N_6303);
nor U10162 (N_10162,N_5731,N_6748);
or U10163 (N_10163,N_5540,N_6910);
and U10164 (N_10164,N_7441,N_9568);
or U10165 (N_10165,N_9495,N_8478);
xnor U10166 (N_10166,N_9988,N_6587);
nand U10167 (N_10167,N_5329,N_5524);
xnor U10168 (N_10168,N_9177,N_5120);
and U10169 (N_10169,N_8698,N_8915);
nor U10170 (N_10170,N_6173,N_7962);
nor U10171 (N_10171,N_6820,N_7773);
xor U10172 (N_10172,N_8898,N_7617);
nor U10173 (N_10173,N_8709,N_7233);
xor U10174 (N_10174,N_8628,N_7136);
and U10175 (N_10175,N_9725,N_8386);
nor U10176 (N_10176,N_9852,N_5921);
or U10177 (N_10177,N_6574,N_5068);
xor U10178 (N_10178,N_5383,N_6389);
or U10179 (N_10179,N_6407,N_8229);
nand U10180 (N_10180,N_5817,N_6210);
and U10181 (N_10181,N_8285,N_5229);
nand U10182 (N_10182,N_5722,N_7159);
xor U10183 (N_10183,N_9017,N_8235);
xnor U10184 (N_10184,N_9807,N_6829);
nor U10185 (N_10185,N_7546,N_9532);
or U10186 (N_10186,N_7046,N_6320);
xor U10187 (N_10187,N_5334,N_6502);
nand U10188 (N_10188,N_8583,N_9511);
or U10189 (N_10189,N_9515,N_8528);
nand U10190 (N_10190,N_6514,N_8877);
and U10191 (N_10191,N_8244,N_8288);
nand U10192 (N_10192,N_6529,N_7952);
nor U10193 (N_10193,N_6301,N_8736);
nor U10194 (N_10194,N_9297,N_7558);
or U10195 (N_10195,N_6374,N_5630);
xor U10196 (N_10196,N_8679,N_9599);
and U10197 (N_10197,N_8572,N_8565);
nor U10198 (N_10198,N_7910,N_6981);
nand U10199 (N_10199,N_7817,N_7354);
or U10200 (N_10200,N_9510,N_6287);
nor U10201 (N_10201,N_9632,N_9152);
nor U10202 (N_10202,N_7495,N_9925);
nor U10203 (N_10203,N_9060,N_6107);
nand U10204 (N_10204,N_8360,N_8424);
nand U10205 (N_10205,N_5205,N_8334);
nand U10206 (N_10206,N_5939,N_9029);
nor U10207 (N_10207,N_9887,N_6866);
or U10208 (N_10208,N_9382,N_8916);
xnor U10209 (N_10209,N_8452,N_9374);
nand U10210 (N_10210,N_9239,N_6410);
xnor U10211 (N_10211,N_9777,N_6472);
nor U10212 (N_10212,N_5124,N_8299);
xnor U10213 (N_10213,N_5877,N_5477);
nand U10214 (N_10214,N_7915,N_7137);
nor U10215 (N_10215,N_7129,N_8191);
and U10216 (N_10216,N_7141,N_5925);
xor U10217 (N_10217,N_6489,N_5889);
xnor U10218 (N_10218,N_8638,N_6954);
nand U10219 (N_10219,N_7368,N_7001);
and U10220 (N_10220,N_8588,N_5434);
nand U10221 (N_10221,N_8393,N_8971);
nand U10222 (N_10222,N_5273,N_7388);
nor U10223 (N_10223,N_7865,N_8570);
nor U10224 (N_10224,N_6874,N_6971);
or U10225 (N_10225,N_8820,N_8416);
and U10226 (N_10226,N_8112,N_9213);
xnor U10227 (N_10227,N_7980,N_7282);
nor U10228 (N_10228,N_8553,N_8443);
nand U10229 (N_10229,N_8317,N_8311);
nand U10230 (N_10230,N_8876,N_7859);
nor U10231 (N_10231,N_8072,N_6707);
or U10232 (N_10232,N_6687,N_9884);
and U10233 (N_10233,N_7278,N_9438);
and U10234 (N_10234,N_7132,N_8687);
nor U10235 (N_10235,N_8521,N_5677);
nand U10236 (N_10236,N_7579,N_9227);
or U10237 (N_10237,N_9776,N_9023);
nor U10238 (N_10238,N_8184,N_6992);
and U10239 (N_10239,N_8430,N_7709);
or U10240 (N_10240,N_9437,N_7011);
nand U10241 (N_10241,N_5881,N_9434);
or U10242 (N_10242,N_9397,N_8338);
xnor U10243 (N_10243,N_5122,N_6640);
xor U10244 (N_10244,N_8688,N_6269);
and U10245 (N_10245,N_6314,N_9541);
or U10246 (N_10246,N_5739,N_6498);
or U10247 (N_10247,N_9323,N_7802);
or U10248 (N_10248,N_6039,N_8165);
or U10249 (N_10249,N_5550,N_5302);
xnor U10250 (N_10250,N_5676,N_9473);
xnor U10251 (N_10251,N_5150,N_7056);
nand U10252 (N_10252,N_9718,N_8657);
or U10253 (N_10253,N_6248,N_5271);
nand U10254 (N_10254,N_8973,N_6486);
nor U10255 (N_10255,N_8232,N_8200);
and U10256 (N_10256,N_6632,N_6842);
xor U10257 (N_10257,N_7912,N_6492);
xor U10258 (N_10258,N_9614,N_5729);
or U10259 (N_10259,N_5084,N_5869);
nor U10260 (N_10260,N_8593,N_9428);
nand U10261 (N_10261,N_6368,N_7300);
xor U10262 (N_10262,N_8312,N_5708);
xor U10263 (N_10263,N_5443,N_5244);
nand U10264 (N_10264,N_9959,N_6154);
xor U10265 (N_10265,N_5620,N_5400);
and U10266 (N_10266,N_9736,N_5836);
xnor U10267 (N_10267,N_5983,N_8217);
nand U10268 (N_10268,N_8703,N_6108);
and U10269 (N_10269,N_7490,N_9835);
and U10270 (N_10270,N_7671,N_7072);
and U10271 (N_10271,N_7004,N_5292);
nand U10272 (N_10272,N_7684,N_7000);
nor U10273 (N_10273,N_5796,N_8800);
nand U10274 (N_10274,N_9595,N_7680);
nor U10275 (N_10275,N_8542,N_5493);
xor U10276 (N_10276,N_9436,N_8378);
or U10277 (N_10277,N_6598,N_8455);
nor U10278 (N_10278,N_5033,N_5417);
nor U10279 (N_10279,N_5180,N_6398);
xor U10280 (N_10280,N_9198,N_9872);
nor U10281 (N_10281,N_7750,N_8541);
nand U10282 (N_10282,N_7760,N_8719);
or U10283 (N_10283,N_6793,N_5855);
xor U10284 (N_10284,N_6776,N_7557);
nor U10285 (N_10285,N_8834,N_5444);
or U10286 (N_10286,N_7450,N_5077);
and U10287 (N_10287,N_8000,N_7181);
nor U10288 (N_10288,N_7735,N_6176);
xor U10289 (N_10289,N_5618,N_7196);
or U10290 (N_10290,N_5651,N_8864);
and U10291 (N_10291,N_6641,N_7687);
xor U10292 (N_10292,N_9547,N_7642);
or U10293 (N_10293,N_7498,N_8233);
or U10294 (N_10294,N_9521,N_8702);
nand U10295 (N_10295,N_5909,N_6315);
and U10296 (N_10296,N_9143,N_9505);
nor U10297 (N_10297,N_8662,N_5036);
xnor U10298 (N_10298,N_7679,N_8585);
nand U10299 (N_10299,N_8036,N_7857);
and U10300 (N_10300,N_8949,N_8196);
xnor U10301 (N_10301,N_5475,N_6698);
xor U10302 (N_10302,N_7798,N_7678);
or U10303 (N_10303,N_8138,N_8004);
and U10304 (N_10304,N_9415,N_7342);
nand U10305 (N_10305,N_5281,N_8535);
or U10306 (N_10306,N_9034,N_8137);
or U10307 (N_10307,N_5961,N_5794);
or U10308 (N_10308,N_7228,N_9999);
and U10309 (N_10309,N_8783,N_9752);
nor U10310 (N_10310,N_8052,N_9543);
xnor U10311 (N_10311,N_9055,N_6834);
xor U10312 (N_10312,N_9086,N_6443);
or U10313 (N_10313,N_6577,N_6704);
or U10314 (N_10314,N_8498,N_5429);
and U10315 (N_10315,N_6230,N_5780);
nand U10316 (N_10316,N_6907,N_6012);
nor U10317 (N_10317,N_9890,N_5834);
or U10318 (N_10318,N_9037,N_5037);
nand U10319 (N_10319,N_7866,N_6739);
nor U10320 (N_10320,N_8906,N_9990);
nor U10321 (N_10321,N_5350,N_8558);
nand U10322 (N_10322,N_8920,N_6830);
and U10323 (N_10323,N_8837,N_6889);
nor U10324 (N_10324,N_6007,N_6382);
or U10325 (N_10325,N_6348,N_5446);
or U10326 (N_10326,N_8094,N_9773);
nand U10327 (N_10327,N_5751,N_6400);
xor U10328 (N_10328,N_7492,N_6887);
nor U10329 (N_10329,N_6718,N_9275);
and U10330 (N_10330,N_6589,N_9983);
and U10331 (N_10331,N_6925,N_8633);
xnor U10332 (N_10332,N_5276,N_6873);
xnor U10333 (N_10333,N_8732,N_7458);
or U10334 (N_10334,N_8919,N_6406);
xnor U10335 (N_10335,N_8392,N_8347);
or U10336 (N_10336,N_9288,N_5319);
nand U10337 (N_10337,N_7363,N_7480);
nor U10338 (N_10338,N_8689,N_9329);
xnor U10339 (N_10339,N_5054,N_9937);
xnor U10340 (N_10340,N_9310,N_5863);
nand U10341 (N_10341,N_6626,N_7239);
and U10342 (N_10342,N_7343,N_9976);
and U10343 (N_10343,N_9403,N_7541);
nor U10344 (N_10344,N_5812,N_8492);
nand U10345 (N_10345,N_7939,N_7059);
nand U10346 (N_10346,N_7886,N_5293);
xnor U10347 (N_10347,N_9262,N_9497);
nand U10348 (N_10348,N_7185,N_8636);
and U10349 (N_10349,N_8626,N_8695);
xnor U10350 (N_10350,N_5225,N_8650);
xnor U10351 (N_10351,N_7504,N_5716);
xor U10352 (N_10352,N_7674,N_7023);
nor U10353 (N_10353,N_7036,N_5656);
xor U10354 (N_10354,N_7006,N_8168);
xnor U10355 (N_10355,N_6342,N_7856);
xnor U10356 (N_10356,N_7744,N_6216);
and U10357 (N_10357,N_9816,N_5134);
nand U10358 (N_10358,N_8637,N_9860);
or U10359 (N_10359,N_9281,N_6917);
nor U10360 (N_10360,N_5502,N_8186);
xnor U10361 (N_10361,N_7968,N_6392);
xor U10362 (N_10362,N_8598,N_7356);
nand U10363 (N_10363,N_9975,N_8105);
or U10364 (N_10364,N_7874,N_9270);
nand U10365 (N_10365,N_8457,N_9387);
nor U10366 (N_10366,N_5669,N_8326);
xnor U10367 (N_10367,N_6055,N_8836);
xor U10368 (N_10368,N_5078,N_6471);
or U10369 (N_10369,N_7281,N_8839);
and U10370 (N_10370,N_5970,N_7177);
nand U10371 (N_10371,N_8135,N_6761);
nand U10372 (N_10372,N_9193,N_5332);
nand U10373 (N_10373,N_6799,N_6844);
or U10374 (N_10374,N_8380,N_6185);
xnor U10375 (N_10375,N_7089,N_6789);
and U10376 (N_10376,N_9877,N_8721);
nor U10377 (N_10377,N_8982,N_6607);
and U10378 (N_10378,N_6884,N_8328);
nand U10379 (N_10379,N_7554,N_7998);
nand U10380 (N_10380,N_5258,N_5250);
nor U10381 (N_10381,N_8641,N_7028);
nand U10382 (N_10382,N_9432,N_9260);
or U10383 (N_10383,N_5029,N_6020);
nand U10384 (N_10384,N_6019,N_5380);
and U10385 (N_10385,N_9164,N_9337);
xnor U10386 (N_10386,N_8379,N_9913);
and U10387 (N_10387,N_7002,N_8020);
xor U10388 (N_10388,N_7176,N_8343);
and U10389 (N_10389,N_5441,N_5014);
or U10390 (N_10390,N_8153,N_9800);
xor U10391 (N_10391,N_7251,N_8824);
nand U10392 (N_10392,N_8419,N_8210);
and U10393 (N_10393,N_5686,N_8976);
or U10394 (N_10394,N_6339,N_9057);
nand U10395 (N_10395,N_5105,N_9817);
and U10396 (N_10396,N_6277,N_9978);
nor U10397 (N_10397,N_6196,N_5952);
nand U10398 (N_10398,N_8175,N_7981);
and U10399 (N_10399,N_6056,N_8056);
or U10400 (N_10400,N_5075,N_5571);
nand U10401 (N_10401,N_7186,N_6986);
and U10402 (N_10402,N_8763,N_7218);
xnor U10403 (N_10403,N_9675,N_8737);
nor U10404 (N_10404,N_5886,N_9970);
or U10405 (N_10405,N_5072,N_5088);
and U10406 (N_10406,N_9040,N_7649);
nor U10407 (N_10407,N_7547,N_9712);
or U10408 (N_10408,N_8938,N_6779);
or U10409 (N_10409,N_6656,N_9615);
and U10410 (N_10410,N_9182,N_5500);
or U10411 (N_10411,N_9254,N_6201);
xor U10412 (N_10412,N_5628,N_5388);
nor U10413 (N_10413,N_8549,N_9989);
nor U10414 (N_10414,N_9246,N_7519);
xnor U10415 (N_10415,N_7899,N_5508);
xor U10416 (N_10416,N_8236,N_6357);
xnor U10417 (N_10417,N_5004,N_9266);
or U10418 (N_10418,N_7613,N_6530);
and U10419 (N_10419,N_8448,N_9813);
nand U10420 (N_10420,N_5975,N_6785);
nor U10421 (N_10421,N_8480,N_6402);
xor U10422 (N_10422,N_9094,N_8123);
nor U10423 (N_10423,N_5215,N_8895);
or U10424 (N_10424,N_6442,N_9731);
or U10425 (N_10425,N_9110,N_9138);
nand U10426 (N_10426,N_5525,N_7467);
and U10427 (N_10427,N_9431,N_6662);
xnor U10428 (N_10428,N_7330,N_7015);
or U10429 (N_10429,N_6165,N_9054);
xnor U10430 (N_10430,N_7139,N_9417);
xor U10431 (N_10431,N_5883,N_9739);
and U10432 (N_10432,N_7958,N_6164);
xnor U10433 (N_10433,N_5506,N_9059);
nand U10434 (N_10434,N_7353,N_5678);
or U10435 (N_10435,N_8403,N_8383);
or U10436 (N_10436,N_6919,N_9896);
nor U10437 (N_10437,N_8799,N_5948);
or U10438 (N_10438,N_6857,N_6304);
nand U10439 (N_10439,N_8741,N_6934);
nor U10440 (N_10440,N_7070,N_8802);
and U10441 (N_10441,N_6229,N_7112);
or U10442 (N_10442,N_6815,N_9823);
xor U10443 (N_10443,N_8557,N_5182);
xnor U10444 (N_10444,N_9588,N_6735);
and U10445 (N_10445,N_5994,N_8048);
nor U10446 (N_10446,N_8446,N_6393);
nor U10447 (N_10447,N_7360,N_9513);
xnor U10448 (N_10448,N_8269,N_8781);
nor U10449 (N_10449,N_6261,N_7106);
or U10450 (N_10450,N_8658,N_7019);
xnor U10451 (N_10451,N_9424,N_5201);
nor U10452 (N_10452,N_9591,N_9036);
or U10453 (N_10453,N_8610,N_5387);
or U10454 (N_10454,N_5510,N_5868);
nor U10455 (N_10455,N_9304,N_8748);
or U10456 (N_10456,N_9664,N_5360);
and U10457 (N_10457,N_6310,N_5342);
and U10458 (N_10458,N_6476,N_9214);
and U10459 (N_10459,N_9700,N_6965);
nor U10460 (N_10460,N_9081,N_9398);
or U10461 (N_10461,N_9419,N_6722);
and U10462 (N_10462,N_5977,N_8977);
and U10463 (N_10463,N_6756,N_7466);
xor U10464 (N_10464,N_6081,N_7147);
and U10465 (N_10465,N_5007,N_6684);
xnor U10466 (N_10466,N_6528,N_6335);
nand U10467 (N_10467,N_6360,N_5112);
xor U10468 (N_10468,N_7913,N_9136);
and U10469 (N_10469,N_7060,N_5935);
nor U10470 (N_10470,N_7785,N_8222);
nor U10471 (N_10471,N_7658,N_9167);
or U10472 (N_10472,N_6197,N_7965);
and U10473 (N_10473,N_5998,N_5170);
nand U10474 (N_10474,N_9871,N_6885);
nand U10475 (N_10475,N_8171,N_8713);
or U10476 (N_10476,N_6549,N_8027);
xor U10477 (N_10477,N_9836,N_8750);
nor U10478 (N_10478,N_9476,N_8532);
nor U10479 (N_10479,N_6939,N_8031);
nor U10480 (N_10480,N_7535,N_9922);
or U10481 (N_10481,N_9694,N_5965);
or U10482 (N_10482,N_8423,N_9215);
and U10483 (N_10483,N_8601,N_7434);
nor U10484 (N_10484,N_9958,N_9366);
or U10485 (N_10485,N_6264,N_6860);
nor U10486 (N_10486,N_8214,N_5269);
or U10487 (N_10487,N_8350,N_6063);
xor U10488 (N_10488,N_9685,N_5228);
and U10489 (N_10489,N_7655,N_5270);
xnor U10490 (N_10490,N_8481,N_9122);
nor U10491 (N_10491,N_6411,N_6791);
or U10492 (N_10492,N_8298,N_5682);
nand U10493 (N_10493,N_5251,N_5027);
nor U10494 (N_10494,N_6646,N_8344);
and U10495 (N_10495,N_5815,N_6161);
nor U10496 (N_10496,N_8707,N_6449);
xor U10497 (N_10497,N_9153,N_8538);
nand U10498 (N_10498,N_8063,N_5827);
nor U10499 (N_10499,N_7428,N_5147);
xnor U10500 (N_10500,N_7763,N_8894);
xor U10501 (N_10501,N_5665,N_6431);
xor U10502 (N_10502,N_7171,N_6157);
or U10503 (N_10503,N_5498,N_8775);
or U10504 (N_10504,N_6711,N_9273);
and U10505 (N_10505,N_8444,N_9255);
or U10506 (N_10506,N_5363,N_8998);
nand U10507 (N_10507,N_7762,N_5890);
or U10508 (N_10508,N_8745,N_9585);
nor U10509 (N_10509,N_7926,N_8293);
xnor U10510 (N_10510,N_9679,N_6697);
and U10511 (N_10511,N_5073,N_7369);
xor U10512 (N_10512,N_7993,N_5547);
or U10513 (N_10513,N_7042,N_7530);
nor U10514 (N_10514,N_7813,N_8447);
or U10515 (N_10515,N_6334,N_6396);
nand U10516 (N_10516,N_5370,N_6403);
nor U10517 (N_10517,N_6322,N_8499);
nand U10518 (N_10518,N_6886,N_7035);
and U10519 (N_10519,N_8625,N_8817);
nor U10520 (N_10520,N_9309,N_7609);
nand U10521 (N_10521,N_7665,N_6028);
xnor U10522 (N_10522,N_8503,N_5186);
xnor U10523 (N_10523,N_7627,N_5987);
nor U10524 (N_10524,N_7851,N_6814);
xor U10525 (N_10525,N_5721,N_9569);
or U10526 (N_10526,N_9762,N_6974);
xor U10527 (N_10527,N_7990,N_6175);
xor U10528 (N_10528,N_6899,N_7374);
xnor U10529 (N_10529,N_8569,N_6363);
and U10530 (N_10530,N_8329,N_6506);
and U10531 (N_10531,N_6325,N_5607);
and U10532 (N_10532,N_7418,N_5950);
xor U10533 (N_10533,N_8795,N_8058);
or U10534 (N_10534,N_5082,N_8673);
nor U10535 (N_10535,N_6057,N_5918);
xnor U10536 (N_10536,N_6810,N_5913);
nor U10537 (N_10537,N_6582,N_7863);
xnor U10538 (N_10538,N_9207,N_8014);
or U10539 (N_10539,N_9601,N_8246);
nor U10540 (N_10540,N_5325,N_8605);
or U10541 (N_10541,N_8482,N_6531);
nor U10542 (N_10542,N_8785,N_8891);
nand U10543 (N_10543,N_7628,N_5754);
xnor U10544 (N_10544,N_6780,N_5356);
nand U10545 (N_10545,N_7151,N_9977);
nand U10546 (N_10546,N_7862,N_9315);
nor U10547 (N_10547,N_7497,N_5655);
nor U10548 (N_10548,N_9025,N_9303);
nor U10549 (N_10549,N_7258,N_7398);
or U10550 (N_10550,N_6126,N_7341);
xnor U10551 (N_10551,N_8675,N_7220);
or U10552 (N_10552,N_6665,N_9558);
nor U10553 (N_10553,N_8681,N_8661);
nand U10554 (N_10554,N_9268,N_8815);
xnor U10555 (N_10555,N_8942,N_9834);
or U10556 (N_10556,N_5956,N_5962);
nand U10557 (N_10557,N_7598,N_6249);
and U10558 (N_10558,N_5592,N_5830);
and U10559 (N_10559,N_8672,N_6080);
nor U10560 (N_10560,N_7979,N_5850);
nand U10561 (N_10561,N_5843,N_5389);
nand U10562 (N_10562,N_7404,N_7487);
xnor U10563 (N_10563,N_8691,N_9621);
and U10564 (N_10564,N_5637,N_9910);
xnor U10565 (N_10565,N_9231,N_7266);
and U10566 (N_10566,N_9381,N_9044);
xnor U10567 (N_10567,N_6584,N_8563);
nor U10568 (N_10568,N_9549,N_7063);
nor U10569 (N_10569,N_5621,N_6772);
nand U10570 (N_10570,N_5597,N_5876);
nand U10571 (N_10571,N_6578,N_5101);
and U10572 (N_10572,N_8204,N_9435);
nand U10573 (N_10573,N_5688,N_6109);
or U10574 (N_10574,N_5603,N_9812);
and U10575 (N_10575,N_9647,N_6155);
or U10576 (N_10576,N_8940,N_7820);
nand U10577 (N_10577,N_8550,N_9572);
nand U10578 (N_10578,N_7957,N_8629);
nand U10579 (N_10579,N_5635,N_9534);
nor U10580 (N_10580,N_7803,N_5420);
nand U10581 (N_10581,N_8941,N_8944);
and U10582 (N_10582,N_9339,N_7486);
and U10583 (N_10583,N_8801,N_6694);
nand U10584 (N_10584,N_9519,N_7606);
nor U10585 (N_10585,N_6747,N_6914);
xor U10586 (N_10586,N_5963,N_5772);
and U10587 (N_10587,N_7118,N_6217);
or U10588 (N_10588,N_8617,N_7041);
nor U10589 (N_10589,N_9997,N_8866);
nor U10590 (N_10590,N_8901,N_8188);
nand U10591 (N_10591,N_5793,N_7277);
or U10592 (N_10592,N_5583,N_8632);
nand U10593 (N_10593,N_5046,N_6732);
or U10594 (N_10594,N_5633,N_6674);
xor U10595 (N_10595,N_8524,N_6262);
xor U10596 (N_10596,N_6331,N_7326);
and U10597 (N_10597,N_8727,N_9248);
or U10598 (N_10598,N_8790,N_6983);
nand U10599 (N_10599,N_8816,N_8127);
nand U10600 (N_10600,N_8692,N_9375);
xor U10601 (N_10601,N_6548,N_9848);
nor U10602 (N_10602,N_8195,N_6058);
and U10603 (N_10603,N_9617,N_7585);
nand U10604 (N_10604,N_7681,N_7876);
and U10605 (N_10605,N_6456,N_6202);
nand U10606 (N_10606,N_9225,N_8653);
nand U10607 (N_10607,N_6890,N_5306);
or U10608 (N_10608,N_9112,N_5548);
nand U10609 (N_10609,N_8243,N_8889);
or U10610 (N_10610,N_9311,N_5567);
nor U10611 (N_10611,N_8885,N_7379);
nand U10612 (N_10612,N_9592,N_9395);
nand U10613 (N_10613,N_7626,N_6218);
nor U10614 (N_10614,N_8220,N_6179);
xnor U10615 (N_10615,N_5880,N_6194);
xor U10616 (N_10616,N_8580,N_8507);
and U10617 (N_10617,N_7325,N_7529);
xor U10618 (N_10618,N_6516,N_5899);
nor U10619 (N_10619,N_5040,N_9673);
or U10620 (N_10620,N_5573,N_8083);
xor U10621 (N_10621,N_6623,N_6811);
xnor U10622 (N_10622,N_5809,N_9801);
and U10623 (N_10623,N_7449,N_9422);
and U10624 (N_10624,N_5725,N_9646);
and U10625 (N_10625,N_8440,N_7875);
nand U10626 (N_10626,N_8950,N_8822);
xnor U10627 (N_10627,N_6333,N_5463);
and U10628 (N_10628,N_8992,N_6383);
nor U10629 (N_10629,N_7025,N_7719);
nand U10630 (N_10630,N_8798,N_8804);
and U10631 (N_10631,N_7443,N_5726);
or U10632 (N_10632,N_7774,N_5010);
or U10633 (N_10633,N_5920,N_5436);
and U10634 (N_10634,N_8435,N_6817);
and U10635 (N_10635,N_6485,N_6242);
nand U10636 (N_10636,N_6072,N_6231);
and U10637 (N_10637,N_5097,N_6022);
nand U10638 (N_10638,N_9453,N_9385);
nand U10639 (N_10639,N_6115,N_7700);
and U10640 (N_10640,N_9965,N_7645);
xnor U10641 (N_10641,N_5941,N_5521);
xnor U10642 (N_10642,N_7651,N_9833);
and U10643 (N_10643,N_9166,N_6533);
and U10644 (N_10644,N_5241,N_8888);
and U10645 (N_10645,N_5039,N_7339);
nor U10646 (N_10646,N_7795,N_8842);
or U10647 (N_10647,N_5728,N_7077);
xor U10648 (N_10648,N_9119,N_9490);
nor U10649 (N_10649,N_7765,N_6945);
and U10650 (N_10650,N_9574,N_5286);
and U10651 (N_10651,N_7088,N_8310);
or U10652 (N_10652,N_8746,N_5242);
or U10653 (N_10653,N_7234,N_7909);
nand U10654 (N_10654,N_9251,N_5406);
or U10655 (N_10655,N_5461,N_9174);
nor U10656 (N_10656,N_6794,N_8240);
and U10657 (N_10657,N_7580,N_7831);
nor U10658 (N_10658,N_6920,N_8261);
or U10659 (N_10659,N_5050,N_5247);
xnor U10660 (N_10660,N_9677,N_5425);
nor U10661 (N_10661,N_7936,N_5430);
xor U10662 (N_10662,N_7576,N_8381);
xnor U10663 (N_10663,N_6592,N_6977);
nor U10664 (N_10664,N_5800,N_6051);
and U10665 (N_10665,N_7331,N_6717);
or U10666 (N_10666,N_8092,N_6180);
nand U10667 (N_10667,N_5062,N_7484);
nor U10668 (N_10668,N_6652,N_9316);
nor U10669 (N_10669,N_6515,N_5574);
nor U10670 (N_10670,N_5552,N_6370);
and U10671 (N_10671,N_5061,N_6673);
nand U10672 (N_10672,N_7100,N_7086);
and U10673 (N_10673,N_9774,N_7463);
and U10674 (N_10674,N_7115,N_7094);
nand U10675 (N_10675,N_6609,N_5462);
nor U10676 (N_10676,N_7878,N_7340);
xnor U10677 (N_10677,N_5870,N_5476);
or U10678 (N_10678,N_7987,N_6215);
nor U10679 (N_10679,N_8227,N_9683);
or U10680 (N_10680,N_6068,N_6430);
or U10681 (N_10681,N_8074,N_8505);
xor U10682 (N_10682,N_9955,N_7378);
nand U10683 (N_10683,N_8007,N_8476);
nand U10684 (N_10684,N_5479,N_6329);
xnor U10685 (N_10685,N_6114,N_7722);
nor U10686 (N_10686,N_9830,N_9850);
nor U10687 (N_10687,N_5456,N_9820);
or U10688 (N_10688,N_6630,N_9105);
xor U10689 (N_10689,N_7991,N_5437);
xor U10690 (N_10690,N_6273,N_5819);
and U10691 (N_10691,N_9336,N_7873);
xor U10692 (N_10692,N_6464,N_8102);
nand U10693 (N_10693,N_9715,N_5736);
and U10694 (N_10694,N_9252,N_9459);
or U10695 (N_10695,N_5702,N_8607);
or U10696 (N_10696,N_7397,N_9555);
or U10697 (N_10697,N_5914,N_8364);
and U10698 (N_10698,N_6460,N_8511);
and U10699 (N_10699,N_8993,N_7116);
or U10700 (N_10700,N_5554,N_7994);
xnor U10701 (N_10701,N_5166,N_8740);
or U10702 (N_10702,N_6637,N_8013);
or U10703 (N_10703,N_9363,N_9600);
nor U10704 (N_10704,N_6425,N_6649);
nand U10705 (N_10705,N_6121,N_5626);
and U10706 (N_10706,N_8693,N_5601);
xor U10707 (N_10707,N_6991,N_9000);
xnor U10708 (N_10708,N_5777,N_7757);
xnor U10709 (N_10709,N_6975,N_9749);
and U10710 (N_10710,N_7032,N_9775);
or U10711 (N_10711,N_7488,N_7109);
or U10712 (N_10712,N_9189,N_8934);
or U10713 (N_10713,N_6603,N_8862);
and U10714 (N_10714,N_8670,N_6953);
or U10715 (N_10715,N_6379,N_6010);
nand U10716 (N_10716,N_8120,N_9706);
nand U10717 (N_10717,N_6353,N_8659);
and U10718 (N_10718,N_8963,N_6677);
and U10719 (N_10719,N_6415,N_8852);
or U10720 (N_10720,N_5519,N_8180);
xor U10721 (N_10721,N_8441,N_6084);
nor U10722 (N_10722,N_6013,N_9245);
xor U10723 (N_10723,N_5232,N_9985);
or U10724 (N_10724,N_6595,N_8865);
nand U10725 (N_10725,N_7638,N_9163);
nor U10726 (N_10726,N_9188,N_9533);
nand U10727 (N_10727,N_7861,N_6347);
nand U10728 (N_10728,N_9849,N_5767);
nor U10729 (N_10729,N_5192,N_9173);
and U10730 (N_10730,N_6579,N_5249);
xor U10731 (N_10731,N_7950,N_6961);
or U10732 (N_10732,N_6413,N_5207);
or U10733 (N_10733,N_5904,N_7782);
nor U10734 (N_10734,N_5392,N_6752);
nand U10735 (N_10735,N_7314,N_8648);
nor U10736 (N_10736,N_9267,N_8367);
nor U10737 (N_10737,N_5458,N_7768);
and U10738 (N_10738,N_7891,N_8099);
xor U10739 (N_10739,N_6127,N_9726);
xnor U10740 (N_10740,N_7372,N_9888);
nand U10741 (N_10741,N_5324,N_8395);
and U10742 (N_10742,N_8983,N_8543);
or U10743 (N_10743,N_6445,N_7753);
and U10744 (N_10744,N_8400,N_5262);
xnor U10745 (N_10745,N_5371,N_8053);
nor U10746 (N_10746,N_8051,N_8342);
and U10747 (N_10747,N_7586,N_9721);
nor U10748 (N_10748,N_7932,N_7951);
and U10749 (N_10749,N_8155,N_8046);
or U10750 (N_10750,N_9179,N_6742);
xnor U10751 (N_10751,N_7667,N_6358);
and U10752 (N_10752,N_7666,N_8514);
nor U10753 (N_10753,N_5418,N_8152);
xnor U10754 (N_10754,N_9563,N_6137);
and U10755 (N_10755,N_7099,N_6628);
and U10756 (N_10756,N_6622,N_5330);
or U10757 (N_10757,N_5311,N_7870);
and U10758 (N_10758,N_5543,N_5658);
nor U10759 (N_10759,N_8087,N_7169);
or U10760 (N_10760,N_6495,N_6300);
and U10761 (N_10761,N_9129,N_9705);
or U10762 (N_10762,N_7984,N_9930);
nand U10763 (N_10763,N_9665,N_8282);
or U10764 (N_10764,N_9405,N_8710);
nand U10765 (N_10765,N_5931,N_6872);
nand U10766 (N_10766,N_9616,N_5298);
xor U10767 (N_10767,N_7302,N_6083);
nand U10768 (N_10768,N_5352,N_7978);
and U10769 (N_10769,N_5145,N_7058);
nor U10770 (N_10770,N_5611,N_7140);
nand U10771 (N_10771,N_6030,N_6354);
or U10772 (N_10772,N_9607,N_9358);
nor U10773 (N_10773,N_7925,N_6151);
xnor U10774 (N_10774,N_6660,N_5168);
xnor U10775 (N_10775,N_5551,N_7696);
and U10776 (N_10776,N_7597,N_6988);
and U10777 (N_10777,N_5240,N_9028);
xor U10778 (N_10778,N_9441,N_5424);
nor U10779 (N_10779,N_9293,N_5117);
or U10780 (N_10780,N_9035,N_7810);
xnor U10781 (N_10781,N_5114,N_8181);
nand U10782 (N_10782,N_5944,N_9481);
and U10783 (N_10783,N_7462,N_8242);
and U10784 (N_10784,N_9373,N_8201);
xnor U10785 (N_10785,N_7506,N_5499);
xor U10786 (N_10786,N_5927,N_9048);
xnor U10787 (N_10787,N_7685,N_5806);
nor U10788 (N_10788,N_6613,N_8882);
or U10789 (N_10789,N_7929,N_9734);
nor U10790 (N_10790,N_8958,N_8128);
and U10791 (N_10791,N_8863,N_8473);
nor U10792 (N_10792,N_8035,N_8257);
or U10793 (N_10793,N_5144,N_7286);
nand U10794 (N_10794,N_5103,N_9113);
and U10795 (N_10795,N_8111,N_7525);
nand U10796 (N_10796,N_9026,N_6198);
nor U10797 (N_10797,N_9659,N_5969);
and U10798 (N_10798,N_7634,N_6564);
nor U10799 (N_10799,N_8032,N_6140);
xor U10800 (N_10800,N_5109,N_8145);
or U10801 (N_10801,N_7726,N_9046);
nor U10802 (N_10802,N_9633,N_6819);
nand U10803 (N_10803,N_7973,N_6937);
nor U10804 (N_10804,N_8846,N_6604);
or U10805 (N_10805,N_7321,N_7328);
and U10806 (N_10806,N_5775,N_6743);
and U10807 (N_10807,N_9221,N_6879);
nor U10808 (N_10808,N_6540,N_7408);
nand U10809 (N_10809,N_9095,N_9886);
or U10810 (N_10810,N_8665,N_7901);
nand U10811 (N_10811,N_7292,N_5709);
xnor U10812 (N_10812,N_6701,N_7167);
nor U10813 (N_10813,N_7727,N_5703);
nor U10814 (N_10814,N_8512,N_5055);
or U10815 (N_10815,N_8272,N_9264);
and U10816 (N_10816,N_8896,N_6015);
and U10817 (N_10817,N_5681,N_8260);
or U10818 (N_10818,N_6494,N_9100);
nand U10819 (N_10819,N_7391,N_9244);
nand U10820 (N_10820,N_9552,N_8113);
and U10821 (N_10821,N_7123,N_6666);
and U10822 (N_10822,N_6054,N_6024);
and U10823 (N_10823,N_7306,N_8537);
and U10824 (N_10824,N_6536,N_8190);
nand U10825 (N_10825,N_9007,N_9645);
and U10826 (N_10826,N_5871,N_9523);
or U10827 (N_10827,N_7456,N_7436);
and U10828 (N_10828,N_8953,N_9618);
nor U10829 (N_10829,N_8621,N_5211);
xor U10830 (N_10830,N_9165,N_8584);
and U10831 (N_10831,N_9560,N_9662);
nor U10832 (N_10832,N_6291,N_6098);
or U10833 (N_10833,N_9702,N_8362);
or U10834 (N_10834,N_6542,N_6740);
nand U10835 (N_10835,N_6457,N_8970);
or U10836 (N_10836,N_8417,N_8552);
nand U10837 (N_10837,N_8567,N_7464);
and U10838 (N_10838,N_6458,N_7552);
and U10839 (N_10839,N_7880,N_5613);
xnor U10840 (N_10840,N_9730,N_6274);
and U10841 (N_10841,N_8952,N_8483);
and U10842 (N_10842,N_6659,N_8060);
xnor U10843 (N_10843,N_7516,N_8140);
nand U10844 (N_10844,N_5001,N_8739);
nor U10845 (N_10845,N_8642,N_7567);
and U10846 (N_10846,N_6426,N_8450);
nor U10847 (N_10847,N_5152,N_8396);
or U10848 (N_10848,N_7829,N_8874);
nor U10849 (N_10849,N_5557,N_6695);
nand U10850 (N_10850,N_7835,N_6428);
and U10851 (N_10851,N_7376,N_7175);
xnor U10852 (N_10852,N_7201,N_9707);
nor U10853 (N_10853,N_6808,N_5119);
xor U10854 (N_10854,N_8301,N_7644);
xor U10855 (N_10855,N_7928,N_6520);
nand U10856 (N_10856,N_8556,N_9171);
and U10857 (N_10857,N_9527,N_5773);
nand U10858 (N_10858,N_9450,N_5469);
or U10859 (N_10859,N_5556,N_8751);
and U10860 (N_10860,N_6852,N_6720);
nand U10861 (N_10861,N_5011,N_7411);
nand U10862 (N_10862,N_5308,N_9482);
nand U10863 (N_10863,N_8907,N_9001);
xnor U10864 (N_10864,N_9584,N_5589);
xnor U10865 (N_10865,N_5372,N_5376);
nor U10866 (N_10866,N_8122,N_7149);
nor U10867 (N_10867,N_8730,N_8151);
nand U10868 (N_10868,N_5653,N_6716);
nor U10869 (N_10869,N_6286,N_7748);
nor U10870 (N_10870,N_6524,N_5856);
or U10871 (N_10871,N_5972,N_8777);
nand U10872 (N_10872,N_8341,N_7563);
or U10873 (N_10873,N_8990,N_7610);
xor U10874 (N_10874,N_8418,N_7697);
xor U10875 (N_10875,N_7390,N_8157);
nand U10876 (N_10876,N_9766,N_5853);
nor U10877 (N_10877,N_6041,N_5181);
nand U10878 (N_10878,N_5527,N_8595);
nand U10879 (N_10879,N_8132,N_6294);
and U10880 (N_10880,N_8722,N_7732);
xor U10881 (N_10881,N_6736,N_8302);
and U10882 (N_10882,N_8097,N_6927);
or U10883 (N_10883,N_9760,N_7165);
xnor U10884 (N_10884,N_5973,N_5813);
nand U10885 (N_10885,N_8245,N_9305);
nand U10886 (N_10886,N_8361,N_9253);
xor U10887 (N_10887,N_8397,N_6786);
nand U10888 (N_10888,N_5995,N_5351);
xor U10889 (N_10889,N_8018,N_8093);
nor U10890 (N_10890,N_6254,N_8162);
nand U10891 (N_10891,N_7888,N_5260);
nand U10892 (N_10892,N_6882,N_7259);
or U10893 (N_10893,N_8321,N_9144);
or U10894 (N_10894,N_7793,N_9356);
xnor U10895 (N_10895,N_7309,N_9903);
nor U10896 (N_10896,N_8280,N_7942);
and U10897 (N_10897,N_5243,N_7587);
nand U10898 (N_10898,N_7512,N_7062);
or U10899 (N_10899,N_5733,N_6744);
nand U10900 (N_10900,N_5175,N_9377);
nand U10901 (N_10901,N_5666,N_5823);
or U10902 (N_10902,N_6926,N_5413);
xor U10903 (N_10903,N_5059,N_6731);
or U10904 (N_10904,N_6721,N_7533);
nor U10905 (N_10905,N_7884,N_8078);
nor U10906 (N_10906,N_9150,N_9626);
nor U10907 (N_10907,N_6130,N_8205);
and U10908 (N_10908,N_9379,N_9791);
nor U10909 (N_10909,N_9413,N_8646);
nand U10910 (N_10910,N_7401,N_5473);
nor U10911 (N_10911,N_6750,N_9684);
nor U10912 (N_10912,N_5882,N_9120);
nand U10913 (N_10913,N_5449,N_5741);
or U10914 (N_10914,N_9795,N_9277);
xor U10915 (N_10915,N_8644,N_8619);
nand U10916 (N_10916,N_9097,N_5047);
nand U10917 (N_10917,N_6517,N_5106);
nand U10918 (N_10918,N_8356,N_8821);
nand U10919 (N_10919,N_9327,N_8811);
xor U10920 (N_10920,N_5277,N_6069);
or U10921 (N_10921,N_8258,N_8742);
nand U10922 (N_10922,N_5284,N_8159);
nor U10923 (N_10923,N_7568,N_9425);
nor U10924 (N_10924,N_9479,N_9973);
or U10925 (N_10925,N_5887,N_7657);
or U10926 (N_10926,N_8794,N_6600);
nor U10927 (N_10927,N_5317,N_9506);
nor U10928 (N_10928,N_8951,N_7333);
nor U10929 (N_10929,N_7599,N_8797);
nand U10930 (N_10930,N_7588,N_8818);
and U10931 (N_10931,N_9831,N_9754);
and U10932 (N_10932,N_7101,N_7791);
xnor U10933 (N_10933,N_5732,N_5515);
nand U10934 (N_10934,N_6893,N_6627);
or U10935 (N_10935,N_5123,N_7298);
nor U10936 (N_10936,N_9137,N_9041);
or U10937 (N_10937,N_6777,N_8119);
nor U10938 (N_10938,N_6523,N_8109);
xor U10939 (N_10939,N_8735,N_7454);
nor U10940 (N_10940,N_6922,N_8061);
nor U10941 (N_10941,N_8716,N_6545);
nand U10942 (N_10942,N_7303,N_9751);
nand U10943 (N_10943,N_9655,N_5590);
xor U10944 (N_10944,N_8855,N_7660);
or U10945 (N_10945,N_8988,N_9728);
and U10946 (N_10946,N_9146,N_7366);
nand U10947 (N_10947,N_5478,N_6050);
or U10948 (N_10948,N_5497,N_8197);
xnor U10949 (N_10949,N_8903,N_6014);
nand U10950 (N_10950,N_5426,N_7031);
nand U10951 (N_10951,N_5706,N_7953);
and U10952 (N_10952,N_8296,N_7210);
or U10953 (N_10953,N_8912,N_8116);
xor U10954 (N_10954,N_7459,N_7896);
xor U10955 (N_10955,N_9669,N_9697);
xnor U10956 (N_10956,N_6391,N_6848);
nand U10957 (N_10957,N_9359,N_6355);
or U10958 (N_10958,N_5171,N_9176);
nand U10959 (N_10959,N_5492,N_9610);
xnor U10960 (N_10960,N_5900,N_7818);
or U10961 (N_10961,N_8398,N_9211);
and U10962 (N_10962,N_5697,N_5785);
nor U10963 (N_10963,N_9865,N_9235);
nor U10964 (N_10964,N_7669,N_6554);
nor U10965 (N_10965,N_6271,N_5696);
or U10966 (N_10966,N_6351,N_9562);
or U10967 (N_10967,N_7387,N_6093);
nand U10968 (N_10968,N_9934,N_8608);
or U10969 (N_10969,N_8623,N_6846);
nor U10970 (N_10970,N_5712,N_9076);
nor U10971 (N_10971,N_9378,N_7986);
nand U10972 (N_10972,N_5933,N_9072);
and U10973 (N_10973,N_8025,N_7066);
and U10974 (N_10974,N_8034,N_5976);
or U10975 (N_10975,N_5647,N_5746);
nand U10976 (N_10976,N_7869,N_7334);
nand U10977 (N_10977,N_6710,N_5711);
nor U10978 (N_10978,N_9032,N_9414);
nor U10979 (N_10979,N_5230,N_8493);
or U10980 (N_10980,N_9943,N_6444);
nand U10981 (N_10981,N_8432,N_6168);
and U10982 (N_10982,N_5564,N_6706);
or U10983 (N_10983,N_5542,N_5787);
xnor U10984 (N_10984,N_9308,N_9446);
nand U10985 (N_10985,N_9370,N_7437);
xor U10986 (N_10986,N_5717,N_9767);
nor U10987 (N_10987,N_9161,N_5140);
xor U10988 (N_10988,N_9771,N_6921);
and U10989 (N_10989,N_8581,N_7584);
or U10990 (N_10990,N_5758,N_5111);
nand U10991 (N_10991,N_6497,N_7045);
nor U10992 (N_10992,N_9987,N_6259);
nor U10993 (N_10993,N_8975,N_8599);
or U10994 (N_10994,N_8861,N_9750);
and U10995 (N_10995,N_9508,N_7766);
nor U10996 (N_10996,N_6146,N_9088);
or U10997 (N_10997,N_8176,N_6679);
xor U10998 (N_10998,N_8705,N_7930);
nor U10999 (N_10999,N_8467,N_7227);
xnor U11000 (N_11000,N_7738,N_6484);
or U11001 (N_11001,N_5996,N_7461);
nand U11002 (N_11002,N_9948,N_9782);
or U11003 (N_11003,N_8513,N_8108);
and U11004 (N_11004,N_7403,N_9545);
nor U11005 (N_11005,N_6467,N_9889);
xnor U11006 (N_11006,N_7809,N_8755);
nor U11007 (N_11007,N_7723,N_6985);
xor U11008 (N_11008,N_9963,N_8597);
xnor U11009 (N_11009,N_8090,N_9287);
nand U11010 (N_11010,N_5558,N_7836);
xnor U11011 (N_11011,N_8978,N_7273);
nor U11012 (N_11012,N_8568,N_6147);
and U11013 (N_11013,N_6699,N_5604);
or U11014 (N_11014,N_6804,N_6004);
xnor U11015 (N_11015,N_9885,N_5423);
and U11016 (N_11016,N_8991,N_8604);
or U11017 (N_11017,N_7113,N_7839);
xnor U11018 (N_11018,N_7355,N_7240);
xor U11019 (N_11019,N_7977,N_9220);
and U11020 (N_11020,N_7799,N_9583);
nand U11021 (N_11021,N_5076,N_6226);
and U11022 (N_11022,N_8375,N_9399);
or U11023 (N_11023,N_6071,N_6340);
nor U11024 (N_11024,N_8129,N_7867);
and U11025 (N_11025,N_7182,N_9440);
nor U11026 (N_11026,N_7560,N_8487);
nor U11027 (N_11027,N_7252,N_5536);
xor U11028 (N_11028,N_7796,N_8490);
nand U11029 (N_11029,N_7184,N_7734);
and U11030 (N_11030,N_5336,N_5783);
nor U11031 (N_11031,N_7941,N_8547);
nor U11032 (N_11032,N_7367,N_5189);
or U11033 (N_11033,N_5538,N_5684);
and U11034 (N_11034,N_5526,N_8671);
and U11035 (N_11035,N_5687,N_6562);
nand U11036 (N_11036,N_7832,N_8613);
xnor U11037 (N_11037,N_6795,N_7788);
nand U11038 (N_11038,N_7284,N_9131);
and U11039 (N_11039,N_9090,N_9430);
xor U11040 (N_11040,N_9867,N_6769);
nand U11041 (N_11041,N_8591,N_6693);
or U11042 (N_11042,N_8926,N_6469);
nand U11043 (N_11043,N_7729,N_8284);
xor U11044 (N_11044,N_7616,N_7916);
nand U11045 (N_11045,N_8796,N_5390);
xor U11046 (N_11046,N_7448,N_5884);
nor U11047 (N_11047,N_9902,N_5403);
nand U11048 (N_11048,N_8526,N_5314);
nand U11049 (N_11049,N_9078,N_6765);
xor U11050 (N_11050,N_6784,N_9577);
nor U11051 (N_11051,N_8696,N_5275);
nor U11052 (N_11052,N_9101,N_5035);
xor U11053 (N_11053,N_5058,N_8331);
and U11054 (N_11054,N_6207,N_8562);
nand U11055 (N_11055,N_5149,N_9998);
nand U11056 (N_11056,N_9429,N_8114);
nand U11057 (N_11057,N_9681,N_6870);
or U11058 (N_11058,N_8539,N_6976);
nor U11059 (N_11059,N_5929,N_6419);
and U11060 (N_11060,N_5172,N_9570);
or U11061 (N_11061,N_8884,N_7160);
xor U11062 (N_11062,N_6581,N_9464);
and U11063 (N_11063,N_7846,N_5608);
nand U11064 (N_11064,N_8464,N_5227);
and U11065 (N_11065,N_7307,N_6299);
xor U11066 (N_11066,N_5224,N_9756);
and U11067 (N_11067,N_9741,N_7920);
nand U11068 (N_11068,N_7223,N_6026);
and U11069 (N_11069,N_8002,N_7410);
and U11070 (N_11070,N_5196,N_8849);
nand U11071 (N_11071,N_6034,N_8831);
xor U11072 (N_11072,N_9127,N_7933);
xnor U11073 (N_11073,N_9643,N_9559);
nand U11074 (N_11074,N_7632,N_7540);
or U11075 (N_11075,N_5086,N_7301);
nand U11076 (N_11076,N_6292,N_9265);
nand U11077 (N_11077,N_9292,N_7073);
nor U11078 (N_11078,N_9307,N_9371);
nor U11079 (N_11079,N_5396,N_8826);
xor U11080 (N_11080,N_6768,N_6691);
and U11081 (N_11081,N_5369,N_8406);
or U11082 (N_11082,N_8055,N_7471);
nor U11083 (N_11083,N_6672,N_5693);
or U11084 (N_11084,N_6131,N_5715);
xnor U11085 (N_11085,N_5384,N_7268);
nand U11086 (N_11086,N_6290,N_7222);
nand U11087 (N_11087,N_6651,N_5202);
xor U11088 (N_11088,N_8471,N_9699);
nor U11089 (N_11089,N_6062,N_5832);
nand U11090 (N_11090,N_6344,N_7518);
nand U11091 (N_11091,N_9149,N_8239);
nor U11092 (N_11092,N_8047,N_8544);
nand U11093 (N_11093,N_8559,N_9014);
or U11094 (N_11094,N_6475,N_5632);
nor U11095 (N_11095,N_8142,N_5294);
or U11096 (N_11096,N_6002,N_5860);
nor U11097 (N_11097,N_7897,N_9313);
nand U11098 (N_11098,N_5017,N_9907);
nand U11099 (N_11099,N_6509,N_8830);
and U11100 (N_11100,N_6302,N_8674);
xnor U11101 (N_11101,N_7200,N_7556);
or U11102 (N_11102,N_9821,N_6260);
nor U11103 (N_11103,N_8491,N_9620);
and U11104 (N_11104,N_5959,N_8879);
xnor U11105 (N_11105,N_9053,N_5735);
or U11106 (N_11106,N_6931,N_7022);
nand U11107 (N_11107,N_6235,N_9118);
nand U11108 (N_11108,N_6505,N_9240);
nor U11109 (N_11109,N_5445,N_5301);
xor U11110 (N_11110,N_6631,N_8304);
or U11111 (N_11111,N_9218,N_7582);
nor U11112 (N_11112,N_5465,N_5431);
nand U11113 (N_11113,N_5679,N_7711);
xnor U11114 (N_11114,N_6236,N_5596);
and U11115 (N_11115,N_8354,N_5968);
xnor U11116 (N_11116,N_8223,N_5907);
nor U11117 (N_11117,N_8835,N_9921);
and U11118 (N_11118,N_7473,N_6067);
nand U11119 (N_11119,N_6960,N_7571);
nor U11120 (N_11120,N_8965,N_9529);
xor U11121 (N_11121,N_9720,N_6408);
nor U11122 (N_11122,N_8530,N_7130);
nand U11123 (N_11123,N_8560,N_6488);
nor U11124 (N_11124,N_7574,N_8611);
or U11125 (N_11125,N_6781,N_9191);
and U11126 (N_11126,N_6856,N_8880);
or U11127 (N_11127,N_5938,N_6800);
xnor U11128 (N_11128,N_9052,N_8345);
and U11129 (N_11129,N_5575,N_9168);
xor U11130 (N_11130,N_5235,N_7776);
nand U11131 (N_11131,N_7076,N_8166);
xnor U11132 (N_11132,N_9114,N_9799);
nor U11133 (N_11133,N_6401,N_8469);
and U11134 (N_11134,N_8928,N_7527);
nor U11135 (N_11135,N_8684,N_5627);
xor U11136 (N_11136,N_6367,N_5263);
xnor U11137 (N_11137,N_7168,N_5902);
or U11138 (N_11138,N_7607,N_6417);
and U11139 (N_11139,N_7944,N_7308);
nor U11140 (N_11140,N_6588,N_7154);
nand U11141 (N_11141,N_6959,N_6465);
nor U11142 (N_11142,N_9916,N_5689);
xor U11143 (N_11143,N_9735,N_7522);
nor U11144 (N_11144,N_9525,N_5087);
and U11145 (N_11145,N_7375,N_7746);
nor U11146 (N_11146,N_7199,N_6990);
and U11147 (N_11147,N_7124,N_7386);
or U11148 (N_11148,N_5737,N_8144);
nand U11149 (N_11149,N_6338,N_7047);
or U11150 (N_11150,N_9966,N_8946);
nor U11151 (N_11151,N_7267,N_8453);
nand U11152 (N_11152,N_5701,N_7652);
or U11153 (N_11153,N_5185,N_8295);
nor U11154 (N_11154,N_7246,N_7682);
and U11155 (N_11155,N_8215,N_8316);
nand U11156 (N_11156,N_6636,N_5505);
nand U11157 (N_11157,N_9704,N_5533);
or U11158 (N_11158,N_7383,N_8508);
xnor U11159 (N_11159,N_5895,N_5138);
nor U11160 (N_11160,N_5710,N_9445);
nand U11161 (N_11161,N_6311,N_7549);
and U11162 (N_11162,N_5690,N_8010);
and U11163 (N_11163,N_9021,N_9458);
and U11164 (N_11164,N_6111,N_9496);
nand U11165 (N_11165,N_9484,N_7668);
or U11166 (N_11166,N_7427,N_5213);
or U11167 (N_11167,N_6326,N_6077);
nand U11168 (N_11168,N_7931,N_5063);
and U11169 (N_11169,N_8178,N_6989);
nand U11170 (N_11170,N_7173,N_7662);
or U11171 (N_11171,N_6908,N_5471);
or U11172 (N_11172,N_6812,N_9935);
xnor U11173 (N_11173,N_7911,N_7714);
or U11174 (N_11174,N_7225,N_9825);
nor U11175 (N_11175,N_9463,N_8780);
xnor U11176 (N_11176,N_5193,N_6316);
nand U11177 (N_11177,N_8289,N_8405);
nand U11178 (N_11178,N_5989,N_5214);
xnor U11179 (N_11179,N_8409,N_7922);
or U11180 (N_11180,N_8057,N_6947);
or U11181 (N_11181,N_5309,N_9126);
or U11182 (N_11182,N_7238,N_9332);
xor U11183 (N_11183,N_7794,N_8011);
or U11184 (N_11184,N_8845,N_6268);
nor U11185 (N_11185,N_6729,N_5074);
nor U11186 (N_11186,N_9347,N_8590);
nor U11187 (N_11187,N_7162,N_5822);
xor U11188 (N_11188,N_5641,N_5980);
nand U11189 (N_11189,N_9067,N_6737);
nand U11190 (N_11190,N_9084,N_7261);
or U11191 (N_11191,N_5835,N_8411);
nor U11192 (N_11192,N_5491,N_6399);
or U11193 (N_11193,N_7974,N_8081);
or U11194 (N_11194,N_7921,N_7213);
nor U11195 (N_11195,N_8333,N_6541);
or U11196 (N_11196,N_7550,N_7447);
xor U11197 (N_11197,N_8021,N_6018);
and U11198 (N_11198,N_5778,N_7204);
xor U11199 (N_11199,N_5799,N_8421);
nor U11200 (N_11200,N_6341,N_8495);
xnor U11201 (N_11201,N_8306,N_9746);
xor U11202 (N_11202,N_7358,N_9911);
nand U11203 (N_11203,N_5053,N_7065);
nor U11204 (N_11204,N_8445,N_6381);
nand U11205 (N_11205,N_7772,N_7128);
or U11206 (N_11206,N_8488,N_7508);
nor U11207 (N_11207,N_9301,N_9261);
nor U11208 (N_11208,N_8724,N_6778);
xor U11209 (N_11209,N_7431,N_7997);
xor U11210 (N_11210,N_5283,N_8844);
and U11211 (N_11211,N_6787,N_5199);
nand U11212 (N_11212,N_5714,N_6094);
or U11213 (N_11213,N_8325,N_8300);
nor U11214 (N_11214,N_5840,N_5142);
nand U11215 (N_11215,N_7422,N_6877);
and U11216 (N_11216,N_6692,N_7797);
and U11217 (N_11217,N_8517,N_8931);
nor U11218 (N_11218,N_8172,N_7975);
nand U11219 (N_11219,N_6023,N_9567);
xnor U11220 (N_11220,N_5442,N_8202);
or U11221 (N_11221,N_5165,N_8192);
nor U11222 (N_11222,N_9345,N_9256);
nand U11223 (N_11223,N_6560,N_7720);
xnor U11224 (N_11224,N_8484,N_6220);
xor U11225 (N_11225,N_7847,N_9883);
or U11226 (N_11226,N_5594,N_7187);
nand U11227 (N_11227,N_8211,N_6755);
nand U11228 (N_11228,N_8373,N_5085);
and U11229 (N_11229,N_5893,N_7751);
nand U11230 (N_11230,N_7914,N_7469);
xnor U11231 (N_11231,N_7206,N_8778);
or U11232 (N_11232,N_5255,N_6385);
nand U11233 (N_11233,N_5997,N_7935);
nand U11234 (N_11234,N_8969,N_7188);
nor U11235 (N_11235,N_5408,N_9899);
xnor U11236 (N_11236,N_8001,N_5316);
nand U11237 (N_11237,N_9780,N_9103);
or U11238 (N_11238,N_7702,N_9951);
nand U11239 (N_11239,N_7715,N_6404);
xor U11240 (N_11240,N_5667,N_6312);
or U11241 (N_11241,N_7971,N_6461);
nor U11242 (N_11242,N_9394,N_5327);
nor U11243 (N_11243,N_8984,N_6635);
nor U11244 (N_11244,N_6670,N_6405);
nand U11245 (N_11245,N_7740,N_8897);
nor U11246 (N_11246,N_6570,N_5742);
xor U11247 (N_11247,N_8247,N_5768);
xor U11248 (N_11248,N_8039,N_9553);
nor U11249 (N_11249,N_7536,N_7413);
and U11250 (N_11250,N_9500,N_5903);
or U11251 (N_11251,N_7068,N_5349);
or U11252 (N_11252,N_7900,N_7402);
and U11253 (N_11253,N_9351,N_7491);
or U11254 (N_11254,N_7242,N_6586);
or U11255 (N_11255,N_7570,N_7117);
or U11256 (N_11256,N_8401,N_5631);
or U11257 (N_11257,N_6941,N_7420);
and U11258 (N_11258,N_5926,N_8600);
and U11259 (N_11259,N_7373,N_5953);
and U11260 (N_11260,N_8757,N_6016);
nand U11261 (N_11261,N_5600,N_5404);
nand U11262 (N_11262,N_5598,N_8812);
nor U11263 (N_11263,N_8390,N_9814);
nor U11264 (N_11264,N_7879,N_7470);
and U11265 (N_11265,N_5056,N_9918);
nand U11266 (N_11266,N_5421,N_5545);
or U11267 (N_11267,N_5194,N_8518);
nor U11268 (N_11268,N_6052,N_9269);
nor U11269 (N_11269,N_9581,N_9880);
and U11270 (N_11270,N_5757,N_8357);
nor U11271 (N_11271,N_9940,N_6343);
or U11272 (N_11272,N_9340,N_8784);
and U11273 (N_11273,N_8680,N_6906);
nor U11274 (N_11274,N_5849,N_5872);
or U11275 (N_11275,N_7209,N_8305);
nor U11276 (N_11276,N_5415,N_7712);
xnor U11277 (N_11277,N_7871,N_8193);
or U11278 (N_11278,N_7451,N_5934);
and U11279 (N_11279,N_8358,N_7752);
nand U11280 (N_11280,N_6644,N_5943);
xnor U11281 (N_11281,N_8095,N_7170);
nor U11282 (N_11282,N_7600,N_7822);
or U11283 (N_11283,N_9444,N_9687);
nand U11284 (N_11284,N_7528,N_9502);
and U11285 (N_11285,N_5981,N_7057);
nand U11286 (N_11286,N_9181,N_5020);
and U11287 (N_11287,N_6702,N_5833);
and U11288 (N_11288,N_5110,N_8649);
and U11289 (N_11289,N_6823,N_7959);
nor U11290 (N_11290,N_6957,N_6189);
nor U11291 (N_11291,N_6078,N_7531);
xnor U11292 (N_11292,N_5864,N_6950);
nand U11293 (N_11293,N_9783,N_6733);
and U11294 (N_11294,N_6076,N_7892);
and U11295 (N_11295,N_9627,N_7265);
and U11296 (N_11296,N_5993,N_9604);
nand U11297 (N_11297,N_6232,N_9503);
nor U11298 (N_11298,N_6463,N_8225);
and U11299 (N_11299,N_5100,N_7429);
or U11300 (N_11300,N_6558,N_8571);
or U11301 (N_11301,N_7153,N_6088);
xnor U11302 (N_11302,N_6568,N_6639);
or U11303 (N_11303,N_7548,N_7098);
nor U11304 (N_11304,N_5928,N_9941);
and U11305 (N_11305,N_6664,N_6493);
nand U11306 (N_11306,N_5842,N_8281);
or U11307 (N_11307,N_8489,N_5405);
or U11308 (N_11308,N_6669,N_9346);
nor U11309 (N_11309,N_5285,N_6553);
xnor U11310 (N_11310,N_6106,N_9979);
or U11311 (N_11311,N_5750,N_7216);
and U11312 (N_11312,N_9178,N_8764);
xnor U11313 (N_11313,N_7841,N_7291);
nor U11314 (N_11314,N_8960,N_5322);
nor U11315 (N_11315,N_9546,N_8587);
xnor U11316 (N_11316,N_5216,N_6073);
or U11317 (N_11317,N_5865,N_5760);
or U11318 (N_11318,N_7725,N_7083);
xor U11319 (N_11319,N_9579,N_8943);
nand U11320 (N_11320,N_7849,N_6741);
xnor U11321 (N_11321,N_6678,N_9142);
xor U11322 (N_11322,N_5501,N_6597);
and U11323 (N_11323,N_9071,N_9318);
nand U11324 (N_11324,N_7804,N_9186);
and U11325 (N_11325,N_8012,N_8267);
nand U11326 (N_11326,N_5991,N_7423);
and U11327 (N_11327,N_9456,N_8762);
xnor U11328 (N_11328,N_5619,N_7332);
xnor U11329 (N_11329,N_7989,N_9717);
or U11330 (N_11330,N_6192,N_8930);
or U11331 (N_11331,N_7611,N_7852);
xor U11332 (N_11332,N_9091,N_7659);
xor U11333 (N_11333,N_5161,N_9593);
or U11334 (N_11334,N_7008,N_9360);
or U11335 (N_11335,N_6366,N_9972);
or U11336 (N_11336,N_9409,N_5738);
and U11337 (N_11337,N_8994,N_7972);
or U11338 (N_11338,N_5485,N_8096);
xor U11339 (N_11339,N_8231,N_9295);
nand U11340 (N_11340,N_7419,N_8808);
or U11341 (N_11341,N_7069,N_5483);
nor U11342 (N_11342,N_5990,N_9342);
xnor U11343 (N_11343,N_6145,N_6021);
and U11344 (N_11344,N_9693,N_9854);
and U11345 (N_11345,N_6642,N_5804);
xnor U11346 (N_11346,N_8427,N_5000);
and U11347 (N_11347,N_6447,N_5846);
xor U11348 (N_11348,N_8273,N_5280);
or U11349 (N_11349,N_7085,N_9031);
nand U11350 (N_11350,N_6713,N_8501);
and U11351 (N_11351,N_7120,N_8023);
nor U11352 (N_11352,N_7615,N_5206);
xor U11353 (N_11353,N_9757,N_8340);
or U11354 (N_11354,N_8622,N_6211);
nand U11355 (N_11355,N_6491,N_9061);
xor U11356 (N_11356,N_7385,N_5640);
and U11357 (N_11357,N_9204,N_7545);
and U11358 (N_11358,N_6074,N_6663);
xnor U11359 (N_11359,N_7483,N_8714);
nand U11360 (N_11360,N_9826,N_9936);
or U11361 (N_11361,N_9489,N_7095);
or U11362 (N_11362,N_6880,N_9272);
xnor U11363 (N_11363,N_5699,N_8566);
or U11364 (N_11364,N_9411,N_7515);
nor U11365 (N_11365,N_8603,N_9824);
nand U11366 (N_11366,N_5440,N_7211);
or U11367 (N_11367,N_7736,N_6293);
xnor U11368 (N_11368,N_9531,N_8460);
and U11369 (N_11369,N_6591,N_9753);
nand U11370 (N_11370,N_9504,N_7553);
and U11371 (N_11371,N_7288,N_7289);
nand U11372 (N_11372,N_6191,N_5734);
and U11373 (N_11373,N_6571,N_7007);
nand U11374 (N_11374,N_6124,N_5026);
nor U11375 (N_11375,N_6773,N_7948);
or U11376 (N_11376,N_9878,N_6618);
nand U11377 (N_11377,N_8283,N_9668);
xor U11378 (N_11378,N_8516,N_8019);
nand U11379 (N_11379,N_7174,N_7310);
xor U11380 (N_11380,N_5291,N_8756);
nor U11381 (N_11381,N_6827,N_5595);
nand U11382 (N_11382,N_8718,N_6647);
and U11383 (N_11383,N_5818,N_5771);
nand U11384 (N_11384,N_9367,N_7290);
or U11385 (N_11385,N_7999,N_6518);
nor U11386 (N_11386,N_7183,N_6323);
xnor U11387 (N_11387,N_6306,N_7287);
nor U11388 (N_11388,N_6102,N_6397);
nor U11389 (N_11389,N_9107,N_9514);
xnor U11390 (N_11390,N_7016,N_7830);
and U11391 (N_11391,N_6029,N_6929);
nor U11392 (N_11392,N_7742,N_9660);
and U11393 (N_11393,N_5565,N_5221);
and U11394 (N_11394,N_6822,N_8758);
or U11395 (N_11395,N_5591,N_6625);
nand U11396 (N_11396,N_8654,N_8415);
nor U11397 (N_11397,N_6655,N_6547);
nor U11398 (N_11398,N_5582,N_5811);
and U11399 (N_11399,N_5654,N_7389);
nand U11400 (N_11400,N_9631,N_7479);
and U11401 (N_11401,N_8857,N_8219);
nor U11402 (N_11402,N_8870,N_8779);
nor U11403 (N_11403,N_6951,N_7416);
nor U11404 (N_11404,N_5915,N_9357);
nor U11405 (N_11405,N_7604,N_8925);
or U11406 (N_11406,N_6556,N_8459);
and U11407 (N_11407,N_5691,N_9383);
or U11408 (N_11408,N_9512,N_8335);
or U11409 (N_11409,N_7400,N_8336);
nor U11410 (N_11410,N_6468,N_9866);
nor U11411 (N_11411,N_7460,N_8100);
and U11412 (N_11412,N_5135,N_7198);
xnor U11413 (N_11413,N_6182,N_6386);
xnor U11414 (N_11414,N_7143,N_5522);
and U11415 (N_11415,N_5234,N_6605);
xor U11416 (N_11416,N_7444,N_5779);
nand U11417 (N_11417,N_7352,N_5022);
nand U11418 (N_11418,N_7614,N_5127);
and U11419 (N_11419,N_5212,N_9769);
nand U11420 (N_11420,N_6305,N_7881);
and U11421 (N_11421,N_7394,N_7275);
nor U11422 (N_11422,N_5639,N_7009);
or U11423 (N_11423,N_6233,N_8404);
nand U11424 (N_11424,N_9641,N_5867);
nor U11425 (N_11425,N_7887,N_7481);
nor U11426 (N_11426,N_8700,N_6968);
and U11427 (N_11427,N_9695,N_5960);
and U11428 (N_11428,N_8723,N_7304);
and U11429 (N_11429,N_5770,N_5344);
xor U11430 (N_11430,N_6423,N_7694);
and U11431 (N_11431,N_5814,N_5896);
xnor U11432 (N_11432,N_8278,N_9859);
xnor U11433 (N_11433,N_5191,N_9386);
nor U11434 (N_11434,N_9486,N_6289);
nor U11435 (N_11435,N_8044,N_9468);
and U11436 (N_11436,N_7430,N_9159);
xnor U11437 (N_11437,N_8803,N_9573);
nand U11438 (N_11438,N_8725,N_7219);
xor U11439 (N_11439,N_6527,N_8711);
nand U11440 (N_11440,N_6105,N_8370);
nand U11441 (N_11441,N_9200,N_5695);
and U11442 (N_11442,N_6205,N_7619);
or U11443 (N_11443,N_9628,N_8923);
nor U11444 (N_11444,N_7247,N_8917);
nand U11445 (N_11445,N_8412,N_5274);
or U11446 (N_11446,N_6387,N_8840);
nor U11447 (N_11447,N_6380,N_7144);
nand U11448 (N_11448,N_9653,N_5888);
nand U11449 (N_11449,N_6504,N_9956);
nor U11450 (N_11450,N_6152,N_9130);
nand U11451 (N_11451,N_9162,N_5071);
nor U11452 (N_11452,N_5885,N_8956);
xor U11453 (N_11453,N_9087,N_6038);
and U11454 (N_11454,N_8237,N_5019);
xnor U11455 (N_11455,N_8754,N_8536);
xnor U11456 (N_11456,N_7465,N_7230);
nand U11457 (N_11457,N_5176,N_9344);
and U11458 (N_11458,N_9045,N_5985);
xnor U11459 (N_11459,N_9020,N_6184);
or U11460 (N_11460,N_8959,N_5588);
nand U11461 (N_11461,N_9960,N_9950);
and U11462 (N_11462,N_9779,N_5051);
xor U11463 (N_11463,N_5474,N_5910);
or U11464 (N_11464,N_9102,N_5482);
nand U11465 (N_11465,N_6583,N_7255);
and U11466 (N_11466,N_5003,N_6394);
nand U11467 (N_11467,N_5769,N_8529);
nand U11468 (N_11468,N_9875,N_6372);
nor U11469 (N_11469,N_5912,N_6144);
nor U11470 (N_11470,N_7096,N_7844);
nor U11471 (N_11471,N_9815,N_9898);
nand U11472 (N_11472,N_7269,N_6964);
xor U11473 (N_11473,N_6681,N_7489);
xnor U11474 (N_11474,N_9488,N_9141);
nor U11475 (N_11475,N_9839,N_6001);
and U11476 (N_11476,N_6318,N_7583);
xnor U11477 (N_11477,N_5949,N_6585);
xnor U11478 (N_11478,N_5315,N_6416);
or U11479 (N_11479,N_5057,N_8254);
xor U11480 (N_11480,N_5204,N_5745);
and U11481 (N_11481,N_5634,N_7248);
nor U11482 (N_11482,N_7767,N_7395);
nor U11483 (N_11483,N_8041,N_5784);
nand U11484 (N_11484,N_9844,N_5031);
nor U11485 (N_11485,N_7157,N_9857);
and U11486 (N_11486,N_5236,N_9388);
nand U11487 (N_11487,N_9286,N_5364);
and U11488 (N_11488,N_5624,N_9442);
or U11489 (N_11489,N_6867,N_9642);
and U11490 (N_11490,N_5116,N_6361);
nor U11491 (N_11491,N_7675,N_5197);
nor U11492 (N_11492,N_9787,N_8899);
or U11493 (N_11493,N_6206,N_6507);
nand U11494 (N_11494,N_8287,N_9901);
and U11495 (N_11495,N_8297,N_8697);
xnor U11496 (N_11496,N_7769,N_5377);
or U11497 (N_11497,N_7532,N_5265);
and U11498 (N_11498,N_7215,N_8596);
xor U11499 (N_11499,N_6847,N_5911);
and U11500 (N_11500,N_7296,N_7110);
and U11501 (N_11501,N_8902,N_7453);
or U11502 (N_11502,N_7191,N_6535);
xnor U11503 (N_11503,N_6923,N_6616);
xor U11504 (N_11504,N_7226,N_9247);
and U11505 (N_11505,N_8147,N_7789);
xor U11506 (N_11506,N_7741,N_5488);
xnor U11507 (N_11507,N_9019,N_9477);
nand U11508 (N_11508,N_8814,N_6141);
and U11509 (N_11509,N_7030,N_5579);
xnor U11510 (N_11510,N_9249,N_6503);
or U11511 (N_11511,N_6913,N_8203);
nand U11512 (N_11512,N_9652,N_7620);
nor U11513 (N_11513,N_7097,N_7510);
or U11514 (N_11514,N_9156,N_9319);
nand U11515 (N_11515,N_5453,N_7044);
nor U11516 (N_11516,N_6046,N_5452);
nand U11517 (N_11517,N_6754,N_8900);
and U11518 (N_11518,N_7257,N_5038);
and U11519 (N_11519,N_9485,N_8586);
nor U11520 (N_11520,N_5340,N_9184);
nand U11521 (N_11521,N_6065,N_7924);
nand U11522 (N_11522,N_5584,N_6709);
xnor U11523 (N_11523,N_8892,N_5487);
or U11524 (N_11524,N_9790,N_5495);
and U11525 (N_11525,N_6686,N_9637);
nor U11526 (N_11526,N_7426,N_5568);
and U11527 (N_11527,N_8234,N_8825);
nor U11528 (N_11528,N_8766,N_9676);
nor U11529 (N_11529,N_8369,N_6483);
nand U11530 (N_11530,N_5064,N_7039);
nor U11531 (N_11531,N_9942,N_6247);
nor U11532 (N_11532,N_8086,N_8337);
or U11533 (N_11533,N_9452,N_9789);
or U11534 (N_11534,N_7728,N_6725);
xor U11535 (N_11535,N_5756,N_6433);
and U11536 (N_11536,N_9722,N_6451);
or U11537 (N_11537,N_9944,N_9024);
xor U11538 (N_11538,N_6128,N_7365);
and U11539 (N_11539,N_6724,N_8848);
or U11540 (N_11540,N_9230,N_7038);
xnor U11541 (N_11541,N_5381,N_5605);
and U11542 (N_11542,N_8314,N_9058);
nor U11543 (N_11543,N_5030,N_6526);
and U11544 (N_11544,N_9396,N_9233);
or U11545 (N_11545,N_5454,N_5331);
or U11546 (N_11546,N_7855,N_9352);
nor U11547 (N_11547,N_9904,N_9784);
and U11548 (N_11548,N_9772,N_6946);
or U11549 (N_11549,N_9049,N_5231);
nand U11550 (N_11550,N_5859,N_7688);
or U11551 (N_11551,N_7551,N_7457);
and U11552 (N_11552,N_7631,N_7947);
and U11553 (N_11553,N_5139,N_7967);
and U11554 (N_11554,N_6708,N_8130);
nor U11555 (N_11555,N_8731,N_6734);
or U11556 (N_11556,N_7433,N_7825);
and U11557 (N_11557,N_6849,N_6832);
xnor U11558 (N_11558,N_5222,N_5321);
xnor U11559 (N_11559,N_6222,N_9043);
and U11560 (N_11560,N_7253,N_8890);
nor U11561 (N_11561,N_5409,N_9501);
xor U11562 (N_11562,N_7145,N_6580);
or U11563 (N_11563,N_9894,N_8643);
nor U11564 (N_11564,N_7221,N_5374);
nor U11565 (N_11565,N_8660,N_9132);
and U11566 (N_11566,N_7407,N_8402);
and U11567 (N_11567,N_6621,N_8909);
or U11568 (N_11568,N_7934,N_7396);
or U11569 (N_11569,N_8682,N_8579);
and U11570 (N_11570,N_9299,N_6481);
nand U11571 (N_11571,N_6612,N_8728);
and U11572 (N_11572,N_6125,N_5534);
nor U11573 (N_11573,N_8216,N_5978);
and U11574 (N_11574,N_9492,N_5674);
nand U11575 (N_11575,N_6881,N_6190);
nor U11576 (N_11576,N_6790,N_9483);
nand U11577 (N_11577,N_6519,N_6511);
or U11578 (N_11578,N_6858,N_8431);
or U11579 (N_11579,N_8470,N_7906);
or U11580 (N_11580,N_9594,N_5821);
xnor U11581 (N_11581,N_5079,N_9209);
or U11582 (N_11582,N_6840,N_7538);
or U11583 (N_11583,N_8620,N_6967);
nand U11584 (N_11584,N_5025,N_7889);
or U11585 (N_11585,N_6149,N_8972);
or U11586 (N_11586,N_7591,N_7755);
or U11587 (N_11587,N_9241,N_5581);
xor U11588 (N_11588,N_9580,N_9540);
xnor U11589 (N_11589,N_5399,N_8045);
or U11590 (N_11590,N_6208,N_9608);
nand U11591 (N_11591,N_9079,N_5762);
nand U11592 (N_11592,N_6006,N_9778);
and U11593 (N_11593,N_8833,N_8883);
nand U11594 (N_11594,N_5028,N_6239);
or U11595 (N_11595,N_9030,N_9644);
xor U11596 (N_11596,N_9372,N_8098);
xor U11597 (N_11597,N_9737,N_5246);
nand U11598 (N_11598,N_7943,N_6763);
xnor U11599 (N_11599,N_6452,N_6204);
nor U11600 (N_11600,N_8458,N_8420);
nand U11601 (N_11601,N_8062,N_8309);
or U11602 (N_11602,N_7650,N_9285);
nor U11603 (N_11603,N_5296,N_8407);
and U11604 (N_11604,N_5359,N_7780);
and U11605 (N_11605,N_8030,N_7904);
xnor U11606 (N_11606,N_6221,N_9300);
nor U11607 (N_11607,N_9051,N_6807);
nor U11608 (N_11608,N_8466,N_9223);
and U11609 (N_11609,N_8394,N_9550);
or U11610 (N_11610,N_9365,N_7311);
or U11611 (N_11611,N_9454,N_9765);
nand U11612 (N_11612,N_5999,N_5906);
or U11613 (N_11613,N_8523,N_9507);
or U11614 (N_11614,N_7771,N_5067);
xnor U11615 (N_11615,N_9881,N_7421);
nand U11616 (N_11616,N_9197,N_5366);
nand U11617 (N_11617,N_6308,N_6924);
nand U11618 (N_11618,N_5852,N_5622);
nor U11619 (N_11619,N_7152,N_7021);
and U11620 (N_11620,N_8871,N_9909);
nand U11621 (N_11621,N_6689,N_6551);
or U11622 (N_11622,N_5208,N_5094);
or U11623 (N_11623,N_8255,N_6284);
nor U11624 (N_11624,N_7601,N_9092);
nor U11625 (N_11625,N_5675,N_6321);
and U11626 (N_11626,N_9542,N_9663);
xnor U11627 (N_11627,N_6948,N_6092);
or U11628 (N_11628,N_9613,N_7877);
nand U11629 (N_11629,N_8110,N_7299);
xor U11630 (N_11630,N_8937,N_8522);
xor U11631 (N_11631,N_7854,N_7907);
and U11632 (N_11632,N_5599,N_7559);
and U11633 (N_11633,N_8540,N_6837);
nand U11634 (N_11634,N_9012,N_6797);
nand U11635 (N_11635,N_7648,N_5749);
and U11636 (N_11636,N_6859,N_6136);
nor U11637 (N_11637,N_7029,N_9840);
and U11638 (N_11638,N_9509,N_8028);
xnor U11639 (N_11639,N_7858,N_5402);
and U11640 (N_11640,N_6253,N_7350);
xnor U11641 (N_11641,N_7514,N_7256);
or U11642 (N_11642,N_7842,N_6963);
or U11643 (N_11643,N_6275,N_6610);
nand U11644 (N_11644,N_7827,N_5338);
nor U11645 (N_11645,N_6862,N_7908);
nor U11646 (N_11646,N_8263,N_6243);
or U11647 (N_11647,N_7872,N_8664);
nor U11648 (N_11648,N_8104,N_9689);
nor U11649 (N_11649,N_9219,N_9206);
xnor U11650 (N_11650,N_7263,N_7399);
and U11651 (N_11651,N_6200,N_9314);
xnor U11652 (N_11652,N_6543,N_5089);
nor U11653 (N_11653,N_7572,N_9093);
nand U11654 (N_11654,N_7119,N_7061);
nand U11655 (N_11655,N_7079,N_7322);
nand U11656 (N_11656,N_5398,N_5451);
and U11657 (N_11657,N_6705,N_6602);
nand U11658 (N_11658,N_9657,N_9847);
and U11659 (N_11659,N_5642,N_9238);
or U11660 (N_11660,N_8259,N_9410);
and U11661 (N_11661,N_7621,N_8987);
nor U11662 (N_11662,N_5878,N_8349);
and U11663 (N_11663,N_9073,N_6930);
and U11664 (N_11664,N_5044,N_6749);
or U11665 (N_11665,N_8077,N_6803);
nor U11666 (N_11666,N_7624,N_9439);
nand U11667 (N_11667,N_7826,N_9873);
or U11668 (N_11668,N_7087,N_9606);
nand U11669 (N_11669,N_6116,N_5379);
nand U11670 (N_11670,N_5788,N_8878);
or U11671 (N_11671,N_8308,N_7983);
nor U11672 (N_11672,N_9688,N_8668);
or U11673 (N_11673,N_5195,N_7502);
and U11674 (N_11674,N_5422,N_6059);
nand U11675 (N_11675,N_5065,N_9355);
xnor U11676 (N_11676,N_7024,N_5042);
nand U11677 (N_11677,N_8592,N_6349);
nand U11678 (N_11678,N_6690,N_6369);
xnor U11679 (N_11679,N_7699,N_6089);
nand U11680 (N_11680,N_8589,N_6935);
nand U11681 (N_11681,N_6928,N_6035);
nor U11682 (N_11682,N_8189,N_6634);
nor U11683 (N_11683,N_6703,N_5288);
nor U11684 (N_11684,N_8594,N_5045);
and U11685 (N_11685,N_5577,N_5700);
and U11686 (N_11686,N_6723,N_6994);
nor U11687 (N_11687,N_9522,N_6087);
nor U11688 (N_11688,N_9612,N_5407);
xnor U11689 (N_11689,N_8156,N_9638);
nor U11690 (N_11690,N_8294,N_9274);
nand U11691 (N_11691,N_8291,N_8699);
nand U11692 (N_11692,N_5795,N_7279);
nor U11693 (N_11693,N_9723,N_6209);
or U11694 (N_11694,N_5662,N_6086);
nand U11695 (N_11695,N_7819,N_8363);
or U11696 (N_11696,N_7770,N_7807);
or U11697 (N_11697,N_9010,N_9317);
xor U11698 (N_11698,N_8841,N_6446);
nor U11699 (N_11699,N_6203,N_5489);
nor U11700 (N_11700,N_7237,N_6267);
nor U11701 (N_11701,N_8022,N_5650);
nor U11702 (N_11702,N_5652,N_5578);
nor U11703 (N_11703,N_6619,N_7472);
and U11704 (N_11704,N_5513,N_6424);
nor U11705 (N_11705,N_5416,N_6567);
nor U11706 (N_11706,N_9157,N_9015);
xnor U11707 (N_11707,N_7731,N_5905);
nor U11708 (N_11708,N_8918,N_7790);
xor U11709 (N_11709,N_8089,N_6162);
or U11710 (N_11710,N_7733,N_9711);
or U11711 (N_11711,N_7730,N_5125);
nand U11712 (N_11712,N_5509,N_9294);
xnor U11713 (N_11713,N_6561,N_9312);
or U11714 (N_11714,N_8968,N_7093);
xnor U11715 (N_11715,N_8126,N_5829);
nand U11716 (N_11716,N_8475,N_8167);
nor U11717 (N_11717,N_6337,N_6336);
and U11718 (N_11718,N_5080,N_5672);
and U11719 (N_11719,N_6508,N_6295);
nor U11720 (N_11720,N_7323,N_7250);
nand U11721 (N_11721,N_9322,N_6510);
or U11722 (N_11722,N_9768,N_9832);
nor U11723 (N_11723,N_8647,N_8199);
xor U11724 (N_11724,N_8185,N_5013);
or U11725 (N_11725,N_9636,N_5572);
xnor U11726 (N_11726,N_9535,N_8685);
nor U11727 (N_11727,N_9349,N_5984);
and U11728 (N_11728,N_9845,N_6223);
xnor U11729 (N_11729,N_5304,N_8853);
nor U11730 (N_11730,N_5839,N_6040);
and U11731 (N_11731,N_8787,N_8163);
or U11732 (N_11732,N_8182,N_7285);
nand U11733 (N_11733,N_6614,N_6462);
or U11734 (N_11734,N_8429,N_6213);
or U11735 (N_11735,N_5720,N_6828);
nor U11736 (N_11736,N_9874,N_9929);
and U11737 (N_11737,N_9743,N_6100);
nand U11738 (N_11738,N_8065,N_7707);
and U11739 (N_11739,N_5034,N_8606);
nand U11740 (N_11740,N_8683,N_7178);
xor U11741 (N_11741,N_9022,N_8635);
or U11742 (N_11742,N_6688,N_9686);
nor U11743 (N_11743,N_9912,N_7377);
or U11744 (N_11744,N_9109,N_6255);
or U11745 (N_11745,N_7414,N_7455);
or U11746 (N_11746,N_5958,N_9404);
or U11747 (N_11747,N_9690,N_6167);
nand U11748 (N_11748,N_5894,N_9134);
nand U11749 (N_11749,N_7923,N_8241);
or U11750 (N_11750,N_5892,N_9962);
nand U11751 (N_11751,N_8015,N_7890);
xor U11752 (N_11752,N_6279,N_6296);
or U11753 (N_11753,N_8561,N_9629);
or U11754 (N_11754,N_5433,N_7254);
xnor U11755 (N_11755,N_6942,N_9624);
xor U11756 (N_11756,N_8150,N_6278);
nand U11757 (N_11757,N_9667,N_7135);
and U11758 (N_11758,N_7747,N_8434);
nand U11759 (N_11759,N_7663,N_6896);
xor U11760 (N_11760,N_8531,N_9895);
nand U11761 (N_11761,N_7594,N_5357);
and U11762 (N_11762,N_6949,N_7158);
xor U11763 (N_11763,N_8947,N_7018);
nand U11764 (N_11764,N_5507,N_5891);
xor U11765 (N_11765,N_8462,N_9400);
or U11766 (N_11766,N_8715,N_7405);
and U11767 (N_11767,N_8873,N_7717);
xnor U11768 (N_11768,N_7806,N_6188);
nor U11769 (N_11769,N_8085,N_5411);
nor U11770 (N_11770,N_7689,N_6099);
nor U11771 (N_11771,N_7082,N_7108);
or U11772 (N_11772,N_8332,N_8686);
nand U11773 (N_11773,N_9967,N_6482);
or U11774 (N_11774,N_6160,N_8170);
nand U11775 (N_11775,N_8854,N_7345);
nand U11776 (N_11776,N_5964,N_7127);
xor U11777 (N_11777,N_5368,N_6437);
nand U11778 (N_11778,N_5382,N_7337);
and U11779 (N_11779,N_6993,N_5386);
nor U11780 (N_11780,N_8743,N_9548);
nor U11781 (N_11781,N_9732,N_9986);
xor U11782 (N_11782,N_9879,N_8911);
xor U11783 (N_11783,N_9851,N_7150);
nand U11784 (N_11784,N_9648,N_5724);
and U11785 (N_11785,N_9947,N_7013);
xor U11786 (N_11786,N_6033,N_7792);
and U11787 (N_11787,N_9961,N_9802);
nand U11788 (N_11788,N_5394,N_5908);
or U11789 (N_11789,N_5816,N_7622);
or U11790 (N_11790,N_7749,N_7940);
xor U11791 (N_11791,N_8867,N_9551);
nand U11792 (N_11792,N_9745,N_7468);
or U11793 (N_11793,N_7357,N_7761);
nand U11794 (N_11794,N_9389,N_8782);
xor U11795 (N_11795,N_6715,N_8838);
nand U11796 (N_11796,N_5923,N_5982);
nand U11797 (N_11797,N_6987,N_7555);
xor U11798 (N_11798,N_6070,N_7992);
nand U11799 (N_11799,N_6714,N_8256);
nand U11800 (N_11800,N_6650,N_7163);
and U11801 (N_11801,N_7125,N_9708);
or U11802 (N_11802,N_5198,N_9893);
nand U11803 (N_11803,N_7581,N_8985);
nor U11804 (N_11804,N_7166,N_5179);
and U11805 (N_11805,N_8810,N_9448);
nand U11806 (N_11806,N_8847,N_7860);
xor U11807 (N_11807,N_6771,N_5837);
xor U11808 (N_11808,N_7595,N_9003);
nand U11809 (N_11809,N_6118,N_6453);
and U11810 (N_11810,N_5560,N_8131);
nor U11811 (N_11811,N_8819,N_5644);
nor U11812 (N_11812,N_7982,N_5897);
and U11813 (N_11813,N_5845,N_7739);
and U11814 (N_11814,N_5966,N_5643);
nand U11815 (N_11815,N_7048,N_6438);
or U11816 (N_11816,N_6569,N_6440);
or U11817 (N_11817,N_8262,N_5765);
and U11818 (N_11818,N_5289,N_9406);
xor U11819 (N_11819,N_7963,N_8645);
and U11820 (N_11820,N_9869,N_7544);
nand U11821 (N_11821,N_8410,N_9931);
and U11822 (N_11822,N_5009,N_8860);
nand U11823 (N_11823,N_7501,N_8805);
or U11824 (N_11824,N_5008,N_5132);
nand U11825 (N_11825,N_9226,N_6936);
and U11826 (N_11826,N_8359,N_8389);
or U11827 (N_11827,N_5312,N_6575);
xnor U11828 (N_11828,N_9609,N_6730);
and U11829 (N_11829,N_9576,N_6199);
or U11830 (N_11830,N_5810,N_8327);
and U11831 (N_11831,N_7156,N_7641);
xnor U11832 (N_11832,N_9897,N_7664);
nand U11833 (N_11833,N_5159,N_9984);
nand U11834 (N_11834,N_7686,N_5267);
nand U11835 (N_11835,N_9471,N_6998);
nor U11836 (N_11836,N_6365,N_9407);
and U11837 (N_11837,N_6876,N_7274);
or U11838 (N_11838,N_5957,N_9747);
nand U11839 (N_11839,N_5272,N_6432);
and U11840 (N_11840,N_6682,N_5561);
xnor U11841 (N_11841,N_8996,N_8160);
or U11842 (N_11842,N_6036,N_5303);
nor U11843 (N_11843,N_6956,N_8813);
or U11844 (N_11844,N_7161,N_5901);
and U11845 (N_11845,N_6841,N_6112);
nor U11846 (N_11846,N_9586,N_8059);
and U11847 (N_11847,N_9192,N_9038);
nor U11848 (N_11848,N_7801,N_6241);
and U11849 (N_11849,N_6429,N_7131);
nor U11850 (N_11850,N_6132,N_8551);
nand U11851 (N_11851,N_5299,N_6900);
and U11852 (N_11852,N_9939,N_7593);
or U11853 (N_11853,N_9713,N_9905);
nand U11854 (N_11854,N_7543,N_8238);
xnor U11855 (N_11855,N_9855,N_7409);
and U11856 (N_11856,N_8527,N_9216);
nand U11857 (N_11857,N_9480,N_6816);
xor U11858 (N_11858,N_9002,N_9096);
or U11859 (N_11859,N_6671,N_5355);
nand U11860 (N_11860,N_6364,N_5638);
nor U11861 (N_11861,N_9980,N_8694);
nand U11862 (N_11862,N_8733,N_5362);
nand U11863 (N_11863,N_8964,N_6435);
or U11864 (N_11864,N_5435,N_5797);
or U11865 (N_11865,N_6806,N_6802);
nand U11866 (N_11866,N_7324,N_9846);
or U11867 (N_11867,N_9075,N_9004);
nor U11868 (N_11868,N_7703,N_8747);
and U11869 (N_11869,N_7945,N_5460);
xnor U11870 (N_11870,N_9528,N_5052);
xnor U11871 (N_11871,N_6775,N_6352);
nor U11872 (N_11872,N_7565,N_7954);
nor U11873 (N_11873,N_8026,N_5683);
or U11874 (N_11874,N_6371,N_5623);
xor U11875 (N_11875,N_8003,N_7647);
nand U11876 (N_11876,N_9964,N_7692);
or U11877 (N_11877,N_5763,N_5290);
or U11878 (N_11878,N_9475,N_8858);
nand U11879 (N_11879,N_8717,N_5873);
xor U11880 (N_11880,N_7050,N_7319);
nand U11881 (N_11881,N_9416,N_5239);
and U11882 (N_11882,N_5587,N_5988);
xnor U11883 (N_11883,N_6499,N_7241);
xnor U11884 (N_11884,N_8666,N_9946);
and U11885 (N_11885,N_9361,N_9282);
nor U11886 (N_11886,N_7197,N_7262);
nand U11887 (N_11887,N_9333,N_6060);
nor U11888 (N_11888,N_8856,N_8436);
nor U11889 (N_11889,N_6978,N_9099);
nor U11890 (N_11890,N_5328,N_7494);
or U11891 (N_11891,N_7520,N_7482);
nor U11892 (N_11892,N_8614,N_7949);
xor U11893 (N_11893,N_9145,N_6661);
nand U11894 (N_11894,N_8290,N_6153);
nor U11895 (N_11895,N_5874,N_7821);
nand U11896 (N_11896,N_7636,N_6667);
nand U11897 (N_11897,N_9809,N_5128);
or U11898 (N_11898,N_9341,N_8667);
nor U11899 (N_11899,N_7919,N_5752);
nor U11900 (N_11900,N_6944,N_7091);
xnor U11901 (N_11901,N_5468,N_5486);
xnor U11902 (N_11902,N_6075,N_6552);
nor U11903 (N_11903,N_9758,N_9923);
or U11904 (N_11904,N_5041,N_9016);
xnor U11905 (N_11905,N_9924,N_7212);
xor U11906 (N_11906,N_6053,N_7280);
or U11907 (N_11907,N_9457,N_6085);
or U11908 (N_11908,N_9487,N_8079);
xnor U11909 (N_11909,N_7499,N_5826);
or U11910 (N_11910,N_5615,N_7676);
or U11911 (N_11911,N_9619,N_6869);
and U11912 (N_11912,N_7485,N_9158);
nor U11913 (N_11913,N_9982,N_6082);
nand U11914 (N_11914,N_8213,N_7439);
and U11915 (N_11915,N_5190,N_7737);
or U11916 (N_11916,N_5490,N_9761);
nand U11917 (N_11917,N_5131,N_7382);
or U11918 (N_11918,N_8029,N_6933);
xor U11919 (N_11919,N_8198,N_7478);
nand U11920 (N_11920,N_5659,N_8564);
nor U11921 (N_11921,N_9420,N_7775);
and U11922 (N_11922,N_9263,N_5803);
nor U11923 (N_11923,N_7612,N_6048);
nand U11924 (N_11924,N_6796,N_8945);
or U11925 (N_11925,N_7505,N_7713);
or U11926 (N_11926,N_9748,N_9284);
or U11927 (N_11927,N_5585,N_5323);
nand U11928 (N_11928,N_5099,N_9709);
nand U11929 (N_11929,N_9822,N_8042);
nand U11930 (N_11930,N_8677,N_7976);
or U11931 (N_11931,N_9013,N_8080);
xnor U11932 (N_11932,N_8275,N_8496);
nor U11933 (N_11933,N_9070,N_6454);
or U11934 (N_11934,N_7305,N_7643);
nand U11935 (N_11935,N_9649,N_8454);
xnor U11936 (N_11936,N_9969,N_5219);
or U11937 (N_11937,N_8248,N_6418);
nor U11938 (N_11938,N_6319,N_6282);
nand U11939 (N_11939,N_9993,N_5747);
xor U11940 (N_11940,N_8313,N_8149);
nor U11941 (N_11941,N_7335,N_7603);
or U11942 (N_11942,N_8708,N_5480);
and U11943 (N_11943,N_6853,N_5121);
nor U11944 (N_11944,N_9696,N_6251);
and U11945 (N_11945,N_8887,N_9467);
nor U11946 (N_11946,N_6825,N_6892);
nand U11947 (N_11947,N_7705,N_6117);
nor U11948 (N_11948,N_5343,N_6008);
nand U11949 (N_11949,N_9306,N_6611);
xnor U11950 (N_11950,N_8773,N_5528);
and U11951 (N_11951,N_9195,N_8631);
nand U11952 (N_11952,N_6156,N_5353);
xor U11953 (N_11953,N_7033,N_9362);
nor U11954 (N_11954,N_6895,N_9376);
nand U11955 (N_11955,N_5776,N_5544);
nor U11956 (N_11956,N_8618,N_6835);
nand U11957 (N_11957,N_8893,N_6120);
nand U11958 (N_11958,N_5824,N_5719);
nor U11959 (N_11959,N_8806,N_7037);
and U11960 (N_11960,N_5848,N_5365);
and U11961 (N_11961,N_9755,N_9625);
xnor U11962 (N_11962,N_7833,N_5898);
and U11963 (N_11963,N_5153,N_7837);
nor U11964 (N_11964,N_9423,N_8922);
or U11965 (N_11965,N_8578,N_8477);
nand U11966 (N_11966,N_8933,N_5070);
or U11967 (N_11967,N_8554,N_8073);
or U11968 (N_11968,N_9674,N_9135);
nand U11969 (N_11969,N_8995,N_5104);
nor U11970 (N_11970,N_6712,N_6270);
xnor U11971 (N_11971,N_8322,N_7511);
xnor U11972 (N_11972,N_6477,N_5108);
xor U11973 (N_11973,N_5164,N_6821);
nand U11974 (N_11974,N_5569,N_7313);
or U11975 (N_11975,N_5808,N_7840);
and U11976 (N_11976,N_8038,N_9449);
or U11977 (N_11977,N_5278,N_9278);
xnor U11978 (N_11978,N_5146,N_6970);
and U11979 (N_11979,N_6958,N_9050);
and U11980 (N_11980,N_8449,N_5789);
xor U11981 (N_11981,N_8033,N_5838);
xnor U11982 (N_11982,N_8509,N_5954);
and U11983 (N_11983,N_7690,N_5335);
and U11984 (N_11984,N_8271,N_9418);
or U11985 (N_11985,N_8384,N_6875);
nor U11986 (N_11986,N_6955,N_8428);
nand U11987 (N_11987,N_6573,N_6512);
and U11988 (N_11988,N_9770,N_8426);
or U11989 (N_11989,N_9868,N_8921);
nor U11990 (N_11990,N_9622,N_9236);
nor U11991 (N_11991,N_7691,N_7245);
xnor U11992 (N_11992,N_9089,N_7027);
nand U11993 (N_11993,N_6032,N_9280);
or U11994 (N_11994,N_9460,N_5704);
nand U11995 (N_11995,N_9639,N_5730);
and U11996 (N_11996,N_8372,N_7561);
nand U11997 (N_11997,N_6066,N_9516);
xor U11998 (N_11998,N_7476,N_7646);
nand U11999 (N_11999,N_7996,N_8832);
or U12000 (N_12000,N_7743,N_7067);
and U12001 (N_12001,N_9008,N_8510);
or U12002 (N_12002,N_6864,N_7442);
nor U12003 (N_12003,N_6633,N_5373);
nand U12004 (N_12004,N_6792,N_9194);
nand U12005 (N_12005,N_6904,N_5016);
or U12006 (N_12006,N_8486,N_8954);
nand U12007 (N_12007,N_8678,N_7961);
and U12008 (N_12008,N_9792,N_9491);
or U12009 (N_12009,N_6805,N_7704);
and U12010 (N_12010,N_9906,N_8307);
or U12011 (N_12011,N_8463,N_7107);
and U12012 (N_12012,N_8054,N_9393);
or U12013 (N_12013,N_7415,N_9443);
and U12014 (N_12014,N_7074,N_9843);
nand U12015 (N_12015,N_7440,N_8320);
xnor U12016 (N_12016,N_9243,N_8957);
nand U12017 (N_12017,N_8268,N_9201);
nor U12018 (N_12018,N_9259,N_9798);
xnor U12019 (N_12019,N_6831,N_5248);
or U12020 (N_12020,N_6898,N_9650);
and U12021 (N_12021,N_5828,N_9992);
and U12022 (N_12022,N_5439,N_9391);
and U12023 (N_12023,N_6158,N_6142);
and U12024 (N_12024,N_6285,N_8146);
or U12025 (N_12025,N_7868,N_7392);
xor U12026 (N_12026,N_9597,N_5151);
and U12027 (N_12027,N_9222,N_9470);
nand U12028 (N_12028,N_5879,N_7329);
xor U12029 (N_12029,N_5496,N_8209);
nand U12030 (N_12030,N_8886,N_7260);
xor U12031 (N_12031,N_9938,N_6911);
nand U12032 (N_12032,N_8124,N_9196);
and U12033 (N_12033,N_5986,N_7406);
nor U12034 (N_12034,N_5307,N_7903);
and U12035 (N_12035,N_7564,N_5807);
xor U12036 (N_12036,N_9125,N_7985);
xnor U12037 (N_12037,N_5514,N_6863);
or U12038 (N_12038,N_5805,N_9169);
and U12039 (N_12039,N_7970,N_6037);
nand U12040 (N_12040,N_9108,N_9421);
nand U12041 (N_12041,N_9806,N_5786);
or U12042 (N_12042,N_7964,N_7708);
nand U12043 (N_12043,N_6005,N_7623);
or U12044 (N_12044,N_6798,N_6064);
and U12045 (N_12045,N_6119,N_6839);
or U12046 (N_12046,N_6309,N_5361);
nand U12047 (N_12047,N_9863,N_6390);
nand U12048 (N_12048,N_5410,N_6788);
nand U12049 (N_12049,N_7823,N_6537);
nand U12050 (N_12050,N_9623,N_9692);
nor U12051 (N_12051,N_7474,N_8793);
nand U12052 (N_12052,N_5233,N_8125);
xnor U12053 (N_12053,N_6246,N_7432);
nand U12054 (N_12054,N_5503,N_7562);
nand U12055 (N_12055,N_7637,N_6566);
nor U12056 (N_12056,N_9006,N_8250);
xnor U12057 (N_12057,N_7969,N_9279);
nor U12058 (N_12058,N_8615,N_9212);
and U12059 (N_12059,N_9493,N_8792);
or U12060 (N_12060,N_9155,N_8043);
xor U12061 (N_12061,N_7787,N_9557);
nor U12062 (N_12062,N_5448,N_7569);
or U12063 (N_12063,N_7017,N_9271);
nor U12064 (N_12064,N_8251,N_9565);
xor U12065 (N_12065,N_7883,N_5048);
or U12066 (N_12066,N_5636,N_9995);
nand U12067 (N_12067,N_9682,N_7122);
and U12068 (N_12068,N_8117,N_6434);
nand U12069 (N_12069,N_5163,N_7625);
and U12070 (N_12070,N_6851,N_6550);
and U12071 (N_12071,N_9957,N_9080);
nor U12072 (N_12072,N_5018,N_7249);
or U12073 (N_12073,N_9232,N_9334);
nand U12074 (N_12074,N_7893,N_5320);
or U12075 (N_12075,N_5820,N_7475);
and U12076 (N_12076,N_6727,N_9027);
xor U12077 (N_12077,N_9764,N_8319);
nand U12078 (N_12078,N_7205,N_8339);
and U12079 (N_12079,N_5936,N_7155);
and U12080 (N_12080,N_7270,N_6384);
nor U12081 (N_12081,N_5755,N_7020);
and U12082 (N_12082,N_5183,N_8324);
and U12083 (N_12083,N_9082,N_5428);
xor U12084 (N_12084,N_5606,N_6843);
or U12085 (N_12085,N_9276,N_5012);
nand U12086 (N_12086,N_5220,N_7293);
nor U12087 (N_12087,N_5015,N_7294);
nand U12088 (N_12088,N_9461,N_7786);
nand U12089 (N_12089,N_9788,N_7937);
xor U12090 (N_12090,N_5024,N_7361);
and U12091 (N_12091,N_5447,N_9738);
xnor U12092 (N_12092,N_5297,N_8208);
and U12093 (N_12093,N_7815,N_8134);
nor U12094 (N_12094,N_6764,N_6280);
xor U12095 (N_12095,N_5261,N_6110);
nand U12096 (N_12096,N_9952,N_6617);
nor U12097 (N_12097,N_7534,N_9590);
and U12098 (N_12098,N_8066,N_7783);
nor U12099 (N_12099,N_8546,N_6868);
nand U12100 (N_12100,N_5268,N_8927);
nand U12101 (N_12101,N_6134,N_9900);
or U12102 (N_12102,N_7316,N_6487);
and U12103 (N_12103,N_5397,N_6101);
and U12104 (N_12104,N_8500,N_5032);
nor U12105 (N_12105,N_6546,N_5358);
or U12106 (N_12106,N_8382,N_8084);
xor U12107 (N_12107,N_5169,N_5354);
xnor U12108 (N_12108,N_9242,N_8049);
xor U12109 (N_12109,N_6940,N_9828);
and U12110 (N_12110,N_9853,N_6307);
or U12111 (N_12111,N_6645,N_8502);
xor U12112 (N_12112,N_9056,N_9666);
xnor U12113 (N_12113,N_5673,N_7297);
nor U12114 (N_12114,N_7905,N_7179);
nor U12115 (N_12115,N_5178,N_5174);
xor U12116 (N_12116,N_5091,N_5782);
nand U12117 (N_12117,N_8388,N_9123);
nand U12118 (N_12118,N_9671,N_9701);
nand U12119 (N_12119,N_9390,N_9932);
and U12120 (N_12120,N_6043,N_7312);
nor U12121 (N_12121,N_9250,N_6177);
xor U12122 (N_12122,N_6313,N_5184);
nor U12123 (N_12123,N_7670,N_7344);
or U12124 (N_12124,N_8979,N_6683);
or U12125 (N_12125,N_5217,N_9598);
nand U12126 (N_12126,N_6938,N_7566);
nor U12127 (N_12127,N_9117,N_5664);
nand U12128 (N_12128,N_5922,N_5951);
nor U12129 (N_12129,N_6751,N_6801);
and U12130 (N_12130,N_7180,N_7995);
nand U12131 (N_12131,N_6854,N_8652);
nor U12132 (N_12132,N_9670,N_8494);
xnor U12133 (N_12133,N_8761,N_6996);
or U12134 (N_12134,N_8574,N_9462);
and U12135 (N_12135,N_9455,N_7371);
xnor U12136 (N_12136,N_7633,N_6648);
xor U12137 (N_12137,N_7590,N_9283);
nand U12138 (N_12138,N_8206,N_5438);
or U12139 (N_12139,N_8634,N_9258);
xnor U12140 (N_12140,N_7513,N_8706);
and U12141 (N_12141,N_9330,N_6770);
nand U12142 (N_12142,N_7452,N_8173);
nand U12143 (N_12143,N_7605,N_8504);
or U12144 (N_12144,N_8612,N_8479);
and U12145 (N_12145,N_9343,N_8174);
nor U12146 (N_12146,N_9954,N_7758);
nor U12147 (N_12147,N_9151,N_9469);
and U12148 (N_12148,N_8164,N_8106);
nor U12149 (N_12149,N_5367,N_6643);
nor U12150 (N_12150,N_7635,N_5333);
or U12151 (N_12151,N_6629,N_9063);
xnor U12152 (N_12152,N_5093,N_6576);
or U12153 (N_12153,N_9069,N_8040);
or U12154 (N_12154,N_6427,N_8270);
nor U12155 (N_12155,N_5919,N_7327);
xor U12156 (N_12156,N_7142,N_6962);
nor U12157 (N_12157,N_7885,N_7960);
or U12158 (N_12158,N_9077,N_5187);
and U12159 (N_12159,N_5346,N_5753);
or U12160 (N_12160,N_9202,N_7092);
and U12161 (N_12161,N_8005,N_8387);
and U12162 (N_12162,N_5971,N_7192);
xor U12163 (N_12163,N_5685,N_7134);
or U12164 (N_12164,N_9187,N_7078);
xnor U12165 (N_12165,N_6376,N_5455);
or U12166 (N_12166,N_5616,N_5167);
and U12167 (N_12167,N_7745,N_7104);
nor U12168 (N_12168,N_9098,N_5512);
nand U12169 (N_12169,N_9927,N_9005);
nand U12170 (N_12170,N_9759,N_6346);
xnor U12171 (N_12171,N_7425,N_5992);
xor U12172 (N_12172,N_9518,N_6359);
or U12173 (N_12173,N_9564,N_5748);
nor U12174 (N_12174,N_9556,N_7351);
nand U12175 (N_12175,N_6474,N_8986);
xnor U12176 (N_12176,N_9605,N_9128);
xnor U12177 (N_12177,N_5155,N_5593);
and U12178 (N_12178,N_5253,N_6984);
xor U12179 (N_12179,N_6972,N_5563);
xnor U12180 (N_12180,N_5537,N_9953);
and U12181 (N_12181,N_6615,N_8924);
or U12182 (N_12182,N_8640,N_8264);
and U12183 (N_12183,N_7190,N_7834);
nor U12184 (N_12184,N_5713,N_5115);
or U12185 (N_12185,N_7438,N_7043);
nor U12186 (N_12186,N_9062,N_5395);
or U12187 (N_12187,N_9289,N_8194);
and U12188 (N_12188,N_5081,N_7778);
xnor U12189 (N_12189,N_9537,N_8765);
xnor U12190 (N_12190,N_9066,N_8468);
and U12191 (N_12191,N_6090,N_6265);
and U12192 (N_12192,N_8024,N_8391);
or U12193 (N_12193,N_9147,N_6544);
xor U12194 (N_12194,N_7126,N_7575);
nand U12195 (N_12195,N_9350,N_6042);
xor U12196 (N_12196,N_5021,N_6818);
nor U12197 (N_12197,N_5287,N_6327);
xor U12198 (N_12198,N_6680,N_8474);
nor U12199 (N_12199,N_9672,N_8807);
xor U12200 (N_12200,N_7848,N_6969);
and U12201 (N_12201,N_7195,N_8904);
or U12202 (N_12202,N_9781,N_7656);
nand U12203 (N_12203,N_6997,N_7064);
xnor U12204 (N_12204,N_6214,N_9864);
xnor U12205 (N_12205,N_7894,N_9402);
nor U12206 (N_12206,N_6590,N_8115);
xor U12207 (N_12207,N_8701,N_7051);
xor U12208 (N_12208,N_8226,N_7500);
xor U12209 (N_12209,N_7654,N_8303);
nor U12210 (N_12210,N_6759,N_7346);
or U12211 (N_12211,N_7938,N_5617);
nor U12212 (N_12212,N_7864,N_9199);
nand U12213 (N_12213,N_8230,N_8936);
nand U12214 (N_12214,N_9719,N_5339);
nor U12215 (N_12215,N_6169,N_6263);
nand U12216 (N_12216,N_8456,N_7244);
nor U12217 (N_12217,N_6980,N_8545);
nand U12218 (N_12218,N_6113,N_7850);
nor U12219 (N_12219,N_7121,N_9065);
and U12220 (N_12220,N_8371,N_6148);
nor U12221 (N_12221,N_9466,N_7698);
xnor U12222 (N_12222,N_5256,N_7224);
and U12223 (N_12223,N_5472,N_5141);
xnor U12224 (N_12224,N_7348,N_6186);
nand U12225 (N_12225,N_8177,N_8827);
or U12226 (N_12226,N_7927,N_6522);
xnor U12227 (N_12227,N_9324,N_6894);
nand U12228 (N_12228,N_7010,N_5802);
xor U12229 (N_12229,N_9237,N_6973);
or U12230 (N_12230,N_6676,N_8224);
nor U12231 (N_12231,N_5156,N_8377);
nor U12232 (N_12232,N_7194,N_5759);
nor U12233 (N_12233,N_8744,N_9785);
xor U12234 (N_12234,N_7207,N_7477);
nand U12235 (N_12235,N_7724,N_6224);
xor U12236 (N_12236,N_5692,N_9602);
or U12237 (N_12237,N_5841,N_7764);
or U12238 (N_12238,N_5645,N_9861);
nand U12239 (N_12239,N_6283,N_9290);
xnor U12240 (N_12240,N_7853,N_6918);
and U12241 (N_12241,N_8506,N_5663);
xor U12242 (N_12242,N_8669,N_8439);
and U12243 (N_12243,N_9744,N_5203);
nor U12244 (N_12244,N_5459,N_9949);
or U12245 (N_12245,N_5259,N_6377);
or U12246 (N_12246,N_9566,N_9338);
nor U12247 (N_12247,N_5313,N_5378);
nand U12248 (N_12248,N_9794,N_8366);
and U12249 (N_12249,N_5393,N_6281);
nand U12250 (N_12250,N_5102,N_5562);
nand U12251 (N_12251,N_9042,N_5844);
nand U12252 (N_12252,N_8749,N_8769);
xnor U12253 (N_12253,N_9742,N_6766);
nand U12254 (N_12254,N_6163,N_7629);
xnor U12255 (N_12255,N_5945,N_5130);
or U12256 (N_12256,N_5523,N_8069);
or U12257 (N_12257,N_8905,N_6227);
and U12258 (N_12258,N_9994,N_7054);
nand U12259 (N_12259,N_5069,N_5095);
nor U12260 (N_12260,N_9917,N_9172);
nand U12261 (N_12261,N_6459,N_7966);
nand U12262 (N_12262,N_6500,N_8534);
xor U12263 (N_12263,N_7812,N_6044);
xor U12264 (N_12264,N_8154,N_8962);
or U12265 (N_12265,N_8770,N_6356);
nor U12266 (N_12266,N_5006,N_6171);
and U12267 (N_12267,N_5974,N_6324);
and U12268 (N_12268,N_6450,N_7236);
xor U12269 (N_12269,N_6245,N_9139);
and U12270 (N_12270,N_9392,N_9320);
nor U12271 (N_12271,N_8602,N_7271);
nor U12272 (N_12272,N_9499,N_8759);
or U12273 (N_12273,N_6212,N_5162);
nor U12274 (N_12274,N_9085,N_7673);
or U12275 (N_12275,N_7578,N_5705);
xor U12276 (N_12276,N_6330,N_8881);
nor U12277 (N_12277,N_5252,N_7503);
or U12278 (N_12278,N_6133,N_8070);
and U12279 (N_12279,N_9047,N_9763);
nor U12280 (N_12280,N_8408,N_6883);
and U12281 (N_12281,N_5414,N_9974);
xor U12282 (N_12282,N_9996,N_5761);
xnor U12283 (N_12283,N_7710,N_5680);
nor U12284 (N_12284,N_8076,N_5005);
nor U12285 (N_12285,N_8948,N_8519);
xnor U12286 (N_12286,N_8016,N_9634);
or U12287 (N_12287,N_5254,N_7596);
and U12288 (N_12288,N_5060,N_7012);
and U12289 (N_12289,N_7693,N_6478);
or U12290 (N_12290,N_7509,N_8276);
nor U12291 (N_12291,N_9703,N_7203);
and U12292 (N_12292,N_5694,N_5137);
nor U12293 (N_12293,N_9160,N_6181);
and U12294 (N_12294,N_8265,N_9210);
xnor U12295 (N_12295,N_9427,N_9124);
nand U12296 (N_12296,N_5173,N_8914);
and U12297 (N_12297,N_8577,N_7523);
xor U12298 (N_12298,N_9727,N_6009);
nand U12299 (N_12299,N_6266,N_5671);
nor U12300 (N_12300,N_9369,N_7049);
nand U12301 (N_12301,N_7608,N_7779);
nand U12302 (N_12302,N_9064,N_5337);
nand U12303 (N_12303,N_6104,N_9302);
or U12304 (N_12304,N_7882,N_7071);
xor U12305 (N_12305,N_5188,N_6654);
nand U12306 (N_12306,N_8788,N_6027);
or U12307 (N_12307,N_8179,N_8980);
and U12308 (N_12308,N_6097,N_6436);
or U12309 (N_12309,N_7898,N_6966);
nand U12310 (N_12310,N_8582,N_6596);
nor U12311 (N_12311,N_8318,N_9011);
xnor U12312 (N_12312,N_7805,N_9175);
nand U12313 (N_12313,N_6559,N_9876);
and U12314 (N_12314,N_8442,N_5516);
and U12315 (N_12315,N_8266,N_5764);
nand U12316 (N_12316,N_6762,N_9838);
xor U12317 (N_12317,N_7320,N_6932);
or U12318 (N_12318,N_7075,N_6728);
nor U12319 (N_12319,N_8843,N_5092);
xor U12320 (N_12320,N_9729,N_5450);
or U12321 (N_12321,N_6252,N_7695);
and U12322 (N_12322,N_5924,N_7381);
nand U12323 (N_12323,N_8974,N_8734);
xnor U12324 (N_12324,N_8872,N_6135);
or U12325 (N_12325,N_8851,N_5727);
and U12326 (N_12326,N_9808,N_8809);
nand U12327 (N_12327,N_6225,N_5831);
nor U12328 (N_12328,N_6000,N_6850);
xor U12329 (N_12329,N_9819,N_7816);
or U12330 (N_12330,N_6031,N_9915);
or U12331 (N_12331,N_8437,N_7276);
nand U12332 (N_12332,N_5226,N_6833);
nor U12333 (N_12333,N_6845,N_8075);
or U12334 (N_12334,N_8829,N_8989);
or U12335 (N_12335,N_6521,N_6601);
xor U12336 (N_12336,N_9325,N_7005);
nand U12337 (N_12337,N_5792,N_7034);
nor U12338 (N_12338,N_7380,N_7384);
and U12339 (N_12339,N_9640,N_8101);
and U12340 (N_12340,N_7264,N_6047);
nand U12341 (N_12341,N_9498,N_9328);
and U12342 (N_12342,N_8868,N_6685);
nor U12343 (N_12343,N_7103,N_7526);
or U12344 (N_12344,N_7359,N_6809);
and U12345 (N_12345,N_8720,N_9691);
xor U12346 (N_12346,N_6999,N_5854);
or U12347 (N_12347,N_6658,N_5470);
xor U12348 (N_12348,N_8277,N_6565);
and U12349 (N_12349,N_8955,N_5494);
and U12350 (N_12350,N_9217,N_8286);
xnor U12351 (N_12351,N_9678,N_9234);
or U12352 (N_12352,N_6422,N_6328);
nand U12353 (N_12353,N_5237,N_5979);
and U12354 (N_12354,N_7084,N_9433);
and U12355 (N_12355,N_6916,N_7138);
and U12356 (N_12356,N_8121,N_6439);
nand U12357 (N_12357,N_8009,N_5942);
nor U12358 (N_12358,N_9009,N_9348);
or U12359 (N_12359,N_6139,N_7445);
or U12360 (N_12360,N_8850,N_8576);
nand U12361 (N_12361,N_9039,N_7417);
xor U12362 (N_12362,N_7661,N_9296);
nor U12363 (N_12363,N_7214,N_9544);
or U12364 (N_12364,N_6448,N_6395);
or U12365 (N_12365,N_5375,N_8071);
xnor U12366 (N_12366,N_8133,N_5798);
or U12367 (N_12367,N_6473,N_7955);
and U12368 (N_12368,N_5774,N_5401);
nor U12369 (N_12369,N_5657,N_5698);
or U12370 (N_12370,N_8348,N_9654);
and U12371 (N_12371,N_9154,N_9224);
xnor U12372 (N_12372,N_6479,N_5541);
or U12373 (N_12373,N_6915,N_8433);
and U12374 (N_12374,N_7014,N_6782);
xnor U12375 (N_12375,N_8006,N_6496);
and U12376 (N_12376,N_7362,N_5801);
and U12377 (N_12377,N_6979,N_9208);
xor U12378 (N_12378,N_7370,N_8376);
nor U12379 (N_12379,N_7814,N_6159);
or U12380 (N_12380,N_8187,N_9841);
nor U12381 (N_12381,N_8961,N_5862);
nor U12382 (N_12382,N_8292,N_9928);
or U12383 (N_12383,N_7317,N_5612);
and U12384 (N_12384,N_5875,N_9121);
nand U12385 (N_12385,N_5937,N_8218);
xnor U12386 (N_12386,N_5661,N_6538);
nor U12387 (N_12387,N_6257,N_6193);
and U12388 (N_12388,N_9658,N_6757);
or U12389 (N_12389,N_5113,N_5107);
or U12390 (N_12390,N_6909,N_8525);
nand U12391 (N_12391,N_9587,N_6555);
and U12392 (N_12392,N_8520,N_9651);
nand U12393 (N_12393,N_8656,N_9908);
and U12394 (N_12394,N_8315,N_6095);
xnor U12395 (N_12395,N_6466,N_8663);
or U12396 (N_12396,N_9331,N_9465);
xor U12397 (N_12397,N_8472,N_6187);
nor U12398 (N_12398,N_7193,N_5847);
xnor U12399 (N_12399,N_6532,N_9575);
nor U12400 (N_12400,N_5858,N_5517);
nand U12401 (N_12401,N_8352,N_9353);
or U12402 (N_12402,N_8143,N_6745);
or U12403 (N_12403,N_6824,N_9710);
or U12404 (N_12404,N_6760,N_9384);
or U12405 (N_12405,N_6719,N_5670);
nand U12406 (N_12406,N_9408,N_8575);
and U12407 (N_12407,N_5866,N_9291);
nor U12408 (N_12408,N_6091,N_6250);
nor U12409 (N_12409,N_5504,N_5539);
or U12410 (N_12410,N_7808,N_7754);
nand U12411 (N_12411,N_5348,N_9426);
nand U12412 (N_12412,N_6599,N_6572);
nor U12413 (N_12413,N_6901,N_8067);
nand U12414 (N_12414,N_5002,N_6025);
or U12415 (N_12415,N_5023,N_9474);
xor U12416 (N_12416,N_5529,N_6668);
nor U12417 (N_12417,N_5559,N_6871);
nor U12418 (N_12418,N_8869,N_9538);
and U12419 (N_12419,N_7114,N_5947);
nand U12420 (N_12420,N_7716,N_8760);
nand U12421 (N_12421,N_6746,N_5609);
nand U12422 (N_12422,N_5200,N_5385);
and U12423 (N_12423,N_8017,N_8274);
xnor U12424 (N_12424,N_5264,N_6903);
nand U12425 (N_12425,N_7640,N_5148);
nor U12426 (N_12426,N_6174,N_5743);
xnor U12427 (N_12427,N_8413,N_5210);
nor U12428 (N_12428,N_6150,N_8616);
and U12429 (N_12429,N_8690,N_7003);
and U12430 (N_12430,N_5154,N_8704);
nand U12431 (N_12431,N_5546,N_5629);
nand U12432 (N_12432,N_9578,N_7917);
nand U12433 (N_12433,N_8353,N_5457);
xor U12434 (N_12434,N_5532,N_9724);
or U12435 (N_12435,N_7235,N_6238);
or U12436 (N_12436,N_5625,N_6362);
nand U12437 (N_12437,N_9656,N_8786);
nand U12438 (N_12438,N_5049,N_7800);
and U12439 (N_12439,N_5766,N_7824);
xnor U12440 (N_12440,N_7435,N_9630);
nor U12441 (N_12441,N_5305,N_7105);
and U12442 (N_12442,N_5930,N_6375);
or U12443 (N_12443,N_9401,N_6237);
nor U12444 (N_12444,N_7537,N_9571);
xnor U12445 (N_12445,N_9589,N_7412);
nor U12446 (N_12446,N_6753,N_7364);
nor U12447 (N_12447,N_9856,N_8107);
xor U12448 (N_12448,N_7542,N_5718);
nor U12449 (N_12449,N_8139,N_9716);
nor U12450 (N_12450,N_7315,N_7602);
xor U12451 (N_12451,N_8726,N_7040);
xor U12452 (N_12452,N_8365,N_7202);
nor U12453 (N_12453,N_5576,N_8533);
xnor U12454 (N_12454,N_5318,N_6726);
nor U12455 (N_12455,N_6657,N_9203);
nor U12456 (N_12456,N_9335,N_9837);
and U12457 (N_12457,N_9083,N_6378);
nand U12458 (N_12458,N_5266,N_9611);
nor U12459 (N_12459,N_7446,N_6345);
nor U12460 (N_12460,N_6700,N_9524);
xor U12461 (N_12461,N_7496,N_5238);
or U12462 (N_12462,N_9115,N_6490);
and U12463 (N_12463,N_8158,N_7672);
nor U12464 (N_12464,N_9680,N_8438);
or U12465 (N_12465,N_5432,N_5223);
and U12466 (N_12466,N_9635,N_9494);
nand U12467 (N_12467,N_5157,N_6525);
xnor U12468 (N_12468,N_6414,N_6096);
xnor U12469 (N_12469,N_8791,N_9536);
nor U12470 (N_12470,N_6758,N_8037);
nand U12471 (N_12471,N_6738,N_7148);
and U12472 (N_12472,N_5646,N_5649);
xnor U12473 (N_12473,N_8767,N_7838);
nor U12474 (N_12474,N_6045,N_5129);
nor U12475 (N_12475,N_6557,N_6172);
or U12476 (N_12476,N_9185,N_6826);
nor U12477 (N_12477,N_8624,N_6412);
or U12478 (N_12478,N_7721,N_8548);
or U12479 (N_12479,N_9205,N_6513);
or U12480 (N_12480,N_8118,N_5610);
xnor U12481 (N_12481,N_9829,N_6624);
nand U12482 (N_12482,N_9714,N_5916);
nor U12483 (N_12483,N_6183,N_6982);
nand U12484 (N_12484,N_9326,N_7918);
or U12485 (N_12485,N_8330,N_7706);
nand U12486 (N_12486,N_6594,N_8935);
nor U12487 (N_12487,N_5158,N_7336);
or U12488 (N_12488,N_7895,N_7349);
or U12489 (N_12489,N_5466,N_8461);
nand U12490 (N_12490,N_6122,N_7111);
or U12491 (N_12491,N_5723,N_8776);
xor U12492 (N_12492,N_6501,N_9554);
and U12493 (N_12493,N_9926,N_9183);
and U12494 (N_12494,N_8932,N_5518);
and U12495 (N_12495,N_5412,N_7539);
nand U12496 (N_12496,N_7811,N_9811);
nand U12497 (N_12497,N_9561,N_5427);
nand U12498 (N_12498,N_8639,N_9796);
nor U12499 (N_12499,N_5648,N_5861);
xnor U12500 (N_12500,N_7189,N_8884);
nor U12501 (N_12501,N_9098,N_7306);
nand U12502 (N_12502,N_7615,N_5302);
and U12503 (N_12503,N_5100,N_5296);
nor U12504 (N_12504,N_5406,N_6629);
nor U12505 (N_12505,N_5112,N_9744);
or U12506 (N_12506,N_6164,N_8238);
nor U12507 (N_12507,N_8638,N_9592);
xnor U12508 (N_12508,N_9951,N_7825);
nor U12509 (N_12509,N_7340,N_9775);
nand U12510 (N_12510,N_9294,N_5182);
or U12511 (N_12511,N_9284,N_8909);
nand U12512 (N_12512,N_6211,N_8225);
nor U12513 (N_12513,N_9808,N_9500);
xnor U12514 (N_12514,N_9862,N_7168);
and U12515 (N_12515,N_5828,N_5577);
nor U12516 (N_12516,N_9495,N_8203);
or U12517 (N_12517,N_9380,N_9575);
or U12518 (N_12518,N_6337,N_9594);
and U12519 (N_12519,N_8622,N_5822);
or U12520 (N_12520,N_9183,N_8508);
nand U12521 (N_12521,N_7319,N_6071);
or U12522 (N_12522,N_6954,N_6598);
xnor U12523 (N_12523,N_8431,N_8695);
and U12524 (N_12524,N_5363,N_5631);
nand U12525 (N_12525,N_6216,N_6019);
or U12526 (N_12526,N_8175,N_9040);
and U12527 (N_12527,N_7875,N_8066);
and U12528 (N_12528,N_7069,N_9016);
or U12529 (N_12529,N_9740,N_9593);
and U12530 (N_12530,N_5895,N_5001);
xor U12531 (N_12531,N_9534,N_9867);
nor U12532 (N_12532,N_5761,N_9364);
and U12533 (N_12533,N_5402,N_8738);
nand U12534 (N_12534,N_6086,N_9942);
xnor U12535 (N_12535,N_5948,N_5687);
xor U12536 (N_12536,N_9978,N_7989);
or U12537 (N_12537,N_7798,N_8444);
nor U12538 (N_12538,N_6472,N_8346);
or U12539 (N_12539,N_6834,N_6097);
nor U12540 (N_12540,N_8734,N_6189);
nor U12541 (N_12541,N_8365,N_8720);
nand U12542 (N_12542,N_7036,N_5659);
xor U12543 (N_12543,N_9038,N_5754);
nor U12544 (N_12544,N_9932,N_7083);
nand U12545 (N_12545,N_6566,N_8516);
or U12546 (N_12546,N_7271,N_9861);
or U12547 (N_12547,N_7998,N_7069);
nor U12548 (N_12548,N_9561,N_8030);
or U12549 (N_12549,N_8542,N_7876);
and U12550 (N_12550,N_5024,N_8320);
or U12551 (N_12551,N_5931,N_5017);
or U12552 (N_12552,N_5782,N_9848);
xnor U12553 (N_12553,N_9504,N_5835);
and U12554 (N_12554,N_9285,N_5864);
xnor U12555 (N_12555,N_7442,N_6079);
nand U12556 (N_12556,N_6564,N_7298);
nor U12557 (N_12557,N_8414,N_8518);
and U12558 (N_12558,N_6777,N_7575);
xor U12559 (N_12559,N_5743,N_7004);
and U12560 (N_12560,N_9596,N_7789);
or U12561 (N_12561,N_7734,N_5179);
xnor U12562 (N_12562,N_5638,N_9523);
nand U12563 (N_12563,N_8898,N_9322);
and U12564 (N_12564,N_6440,N_7072);
nand U12565 (N_12565,N_6263,N_7288);
and U12566 (N_12566,N_6506,N_9722);
nand U12567 (N_12567,N_7359,N_6754);
or U12568 (N_12568,N_8845,N_8877);
nand U12569 (N_12569,N_5034,N_9180);
xor U12570 (N_12570,N_6153,N_5391);
nor U12571 (N_12571,N_5958,N_6296);
and U12572 (N_12572,N_9868,N_6677);
nand U12573 (N_12573,N_6050,N_9714);
nor U12574 (N_12574,N_8270,N_8145);
nand U12575 (N_12575,N_9320,N_9639);
nand U12576 (N_12576,N_9069,N_8851);
or U12577 (N_12577,N_7174,N_9974);
or U12578 (N_12578,N_5832,N_7286);
and U12579 (N_12579,N_5329,N_6009);
nor U12580 (N_12580,N_9159,N_6510);
and U12581 (N_12581,N_9342,N_5963);
nor U12582 (N_12582,N_6139,N_8543);
or U12583 (N_12583,N_9211,N_8533);
xnor U12584 (N_12584,N_5464,N_5487);
or U12585 (N_12585,N_6152,N_5238);
nand U12586 (N_12586,N_5061,N_5387);
and U12587 (N_12587,N_7125,N_9711);
or U12588 (N_12588,N_6302,N_6327);
xor U12589 (N_12589,N_8441,N_5672);
nand U12590 (N_12590,N_5690,N_5227);
nand U12591 (N_12591,N_7673,N_7042);
xor U12592 (N_12592,N_5600,N_8746);
xor U12593 (N_12593,N_6607,N_6881);
xnor U12594 (N_12594,N_8290,N_6730);
nor U12595 (N_12595,N_8494,N_7540);
and U12596 (N_12596,N_8901,N_7393);
nor U12597 (N_12597,N_6532,N_7091);
or U12598 (N_12598,N_9915,N_9558);
xnor U12599 (N_12599,N_8940,N_6570);
and U12600 (N_12600,N_8719,N_5816);
nand U12601 (N_12601,N_5365,N_9899);
nor U12602 (N_12602,N_6810,N_8376);
nand U12603 (N_12603,N_8084,N_7588);
nor U12604 (N_12604,N_7927,N_6807);
or U12605 (N_12605,N_6266,N_7996);
nand U12606 (N_12606,N_6934,N_9811);
nor U12607 (N_12607,N_9850,N_7903);
or U12608 (N_12608,N_9111,N_6800);
and U12609 (N_12609,N_6779,N_5592);
or U12610 (N_12610,N_9519,N_9595);
or U12611 (N_12611,N_6186,N_9572);
or U12612 (N_12612,N_8919,N_9664);
and U12613 (N_12613,N_6750,N_8013);
xnor U12614 (N_12614,N_6451,N_5800);
nand U12615 (N_12615,N_9407,N_6130);
or U12616 (N_12616,N_7201,N_8604);
and U12617 (N_12617,N_6002,N_8281);
nor U12618 (N_12618,N_9583,N_7536);
nand U12619 (N_12619,N_7902,N_5967);
xor U12620 (N_12620,N_7487,N_7161);
and U12621 (N_12621,N_6539,N_8243);
nor U12622 (N_12622,N_9527,N_8151);
nor U12623 (N_12623,N_6681,N_5825);
nor U12624 (N_12624,N_8234,N_7565);
nand U12625 (N_12625,N_7256,N_9708);
or U12626 (N_12626,N_5768,N_8768);
and U12627 (N_12627,N_7118,N_7669);
or U12628 (N_12628,N_5076,N_9930);
and U12629 (N_12629,N_5031,N_6891);
nor U12630 (N_12630,N_8365,N_9105);
nand U12631 (N_12631,N_7882,N_8744);
nor U12632 (N_12632,N_9840,N_8905);
xnor U12633 (N_12633,N_6485,N_9239);
or U12634 (N_12634,N_7040,N_9045);
xnor U12635 (N_12635,N_9124,N_7130);
or U12636 (N_12636,N_8699,N_9954);
nand U12637 (N_12637,N_9549,N_7719);
or U12638 (N_12638,N_5985,N_5096);
and U12639 (N_12639,N_8262,N_7990);
nor U12640 (N_12640,N_7241,N_8125);
and U12641 (N_12641,N_5554,N_7646);
or U12642 (N_12642,N_6797,N_6325);
or U12643 (N_12643,N_9974,N_9671);
or U12644 (N_12644,N_8599,N_9007);
nor U12645 (N_12645,N_6579,N_7611);
nor U12646 (N_12646,N_6335,N_7063);
or U12647 (N_12647,N_7857,N_8092);
nand U12648 (N_12648,N_6971,N_8717);
or U12649 (N_12649,N_6551,N_7797);
xor U12650 (N_12650,N_7024,N_8832);
or U12651 (N_12651,N_5422,N_7626);
and U12652 (N_12652,N_7384,N_8314);
and U12653 (N_12653,N_8153,N_5593);
nand U12654 (N_12654,N_7228,N_6826);
nand U12655 (N_12655,N_5502,N_6858);
or U12656 (N_12656,N_6044,N_8905);
nand U12657 (N_12657,N_5136,N_8799);
nor U12658 (N_12658,N_5804,N_7278);
xnor U12659 (N_12659,N_8616,N_6910);
or U12660 (N_12660,N_7091,N_7758);
xnor U12661 (N_12661,N_7776,N_8748);
or U12662 (N_12662,N_8519,N_5226);
nand U12663 (N_12663,N_9443,N_7727);
or U12664 (N_12664,N_8889,N_6247);
nand U12665 (N_12665,N_7789,N_8511);
nand U12666 (N_12666,N_5989,N_7224);
nor U12667 (N_12667,N_8214,N_5149);
nor U12668 (N_12668,N_9003,N_8820);
or U12669 (N_12669,N_6261,N_5511);
or U12670 (N_12670,N_9940,N_8672);
nor U12671 (N_12671,N_8563,N_5553);
or U12672 (N_12672,N_5872,N_9802);
nor U12673 (N_12673,N_7967,N_9287);
xnor U12674 (N_12674,N_8020,N_8424);
and U12675 (N_12675,N_5232,N_9962);
or U12676 (N_12676,N_8600,N_6486);
and U12677 (N_12677,N_6091,N_5845);
nand U12678 (N_12678,N_6029,N_7245);
xor U12679 (N_12679,N_6694,N_7031);
xnor U12680 (N_12680,N_5167,N_6334);
nand U12681 (N_12681,N_7410,N_7581);
nand U12682 (N_12682,N_5401,N_9482);
and U12683 (N_12683,N_7139,N_9428);
and U12684 (N_12684,N_6812,N_5495);
and U12685 (N_12685,N_7240,N_9725);
nand U12686 (N_12686,N_5196,N_6914);
xnor U12687 (N_12687,N_8435,N_9127);
and U12688 (N_12688,N_6528,N_5493);
nor U12689 (N_12689,N_8264,N_9278);
nand U12690 (N_12690,N_8495,N_7486);
and U12691 (N_12691,N_5861,N_5014);
xnor U12692 (N_12692,N_5876,N_6063);
or U12693 (N_12693,N_9589,N_9347);
nand U12694 (N_12694,N_9938,N_6266);
or U12695 (N_12695,N_7576,N_8172);
nor U12696 (N_12696,N_7593,N_8255);
or U12697 (N_12697,N_7727,N_5963);
or U12698 (N_12698,N_5077,N_6053);
xor U12699 (N_12699,N_9257,N_6122);
nand U12700 (N_12700,N_5317,N_9468);
xor U12701 (N_12701,N_9925,N_5289);
and U12702 (N_12702,N_9700,N_9988);
or U12703 (N_12703,N_8199,N_6311);
and U12704 (N_12704,N_7348,N_5240);
and U12705 (N_12705,N_9946,N_8908);
and U12706 (N_12706,N_8454,N_9814);
xor U12707 (N_12707,N_5289,N_6381);
or U12708 (N_12708,N_8715,N_7983);
nor U12709 (N_12709,N_5416,N_6617);
xnor U12710 (N_12710,N_9687,N_8036);
or U12711 (N_12711,N_9543,N_5368);
or U12712 (N_12712,N_5574,N_5299);
nand U12713 (N_12713,N_5265,N_9570);
nor U12714 (N_12714,N_6631,N_7371);
and U12715 (N_12715,N_6932,N_9890);
or U12716 (N_12716,N_5540,N_6709);
nand U12717 (N_12717,N_7166,N_9949);
nand U12718 (N_12718,N_5413,N_5822);
nand U12719 (N_12719,N_8417,N_8391);
nor U12720 (N_12720,N_8318,N_9131);
nand U12721 (N_12721,N_7964,N_7781);
nor U12722 (N_12722,N_8471,N_8355);
or U12723 (N_12723,N_7193,N_9921);
or U12724 (N_12724,N_8822,N_8215);
nor U12725 (N_12725,N_8801,N_6460);
nand U12726 (N_12726,N_9455,N_8971);
nand U12727 (N_12727,N_7561,N_8630);
or U12728 (N_12728,N_6846,N_9148);
xnor U12729 (N_12729,N_7171,N_9903);
or U12730 (N_12730,N_8427,N_7729);
nor U12731 (N_12731,N_8043,N_9056);
nand U12732 (N_12732,N_6667,N_8634);
xnor U12733 (N_12733,N_8615,N_7089);
xnor U12734 (N_12734,N_9606,N_6913);
nand U12735 (N_12735,N_7778,N_5461);
or U12736 (N_12736,N_7955,N_6208);
nand U12737 (N_12737,N_9026,N_6764);
nand U12738 (N_12738,N_7928,N_6497);
xnor U12739 (N_12739,N_9825,N_8467);
nor U12740 (N_12740,N_8293,N_7253);
xor U12741 (N_12741,N_5345,N_9611);
nor U12742 (N_12742,N_6430,N_8256);
and U12743 (N_12743,N_7255,N_5452);
and U12744 (N_12744,N_9841,N_5518);
nand U12745 (N_12745,N_9137,N_7587);
or U12746 (N_12746,N_7828,N_5542);
nand U12747 (N_12747,N_6005,N_5329);
or U12748 (N_12748,N_5258,N_6543);
nor U12749 (N_12749,N_5742,N_6979);
nand U12750 (N_12750,N_7008,N_5547);
and U12751 (N_12751,N_5447,N_5693);
nor U12752 (N_12752,N_7204,N_5932);
xnor U12753 (N_12753,N_5132,N_9066);
nand U12754 (N_12754,N_9056,N_9739);
or U12755 (N_12755,N_5189,N_9707);
nand U12756 (N_12756,N_6878,N_9123);
xnor U12757 (N_12757,N_8235,N_9626);
or U12758 (N_12758,N_5816,N_9730);
or U12759 (N_12759,N_7004,N_8133);
or U12760 (N_12760,N_7005,N_8992);
or U12761 (N_12761,N_8759,N_9095);
nor U12762 (N_12762,N_6587,N_5282);
nor U12763 (N_12763,N_5040,N_9072);
and U12764 (N_12764,N_8087,N_8908);
nand U12765 (N_12765,N_7824,N_9802);
nand U12766 (N_12766,N_7900,N_5148);
and U12767 (N_12767,N_5683,N_8536);
nand U12768 (N_12768,N_9604,N_5203);
and U12769 (N_12769,N_9637,N_9707);
nand U12770 (N_12770,N_9089,N_7768);
nand U12771 (N_12771,N_7027,N_8273);
nand U12772 (N_12772,N_6271,N_5665);
and U12773 (N_12773,N_8459,N_5216);
nand U12774 (N_12774,N_7065,N_7041);
and U12775 (N_12775,N_6573,N_9267);
or U12776 (N_12776,N_7346,N_9147);
and U12777 (N_12777,N_8048,N_9426);
xor U12778 (N_12778,N_6266,N_5104);
nor U12779 (N_12779,N_5059,N_8715);
and U12780 (N_12780,N_9458,N_6956);
xnor U12781 (N_12781,N_8199,N_5657);
xor U12782 (N_12782,N_9501,N_8881);
nor U12783 (N_12783,N_7731,N_7596);
xnor U12784 (N_12784,N_9277,N_5542);
nand U12785 (N_12785,N_5054,N_5522);
nor U12786 (N_12786,N_8272,N_6345);
or U12787 (N_12787,N_9675,N_5152);
and U12788 (N_12788,N_6155,N_7704);
nand U12789 (N_12789,N_7151,N_9467);
or U12790 (N_12790,N_5017,N_7529);
and U12791 (N_12791,N_8338,N_7246);
and U12792 (N_12792,N_6726,N_5827);
and U12793 (N_12793,N_6175,N_7767);
nand U12794 (N_12794,N_6488,N_9542);
nor U12795 (N_12795,N_7959,N_8442);
or U12796 (N_12796,N_7441,N_9925);
xnor U12797 (N_12797,N_5087,N_6271);
or U12798 (N_12798,N_6016,N_7964);
nand U12799 (N_12799,N_8273,N_8754);
nand U12800 (N_12800,N_5736,N_7510);
or U12801 (N_12801,N_7054,N_6096);
nor U12802 (N_12802,N_9656,N_5442);
and U12803 (N_12803,N_5324,N_9103);
nand U12804 (N_12804,N_6058,N_9935);
nor U12805 (N_12805,N_9841,N_8258);
nand U12806 (N_12806,N_9876,N_8658);
xor U12807 (N_12807,N_6522,N_7945);
or U12808 (N_12808,N_9728,N_7681);
or U12809 (N_12809,N_5190,N_7820);
and U12810 (N_12810,N_6511,N_6936);
nand U12811 (N_12811,N_6551,N_7679);
nand U12812 (N_12812,N_5055,N_9527);
nand U12813 (N_12813,N_8627,N_9848);
or U12814 (N_12814,N_6436,N_6297);
nand U12815 (N_12815,N_8776,N_6361);
nand U12816 (N_12816,N_5479,N_8555);
nand U12817 (N_12817,N_5003,N_5822);
xnor U12818 (N_12818,N_9141,N_5055);
or U12819 (N_12819,N_6516,N_7498);
or U12820 (N_12820,N_9871,N_6203);
nor U12821 (N_12821,N_5168,N_7195);
nor U12822 (N_12822,N_9353,N_5939);
xnor U12823 (N_12823,N_8916,N_9412);
nor U12824 (N_12824,N_8224,N_8688);
xor U12825 (N_12825,N_8145,N_8194);
nor U12826 (N_12826,N_8894,N_5867);
nor U12827 (N_12827,N_7114,N_7758);
nor U12828 (N_12828,N_8737,N_7126);
nor U12829 (N_12829,N_7843,N_8146);
nor U12830 (N_12830,N_9793,N_5268);
or U12831 (N_12831,N_9388,N_8810);
nor U12832 (N_12832,N_9924,N_7740);
nand U12833 (N_12833,N_8294,N_5288);
xnor U12834 (N_12834,N_6958,N_5450);
and U12835 (N_12835,N_8429,N_9455);
nand U12836 (N_12836,N_6009,N_6222);
nand U12837 (N_12837,N_9304,N_7510);
nand U12838 (N_12838,N_8642,N_6264);
or U12839 (N_12839,N_9656,N_8864);
xor U12840 (N_12840,N_5395,N_5944);
xor U12841 (N_12841,N_7543,N_5783);
nand U12842 (N_12842,N_5065,N_5931);
and U12843 (N_12843,N_8981,N_6262);
nand U12844 (N_12844,N_7197,N_6504);
or U12845 (N_12845,N_8566,N_9268);
and U12846 (N_12846,N_6546,N_9904);
and U12847 (N_12847,N_5267,N_7581);
nand U12848 (N_12848,N_5871,N_9502);
nor U12849 (N_12849,N_9547,N_5360);
xnor U12850 (N_12850,N_8480,N_9281);
or U12851 (N_12851,N_6269,N_6969);
or U12852 (N_12852,N_9640,N_5263);
xnor U12853 (N_12853,N_8539,N_8275);
or U12854 (N_12854,N_6357,N_8399);
xnor U12855 (N_12855,N_8854,N_8188);
and U12856 (N_12856,N_5127,N_9118);
nand U12857 (N_12857,N_8134,N_5304);
xor U12858 (N_12858,N_5724,N_6697);
or U12859 (N_12859,N_7843,N_6060);
and U12860 (N_12860,N_9617,N_6612);
xor U12861 (N_12861,N_9210,N_6400);
nand U12862 (N_12862,N_7132,N_9750);
xnor U12863 (N_12863,N_7765,N_6951);
and U12864 (N_12864,N_7106,N_9609);
nand U12865 (N_12865,N_6411,N_7118);
nor U12866 (N_12866,N_6201,N_5110);
or U12867 (N_12867,N_5090,N_5155);
xor U12868 (N_12868,N_5874,N_6159);
nor U12869 (N_12869,N_6079,N_7133);
xnor U12870 (N_12870,N_6781,N_5756);
or U12871 (N_12871,N_9921,N_8456);
nor U12872 (N_12872,N_5569,N_7073);
xor U12873 (N_12873,N_5049,N_5849);
nand U12874 (N_12874,N_5918,N_7260);
and U12875 (N_12875,N_7199,N_5720);
nor U12876 (N_12876,N_6475,N_5985);
and U12877 (N_12877,N_7974,N_9023);
nor U12878 (N_12878,N_8248,N_9210);
and U12879 (N_12879,N_6013,N_7171);
nand U12880 (N_12880,N_7188,N_8198);
nand U12881 (N_12881,N_5868,N_5594);
nand U12882 (N_12882,N_8128,N_9948);
or U12883 (N_12883,N_8765,N_7596);
nor U12884 (N_12884,N_6569,N_6002);
and U12885 (N_12885,N_6716,N_9317);
nor U12886 (N_12886,N_5148,N_6766);
nand U12887 (N_12887,N_6064,N_7317);
or U12888 (N_12888,N_5292,N_9359);
nand U12889 (N_12889,N_5915,N_6634);
nor U12890 (N_12890,N_7038,N_9787);
or U12891 (N_12891,N_5061,N_8158);
and U12892 (N_12892,N_9494,N_8101);
nor U12893 (N_12893,N_5350,N_5211);
and U12894 (N_12894,N_8141,N_5965);
and U12895 (N_12895,N_9422,N_6158);
or U12896 (N_12896,N_7323,N_8530);
xor U12897 (N_12897,N_6394,N_9270);
or U12898 (N_12898,N_8247,N_7978);
nand U12899 (N_12899,N_8794,N_7087);
nor U12900 (N_12900,N_9501,N_8967);
nand U12901 (N_12901,N_7447,N_6081);
and U12902 (N_12902,N_7821,N_5925);
nand U12903 (N_12903,N_9882,N_5934);
and U12904 (N_12904,N_9026,N_5926);
nand U12905 (N_12905,N_6683,N_7716);
or U12906 (N_12906,N_5495,N_5978);
xnor U12907 (N_12907,N_6381,N_9092);
xnor U12908 (N_12908,N_5978,N_8665);
xor U12909 (N_12909,N_8425,N_8807);
nor U12910 (N_12910,N_5709,N_9240);
or U12911 (N_12911,N_6299,N_9657);
and U12912 (N_12912,N_5158,N_8900);
nand U12913 (N_12913,N_5545,N_7149);
or U12914 (N_12914,N_5919,N_8650);
or U12915 (N_12915,N_5402,N_8509);
or U12916 (N_12916,N_9141,N_7804);
or U12917 (N_12917,N_8748,N_6600);
xnor U12918 (N_12918,N_5855,N_7930);
xnor U12919 (N_12919,N_7439,N_6021);
or U12920 (N_12920,N_9392,N_5405);
or U12921 (N_12921,N_8730,N_8433);
xnor U12922 (N_12922,N_7731,N_8330);
xnor U12923 (N_12923,N_9890,N_8673);
xor U12924 (N_12924,N_9126,N_6581);
nand U12925 (N_12925,N_7326,N_6159);
nor U12926 (N_12926,N_7103,N_9655);
nor U12927 (N_12927,N_5906,N_7582);
and U12928 (N_12928,N_6869,N_8698);
or U12929 (N_12929,N_7497,N_6247);
nand U12930 (N_12930,N_7199,N_7917);
nor U12931 (N_12931,N_9353,N_8009);
xor U12932 (N_12932,N_9519,N_6074);
nand U12933 (N_12933,N_8445,N_9385);
nor U12934 (N_12934,N_8728,N_5386);
or U12935 (N_12935,N_9197,N_9395);
nor U12936 (N_12936,N_9535,N_6001);
nor U12937 (N_12937,N_6677,N_9805);
or U12938 (N_12938,N_6319,N_8367);
xnor U12939 (N_12939,N_9933,N_9659);
or U12940 (N_12940,N_5744,N_6594);
nor U12941 (N_12941,N_5587,N_6672);
nor U12942 (N_12942,N_9405,N_6043);
or U12943 (N_12943,N_6361,N_6176);
nor U12944 (N_12944,N_6970,N_5533);
and U12945 (N_12945,N_6669,N_7462);
nor U12946 (N_12946,N_5663,N_7016);
xnor U12947 (N_12947,N_5797,N_8706);
nand U12948 (N_12948,N_6585,N_9492);
nand U12949 (N_12949,N_6143,N_9579);
nor U12950 (N_12950,N_8017,N_6056);
nand U12951 (N_12951,N_5462,N_7060);
xor U12952 (N_12952,N_6243,N_7298);
nand U12953 (N_12953,N_8449,N_8390);
nand U12954 (N_12954,N_9039,N_5463);
xnor U12955 (N_12955,N_8344,N_7243);
xor U12956 (N_12956,N_7521,N_9670);
nor U12957 (N_12957,N_6300,N_7654);
nand U12958 (N_12958,N_8204,N_6486);
nor U12959 (N_12959,N_7259,N_8849);
nand U12960 (N_12960,N_5294,N_6237);
and U12961 (N_12961,N_5996,N_7160);
and U12962 (N_12962,N_9994,N_9472);
xor U12963 (N_12963,N_7726,N_7709);
xor U12964 (N_12964,N_9870,N_6880);
xnor U12965 (N_12965,N_9155,N_8067);
nor U12966 (N_12966,N_8810,N_8756);
nand U12967 (N_12967,N_5818,N_8747);
xor U12968 (N_12968,N_5528,N_7950);
nand U12969 (N_12969,N_7836,N_5927);
and U12970 (N_12970,N_5885,N_5238);
nor U12971 (N_12971,N_9166,N_9334);
xor U12972 (N_12972,N_6540,N_6912);
and U12973 (N_12973,N_7096,N_7952);
or U12974 (N_12974,N_8364,N_6909);
xor U12975 (N_12975,N_9839,N_6364);
nor U12976 (N_12976,N_8910,N_5380);
nor U12977 (N_12977,N_6376,N_9196);
nor U12978 (N_12978,N_7462,N_7419);
nand U12979 (N_12979,N_6432,N_8253);
xor U12980 (N_12980,N_7840,N_5513);
xor U12981 (N_12981,N_7054,N_8262);
or U12982 (N_12982,N_8838,N_6190);
or U12983 (N_12983,N_8301,N_8932);
or U12984 (N_12984,N_5837,N_6519);
nand U12985 (N_12985,N_5871,N_5825);
nor U12986 (N_12986,N_8576,N_8151);
nor U12987 (N_12987,N_7486,N_7830);
nor U12988 (N_12988,N_9911,N_8805);
xor U12989 (N_12989,N_9689,N_9966);
nand U12990 (N_12990,N_5769,N_7943);
nand U12991 (N_12991,N_6003,N_6034);
and U12992 (N_12992,N_9310,N_7377);
xor U12993 (N_12993,N_8403,N_9687);
nand U12994 (N_12994,N_7848,N_9158);
or U12995 (N_12995,N_7211,N_9114);
and U12996 (N_12996,N_9830,N_8874);
xor U12997 (N_12997,N_8845,N_7214);
or U12998 (N_12998,N_9219,N_5141);
nand U12999 (N_12999,N_6551,N_5758);
xor U13000 (N_13000,N_6621,N_9590);
xnor U13001 (N_13001,N_8842,N_6884);
and U13002 (N_13002,N_9975,N_8475);
xor U13003 (N_13003,N_6174,N_8066);
nor U13004 (N_13004,N_7886,N_6107);
nor U13005 (N_13005,N_9004,N_6348);
xor U13006 (N_13006,N_9872,N_5388);
and U13007 (N_13007,N_9332,N_8224);
xnor U13008 (N_13008,N_7243,N_9296);
and U13009 (N_13009,N_8237,N_8332);
nand U13010 (N_13010,N_8672,N_9059);
nor U13011 (N_13011,N_5078,N_9733);
or U13012 (N_13012,N_6573,N_9947);
xnor U13013 (N_13013,N_7578,N_6149);
or U13014 (N_13014,N_8567,N_8171);
xor U13015 (N_13015,N_8110,N_8613);
nor U13016 (N_13016,N_9966,N_7867);
and U13017 (N_13017,N_5615,N_6177);
nand U13018 (N_13018,N_9565,N_6374);
and U13019 (N_13019,N_9514,N_5007);
nand U13020 (N_13020,N_9927,N_8753);
and U13021 (N_13021,N_6774,N_9933);
nand U13022 (N_13022,N_6906,N_9110);
and U13023 (N_13023,N_8951,N_8529);
nand U13024 (N_13024,N_7420,N_9279);
and U13025 (N_13025,N_8643,N_5095);
nand U13026 (N_13026,N_7482,N_7334);
xor U13027 (N_13027,N_9249,N_9251);
xor U13028 (N_13028,N_9719,N_8555);
and U13029 (N_13029,N_7684,N_6027);
xnor U13030 (N_13030,N_8601,N_8688);
or U13031 (N_13031,N_5855,N_7539);
and U13032 (N_13032,N_5843,N_9941);
nand U13033 (N_13033,N_7233,N_8512);
nand U13034 (N_13034,N_8580,N_7377);
nor U13035 (N_13035,N_5040,N_6389);
nor U13036 (N_13036,N_7926,N_8267);
nand U13037 (N_13037,N_6653,N_6736);
nor U13038 (N_13038,N_5768,N_6613);
or U13039 (N_13039,N_8759,N_8770);
or U13040 (N_13040,N_7822,N_7079);
nand U13041 (N_13041,N_8195,N_5808);
xor U13042 (N_13042,N_6348,N_9880);
nor U13043 (N_13043,N_9585,N_5616);
nand U13044 (N_13044,N_5220,N_8516);
nand U13045 (N_13045,N_6116,N_6099);
xnor U13046 (N_13046,N_6733,N_7307);
xnor U13047 (N_13047,N_5938,N_8224);
nand U13048 (N_13048,N_8931,N_6217);
nor U13049 (N_13049,N_5718,N_5785);
nor U13050 (N_13050,N_7145,N_9450);
nand U13051 (N_13051,N_9973,N_8824);
nor U13052 (N_13052,N_8705,N_9640);
or U13053 (N_13053,N_6165,N_7794);
nand U13054 (N_13054,N_8662,N_7681);
xor U13055 (N_13055,N_8099,N_6125);
nor U13056 (N_13056,N_5020,N_5970);
nand U13057 (N_13057,N_5371,N_7365);
nor U13058 (N_13058,N_6091,N_6760);
nor U13059 (N_13059,N_9180,N_6969);
xnor U13060 (N_13060,N_6770,N_9641);
nor U13061 (N_13061,N_5364,N_7705);
xnor U13062 (N_13062,N_9410,N_8483);
nand U13063 (N_13063,N_9776,N_6733);
and U13064 (N_13064,N_5354,N_8885);
xor U13065 (N_13065,N_8776,N_9421);
or U13066 (N_13066,N_7874,N_9728);
xnor U13067 (N_13067,N_7608,N_9256);
xor U13068 (N_13068,N_9177,N_9127);
nand U13069 (N_13069,N_6442,N_6121);
xnor U13070 (N_13070,N_9691,N_8862);
nor U13071 (N_13071,N_7646,N_7738);
or U13072 (N_13072,N_7143,N_8295);
nor U13073 (N_13073,N_8711,N_7096);
or U13074 (N_13074,N_5968,N_5413);
nor U13075 (N_13075,N_5548,N_7765);
nor U13076 (N_13076,N_6179,N_5256);
nor U13077 (N_13077,N_8377,N_6391);
nor U13078 (N_13078,N_8581,N_9510);
and U13079 (N_13079,N_7789,N_9948);
xnor U13080 (N_13080,N_8454,N_9825);
xnor U13081 (N_13081,N_6356,N_8042);
and U13082 (N_13082,N_8503,N_8991);
nor U13083 (N_13083,N_6040,N_7331);
nor U13084 (N_13084,N_6165,N_8716);
and U13085 (N_13085,N_5830,N_5657);
and U13086 (N_13086,N_6037,N_5555);
and U13087 (N_13087,N_8812,N_8390);
or U13088 (N_13088,N_5175,N_8026);
xor U13089 (N_13089,N_9483,N_9877);
nand U13090 (N_13090,N_9418,N_7475);
nor U13091 (N_13091,N_5890,N_5158);
nand U13092 (N_13092,N_6862,N_8265);
xor U13093 (N_13093,N_5308,N_8458);
and U13094 (N_13094,N_8916,N_5866);
nand U13095 (N_13095,N_6959,N_8727);
nor U13096 (N_13096,N_9080,N_5307);
xnor U13097 (N_13097,N_9209,N_6837);
nand U13098 (N_13098,N_7327,N_9626);
xnor U13099 (N_13099,N_7697,N_6979);
and U13100 (N_13100,N_6140,N_5230);
nor U13101 (N_13101,N_7764,N_7508);
xnor U13102 (N_13102,N_7146,N_9683);
nand U13103 (N_13103,N_7794,N_9916);
and U13104 (N_13104,N_5228,N_5320);
and U13105 (N_13105,N_6744,N_7056);
or U13106 (N_13106,N_7130,N_7920);
nor U13107 (N_13107,N_8652,N_8373);
xnor U13108 (N_13108,N_7597,N_8365);
xnor U13109 (N_13109,N_6970,N_8683);
nand U13110 (N_13110,N_5969,N_7737);
xor U13111 (N_13111,N_7232,N_5063);
nand U13112 (N_13112,N_6892,N_9722);
nor U13113 (N_13113,N_6473,N_6696);
and U13114 (N_13114,N_6618,N_5394);
or U13115 (N_13115,N_9108,N_6160);
nand U13116 (N_13116,N_8022,N_5640);
and U13117 (N_13117,N_5635,N_7514);
xnor U13118 (N_13118,N_9992,N_5429);
nor U13119 (N_13119,N_8914,N_6599);
and U13120 (N_13120,N_5629,N_5406);
or U13121 (N_13121,N_9988,N_7865);
nor U13122 (N_13122,N_5579,N_6780);
nand U13123 (N_13123,N_5148,N_9617);
nand U13124 (N_13124,N_9973,N_6094);
or U13125 (N_13125,N_6299,N_8979);
and U13126 (N_13126,N_6110,N_9129);
and U13127 (N_13127,N_5634,N_6122);
and U13128 (N_13128,N_8935,N_8618);
nand U13129 (N_13129,N_5246,N_8448);
nand U13130 (N_13130,N_5273,N_7491);
or U13131 (N_13131,N_6202,N_5903);
nand U13132 (N_13132,N_9327,N_9250);
nor U13133 (N_13133,N_6827,N_6436);
nor U13134 (N_13134,N_7549,N_6830);
nor U13135 (N_13135,N_7552,N_8947);
or U13136 (N_13136,N_7585,N_9127);
and U13137 (N_13137,N_5078,N_9086);
or U13138 (N_13138,N_6523,N_5467);
and U13139 (N_13139,N_6430,N_5024);
or U13140 (N_13140,N_9871,N_8076);
or U13141 (N_13141,N_9778,N_5617);
nor U13142 (N_13142,N_7238,N_6657);
nand U13143 (N_13143,N_6918,N_9657);
and U13144 (N_13144,N_5951,N_6876);
or U13145 (N_13145,N_5806,N_5761);
nor U13146 (N_13146,N_8795,N_8988);
or U13147 (N_13147,N_8947,N_6315);
xor U13148 (N_13148,N_9034,N_8721);
nand U13149 (N_13149,N_6129,N_5450);
nand U13150 (N_13150,N_9471,N_5040);
xor U13151 (N_13151,N_6470,N_9762);
nor U13152 (N_13152,N_6992,N_5933);
and U13153 (N_13153,N_9091,N_5552);
and U13154 (N_13154,N_6386,N_9443);
xor U13155 (N_13155,N_9788,N_7800);
nand U13156 (N_13156,N_6406,N_6861);
and U13157 (N_13157,N_7540,N_8728);
or U13158 (N_13158,N_7149,N_8022);
xor U13159 (N_13159,N_8824,N_6661);
xnor U13160 (N_13160,N_5904,N_9091);
nor U13161 (N_13161,N_9762,N_6187);
nand U13162 (N_13162,N_8097,N_5851);
or U13163 (N_13163,N_5623,N_7315);
and U13164 (N_13164,N_6826,N_6396);
nor U13165 (N_13165,N_5035,N_6343);
or U13166 (N_13166,N_6007,N_5247);
nand U13167 (N_13167,N_6700,N_9508);
nor U13168 (N_13168,N_8156,N_7248);
nand U13169 (N_13169,N_6478,N_7705);
xor U13170 (N_13170,N_5242,N_7702);
and U13171 (N_13171,N_8527,N_8784);
xor U13172 (N_13172,N_9714,N_7062);
xor U13173 (N_13173,N_6989,N_5185);
and U13174 (N_13174,N_9557,N_8402);
or U13175 (N_13175,N_6582,N_5349);
nand U13176 (N_13176,N_5821,N_9399);
or U13177 (N_13177,N_6783,N_7758);
nand U13178 (N_13178,N_5412,N_9736);
or U13179 (N_13179,N_5633,N_5318);
or U13180 (N_13180,N_6579,N_5013);
or U13181 (N_13181,N_8183,N_8634);
or U13182 (N_13182,N_7295,N_5455);
xor U13183 (N_13183,N_5286,N_5297);
xor U13184 (N_13184,N_6093,N_9668);
xor U13185 (N_13185,N_5227,N_9823);
xnor U13186 (N_13186,N_6821,N_9857);
and U13187 (N_13187,N_5707,N_5449);
and U13188 (N_13188,N_5169,N_5745);
and U13189 (N_13189,N_5330,N_5432);
nor U13190 (N_13190,N_6089,N_6661);
nor U13191 (N_13191,N_7756,N_6468);
xnor U13192 (N_13192,N_8288,N_6437);
nor U13193 (N_13193,N_5733,N_6954);
xor U13194 (N_13194,N_7481,N_5983);
xor U13195 (N_13195,N_6216,N_9509);
and U13196 (N_13196,N_7574,N_7224);
and U13197 (N_13197,N_5565,N_9951);
xnor U13198 (N_13198,N_6233,N_8292);
and U13199 (N_13199,N_9189,N_7935);
nand U13200 (N_13200,N_8482,N_9479);
and U13201 (N_13201,N_8261,N_8783);
nand U13202 (N_13202,N_8992,N_6422);
nor U13203 (N_13203,N_5938,N_6299);
nor U13204 (N_13204,N_8548,N_9625);
or U13205 (N_13205,N_8101,N_9491);
or U13206 (N_13206,N_8836,N_5375);
nor U13207 (N_13207,N_6975,N_9330);
or U13208 (N_13208,N_5116,N_9259);
or U13209 (N_13209,N_8912,N_9871);
nor U13210 (N_13210,N_6560,N_5309);
nand U13211 (N_13211,N_5717,N_6531);
nand U13212 (N_13212,N_6075,N_6821);
nand U13213 (N_13213,N_8150,N_6758);
nand U13214 (N_13214,N_5721,N_9242);
nand U13215 (N_13215,N_9292,N_5316);
and U13216 (N_13216,N_9742,N_6486);
and U13217 (N_13217,N_6053,N_9134);
nand U13218 (N_13218,N_5188,N_8823);
and U13219 (N_13219,N_9740,N_7138);
xnor U13220 (N_13220,N_7800,N_9117);
and U13221 (N_13221,N_9776,N_6622);
nor U13222 (N_13222,N_9404,N_6761);
or U13223 (N_13223,N_7897,N_6246);
nor U13224 (N_13224,N_9071,N_5842);
nor U13225 (N_13225,N_7550,N_7928);
or U13226 (N_13226,N_5355,N_9296);
nor U13227 (N_13227,N_7509,N_8081);
xor U13228 (N_13228,N_9607,N_9153);
xor U13229 (N_13229,N_6051,N_8658);
or U13230 (N_13230,N_7908,N_9379);
nand U13231 (N_13231,N_8963,N_7844);
and U13232 (N_13232,N_8522,N_9904);
nor U13233 (N_13233,N_8366,N_5591);
or U13234 (N_13234,N_6987,N_6023);
and U13235 (N_13235,N_5457,N_9564);
nor U13236 (N_13236,N_5284,N_5863);
and U13237 (N_13237,N_9928,N_7409);
nand U13238 (N_13238,N_6837,N_6273);
nand U13239 (N_13239,N_7913,N_5473);
or U13240 (N_13240,N_6043,N_7461);
xnor U13241 (N_13241,N_5990,N_8856);
nor U13242 (N_13242,N_6012,N_6950);
xnor U13243 (N_13243,N_8805,N_6803);
nand U13244 (N_13244,N_8429,N_8761);
nand U13245 (N_13245,N_6257,N_6509);
and U13246 (N_13246,N_8636,N_6608);
nor U13247 (N_13247,N_6688,N_7456);
xnor U13248 (N_13248,N_5622,N_5462);
nand U13249 (N_13249,N_9351,N_6774);
and U13250 (N_13250,N_6187,N_8906);
or U13251 (N_13251,N_6449,N_6422);
and U13252 (N_13252,N_9424,N_7682);
xnor U13253 (N_13253,N_8534,N_6314);
nand U13254 (N_13254,N_6394,N_6602);
xnor U13255 (N_13255,N_5914,N_7673);
nor U13256 (N_13256,N_8510,N_5808);
xor U13257 (N_13257,N_6918,N_7406);
or U13258 (N_13258,N_5407,N_8065);
nor U13259 (N_13259,N_7690,N_6452);
and U13260 (N_13260,N_9427,N_6569);
nor U13261 (N_13261,N_6565,N_6501);
and U13262 (N_13262,N_5076,N_7500);
and U13263 (N_13263,N_5770,N_9030);
and U13264 (N_13264,N_8833,N_6699);
nor U13265 (N_13265,N_9970,N_5624);
nand U13266 (N_13266,N_6334,N_7227);
xnor U13267 (N_13267,N_9249,N_8706);
and U13268 (N_13268,N_6271,N_9105);
xor U13269 (N_13269,N_6248,N_7116);
or U13270 (N_13270,N_8129,N_8833);
xor U13271 (N_13271,N_5176,N_7550);
and U13272 (N_13272,N_7487,N_5826);
nand U13273 (N_13273,N_7672,N_6447);
xor U13274 (N_13274,N_6561,N_8635);
or U13275 (N_13275,N_5892,N_9238);
xor U13276 (N_13276,N_6361,N_8198);
or U13277 (N_13277,N_8587,N_6396);
nor U13278 (N_13278,N_6284,N_8837);
or U13279 (N_13279,N_5496,N_8614);
xnor U13280 (N_13280,N_6075,N_9983);
nand U13281 (N_13281,N_5915,N_6164);
xnor U13282 (N_13282,N_9241,N_6638);
nor U13283 (N_13283,N_6918,N_5220);
or U13284 (N_13284,N_5343,N_8703);
nor U13285 (N_13285,N_6056,N_5288);
and U13286 (N_13286,N_9205,N_8481);
nand U13287 (N_13287,N_9325,N_8484);
and U13288 (N_13288,N_6889,N_6156);
nor U13289 (N_13289,N_6667,N_6482);
nand U13290 (N_13290,N_5256,N_5972);
nor U13291 (N_13291,N_8924,N_5848);
nor U13292 (N_13292,N_7771,N_7807);
nand U13293 (N_13293,N_6239,N_7910);
or U13294 (N_13294,N_7346,N_8918);
or U13295 (N_13295,N_9383,N_8878);
nor U13296 (N_13296,N_5758,N_5438);
nor U13297 (N_13297,N_6162,N_8632);
nand U13298 (N_13298,N_5317,N_5032);
xor U13299 (N_13299,N_5031,N_6089);
or U13300 (N_13300,N_5721,N_8472);
or U13301 (N_13301,N_7125,N_6205);
and U13302 (N_13302,N_5301,N_7272);
xor U13303 (N_13303,N_5130,N_5565);
nand U13304 (N_13304,N_9053,N_8684);
xor U13305 (N_13305,N_5723,N_6479);
xnor U13306 (N_13306,N_5194,N_8963);
xor U13307 (N_13307,N_8132,N_9519);
nand U13308 (N_13308,N_6982,N_5082);
or U13309 (N_13309,N_5016,N_7643);
or U13310 (N_13310,N_7919,N_9419);
and U13311 (N_13311,N_9468,N_6240);
xor U13312 (N_13312,N_8068,N_8751);
nand U13313 (N_13313,N_7118,N_9791);
and U13314 (N_13314,N_8145,N_6160);
nor U13315 (N_13315,N_6749,N_9471);
nand U13316 (N_13316,N_5138,N_9140);
nand U13317 (N_13317,N_9202,N_5955);
and U13318 (N_13318,N_7286,N_9680);
xor U13319 (N_13319,N_6710,N_9949);
or U13320 (N_13320,N_5050,N_8356);
or U13321 (N_13321,N_9482,N_6001);
nand U13322 (N_13322,N_7188,N_5795);
nand U13323 (N_13323,N_7301,N_9472);
nand U13324 (N_13324,N_5099,N_9205);
nor U13325 (N_13325,N_8387,N_6757);
or U13326 (N_13326,N_5533,N_8750);
xor U13327 (N_13327,N_6180,N_6654);
xnor U13328 (N_13328,N_8770,N_8594);
or U13329 (N_13329,N_5349,N_8739);
and U13330 (N_13330,N_8026,N_6957);
and U13331 (N_13331,N_8833,N_5327);
and U13332 (N_13332,N_5791,N_8657);
nand U13333 (N_13333,N_9957,N_7140);
nor U13334 (N_13334,N_8070,N_7364);
xnor U13335 (N_13335,N_5045,N_9250);
and U13336 (N_13336,N_6389,N_7329);
and U13337 (N_13337,N_9702,N_7537);
or U13338 (N_13338,N_8200,N_7483);
nand U13339 (N_13339,N_8660,N_8819);
nand U13340 (N_13340,N_8497,N_7007);
and U13341 (N_13341,N_9104,N_5652);
xor U13342 (N_13342,N_5964,N_5821);
nand U13343 (N_13343,N_7724,N_6445);
and U13344 (N_13344,N_6500,N_7451);
or U13345 (N_13345,N_6978,N_8011);
xnor U13346 (N_13346,N_7913,N_6132);
nor U13347 (N_13347,N_8161,N_5337);
nor U13348 (N_13348,N_5656,N_9524);
or U13349 (N_13349,N_8091,N_5560);
and U13350 (N_13350,N_6890,N_8471);
xnor U13351 (N_13351,N_5561,N_8101);
or U13352 (N_13352,N_6188,N_8389);
and U13353 (N_13353,N_9227,N_6024);
or U13354 (N_13354,N_8664,N_8782);
or U13355 (N_13355,N_7771,N_8626);
or U13356 (N_13356,N_8589,N_6454);
xor U13357 (N_13357,N_6146,N_6168);
xnor U13358 (N_13358,N_9832,N_5950);
xor U13359 (N_13359,N_7492,N_7959);
and U13360 (N_13360,N_7625,N_7594);
or U13361 (N_13361,N_8167,N_8981);
nand U13362 (N_13362,N_7739,N_7994);
nand U13363 (N_13363,N_8481,N_9337);
and U13364 (N_13364,N_9916,N_6788);
or U13365 (N_13365,N_9433,N_7231);
or U13366 (N_13366,N_8443,N_7417);
nand U13367 (N_13367,N_7761,N_9259);
and U13368 (N_13368,N_9706,N_7411);
or U13369 (N_13369,N_5722,N_9151);
nand U13370 (N_13370,N_7508,N_5786);
or U13371 (N_13371,N_8250,N_5904);
and U13372 (N_13372,N_7812,N_5372);
and U13373 (N_13373,N_8639,N_7769);
nand U13374 (N_13374,N_7187,N_5750);
nor U13375 (N_13375,N_7859,N_9152);
and U13376 (N_13376,N_6556,N_8755);
xor U13377 (N_13377,N_8568,N_5248);
xor U13378 (N_13378,N_5628,N_5534);
and U13379 (N_13379,N_5917,N_9756);
or U13380 (N_13380,N_8801,N_9729);
or U13381 (N_13381,N_6920,N_5789);
xnor U13382 (N_13382,N_8398,N_7371);
nand U13383 (N_13383,N_6133,N_8579);
xnor U13384 (N_13384,N_6193,N_7991);
or U13385 (N_13385,N_7747,N_9912);
xnor U13386 (N_13386,N_8746,N_5683);
and U13387 (N_13387,N_8606,N_5522);
nand U13388 (N_13388,N_6263,N_6229);
nand U13389 (N_13389,N_7442,N_5471);
or U13390 (N_13390,N_8407,N_5103);
xnor U13391 (N_13391,N_5822,N_9210);
nand U13392 (N_13392,N_9794,N_7617);
nor U13393 (N_13393,N_6797,N_7536);
and U13394 (N_13394,N_6867,N_7407);
and U13395 (N_13395,N_5623,N_7467);
nand U13396 (N_13396,N_5480,N_8498);
nor U13397 (N_13397,N_7322,N_8938);
or U13398 (N_13398,N_7057,N_7700);
or U13399 (N_13399,N_6188,N_9927);
nand U13400 (N_13400,N_6841,N_7645);
or U13401 (N_13401,N_6197,N_6083);
or U13402 (N_13402,N_5358,N_9875);
or U13403 (N_13403,N_5968,N_6869);
nor U13404 (N_13404,N_6877,N_8283);
or U13405 (N_13405,N_5819,N_5760);
or U13406 (N_13406,N_7551,N_5026);
xor U13407 (N_13407,N_7384,N_8757);
or U13408 (N_13408,N_8803,N_5061);
and U13409 (N_13409,N_7810,N_5720);
and U13410 (N_13410,N_9998,N_5533);
nand U13411 (N_13411,N_5388,N_6806);
xor U13412 (N_13412,N_5189,N_8926);
and U13413 (N_13413,N_9833,N_8107);
and U13414 (N_13414,N_9893,N_5987);
xnor U13415 (N_13415,N_7361,N_9661);
and U13416 (N_13416,N_7238,N_8334);
nor U13417 (N_13417,N_5095,N_5169);
nor U13418 (N_13418,N_8641,N_9941);
and U13419 (N_13419,N_9923,N_9834);
nand U13420 (N_13420,N_8082,N_9475);
and U13421 (N_13421,N_5390,N_5639);
nor U13422 (N_13422,N_5019,N_5084);
or U13423 (N_13423,N_7511,N_7138);
and U13424 (N_13424,N_5188,N_7030);
nor U13425 (N_13425,N_9301,N_6328);
and U13426 (N_13426,N_9955,N_7995);
and U13427 (N_13427,N_7273,N_7868);
or U13428 (N_13428,N_7671,N_9360);
nand U13429 (N_13429,N_7795,N_9977);
nand U13430 (N_13430,N_5676,N_5666);
nand U13431 (N_13431,N_9031,N_7025);
xnor U13432 (N_13432,N_6266,N_9484);
nand U13433 (N_13433,N_8992,N_8317);
xnor U13434 (N_13434,N_9292,N_8798);
and U13435 (N_13435,N_6548,N_6378);
nand U13436 (N_13436,N_7023,N_9955);
and U13437 (N_13437,N_9786,N_6297);
and U13438 (N_13438,N_5958,N_5167);
nor U13439 (N_13439,N_5377,N_7790);
and U13440 (N_13440,N_6546,N_5539);
and U13441 (N_13441,N_5177,N_9678);
nand U13442 (N_13442,N_5419,N_7966);
or U13443 (N_13443,N_6546,N_8484);
xnor U13444 (N_13444,N_9707,N_8241);
and U13445 (N_13445,N_6944,N_8286);
nor U13446 (N_13446,N_9928,N_6650);
or U13447 (N_13447,N_9356,N_7723);
or U13448 (N_13448,N_7649,N_8786);
or U13449 (N_13449,N_7297,N_5475);
nand U13450 (N_13450,N_6427,N_7282);
and U13451 (N_13451,N_5943,N_9099);
or U13452 (N_13452,N_8370,N_9529);
nor U13453 (N_13453,N_5411,N_5670);
nor U13454 (N_13454,N_9219,N_6796);
nor U13455 (N_13455,N_9829,N_6216);
nor U13456 (N_13456,N_8445,N_9153);
or U13457 (N_13457,N_8123,N_7598);
nand U13458 (N_13458,N_8191,N_9487);
nor U13459 (N_13459,N_5114,N_7310);
xnor U13460 (N_13460,N_6410,N_9589);
and U13461 (N_13461,N_5108,N_9675);
or U13462 (N_13462,N_8766,N_8611);
and U13463 (N_13463,N_9048,N_6422);
and U13464 (N_13464,N_7199,N_7176);
xnor U13465 (N_13465,N_6994,N_7161);
or U13466 (N_13466,N_8045,N_7325);
and U13467 (N_13467,N_9909,N_5075);
or U13468 (N_13468,N_9749,N_5781);
or U13469 (N_13469,N_7792,N_5343);
nand U13470 (N_13470,N_5337,N_5436);
or U13471 (N_13471,N_5707,N_8451);
nor U13472 (N_13472,N_8529,N_9635);
xor U13473 (N_13473,N_6030,N_8007);
nor U13474 (N_13474,N_8182,N_9888);
or U13475 (N_13475,N_6556,N_9140);
xor U13476 (N_13476,N_8130,N_9089);
nor U13477 (N_13477,N_9520,N_6701);
or U13478 (N_13478,N_5989,N_5905);
xor U13479 (N_13479,N_9404,N_6802);
nand U13480 (N_13480,N_7295,N_5544);
nand U13481 (N_13481,N_6296,N_7457);
and U13482 (N_13482,N_9119,N_5359);
nand U13483 (N_13483,N_7962,N_6562);
and U13484 (N_13484,N_8883,N_5013);
and U13485 (N_13485,N_5443,N_8894);
xnor U13486 (N_13486,N_6595,N_6647);
xor U13487 (N_13487,N_6149,N_7153);
nand U13488 (N_13488,N_9475,N_5007);
or U13489 (N_13489,N_7775,N_8389);
xnor U13490 (N_13490,N_9814,N_5806);
and U13491 (N_13491,N_8302,N_6535);
xor U13492 (N_13492,N_7137,N_6713);
and U13493 (N_13493,N_5390,N_9431);
and U13494 (N_13494,N_7967,N_7763);
nand U13495 (N_13495,N_7300,N_7503);
or U13496 (N_13496,N_5762,N_8306);
xor U13497 (N_13497,N_9455,N_7383);
nor U13498 (N_13498,N_8349,N_6888);
xor U13499 (N_13499,N_5502,N_8917);
xor U13500 (N_13500,N_9033,N_6387);
and U13501 (N_13501,N_5663,N_9936);
nand U13502 (N_13502,N_6425,N_7667);
or U13503 (N_13503,N_9476,N_7225);
nand U13504 (N_13504,N_5541,N_6915);
or U13505 (N_13505,N_7477,N_9066);
nor U13506 (N_13506,N_5608,N_7068);
and U13507 (N_13507,N_9601,N_7371);
nor U13508 (N_13508,N_9886,N_8636);
or U13509 (N_13509,N_9735,N_6532);
and U13510 (N_13510,N_9079,N_6356);
and U13511 (N_13511,N_8094,N_8585);
or U13512 (N_13512,N_5346,N_7639);
nand U13513 (N_13513,N_8857,N_8436);
xor U13514 (N_13514,N_6574,N_5071);
xor U13515 (N_13515,N_5068,N_5645);
xor U13516 (N_13516,N_5944,N_7965);
and U13517 (N_13517,N_9504,N_6536);
nor U13518 (N_13518,N_5562,N_8988);
nand U13519 (N_13519,N_5981,N_5896);
and U13520 (N_13520,N_5725,N_6578);
nor U13521 (N_13521,N_5945,N_9131);
nand U13522 (N_13522,N_7593,N_7881);
and U13523 (N_13523,N_8102,N_9059);
nand U13524 (N_13524,N_5421,N_7572);
nand U13525 (N_13525,N_8197,N_6666);
nor U13526 (N_13526,N_9351,N_6161);
nor U13527 (N_13527,N_9414,N_5524);
xor U13528 (N_13528,N_7069,N_5286);
and U13529 (N_13529,N_8970,N_6582);
xnor U13530 (N_13530,N_7523,N_9499);
nand U13531 (N_13531,N_5388,N_5918);
nor U13532 (N_13532,N_5691,N_9864);
nor U13533 (N_13533,N_5289,N_9995);
nor U13534 (N_13534,N_9668,N_8888);
nor U13535 (N_13535,N_7439,N_9089);
nand U13536 (N_13536,N_8108,N_6563);
nor U13537 (N_13537,N_9207,N_6268);
xor U13538 (N_13538,N_5997,N_9935);
nand U13539 (N_13539,N_7464,N_6916);
nor U13540 (N_13540,N_6064,N_7949);
nor U13541 (N_13541,N_5692,N_6383);
nor U13542 (N_13542,N_9148,N_8791);
and U13543 (N_13543,N_7441,N_7749);
and U13544 (N_13544,N_6841,N_6524);
xor U13545 (N_13545,N_5578,N_5306);
xor U13546 (N_13546,N_8361,N_7521);
nor U13547 (N_13547,N_6842,N_7809);
nor U13548 (N_13548,N_9785,N_9040);
and U13549 (N_13549,N_5690,N_7872);
or U13550 (N_13550,N_5147,N_7576);
and U13551 (N_13551,N_8376,N_7411);
and U13552 (N_13552,N_6080,N_8264);
nand U13553 (N_13553,N_9937,N_5202);
and U13554 (N_13554,N_7254,N_6368);
nor U13555 (N_13555,N_9541,N_5295);
or U13556 (N_13556,N_6990,N_9192);
and U13557 (N_13557,N_6677,N_9667);
xor U13558 (N_13558,N_5647,N_5062);
or U13559 (N_13559,N_8066,N_8840);
nand U13560 (N_13560,N_7420,N_7078);
or U13561 (N_13561,N_5158,N_6215);
nand U13562 (N_13562,N_5654,N_7714);
xnor U13563 (N_13563,N_6847,N_5726);
nor U13564 (N_13564,N_8409,N_6812);
nor U13565 (N_13565,N_7915,N_5837);
nor U13566 (N_13566,N_6260,N_9066);
nand U13567 (N_13567,N_9782,N_9977);
nand U13568 (N_13568,N_6172,N_5847);
and U13569 (N_13569,N_9406,N_5834);
xnor U13570 (N_13570,N_9355,N_7762);
xnor U13571 (N_13571,N_6677,N_5999);
nand U13572 (N_13572,N_8445,N_5623);
or U13573 (N_13573,N_7423,N_9355);
nor U13574 (N_13574,N_7295,N_5619);
nand U13575 (N_13575,N_8105,N_6319);
or U13576 (N_13576,N_8616,N_6165);
nand U13577 (N_13577,N_5810,N_5983);
nor U13578 (N_13578,N_7973,N_9399);
nand U13579 (N_13579,N_7603,N_5834);
xor U13580 (N_13580,N_6145,N_9125);
nand U13581 (N_13581,N_8212,N_9228);
nor U13582 (N_13582,N_5622,N_8926);
nand U13583 (N_13583,N_8065,N_7718);
nand U13584 (N_13584,N_5346,N_9896);
xnor U13585 (N_13585,N_9020,N_7670);
nand U13586 (N_13586,N_9282,N_5223);
nand U13587 (N_13587,N_6800,N_9397);
nand U13588 (N_13588,N_7477,N_7120);
nor U13589 (N_13589,N_5625,N_9209);
or U13590 (N_13590,N_6968,N_7602);
xnor U13591 (N_13591,N_6775,N_6535);
nand U13592 (N_13592,N_9059,N_8227);
xor U13593 (N_13593,N_8032,N_5063);
and U13594 (N_13594,N_5909,N_6783);
xnor U13595 (N_13595,N_7850,N_5385);
nor U13596 (N_13596,N_5945,N_9611);
and U13597 (N_13597,N_6359,N_5245);
nor U13598 (N_13598,N_7587,N_9933);
or U13599 (N_13599,N_9961,N_7188);
nand U13600 (N_13600,N_8458,N_5790);
nand U13601 (N_13601,N_7486,N_6737);
and U13602 (N_13602,N_5571,N_7517);
or U13603 (N_13603,N_9101,N_7766);
xor U13604 (N_13604,N_5858,N_6516);
and U13605 (N_13605,N_8839,N_6572);
and U13606 (N_13606,N_5489,N_9292);
or U13607 (N_13607,N_7150,N_8783);
nor U13608 (N_13608,N_9088,N_6726);
nand U13609 (N_13609,N_7247,N_5745);
nor U13610 (N_13610,N_7450,N_8331);
and U13611 (N_13611,N_7878,N_7750);
xor U13612 (N_13612,N_9233,N_6962);
or U13613 (N_13613,N_6923,N_8839);
and U13614 (N_13614,N_7743,N_5414);
nor U13615 (N_13615,N_7137,N_8502);
and U13616 (N_13616,N_8308,N_8320);
or U13617 (N_13617,N_7003,N_5920);
nand U13618 (N_13618,N_8452,N_7757);
nand U13619 (N_13619,N_8540,N_9048);
and U13620 (N_13620,N_7751,N_6832);
nand U13621 (N_13621,N_5125,N_7719);
xnor U13622 (N_13622,N_6775,N_8621);
nand U13623 (N_13623,N_6265,N_5715);
nor U13624 (N_13624,N_8753,N_8827);
or U13625 (N_13625,N_5873,N_9757);
nand U13626 (N_13626,N_8529,N_8824);
and U13627 (N_13627,N_6391,N_7639);
xor U13628 (N_13628,N_7219,N_6548);
nor U13629 (N_13629,N_8361,N_9525);
and U13630 (N_13630,N_5856,N_5258);
nor U13631 (N_13631,N_5652,N_7922);
or U13632 (N_13632,N_9396,N_7050);
or U13633 (N_13633,N_7357,N_8127);
or U13634 (N_13634,N_7918,N_8164);
or U13635 (N_13635,N_9040,N_8098);
nand U13636 (N_13636,N_6439,N_5379);
or U13637 (N_13637,N_7130,N_8252);
nor U13638 (N_13638,N_9432,N_5244);
and U13639 (N_13639,N_8808,N_5009);
nor U13640 (N_13640,N_7134,N_7799);
nand U13641 (N_13641,N_5372,N_8368);
and U13642 (N_13642,N_9198,N_8179);
and U13643 (N_13643,N_6286,N_8429);
nor U13644 (N_13644,N_5760,N_7075);
nor U13645 (N_13645,N_6503,N_9582);
nor U13646 (N_13646,N_8524,N_7639);
xnor U13647 (N_13647,N_6714,N_5721);
nor U13648 (N_13648,N_8786,N_8007);
nand U13649 (N_13649,N_7296,N_5890);
nand U13650 (N_13650,N_7752,N_9299);
and U13651 (N_13651,N_7418,N_5811);
and U13652 (N_13652,N_6219,N_8244);
and U13653 (N_13653,N_9451,N_9675);
xor U13654 (N_13654,N_6040,N_5480);
or U13655 (N_13655,N_7203,N_7584);
or U13656 (N_13656,N_9465,N_8190);
xor U13657 (N_13657,N_9153,N_6171);
or U13658 (N_13658,N_5514,N_8743);
nand U13659 (N_13659,N_7440,N_9175);
nor U13660 (N_13660,N_6418,N_6551);
nand U13661 (N_13661,N_8815,N_9111);
or U13662 (N_13662,N_7703,N_7455);
or U13663 (N_13663,N_5606,N_7219);
nor U13664 (N_13664,N_6388,N_7196);
or U13665 (N_13665,N_9392,N_5882);
xor U13666 (N_13666,N_5251,N_8370);
and U13667 (N_13667,N_5858,N_8478);
xnor U13668 (N_13668,N_7492,N_8210);
and U13669 (N_13669,N_8312,N_7998);
xor U13670 (N_13670,N_5154,N_8533);
or U13671 (N_13671,N_7219,N_6131);
nor U13672 (N_13672,N_9471,N_9277);
and U13673 (N_13673,N_5936,N_9669);
nand U13674 (N_13674,N_9978,N_7358);
nand U13675 (N_13675,N_8545,N_5050);
or U13676 (N_13676,N_9899,N_7025);
xor U13677 (N_13677,N_9227,N_5840);
nor U13678 (N_13678,N_6997,N_5863);
or U13679 (N_13679,N_9455,N_7917);
nor U13680 (N_13680,N_6114,N_9709);
nor U13681 (N_13681,N_9335,N_7122);
and U13682 (N_13682,N_7045,N_9557);
or U13683 (N_13683,N_6795,N_6345);
or U13684 (N_13684,N_5440,N_8299);
nor U13685 (N_13685,N_7999,N_5540);
or U13686 (N_13686,N_7985,N_5556);
and U13687 (N_13687,N_8773,N_9874);
nand U13688 (N_13688,N_7507,N_5454);
nor U13689 (N_13689,N_6980,N_9259);
or U13690 (N_13690,N_8632,N_6224);
and U13691 (N_13691,N_9826,N_6409);
nand U13692 (N_13692,N_5946,N_5592);
or U13693 (N_13693,N_9490,N_6479);
nor U13694 (N_13694,N_6585,N_6255);
nor U13695 (N_13695,N_5193,N_8934);
or U13696 (N_13696,N_8113,N_6927);
or U13697 (N_13697,N_6500,N_8342);
and U13698 (N_13698,N_8460,N_6636);
or U13699 (N_13699,N_8835,N_7166);
nor U13700 (N_13700,N_5465,N_6962);
nor U13701 (N_13701,N_9591,N_9939);
and U13702 (N_13702,N_7973,N_9716);
and U13703 (N_13703,N_8070,N_6268);
nor U13704 (N_13704,N_6187,N_9818);
or U13705 (N_13705,N_9512,N_7014);
nand U13706 (N_13706,N_6876,N_8747);
xnor U13707 (N_13707,N_9169,N_7571);
nor U13708 (N_13708,N_8184,N_8403);
and U13709 (N_13709,N_8671,N_9611);
or U13710 (N_13710,N_9537,N_9038);
xor U13711 (N_13711,N_8976,N_8127);
or U13712 (N_13712,N_7223,N_7087);
nor U13713 (N_13713,N_7996,N_7210);
nand U13714 (N_13714,N_8026,N_5512);
nand U13715 (N_13715,N_8177,N_6953);
or U13716 (N_13716,N_6890,N_7170);
nand U13717 (N_13717,N_9897,N_8700);
nand U13718 (N_13718,N_6221,N_8881);
xor U13719 (N_13719,N_7506,N_8908);
nor U13720 (N_13720,N_9884,N_8319);
nor U13721 (N_13721,N_9008,N_8445);
nand U13722 (N_13722,N_5969,N_7905);
or U13723 (N_13723,N_5196,N_8376);
or U13724 (N_13724,N_9736,N_8061);
xnor U13725 (N_13725,N_8662,N_9073);
nor U13726 (N_13726,N_7884,N_8165);
xnor U13727 (N_13727,N_8845,N_9962);
xnor U13728 (N_13728,N_9946,N_8763);
nor U13729 (N_13729,N_8612,N_6481);
and U13730 (N_13730,N_9584,N_8022);
and U13731 (N_13731,N_7045,N_6387);
nand U13732 (N_13732,N_9729,N_8456);
xnor U13733 (N_13733,N_9144,N_9399);
or U13734 (N_13734,N_9101,N_7519);
nand U13735 (N_13735,N_7503,N_8951);
and U13736 (N_13736,N_5839,N_5101);
or U13737 (N_13737,N_8699,N_6806);
nand U13738 (N_13738,N_5339,N_9343);
nor U13739 (N_13739,N_9607,N_8041);
and U13740 (N_13740,N_8899,N_9679);
nor U13741 (N_13741,N_9938,N_6102);
or U13742 (N_13742,N_6931,N_6897);
and U13743 (N_13743,N_5513,N_5594);
and U13744 (N_13744,N_7894,N_9824);
xnor U13745 (N_13745,N_5541,N_8492);
and U13746 (N_13746,N_9396,N_5857);
xnor U13747 (N_13747,N_7230,N_5256);
nor U13748 (N_13748,N_8150,N_6093);
and U13749 (N_13749,N_7426,N_9146);
xor U13750 (N_13750,N_7184,N_5446);
or U13751 (N_13751,N_8958,N_6553);
and U13752 (N_13752,N_8768,N_8546);
nand U13753 (N_13753,N_7019,N_6201);
and U13754 (N_13754,N_6785,N_8051);
xnor U13755 (N_13755,N_5837,N_6561);
nand U13756 (N_13756,N_5249,N_6641);
xor U13757 (N_13757,N_7084,N_7426);
nor U13758 (N_13758,N_9982,N_6913);
and U13759 (N_13759,N_9807,N_7793);
xor U13760 (N_13760,N_8732,N_5736);
or U13761 (N_13761,N_7589,N_6734);
and U13762 (N_13762,N_9992,N_8282);
nand U13763 (N_13763,N_9431,N_7849);
or U13764 (N_13764,N_5437,N_7833);
xnor U13765 (N_13765,N_7877,N_7385);
nand U13766 (N_13766,N_6828,N_6251);
nor U13767 (N_13767,N_5404,N_5368);
or U13768 (N_13768,N_6964,N_7149);
nand U13769 (N_13769,N_7207,N_5118);
xnor U13770 (N_13770,N_8626,N_7493);
or U13771 (N_13771,N_8777,N_7404);
and U13772 (N_13772,N_6373,N_9521);
nand U13773 (N_13773,N_5173,N_6482);
nor U13774 (N_13774,N_6079,N_6687);
nand U13775 (N_13775,N_6140,N_7597);
nand U13776 (N_13776,N_5365,N_9093);
nor U13777 (N_13777,N_5250,N_9900);
xor U13778 (N_13778,N_8652,N_9567);
and U13779 (N_13779,N_5109,N_5304);
and U13780 (N_13780,N_6578,N_6147);
nand U13781 (N_13781,N_7377,N_8766);
or U13782 (N_13782,N_9299,N_8200);
xor U13783 (N_13783,N_6949,N_5530);
nand U13784 (N_13784,N_8930,N_5297);
nand U13785 (N_13785,N_5582,N_8567);
nor U13786 (N_13786,N_5025,N_6092);
xnor U13787 (N_13787,N_8265,N_5848);
xor U13788 (N_13788,N_8227,N_6785);
or U13789 (N_13789,N_6820,N_7723);
or U13790 (N_13790,N_8726,N_7396);
xnor U13791 (N_13791,N_6272,N_9728);
or U13792 (N_13792,N_5528,N_9680);
nor U13793 (N_13793,N_7853,N_6961);
or U13794 (N_13794,N_7511,N_8558);
and U13795 (N_13795,N_7794,N_8277);
nor U13796 (N_13796,N_5703,N_6166);
nor U13797 (N_13797,N_9813,N_7658);
xor U13798 (N_13798,N_9063,N_6438);
nor U13799 (N_13799,N_6827,N_9849);
nand U13800 (N_13800,N_6396,N_7134);
xor U13801 (N_13801,N_6954,N_7210);
and U13802 (N_13802,N_6131,N_7787);
or U13803 (N_13803,N_9822,N_7548);
or U13804 (N_13804,N_7133,N_7235);
xnor U13805 (N_13805,N_6135,N_6122);
or U13806 (N_13806,N_9940,N_5473);
or U13807 (N_13807,N_9747,N_9141);
or U13808 (N_13808,N_6203,N_6922);
xor U13809 (N_13809,N_7279,N_7387);
or U13810 (N_13810,N_8021,N_8181);
xnor U13811 (N_13811,N_8536,N_5096);
nand U13812 (N_13812,N_9990,N_5562);
xor U13813 (N_13813,N_9613,N_9183);
xnor U13814 (N_13814,N_7188,N_5992);
and U13815 (N_13815,N_9746,N_9622);
xnor U13816 (N_13816,N_6172,N_7050);
and U13817 (N_13817,N_9410,N_8961);
xnor U13818 (N_13818,N_6713,N_6946);
xor U13819 (N_13819,N_7337,N_6308);
nand U13820 (N_13820,N_6297,N_7039);
xnor U13821 (N_13821,N_8693,N_6310);
nand U13822 (N_13822,N_5728,N_5376);
nor U13823 (N_13823,N_7766,N_6988);
or U13824 (N_13824,N_5871,N_9222);
and U13825 (N_13825,N_7292,N_8552);
and U13826 (N_13826,N_5839,N_5006);
xor U13827 (N_13827,N_9332,N_6684);
nand U13828 (N_13828,N_5798,N_6448);
xor U13829 (N_13829,N_9597,N_5460);
and U13830 (N_13830,N_8863,N_5915);
nor U13831 (N_13831,N_9217,N_7098);
nand U13832 (N_13832,N_8145,N_9391);
and U13833 (N_13833,N_5619,N_8336);
xnor U13834 (N_13834,N_5747,N_6486);
xor U13835 (N_13835,N_7675,N_8723);
or U13836 (N_13836,N_9399,N_7118);
or U13837 (N_13837,N_8390,N_8544);
or U13838 (N_13838,N_5657,N_6215);
xnor U13839 (N_13839,N_6213,N_6235);
or U13840 (N_13840,N_5400,N_6844);
nand U13841 (N_13841,N_5714,N_5968);
nor U13842 (N_13842,N_5928,N_7422);
or U13843 (N_13843,N_5746,N_7455);
and U13844 (N_13844,N_8284,N_7808);
and U13845 (N_13845,N_7889,N_5205);
nand U13846 (N_13846,N_7279,N_6592);
nand U13847 (N_13847,N_5927,N_7624);
nand U13848 (N_13848,N_9447,N_7023);
nor U13849 (N_13849,N_8015,N_9385);
and U13850 (N_13850,N_5998,N_8282);
and U13851 (N_13851,N_9780,N_8983);
nor U13852 (N_13852,N_9177,N_7490);
or U13853 (N_13853,N_6807,N_8590);
nor U13854 (N_13854,N_6459,N_9247);
xor U13855 (N_13855,N_7532,N_6803);
nor U13856 (N_13856,N_6220,N_9461);
or U13857 (N_13857,N_9807,N_7311);
nor U13858 (N_13858,N_8534,N_9482);
nand U13859 (N_13859,N_6700,N_6232);
nand U13860 (N_13860,N_5121,N_8289);
and U13861 (N_13861,N_9713,N_7871);
nor U13862 (N_13862,N_9638,N_7965);
and U13863 (N_13863,N_8183,N_7688);
xor U13864 (N_13864,N_9000,N_7193);
xor U13865 (N_13865,N_6274,N_8849);
nor U13866 (N_13866,N_9655,N_9632);
nor U13867 (N_13867,N_9448,N_7862);
xor U13868 (N_13868,N_8035,N_7818);
nand U13869 (N_13869,N_7288,N_8156);
nand U13870 (N_13870,N_7817,N_6861);
nor U13871 (N_13871,N_9164,N_9116);
xor U13872 (N_13872,N_5410,N_8810);
or U13873 (N_13873,N_8571,N_8654);
and U13874 (N_13874,N_8484,N_7959);
nand U13875 (N_13875,N_6826,N_7830);
nand U13876 (N_13876,N_5985,N_8225);
xnor U13877 (N_13877,N_9075,N_7277);
nand U13878 (N_13878,N_7777,N_7812);
and U13879 (N_13879,N_7213,N_7746);
or U13880 (N_13880,N_7772,N_9555);
nand U13881 (N_13881,N_6348,N_8465);
and U13882 (N_13882,N_6325,N_6108);
or U13883 (N_13883,N_9506,N_8391);
and U13884 (N_13884,N_9778,N_7940);
and U13885 (N_13885,N_5354,N_6186);
xnor U13886 (N_13886,N_8275,N_5084);
and U13887 (N_13887,N_7078,N_8126);
or U13888 (N_13888,N_5734,N_5717);
and U13889 (N_13889,N_8649,N_7451);
nand U13890 (N_13890,N_5437,N_7860);
nor U13891 (N_13891,N_7213,N_8046);
nand U13892 (N_13892,N_6137,N_9036);
nor U13893 (N_13893,N_8237,N_8763);
xor U13894 (N_13894,N_9702,N_5575);
xor U13895 (N_13895,N_8949,N_7743);
nand U13896 (N_13896,N_9224,N_7890);
nand U13897 (N_13897,N_8851,N_5206);
nand U13898 (N_13898,N_8003,N_8318);
nand U13899 (N_13899,N_7662,N_8572);
xnor U13900 (N_13900,N_7838,N_8428);
nand U13901 (N_13901,N_5343,N_7647);
nor U13902 (N_13902,N_5296,N_5323);
and U13903 (N_13903,N_6784,N_8172);
xnor U13904 (N_13904,N_9595,N_8106);
nor U13905 (N_13905,N_6485,N_7387);
or U13906 (N_13906,N_7628,N_8080);
nor U13907 (N_13907,N_9758,N_8291);
nor U13908 (N_13908,N_7367,N_8920);
nor U13909 (N_13909,N_9884,N_9760);
and U13910 (N_13910,N_8173,N_9010);
and U13911 (N_13911,N_9519,N_8049);
nor U13912 (N_13912,N_6900,N_6796);
nor U13913 (N_13913,N_7095,N_7795);
nand U13914 (N_13914,N_7351,N_5782);
and U13915 (N_13915,N_7476,N_6510);
nor U13916 (N_13916,N_7312,N_5372);
xnor U13917 (N_13917,N_8086,N_5653);
or U13918 (N_13918,N_8798,N_8540);
nand U13919 (N_13919,N_5682,N_9813);
and U13920 (N_13920,N_6103,N_5553);
or U13921 (N_13921,N_8183,N_9389);
or U13922 (N_13922,N_5753,N_7683);
and U13923 (N_13923,N_9000,N_5333);
nand U13924 (N_13924,N_8894,N_5370);
nor U13925 (N_13925,N_6440,N_7042);
and U13926 (N_13926,N_6067,N_8778);
xor U13927 (N_13927,N_6178,N_5058);
nand U13928 (N_13928,N_9851,N_5632);
nand U13929 (N_13929,N_5236,N_9589);
and U13930 (N_13930,N_6621,N_8053);
nor U13931 (N_13931,N_8875,N_5356);
nor U13932 (N_13932,N_6614,N_7384);
and U13933 (N_13933,N_7489,N_9776);
or U13934 (N_13934,N_6241,N_6663);
nor U13935 (N_13935,N_8518,N_5311);
xor U13936 (N_13936,N_5981,N_5362);
nor U13937 (N_13937,N_8792,N_8624);
xnor U13938 (N_13938,N_5797,N_5220);
or U13939 (N_13939,N_8743,N_6647);
xor U13940 (N_13940,N_5913,N_9966);
nor U13941 (N_13941,N_9937,N_9390);
xor U13942 (N_13942,N_8340,N_9799);
and U13943 (N_13943,N_6368,N_9891);
nand U13944 (N_13944,N_8020,N_6151);
nand U13945 (N_13945,N_5100,N_7788);
or U13946 (N_13946,N_5188,N_8636);
nand U13947 (N_13947,N_7670,N_5908);
xor U13948 (N_13948,N_6132,N_5339);
and U13949 (N_13949,N_5750,N_7305);
or U13950 (N_13950,N_5623,N_8706);
or U13951 (N_13951,N_8217,N_6089);
nand U13952 (N_13952,N_7358,N_9557);
nor U13953 (N_13953,N_9791,N_6320);
nor U13954 (N_13954,N_6745,N_9921);
or U13955 (N_13955,N_8411,N_9927);
nand U13956 (N_13956,N_7969,N_8010);
and U13957 (N_13957,N_9337,N_7459);
nor U13958 (N_13958,N_9116,N_7329);
nand U13959 (N_13959,N_9993,N_8117);
nand U13960 (N_13960,N_7595,N_9364);
xor U13961 (N_13961,N_5729,N_8082);
xor U13962 (N_13962,N_7726,N_6100);
xor U13963 (N_13963,N_7104,N_5341);
and U13964 (N_13964,N_7342,N_6779);
or U13965 (N_13965,N_9249,N_9216);
nor U13966 (N_13966,N_9644,N_9602);
or U13967 (N_13967,N_5947,N_5915);
nor U13968 (N_13968,N_5097,N_9194);
nand U13969 (N_13969,N_7504,N_8616);
and U13970 (N_13970,N_5533,N_8295);
nand U13971 (N_13971,N_6448,N_7328);
and U13972 (N_13972,N_9343,N_6622);
nor U13973 (N_13973,N_9600,N_5084);
and U13974 (N_13974,N_9299,N_8825);
xnor U13975 (N_13975,N_8355,N_9696);
and U13976 (N_13976,N_7335,N_6104);
or U13977 (N_13977,N_9182,N_7724);
and U13978 (N_13978,N_7752,N_9172);
and U13979 (N_13979,N_9300,N_9000);
and U13980 (N_13980,N_9636,N_9316);
xor U13981 (N_13981,N_8688,N_6314);
and U13982 (N_13982,N_6450,N_5296);
nand U13983 (N_13983,N_6155,N_8141);
or U13984 (N_13984,N_8140,N_9148);
or U13985 (N_13985,N_7902,N_7422);
nor U13986 (N_13986,N_8768,N_5929);
nand U13987 (N_13987,N_5882,N_9352);
or U13988 (N_13988,N_9173,N_9899);
or U13989 (N_13989,N_5468,N_5204);
and U13990 (N_13990,N_7347,N_8725);
xor U13991 (N_13991,N_8934,N_7217);
nand U13992 (N_13992,N_7182,N_6103);
or U13993 (N_13993,N_6584,N_8092);
nand U13994 (N_13994,N_9261,N_6134);
nand U13995 (N_13995,N_6350,N_9562);
or U13996 (N_13996,N_7025,N_6265);
or U13997 (N_13997,N_6385,N_5470);
nand U13998 (N_13998,N_7300,N_7037);
nand U13999 (N_13999,N_9243,N_9965);
nor U14000 (N_14000,N_7656,N_7435);
and U14001 (N_14001,N_5076,N_6445);
nand U14002 (N_14002,N_6627,N_8926);
or U14003 (N_14003,N_5104,N_9437);
nor U14004 (N_14004,N_6115,N_5992);
nor U14005 (N_14005,N_6159,N_8315);
nor U14006 (N_14006,N_6656,N_9453);
or U14007 (N_14007,N_6973,N_9300);
nand U14008 (N_14008,N_5871,N_6891);
and U14009 (N_14009,N_8732,N_8475);
or U14010 (N_14010,N_5192,N_5559);
and U14011 (N_14011,N_7254,N_6757);
or U14012 (N_14012,N_8586,N_5784);
nor U14013 (N_14013,N_7880,N_7087);
nand U14014 (N_14014,N_5638,N_7332);
or U14015 (N_14015,N_8155,N_9049);
nor U14016 (N_14016,N_6637,N_9406);
nand U14017 (N_14017,N_5609,N_8827);
nand U14018 (N_14018,N_9592,N_5539);
nand U14019 (N_14019,N_5585,N_9771);
nor U14020 (N_14020,N_8059,N_7547);
xnor U14021 (N_14021,N_6498,N_8805);
or U14022 (N_14022,N_7573,N_9184);
nor U14023 (N_14023,N_8016,N_9454);
nor U14024 (N_14024,N_9445,N_7084);
nand U14025 (N_14025,N_7784,N_8648);
xor U14026 (N_14026,N_9967,N_9997);
xnor U14027 (N_14027,N_7104,N_9802);
and U14028 (N_14028,N_6576,N_9461);
and U14029 (N_14029,N_7013,N_8369);
or U14030 (N_14030,N_7381,N_6150);
nand U14031 (N_14031,N_7210,N_7500);
nand U14032 (N_14032,N_9459,N_5897);
or U14033 (N_14033,N_6554,N_5053);
and U14034 (N_14034,N_9647,N_5983);
or U14035 (N_14035,N_7029,N_9918);
nor U14036 (N_14036,N_9011,N_9496);
nor U14037 (N_14037,N_6489,N_7070);
or U14038 (N_14038,N_5147,N_8832);
and U14039 (N_14039,N_7521,N_5319);
nand U14040 (N_14040,N_5565,N_7129);
or U14041 (N_14041,N_6131,N_9507);
nor U14042 (N_14042,N_9764,N_7746);
nand U14043 (N_14043,N_8868,N_6388);
nor U14044 (N_14044,N_5023,N_5283);
and U14045 (N_14045,N_9525,N_5642);
nand U14046 (N_14046,N_7048,N_7886);
or U14047 (N_14047,N_6458,N_7834);
or U14048 (N_14048,N_8145,N_6583);
nand U14049 (N_14049,N_7800,N_7614);
nor U14050 (N_14050,N_7410,N_8864);
nand U14051 (N_14051,N_7719,N_6725);
xnor U14052 (N_14052,N_5483,N_9810);
and U14053 (N_14053,N_9018,N_9855);
or U14054 (N_14054,N_6612,N_9300);
nor U14055 (N_14055,N_8224,N_7839);
nand U14056 (N_14056,N_5499,N_7627);
nand U14057 (N_14057,N_6544,N_5904);
and U14058 (N_14058,N_7127,N_5883);
nor U14059 (N_14059,N_7016,N_8574);
and U14060 (N_14060,N_5676,N_7933);
nand U14061 (N_14061,N_7550,N_8918);
or U14062 (N_14062,N_9321,N_8333);
xnor U14063 (N_14063,N_8130,N_9185);
nor U14064 (N_14064,N_9626,N_6285);
nor U14065 (N_14065,N_6957,N_9105);
xnor U14066 (N_14066,N_8813,N_5197);
xor U14067 (N_14067,N_5935,N_8165);
nor U14068 (N_14068,N_8555,N_8367);
nor U14069 (N_14069,N_6437,N_6349);
xor U14070 (N_14070,N_6056,N_6969);
nand U14071 (N_14071,N_8577,N_8556);
or U14072 (N_14072,N_7783,N_6366);
and U14073 (N_14073,N_5047,N_6275);
nor U14074 (N_14074,N_7518,N_8591);
or U14075 (N_14075,N_8546,N_9032);
nand U14076 (N_14076,N_5866,N_8084);
nand U14077 (N_14077,N_8612,N_7759);
and U14078 (N_14078,N_5977,N_7216);
nor U14079 (N_14079,N_9170,N_5755);
nor U14080 (N_14080,N_6619,N_8272);
xnor U14081 (N_14081,N_5969,N_8122);
or U14082 (N_14082,N_8941,N_5677);
or U14083 (N_14083,N_5049,N_5026);
or U14084 (N_14084,N_6300,N_5678);
and U14085 (N_14085,N_9670,N_7072);
or U14086 (N_14086,N_8438,N_8584);
and U14087 (N_14087,N_6248,N_5575);
and U14088 (N_14088,N_6906,N_9560);
nand U14089 (N_14089,N_7701,N_6443);
or U14090 (N_14090,N_5947,N_6105);
nor U14091 (N_14091,N_6537,N_5717);
xnor U14092 (N_14092,N_6225,N_8512);
nor U14093 (N_14093,N_8698,N_5191);
or U14094 (N_14094,N_6852,N_6662);
nor U14095 (N_14095,N_7507,N_6199);
or U14096 (N_14096,N_9949,N_6106);
nor U14097 (N_14097,N_6464,N_6951);
nor U14098 (N_14098,N_6059,N_8954);
nor U14099 (N_14099,N_6513,N_8051);
or U14100 (N_14100,N_7772,N_9366);
nand U14101 (N_14101,N_9857,N_8978);
nor U14102 (N_14102,N_7507,N_9496);
xor U14103 (N_14103,N_8623,N_7952);
or U14104 (N_14104,N_7728,N_7285);
xor U14105 (N_14105,N_9976,N_8987);
nand U14106 (N_14106,N_8402,N_6420);
or U14107 (N_14107,N_8874,N_9475);
nor U14108 (N_14108,N_6865,N_6108);
or U14109 (N_14109,N_7763,N_5471);
and U14110 (N_14110,N_7091,N_9419);
or U14111 (N_14111,N_8876,N_9870);
xnor U14112 (N_14112,N_9781,N_8576);
nor U14113 (N_14113,N_9096,N_8116);
nor U14114 (N_14114,N_7383,N_9415);
or U14115 (N_14115,N_8305,N_5786);
nand U14116 (N_14116,N_6372,N_9150);
nor U14117 (N_14117,N_6146,N_8394);
or U14118 (N_14118,N_9009,N_7213);
xnor U14119 (N_14119,N_8508,N_9992);
and U14120 (N_14120,N_7686,N_8488);
xor U14121 (N_14121,N_9333,N_6935);
or U14122 (N_14122,N_9261,N_5205);
and U14123 (N_14123,N_9932,N_7133);
and U14124 (N_14124,N_6093,N_5949);
and U14125 (N_14125,N_7579,N_9430);
xnor U14126 (N_14126,N_9994,N_5998);
and U14127 (N_14127,N_8335,N_6668);
nor U14128 (N_14128,N_7182,N_9664);
and U14129 (N_14129,N_6542,N_6833);
nor U14130 (N_14130,N_6239,N_6335);
and U14131 (N_14131,N_7705,N_8699);
or U14132 (N_14132,N_6827,N_8017);
and U14133 (N_14133,N_8977,N_9101);
or U14134 (N_14134,N_7711,N_7554);
nor U14135 (N_14135,N_7713,N_7139);
or U14136 (N_14136,N_8886,N_5697);
or U14137 (N_14137,N_9219,N_7862);
xnor U14138 (N_14138,N_5902,N_8400);
or U14139 (N_14139,N_8175,N_7031);
nand U14140 (N_14140,N_7673,N_9840);
nand U14141 (N_14141,N_8322,N_5888);
nand U14142 (N_14142,N_8849,N_7391);
nand U14143 (N_14143,N_6227,N_5341);
nand U14144 (N_14144,N_9598,N_6649);
nand U14145 (N_14145,N_5183,N_8637);
and U14146 (N_14146,N_9695,N_6742);
or U14147 (N_14147,N_7795,N_5508);
nor U14148 (N_14148,N_6510,N_9050);
and U14149 (N_14149,N_5962,N_8506);
and U14150 (N_14150,N_8504,N_8678);
nor U14151 (N_14151,N_9135,N_7419);
and U14152 (N_14152,N_7857,N_6084);
nand U14153 (N_14153,N_5907,N_7000);
and U14154 (N_14154,N_9478,N_6355);
xor U14155 (N_14155,N_9931,N_8526);
and U14156 (N_14156,N_5262,N_5891);
xor U14157 (N_14157,N_6947,N_5645);
nand U14158 (N_14158,N_7942,N_8851);
nand U14159 (N_14159,N_8270,N_5033);
xnor U14160 (N_14160,N_7215,N_5930);
and U14161 (N_14161,N_6043,N_9963);
nand U14162 (N_14162,N_9007,N_9205);
or U14163 (N_14163,N_5026,N_6270);
nand U14164 (N_14164,N_8341,N_7057);
xor U14165 (N_14165,N_5727,N_6050);
nand U14166 (N_14166,N_9334,N_5137);
nor U14167 (N_14167,N_8892,N_6703);
or U14168 (N_14168,N_6146,N_6348);
and U14169 (N_14169,N_7668,N_7120);
or U14170 (N_14170,N_8367,N_5003);
nand U14171 (N_14171,N_7248,N_9401);
xnor U14172 (N_14172,N_7514,N_6070);
nor U14173 (N_14173,N_8167,N_6692);
nor U14174 (N_14174,N_7846,N_9626);
xor U14175 (N_14175,N_9594,N_9051);
nand U14176 (N_14176,N_8160,N_9908);
nand U14177 (N_14177,N_6176,N_8133);
nand U14178 (N_14178,N_7068,N_7365);
or U14179 (N_14179,N_7031,N_9441);
nand U14180 (N_14180,N_8177,N_9096);
or U14181 (N_14181,N_6982,N_8661);
or U14182 (N_14182,N_8217,N_5379);
nor U14183 (N_14183,N_5753,N_8650);
or U14184 (N_14184,N_9440,N_8469);
nand U14185 (N_14185,N_6257,N_9891);
or U14186 (N_14186,N_7688,N_9535);
or U14187 (N_14187,N_6161,N_6513);
nand U14188 (N_14188,N_5751,N_9867);
or U14189 (N_14189,N_7298,N_8279);
or U14190 (N_14190,N_9666,N_5589);
and U14191 (N_14191,N_7781,N_9148);
nor U14192 (N_14192,N_7991,N_6006);
xnor U14193 (N_14193,N_6278,N_8676);
nor U14194 (N_14194,N_7145,N_5242);
nand U14195 (N_14195,N_9747,N_8174);
and U14196 (N_14196,N_6159,N_7450);
nand U14197 (N_14197,N_7945,N_7379);
xor U14198 (N_14198,N_7136,N_5369);
nand U14199 (N_14199,N_7993,N_9011);
nor U14200 (N_14200,N_6642,N_7327);
or U14201 (N_14201,N_7749,N_5362);
and U14202 (N_14202,N_9604,N_6841);
xnor U14203 (N_14203,N_5104,N_9611);
and U14204 (N_14204,N_7027,N_9946);
nor U14205 (N_14205,N_9133,N_7071);
or U14206 (N_14206,N_9341,N_9535);
nor U14207 (N_14207,N_8187,N_7675);
nand U14208 (N_14208,N_8938,N_5311);
nor U14209 (N_14209,N_9753,N_8103);
and U14210 (N_14210,N_9375,N_5477);
nand U14211 (N_14211,N_5080,N_6979);
nand U14212 (N_14212,N_8183,N_5600);
xor U14213 (N_14213,N_7260,N_7167);
nand U14214 (N_14214,N_5864,N_6781);
nand U14215 (N_14215,N_5048,N_9246);
xor U14216 (N_14216,N_7559,N_7616);
nor U14217 (N_14217,N_6751,N_8071);
and U14218 (N_14218,N_8009,N_7881);
xnor U14219 (N_14219,N_5761,N_8581);
nand U14220 (N_14220,N_7984,N_9433);
xnor U14221 (N_14221,N_9636,N_6033);
or U14222 (N_14222,N_8195,N_7255);
or U14223 (N_14223,N_8129,N_7041);
xor U14224 (N_14224,N_5100,N_7413);
and U14225 (N_14225,N_8247,N_8858);
and U14226 (N_14226,N_9947,N_8358);
nand U14227 (N_14227,N_8565,N_9832);
xnor U14228 (N_14228,N_5082,N_8400);
nand U14229 (N_14229,N_6066,N_8969);
nand U14230 (N_14230,N_9651,N_9762);
nor U14231 (N_14231,N_9691,N_7030);
and U14232 (N_14232,N_5813,N_7521);
xor U14233 (N_14233,N_8912,N_5747);
and U14234 (N_14234,N_8623,N_6569);
and U14235 (N_14235,N_9597,N_7804);
or U14236 (N_14236,N_9366,N_7620);
xor U14237 (N_14237,N_9957,N_5208);
nand U14238 (N_14238,N_8433,N_5594);
xnor U14239 (N_14239,N_5583,N_9006);
xnor U14240 (N_14240,N_5978,N_7420);
and U14241 (N_14241,N_5488,N_9592);
nor U14242 (N_14242,N_5915,N_8464);
xnor U14243 (N_14243,N_5288,N_5492);
nand U14244 (N_14244,N_6004,N_9894);
nand U14245 (N_14245,N_9576,N_7498);
nor U14246 (N_14246,N_9624,N_6929);
nor U14247 (N_14247,N_7009,N_5806);
nand U14248 (N_14248,N_6386,N_5558);
xor U14249 (N_14249,N_9200,N_7331);
xor U14250 (N_14250,N_8010,N_8105);
and U14251 (N_14251,N_5890,N_6041);
and U14252 (N_14252,N_5004,N_7438);
or U14253 (N_14253,N_8024,N_5051);
nor U14254 (N_14254,N_5958,N_5558);
and U14255 (N_14255,N_7767,N_5097);
nand U14256 (N_14256,N_5005,N_8700);
or U14257 (N_14257,N_7131,N_8543);
nor U14258 (N_14258,N_6586,N_8921);
or U14259 (N_14259,N_6642,N_7371);
nand U14260 (N_14260,N_6500,N_9650);
nand U14261 (N_14261,N_6149,N_6013);
xnor U14262 (N_14262,N_6806,N_7037);
or U14263 (N_14263,N_8045,N_6750);
nand U14264 (N_14264,N_9849,N_5846);
nand U14265 (N_14265,N_7624,N_9622);
and U14266 (N_14266,N_7286,N_7413);
xnor U14267 (N_14267,N_6047,N_9197);
or U14268 (N_14268,N_6688,N_6986);
or U14269 (N_14269,N_6162,N_7293);
or U14270 (N_14270,N_7776,N_8799);
nand U14271 (N_14271,N_9179,N_5467);
and U14272 (N_14272,N_8183,N_9801);
xor U14273 (N_14273,N_5780,N_9726);
nor U14274 (N_14274,N_5315,N_9498);
nand U14275 (N_14275,N_5373,N_8762);
nand U14276 (N_14276,N_9657,N_6499);
nor U14277 (N_14277,N_7043,N_5973);
and U14278 (N_14278,N_6973,N_9094);
and U14279 (N_14279,N_5887,N_8776);
xnor U14280 (N_14280,N_6031,N_8577);
nand U14281 (N_14281,N_5917,N_6496);
nor U14282 (N_14282,N_8878,N_6483);
nand U14283 (N_14283,N_7990,N_7156);
nand U14284 (N_14284,N_8412,N_6997);
and U14285 (N_14285,N_5576,N_5707);
xnor U14286 (N_14286,N_5123,N_5971);
and U14287 (N_14287,N_6981,N_5782);
or U14288 (N_14288,N_6967,N_6859);
and U14289 (N_14289,N_9721,N_9790);
nor U14290 (N_14290,N_8452,N_5560);
xor U14291 (N_14291,N_8039,N_9950);
or U14292 (N_14292,N_5669,N_6456);
nand U14293 (N_14293,N_5551,N_9824);
nor U14294 (N_14294,N_8295,N_5148);
or U14295 (N_14295,N_5530,N_7091);
and U14296 (N_14296,N_5640,N_6944);
and U14297 (N_14297,N_8287,N_6421);
xnor U14298 (N_14298,N_9631,N_5399);
nand U14299 (N_14299,N_5723,N_8135);
xnor U14300 (N_14300,N_8050,N_6294);
or U14301 (N_14301,N_7074,N_5642);
xnor U14302 (N_14302,N_8534,N_6916);
xnor U14303 (N_14303,N_9232,N_5091);
nand U14304 (N_14304,N_6928,N_6181);
and U14305 (N_14305,N_6920,N_8249);
and U14306 (N_14306,N_8970,N_6815);
nor U14307 (N_14307,N_8367,N_9494);
or U14308 (N_14308,N_8118,N_7695);
nand U14309 (N_14309,N_5012,N_7347);
nand U14310 (N_14310,N_6353,N_7666);
nor U14311 (N_14311,N_5557,N_5721);
and U14312 (N_14312,N_8568,N_8227);
xor U14313 (N_14313,N_8303,N_8507);
and U14314 (N_14314,N_8891,N_7725);
nand U14315 (N_14315,N_8695,N_7190);
or U14316 (N_14316,N_7629,N_6411);
xor U14317 (N_14317,N_6064,N_9013);
or U14318 (N_14318,N_7365,N_9151);
and U14319 (N_14319,N_6011,N_8570);
nand U14320 (N_14320,N_7979,N_9700);
nor U14321 (N_14321,N_8473,N_8761);
xnor U14322 (N_14322,N_5142,N_9256);
xor U14323 (N_14323,N_7186,N_7112);
or U14324 (N_14324,N_5473,N_7421);
nor U14325 (N_14325,N_8218,N_6722);
nor U14326 (N_14326,N_8161,N_6137);
and U14327 (N_14327,N_8557,N_7077);
nand U14328 (N_14328,N_9721,N_5862);
or U14329 (N_14329,N_9793,N_5088);
and U14330 (N_14330,N_6713,N_9527);
or U14331 (N_14331,N_5717,N_8530);
nand U14332 (N_14332,N_9155,N_5696);
and U14333 (N_14333,N_5218,N_5097);
xnor U14334 (N_14334,N_7342,N_9043);
and U14335 (N_14335,N_5976,N_7874);
xnor U14336 (N_14336,N_7096,N_5690);
or U14337 (N_14337,N_6284,N_8243);
nor U14338 (N_14338,N_9971,N_5111);
nand U14339 (N_14339,N_7563,N_6669);
and U14340 (N_14340,N_9420,N_9198);
or U14341 (N_14341,N_8282,N_9047);
and U14342 (N_14342,N_6433,N_7714);
or U14343 (N_14343,N_5413,N_8744);
nor U14344 (N_14344,N_7515,N_9142);
nand U14345 (N_14345,N_6911,N_6769);
nor U14346 (N_14346,N_9962,N_6907);
nand U14347 (N_14347,N_8153,N_5903);
or U14348 (N_14348,N_5524,N_5281);
and U14349 (N_14349,N_5776,N_6889);
nand U14350 (N_14350,N_8207,N_9586);
and U14351 (N_14351,N_6542,N_5469);
xnor U14352 (N_14352,N_8004,N_6244);
or U14353 (N_14353,N_6079,N_9387);
nor U14354 (N_14354,N_9183,N_8679);
nand U14355 (N_14355,N_5995,N_8814);
and U14356 (N_14356,N_9748,N_7854);
or U14357 (N_14357,N_9322,N_8950);
nand U14358 (N_14358,N_9390,N_9969);
and U14359 (N_14359,N_5810,N_7975);
or U14360 (N_14360,N_7345,N_8465);
nand U14361 (N_14361,N_7715,N_6313);
nor U14362 (N_14362,N_6981,N_6687);
and U14363 (N_14363,N_6845,N_6446);
and U14364 (N_14364,N_6106,N_6122);
and U14365 (N_14365,N_7454,N_7865);
or U14366 (N_14366,N_9614,N_6096);
or U14367 (N_14367,N_6753,N_6914);
or U14368 (N_14368,N_6234,N_5871);
and U14369 (N_14369,N_8700,N_5840);
or U14370 (N_14370,N_9181,N_7637);
and U14371 (N_14371,N_9816,N_6942);
nor U14372 (N_14372,N_7681,N_5208);
nor U14373 (N_14373,N_7944,N_8501);
and U14374 (N_14374,N_9237,N_9896);
xor U14375 (N_14375,N_8899,N_9398);
nor U14376 (N_14376,N_5164,N_6105);
or U14377 (N_14377,N_5331,N_5938);
or U14378 (N_14378,N_8174,N_9456);
xnor U14379 (N_14379,N_9832,N_5415);
and U14380 (N_14380,N_9679,N_6349);
and U14381 (N_14381,N_8973,N_5707);
xor U14382 (N_14382,N_8197,N_5861);
and U14383 (N_14383,N_7105,N_8564);
nand U14384 (N_14384,N_9099,N_7949);
and U14385 (N_14385,N_9881,N_9644);
and U14386 (N_14386,N_9867,N_9948);
nand U14387 (N_14387,N_8529,N_6116);
nor U14388 (N_14388,N_7671,N_9150);
and U14389 (N_14389,N_7772,N_7711);
nor U14390 (N_14390,N_8264,N_7631);
nand U14391 (N_14391,N_8624,N_6662);
or U14392 (N_14392,N_5508,N_5478);
and U14393 (N_14393,N_9035,N_8595);
or U14394 (N_14394,N_6103,N_5194);
and U14395 (N_14395,N_9833,N_7581);
xor U14396 (N_14396,N_8719,N_8842);
nand U14397 (N_14397,N_9695,N_8861);
nor U14398 (N_14398,N_8701,N_8847);
nor U14399 (N_14399,N_5087,N_5646);
xnor U14400 (N_14400,N_8575,N_8110);
or U14401 (N_14401,N_8061,N_5922);
xnor U14402 (N_14402,N_7901,N_8994);
nor U14403 (N_14403,N_9302,N_8810);
and U14404 (N_14404,N_9767,N_9879);
nor U14405 (N_14405,N_6062,N_8545);
and U14406 (N_14406,N_7753,N_7782);
xnor U14407 (N_14407,N_8933,N_6596);
and U14408 (N_14408,N_8455,N_5266);
nor U14409 (N_14409,N_8672,N_9639);
or U14410 (N_14410,N_7853,N_6413);
and U14411 (N_14411,N_6223,N_5067);
xnor U14412 (N_14412,N_7449,N_7325);
xnor U14413 (N_14413,N_6330,N_8669);
xnor U14414 (N_14414,N_5711,N_5119);
nor U14415 (N_14415,N_5386,N_6168);
and U14416 (N_14416,N_5311,N_5797);
and U14417 (N_14417,N_9333,N_9465);
xnor U14418 (N_14418,N_5973,N_8993);
or U14419 (N_14419,N_7564,N_8869);
or U14420 (N_14420,N_7440,N_9691);
xor U14421 (N_14421,N_7922,N_8276);
nand U14422 (N_14422,N_6934,N_5802);
xor U14423 (N_14423,N_7756,N_8031);
and U14424 (N_14424,N_5472,N_6119);
or U14425 (N_14425,N_6022,N_7317);
nand U14426 (N_14426,N_8624,N_9116);
xor U14427 (N_14427,N_6356,N_5907);
nand U14428 (N_14428,N_6203,N_9376);
nand U14429 (N_14429,N_9869,N_8285);
nand U14430 (N_14430,N_8076,N_8786);
xor U14431 (N_14431,N_9515,N_7060);
xor U14432 (N_14432,N_5591,N_7103);
xnor U14433 (N_14433,N_9656,N_6518);
xor U14434 (N_14434,N_7184,N_5393);
nor U14435 (N_14435,N_7580,N_6366);
or U14436 (N_14436,N_5811,N_8745);
nand U14437 (N_14437,N_7208,N_6121);
or U14438 (N_14438,N_6574,N_8222);
nand U14439 (N_14439,N_7410,N_7069);
nor U14440 (N_14440,N_7229,N_9252);
nand U14441 (N_14441,N_6979,N_8651);
nor U14442 (N_14442,N_9226,N_5600);
nor U14443 (N_14443,N_5862,N_9244);
or U14444 (N_14444,N_5572,N_7043);
or U14445 (N_14445,N_7215,N_7304);
nor U14446 (N_14446,N_7916,N_9518);
nand U14447 (N_14447,N_8948,N_6781);
nor U14448 (N_14448,N_9296,N_6721);
and U14449 (N_14449,N_5400,N_6712);
or U14450 (N_14450,N_6195,N_7853);
and U14451 (N_14451,N_8887,N_9513);
nor U14452 (N_14452,N_8644,N_7033);
and U14453 (N_14453,N_5020,N_6492);
nor U14454 (N_14454,N_6563,N_6720);
nand U14455 (N_14455,N_9264,N_9887);
and U14456 (N_14456,N_8804,N_9012);
xor U14457 (N_14457,N_6007,N_6116);
and U14458 (N_14458,N_9753,N_8724);
or U14459 (N_14459,N_6892,N_7398);
and U14460 (N_14460,N_5113,N_7157);
and U14461 (N_14461,N_9700,N_8044);
and U14462 (N_14462,N_8083,N_8521);
nor U14463 (N_14463,N_6924,N_9361);
and U14464 (N_14464,N_7291,N_5424);
and U14465 (N_14465,N_7253,N_5333);
nand U14466 (N_14466,N_7187,N_8844);
nand U14467 (N_14467,N_8035,N_7752);
and U14468 (N_14468,N_7527,N_9666);
and U14469 (N_14469,N_5747,N_6390);
or U14470 (N_14470,N_6074,N_5239);
xnor U14471 (N_14471,N_6112,N_5498);
nand U14472 (N_14472,N_7250,N_9454);
xor U14473 (N_14473,N_6036,N_5887);
or U14474 (N_14474,N_5955,N_5210);
and U14475 (N_14475,N_8278,N_9196);
and U14476 (N_14476,N_6706,N_9941);
xnor U14477 (N_14477,N_6205,N_9349);
nand U14478 (N_14478,N_7893,N_8624);
xnor U14479 (N_14479,N_8185,N_7087);
nor U14480 (N_14480,N_8542,N_8343);
and U14481 (N_14481,N_6307,N_6625);
or U14482 (N_14482,N_8961,N_8037);
nand U14483 (N_14483,N_8385,N_7095);
nor U14484 (N_14484,N_8743,N_5017);
xnor U14485 (N_14485,N_9186,N_9610);
nand U14486 (N_14486,N_8404,N_9286);
nor U14487 (N_14487,N_5063,N_7053);
nor U14488 (N_14488,N_9477,N_9846);
and U14489 (N_14489,N_5787,N_6921);
nor U14490 (N_14490,N_9828,N_6732);
nor U14491 (N_14491,N_9776,N_6378);
nand U14492 (N_14492,N_9459,N_7659);
xnor U14493 (N_14493,N_9237,N_7318);
or U14494 (N_14494,N_5540,N_8631);
or U14495 (N_14495,N_8656,N_7446);
xnor U14496 (N_14496,N_9221,N_7122);
or U14497 (N_14497,N_6978,N_8986);
xor U14498 (N_14498,N_7796,N_5803);
and U14499 (N_14499,N_7493,N_7663);
and U14500 (N_14500,N_7574,N_8270);
nand U14501 (N_14501,N_8973,N_7743);
nand U14502 (N_14502,N_8642,N_6844);
nor U14503 (N_14503,N_8161,N_6786);
and U14504 (N_14504,N_6956,N_5350);
xnor U14505 (N_14505,N_8787,N_8491);
and U14506 (N_14506,N_5398,N_6344);
nor U14507 (N_14507,N_5024,N_7195);
xnor U14508 (N_14508,N_7796,N_7033);
nor U14509 (N_14509,N_8803,N_6931);
or U14510 (N_14510,N_5656,N_7562);
xnor U14511 (N_14511,N_9896,N_7044);
xor U14512 (N_14512,N_7717,N_8483);
nand U14513 (N_14513,N_9091,N_7425);
nand U14514 (N_14514,N_5387,N_7879);
nor U14515 (N_14515,N_7674,N_9942);
xnor U14516 (N_14516,N_7930,N_5483);
nand U14517 (N_14517,N_8261,N_8246);
nor U14518 (N_14518,N_7625,N_5119);
xnor U14519 (N_14519,N_6723,N_6270);
nand U14520 (N_14520,N_5087,N_5011);
xor U14521 (N_14521,N_6905,N_9319);
and U14522 (N_14522,N_9764,N_5790);
or U14523 (N_14523,N_7355,N_5982);
nand U14524 (N_14524,N_9559,N_9288);
xor U14525 (N_14525,N_9813,N_9891);
or U14526 (N_14526,N_8734,N_6553);
nor U14527 (N_14527,N_8950,N_8232);
nand U14528 (N_14528,N_8444,N_5621);
xnor U14529 (N_14529,N_6709,N_8909);
and U14530 (N_14530,N_9109,N_5338);
nor U14531 (N_14531,N_7619,N_6947);
nand U14532 (N_14532,N_9618,N_5341);
xor U14533 (N_14533,N_9149,N_7487);
nor U14534 (N_14534,N_9120,N_7273);
nor U14535 (N_14535,N_9053,N_6091);
and U14536 (N_14536,N_8205,N_5528);
nor U14537 (N_14537,N_5969,N_5096);
nand U14538 (N_14538,N_9863,N_6297);
and U14539 (N_14539,N_5847,N_8517);
or U14540 (N_14540,N_5165,N_6462);
nand U14541 (N_14541,N_7380,N_9015);
or U14542 (N_14542,N_5159,N_9465);
or U14543 (N_14543,N_5203,N_6135);
xnor U14544 (N_14544,N_7848,N_9763);
nand U14545 (N_14545,N_9090,N_5120);
nand U14546 (N_14546,N_8738,N_6461);
nor U14547 (N_14547,N_6573,N_6288);
xor U14548 (N_14548,N_8148,N_7475);
and U14549 (N_14549,N_7011,N_7154);
nor U14550 (N_14550,N_9271,N_7891);
nor U14551 (N_14551,N_6658,N_5401);
or U14552 (N_14552,N_5067,N_5646);
or U14553 (N_14553,N_8308,N_5048);
or U14554 (N_14554,N_7807,N_5883);
and U14555 (N_14555,N_8040,N_8920);
nor U14556 (N_14556,N_9155,N_8343);
xnor U14557 (N_14557,N_8492,N_6763);
nand U14558 (N_14558,N_5293,N_8302);
or U14559 (N_14559,N_6391,N_6204);
nand U14560 (N_14560,N_6253,N_9860);
xor U14561 (N_14561,N_5451,N_5527);
or U14562 (N_14562,N_7394,N_9557);
nor U14563 (N_14563,N_6424,N_7637);
or U14564 (N_14564,N_7688,N_5355);
and U14565 (N_14565,N_9994,N_5429);
nand U14566 (N_14566,N_7420,N_8770);
nor U14567 (N_14567,N_5399,N_6351);
nand U14568 (N_14568,N_5754,N_8742);
nand U14569 (N_14569,N_7195,N_5406);
or U14570 (N_14570,N_7125,N_9159);
xor U14571 (N_14571,N_8778,N_9245);
or U14572 (N_14572,N_8965,N_8870);
xnor U14573 (N_14573,N_5646,N_8708);
nand U14574 (N_14574,N_8268,N_5591);
nor U14575 (N_14575,N_8187,N_6977);
or U14576 (N_14576,N_8107,N_5158);
or U14577 (N_14577,N_9690,N_6512);
and U14578 (N_14578,N_9530,N_6156);
nor U14579 (N_14579,N_8720,N_5032);
xnor U14580 (N_14580,N_7445,N_6503);
and U14581 (N_14581,N_7365,N_6441);
xor U14582 (N_14582,N_8038,N_8234);
nor U14583 (N_14583,N_8332,N_5272);
nor U14584 (N_14584,N_5974,N_9019);
and U14585 (N_14585,N_7824,N_9067);
and U14586 (N_14586,N_7226,N_9464);
or U14587 (N_14587,N_6601,N_8193);
xor U14588 (N_14588,N_9155,N_7404);
nand U14589 (N_14589,N_5007,N_5431);
xor U14590 (N_14590,N_6015,N_6231);
nand U14591 (N_14591,N_9071,N_6552);
xor U14592 (N_14592,N_7666,N_5014);
xor U14593 (N_14593,N_5125,N_8345);
nor U14594 (N_14594,N_5738,N_8960);
xor U14595 (N_14595,N_6234,N_5834);
and U14596 (N_14596,N_6355,N_8985);
or U14597 (N_14597,N_9040,N_7057);
or U14598 (N_14598,N_8904,N_9166);
nand U14599 (N_14599,N_8221,N_6475);
or U14600 (N_14600,N_5012,N_8233);
or U14601 (N_14601,N_6317,N_5633);
nor U14602 (N_14602,N_9760,N_6408);
or U14603 (N_14603,N_5565,N_6372);
xnor U14604 (N_14604,N_6528,N_5868);
or U14605 (N_14605,N_9238,N_6123);
nand U14606 (N_14606,N_8620,N_8228);
or U14607 (N_14607,N_9294,N_9473);
nand U14608 (N_14608,N_5011,N_9549);
or U14609 (N_14609,N_8376,N_8243);
nor U14610 (N_14610,N_5092,N_9376);
nand U14611 (N_14611,N_5722,N_8760);
or U14612 (N_14612,N_5965,N_9439);
nor U14613 (N_14613,N_7513,N_8610);
nand U14614 (N_14614,N_8109,N_9583);
xnor U14615 (N_14615,N_8800,N_6175);
xor U14616 (N_14616,N_9538,N_7058);
nand U14617 (N_14617,N_5650,N_5113);
nand U14618 (N_14618,N_8035,N_8073);
nor U14619 (N_14619,N_8812,N_5804);
and U14620 (N_14620,N_6795,N_8167);
and U14621 (N_14621,N_7244,N_9798);
and U14622 (N_14622,N_8038,N_5815);
nor U14623 (N_14623,N_7159,N_9702);
and U14624 (N_14624,N_6658,N_8260);
xor U14625 (N_14625,N_6463,N_6007);
xnor U14626 (N_14626,N_6004,N_9019);
and U14627 (N_14627,N_8581,N_8702);
nor U14628 (N_14628,N_9969,N_8731);
nor U14629 (N_14629,N_9956,N_5958);
and U14630 (N_14630,N_7187,N_6920);
or U14631 (N_14631,N_9150,N_8298);
and U14632 (N_14632,N_8392,N_7629);
nor U14633 (N_14633,N_9991,N_9434);
nand U14634 (N_14634,N_6617,N_9743);
nor U14635 (N_14635,N_5075,N_9212);
or U14636 (N_14636,N_8976,N_5638);
xor U14637 (N_14637,N_9465,N_8129);
nor U14638 (N_14638,N_9427,N_5292);
xor U14639 (N_14639,N_7954,N_8164);
and U14640 (N_14640,N_9698,N_8967);
xor U14641 (N_14641,N_9096,N_5761);
nor U14642 (N_14642,N_9147,N_6030);
and U14643 (N_14643,N_5470,N_7355);
nand U14644 (N_14644,N_7963,N_9153);
nand U14645 (N_14645,N_8733,N_8355);
xor U14646 (N_14646,N_6659,N_7156);
nand U14647 (N_14647,N_7168,N_9035);
and U14648 (N_14648,N_7788,N_8509);
and U14649 (N_14649,N_7458,N_9247);
nor U14650 (N_14650,N_5620,N_5498);
nor U14651 (N_14651,N_8376,N_6315);
or U14652 (N_14652,N_7840,N_6870);
and U14653 (N_14653,N_8673,N_9380);
nand U14654 (N_14654,N_6406,N_6906);
nand U14655 (N_14655,N_7657,N_5875);
nand U14656 (N_14656,N_9938,N_7590);
or U14657 (N_14657,N_8361,N_9022);
and U14658 (N_14658,N_9883,N_7684);
or U14659 (N_14659,N_9946,N_9603);
and U14660 (N_14660,N_5024,N_9491);
or U14661 (N_14661,N_5576,N_5181);
and U14662 (N_14662,N_9641,N_7131);
and U14663 (N_14663,N_5048,N_6387);
or U14664 (N_14664,N_5705,N_9920);
xnor U14665 (N_14665,N_8568,N_6835);
or U14666 (N_14666,N_7388,N_8050);
nor U14667 (N_14667,N_8429,N_7956);
or U14668 (N_14668,N_8793,N_7031);
nor U14669 (N_14669,N_6561,N_5213);
and U14670 (N_14670,N_6396,N_6292);
and U14671 (N_14671,N_7818,N_5083);
xnor U14672 (N_14672,N_5276,N_6681);
nor U14673 (N_14673,N_5482,N_9284);
xor U14674 (N_14674,N_5401,N_5404);
xnor U14675 (N_14675,N_6185,N_5933);
nand U14676 (N_14676,N_5680,N_5111);
nand U14677 (N_14677,N_6963,N_5261);
nor U14678 (N_14678,N_6891,N_7685);
nor U14679 (N_14679,N_6923,N_6259);
and U14680 (N_14680,N_6073,N_5873);
nor U14681 (N_14681,N_7109,N_6684);
nand U14682 (N_14682,N_5251,N_5778);
nor U14683 (N_14683,N_6442,N_8411);
nand U14684 (N_14684,N_7177,N_8505);
and U14685 (N_14685,N_6908,N_7471);
and U14686 (N_14686,N_8525,N_9447);
and U14687 (N_14687,N_9729,N_6552);
nand U14688 (N_14688,N_6438,N_8903);
nand U14689 (N_14689,N_8964,N_6138);
xnor U14690 (N_14690,N_7201,N_7518);
or U14691 (N_14691,N_8834,N_5995);
and U14692 (N_14692,N_7877,N_8126);
and U14693 (N_14693,N_6519,N_9958);
nand U14694 (N_14694,N_6252,N_7914);
nand U14695 (N_14695,N_5642,N_8085);
and U14696 (N_14696,N_7718,N_7589);
xnor U14697 (N_14697,N_7133,N_7321);
or U14698 (N_14698,N_6674,N_9069);
nand U14699 (N_14699,N_7558,N_9825);
xnor U14700 (N_14700,N_6754,N_6058);
and U14701 (N_14701,N_7172,N_9129);
nor U14702 (N_14702,N_6308,N_6792);
xor U14703 (N_14703,N_6530,N_7687);
nor U14704 (N_14704,N_8486,N_6449);
xnor U14705 (N_14705,N_9993,N_8892);
xnor U14706 (N_14706,N_9658,N_5210);
or U14707 (N_14707,N_7343,N_8614);
nand U14708 (N_14708,N_7261,N_8587);
xnor U14709 (N_14709,N_8981,N_5141);
nor U14710 (N_14710,N_8434,N_7901);
and U14711 (N_14711,N_5147,N_7241);
nand U14712 (N_14712,N_9033,N_7627);
nand U14713 (N_14713,N_5508,N_6817);
or U14714 (N_14714,N_9909,N_9669);
or U14715 (N_14715,N_5232,N_6820);
xnor U14716 (N_14716,N_8372,N_8996);
and U14717 (N_14717,N_5151,N_5279);
xor U14718 (N_14718,N_8027,N_8822);
xnor U14719 (N_14719,N_7297,N_8834);
nand U14720 (N_14720,N_7073,N_5776);
nor U14721 (N_14721,N_5699,N_9483);
or U14722 (N_14722,N_5819,N_5517);
and U14723 (N_14723,N_6038,N_7934);
nor U14724 (N_14724,N_9357,N_8169);
or U14725 (N_14725,N_8212,N_7390);
xor U14726 (N_14726,N_6329,N_8171);
nor U14727 (N_14727,N_6264,N_6427);
xor U14728 (N_14728,N_6766,N_5703);
or U14729 (N_14729,N_7966,N_8719);
nand U14730 (N_14730,N_7690,N_5087);
nor U14731 (N_14731,N_9130,N_7482);
nor U14732 (N_14732,N_7428,N_6661);
xnor U14733 (N_14733,N_5424,N_7157);
nand U14734 (N_14734,N_6831,N_8586);
xnor U14735 (N_14735,N_8280,N_6592);
xor U14736 (N_14736,N_6889,N_5024);
nor U14737 (N_14737,N_6528,N_8860);
xnor U14738 (N_14738,N_9211,N_5806);
nand U14739 (N_14739,N_5950,N_9240);
nor U14740 (N_14740,N_7527,N_8015);
nor U14741 (N_14741,N_8525,N_5067);
nor U14742 (N_14742,N_7118,N_9871);
nor U14743 (N_14743,N_7805,N_5964);
or U14744 (N_14744,N_7867,N_9528);
or U14745 (N_14745,N_9793,N_8625);
and U14746 (N_14746,N_5286,N_8574);
nand U14747 (N_14747,N_7412,N_6159);
xor U14748 (N_14748,N_9943,N_5429);
nor U14749 (N_14749,N_5118,N_5309);
and U14750 (N_14750,N_5378,N_6573);
nand U14751 (N_14751,N_8359,N_6114);
nor U14752 (N_14752,N_7148,N_8472);
xnor U14753 (N_14753,N_5029,N_5981);
or U14754 (N_14754,N_7272,N_7928);
nor U14755 (N_14755,N_6708,N_9502);
and U14756 (N_14756,N_8348,N_5780);
nor U14757 (N_14757,N_8144,N_8280);
nor U14758 (N_14758,N_6482,N_6925);
or U14759 (N_14759,N_8938,N_8099);
or U14760 (N_14760,N_9386,N_7572);
or U14761 (N_14761,N_8131,N_7732);
and U14762 (N_14762,N_6327,N_9253);
nand U14763 (N_14763,N_7558,N_7660);
xnor U14764 (N_14764,N_5819,N_6483);
nand U14765 (N_14765,N_9449,N_8597);
or U14766 (N_14766,N_6837,N_9254);
nor U14767 (N_14767,N_8679,N_8101);
xor U14768 (N_14768,N_8214,N_7708);
or U14769 (N_14769,N_6005,N_5175);
nor U14770 (N_14770,N_7449,N_8501);
or U14771 (N_14771,N_7502,N_6048);
or U14772 (N_14772,N_9312,N_5537);
and U14773 (N_14773,N_8559,N_5188);
nand U14774 (N_14774,N_6271,N_9183);
xor U14775 (N_14775,N_8275,N_9660);
xnor U14776 (N_14776,N_9515,N_6436);
nand U14777 (N_14777,N_7548,N_7373);
or U14778 (N_14778,N_5837,N_5005);
xor U14779 (N_14779,N_6747,N_5415);
nand U14780 (N_14780,N_8872,N_5297);
xor U14781 (N_14781,N_9145,N_9237);
and U14782 (N_14782,N_5245,N_9637);
and U14783 (N_14783,N_7687,N_6856);
or U14784 (N_14784,N_9735,N_8539);
xnor U14785 (N_14785,N_7377,N_5150);
nor U14786 (N_14786,N_6050,N_5491);
nor U14787 (N_14787,N_7500,N_9579);
xor U14788 (N_14788,N_5851,N_8837);
nor U14789 (N_14789,N_9190,N_6204);
nor U14790 (N_14790,N_7445,N_7557);
nor U14791 (N_14791,N_6826,N_6327);
and U14792 (N_14792,N_8145,N_6080);
or U14793 (N_14793,N_5307,N_7475);
xor U14794 (N_14794,N_5170,N_9311);
and U14795 (N_14795,N_7414,N_7740);
or U14796 (N_14796,N_6331,N_7761);
xor U14797 (N_14797,N_6242,N_9494);
nand U14798 (N_14798,N_9885,N_7910);
and U14799 (N_14799,N_5452,N_8586);
nand U14800 (N_14800,N_5461,N_5007);
or U14801 (N_14801,N_8418,N_7283);
and U14802 (N_14802,N_8796,N_6449);
and U14803 (N_14803,N_5332,N_8136);
nor U14804 (N_14804,N_7232,N_9876);
or U14805 (N_14805,N_7689,N_6065);
nor U14806 (N_14806,N_9960,N_7537);
or U14807 (N_14807,N_7857,N_9638);
and U14808 (N_14808,N_6926,N_8923);
or U14809 (N_14809,N_5907,N_6615);
or U14810 (N_14810,N_6702,N_9746);
xnor U14811 (N_14811,N_8847,N_7205);
nor U14812 (N_14812,N_8880,N_9284);
nand U14813 (N_14813,N_8204,N_8690);
xnor U14814 (N_14814,N_8505,N_6825);
xnor U14815 (N_14815,N_7078,N_9057);
nor U14816 (N_14816,N_7398,N_7466);
nand U14817 (N_14817,N_6362,N_8736);
and U14818 (N_14818,N_6460,N_9207);
nand U14819 (N_14819,N_7051,N_6701);
xor U14820 (N_14820,N_7084,N_9073);
or U14821 (N_14821,N_8423,N_7835);
xor U14822 (N_14822,N_5060,N_7794);
or U14823 (N_14823,N_9819,N_6949);
xor U14824 (N_14824,N_6146,N_6441);
or U14825 (N_14825,N_8669,N_5569);
nand U14826 (N_14826,N_5225,N_9929);
nand U14827 (N_14827,N_5301,N_6871);
and U14828 (N_14828,N_6801,N_6480);
and U14829 (N_14829,N_7290,N_8991);
nand U14830 (N_14830,N_6854,N_6847);
nand U14831 (N_14831,N_5500,N_7438);
xor U14832 (N_14832,N_8844,N_8181);
nor U14833 (N_14833,N_6407,N_7152);
or U14834 (N_14834,N_8581,N_6088);
xnor U14835 (N_14835,N_7061,N_5453);
nor U14836 (N_14836,N_5437,N_5923);
nor U14837 (N_14837,N_9022,N_7236);
nor U14838 (N_14838,N_8466,N_8114);
nand U14839 (N_14839,N_7616,N_7208);
or U14840 (N_14840,N_5019,N_6823);
and U14841 (N_14841,N_6289,N_5080);
xnor U14842 (N_14842,N_7312,N_8654);
xor U14843 (N_14843,N_6940,N_9627);
and U14844 (N_14844,N_7093,N_8377);
or U14845 (N_14845,N_5658,N_6144);
or U14846 (N_14846,N_5761,N_9724);
nand U14847 (N_14847,N_5774,N_6784);
nor U14848 (N_14848,N_6345,N_6825);
nor U14849 (N_14849,N_8720,N_7013);
or U14850 (N_14850,N_9193,N_5002);
nand U14851 (N_14851,N_9143,N_6466);
and U14852 (N_14852,N_8431,N_5934);
or U14853 (N_14853,N_5517,N_6441);
and U14854 (N_14854,N_8739,N_9999);
nor U14855 (N_14855,N_8698,N_9465);
and U14856 (N_14856,N_5923,N_6491);
xor U14857 (N_14857,N_6165,N_5488);
xnor U14858 (N_14858,N_8579,N_8997);
nand U14859 (N_14859,N_8074,N_7229);
or U14860 (N_14860,N_5335,N_7377);
nand U14861 (N_14861,N_6331,N_8951);
or U14862 (N_14862,N_5006,N_9143);
and U14863 (N_14863,N_5148,N_5029);
nand U14864 (N_14864,N_9820,N_5746);
nor U14865 (N_14865,N_5793,N_6759);
xnor U14866 (N_14866,N_8591,N_8212);
and U14867 (N_14867,N_8782,N_6890);
nor U14868 (N_14868,N_9100,N_6721);
nor U14869 (N_14869,N_8691,N_9121);
xor U14870 (N_14870,N_5497,N_9267);
xnor U14871 (N_14871,N_5878,N_8807);
or U14872 (N_14872,N_8556,N_9463);
or U14873 (N_14873,N_7708,N_6346);
and U14874 (N_14874,N_7237,N_7488);
and U14875 (N_14875,N_6081,N_7256);
or U14876 (N_14876,N_7885,N_9625);
or U14877 (N_14877,N_9545,N_7832);
or U14878 (N_14878,N_9313,N_5198);
or U14879 (N_14879,N_7964,N_9193);
nor U14880 (N_14880,N_8740,N_5812);
and U14881 (N_14881,N_9324,N_5820);
or U14882 (N_14882,N_6947,N_5348);
xor U14883 (N_14883,N_8082,N_9054);
xnor U14884 (N_14884,N_6054,N_9014);
nand U14885 (N_14885,N_8012,N_7601);
or U14886 (N_14886,N_8435,N_7383);
nand U14887 (N_14887,N_7516,N_5979);
or U14888 (N_14888,N_9846,N_9195);
nor U14889 (N_14889,N_6920,N_7927);
and U14890 (N_14890,N_6969,N_7112);
xor U14891 (N_14891,N_9743,N_8686);
nor U14892 (N_14892,N_5472,N_8351);
or U14893 (N_14893,N_7514,N_8197);
nand U14894 (N_14894,N_8178,N_9693);
nand U14895 (N_14895,N_6011,N_6190);
nor U14896 (N_14896,N_9735,N_8962);
nand U14897 (N_14897,N_8782,N_7055);
nand U14898 (N_14898,N_6336,N_5165);
and U14899 (N_14899,N_5817,N_6756);
or U14900 (N_14900,N_5631,N_6998);
and U14901 (N_14901,N_5139,N_8651);
nand U14902 (N_14902,N_9551,N_9366);
or U14903 (N_14903,N_9470,N_9383);
or U14904 (N_14904,N_6954,N_9717);
and U14905 (N_14905,N_6172,N_6340);
nand U14906 (N_14906,N_9650,N_6667);
nor U14907 (N_14907,N_6112,N_7047);
nor U14908 (N_14908,N_5929,N_9434);
nor U14909 (N_14909,N_7308,N_9036);
nand U14910 (N_14910,N_9773,N_8691);
xor U14911 (N_14911,N_9461,N_7155);
nand U14912 (N_14912,N_9228,N_8107);
nor U14913 (N_14913,N_6089,N_9905);
nor U14914 (N_14914,N_7845,N_9307);
nor U14915 (N_14915,N_8038,N_9260);
xnor U14916 (N_14916,N_5441,N_7240);
nand U14917 (N_14917,N_7857,N_5216);
nand U14918 (N_14918,N_7208,N_7369);
nand U14919 (N_14919,N_9645,N_9233);
or U14920 (N_14920,N_9556,N_6584);
nor U14921 (N_14921,N_9724,N_9068);
nand U14922 (N_14922,N_5296,N_6502);
xor U14923 (N_14923,N_5940,N_7620);
and U14924 (N_14924,N_7826,N_9716);
and U14925 (N_14925,N_7705,N_6717);
nor U14926 (N_14926,N_9721,N_8224);
nor U14927 (N_14927,N_5747,N_6185);
nor U14928 (N_14928,N_5633,N_5215);
nor U14929 (N_14929,N_5266,N_5968);
nor U14930 (N_14930,N_7445,N_9146);
and U14931 (N_14931,N_5626,N_6837);
nor U14932 (N_14932,N_8448,N_9469);
and U14933 (N_14933,N_5637,N_7208);
and U14934 (N_14934,N_7400,N_6566);
xor U14935 (N_14935,N_5019,N_5620);
or U14936 (N_14936,N_7977,N_6407);
nand U14937 (N_14937,N_9167,N_8363);
nand U14938 (N_14938,N_6344,N_6551);
nand U14939 (N_14939,N_5807,N_6413);
nor U14940 (N_14940,N_7970,N_7506);
and U14941 (N_14941,N_6625,N_9755);
and U14942 (N_14942,N_8238,N_8701);
nand U14943 (N_14943,N_9744,N_7883);
nor U14944 (N_14944,N_6269,N_8755);
nand U14945 (N_14945,N_8229,N_6934);
xnor U14946 (N_14946,N_8508,N_6140);
xor U14947 (N_14947,N_8889,N_9805);
and U14948 (N_14948,N_6646,N_7679);
nand U14949 (N_14949,N_7480,N_6033);
and U14950 (N_14950,N_6682,N_8587);
and U14951 (N_14951,N_9574,N_9971);
xor U14952 (N_14952,N_9568,N_6615);
or U14953 (N_14953,N_5526,N_5836);
nand U14954 (N_14954,N_7828,N_6459);
xor U14955 (N_14955,N_9419,N_9600);
or U14956 (N_14956,N_5839,N_5854);
or U14957 (N_14957,N_8415,N_5222);
or U14958 (N_14958,N_8569,N_9823);
nand U14959 (N_14959,N_9643,N_6876);
nand U14960 (N_14960,N_8048,N_8913);
nor U14961 (N_14961,N_8140,N_8103);
xnor U14962 (N_14962,N_7288,N_8833);
nand U14963 (N_14963,N_8469,N_9165);
xnor U14964 (N_14964,N_9719,N_6270);
xnor U14965 (N_14965,N_6061,N_8500);
nor U14966 (N_14966,N_8086,N_5398);
xnor U14967 (N_14967,N_7345,N_5724);
nand U14968 (N_14968,N_7697,N_6450);
and U14969 (N_14969,N_7217,N_8480);
and U14970 (N_14970,N_7304,N_9396);
nand U14971 (N_14971,N_8600,N_5531);
nand U14972 (N_14972,N_6412,N_9608);
or U14973 (N_14973,N_8891,N_5641);
xnor U14974 (N_14974,N_9467,N_5814);
nand U14975 (N_14975,N_6966,N_7052);
and U14976 (N_14976,N_5848,N_6835);
and U14977 (N_14977,N_5233,N_7323);
nor U14978 (N_14978,N_6878,N_9266);
nor U14979 (N_14979,N_9669,N_7527);
nand U14980 (N_14980,N_6244,N_7844);
nor U14981 (N_14981,N_5045,N_9783);
and U14982 (N_14982,N_6577,N_5310);
nand U14983 (N_14983,N_9193,N_8816);
or U14984 (N_14984,N_5020,N_9266);
nor U14985 (N_14985,N_6442,N_7700);
xnor U14986 (N_14986,N_5500,N_7977);
and U14987 (N_14987,N_8774,N_8028);
nand U14988 (N_14988,N_9226,N_6988);
nand U14989 (N_14989,N_9012,N_5605);
and U14990 (N_14990,N_8835,N_9353);
or U14991 (N_14991,N_7007,N_7757);
nand U14992 (N_14992,N_7607,N_6170);
and U14993 (N_14993,N_5045,N_7639);
or U14994 (N_14994,N_7196,N_6521);
and U14995 (N_14995,N_5714,N_9293);
nor U14996 (N_14996,N_7489,N_8286);
or U14997 (N_14997,N_6736,N_6532);
xor U14998 (N_14998,N_7842,N_9917);
xor U14999 (N_14999,N_7728,N_8795);
xnor U15000 (N_15000,N_13442,N_12277);
nor U15001 (N_15001,N_12755,N_10653);
nand U15002 (N_15002,N_10583,N_11091);
and U15003 (N_15003,N_14255,N_14437);
or U15004 (N_15004,N_10499,N_14576);
nand U15005 (N_15005,N_13959,N_12700);
or U15006 (N_15006,N_13133,N_13154);
and U15007 (N_15007,N_10909,N_14948);
and U15008 (N_15008,N_10315,N_13576);
nor U15009 (N_15009,N_14814,N_11374);
or U15010 (N_15010,N_11808,N_13951);
xnor U15011 (N_15011,N_14248,N_12563);
and U15012 (N_15012,N_11783,N_10688);
nand U15013 (N_15013,N_12168,N_10343);
nor U15014 (N_15014,N_13157,N_14602);
or U15015 (N_15015,N_14568,N_14736);
and U15016 (N_15016,N_10391,N_11725);
and U15017 (N_15017,N_10427,N_14941);
xor U15018 (N_15018,N_14101,N_13135);
nand U15019 (N_15019,N_10994,N_12011);
nor U15020 (N_15020,N_14351,N_12558);
or U15021 (N_15021,N_14543,N_14624);
xor U15022 (N_15022,N_11813,N_13118);
and U15023 (N_15023,N_12679,N_12726);
nor U15024 (N_15024,N_12969,N_12974);
nand U15025 (N_15025,N_14368,N_13469);
or U15026 (N_15026,N_10516,N_12286);
and U15027 (N_15027,N_11582,N_14785);
nand U15028 (N_15028,N_11310,N_10323);
nand U15029 (N_15029,N_11316,N_11908);
xnor U15030 (N_15030,N_10594,N_10749);
or U15031 (N_15031,N_13144,N_12920);
nand U15032 (N_15032,N_12473,N_14607);
nor U15033 (N_15033,N_14170,N_14415);
nand U15034 (N_15034,N_12963,N_12228);
nor U15035 (N_15035,N_12701,N_11919);
and U15036 (N_15036,N_14837,N_13239);
or U15037 (N_15037,N_13603,N_12347);
nand U15038 (N_15038,N_14540,N_12371);
nor U15039 (N_15039,N_10924,N_11361);
and U15040 (N_15040,N_13030,N_12926);
xnor U15041 (N_15041,N_11731,N_14420);
and U15042 (N_15042,N_12155,N_13685);
nand U15043 (N_15043,N_14601,N_13493);
nor U15044 (N_15044,N_10109,N_14181);
nor U15045 (N_15045,N_13669,N_13424);
nor U15046 (N_15046,N_11454,N_13209);
and U15047 (N_15047,N_13005,N_12145);
and U15048 (N_15048,N_14995,N_10941);
nand U15049 (N_15049,N_13158,N_14413);
and U15050 (N_15050,N_13969,N_13599);
or U15051 (N_15051,N_10958,N_11327);
or U15052 (N_15052,N_11460,N_11542);
xnor U15053 (N_15053,N_12122,N_12084);
nand U15054 (N_15054,N_10366,N_14986);
and U15055 (N_15055,N_13379,N_10769);
or U15056 (N_15056,N_12330,N_11094);
nor U15057 (N_15057,N_12635,N_11786);
and U15058 (N_15058,N_11475,N_10944);
and U15059 (N_15059,N_13869,N_12045);
and U15060 (N_15060,N_14066,N_14581);
nor U15061 (N_15061,N_14093,N_10827);
or U15062 (N_15062,N_10189,N_11947);
nor U15063 (N_15063,N_10683,N_13280);
nor U15064 (N_15064,N_14769,N_13872);
and U15065 (N_15065,N_13911,N_11569);
nand U15066 (N_15066,N_12464,N_12801);
xor U15067 (N_15067,N_10218,N_11009);
nand U15068 (N_15068,N_14214,N_13713);
and U15069 (N_15069,N_12375,N_12170);
and U15070 (N_15070,N_12631,N_10470);
or U15071 (N_15071,N_11155,N_12249);
nor U15072 (N_15072,N_12208,N_12587);
nor U15073 (N_15073,N_11780,N_11660);
xor U15074 (N_15074,N_13568,N_14606);
or U15075 (N_15075,N_12067,N_12958);
or U15076 (N_15076,N_14094,N_13261);
nand U15077 (N_15077,N_11029,N_11358);
xor U15078 (N_15078,N_12555,N_13043);
nand U15079 (N_15079,N_14155,N_14844);
nor U15080 (N_15080,N_14777,N_10217);
or U15081 (N_15081,N_10585,N_10076);
nand U15082 (N_15082,N_10817,N_11942);
xnor U15083 (N_15083,N_11283,N_12935);
nand U15084 (N_15084,N_10955,N_10643);
nand U15085 (N_15085,N_14538,N_14697);
or U15086 (N_15086,N_11382,N_11722);
and U15087 (N_15087,N_13232,N_14300);
nand U15088 (N_15088,N_14726,N_10182);
xor U15089 (N_15089,N_13907,N_13765);
nor U15090 (N_15090,N_14104,N_13919);
and U15091 (N_15091,N_14201,N_10490);
and U15092 (N_15092,N_14627,N_11240);
and U15093 (N_15093,N_11812,N_14085);
nand U15094 (N_15094,N_11644,N_11761);
or U15095 (N_15095,N_13958,N_10649);
nand U15096 (N_15096,N_11863,N_12000);
xnor U15097 (N_15097,N_10259,N_14106);
and U15098 (N_15098,N_13640,N_14553);
xnor U15099 (N_15099,N_14482,N_10146);
nand U15100 (N_15100,N_11206,N_14667);
xnor U15101 (N_15101,N_10111,N_12560);
nor U15102 (N_15102,N_11377,N_13647);
nand U15103 (N_15103,N_13878,N_14889);
nand U15104 (N_15104,N_12303,N_13884);
and U15105 (N_15105,N_10050,N_14779);
xor U15106 (N_15106,N_14706,N_11690);
xor U15107 (N_15107,N_12811,N_11898);
nand U15108 (N_15108,N_12344,N_11597);
or U15109 (N_15109,N_11529,N_14565);
and U15110 (N_15110,N_14324,N_12281);
or U15111 (N_15111,N_11719,N_13539);
or U15112 (N_15112,N_11152,N_11504);
nand U15113 (N_15113,N_12254,N_13826);
and U15114 (N_15114,N_13026,N_10153);
nor U15115 (N_15115,N_13590,N_11464);
nor U15116 (N_15116,N_11553,N_11929);
or U15117 (N_15117,N_13031,N_10498);
or U15118 (N_15118,N_11395,N_11732);
nor U15119 (N_15119,N_13429,N_13347);
nor U15120 (N_15120,N_14906,N_14648);
xnor U15121 (N_15121,N_14856,N_12112);
nor U15122 (N_15122,N_13695,N_14866);
nand U15123 (N_15123,N_12317,N_14940);
and U15124 (N_15124,N_14829,N_14491);
nor U15125 (N_15125,N_14037,N_14325);
nand U15126 (N_15126,N_13012,N_10560);
nand U15127 (N_15127,N_14847,N_10266);
nor U15128 (N_15128,N_13794,N_12175);
xnor U15129 (N_15129,N_11595,N_10602);
or U15130 (N_15130,N_12754,N_14994);
xnor U15131 (N_15131,N_14111,N_10588);
nand U15132 (N_15132,N_14359,N_13314);
and U15133 (N_15133,N_13771,N_12841);
or U15134 (N_15134,N_12648,N_13824);
nand U15135 (N_15135,N_11443,N_12676);
xor U15136 (N_15136,N_10098,N_14382);
xor U15137 (N_15137,N_11585,N_11090);
nand U15138 (N_15138,N_14291,N_14926);
or U15139 (N_15139,N_13077,N_11445);
or U15140 (N_15140,N_12188,N_14310);
nor U15141 (N_15141,N_12750,N_10996);
and U15142 (N_15142,N_12906,N_10440);
nand U15143 (N_15143,N_10547,N_13104);
and U15144 (N_15144,N_13271,N_12026);
or U15145 (N_15145,N_10879,N_12260);
nor U15146 (N_15146,N_13777,N_11050);
and U15147 (N_15147,N_11389,N_10397);
xnor U15148 (N_15148,N_13392,N_12193);
xnor U15149 (N_15149,N_13793,N_10365);
and U15150 (N_15150,N_12034,N_11872);
nand U15151 (N_15151,N_13578,N_10057);
nor U15152 (N_15152,N_10243,N_11698);
nor U15153 (N_15153,N_10957,N_11753);
xor U15154 (N_15154,N_12753,N_13701);
nor U15155 (N_15155,N_11736,N_13384);
nand U15156 (N_15156,N_10745,N_12605);
or U15157 (N_15157,N_11794,N_12348);
nand U15158 (N_15158,N_13899,N_10822);
or U15159 (N_15159,N_12320,N_11914);
and U15160 (N_15160,N_10581,N_13002);
nor U15161 (N_15161,N_14566,N_14100);
nand U15162 (N_15162,N_14259,N_14921);
xnor U15163 (N_15163,N_13003,N_13054);
and U15164 (N_15164,N_11613,N_10389);
xnor U15165 (N_15165,N_11498,N_10080);
or U15166 (N_15166,N_11227,N_14409);
nor U15167 (N_15167,N_11833,N_12394);
xor U15168 (N_15168,N_12198,N_12730);
xor U15169 (N_15169,N_11079,N_10515);
nor U15170 (N_15170,N_10424,N_12670);
nor U15171 (N_15171,N_13885,N_10874);
nor U15172 (N_15172,N_10782,N_14452);
nor U15173 (N_15173,N_10043,N_12486);
nand U15174 (N_15174,N_13452,N_10068);
nor U15175 (N_15175,N_14250,N_12722);
or U15176 (N_15176,N_10964,N_14298);
or U15177 (N_15177,N_12781,N_12436);
xor U15178 (N_15178,N_10796,N_11583);
nand U15179 (N_15179,N_14812,N_14805);
nand U15180 (N_15180,N_14901,N_12385);
nand U15181 (N_15181,N_14247,N_11737);
and U15182 (N_15182,N_12247,N_14447);
nor U15183 (N_15183,N_10691,N_13119);
nand U15184 (N_15184,N_12036,N_14603);
xnor U15185 (N_15185,N_12187,N_12955);
nor U15186 (N_15186,N_11624,N_14330);
nor U15187 (N_15187,N_12884,N_12176);
and U15188 (N_15188,N_14421,N_12567);
xnor U15189 (N_15189,N_13788,N_11654);
nor U15190 (N_15190,N_10381,N_10219);
nand U15191 (N_15191,N_12923,N_11564);
and U15192 (N_15192,N_14362,N_11894);
nand U15193 (N_15193,N_11512,N_14992);
nand U15194 (N_15194,N_13141,N_12691);
or U15195 (N_15195,N_10985,N_13830);
nor U15196 (N_15196,N_11941,N_10661);
or U15197 (N_15197,N_11436,N_12651);
or U15198 (N_15198,N_11008,N_11384);
xnor U15199 (N_15199,N_10064,N_11423);
and U15200 (N_15200,N_13421,N_13061);
nand U15201 (N_15201,N_10304,N_14279);
or U15202 (N_15202,N_11940,N_11349);
nor U15203 (N_15203,N_11554,N_13858);
nor U15204 (N_15204,N_11406,N_11478);
and U15205 (N_15205,N_11267,N_13883);
nand U15206 (N_15206,N_12874,N_10654);
or U15207 (N_15207,N_10695,N_14830);
nor U15208 (N_15208,N_12017,N_14384);
xnor U15209 (N_15209,N_10067,N_11393);
or U15210 (N_15210,N_13938,N_12132);
xor U15211 (N_15211,N_10980,N_12196);
xnor U15212 (N_15212,N_10942,N_14001);
nor U15213 (N_15213,N_13863,N_11902);
nor U15214 (N_15214,N_13089,N_10419);
nand U15215 (N_15215,N_10326,N_13370);
nor U15216 (N_15216,N_11196,N_11258);
xor U15217 (N_15217,N_13170,N_12009);
nand U15218 (N_15218,N_14458,N_12305);
xnor U15219 (N_15219,N_13246,N_14154);
xnor U15220 (N_15220,N_13671,N_13386);
or U15221 (N_15221,N_11648,N_14680);
or U15222 (N_15222,N_10712,N_14700);
or U15223 (N_15223,N_12046,N_12798);
nand U15224 (N_15224,N_11727,N_12250);
and U15225 (N_15225,N_11183,N_13966);
nor U15226 (N_15226,N_12027,N_14717);
nand U15227 (N_15227,N_10267,N_14551);
or U15228 (N_15228,N_14761,N_14164);
and U15229 (N_15229,N_12620,N_13484);
and U15230 (N_15230,N_13902,N_14753);
nand U15231 (N_15231,N_11237,N_10220);
and U15232 (N_15232,N_12994,N_14897);
or U15233 (N_15233,N_11869,N_13790);
and U15234 (N_15234,N_11999,N_12513);
nand U15235 (N_15235,N_10681,N_11122);
xnor U15236 (N_15236,N_14723,N_12349);
nor U15237 (N_15237,N_12352,N_14006);
nand U15238 (N_15238,N_11667,N_12267);
and U15239 (N_15239,N_14712,N_12446);
xnor U15240 (N_15240,N_11527,N_12268);
nand U15241 (N_15241,N_12904,N_12695);
and U15242 (N_15242,N_10034,N_14072);
nand U15243 (N_15243,N_11659,N_10033);
nand U15244 (N_15244,N_12483,N_11205);
nor U15245 (N_15245,N_13307,N_11486);
or U15246 (N_15246,N_10270,N_11016);
nand U15247 (N_15247,N_12339,N_12769);
xnor U15248 (N_15248,N_10108,N_14744);
xnor U15249 (N_15249,N_10203,N_12202);
nor U15250 (N_15250,N_11822,N_10009);
or U15251 (N_15251,N_14560,N_11433);
and U15252 (N_15252,N_13874,N_12076);
or U15253 (N_15253,N_14931,N_12578);
xnor U15254 (N_15254,N_10761,N_13728);
xor U15255 (N_15255,N_13663,N_10598);
nand U15256 (N_15256,N_11980,N_10377);
or U15257 (N_15257,N_10977,N_13029);
nand U15258 (N_15258,N_12624,N_14886);
nor U15259 (N_15259,N_13876,N_10718);
nand U15260 (N_15260,N_14092,N_12592);
xnor U15261 (N_15261,N_14227,N_11077);
and U15262 (N_15262,N_10508,N_13335);
and U15263 (N_15263,N_13717,N_14786);
or U15264 (N_15264,N_10300,N_11288);
nand U15265 (N_15265,N_12859,N_14582);
xnor U15266 (N_15266,N_14719,N_10122);
and U15267 (N_15267,N_10013,N_14463);
or U15268 (N_15268,N_12448,N_13460);
nand U15269 (N_15269,N_11154,N_12181);
or U15270 (N_15270,N_14150,N_14879);
and U15271 (N_15271,N_14394,N_14268);
nand U15272 (N_15272,N_10903,N_14890);
and U15273 (N_15273,N_12912,N_11345);
nor U15274 (N_15274,N_11663,N_11805);
xnor U15275 (N_15275,N_11533,N_10071);
or U15276 (N_15276,N_12301,N_14398);
or U15277 (N_15277,N_14393,N_11230);
nor U15278 (N_15278,N_14859,N_13120);
xor U15279 (N_15279,N_13477,N_11972);
xor U15280 (N_15280,N_14058,N_12746);
nand U15281 (N_15281,N_10674,N_14999);
nor U15282 (N_15282,N_11166,N_11388);
or U15283 (N_15283,N_14872,N_11601);
nand U15284 (N_15284,N_14580,N_12715);
nor U15285 (N_15285,N_14915,N_13354);
and U15286 (N_15286,N_10472,N_13709);
and U15287 (N_15287,N_13451,N_10951);
nor U15288 (N_15288,N_13742,N_11189);
xor U15289 (N_15289,N_14764,N_14173);
xor U15290 (N_15290,N_11193,N_10321);
nor U15291 (N_15291,N_13572,N_14524);
and U15292 (N_15292,N_10505,N_14533);
or U15293 (N_15293,N_11591,N_11562);
nor U15294 (N_15294,N_14056,N_11238);
and U15295 (N_15295,N_13650,N_10757);
and U15296 (N_15296,N_14913,N_12510);
and U15297 (N_15297,N_12931,N_13795);
nor U15298 (N_15298,N_14817,N_12365);
and U15299 (N_15299,N_10734,N_12291);
or U15300 (N_15300,N_11068,N_10597);
nor U15301 (N_15301,N_11211,N_11359);
xor U15302 (N_15302,N_12805,N_10274);
and U15303 (N_15303,N_13300,N_13256);
or U15304 (N_15304,N_12094,N_14287);
nor U15305 (N_15305,N_10252,N_13333);
and U15306 (N_15306,N_11015,N_12119);
nand U15307 (N_15307,N_13413,N_13616);
nor U15308 (N_15308,N_13143,N_12870);
and U15309 (N_15309,N_10636,N_11774);
xnor U15310 (N_15310,N_11130,N_14123);
nand U15311 (N_15311,N_10194,N_13823);
or U15312 (N_15312,N_12516,N_14677);
and U15313 (N_15313,N_11847,N_13110);
or U15314 (N_15314,N_13506,N_12013);
and U15315 (N_15315,N_11579,N_11386);
nor U15316 (N_15316,N_13562,N_12653);
nand U15317 (N_15317,N_10156,N_13900);
nand U15318 (N_15318,N_10821,N_12269);
nor U15319 (N_15319,N_13918,N_13913);
nor U15320 (N_15320,N_13664,N_13566);
nor U15321 (N_15321,N_13980,N_13136);
and U15322 (N_15322,N_12321,N_13199);
or U15323 (N_15323,N_10595,N_14755);
and U15324 (N_15324,N_13147,N_13646);
or U15325 (N_15325,N_14609,N_11816);
nor U15326 (N_15326,N_12962,N_14787);
nor U15327 (N_15327,N_12490,N_14230);
xnor U15328 (N_15328,N_12495,N_10434);
nand U15329 (N_15329,N_11242,N_12388);
and U15330 (N_15330,N_11629,N_10387);
nor U15331 (N_15331,N_11045,N_14682);
and U15332 (N_15332,N_14171,N_14065);
nor U15333 (N_15333,N_13838,N_12530);
or U15334 (N_15334,N_12766,N_10298);
nor U15335 (N_15335,N_13142,N_13584);
xnor U15336 (N_15336,N_13503,N_14574);
nand U15337 (N_15337,N_14443,N_10268);
and U15338 (N_15338,N_13797,N_10234);
or U15339 (N_15339,N_13871,N_12785);
nor U15340 (N_15340,N_11372,N_10934);
and U15341 (N_15341,N_13567,N_12395);
nand U15342 (N_15342,N_14966,N_11437);
xnor U15343 (N_15343,N_14741,N_13614);
and U15344 (N_15344,N_11936,N_10342);
nor U15345 (N_15345,N_10041,N_13955);
xnor U15346 (N_15346,N_12989,N_10264);
or U15347 (N_15347,N_13049,N_10392);
nor U15348 (N_15348,N_11730,N_14046);
and U15349 (N_15349,N_10592,N_12796);
or U15350 (N_15350,N_13294,N_13723);
xnor U15351 (N_15351,N_12271,N_11302);
nand U15352 (N_15352,N_13815,N_14508);
or U15353 (N_15353,N_13456,N_14142);
and U15354 (N_15354,N_10437,N_10288);
nand U15355 (N_15355,N_13057,N_12134);
or U15356 (N_15356,N_12265,N_12693);
nand U15357 (N_15357,N_12609,N_14924);
xor U15358 (N_15358,N_13799,N_12054);
nand U15359 (N_15359,N_11461,N_10305);
nor U15360 (N_15360,N_11485,N_11912);
and U15361 (N_15361,N_13984,N_13322);
and U15362 (N_15362,N_14470,N_10330);
xor U15363 (N_15363,N_11023,N_11368);
nand U15364 (N_15364,N_12543,N_14469);
or U15365 (N_15365,N_13882,N_14851);
xnor U15366 (N_15366,N_10077,N_10173);
or U15367 (N_15367,N_10946,N_13625);
xor U15368 (N_15368,N_13000,N_12456);
and U15369 (N_15369,N_10639,N_11303);
and U15370 (N_15370,N_10279,N_14246);
and U15371 (N_15371,N_12217,N_14858);
xor U15372 (N_15372,N_14823,N_13930);
nand U15373 (N_15373,N_10312,N_12553);
nor U15374 (N_15374,N_12392,N_12400);
xnor U15375 (N_15375,N_12574,N_12501);
xor U15376 (N_15376,N_10341,N_13166);
and U15377 (N_15377,N_13324,N_13639);
xor U15378 (N_15378,N_11876,N_11138);
nor U15379 (N_15379,N_12058,N_12856);
xnor U15380 (N_15380,N_13798,N_14947);
or U15381 (N_15381,N_14365,N_14539);
nand U15382 (N_15382,N_12647,N_13948);
or U15383 (N_15383,N_13420,N_11621);
and U15384 (N_15384,N_14780,N_13373);
or U15385 (N_15385,N_10040,N_11208);
nand U15386 (N_15386,N_10754,N_10107);
nand U15387 (N_15387,N_12396,N_10963);
nor U15388 (N_15388,N_13100,N_10245);
nand U15389 (N_15389,N_11984,N_11650);
xor U15390 (N_15390,N_11124,N_10700);
or U15391 (N_15391,N_12041,N_13768);
nand U15392 (N_15392,N_10078,N_11546);
xnor U15393 (N_15393,N_14379,N_12779);
nor U15394 (N_15394,N_10390,N_10604);
nand U15395 (N_15395,N_10936,N_10866);
nor U15396 (N_15396,N_13459,N_14997);
xnor U15397 (N_15397,N_12171,N_11466);
xor U15398 (N_15398,N_10354,N_10899);
xnor U15399 (N_15399,N_12678,N_11260);
and U15400 (N_15400,N_14481,N_10195);
or U15401 (N_15401,N_11688,N_11599);
xnor U15402 (N_15402,N_10709,N_14651);
or U15403 (N_15403,N_12421,N_11144);
and U15404 (N_15404,N_10623,N_12556);
or U15405 (N_15405,N_10786,N_14802);
and U15406 (N_15406,N_12600,N_14135);
nand U15407 (N_15407,N_14262,N_10303);
nor U15408 (N_15408,N_13086,N_14860);
nor U15409 (N_15409,N_10458,N_13518);
and U15410 (N_15410,N_13299,N_11140);
or U15411 (N_15411,N_14874,N_14028);
nand U15412 (N_15412,N_13702,N_10586);
xor U15413 (N_15413,N_10172,N_12470);
nor U15414 (N_15414,N_10014,N_13780);
xnor U15415 (N_15415,N_13453,N_10738);
xnor U15416 (N_15416,N_10522,N_12873);
nand U15417 (N_15417,N_14243,N_13602);
xnor U15418 (N_15418,N_14190,N_11202);
or U15419 (N_15419,N_11516,N_10704);
nand U15420 (N_15420,N_12869,N_14088);
nand U15421 (N_15421,N_14483,N_13315);
nor U15422 (N_15422,N_10965,N_14099);
xor U15423 (N_15423,N_11534,N_10692);
nand U15424 (N_15424,N_13528,N_13781);
xnor U15425 (N_15425,N_11199,N_11181);
and U15426 (N_15426,N_14238,N_12242);
nand U15427 (N_15427,N_12139,N_14537);
and U15428 (N_15428,N_12985,N_10823);
xor U15429 (N_15429,N_11220,N_13637);
and U15430 (N_15430,N_13517,N_13090);
nor U15431 (N_15431,N_12223,N_13809);
nor U15432 (N_15432,N_14510,N_10410);
nor U15433 (N_15433,N_12472,N_12474);
nor U15434 (N_15434,N_14988,N_12740);
and U15435 (N_15435,N_11210,N_12724);
nand U15436 (N_15436,N_12459,N_13048);
and U15437 (N_15437,N_14086,N_10686);
xnor U15438 (N_15438,N_13582,N_10185);
nor U15439 (N_15439,N_10269,N_10716);
xnor U15440 (N_15440,N_11851,N_10814);
or U15441 (N_15441,N_11699,N_11059);
and U15442 (N_15442,N_14548,N_13444);
nor U15443 (N_15443,N_14919,N_13733);
nor U15444 (N_15444,N_11061,N_13761);
or U15445 (N_15445,N_12021,N_14253);
nor U15446 (N_15446,N_11759,N_12972);
and U15447 (N_15447,N_13970,N_13082);
nand U15448 (N_15448,N_12314,N_10930);
or U15449 (N_15449,N_10698,N_10948);
and U15450 (N_15450,N_12370,N_12404);
xor U15451 (N_15451,N_14450,N_13435);
and U15452 (N_15452,N_12732,N_10409);
nor U15453 (N_15453,N_10912,N_13221);
xnor U15454 (N_15454,N_10338,N_13731);
nor U15455 (N_15455,N_11294,N_12623);
xnor U15456 (N_15456,N_14563,N_14442);
xor U15457 (N_15457,N_10311,N_14321);
or U15458 (N_15458,N_11013,N_14654);
xor U15459 (N_15459,N_13466,N_11704);
nand U15460 (N_15460,N_13811,N_12520);
or U15461 (N_15461,N_10666,N_12737);
nor U15462 (N_15462,N_14411,N_14699);
xor U15463 (N_15463,N_14119,N_12437);
or U15464 (N_15464,N_11666,N_13191);
or U15465 (N_15465,N_14030,N_13740);
or U15466 (N_15466,N_13266,N_11452);
xnor U15467 (N_15467,N_10740,N_13016);
xnor U15468 (N_15468,N_11665,N_11706);
nand U15469 (N_15469,N_13954,N_11933);
xnor U15470 (N_15470,N_11491,N_11588);
and U15471 (N_15471,N_13792,N_11906);
and U15472 (N_15472,N_10500,N_11768);
nand U15473 (N_15473,N_13628,N_13137);
xnor U15474 (N_15474,N_14727,N_14575);
xnor U15475 (N_15475,N_13174,N_13536);
or U15476 (N_15476,N_14742,N_10404);
nor U15477 (N_15477,N_14898,N_11080);
or U15478 (N_15478,N_13028,N_13362);
nor U15479 (N_15479,N_12696,N_10618);
nand U15480 (N_15480,N_10011,N_10774);
nor U15481 (N_15481,N_12794,N_12731);
and U15482 (N_15482,N_14993,N_14431);
and U15483 (N_15483,N_12442,N_12895);
nor U15484 (N_15484,N_10635,N_11284);
and U15485 (N_15485,N_12776,N_14690);
and U15486 (N_15486,N_14485,N_10421);
nand U15487 (N_15487,N_10178,N_10641);
xor U15488 (N_15488,N_13285,N_12420);
nor U15489 (N_15489,N_12993,N_14731);
nand U15490 (N_15490,N_10663,N_10830);
nand U15491 (N_15491,N_10650,N_12398);
xor U15492 (N_15492,N_11934,N_11320);
and U15493 (N_15493,N_11473,N_11339);
nand U15494 (N_15494,N_13204,N_12368);
nor U15495 (N_15495,N_10070,N_10346);
nand U15496 (N_15496,N_14022,N_12864);
nand U15497 (N_15497,N_13004,N_10152);
and U15498 (N_15498,N_12862,N_11705);
nor U15499 (N_15499,N_12307,N_14599);
nor U15500 (N_15500,N_10171,N_10968);
nor U15501 (N_15501,N_13437,N_11713);
nand U15502 (N_15502,N_14448,N_14775);
or U15503 (N_15503,N_14282,N_10372);
nand U15504 (N_15504,N_11317,N_11781);
xnor U15505 (N_15505,N_11572,N_10620);
or U15506 (N_15506,N_14156,N_14468);
nand U15507 (N_15507,N_10084,N_12821);
xnor U15508 (N_15508,N_14363,N_12511);
nand U15509 (N_15509,N_13409,N_14370);
nor U15510 (N_15510,N_14748,N_14702);
nand U15511 (N_15511,N_14010,N_14040);
and U15512 (N_15512,N_12359,N_10792);
nand U15513 (N_15513,N_11111,N_13624);
nand U15514 (N_15514,N_13648,N_10911);
nand U15515 (N_15515,N_13563,N_10923);
and U15516 (N_15516,N_13123,N_10017);
nor U15517 (N_15517,N_13845,N_14972);
and U15518 (N_15518,N_13485,N_11156);
or U15519 (N_15519,N_11749,N_10507);
xor U15520 (N_15520,N_11790,N_14567);
and U15521 (N_15521,N_10356,N_12052);
or U15522 (N_15522,N_12062,N_14678);
nand U15523 (N_15523,N_13994,N_14794);
nand U15524 (N_15524,N_11958,N_13925);
nand U15525 (N_15525,N_10887,N_13181);
or U15526 (N_15526,N_11129,N_12603);
nand U15527 (N_15527,N_12621,N_13796);
or U15528 (N_15528,N_11048,N_11769);
and U15529 (N_15529,N_10227,N_13069);
and U15530 (N_15530,N_11297,N_12716);
xor U15531 (N_15531,N_11577,N_10134);
nand U15532 (N_15532,N_10362,N_11517);
xor U15533 (N_15533,N_14715,N_10664);
xnor U15534 (N_15534,N_12144,N_11712);
nor U15535 (N_15535,N_10369,N_14883);
and U15536 (N_15536,N_13555,N_13498);
nor U15537 (N_15537,N_10726,N_14345);
xnor U15538 (N_15538,N_14047,N_12951);
xnor U15539 (N_15539,N_10110,N_11484);
xnor U15540 (N_15540,N_14277,N_12506);
or U15541 (N_15541,N_14735,N_10052);
or U15542 (N_15542,N_12149,N_14003);
and U15543 (N_15543,N_14808,N_11823);
xnor U15544 (N_15544,N_10523,N_13682);
xor U15545 (N_15545,N_10406,N_12934);
xnor U15546 (N_15546,N_14798,N_12406);
xnor U15547 (N_15547,N_13806,N_14990);
or U15548 (N_15548,N_14534,N_13953);
nand U15549 (N_15549,N_10471,N_10573);
nand U15550 (N_15550,N_14863,N_13787);
nor U15551 (N_15551,N_11837,N_12077);
and U15552 (N_15552,N_11890,N_12476);
or U15553 (N_15553,N_10552,N_12789);
and U15554 (N_15554,N_14406,N_10430);
nor U15555 (N_15555,N_14953,N_10564);
nor U15556 (N_15556,N_13269,N_12319);
xnor U15557 (N_15557,N_13720,N_12327);
nor U15558 (N_15558,N_14888,N_13504);
nand U15559 (N_15559,N_11563,N_10232);
nor U15560 (N_15560,N_11085,N_14313);
xor U15561 (N_15561,N_13398,N_12829);
nand U15562 (N_15562,N_14896,N_11901);
nor U15563 (N_15563,N_12128,N_11605);
or U15564 (N_15564,N_13301,N_10089);
xor U15565 (N_15565,N_14710,N_12995);
nand U15566 (N_15566,N_10819,N_13950);
nor U15567 (N_15567,N_13064,N_10157);
nor U15568 (N_15568,N_12979,N_13641);
or U15569 (N_15569,N_10538,N_13546);
or U15570 (N_15570,N_12415,N_10841);
nor U15571 (N_15571,N_13693,N_13193);
xor U15572 (N_15572,N_10915,N_12667);
or U15573 (N_15573,N_11499,N_10877);
nor U15574 (N_15574,N_11022,N_14623);
xnor U15575 (N_15575,N_12331,N_12932);
and U15576 (N_15576,N_11514,N_13513);
xor U15577 (N_15577,N_10806,N_10898);
nand U15578 (N_15578,N_13464,N_14705);
nand U15579 (N_15579,N_12218,N_13835);
nor U15580 (N_15580,N_10867,N_11689);
and U15581 (N_15581,N_11070,N_10150);
and U15582 (N_15582,N_10609,N_10005);
nand U15583 (N_15583,N_13180,N_12068);
xor U15584 (N_15584,N_10363,N_14781);
nand U15585 (N_15585,N_12123,N_11944);
nand U15586 (N_15586,N_13011,N_11615);
nor U15587 (N_15587,N_12826,N_13652);
nor U15588 (N_15588,N_12657,N_12847);
or U15589 (N_15589,N_11381,N_13165);
nand U15590 (N_15590,N_13318,N_12714);
and U15591 (N_15591,N_12061,N_11121);
nor U15592 (N_15592,N_11357,N_12548);
or U15593 (N_15593,N_13957,N_12407);
nand U15594 (N_15594,N_13062,N_13406);
nor U15595 (N_15595,N_13627,N_14434);
and U15596 (N_15596,N_13345,N_12227);
nor U15597 (N_15597,N_13293,N_13275);
nor U15598 (N_15598,N_12180,N_10439);
nand U15599 (N_15599,N_13943,N_11469);
xnor U15600 (N_15600,N_12292,N_11946);
nand U15601 (N_15601,N_10479,N_11684);
xnor U15602 (N_15602,N_10337,N_10622);
xnor U15603 (N_15603,N_13184,N_14473);
xnor U15604 (N_15604,N_10937,N_10524);
nor U15605 (N_15605,N_11247,N_12739);
and U15606 (N_15606,N_12081,N_10875);
xnor U15607 (N_15607,N_10015,N_11405);
nor U15608 (N_15608,N_12075,N_10204);
nand U15609 (N_15609,N_14952,N_11429);
nand U15610 (N_15610,N_14881,N_10393);
xor U15611 (N_15611,N_13185,N_14809);
and U15612 (N_15612,N_13058,N_13831);
nand U15613 (N_15613,N_12475,N_10561);
and U15614 (N_15614,N_14424,N_14950);
or U15615 (N_15615,N_10349,N_11043);
or U15616 (N_15616,N_11883,N_14987);
and U15617 (N_15617,N_11834,N_13457);
and U15618 (N_15618,N_13486,N_12257);
or U15619 (N_15619,N_12588,N_13716);
and U15620 (N_15620,N_11600,N_10682);
and U15621 (N_15621,N_12231,N_13618);
or U15622 (N_15622,N_14836,N_10139);
xnor U15623 (N_15623,N_13915,N_11882);
and U15624 (N_15624,N_13622,N_13292);
nor U15625 (N_15625,N_13851,N_14634);
nand U15626 (N_15626,N_12778,N_11264);
xor U15627 (N_15627,N_13272,N_13644);
xnor U15628 (N_15628,N_10771,N_12424);
nor U15629 (N_15629,N_11158,N_11159);
and U15630 (N_15630,N_13055,N_10450);
nand U15631 (N_15631,N_10127,N_13334);
nand U15632 (N_15632,N_10918,N_10891);
xnor U15633 (N_15633,N_11798,N_10082);
or U15634 (N_15634,N_10840,N_11856);
or U15635 (N_15635,N_12840,N_10732);
nand U15636 (N_15636,N_10074,N_12059);
and U15637 (N_15637,N_11682,N_14824);
nand U15638 (N_15638,N_14143,N_10568);
nor U15639 (N_15639,N_14506,N_12580);
or U15640 (N_15640,N_14200,N_11006);
nor U15641 (N_15641,N_12019,N_11505);
nand U15642 (N_15642,N_10625,N_11253);
and U15643 (N_15643,N_10301,N_10739);
and U15644 (N_15644,N_13465,N_14970);
nand U15645 (N_15645,N_14136,N_14718);
and U15646 (N_15646,N_14439,N_14062);
nand U15647 (N_15647,N_13659,N_14819);
or U15648 (N_15648,N_11904,N_10646);
and U15649 (N_15649,N_12749,N_12391);
nand U15650 (N_15650,N_11829,N_12956);
and U15651 (N_15651,N_14958,N_12659);
nor U15652 (N_15652,N_14762,N_11408);
nand U15653 (N_15653,N_13371,N_13346);
xor U15654 (N_15654,N_12689,N_11559);
and U15655 (N_15655,N_12752,N_14404);
or U15656 (N_15656,N_13297,N_10548);
xnor U15657 (N_15657,N_13240,N_13615);
xor U15658 (N_15658,N_11596,N_13078);
nand U15659 (N_15659,N_14936,N_12345);
xor U15660 (N_15660,N_14635,N_11126);
or U15661 (N_15661,N_10873,N_11593);
nor U15662 (N_15662,N_13416,N_14976);
nand U15663 (N_15663,N_14895,N_13156);
nand U15664 (N_15664,N_12312,N_14893);
nand U15665 (N_15665,N_13554,N_12089);
and U15666 (N_15666,N_11213,N_13556);
or U15667 (N_15667,N_14134,N_11239);
and U15668 (N_15668,N_10449,N_12827);
and U15669 (N_15669,N_12362,N_14407);
and U15670 (N_15670,N_14646,N_11677);
and U15671 (N_15671,N_12147,N_14825);
and U15672 (N_15672,N_12542,N_13441);
or U15673 (N_15673,N_10910,N_12358);
nor U15674 (N_15674,N_14649,N_13993);
nor U15675 (N_15675,N_13366,N_11106);
or U15676 (N_15676,N_13786,N_12086);
or U15677 (N_15677,N_13535,N_12509);
or U15678 (N_15678,N_12713,N_10447);
nand U15679 (N_15679,N_12353,N_14038);
and U15680 (N_15680,N_14572,N_10659);
and U15681 (N_15681,N_14520,N_12412);
xor U15682 (N_15682,N_12182,N_14122);
nand U15683 (N_15683,N_13710,N_14275);
nand U15684 (N_15684,N_14271,N_12355);
nand U15685 (N_15685,N_14340,N_11745);
xor U15686 (N_15686,N_10895,N_14908);
nand U15687 (N_15687,N_10714,N_11173);
and U15688 (N_15688,N_13672,N_13629);
and U15689 (N_15689,N_13758,N_10928);
and U15690 (N_15690,N_10986,N_12453);
or U15691 (N_15691,N_10532,N_14701);
nand U15692 (N_15692,N_11968,N_12403);
and U15693 (N_15693,N_10816,N_14523);
nand U15694 (N_15694,N_13532,N_10960);
nand U15695 (N_15695,N_10812,N_14975);
and U15696 (N_15696,N_13258,N_11164);
nand U15697 (N_15697,N_13313,N_14935);
nand U15698 (N_15698,N_10023,N_10431);
and U15699 (N_15699,N_10058,N_11603);
xor U15700 (N_15700,N_12356,N_13474);
nand U15701 (N_15701,N_10095,N_13841);
or U15702 (N_15702,N_14662,N_10175);
xnor U15703 (N_15703,N_14498,N_14412);
nand U15704 (N_15704,N_14594,N_10848);
nor U15705 (N_15705,N_11336,N_13047);
or U15706 (N_15706,N_10897,N_13501);
or U15707 (N_15707,N_11184,N_13245);
nand U15708 (N_15708,N_14907,N_10558);
and U15709 (N_15709,N_12708,N_13033);
xnor U15710 (N_15710,N_14722,N_13044);
nand U15711 (N_15711,N_11935,N_14069);
nand U15712 (N_15712,N_10004,N_11627);
nand U15713 (N_15713,N_13227,N_11616);
or U15714 (N_15714,N_13231,N_11030);
nor U15715 (N_15715,N_12612,N_13288);
and U15716 (N_15716,N_11841,N_14445);
and U15717 (N_15717,N_14016,N_13414);
nor U15718 (N_15718,N_11379,N_14358);
or U15719 (N_15719,N_10168,N_12439);
or U15720 (N_15720,N_14578,N_14344);
nand U15721 (N_15721,N_14254,N_14035);
and U15722 (N_15722,N_13638,N_10251);
or U15723 (N_15723,N_14269,N_12694);
xor U15724 (N_15724,N_14998,N_11793);
nand U15725 (N_15725,N_11649,N_11474);
or U15726 (N_15726,N_11584,N_13046);
or U15727 (N_15727,N_10794,N_11620);
nor U15728 (N_15728,N_10187,N_13891);
nor U15729 (N_15729,N_12517,N_10436);
nand U15730 (N_15730,N_10803,N_13952);
and U15731 (N_15731,N_14713,N_13817);
nand U15732 (N_15732,N_12589,N_14236);
nand U15733 (N_15733,N_14303,N_11861);
or U15734 (N_15734,N_10901,N_13175);
nor U15735 (N_15735,N_13115,N_14373);
nand U15736 (N_15736,N_11545,N_11862);
nand U15737 (N_15737,N_10962,N_11960);
xor U15738 (N_15738,N_10035,N_14880);
or U15739 (N_15739,N_14869,N_10101);
and U15740 (N_15740,N_11257,N_11807);
nand U15741 (N_15741,N_11226,N_11859);
or U15742 (N_15742,N_11244,N_11877);
or U15743 (N_15743,N_11740,N_12029);
and U15744 (N_15744,N_11020,N_12702);
and U15745 (N_15745,N_11773,N_11843);
nand U15746 (N_15746,N_14904,N_11776);
or U15747 (N_15747,N_14178,N_10262);
and U15748 (N_15748,N_12711,N_12240);
xnor U15749 (N_15749,N_13691,N_12252);
nand U15750 (N_15750,N_12369,N_10494);
nor U15751 (N_15751,N_14288,N_10126);
or U15752 (N_15752,N_13631,N_11252);
and U15753 (N_15753,N_13801,N_13481);
xor U15754 (N_15754,N_11455,N_12458);
and U15755 (N_15755,N_12288,N_11978);
nand U15756 (N_15756,N_13068,N_10278);
nand U15757 (N_15757,N_10348,N_14018);
nand U15758 (N_15758,N_14655,N_13260);
xnor U15759 (N_15759,N_14664,N_13213);
or U15760 (N_15760,N_13151,N_14850);
xnor U15761 (N_15761,N_13686,N_12660);
and U15762 (N_15762,N_11040,N_10633);
xnor U15763 (N_15763,N_10810,N_11679);
xnor U15764 (N_15764,N_11439,N_14598);
nor U15765 (N_15765,N_12505,N_14017);
nor U15766 (N_15766,N_10616,N_13662);
nand U15767 (N_15767,N_12377,N_13045);
or U15768 (N_15768,N_11410,N_13932);
nand U15769 (N_15769,N_13502,N_13310);
nor U15770 (N_15770,N_14159,N_10590);
nor U15771 (N_15771,N_10741,N_11567);
xor U15772 (N_15772,N_11900,N_14041);
or U15773 (N_15773,N_12721,N_11453);
xnor U15774 (N_15774,N_10989,N_11192);
nand U15775 (N_15775,N_11092,N_12540);
nand U15776 (N_15776,N_10466,N_10257);
or U15777 (N_15777,N_12361,N_12611);
and U15778 (N_15778,N_13341,N_12350);
nand U15779 (N_15779,N_12809,N_10407);
xor U15780 (N_15780,N_10221,N_10088);
and U15781 (N_15781,N_11871,N_14650);
nand U15782 (N_15782,N_10637,N_10256);
nand U15783 (N_15783,N_11432,N_12326);
and U15784 (N_15784,N_10207,N_11905);
nor U15785 (N_15785,N_11038,N_13489);
nand U15786 (N_15786,N_12759,N_14930);
nand U15787 (N_15787,N_10367,N_13010);
and U15788 (N_15788,N_13140,N_12329);
nor U15789 (N_15789,N_14301,N_14385);
or U15790 (N_15790,N_14905,N_12239);
xor U15791 (N_15791,N_12531,N_13402);
or U15792 (N_15792,N_14044,N_12195);
nor U15793 (N_15793,N_10008,N_10603);
and U15794 (N_15794,N_11133,N_10991);
nor U15795 (N_15795,N_11235,N_12216);
and U15796 (N_15796,N_10863,N_13253);
nor U15797 (N_15797,N_11292,N_12340);
and U15798 (N_15798,N_12717,N_13169);
nor U15799 (N_15799,N_12005,N_11508);
nor U15800 (N_15800,N_14273,N_14928);
nor U15801 (N_15801,N_12050,N_14388);
or U15802 (N_15802,N_11709,N_10468);
xnor U15803 (N_15803,N_12210,N_11932);
xnor U15804 (N_15804,N_13819,N_14339);
and U15805 (N_15805,N_13325,N_11426);
or U15806 (N_15806,N_13385,N_12422);
nand U15807 (N_15807,N_12961,N_11127);
nand U15808 (N_15808,N_13393,N_10132);
nand U15809 (N_15809,N_11403,N_12817);
xor U15810 (N_15810,N_11028,N_13692);
and U15811 (N_15811,N_14676,N_11131);
xor U15812 (N_15812,N_11067,N_14077);
nor U15813 (N_15813,N_14380,N_14270);
nand U15814 (N_15814,N_13920,N_12283);
nand U15815 (N_15815,N_13201,N_12383);
nand U15816 (N_15816,N_12836,N_11026);
nand U15817 (N_15817,N_12544,N_11396);
or U15818 (N_15818,N_12642,N_10517);
or U15819 (N_15819,N_10336,N_14308);
and U15820 (N_15820,N_11412,N_10805);
nand U15821 (N_15821,N_13997,N_10402);
nor U15822 (N_15822,N_13510,N_10316);
xor U15823 (N_15823,N_10066,N_11400);
and U15824 (N_15824,N_10214,N_13132);
nor U15825 (N_15825,N_12547,N_14558);
and U15826 (N_15826,N_12680,N_14961);
nand U15827 (N_15827,N_13881,N_13726);
and U15828 (N_15828,N_13192,N_11797);
nor U15829 (N_15829,N_13017,N_12703);
nand U15830 (N_15830,N_11263,N_13277);
and U15831 (N_15831,N_12169,N_12479);
xnor U15832 (N_15832,N_11113,N_13757);
or U15833 (N_15833,N_12440,N_11686);
xnor U15834 (N_15834,N_14292,N_10420);
nand U15835 (N_15835,N_13383,N_14818);
nor U15836 (N_15836,N_13597,N_14920);
nand U15837 (N_15837,N_13642,N_12839);
nor U15838 (N_15838,N_12380,N_14628);
or U15839 (N_15839,N_14149,N_12477);
nand U15840 (N_15840,N_10600,N_13812);
xor U15841 (N_15841,N_12976,N_14688);
or U15842 (N_15842,N_11215,N_12607);
nor U15843 (N_15843,N_13212,N_10973);
nor U15844 (N_15844,N_10112,N_10131);
and U15845 (N_15845,N_12593,N_10780);
nand U15846 (N_15846,N_10837,N_14938);
and U15847 (N_15847,N_13523,N_14341);
xnor U15848 (N_15848,N_14327,N_12289);
or U15849 (N_15849,N_10412,N_11463);
xor U15850 (N_15850,N_14927,N_12616);
nor U15851 (N_15851,N_11128,N_12306);
nor U15852 (N_15852,N_13244,N_12929);
and U15853 (N_15853,N_11483,N_14899);
nand U15854 (N_15854,N_10121,N_10521);
and U15855 (N_15855,N_11307,N_11509);
or U15856 (N_15856,N_13179,N_10396);
or U15857 (N_15857,N_14169,N_13750);
and U15858 (N_15858,N_11250,N_12725);
xor U15859 (N_15859,N_12489,N_10563);
and U15860 (N_15860,N_10467,N_14078);
nor U15861 (N_15861,N_14432,N_12296);
or U15862 (N_15862,N_11513,N_10744);
and U15863 (N_15863,N_11322,N_12538);
xor U15864 (N_15864,N_10708,N_11870);
nand U15865 (N_15865,N_13381,N_12335);
xnor U15866 (N_15866,N_13982,N_11983);
and U15867 (N_15867,N_10921,N_10091);
or U15868 (N_15868,N_13106,N_14163);
and U15869 (N_15869,N_10291,N_10465);
nand U15870 (N_15870,N_11637,N_13776);
nand U15871 (N_15871,N_13917,N_14272);
xnor U15872 (N_15872,N_11341,N_14438);
nand U15873 (N_15873,N_10518,N_12823);
nor U15874 (N_15874,N_11959,N_11318);
or U15875 (N_15875,N_12140,N_12806);
or U15876 (N_15876,N_11204,N_13861);
or U15877 (N_15877,N_11695,N_13241);
nor U15878 (N_15878,N_13607,N_11974);
nand U15879 (N_15879,N_14167,N_12270);
nand U15880 (N_15880,N_10166,N_14132);
nand U15881 (N_15881,N_11018,N_14317);
nand U15882 (N_15882,N_10730,N_11568);
xnor U15883 (N_15883,N_11835,N_12131);
and U15884 (N_15884,N_11708,N_12338);
nor U15885 (N_15885,N_14792,N_11063);
nor U15886 (N_15886,N_12497,N_13526);
nor U15887 (N_15887,N_11081,N_10025);
nand U15888 (N_15888,N_13284,N_12743);
and U15889 (N_15889,N_12893,N_13079);
or U15890 (N_15890,N_13852,N_14416);
nand U15891 (N_15891,N_11082,N_13834);
or U15892 (N_15892,N_11223,N_13700);
nor U15893 (N_15893,N_14068,N_14105);
nor U15894 (N_15894,N_10193,N_14771);
nor U15895 (N_15895,N_11632,N_14000);
nor U15896 (N_15896,N_12135,N_12728);
nand U15897 (N_15897,N_12900,N_11401);
nand U15898 (N_15898,N_10247,N_13470);
and U15899 (N_15899,N_10275,N_13697);
nor U15900 (N_15900,N_13992,N_12886);
nor U15901 (N_15901,N_10787,N_12656);
nor U15902 (N_15902,N_13810,N_10128);
or U15903 (N_15903,N_14075,N_11224);
and U15904 (N_15904,N_10216,N_12279);
and U15905 (N_15905,N_10673,N_11633);
or U15906 (N_15906,N_13940,N_12787);
and U15907 (N_15907,N_13194,N_13367);
nand U15908 (N_15908,N_10092,N_12299);
nor U15909 (N_15909,N_11489,N_11225);
nand U15910 (N_15910,N_12529,N_11779);
nand U15911 (N_15911,N_11145,N_11910);
nor U15912 (N_15912,N_12668,N_14264);
or U15913 (N_15913,N_13434,N_13189);
or U15914 (N_15914,N_14055,N_11103);
xor U15915 (N_15915,N_11179,N_14674);
nand U15916 (N_15916,N_11036,N_10451);
xor U15917 (N_15917,N_11169,N_12016);
nand U15918 (N_15918,N_11456,N_11440);
nor U15919 (N_15919,N_14918,N_12212);
nor U15920 (N_15920,N_13247,N_11685);
and U15921 (N_15921,N_12300,N_14846);
and U15922 (N_15922,N_10296,N_10657);
or U15923 (N_15923,N_12493,N_11290);
nand U15924 (N_15924,N_10723,N_12194);
or U15925 (N_15925,N_14322,N_14224);
and U15926 (N_15926,N_11720,N_14256);
nand U15927 (N_15927,N_13395,N_10815);
nand U15928 (N_15928,N_12295,N_12367);
xnor U15929 (N_15929,N_13537,N_12535);
nor U15930 (N_15930,N_12537,N_10133);
or U15931 (N_15931,N_10990,N_13808);
or U15932 (N_15932,N_12919,N_14426);
and U15933 (N_15933,N_11523,N_12665);
xor U15934 (N_15934,N_13748,N_11628);
and U15935 (N_15935,N_13636,N_13375);
nand U15936 (N_15936,N_14620,N_11217);
and U15937 (N_15937,N_11419,N_14969);
xnor U15938 (N_15938,N_11765,N_10506);
nand U15939 (N_15939,N_14386,N_11241);
and U15940 (N_15940,N_14285,N_13094);
xor U15941 (N_15941,N_10501,N_10826);
nand U15942 (N_15942,N_13431,N_11168);
or U15943 (N_15943,N_10756,N_10702);
xor U15944 (N_15944,N_12568,N_10167);
nand U15945 (N_15945,N_13391,N_10705);
and U15946 (N_15946,N_13358,N_14444);
nand U15947 (N_15947,N_13080,N_12243);
nor U15948 (N_15948,N_13844,N_13473);
nand U15949 (N_15949,N_11681,N_11084);
and U15950 (N_15950,N_12673,N_10886);
or U15951 (N_15951,N_11034,N_13330);
nor U15952 (N_15952,N_12297,N_13238);
xor U15953 (N_15953,N_13668,N_13989);
or U15954 (N_15954,N_13146,N_11556);
nor U15955 (N_15955,N_12427,N_13202);
and U15956 (N_15956,N_10164,N_10872);
and U15957 (N_15957,N_14391,N_10993);
or U15958 (N_15958,N_12871,N_14453);
nor U15959 (N_15959,N_11175,N_11269);
nor U15960 (N_15960,N_11818,N_13363);
or U15961 (N_15961,N_13859,N_10141);
and U15962 (N_15962,N_10531,N_11525);
nand U15963 (N_15963,N_10308,N_11638);
xor U15964 (N_15964,N_11928,N_11409);
nor U15965 (N_15965,N_14032,N_13021);
nand U15966 (N_15966,N_14756,N_13236);
or U15967 (N_15967,N_12784,N_14789);
nand U15968 (N_15968,N_11096,N_10473);
or U15969 (N_15969,N_10464,N_10706);
or U15970 (N_15970,N_14503,N_10229);
or U15971 (N_15971,N_12897,N_14917);
or U15972 (N_15972,N_14472,N_11548);
or U15973 (N_15973,N_10250,N_12430);
nand U15974 (N_15974,N_13368,N_14937);
nand U15975 (N_15975,N_12571,N_11172);
nor U15976 (N_15976,N_10519,N_12018);
nand U15977 (N_15977,N_11037,N_12346);
nand U15978 (N_15978,N_12853,N_14180);
and U15979 (N_15979,N_14695,N_13975);
nor U15980 (N_15980,N_13487,N_14129);
or U15981 (N_15981,N_12200,N_14589);
nor U15982 (N_15982,N_13928,N_14486);
and U15983 (N_15983,N_10159,N_12682);
and U15984 (N_15984,N_11707,N_13505);
and U15985 (N_15985,N_11503,N_14500);
nand U15986 (N_15986,N_12111,N_14220);
nor U15987 (N_15987,N_12772,N_10995);
nor U15988 (N_15988,N_11828,N_12819);
nor U15989 (N_15989,N_14884,N_12078);
xor U15990 (N_15990,N_14799,N_13573);
or U15991 (N_15991,N_14725,N_10798);
xnor U15992 (N_15992,N_11014,N_12113);
nand U15993 (N_15993,N_14405,N_13461);
nand U15994 (N_15994,N_14885,N_13215);
nor U15995 (N_15995,N_13274,N_14530);
and U15996 (N_15996,N_12899,N_12150);
and U15997 (N_15997,N_12803,N_11492);
xnor U15998 (N_15998,N_10902,N_11100);
nor U15999 (N_15999,N_11442,N_11203);
xor U16000 (N_16000,N_11598,N_12071);
and U16001 (N_16001,N_12883,N_13312);
xnor U16002 (N_16002,N_12965,N_12126);
xnor U16003 (N_16003,N_12602,N_10855);
nand U16004 (N_16004,N_10820,N_12133);
and U16005 (N_16005,N_11825,N_10888);
xor U16006 (N_16006,N_12581,N_12590);
nor U16007 (N_16007,N_14318,N_12692);
nor U16008 (N_16008,N_14488,N_11487);
and U16009 (N_16009,N_14141,N_11479);
xor U16010 (N_16010,N_13619,N_12154);
nand U16011 (N_16011,N_14206,N_10781);
xnor U16012 (N_16012,N_13263,N_13756);
nand U16013 (N_16013,N_14235,N_12460);
nand U16014 (N_16014,N_11506,N_11375);
nor U16015 (N_16015,N_11985,N_10331);
nor U16016 (N_16016,N_13176,N_12386);
or U16017 (N_16017,N_12688,N_14103);
or U16018 (N_16018,N_12832,N_12191);
xor U16019 (N_16019,N_11472,N_11470);
or U16020 (N_16020,N_11535,N_12015);
or U16021 (N_16021,N_14179,N_13655);
or U16022 (N_16022,N_11441,N_13203);
nand U16023 (N_16023,N_14618,N_12984);
xor U16024 (N_16024,N_11275,N_13447);
xnor U16025 (N_16025,N_13888,N_12409);
nor U16026 (N_16026,N_12310,N_11186);
nor U16027 (N_16027,N_11889,N_11174);
nor U16028 (N_16028,N_11012,N_14659);
xnor U16029 (N_16029,N_12908,N_11364);
or U16030 (N_16030,N_13942,N_12549);
nor U16031 (N_16031,N_14853,N_14263);
and U16032 (N_16032,N_11019,N_10534);
nand U16033 (N_16033,N_11966,N_14061);
nand U16034 (N_16034,N_12066,N_11971);
or U16035 (N_16035,N_11515,N_13088);
nand U16036 (N_16036,N_12073,N_10445);
xnor U16037 (N_16037,N_12924,N_14466);
or U16038 (N_16038,N_10589,N_11853);
or U16039 (N_16039,N_11150,N_13355);
xnor U16040 (N_16040,N_10770,N_14203);
nand U16041 (N_16041,N_10188,N_11750);
and U16042 (N_16042,N_13564,N_11136);
xnor U16043 (N_16043,N_11104,N_14597);
xor U16044 (N_16044,N_12814,N_14636);
and U16045 (N_16045,N_12828,N_13507);
xor U16046 (N_16046,N_12251,N_11233);
or U16047 (N_16047,N_10432,N_14192);
nand U16048 (N_16048,N_11662,N_13675);
nand U16049 (N_16049,N_10334,N_14007);
and U16050 (N_16050,N_12025,N_12774);
nand U16051 (N_16051,N_11758,N_10950);
nand U16052 (N_16052,N_13508,N_10380);
or U16053 (N_16053,N_14977,N_11752);
and U16054 (N_16054,N_11007,N_14687);
or U16055 (N_16055,N_11550,N_12120);
nor U16056 (N_16056,N_11279,N_12852);
nor U16057 (N_16057,N_14683,N_11392);
xor U16058 (N_16058,N_12903,N_12861);
nor U16059 (N_16059,N_12190,N_10533);
xor U16060 (N_16060,N_12882,N_10302);
nand U16061 (N_16061,N_13791,N_11907);
and U16062 (N_16062,N_13428,N_13443);
and U16063 (N_16063,N_12559,N_12152);
nor U16064 (N_16064,N_14774,N_13162);
xor U16065 (N_16065,N_12788,N_11430);
nor U16066 (N_16066,N_13738,N_12039);
and U16067 (N_16067,N_13138,N_14584);
and U16068 (N_16068,N_13722,N_13867);
xnor U16069 (N_16069,N_10002,N_14118);
or U16070 (N_16070,N_12498,N_12387);
xor U16071 (N_16071,N_12698,N_13689);
or U16072 (N_16072,N_10772,N_12037);
nor U16073 (N_16073,N_14502,N_10789);
nand U16074 (N_16074,N_13449,N_13929);
nand U16075 (N_16075,N_11097,N_13931);
nand U16076 (N_16076,N_11011,N_11520);
nor U16077 (N_16077,N_10161,N_10969);
nor U16078 (N_16078,N_10880,N_13134);
or U16079 (N_16079,N_13525,N_14542);
and U16080 (N_16080,N_10212,N_14402);
and U16081 (N_16081,N_12333,N_12177);
nand U16082 (N_16082,N_14493,N_12173);
or U16083 (N_16083,N_10297,N_14475);
or U16084 (N_16084,N_12484,N_11717);
xnor U16085 (N_16085,N_14008,N_14052);
or U16086 (N_16086,N_12896,N_13248);
or U16087 (N_16087,N_13736,N_11274);
nand U16088 (N_16088,N_13490,N_14640);
nor U16089 (N_16089,N_11064,N_10808);
or U16090 (N_16090,N_11751,N_14875);
nor U16091 (N_16091,N_14131,N_10038);
xor U16092 (N_16092,N_11763,N_12146);
and U16093 (N_16093,N_11278,N_11062);
nand U16094 (N_16094,N_12639,N_12554);
nor U16095 (N_16095,N_12097,N_11161);
or U16096 (N_16096,N_13195,N_14261);
or U16097 (N_16097,N_13255,N_11537);
or U16098 (N_16098,N_14013,N_13197);
nor U16099 (N_16099,N_10069,N_13609);
or U16100 (N_16100,N_13059,N_12950);
xnor U16101 (N_16101,N_14728,N_13276);
nor U16102 (N_16102,N_13305,N_13956);
nor U16103 (N_16103,N_11369,N_13559);
xor U16104 (N_16104,N_12780,N_14949);
nand U16105 (N_16105,N_14951,N_10378);
or U16106 (N_16106,N_11271,N_12163);
and U16107 (N_16107,N_11259,N_11194);
and U16108 (N_16108,N_10246,N_10106);
nor U16109 (N_16109,N_10018,N_10970);
and U16110 (N_16110,N_13515,N_14334);
nor U16111 (N_16111,N_11897,N_10137);
nand U16112 (N_16112,N_12290,N_13372);
and U16113 (N_16113,N_14693,N_14996);
nor U16114 (N_16114,N_10576,N_13415);
or U16115 (N_16115,N_11635,N_10183);
xnor U16116 (N_16116,N_14782,N_14660);
xnor U16117 (N_16117,N_12083,N_13200);
and U16118 (N_16118,N_10540,N_13544);
nand U16119 (N_16119,N_10783,N_11714);
xor U16120 (N_16120,N_14673,N_10382);
nor U16121 (N_16121,N_10345,N_10003);
or U16122 (N_16122,N_11973,N_11343);
and U16123 (N_16123,N_11229,N_11243);
or U16124 (N_16124,N_10086,N_11702);
or U16125 (N_16125,N_10889,N_12876);
and U16126 (N_16126,N_10293,N_10914);
or U16127 (N_16127,N_12411,N_11561);
nand U16128 (N_16128,N_12055,N_11355);
and U16129 (N_16129,N_12309,N_14217);
nor U16130 (N_16130,N_12619,N_13968);
and U16131 (N_16131,N_11119,N_11955);
and U16132 (N_16132,N_10055,N_14219);
and U16133 (N_16133,N_14577,N_12313);
nor U16134 (N_16134,N_14826,N_13816);
xor U16135 (N_16135,N_13050,N_11587);
nand U16136 (N_16136,N_13218,N_13978);
nor U16137 (N_16137,N_12863,N_10032);
nand U16138 (N_16138,N_14377,N_11996);
or U16139 (N_16139,N_11915,N_12585);
xor U16140 (N_16140,N_12485,N_11716);
and U16141 (N_16141,N_14144,N_14831);
or U16142 (N_16142,N_12230,N_12536);
nand U16143 (N_16143,N_10566,N_11495);
xor U16144 (N_16144,N_11850,N_12744);
and U16145 (N_16145,N_12921,N_10162);
xnor U16146 (N_16146,N_10388,N_11298);
and U16147 (N_16147,N_10883,N_11471);
xnor U16148 (N_16148,N_11394,N_11937);
nor U16149 (N_16149,N_14338,N_10029);
nand U16150 (N_16150,N_11212,N_13446);
and U16151 (N_16151,N_13417,N_10913);
and U16152 (N_16152,N_13206,N_14231);
xor U16153 (N_16153,N_14868,N_14364);
and U16154 (N_16154,N_11547,N_13149);
and U16155 (N_16155,N_11887,N_13530);
and U16156 (N_16156,N_11295,N_12891);
xnor U16157 (N_16157,N_10842,N_12162);
or U16158 (N_16158,N_12618,N_10324);
nand U16159 (N_16159,N_12504,N_12298);
nor U16160 (N_16160,N_12569,N_13351);
xnor U16161 (N_16161,N_14955,N_11977);
and U16162 (N_16162,N_10711,N_12064);
nand U16163 (N_16163,N_12454,N_13893);
or U16164 (N_16164,N_13906,N_14392);
nor U16165 (N_16165,N_10281,N_10927);
nor U16166 (N_16166,N_10254,N_14296);
nand U16167 (N_16167,N_12655,N_14297);
and U16168 (N_16168,N_13921,N_11544);
nor U16169 (N_16169,N_10851,N_10205);
and U16170 (N_16170,N_12366,N_10513);
and U16171 (N_16171,N_14039,N_10113);
nand U16172 (N_16172,N_14371,N_12677);
xor U16173 (N_16173,N_11655,N_12253);
nor U16174 (N_16174,N_13813,N_12085);
nand U16175 (N_16175,N_13264,N_14125);
xor U16176 (N_16176,N_13965,N_10685);
nor U16177 (N_16177,N_12098,N_13613);
nor U16178 (N_16178,N_13405,N_11571);
nor U16179 (N_16179,N_13849,N_12996);
or U16180 (N_16180,N_10019,N_10399);
or U16181 (N_16181,N_10119,N_11687);
xnor U16182 (N_16182,N_11939,N_13986);
nor U16183 (N_16183,N_13587,N_13981);
nor U16184 (N_16184,N_11590,N_10502);
or U16185 (N_16185,N_11994,N_11868);
or U16186 (N_16186,N_12201,N_10640);
nand U16187 (N_16187,N_13558,N_10629);
or U16188 (N_16188,N_10114,N_10422);
and U16189 (N_16189,N_14189,N_13739);
or U16190 (N_16190,N_10176,N_14637);
nand U16191 (N_16191,N_10325,N_11770);
or U16192 (N_16192,N_10849,N_11643);
and U16193 (N_16193,N_10230,N_11338);
nor U16194 (N_16194,N_14670,N_11049);
nor U16195 (N_16195,N_11943,N_14465);
nand U16196 (N_16196,N_11221,N_11398);
nor U16197 (N_16197,N_13019,N_14588);
nor U16198 (N_16198,N_13751,N_11927);
and U16199 (N_16199,N_13540,N_13856);
nor U16200 (N_16200,N_14583,N_14776);
and U16201 (N_16201,N_10608,N_13377);
nand U16202 (N_16202,N_10621,N_14307);
nand U16203 (N_16203,N_11913,N_14198);
nand U16204 (N_16204,N_13890,N_13516);
nor U16205 (N_16205,N_10530,N_11981);
and U16206 (N_16206,N_13388,N_10192);
nor U16207 (N_16207,N_14009,N_10601);
xor U16208 (N_16208,N_13067,N_14350);
and U16209 (N_16209,N_12645,N_11724);
nand U16210 (N_16210,N_12938,N_13328);
nand U16211 (N_16211,N_13178,N_13727);
xnor U16212 (N_16212,N_12137,N_12608);
xor U16213 (N_16213,N_10495,N_13101);
nor U16214 (N_16214,N_10612,N_10242);
and U16215 (N_16215,N_12953,N_14257);
or U16216 (N_16216,N_13163,N_10943);
nor U16217 (N_16217,N_11723,N_12981);
xor U16218 (N_16218,N_14241,N_14333);
nand U16219 (N_16219,N_11321,N_14494);
or U16220 (N_16220,N_14315,N_12116);
or U16221 (N_16221,N_14095,N_12160);
nand U16222 (N_16222,N_11618,N_10998);
or U16223 (N_16223,N_11657,N_11041);
and U16224 (N_16224,N_11052,N_12100);
nand U16225 (N_16225,N_12248,N_13680);
and U16226 (N_16226,N_11139,N_10610);
and U16227 (N_16227,N_10031,N_11060);
xnor U16228 (N_16228,N_10571,N_10287);
and U16229 (N_16229,N_11120,N_10010);
nor U16230 (N_16230,N_10747,N_11232);
nor U16231 (N_16231,N_10469,N_11858);
xnor U16232 (N_16232,N_10557,N_10735);
xnor U16233 (N_16233,N_14903,N_11480);
and U16234 (N_16234,N_10862,N_13825);
and U16235 (N_16235,N_13408,N_14614);
and U16236 (N_16236,N_10319,N_14429);
and U16237 (N_16237,N_14076,N_11810);
and U16238 (N_16238,N_12006,N_13914);
and U16239 (N_16239,N_13923,N_13960);
and U16240 (N_16240,N_13879,N_13865);
or U16241 (N_16241,N_13374,N_10582);
nor U16242 (N_16242,N_14274,N_13894);
nor U16243 (N_16243,N_12381,N_11325);
nand U16244 (N_16244,N_14096,N_10240);
and U16245 (N_16245,N_11578,N_12905);
and U16246 (N_16246,N_12360,N_14352);
or U16247 (N_16247,N_11742,N_11160);
or U16248 (N_16248,N_14228,N_13356);
or U16249 (N_16249,N_14126,N_12804);
or U16250 (N_16250,N_12438,N_13267);
or U16251 (N_16251,N_13549,N_13553);
and U16252 (N_16252,N_14681,N_14319);
nor U16253 (N_16253,N_13496,N_12675);
nand U16254 (N_16254,N_14115,N_10959);
or U16255 (N_16255,N_12192,N_10438);
nand U16256 (N_16256,N_14348,N_14720);
or U16257 (N_16257,N_11123,N_14064);
or U16258 (N_16258,N_11228,N_11541);
and U16259 (N_16259,N_13829,N_14513);
nand U16260 (N_16260,N_11819,N_11879);
and U16261 (N_16261,N_13698,N_10611);
xor U16262 (N_16262,N_10667,N_13676);
xnor U16263 (N_16263,N_13630,N_13654);
nor U16264 (N_16264,N_10329,N_12276);
nor U16265 (N_16265,N_12723,N_12401);
or U16266 (N_16266,N_10949,N_12393);
and U16267 (N_16267,N_10280,N_14734);
or U16268 (N_16268,N_14216,N_10045);
or U16269 (N_16269,N_11800,N_11177);
nor U16270 (N_16270,N_10158,N_13152);
xnor U16271 (N_16271,N_10125,N_11313);
or U16272 (N_16272,N_12390,N_11468);
nand U16273 (N_16273,N_12014,N_11270);
nand U16274 (N_16274,N_12550,N_10755);
xor U16275 (N_16275,N_11306,N_10322);
and U16276 (N_16276,N_11420,N_10939);
nor U16277 (N_16277,N_14489,N_14729);
and U16278 (N_16278,N_11268,N_11875);
nand U16279 (N_16279,N_10850,N_11110);
xnor U16280 (N_16280,N_14290,N_13440);
or U16281 (N_16281,N_14337,N_14845);
nor U16282 (N_16282,N_12683,N_12204);
or U16283 (N_16283,N_10778,N_12615);
or U16284 (N_16284,N_10763,N_10028);
and U16285 (N_16285,N_12125,N_14021);
nand U16286 (N_16286,N_13935,N_10059);
nor U16287 (N_16287,N_11979,N_11458);
and U16288 (N_16288,N_11222,N_11874);
nor U16289 (N_16289,N_12964,N_12070);
nor U16290 (N_16290,N_14240,N_12519);
xnor U16291 (N_16291,N_10859,N_14922);
and U16292 (N_16292,N_11796,N_12848);
or U16293 (N_16293,N_13494,N_14546);
or U16294 (N_16294,N_10766,N_13715);
or U16295 (N_16295,N_13976,N_12416);
and U16296 (N_16296,N_13349,N_10765);
nor U16297 (N_16297,N_10100,N_14767);
xnor U16298 (N_16298,N_13418,N_10263);
xor U16299 (N_16299,N_14759,N_11025);
or U16300 (N_16300,N_12943,N_14005);
nor U16301 (N_16301,N_11365,N_14185);
nor U16302 (N_16302,N_12586,N_13538);
and U16303 (N_16303,N_11852,N_13836);
and U16304 (N_16304,N_13155,N_11234);
or U16305 (N_16305,N_13575,N_11814);
xor U16306 (N_16306,N_11299,N_13472);
and U16307 (N_16307,N_12213,N_12263);
xnor U16308 (N_16308,N_13905,N_14617);
or U16309 (N_16309,N_14852,N_12846);
xnor U16310 (N_16310,N_10186,N_11069);
or U16311 (N_16311,N_11820,N_11570);
xor U16312 (N_16312,N_12637,N_11088);
and U16313 (N_16313,N_11965,N_14067);
and U16314 (N_16314,N_14981,N_12786);
or U16315 (N_16315,N_14790,N_11017);
nor U16316 (N_16316,N_14586,N_13832);
nand U16317 (N_16317,N_11114,N_14616);
xor U16318 (N_16318,N_10931,N_10130);
or U16319 (N_16319,N_10555,N_14526);
or U16320 (N_16320,N_10454,N_14223);
and U16321 (N_16321,N_13220,N_14933);
or U16322 (N_16322,N_13706,N_11950);
nor U16323 (N_16323,N_14684,N_14459);
or U16324 (N_16324,N_13139,N_12532);
nand U16325 (N_16325,N_10658,N_10260);
and U16326 (N_16326,N_12813,N_12278);
nand U16327 (N_16327,N_12941,N_13807);
and U16328 (N_16328,N_13024,N_12528);
nand U16329 (N_16329,N_10020,N_10896);
nor U16330 (N_16330,N_12551,N_10938);
and U16331 (N_16331,N_10736,N_14260);
xor U16332 (N_16332,N_12432,N_13394);
nand U16333 (N_16333,N_14356,N_11953);
xnor U16334 (N_16334,N_12782,N_13198);
nor U16335 (N_16335,N_10791,N_10760);
nand U16336 (N_16336,N_14515,N_14020);
nand U16337 (N_16337,N_11185,N_11287);
or U16338 (N_16338,N_12596,N_14621);
or U16339 (N_16339,N_10272,N_10832);
and U16340 (N_16340,N_10413,N_11566);
or U16341 (N_16341,N_14029,N_10140);
and U16342 (N_16342,N_13579,N_14642);
or U16343 (N_16343,N_10118,N_13182);
nand U16344 (N_16344,N_12101,N_11314);
nor U16345 (N_16345,N_12527,N_14801);
nand U16346 (N_16346,N_14848,N_10715);
and U16347 (N_16347,N_14367,N_12644);
nand U16348 (N_16348,N_11676,N_12105);
or U16349 (N_16349,N_10284,N_14140);
and U16350 (N_16350,N_14436,N_11304);
or U16351 (N_16351,N_11099,N_13216);
or U16352 (N_16352,N_10097,N_12164);
nor U16353 (N_16353,N_10075,N_11715);
nor U16354 (N_16354,N_13974,N_13411);
and U16355 (N_16355,N_11108,N_13327);
or U16356 (N_16356,N_13683,N_12706);
or U16357 (N_16357,N_10249,N_13846);
nor U16358 (N_16358,N_14854,N_10539);
nor U16359 (N_16359,N_14611,N_14822);
nor U16360 (N_16360,N_10572,N_10799);
and U16361 (N_16361,N_11909,N_10813);
nand U16362 (N_16362,N_11532,N_10053);
nand U16363 (N_16363,N_11116,N_13230);
nand U16364 (N_16364,N_12562,N_10426);
nand U16365 (N_16365,N_11488,N_10147);
and U16366 (N_16366,N_10138,N_12389);
nand U16367 (N_16367,N_14193,N_10400);
or U16368 (N_16368,N_10486,N_14355);
and U16369 (N_16369,N_12468,N_13168);
and U16370 (N_16370,N_13961,N_12433);
nand U16371 (N_16371,N_12293,N_11281);
nor U16372 (N_16372,N_14692,N_10679);
nand U16373 (N_16373,N_11911,N_14529);
or U16374 (N_16374,N_11832,N_13511);
and U16375 (N_16375,N_12148,N_11353);
nor U16376 (N_16376,N_14211,N_10048);
nand U16377 (N_16377,N_11511,N_13548);
or U16378 (N_16378,N_11703,N_11051);
xor U16379 (N_16379,N_10083,N_13015);
or U16380 (N_16380,N_14089,N_14346);
xnor U16381 (N_16381,N_14492,N_11538);
nor U16382 (N_16382,N_11214,N_11697);
xor U16383 (N_16383,N_12911,N_13287);
xnor U16384 (N_16384,N_11631,N_10834);
xor U16385 (N_16385,N_10797,N_11614);
nand U16386 (N_16386,N_14911,N_13083);
or U16387 (N_16387,N_14979,N_12091);
or U16388 (N_16388,N_14556,N_10117);
or U16389 (N_16389,N_12837,N_13926);
nand U16390 (N_16390,N_11132,N_12552);
and U16391 (N_16391,N_11917,N_10480);
and U16392 (N_16392,N_14237,N_13743);
and U16393 (N_16393,N_12617,N_11344);
xnor U16394 (N_16394,N_14417,N_12830);
nor U16395 (N_16395,N_10371,N_10001);
nor U16396 (N_16396,N_11526,N_10882);
xnor U16397 (N_16397,N_10719,N_11784);
xor U16398 (N_16398,N_13977,N_11448);
and U16399 (N_16399,N_14120,N_11842);
or U16400 (N_16400,N_13592,N_11507);
nor U16401 (N_16401,N_12282,N_11065);
xor U16402 (N_16402,N_10226,N_10885);
xor U16403 (N_16403,N_11351,N_12429);
nor U16404 (N_16404,N_10144,N_13309);
nand U16405 (N_16405,N_13571,N_12844);
and U16406 (N_16406,N_14512,N_10619);
nand U16407 (N_16407,N_12328,N_10565);
nor U16408 (N_16408,N_12482,N_13344);
xor U16409 (N_16409,N_10856,N_13439);
nor U16410 (N_16410,N_11848,N_14423);
or U16411 (N_16411,N_10049,N_12992);
or U16412 (N_16412,N_10978,N_14462);
or U16413 (N_16413,N_12471,N_14521);
nor U16414 (N_16414,N_10094,N_13432);
xnor U16415 (N_16415,N_14738,N_11671);
and U16416 (N_16416,N_10414,N_11612);
xnor U16417 (N_16417,N_14983,N_11664);
and U16418 (N_16418,N_11402,N_12597);
xnor U16419 (N_16419,N_13357,N_10728);
or U16420 (N_16420,N_13674,N_13022);
xor U16421 (N_16421,N_12583,N_11539);
or U16422 (N_16422,N_10492,N_14711);
and U16423 (N_16423,N_12777,N_12178);
xor U16424 (N_16424,N_14049,N_14686);
nand U16425 (N_16425,N_13649,N_12627);
or U16426 (N_16426,N_13226,N_13749);
nand U16427 (N_16427,N_11885,N_10213);
xnor U16428 (N_16428,N_13454,N_12613);
nor U16429 (N_16429,N_12138,N_11397);
nand U16430 (N_16430,N_11447,N_14082);
and U16431 (N_16431,N_11760,N_11831);
and U16432 (N_16432,N_14289,N_12219);
nand U16433 (N_16433,N_12909,N_11524);
nor U16434 (N_16434,N_11767,N_14765);
nor U16435 (N_16435,N_13171,N_10503);
nor U16436 (N_16436,N_13998,N_10235);
nand U16437 (N_16437,N_12341,N_11692);
and U16438 (N_16438,N_10318,N_14369);
or U16439 (N_16439,N_13364,N_11027);
xnor U16440 (N_16440,N_10056,N_13326);
nand U16441 (N_16441,N_12318,N_14353);
nor U16442 (N_16442,N_10742,N_12004);
nor U16443 (N_16443,N_14932,N_10838);
and U16444 (N_16444,N_13617,N_12461);
or U16445 (N_16445,N_11449,N_11141);
xor U16446 (N_16446,N_10333,N_10545);
xor U16447 (N_16447,N_11073,N_11622);
xor U16448 (N_16448,N_14663,N_12332);
xor U16449 (N_16449,N_14266,N_13041);
xnor U16450 (N_16450,N_11309,N_12273);
nor U16451 (N_16451,N_13455,N_14293);
nand U16452 (N_16452,N_12214,N_10292);
and U16453 (N_16453,N_12379,N_11334);
nand U16454 (N_16454,N_10258,N_12480);
nor U16455 (N_16455,N_10809,N_11107);
nor U16456 (N_16456,N_13020,N_13862);
or U16457 (N_16457,N_13483,N_13703);
nand U16458 (N_16458,N_11165,N_12095);
nor U16459 (N_16459,N_11646,N_12757);
nand U16460 (N_16460,N_14070,N_12741);
nor U16461 (N_16461,N_13036,N_12854);
or U16462 (N_16462,N_11951,N_11647);
and U16463 (N_16463,N_10211,N_10120);
and U16464 (N_16464,N_11986,N_11291);
nand U16465 (N_16465,N_10411,N_14408);
or U16466 (N_16466,N_14080,N_12835);
nor U16467 (N_16467,N_14376,N_13009);
and U16468 (N_16468,N_14107,N_14441);
nor U16469 (N_16469,N_14600,N_11330);
nor U16470 (N_16470,N_12466,N_12092);
and U16471 (N_16471,N_12234,N_13895);
and U16472 (N_16472,N_12507,N_11190);
nor U16473 (N_16473,N_14130,N_11549);
nand U16474 (N_16474,N_12975,N_10824);
nand U16475 (N_16475,N_13008,N_10511);
nor U16476 (N_16476,N_14202,N_14559);
nor U16477 (N_16477,N_10892,N_11425);
nor U16478 (N_16478,N_11821,N_12887);
nor U16479 (N_16479,N_12334,N_11021);
nand U16480 (N_16480,N_12236,N_14019);
and U16481 (N_16481,N_13348,N_12918);
or U16482 (N_16482,N_11645,N_10975);
nor U16483 (N_16483,N_10725,N_10418);
nand U16484 (N_16484,N_14810,N_11608);
xor U16485 (N_16485,N_14517,N_11118);
nand U16486 (N_16486,N_14967,N_11356);
and U16487 (N_16487,N_14161,N_14414);
or U16488 (N_16488,N_14569,N_12156);
and U16489 (N_16489,N_14464,N_11417);
nor U16490 (N_16490,N_12890,N_13316);
or U16491 (N_16491,N_14827,N_13560);
nand U16492 (N_16492,N_11961,N_14207);
and U16493 (N_16493,N_11543,N_14925);
or U16494 (N_16494,N_13545,N_10972);
nand U16495 (N_16495,N_13210,N_10209);
and U16496 (N_16496,N_14053,N_10751);
or U16497 (N_16497,N_14873,N_13665);
xnor U16498 (N_16498,N_12928,N_13707);
or U16499 (N_16499,N_11467,N_13877);
xor U16500 (N_16500,N_11923,N_12508);
nand U16501 (N_16501,N_14433,N_10415);
and U16502 (N_16502,N_13099,N_12274);
nor U16503 (N_16503,N_13745,N_12881);
or U16504 (N_16504,N_14803,N_14887);
or U16505 (N_16505,N_11245,N_12354);
xor U16506 (N_16506,N_11261,N_13109);
and U16507 (N_16507,N_13196,N_14870);
and U16508 (N_16508,N_14204,N_10320);
nor U16509 (N_16509,N_10577,N_12927);
nor U16510 (N_16510,N_12402,N_10829);
xnor U16511 (N_16511,N_10758,N_10497);
xor U16512 (N_16512,N_13527,N_13387);
nand U16513 (N_16513,N_13670,N_10370);
nor U16514 (N_16514,N_13492,N_14194);
or U16515 (N_16515,N_11987,N_14914);
and U16516 (N_16516,N_13187,N_12764);
xor U16517 (N_16517,N_10916,N_13574);
nor U16518 (N_16518,N_11778,N_12646);
xnor U16519 (N_16519,N_10228,N_14116);
xnor U16520 (N_16520,N_14647,N_10417);
and U16521 (N_16521,N_13551,N_11200);
or U16522 (N_16522,N_14796,N_10081);
and U16523 (N_16523,N_11873,N_13557);
nand U16524 (N_16524,N_10435,N_10065);
xnor U16525 (N_16525,N_10253,N_14090);
xnor U16526 (N_16526,N_11576,N_14957);
or U16527 (N_16527,N_10878,N_13265);
and U16528 (N_16528,N_11552,N_14876);
xor U16529 (N_16529,N_11838,N_14772);
xor U16530 (N_16530,N_10737,N_12684);
and U16531 (N_16531,N_13066,N_13873);
nand U16532 (N_16532,N_13268,N_10767);
nor U16533 (N_16533,N_12072,N_10493);
or U16534 (N_16534,N_11809,N_11865);
xnor U16535 (N_16535,N_13610,N_10680);
nand U16536 (N_16536,N_10893,N_10357);
or U16537 (N_16537,N_10559,N_11782);
nor U16538 (N_16538,N_11652,N_13056);
and U16539 (N_16539,N_13376,N_14281);
nand U16540 (N_16540,N_13480,N_11728);
xor U16541 (N_16541,N_14397,N_12028);
xor U16542 (N_16542,N_10701,N_13889);
and U16543 (N_16543,N_12408,N_12118);
nor U16544 (N_16544,N_14184,N_11182);
and U16545 (N_16545,N_10474,N_12997);
nand U16546 (N_16546,N_13121,N_13060);
nand U16547 (N_16547,N_14746,N_12867);
or U16548 (N_16548,N_10223,N_14843);
nor U16549 (N_16549,N_10746,N_11001);
nor U16550 (N_16550,N_13295,N_14267);
and U16551 (N_16551,N_11970,N_10394);
nor U16552 (N_16552,N_13705,N_10317);
nor U16553 (N_16553,N_11493,N_10376);
and U16554 (N_16554,N_10231,N_13337);
and U16555 (N_16555,N_14449,N_11421);
nor U16556 (N_16556,N_13278,N_14316);
and U16557 (N_16557,N_14045,N_10491);
or U16558 (N_16558,N_10462,N_11387);
and U16559 (N_16559,N_13114,N_10222);
xnor U16560 (N_16560,N_13755,N_11604);
and U16561 (N_16561,N_13102,N_10206);
nand U16562 (N_16562,N_12834,N_13339);
or U16563 (N_16563,N_12494,N_11993);
or U16564 (N_16564,N_14797,N_11438);
nand U16565 (N_16565,N_12982,N_12719);
xor U16566 (N_16566,N_12087,N_14864);
nor U16567 (N_16567,N_10290,N_10788);
and U16568 (N_16568,N_14175,N_14188);
and U16569 (N_16569,N_14063,N_10759);
nand U16570 (N_16570,N_14378,N_12235);
and U16571 (N_16571,N_14954,N_10452);
xnor U16572 (N_16572,N_13857,N_11930);
nor U16573 (N_16573,N_10543,N_13688);
xnor U16574 (N_16574,N_13661,N_13273);
and U16575 (N_16575,N_10900,N_10656);
nand U16576 (N_16576,N_14455,N_11574);
xor U16577 (N_16577,N_14573,N_10828);
xor U16578 (N_16578,N_11266,N_10085);
xnor U16579 (N_16579,N_11286,N_11744);
nand U16580 (N_16580,N_14800,N_13126);
nor U16581 (N_16581,N_13032,N_12384);
or U16582 (N_16582,N_14186,N_12738);
and U16583 (N_16583,N_13843,N_11354);
nand U16584 (N_16584,N_13803,N_12577);
nand U16585 (N_16585,N_14215,N_12685);
nor U16586 (N_16586,N_12462,N_14177);
and U16587 (N_16587,N_14832,N_10416);
and U16588 (N_16588,N_13173,N_13947);
nor U16589 (N_16589,N_14571,N_13910);
and U16590 (N_16590,N_10177,N_11350);
xor U16591 (N_16591,N_13621,N_10282);
and U16592 (N_16592,N_14544,N_11661);
nor U16593 (N_16593,N_13611,N_14507);
nand U16594 (N_16594,N_11273,N_12812);
nor U16595 (N_16595,N_13071,N_11888);
nor U16596 (N_16596,N_14754,N_11076);
nor U16597 (N_16597,N_11521,N_10386);
nand U16598 (N_16598,N_12124,N_10626);
or U16599 (N_16599,N_10864,N_12515);
nand U16600 (N_16600,N_12323,N_13561);
or U16601 (N_16601,N_11669,N_11860);
xnor U16602 (N_16602,N_12622,N_11594);
nor U16603 (N_16603,N_10482,N_13596);
nor U16604 (N_16604,N_11231,N_13257);
and U16605 (N_16605,N_11362,N_10724);
xor U16606 (N_16606,N_13235,N_10541);
xnor U16607 (N_16607,N_14251,N_13433);
nand U16608 (N_16608,N_13854,N_14795);
xnor U16609 (N_16609,N_12582,N_12872);
nand U16610 (N_16610,N_11948,N_13524);
nor U16611 (N_16611,N_14749,N_11277);
nand U16612 (N_16612,N_11817,N_11282);
nor U16613 (N_16613,N_13482,N_13075);
nor U16614 (N_16614,N_11251,N_12373);
or U16615 (N_16615,N_13072,N_11880);
xnor U16616 (N_16616,N_11866,N_10143);
nor U16617 (N_16617,N_14629,N_14653);
xor U16618 (N_16618,N_11696,N_14428);
or U16619 (N_16619,N_10487,N_12336);
and U16620 (N_16620,N_11146,N_13188);
nand U16621 (N_16621,N_13708,N_10665);
nand U16622 (N_16622,N_12792,N_12987);
nand U16623 (N_16623,N_14074,N_14212);
nand U16624 (N_16624,N_14545,N_13673);
nand U16625 (N_16625,N_11342,N_13430);
nor U16626 (N_16626,N_13684,N_13458);
and U16627 (N_16627,N_11066,N_13512);
and U16628 (N_16628,N_12205,N_13093);
or U16629 (N_16629,N_11903,N_14110);
nand U16630 (N_16630,N_12636,N_12063);
and U16631 (N_16631,N_10988,N_11328);
and U16632 (N_16632,N_14518,N_10868);
or U16633 (N_16633,N_13842,N_10054);
and U16634 (N_16634,N_14758,N_10332);
or U16635 (N_16635,N_13820,N_13013);
nor U16636 (N_16636,N_14643,N_14461);
xnor U16637 (N_16637,N_13186,N_11896);
nand U16638 (N_16638,N_13774,N_14971);
nor U16639 (N_16639,N_13937,N_10210);
nor U16640 (N_16640,N_10061,N_13896);
nand U16641 (N_16641,N_11024,N_11573);
and U16642 (N_16642,N_12767,N_10535);
nor U16643 (N_16643,N_11606,N_10669);
nand U16644 (N_16644,N_13909,N_10549);
and U16645 (N_16645,N_12419,N_11575);
xnor U16646 (N_16646,N_11766,N_10865);
or U16647 (N_16647,N_12967,N_10699);
nor U16648 (N_16648,N_11824,N_11335);
nand U16649 (N_16649,N_14519,N_10233);
and U16650 (N_16650,N_14739,N_14233);
or U16651 (N_16651,N_10655,N_14834);
or U16652 (N_16652,N_13338,N_13934);
xnor U16653 (N_16653,N_13234,N_12539);
xor U16654 (N_16654,N_14760,N_13249);
or U16655 (N_16655,N_12795,N_11673);
and U16656 (N_16656,N_14978,N_11954);
and U16657 (N_16657,N_12857,N_12747);
and U16658 (N_16658,N_13042,N_13927);
xor U16659 (N_16659,N_14357,N_11674);
and U16660 (N_16660,N_12457,N_10811);
nor U16661 (N_16661,N_11340,N_13772);
nor U16662 (N_16662,N_11799,N_13746);
nand U16663 (N_16663,N_12773,N_14025);
xnor U16664 (N_16664,N_13329,N_11151);
and U16665 (N_16665,N_11326,N_13853);
nor U16666 (N_16666,N_14314,N_10309);
nor U16667 (N_16667,N_13901,N_12363);
nor U16668 (N_16668,N_13145,N_11035);
xor U16669 (N_16669,N_12153,N_11658);
nand U16670 (N_16670,N_14027,N_10453);
or U16671 (N_16671,N_11105,N_12825);
and U16672 (N_16672,N_13131,N_10707);
and U16673 (N_16673,N_11236,N_13747);
xor U16674 (N_16674,N_10191,N_12167);
xor U16675 (N_16675,N_11367,N_10917);
and U16676 (N_16676,N_12991,N_14374);
or U16677 (N_16677,N_13550,N_12960);
nand U16678 (N_16678,N_14547,N_14968);
nor U16679 (N_16679,N_10225,N_12971);
or U16680 (N_16680,N_14704,N_10285);
and U16681 (N_16681,N_10405,N_10800);
or U16682 (N_16682,N_11115,N_12573);
nand U16683 (N_16683,N_10339,N_13468);
xnor U16684 (N_16684,N_13361,N_10456);
and U16685 (N_16685,N_14505,N_10672);
or U16686 (N_16686,N_10671,N_14793);
nor U16687 (N_16687,N_14991,N_12033);
nor U16688 (N_16688,N_14057,N_12561);
or U16689 (N_16689,N_12246,N_13222);
and U16690 (N_16690,N_12915,N_14456);
and U16691 (N_16691,N_13987,N_12096);
nor U16692 (N_16692,N_13626,N_10174);
and U16693 (N_16693,N_13190,N_13892);
and U16694 (N_16694,N_11748,N_11301);
or U16695 (N_16695,N_14694,N_11075);
nor U16696 (N_16696,N_12417,N_12649);
xor U16697 (N_16697,N_13095,N_13660);
and U16698 (N_16698,N_13336,N_14480);
nor U16699 (N_16699,N_11053,N_14210);
xor U16700 (N_16700,N_13908,N_13595);
and U16701 (N_16701,N_12423,N_13967);
xnor U16702 (N_16702,N_12069,N_14479);
or U16703 (N_16703,N_14446,N_13734);
nand U16704 (N_16704,N_14043,N_11089);
nand U16705 (N_16705,N_14806,N_11565);
nor U16706 (N_16706,N_13591,N_13711);
and U16707 (N_16707,N_11276,N_10981);
nand U16708 (N_16708,N_11964,N_14939);
nand U16709 (N_16709,N_10123,N_13522);
and U16710 (N_16710,N_14716,N_13167);
nor U16711 (N_16711,N_10845,N_13427);
and U16712 (N_16712,N_13038,N_12718);
nor U16713 (N_16713,N_10429,N_11450);
and U16714 (N_16714,N_14218,N_12110);
nor U16715 (N_16715,N_13946,N_11710);
nand U16716 (N_16716,N_12643,N_11219);
nor U16717 (N_16717,N_10703,N_12065);
nand U16718 (N_16718,N_12074,N_11846);
nand U16719 (N_16719,N_11125,N_14657);
and U16720 (N_16720,N_14360,N_10375);
and U16721 (N_16721,N_10358,N_11087);
nor U16722 (N_16722,N_11086,N_13833);
nor U16723 (N_16723,N_12399,N_11319);
or U16724 (N_16724,N_14221,N_11083);
and U16725 (N_16725,N_10933,N_11427);
nand U16726 (N_16726,N_10307,N_10170);
xnor U16727 (N_16727,N_13296,N_11680);
nor U16728 (N_16728,N_10239,N_10731);
xor U16729 (N_16729,N_10690,N_11931);
nor U16730 (N_16730,N_11046,N_14608);
and U16731 (N_16731,N_11347,N_10477);
nand U16732 (N_16732,N_13767,N_14849);
or U16733 (N_16733,N_10676,N_14320);
and U16734 (N_16734,N_12001,N_10971);
and U16735 (N_16735,N_12933,N_13448);
xor U16736 (N_16736,N_11482,N_11329);
xor U16737 (N_16737,N_11952,N_13699);
nor U16738 (N_16738,N_12102,N_13840);
or U16739 (N_16739,N_13850,N_12183);
xor U16740 (N_16740,N_14842,N_14165);
xor U16741 (N_16741,N_13593,N_14525);
nor U16742 (N_16742,N_10310,N_10461);
nand U16743 (N_16743,N_14784,N_12632);
nor U16744 (N_16744,N_12629,N_13581);
nand U16745 (N_16745,N_13818,N_12469);
nor U16746 (N_16746,N_13847,N_11134);
xor U16747 (N_16747,N_13225,N_14732);
nand U16748 (N_16748,N_14430,N_11331);
and U16749 (N_16749,N_12351,N_11348);
and U16750 (N_16750,N_12197,N_11701);
nor U16751 (N_16751,N_10675,N_12745);
or U16752 (N_16752,N_11630,N_10155);
and U16753 (N_16753,N_11518,N_13023);
xnor U16754 (N_16754,N_10651,N_11801);
and U16755 (N_16755,N_12030,N_10087);
or U16756 (N_16756,N_13113,N_13153);
xnor U16757 (N_16757,N_13753,N_13962);
or U16758 (N_16758,N_13159,N_14033);
xor U16759 (N_16759,N_11803,N_13719);
nor U16760 (N_16760,N_11792,N_12614);
nand U16761 (N_16761,N_14527,N_13679);
xor U16762 (N_16762,N_14730,N_10441);
or U16763 (N_16763,N_12858,N_11363);
nor U16764 (N_16764,N_10982,N_13939);
or U16765 (N_16765,N_10881,N_12158);
nor U16766 (N_16766,N_12244,N_14048);
or U16767 (N_16767,N_13040,N_13001);
or U16768 (N_16768,N_12141,N_12599);
or U16769 (N_16769,N_11098,N_10145);
or U16770 (N_16770,N_12916,N_12672);
or U16771 (N_16771,N_10940,N_13125);
nand U16772 (N_16772,N_13500,N_10244);
or U16773 (N_16773,N_14610,N_11191);
or U16774 (N_16774,N_12142,N_11700);
nand U16775 (N_16775,N_14745,N_13509);
nand U16776 (N_16776,N_10353,N_11246);
or U16777 (N_16777,N_10536,N_11143);
and U16778 (N_16778,N_13633,N_13034);
xnor U16779 (N_16779,N_11249,N_12226);
or U16780 (N_16780,N_12259,N_14841);
nor U16781 (N_16781,N_14166,N_10935);
xor U16782 (N_16782,N_12324,N_12047);
nor U16783 (N_16783,N_14283,N_14561);
or U16784 (N_16784,N_12413,N_10102);
nand U16785 (N_16785,N_12954,N_12610);
nor U16786 (N_16786,N_10238,N_13985);
nand U16787 (N_16787,N_14026,N_12093);
nor U16788 (N_16788,N_12049,N_11771);
nand U16789 (N_16789,N_11216,N_12630);
and U16790 (N_16790,N_10876,N_11149);
xor U16791 (N_16791,N_10277,N_14974);
nor U16792 (N_16792,N_11580,N_12127);
nand U16793 (N_16793,N_12720,N_11718);
nor U16794 (N_16794,N_12056,N_13822);
nand U16795 (N_16795,N_14733,N_13463);
or U16796 (N_16796,N_14023,N_10599);
nor U16797 (N_16797,N_11757,N_13111);
and U16798 (N_16798,N_13519,N_13759);
or U16799 (N_16799,N_14323,N_11857);
xnor U16800 (N_16800,N_13694,N_11626);
xnor U16801 (N_16801,N_12998,N_13588);
nand U16802 (N_16802,N_13475,N_13804);
and U16803 (N_16803,N_12038,N_10520);
and U16804 (N_16804,N_13828,N_12031);
and U16805 (N_16805,N_14945,N_12185);
and U16806 (N_16806,N_11494,N_13380);
nor U16807 (N_16807,N_14176,N_13108);
nor U16808 (N_16808,N_13821,N_12849);
nand U16809 (N_16809,N_10327,N_10514);
and U16810 (N_16810,N_12533,N_10455);
nor U16811 (N_16811,N_12658,N_11265);
nor U16812 (N_16812,N_14666,N_11726);
and U16813 (N_16813,N_11167,N_10795);
or U16814 (N_16814,N_10104,N_12591);
or U16815 (N_16815,N_10276,N_10344);
xor U16816 (N_16816,N_13903,N_14696);
nand U16817 (N_16817,N_14807,N_10890);
or U16818 (N_16818,N_12463,N_13875);
nor U16819 (N_16819,N_14595,N_12465);
nor U16820 (N_16820,N_12104,N_12241);
and U16821 (N_16821,N_14354,N_14139);
xor U16822 (N_16822,N_10036,N_12626);
or U16823 (N_16823,N_12357,N_10550);
or U16824 (N_16824,N_10401,N_11153);
or U16825 (N_16825,N_14675,N_12088);
and U16826 (N_16826,N_11610,N_11826);
and U16827 (N_16827,N_10425,N_14934);
or U16828 (N_16828,N_14147,N_12179);
xor U16829 (N_16829,N_13542,N_10163);
or U16830 (N_16830,N_12566,N_14839);
nor U16831 (N_16831,N_11756,N_11795);
or U16832 (N_16832,N_14467,N_10255);
nand U16833 (N_16833,N_13495,N_11385);
nor U16834 (N_16834,N_12793,N_10908);
nor U16835 (N_16835,N_11201,N_12733);
nand U16836 (N_16836,N_13491,N_14757);
nor U16837 (N_16837,N_12930,N_10720);
nand U16838 (N_16838,N_12238,N_12579);
nor U16839 (N_16839,N_13990,N_12266);
xor U16840 (N_16840,N_14751,N_11416);
xor U16841 (N_16841,N_10831,N_10528);
nand U16842 (N_16842,N_14396,N_12500);
xor U16843 (N_16843,N_13091,N_13855);
or U16844 (N_16844,N_13039,N_13399);
or U16845 (N_16845,N_13541,N_14878);
or U16846 (N_16846,N_12189,N_14422);
and U16847 (N_16847,N_11033,N_14516);
nor U16848 (N_16848,N_14183,N_11187);
nor U16849 (N_16849,N_11670,N_10124);
nand U16850 (N_16850,N_11435,N_12166);
and U16851 (N_16851,N_13332,N_11459);
and U16852 (N_16852,N_14419,N_12481);
xnor U16853 (N_16853,N_12512,N_10999);
xnor U16854 (N_16854,N_10184,N_12444);
nand U16855 (N_16855,N_10030,N_12727);
or U16856 (N_16856,N_10537,N_10062);
xnor U16857 (N_16857,N_10443,N_11827);
nor U16858 (N_16858,N_12428,N_13205);
and U16859 (N_16859,N_14387,N_12382);
nor U16860 (N_16860,N_10945,N_10696);
xnor U16861 (N_16861,N_10289,N_14349);
nand U16862 (N_16862,N_13533,N_13107);
nand U16863 (N_16863,N_14671,N_10428);
xor U16864 (N_16864,N_10644,N_10103);
nand U16865 (N_16865,N_14587,N_12233);
nand U16866 (N_16866,N_10403,N_13924);
nand U16867 (N_16867,N_13177,N_10627);
nor U16868 (N_16868,N_14306,N_12843);
and U16869 (N_16869,N_10861,N_10021);
nor U16870 (N_16870,N_12280,N_11197);
xor U16871 (N_16871,N_11558,N_12865);
xnor U16872 (N_16872,N_10729,N_12704);
and U16873 (N_16873,N_11721,N_13074);
nor U16874 (N_16874,N_10694,N_14641);
nor U16875 (N_16875,N_10584,N_14912);
nand U16876 (N_16876,N_13208,N_12584);
xnor U16877 (N_16877,N_14536,N_14669);
and U16878 (N_16878,N_14403,N_12308);
nand U16879 (N_16879,N_14691,N_13570);
or U16880 (N_16880,N_14197,N_14451);
nand U16881 (N_16881,N_11465,N_10460);
xnor U16882 (N_16882,N_10295,N_10596);
or U16883 (N_16883,N_12748,N_12888);
xnor U16884 (N_16884,N_10947,N_11560);
or U16885 (N_16885,N_14153,N_14425);
xor U16886 (N_16886,N_12949,N_12325);
and U16887 (N_16887,N_13488,N_12258);
xnor U16888 (N_16888,N_11881,N_10012);
or U16889 (N_16889,N_10954,N_10591);
or U16890 (N_16890,N_10116,N_13400);
and U16891 (N_16891,N_13007,N_10457);
or U16892 (N_16892,N_10920,N_11775);
xor U16893 (N_16893,N_12557,N_12316);
and U16894 (N_16894,N_12035,N_12986);
nor U16895 (N_16895,N_12435,N_12048);
nor U16896 (N_16896,N_13014,N_11280);
nand U16897 (N_16897,N_14747,N_13340);
and U16898 (N_16898,N_12681,N_13949);
xor U16899 (N_16899,N_11519,N_14707);
nor U16900 (N_16900,N_12322,N_14541);
or U16901 (N_16901,N_12973,N_12264);
and U16902 (N_16902,N_10090,N_10236);
and U16903 (N_16903,N_13778,N_10136);
and U16904 (N_16904,N_13148,N_10079);
and U16905 (N_16905,N_11315,N_13864);
nand U16906 (N_16906,N_14652,N_10481);
nor U16907 (N_16907,N_13766,N_13359);
nor U16908 (N_16908,N_14454,N_11607);
xnor U16909 (N_16909,N_11502,N_10775);
xor U16910 (N_16910,N_12907,N_11691);
nand U16911 (N_16911,N_11625,N_11497);
xnor U16912 (N_16912,N_14127,N_12378);
and U16913 (N_16913,N_13732,N_10142);
nor U16914 (N_16914,N_10544,N_11163);
and U16915 (N_16915,N_14821,N_12199);
and U16916 (N_16916,N_12499,N_13775);
or U16917 (N_16917,N_10574,N_12790);
xor U16918 (N_16918,N_12735,N_12002);
nor U16919 (N_16919,N_12117,N_11988);
nor U16920 (N_16920,N_12822,N_14399);
and U16921 (N_16921,N_12541,N_11747);
nand U16922 (N_16922,N_11619,N_10350);
nand U16923 (N_16923,N_12937,N_12952);
and U16924 (N_16924,N_14916,N_11093);
xor U16925 (N_16925,N_13784,N_11457);
or U16926 (N_16926,N_12833,N_13577);
nor U16927 (N_16927,N_13281,N_14091);
xnor U16928 (N_16928,N_13289,N_12808);
xor U16929 (N_16929,N_14191,N_14882);
nor U16930 (N_16930,N_11476,N_14435);
nor U16931 (N_16931,N_12522,N_14564);
nor U16932 (N_16932,N_12734,N_13653);
and U16933 (N_16933,N_11555,N_13419);
or U16934 (N_16934,N_11293,N_10374);
or U16935 (N_16935,N_14071,N_13580);
nand U16936 (N_16936,N_11162,N_13623);
or U16937 (N_16937,N_13237,N_11675);
and U16938 (N_16938,N_14549,N_12606);
and U16939 (N_16939,N_14366,N_11057);
nor U16940 (N_16940,N_14014,N_10328);
xnor U16941 (N_16941,N_12051,N_12885);
nand U16942 (N_16942,N_14501,N_11117);
nand U16943 (N_16943,N_11010,N_10463);
or U16944 (N_16944,N_11845,N_11324);
nand U16945 (N_16945,N_11849,N_10773);
xnor U16946 (N_16946,N_10093,N_10804);
and U16947 (N_16947,N_10135,N_12020);
xor U16948 (N_16948,N_13262,N_10224);
nor U16949 (N_16949,N_10802,N_13037);
nand U16950 (N_16950,N_10007,N_14060);
xnor U16951 (N_16951,N_11074,N_14509);
and U16952 (N_16952,N_12990,N_14943);
nor U16953 (N_16953,N_12707,N_13116);
nor U16954 (N_16954,N_12455,N_12222);
xor U16955 (N_16955,N_14615,N_12496);
and U16956 (N_16956,N_12304,N_10199);
or U16957 (N_16957,N_11188,N_12690);
nor U16958 (N_16958,N_11789,N_11735);
and U16959 (N_16959,N_14956,N_13898);
or U16960 (N_16960,N_10475,N_12397);
nand U16961 (N_16961,N_11522,N_11272);
and U16962 (N_16962,N_12705,N_11422);
or U16963 (N_16963,N_14622,N_13677);
nand U16964 (N_16964,N_14522,N_11528);
nor U16965 (N_16965,N_12342,N_12654);
nor U16966 (N_16966,N_11886,N_11855);
nor U16967 (N_16967,N_14857,N_10953);
xnor U16968 (N_16968,N_12902,N_11446);
xor U16969 (N_16969,N_11003,N_13160);
nor U16970 (N_16970,N_14079,N_12977);
xnor U16971 (N_16971,N_14788,N_11867);
and U16972 (N_16972,N_12710,N_12783);
nor U16973 (N_16973,N_10360,N_13666);
xnor U16974 (N_16974,N_12802,N_14168);
nor U16975 (N_16975,N_11642,N_11414);
and U16976 (N_16976,N_10525,N_12114);
and U16977 (N_16977,N_13936,N_14145);
nand U16978 (N_16978,N_14596,N_12082);
nand U16979 (N_16979,N_11032,N_11785);
nand U16980 (N_16980,N_11804,N_11586);
nor U16981 (N_16981,N_10512,N_14372);
and U16982 (N_16982,N_13565,N_14828);
nand U16983 (N_16983,N_14234,N_13150);
nor U16984 (N_16984,N_12820,N_10006);
xnor U16985 (N_16985,N_13450,N_12669);
nand U16986 (N_16986,N_13426,N_12445);
or U16987 (N_16987,N_11922,N_11962);
nand U16988 (N_16988,N_10697,N_12157);
nor U16989 (N_16989,N_10215,N_10299);
nand U16990 (N_16990,N_14703,N_14965);
nor U16991 (N_16991,N_14024,N_11424);
xnor U16992 (N_16992,N_11976,N_12003);
nor U16993 (N_16993,N_12012,N_14383);
xnor U16994 (N_16994,N_10790,N_14813);
nand U16995 (N_16995,N_13211,N_13870);
or U16996 (N_16996,N_10051,N_12712);
nand U16997 (N_16997,N_13343,N_14490);
nor U16998 (N_16998,N_14158,N_11296);
xor U16999 (N_16999,N_13320,N_12256);
or U17000 (N_17000,N_12040,N_10546);
nor U17001 (N_17001,N_13369,N_14511);
nand U17002 (N_17002,N_13098,N_12414);
or U17003 (N_17003,N_12434,N_10542);
xnor U17004 (N_17004,N_13467,N_13438);
and U17005 (N_17005,N_14658,N_10617);
nor U17006 (N_17006,N_11982,N_13762);
and U17007 (N_17007,N_12771,N_13667);
and U17008 (N_17008,N_11444,N_13352);
and U17009 (N_17009,N_13802,N_13529);
or U17010 (N_17010,N_13814,N_13317);
or U17011 (N_17011,N_10843,N_10932);
xnor U17012 (N_17012,N_14672,N_14644);
or U17013 (N_17013,N_11815,N_14604);
or U17014 (N_17014,N_13497,N_12564);
nor U17015 (N_17015,N_13729,N_14117);
xor U17016 (N_17016,N_14182,N_13724);
xnor U17017 (N_17017,N_14902,N_12988);
and U17018 (N_17018,N_10762,N_12487);
and U17019 (N_17019,N_14054,N_12023);
nor U17020 (N_17020,N_10489,N_12565);
xnor U17021 (N_17021,N_11967,N_13744);
nand U17022 (N_17022,N_14138,N_14773);
nor U17023 (N_17023,N_14102,N_13471);
nor U17024 (N_17024,N_10979,N_10904);
nand U17025 (N_17025,N_13589,N_14311);
or U17026 (N_17026,N_14960,N_11938);
or U17027 (N_17027,N_10632,N_14157);
xnor U17028 (N_17028,N_11741,N_13404);
and U17029 (N_17029,N_14562,N_12758);
nand U17030 (N_17030,N_11366,N_10605);
nand U17031 (N_17031,N_14638,N_12452);
nor U17032 (N_17032,N_10154,N_11925);
nand U17033 (N_17033,N_14891,N_14964);
nor U17034 (N_17034,N_14042,N_10615);
xor U17035 (N_17035,N_10752,N_10554);
xor U17036 (N_17036,N_12060,N_13025);
xnor U17037 (N_17037,N_10987,N_13681);
and U17038 (N_17038,N_13223,N_13407);
or U17039 (N_17039,N_11924,N_11918);
nand U17040 (N_17040,N_10529,N_14985);
or U17041 (N_17041,N_10444,N_10722);
and U17042 (N_17042,N_13785,N_14528);
and U17043 (N_17043,N_10340,N_13735);
xnor U17044 (N_17044,N_10379,N_12850);
and U17045 (N_17045,N_13425,N_14015);
nand U17046 (N_17046,N_14766,N_13612);
or U17047 (N_17047,N_14555,N_10717);
and U17048 (N_17048,N_14112,N_11413);
nand U17049 (N_17049,N_12598,N_10871);
xnor U17050 (N_17050,N_10527,N_12425);
or U17051 (N_17051,N_13436,N_14531);
nand U17052 (N_17052,N_10271,N_14162);
or U17053 (N_17053,N_10351,N_12879);
xor U17054 (N_17054,N_11056,N_11308);
nand U17055 (N_17055,N_11071,N_12939);
nand U17056 (N_17056,N_12042,N_14199);
nor U17057 (N_17057,N_12968,N_12521);
or U17058 (N_17058,N_14208,N_11102);
nand U17059 (N_17059,N_13521,N_10967);
nand U17060 (N_17060,N_12983,N_13403);
nor U17061 (N_17061,N_10713,N_11609);
nand U17062 (N_17062,N_12080,N_13378);
nor U17063 (N_17063,N_14034,N_10852);
nor U17064 (N_17064,N_13219,N_14894);
nand U17065 (N_17065,N_13279,N_10151);
nand U17066 (N_17066,N_11055,N_12760);
xor U17067 (N_17067,N_11651,N_14329);
and U17068 (N_17068,N_12109,N_10743);
xor U17069 (N_17069,N_12372,N_11311);
and U17070 (N_17070,N_12810,N_14249);
and U17071 (N_17071,N_10408,N_14400);
nand U17072 (N_17072,N_11147,N_13360);
and U17073 (N_17073,N_12534,N_12207);
xor U17074 (N_17074,N_14160,N_14625);
nor U17075 (N_17075,N_14783,N_14959);
xor U17076 (N_17076,N_10613,N_11054);
xor U17077 (N_17077,N_11170,N_14877);
or U17078 (N_17078,N_11047,N_14685);
or U17079 (N_17079,N_14626,N_13105);
nor U17080 (N_17080,N_11743,N_13397);
and U17081 (N_17081,N_13718,N_14804);
or U17082 (N_17082,N_12845,N_12057);
nor U17083 (N_17083,N_13687,N_13941);
and U17084 (N_17084,N_14474,N_11844);
or U17085 (N_17085,N_12775,N_11916);
and U17086 (N_17086,N_13311,N_12917);
nor U17087 (N_17087,N_10628,N_13608);
nor U17088 (N_17088,N_13620,N_14213);
nand U17089 (N_17089,N_10261,N_13634);
xor U17090 (N_17090,N_12467,N_13350);
xnor U17091 (N_17091,N_14605,N_14689);
and U17092 (N_17092,N_13543,N_10181);
or U17093 (N_17093,N_14942,N_13243);
nand U17094 (N_17094,N_14245,N_12945);
or U17095 (N_17095,N_12666,N_10241);
nand U17096 (N_17096,N_11407,N_11300);
and U17097 (N_17097,N_13217,N_14973);
or U17098 (N_17098,N_13712,N_10364);
nor U17099 (N_17099,N_10575,N_10606);
and U17100 (N_17100,N_13534,N_13658);
nor U17101 (N_17101,N_10072,N_11371);
nor U17102 (N_17102,N_12524,N_11531);
xor U17103 (N_17103,N_10383,N_10016);
and U17104 (N_17104,N_12797,N_10894);
nor U17105 (N_17105,N_11602,N_12815);
xnor U17106 (N_17106,N_12638,N_11004);
nor U17107 (N_17107,N_12203,N_13972);
nor U17108 (N_17108,N_14152,N_10368);
nand U17109 (N_17109,N_13860,N_12151);
xor U17110 (N_17110,N_11399,N_14073);
nor U17111 (N_17111,N_13298,N_11333);
or U17112 (N_17112,N_12594,N_14087);
nor U17113 (N_17113,N_12868,N_11000);
nand U17114 (N_17114,N_10208,N_14294);
or U17115 (N_17115,N_12855,N_10352);
and U17116 (N_17116,N_11581,N_12488);
or U17117 (N_17117,N_14593,N_11895);
or U17118 (N_17118,N_13773,N_11683);
and U17119 (N_17119,N_13944,N_13585);
and U17120 (N_17120,N_10569,N_13973);
and U17121 (N_17121,N_11415,N_12090);
nand U17122 (N_17122,N_14698,N_12159);
and U17123 (N_17123,N_12130,N_13586);
nor U17124 (N_17124,N_11656,N_10562);
and U17125 (N_17125,N_10687,N_12311);
nor U17126 (N_17126,N_11733,N_10777);
nor U17127 (N_17127,N_12115,N_10553);
and U17128 (N_17128,N_13081,N_14752);
nor U17129 (N_17129,N_12161,N_10905);
nand U17130 (N_17130,N_14591,N_11694);
or U17131 (N_17131,N_12729,N_10870);
or U17132 (N_17132,N_10096,N_10727);
and U17133 (N_17133,N_13319,N_10844);
nor U17134 (N_17134,N_14613,N_11878);
nor U17135 (N_17135,N_14816,N_10169);
xor U17136 (N_17136,N_10853,N_13604);
nor U17137 (N_17137,N_12572,N_14342);
nand U17138 (N_17138,N_14280,N_13085);
nor U17139 (N_17139,N_13933,N_14258);
nand U17140 (N_17140,N_12225,N_12491);
nand U17141 (N_17141,N_13172,N_12663);
or U17142 (N_17142,N_10037,N_13945);
xor U17143 (N_17143,N_14284,N_12866);
xnor U17144 (N_17144,N_10642,N_10000);
nor U17145 (N_17145,N_13704,N_14196);
xor U17146 (N_17146,N_13308,N_14418);
or U17147 (N_17147,N_12285,N_12625);
nor U17148 (N_17148,N_11734,N_12936);
and U17149 (N_17149,N_13396,N_11042);
or U17150 (N_17150,N_12947,N_14108);
xnor U17151 (N_17151,N_10160,N_13462);
xnor U17152 (N_17152,N_10836,N_13183);
xor U17153 (N_17153,N_11998,N_10733);
or U17154 (N_17154,N_13983,N_12044);
or U17155 (N_17155,N_13866,N_13306);
nor U17156 (N_17156,N_14299,N_13645);
nand U17157 (N_17157,N_12374,N_12526);
xnor U17158 (N_17158,N_13053,N_14778);
nand U17159 (N_17159,N_13476,N_14639);
xor U17160 (N_17160,N_11668,N_13096);
nor U17161 (N_17161,N_11195,N_13988);
xnor U17162 (N_17162,N_13445,N_13323);
or U17163 (N_17163,N_10678,N_10485);
and U17164 (N_17164,N_13991,N_14187);
nor U17165 (N_17165,N_10483,N_14128);
nand U17166 (N_17166,N_10926,N_11969);
and U17167 (N_17167,N_14724,N_14059);
nand U17168 (N_17168,N_11135,N_11176);
nor U17169 (N_17169,N_12751,N_11360);
and U17170 (N_17170,N_11891,N_11739);
or U17171 (N_17171,N_14740,N_11171);
nor U17172 (N_17172,N_10668,N_11072);
xor U17173 (N_17173,N_12107,N_12816);
nand U17174 (N_17174,N_10638,N_14984);
nor U17175 (N_17175,N_13124,N_10478);
and U17176 (N_17176,N_11777,N_10721);
xor U17177 (N_17177,N_10149,N_10670);
nand U17178 (N_17178,N_11956,N_14226);
and U17179 (N_17179,N_10024,N_13995);
xnor U17180 (N_17180,N_12709,N_13690);
or U17181 (N_17181,N_12838,N_11383);
xor U17182 (N_17182,N_13764,N_12978);
and U17183 (N_17183,N_13070,N_13601);
xor U17184 (N_17184,N_13886,N_14946);
nor U17185 (N_17185,N_10784,N_11404);
xnor U17186 (N_17186,N_11641,N_14252);
nor U17187 (N_17187,N_11920,N_10448);
xor U17188 (N_17188,N_14982,N_11255);
and U17189 (N_17189,N_11207,N_14495);
nand U17190 (N_17190,N_13837,N_14401);
nand U17191 (N_17191,N_10570,N_12662);
nand U17192 (N_17192,N_12942,N_14892);
nand U17193 (N_17193,N_14328,N_11337);
nand U17194 (N_17194,N_13479,N_11892);
or U17195 (N_17195,N_11787,N_10073);
nor U17196 (N_17196,N_10662,N_13999);
nand U17197 (N_17197,N_14146,N_12343);
xnor U17198 (N_17198,N_14232,N_10347);
or U17199 (N_17199,N_11729,N_13800);
nor U17200 (N_17200,N_11031,N_11428);
nor U17201 (N_17201,N_12032,N_12099);
and U17202 (N_17202,N_12410,N_14743);
nand U17203 (N_17203,N_11738,N_11997);
xor U17204 (N_17204,N_12761,N_11551);
and U17205 (N_17205,N_11754,N_12272);
nor U17206 (N_17206,N_11762,N_10313);
xor U17207 (N_17207,N_11746,N_11592);
nand U17208 (N_17208,N_11101,N_11500);
xor U17209 (N_17209,N_10634,N_10039);
and U17210 (N_17210,N_14665,N_13084);
nor U17211 (N_17211,N_10907,N_11854);
nand U17212 (N_17212,N_10180,N_14265);
or U17213 (N_17213,N_14137,N_11418);
nor U17214 (N_17214,N_11884,N_11764);
nand U17215 (N_17215,N_13290,N_11198);
nor U17216 (N_17216,N_10925,N_10858);
and U17217 (N_17217,N_14222,N_12215);
nor U17218 (N_17218,N_11957,N_14592);
nor U17219 (N_17219,N_12894,N_14304);
or U17220 (N_17220,N_10306,N_14554);
xnor U17221 (N_17221,N_11434,N_12860);
xnor U17222 (N_17222,N_14036,N_12284);
or U17223 (N_17223,N_12008,N_14815);
or U17224 (N_17224,N_13880,N_11678);
or U17225 (N_17225,N_13782,N_14679);
nor U17226 (N_17226,N_13752,N_13302);
and U17227 (N_17227,N_14395,N_12824);
nand U17228 (N_17228,N_13389,N_11180);
or U17229 (N_17229,N_14590,N_11788);
nand U17230 (N_17230,N_12224,N_14361);
xor U17231 (N_17231,N_10919,N_10952);
and U17232 (N_17232,N_12946,N_11926);
nand U17233 (N_17233,N_14244,N_10265);
and U17234 (N_17234,N_11830,N_14278);
and U17235 (N_17235,N_12010,N_10693);
or U17236 (N_17236,N_10190,N_12136);
and U17237 (N_17237,N_14011,N_14923);
xnor U17238 (N_17238,N_12443,N_13594);
xnor U17239 (N_17239,N_13760,N_13224);
or U17240 (N_17240,N_10785,N_12221);
xor U17241 (N_17241,N_10648,N_10026);
or U17242 (N_17242,N_11218,N_11254);
and U17243 (N_17243,N_12172,N_13214);
or U17244 (N_17244,N_13552,N_12108);
nand U17245 (N_17245,N_13282,N_11791);
xnor U17246 (N_17246,N_10793,N_11840);
or U17247 (N_17247,N_13569,N_10027);
nor U17248 (N_17248,N_10046,N_12315);
xor U17249 (N_17249,N_10833,N_13092);
xor U17250 (N_17250,N_13076,N_14910);
and U17251 (N_17251,N_13128,N_12121);
or U17252 (N_17252,N_10580,N_14962);
nand U17253 (N_17253,N_14051,N_12791);
and U17254 (N_17254,N_13971,N_13207);
nor U17255 (N_17255,N_13520,N_14427);
nand U17256 (N_17256,N_10922,N_10335);
and U17257 (N_17257,N_10042,N_11975);
or U17258 (N_17258,N_10645,N_11391);
or U17259 (N_17259,N_14343,N_12736);
or U17260 (N_17260,N_10860,N_14335);
nor U17261 (N_17261,N_13531,N_10983);
nor U17262 (N_17262,N_12545,N_13478);
nor U17263 (N_17263,N_14031,N_10248);
nand U17264 (N_17264,N_12451,N_13606);
or U17265 (N_17265,N_12889,N_10835);
or U17266 (N_17266,N_14840,N_10510);
nand U17267 (N_17267,N_12364,N_14229);
and U17268 (N_17268,N_12525,N_13410);
nand U17269 (N_17269,N_14309,N_13353);
nor U17270 (N_17270,N_11611,N_14645);
nor U17271 (N_17271,N_14050,N_13721);
xnor U17272 (N_17272,N_10099,N_11002);
or U17273 (N_17273,N_14871,N_12245);
nand U17274 (N_17274,N_13657,N_10748);
nand U17275 (N_17275,N_13770,N_13964);
and U17276 (N_17276,N_13291,N_11481);
nor U17277 (N_17277,N_13283,N_14305);
or U17278 (N_17278,N_10764,N_10395);
nand U17279 (N_17279,N_12959,N_13229);
or U17280 (N_17280,N_13254,N_11005);
or U17281 (N_17281,N_13303,N_13643);
or U17282 (N_17282,N_13321,N_10614);
nand U17283 (N_17283,N_10488,N_10022);
nand U17284 (N_17284,N_10818,N_12237);
xnor U17285 (N_17285,N_11921,N_13233);
nor U17286 (N_17286,N_10884,N_11352);
or U17287 (N_17287,N_10630,N_12650);
and U17288 (N_17288,N_12184,N_14833);
nand U17289 (N_17289,N_14862,N_10423);
nor U17290 (N_17290,N_11142,N_12576);
or U17291 (N_17291,N_14083,N_14557);
and U17292 (N_17292,N_10976,N_14865);
nor U17293 (N_17293,N_12634,N_13270);
or U17294 (N_17294,N_12831,N_14172);
nor U17295 (N_17295,N_11431,N_11949);
nand U17296 (N_17296,N_12232,N_12186);
xor U17297 (N_17297,N_12878,N_10753);
and U17298 (N_17298,N_12022,N_11078);
nand U17299 (N_17299,N_14900,N_12546);
nor U17300 (N_17300,N_13547,N_13365);
nor U17301 (N_17301,N_13304,N_13129);
xor U17302 (N_17302,N_10200,N_11839);
nand U17303 (N_17303,N_11373,N_10906);
nor U17304 (N_17304,N_13401,N_13714);
or U17305 (N_17305,N_12053,N_10201);
or U17306 (N_17306,N_13252,N_14114);
xor U17307 (N_17307,N_14121,N_11112);
nor U17308 (N_17308,N_13130,N_13979);
xnor U17309 (N_17309,N_13117,N_12426);
xor U17310 (N_17310,N_11991,N_10060);
or U17311 (N_17311,N_13087,N_14410);
xnor U17312 (N_17312,N_12209,N_12892);
and U17313 (N_17313,N_13331,N_11248);
and U17314 (N_17314,N_10044,N_12103);
and U17315 (N_17315,N_14326,N_14980);
or U17316 (N_17316,N_12514,N_10551);
or U17317 (N_17317,N_14835,N_10314);
xor U17318 (N_17318,N_11044,N_10484);
nor U17319 (N_17319,N_14579,N_14209);
nand U17320 (N_17320,N_10459,N_12633);
nand U17321 (N_17321,N_10361,N_14820);
nand U17322 (N_17322,N_13805,N_11490);
nor U17323 (N_17323,N_11530,N_14098);
and U17324 (N_17324,N_12999,N_14944);
and U17325 (N_17325,N_13737,N_13904);
and U17326 (N_17326,N_14550,N_10684);
nand U17327 (N_17327,N_12478,N_12948);
and U17328 (N_17328,N_14302,N_14619);
and U17329 (N_17329,N_12450,N_14709);
and U17330 (N_17330,N_10997,N_14633);
and U17331 (N_17331,N_10750,N_11899);
and U17332 (N_17332,N_11995,N_14457);
and U17333 (N_17333,N_11634,N_14460);
xor U17334 (N_17334,N_12697,N_12441);
and U17335 (N_17335,N_11209,N_14239);
and U17336 (N_17336,N_10807,N_14630);
nand U17337 (N_17337,N_14331,N_13763);
nand U17338 (N_17338,N_14151,N_12674);
xnor U17339 (N_17339,N_12174,N_14855);
and U17340 (N_17340,N_10992,N_13922);
and U17341 (N_17341,N_11305,N_14867);
nor U17342 (N_17342,N_14004,N_14909);
nor U17343 (N_17343,N_13499,N_12880);
and U17344 (N_17344,N_10660,N_12601);
and U17345 (N_17345,N_13789,N_13052);
or U17346 (N_17346,N_13250,N_11672);
nand U17347 (N_17347,N_13996,N_12770);
xnor U17348 (N_17348,N_11636,N_13027);
or U17349 (N_17349,N_11256,N_10115);
and U17350 (N_17350,N_11893,N_12898);
xnor U17351 (N_17351,N_12294,N_10047);
nor U17352 (N_17352,N_14811,N_11157);
xnor U17353 (N_17353,N_11058,N_13887);
nand U17354 (N_17354,N_10956,N_13605);
nand U17355 (N_17355,N_10631,N_14312);
nor U17356 (N_17356,N_12024,N_12628);
nor U17357 (N_17357,N_12449,N_14668);
nand U17358 (N_17358,N_12756,N_11640);
nand U17359 (N_17359,N_12914,N_11989);
and U17360 (N_17360,N_12595,N_10373);
or U17361 (N_17361,N_14656,N_12671);
or U17362 (N_17362,N_13678,N_12877);
nor U17363 (N_17363,N_14389,N_14570);
and U17364 (N_17364,N_10839,N_14336);
xor U17365 (N_17365,N_14477,N_14552);
and U17366 (N_17366,N_10578,N_11451);
and U17367 (N_17367,N_14012,N_14113);
nor U17368 (N_17368,N_12768,N_11693);
and U17369 (N_17369,N_12007,N_12275);
nor U17370 (N_17370,N_13259,N_12970);
nor U17371 (N_17371,N_14276,N_12502);
and U17372 (N_17372,N_10974,N_11332);
xor U17373 (N_17373,N_10433,N_12687);
nor U17374 (N_17374,N_10607,N_12800);
and U17375 (N_17375,N_12518,N_14532);
nor U17376 (N_17376,N_11378,N_12570);
nor U17377 (N_17377,N_14148,N_12641);
xor U17378 (N_17378,N_13073,N_12901);
or U17379 (N_17379,N_12807,N_14721);
xor U17380 (N_17380,N_12910,N_13286);
or U17381 (N_17381,N_13912,N_10961);
nor U17382 (N_17382,N_14763,N_14347);
xnor U17383 (N_17383,N_13754,N_10776);
and U17384 (N_17384,N_12262,N_10202);
xor U17385 (N_17385,N_11312,N_12925);
nand U17386 (N_17386,N_12765,N_10442);
or U17387 (N_17387,N_11653,N_10359);
or U17388 (N_17388,N_11496,N_14390);
nand U17389 (N_17389,N_10768,N_10689);
and U17390 (N_17390,N_10587,N_13006);
and U17391 (N_17391,N_11811,N_10496);
nand U17392 (N_17392,N_12447,N_12664);
nor U17393 (N_17393,N_14295,N_14499);
nor U17394 (N_17394,N_12405,N_14286);
and U17395 (N_17395,N_11137,N_13741);
xor U17396 (N_17396,N_12503,N_11285);
xnor U17397 (N_17397,N_11755,N_10593);
and U17398 (N_17398,N_12129,N_13251);
nand U17399 (N_17399,N_12418,N_12337);
or U17400 (N_17400,N_14109,N_11380);
nand U17401 (N_17401,N_12079,N_10647);
nor U17402 (N_17402,N_12229,N_12661);
and U17403 (N_17403,N_12287,N_10677);
nor U17404 (N_17404,N_13600,N_11148);
nand U17405 (N_17405,N_11639,N_12842);
nor U17406 (N_17406,N_10579,N_14133);
xor U17407 (N_17407,N_14097,N_12851);
nor U17408 (N_17408,N_10385,N_14632);
nand U17409 (N_17409,N_13514,N_10286);
xor U17410 (N_17410,N_14612,N_12431);
nand U17411 (N_17411,N_10567,N_14737);
or U17412 (N_17412,N_14205,N_11623);
and U17413 (N_17413,N_12523,N_11289);
nor U17414 (N_17414,N_12944,N_11557);
or U17415 (N_17415,N_13632,N_13779);
or U17416 (N_17416,N_12762,N_10179);
and U17417 (N_17417,N_10556,N_11390);
or U17418 (N_17418,N_13963,N_13598);
and U17419 (N_17419,N_10384,N_14497);
xor U17420 (N_17420,N_13228,N_13583);
nand U17421 (N_17421,N_10847,N_12211);
nand U17422 (N_17422,N_11477,N_10446);
and U17423 (N_17423,N_14124,N_11411);
xnor U17424 (N_17424,N_10966,N_10196);
nor U17425 (N_17425,N_14989,N_12818);
and U17426 (N_17426,N_14332,N_14770);
nand U17427 (N_17427,N_14496,N_12261);
xor U17428 (N_17428,N_11323,N_10063);
nor U17429 (N_17429,N_10984,N_10398);
xor U17430 (N_17430,N_12980,N_13422);
or U17431 (N_17431,N_11262,N_12799);
nor U17432 (N_17432,N_12742,N_13164);
xnor U17433 (N_17433,N_13868,N_14750);
nand U17434 (N_17434,N_14768,N_13382);
or U17435 (N_17435,N_11836,N_11536);
or U17436 (N_17436,N_14963,N_12106);
and U17437 (N_17437,N_14225,N_14535);
or U17438 (N_17438,N_13112,N_10846);
or U17439 (N_17439,N_10857,N_11990);
and U17440 (N_17440,N_11039,N_10355);
nor U17441 (N_17441,N_13051,N_13423);
and U17442 (N_17442,N_13730,N_12206);
nor U17443 (N_17443,N_14487,N_12604);
and U17444 (N_17444,N_11178,N_11963);
or U17445 (N_17445,N_12940,N_10105);
nand U17446 (N_17446,N_13769,N_14476);
and U17447 (N_17447,N_14585,N_11711);
or U17448 (N_17448,N_11462,N_12652);
and U17449 (N_17449,N_10869,N_10197);
or U17450 (N_17450,N_10652,N_13916);
nand U17451 (N_17451,N_13651,N_12913);
xor U17452 (N_17452,N_13035,N_13063);
and U17453 (N_17453,N_14440,N_11945);
nor U17454 (N_17454,N_11501,N_10801);
nand U17455 (N_17455,N_13018,N_13342);
or U17456 (N_17456,N_12922,N_14514);
xor U17457 (N_17457,N_10198,N_10509);
or U17458 (N_17458,N_14838,N_13127);
or U17459 (N_17459,N_14381,N_10710);
nand U17460 (N_17460,N_11617,N_13103);
and U17461 (N_17461,N_14504,N_11370);
nor U17462 (N_17462,N_13827,N_13725);
nor U17463 (N_17463,N_12043,N_10854);
or U17464 (N_17464,N_10476,N_14861);
nor U17465 (N_17465,N_14174,N_10624);
xnor U17466 (N_17466,N_13897,N_12302);
xor U17467 (N_17467,N_12575,N_14002);
nand U17468 (N_17468,N_11772,N_13839);
xor U17469 (N_17469,N_10283,N_14714);
or U17470 (N_17470,N_14375,N_14471);
xnor U17471 (N_17471,N_10148,N_14708);
nor U17472 (N_17472,N_10526,N_14242);
xnor U17473 (N_17473,N_13122,N_14081);
xor U17474 (N_17474,N_14791,N_14084);
or U17475 (N_17475,N_12143,N_11589);
nand U17476 (N_17476,N_11376,N_13635);
xnor U17477 (N_17477,N_13412,N_11802);
and U17478 (N_17478,N_10129,N_11510);
xnor U17479 (N_17479,N_12255,N_13097);
xnor U17480 (N_17480,N_12699,N_10273);
or U17481 (N_17481,N_11540,N_13656);
nand U17482 (N_17482,N_11806,N_14929);
nand U17483 (N_17483,N_14478,N_14631);
or U17484 (N_17484,N_12640,N_12957);
or U17485 (N_17485,N_14195,N_11095);
xor U17486 (N_17486,N_13390,N_10929);
nand U17487 (N_17487,N_11992,N_12220);
nand U17488 (N_17488,N_11109,N_14484);
or U17489 (N_17489,N_13848,N_10294);
xor U17490 (N_17490,N_12376,N_10825);
nand U17491 (N_17491,N_13242,N_11346);
and U17492 (N_17492,N_13065,N_10237);
and U17493 (N_17493,N_13696,N_14661);
nor U17494 (N_17494,N_12875,N_12492);
nand U17495 (N_17495,N_10165,N_11864);
and U17496 (N_17496,N_12165,N_13783);
xor U17497 (N_17497,N_12763,N_12966);
and U17498 (N_17498,N_10779,N_13161);
nor U17499 (N_17499,N_12686,N_10504);
nand U17500 (N_17500,N_10157,N_13551);
xnor U17501 (N_17501,N_10405,N_12575);
xor U17502 (N_17502,N_12426,N_12100);
and U17503 (N_17503,N_14939,N_10599);
or U17504 (N_17504,N_13024,N_10156);
nand U17505 (N_17505,N_10293,N_12633);
or U17506 (N_17506,N_14048,N_11123);
or U17507 (N_17507,N_13410,N_11727);
or U17508 (N_17508,N_12282,N_14705);
or U17509 (N_17509,N_11125,N_10148);
xor U17510 (N_17510,N_10513,N_12357);
nand U17511 (N_17511,N_13201,N_14235);
xnor U17512 (N_17512,N_10055,N_12886);
nand U17513 (N_17513,N_12101,N_14646);
and U17514 (N_17514,N_12584,N_11517);
and U17515 (N_17515,N_13934,N_11337);
nor U17516 (N_17516,N_14631,N_13935);
nor U17517 (N_17517,N_12561,N_11358);
or U17518 (N_17518,N_11131,N_10610);
nor U17519 (N_17519,N_14406,N_12092);
nand U17520 (N_17520,N_12192,N_10660);
or U17521 (N_17521,N_14715,N_14749);
xnor U17522 (N_17522,N_13142,N_12764);
nor U17523 (N_17523,N_14481,N_12150);
nor U17524 (N_17524,N_10281,N_11969);
or U17525 (N_17525,N_10704,N_11723);
nor U17526 (N_17526,N_11295,N_12227);
or U17527 (N_17527,N_10539,N_13805);
and U17528 (N_17528,N_12039,N_13871);
xor U17529 (N_17529,N_11015,N_12896);
xnor U17530 (N_17530,N_10453,N_14283);
nand U17531 (N_17531,N_14413,N_14241);
xor U17532 (N_17532,N_13971,N_14257);
nand U17533 (N_17533,N_12053,N_12292);
or U17534 (N_17534,N_12331,N_13923);
or U17535 (N_17535,N_11194,N_11115);
nand U17536 (N_17536,N_13221,N_11429);
xor U17537 (N_17537,N_12524,N_10997);
nor U17538 (N_17538,N_10137,N_13473);
or U17539 (N_17539,N_11338,N_13623);
or U17540 (N_17540,N_12238,N_14191);
and U17541 (N_17541,N_14606,N_14718);
nor U17542 (N_17542,N_11032,N_12349);
nand U17543 (N_17543,N_12612,N_14991);
nand U17544 (N_17544,N_14255,N_14061);
and U17545 (N_17545,N_14065,N_14827);
xnor U17546 (N_17546,N_14733,N_11198);
nor U17547 (N_17547,N_11613,N_12887);
and U17548 (N_17548,N_11805,N_13631);
nor U17549 (N_17549,N_12771,N_13394);
and U17550 (N_17550,N_12671,N_13528);
nand U17551 (N_17551,N_14287,N_12608);
and U17552 (N_17552,N_12600,N_12473);
or U17553 (N_17553,N_11036,N_10575);
or U17554 (N_17554,N_10017,N_14605);
nand U17555 (N_17555,N_10966,N_13186);
or U17556 (N_17556,N_13259,N_14679);
nor U17557 (N_17557,N_14312,N_12188);
or U17558 (N_17558,N_12836,N_11605);
xnor U17559 (N_17559,N_12416,N_12362);
nor U17560 (N_17560,N_12382,N_14054);
or U17561 (N_17561,N_13902,N_14835);
and U17562 (N_17562,N_14014,N_11274);
and U17563 (N_17563,N_10491,N_10316);
and U17564 (N_17564,N_13277,N_11677);
xor U17565 (N_17565,N_14016,N_11568);
and U17566 (N_17566,N_10870,N_12900);
xnor U17567 (N_17567,N_12136,N_13015);
xnor U17568 (N_17568,N_11346,N_11492);
xor U17569 (N_17569,N_14681,N_14241);
nand U17570 (N_17570,N_12884,N_11756);
xor U17571 (N_17571,N_12330,N_11841);
nand U17572 (N_17572,N_13024,N_13188);
and U17573 (N_17573,N_13056,N_10349);
nor U17574 (N_17574,N_14469,N_10537);
xnor U17575 (N_17575,N_14324,N_10680);
or U17576 (N_17576,N_13208,N_13127);
xor U17577 (N_17577,N_14721,N_14190);
xor U17578 (N_17578,N_13476,N_12291);
nor U17579 (N_17579,N_14460,N_10227);
or U17580 (N_17580,N_12030,N_11295);
xor U17581 (N_17581,N_14477,N_13301);
xor U17582 (N_17582,N_10710,N_13003);
and U17583 (N_17583,N_14756,N_14132);
xor U17584 (N_17584,N_14044,N_11521);
nor U17585 (N_17585,N_14570,N_11809);
nand U17586 (N_17586,N_10129,N_14789);
or U17587 (N_17587,N_12573,N_13056);
and U17588 (N_17588,N_14112,N_11098);
and U17589 (N_17589,N_10307,N_12710);
xnor U17590 (N_17590,N_10282,N_14536);
or U17591 (N_17591,N_12227,N_12384);
or U17592 (N_17592,N_14753,N_13372);
nor U17593 (N_17593,N_10645,N_10864);
and U17594 (N_17594,N_13961,N_10815);
nand U17595 (N_17595,N_11786,N_13514);
nor U17596 (N_17596,N_12151,N_10689);
nand U17597 (N_17597,N_12318,N_14363);
and U17598 (N_17598,N_12200,N_12743);
or U17599 (N_17599,N_11252,N_13970);
or U17600 (N_17600,N_14009,N_13760);
and U17601 (N_17601,N_14663,N_14904);
xor U17602 (N_17602,N_14216,N_14073);
and U17603 (N_17603,N_10649,N_13731);
or U17604 (N_17604,N_12929,N_13680);
and U17605 (N_17605,N_12637,N_12838);
and U17606 (N_17606,N_13179,N_14260);
or U17607 (N_17607,N_14552,N_12538);
nor U17608 (N_17608,N_10174,N_10848);
or U17609 (N_17609,N_12139,N_12663);
xor U17610 (N_17610,N_11746,N_10869);
nor U17611 (N_17611,N_14582,N_14930);
xor U17612 (N_17612,N_11918,N_12810);
nand U17613 (N_17613,N_12374,N_10995);
xor U17614 (N_17614,N_11513,N_12973);
xor U17615 (N_17615,N_13787,N_12569);
xnor U17616 (N_17616,N_11164,N_13140);
and U17617 (N_17617,N_13833,N_13683);
nor U17618 (N_17618,N_11275,N_14751);
nand U17619 (N_17619,N_11187,N_10500);
nand U17620 (N_17620,N_14694,N_12438);
and U17621 (N_17621,N_10380,N_12831);
nor U17622 (N_17622,N_10352,N_14527);
xnor U17623 (N_17623,N_13370,N_12886);
xnor U17624 (N_17624,N_13384,N_10835);
xor U17625 (N_17625,N_14881,N_13531);
xnor U17626 (N_17626,N_11023,N_10018);
xnor U17627 (N_17627,N_14666,N_13958);
or U17628 (N_17628,N_14008,N_10261);
or U17629 (N_17629,N_10590,N_14446);
nand U17630 (N_17630,N_14628,N_14939);
nand U17631 (N_17631,N_14625,N_12935);
or U17632 (N_17632,N_12885,N_13685);
xor U17633 (N_17633,N_14484,N_13294);
and U17634 (N_17634,N_10243,N_14760);
xnor U17635 (N_17635,N_13851,N_12700);
xor U17636 (N_17636,N_13970,N_13279);
nand U17637 (N_17637,N_13591,N_13423);
nand U17638 (N_17638,N_10850,N_10462);
or U17639 (N_17639,N_13613,N_12480);
and U17640 (N_17640,N_14280,N_13212);
or U17641 (N_17641,N_11502,N_14344);
or U17642 (N_17642,N_11763,N_14837);
xnor U17643 (N_17643,N_10319,N_14834);
xor U17644 (N_17644,N_13694,N_12552);
nor U17645 (N_17645,N_10342,N_11028);
and U17646 (N_17646,N_14965,N_13287);
nand U17647 (N_17647,N_14454,N_10168);
nand U17648 (N_17648,N_11418,N_13274);
nand U17649 (N_17649,N_10716,N_12647);
nor U17650 (N_17650,N_14949,N_11185);
xor U17651 (N_17651,N_12233,N_14917);
nand U17652 (N_17652,N_12031,N_10212);
and U17653 (N_17653,N_14330,N_10402);
and U17654 (N_17654,N_14972,N_12024);
and U17655 (N_17655,N_10968,N_14529);
nor U17656 (N_17656,N_12004,N_13236);
nand U17657 (N_17657,N_10560,N_14614);
nand U17658 (N_17658,N_12007,N_12831);
or U17659 (N_17659,N_14538,N_11635);
and U17660 (N_17660,N_14439,N_11958);
or U17661 (N_17661,N_11675,N_10383);
nor U17662 (N_17662,N_12741,N_14877);
nor U17663 (N_17663,N_13191,N_13074);
nand U17664 (N_17664,N_14386,N_12009);
nor U17665 (N_17665,N_12702,N_11251);
nand U17666 (N_17666,N_14647,N_14626);
and U17667 (N_17667,N_11653,N_12857);
or U17668 (N_17668,N_14977,N_11280);
nor U17669 (N_17669,N_13656,N_12367);
or U17670 (N_17670,N_11334,N_10773);
nand U17671 (N_17671,N_13055,N_10889);
nor U17672 (N_17672,N_13843,N_13865);
nor U17673 (N_17673,N_11927,N_10894);
nor U17674 (N_17674,N_14919,N_13455);
nor U17675 (N_17675,N_14027,N_10459);
xor U17676 (N_17676,N_13200,N_11787);
xnor U17677 (N_17677,N_14568,N_12411);
and U17678 (N_17678,N_14689,N_13875);
nor U17679 (N_17679,N_14760,N_14575);
nor U17680 (N_17680,N_11321,N_11166);
or U17681 (N_17681,N_11974,N_10612);
xnor U17682 (N_17682,N_14474,N_14256);
and U17683 (N_17683,N_12386,N_14945);
or U17684 (N_17684,N_11670,N_13515);
and U17685 (N_17685,N_14405,N_10179);
nand U17686 (N_17686,N_14722,N_12683);
or U17687 (N_17687,N_12225,N_11096);
xor U17688 (N_17688,N_10430,N_14239);
or U17689 (N_17689,N_14742,N_10655);
nor U17690 (N_17690,N_13829,N_12530);
nand U17691 (N_17691,N_11690,N_12757);
and U17692 (N_17692,N_11559,N_12102);
or U17693 (N_17693,N_11065,N_12337);
xnor U17694 (N_17694,N_11866,N_11959);
nor U17695 (N_17695,N_14190,N_14363);
or U17696 (N_17696,N_10077,N_12987);
xnor U17697 (N_17697,N_12225,N_10260);
and U17698 (N_17698,N_11843,N_10032);
and U17699 (N_17699,N_12198,N_10473);
or U17700 (N_17700,N_13552,N_10332);
nand U17701 (N_17701,N_11906,N_13684);
nor U17702 (N_17702,N_14377,N_11005);
nor U17703 (N_17703,N_10784,N_11987);
and U17704 (N_17704,N_14835,N_10543);
nor U17705 (N_17705,N_13053,N_14168);
and U17706 (N_17706,N_14103,N_11822);
nor U17707 (N_17707,N_12881,N_14461);
xnor U17708 (N_17708,N_12999,N_11157);
nand U17709 (N_17709,N_11018,N_11923);
or U17710 (N_17710,N_10419,N_12789);
or U17711 (N_17711,N_11426,N_14427);
nand U17712 (N_17712,N_12013,N_10167);
nand U17713 (N_17713,N_12446,N_12217);
xor U17714 (N_17714,N_13723,N_13375);
and U17715 (N_17715,N_13636,N_11337);
xnor U17716 (N_17716,N_12672,N_10394);
nor U17717 (N_17717,N_13114,N_13625);
or U17718 (N_17718,N_11953,N_14367);
nand U17719 (N_17719,N_13370,N_12728);
nand U17720 (N_17720,N_11504,N_12643);
xor U17721 (N_17721,N_12186,N_10654);
and U17722 (N_17722,N_12785,N_11516);
nor U17723 (N_17723,N_14764,N_12321);
or U17724 (N_17724,N_10743,N_13415);
nand U17725 (N_17725,N_11343,N_11770);
nor U17726 (N_17726,N_14902,N_14844);
nor U17727 (N_17727,N_13030,N_14372);
or U17728 (N_17728,N_13021,N_11518);
xnor U17729 (N_17729,N_10190,N_12650);
nand U17730 (N_17730,N_14267,N_13558);
nor U17731 (N_17731,N_13288,N_11270);
or U17732 (N_17732,N_14842,N_12645);
nand U17733 (N_17733,N_14450,N_13758);
nand U17734 (N_17734,N_11807,N_10717);
and U17735 (N_17735,N_10274,N_10285);
xor U17736 (N_17736,N_12791,N_11801);
nand U17737 (N_17737,N_11558,N_11403);
nor U17738 (N_17738,N_12393,N_12232);
nand U17739 (N_17739,N_10630,N_13270);
nor U17740 (N_17740,N_12716,N_12586);
nor U17741 (N_17741,N_12172,N_10007);
and U17742 (N_17742,N_10410,N_12398);
xor U17743 (N_17743,N_12500,N_13263);
nand U17744 (N_17744,N_13583,N_10729);
nor U17745 (N_17745,N_12969,N_11211);
xor U17746 (N_17746,N_13187,N_14994);
and U17747 (N_17747,N_11751,N_10886);
xor U17748 (N_17748,N_11512,N_10861);
nand U17749 (N_17749,N_14902,N_12346);
nor U17750 (N_17750,N_11872,N_12149);
and U17751 (N_17751,N_13815,N_11566);
nor U17752 (N_17752,N_11065,N_13350);
and U17753 (N_17753,N_13718,N_13325);
and U17754 (N_17754,N_12277,N_11116);
nand U17755 (N_17755,N_13991,N_10284);
xor U17756 (N_17756,N_11527,N_13741);
nor U17757 (N_17757,N_14097,N_14413);
nand U17758 (N_17758,N_14496,N_10974);
xor U17759 (N_17759,N_14443,N_13462);
and U17760 (N_17760,N_12974,N_12450);
xor U17761 (N_17761,N_13114,N_13986);
nand U17762 (N_17762,N_13886,N_11145);
and U17763 (N_17763,N_13611,N_10895);
nor U17764 (N_17764,N_12040,N_12664);
nor U17765 (N_17765,N_10267,N_13527);
nor U17766 (N_17766,N_12528,N_11212);
nor U17767 (N_17767,N_10027,N_12196);
nor U17768 (N_17768,N_12745,N_10841);
or U17769 (N_17769,N_14715,N_11451);
nand U17770 (N_17770,N_11562,N_14953);
nor U17771 (N_17771,N_11029,N_11318);
nand U17772 (N_17772,N_10485,N_12272);
nor U17773 (N_17773,N_10981,N_12142);
or U17774 (N_17774,N_12049,N_10353);
and U17775 (N_17775,N_13513,N_12467);
nor U17776 (N_17776,N_13095,N_10401);
nor U17777 (N_17777,N_14411,N_12070);
xnor U17778 (N_17778,N_14812,N_13292);
or U17779 (N_17779,N_14344,N_12288);
xnor U17780 (N_17780,N_10926,N_12094);
nor U17781 (N_17781,N_10758,N_10145);
nor U17782 (N_17782,N_11797,N_14225);
xnor U17783 (N_17783,N_10520,N_10876);
nor U17784 (N_17784,N_12006,N_11382);
nand U17785 (N_17785,N_13530,N_11091);
and U17786 (N_17786,N_13607,N_12955);
xor U17787 (N_17787,N_14541,N_13047);
nor U17788 (N_17788,N_10607,N_11558);
or U17789 (N_17789,N_11700,N_10766);
xnor U17790 (N_17790,N_13972,N_12526);
or U17791 (N_17791,N_14981,N_11509);
nor U17792 (N_17792,N_12591,N_11993);
nand U17793 (N_17793,N_14664,N_10772);
or U17794 (N_17794,N_11733,N_12554);
nand U17795 (N_17795,N_10696,N_10176);
nor U17796 (N_17796,N_12565,N_11465);
nand U17797 (N_17797,N_12928,N_11089);
or U17798 (N_17798,N_10971,N_10880);
nand U17799 (N_17799,N_10577,N_11958);
and U17800 (N_17800,N_11540,N_11658);
nor U17801 (N_17801,N_12852,N_14406);
and U17802 (N_17802,N_14343,N_11445);
and U17803 (N_17803,N_11438,N_14405);
nor U17804 (N_17804,N_11662,N_10271);
xor U17805 (N_17805,N_12177,N_13776);
nand U17806 (N_17806,N_10292,N_13179);
or U17807 (N_17807,N_10773,N_12506);
nor U17808 (N_17808,N_14884,N_13572);
or U17809 (N_17809,N_11556,N_13519);
xnor U17810 (N_17810,N_11565,N_14343);
and U17811 (N_17811,N_14145,N_12557);
and U17812 (N_17812,N_10293,N_10550);
and U17813 (N_17813,N_14509,N_11059);
or U17814 (N_17814,N_13280,N_12150);
or U17815 (N_17815,N_13728,N_11419);
xnor U17816 (N_17816,N_12774,N_14253);
or U17817 (N_17817,N_14143,N_13615);
xor U17818 (N_17818,N_13678,N_11300);
nor U17819 (N_17819,N_11928,N_11331);
or U17820 (N_17820,N_13910,N_14685);
nand U17821 (N_17821,N_11243,N_11292);
xor U17822 (N_17822,N_11077,N_12577);
or U17823 (N_17823,N_12144,N_14836);
nor U17824 (N_17824,N_14134,N_13303);
nand U17825 (N_17825,N_11122,N_10075);
nand U17826 (N_17826,N_13416,N_12728);
xor U17827 (N_17827,N_13671,N_10189);
and U17828 (N_17828,N_14455,N_10799);
nor U17829 (N_17829,N_10460,N_14091);
nor U17830 (N_17830,N_14338,N_12237);
xor U17831 (N_17831,N_14100,N_14162);
nor U17832 (N_17832,N_14940,N_14105);
nor U17833 (N_17833,N_13748,N_13099);
nor U17834 (N_17834,N_12861,N_12849);
xor U17835 (N_17835,N_11501,N_12043);
and U17836 (N_17836,N_12272,N_13656);
or U17837 (N_17837,N_10561,N_10932);
nor U17838 (N_17838,N_10209,N_12159);
xor U17839 (N_17839,N_11523,N_10069);
or U17840 (N_17840,N_10844,N_13425);
nand U17841 (N_17841,N_14435,N_14807);
xor U17842 (N_17842,N_13177,N_11630);
or U17843 (N_17843,N_10355,N_13431);
nand U17844 (N_17844,N_11157,N_11911);
nor U17845 (N_17845,N_10313,N_10546);
xnor U17846 (N_17846,N_10082,N_11570);
or U17847 (N_17847,N_13423,N_14000);
or U17848 (N_17848,N_13176,N_11595);
xor U17849 (N_17849,N_14280,N_10458);
xor U17850 (N_17850,N_11191,N_11618);
or U17851 (N_17851,N_13760,N_10248);
nand U17852 (N_17852,N_12236,N_11765);
and U17853 (N_17853,N_12680,N_12476);
and U17854 (N_17854,N_14911,N_12128);
nor U17855 (N_17855,N_11306,N_14062);
nand U17856 (N_17856,N_14044,N_13409);
xor U17857 (N_17857,N_11410,N_12630);
nand U17858 (N_17858,N_11427,N_13241);
and U17859 (N_17859,N_14515,N_11821);
and U17860 (N_17860,N_13590,N_10261);
nand U17861 (N_17861,N_13530,N_10336);
xor U17862 (N_17862,N_12374,N_13401);
nor U17863 (N_17863,N_13330,N_13447);
or U17864 (N_17864,N_10508,N_14785);
or U17865 (N_17865,N_12491,N_10161);
or U17866 (N_17866,N_10388,N_11121);
and U17867 (N_17867,N_13927,N_11803);
xnor U17868 (N_17868,N_11365,N_12997);
nor U17869 (N_17869,N_11645,N_10765);
and U17870 (N_17870,N_10150,N_12412);
nor U17871 (N_17871,N_10590,N_10755);
nand U17872 (N_17872,N_11420,N_10455);
nor U17873 (N_17873,N_11913,N_14067);
xor U17874 (N_17874,N_14269,N_14145);
nor U17875 (N_17875,N_11345,N_14381);
xnor U17876 (N_17876,N_10210,N_14735);
and U17877 (N_17877,N_13464,N_14842);
nor U17878 (N_17878,N_13836,N_10124);
nand U17879 (N_17879,N_13711,N_14031);
or U17880 (N_17880,N_11410,N_14787);
xnor U17881 (N_17881,N_11366,N_12747);
nor U17882 (N_17882,N_14781,N_11987);
nand U17883 (N_17883,N_12168,N_14241);
nor U17884 (N_17884,N_11376,N_13530);
and U17885 (N_17885,N_13987,N_12086);
or U17886 (N_17886,N_14098,N_12854);
and U17887 (N_17887,N_10992,N_11064);
xnor U17888 (N_17888,N_13511,N_10558);
nor U17889 (N_17889,N_14596,N_14933);
or U17890 (N_17890,N_12558,N_12773);
or U17891 (N_17891,N_12316,N_13893);
nand U17892 (N_17892,N_13707,N_14642);
xor U17893 (N_17893,N_11248,N_12256);
nor U17894 (N_17894,N_13165,N_13855);
xor U17895 (N_17895,N_14703,N_13292);
nand U17896 (N_17896,N_12815,N_12999);
nor U17897 (N_17897,N_11186,N_11204);
xnor U17898 (N_17898,N_13306,N_12839);
xnor U17899 (N_17899,N_10448,N_11333);
xnor U17900 (N_17900,N_14657,N_12710);
or U17901 (N_17901,N_13232,N_10839);
and U17902 (N_17902,N_11048,N_10215);
or U17903 (N_17903,N_12413,N_10496);
or U17904 (N_17904,N_10309,N_13140);
nor U17905 (N_17905,N_13702,N_11224);
xnor U17906 (N_17906,N_12166,N_14414);
nor U17907 (N_17907,N_13773,N_13902);
or U17908 (N_17908,N_12158,N_13347);
or U17909 (N_17909,N_12621,N_11125);
and U17910 (N_17910,N_11785,N_10474);
xnor U17911 (N_17911,N_12283,N_10295);
xnor U17912 (N_17912,N_14738,N_11952);
nor U17913 (N_17913,N_11826,N_13104);
and U17914 (N_17914,N_14527,N_13626);
and U17915 (N_17915,N_14449,N_13798);
nand U17916 (N_17916,N_10000,N_12843);
and U17917 (N_17917,N_14352,N_10647);
or U17918 (N_17918,N_11644,N_14621);
nand U17919 (N_17919,N_14331,N_10761);
and U17920 (N_17920,N_14614,N_11970);
xnor U17921 (N_17921,N_12367,N_10536);
nor U17922 (N_17922,N_14585,N_14883);
or U17923 (N_17923,N_13042,N_12309);
or U17924 (N_17924,N_13038,N_10075);
and U17925 (N_17925,N_12267,N_11673);
xnor U17926 (N_17926,N_11652,N_14172);
nor U17927 (N_17927,N_12652,N_14086);
xor U17928 (N_17928,N_14013,N_14031);
nor U17929 (N_17929,N_14752,N_13495);
nand U17930 (N_17930,N_13455,N_12112);
xor U17931 (N_17931,N_13898,N_12122);
and U17932 (N_17932,N_11999,N_10026);
xor U17933 (N_17933,N_13200,N_12790);
nor U17934 (N_17934,N_13171,N_12009);
and U17935 (N_17935,N_10806,N_11480);
and U17936 (N_17936,N_10812,N_13148);
and U17937 (N_17937,N_10457,N_12729);
xnor U17938 (N_17938,N_14572,N_12340);
or U17939 (N_17939,N_10864,N_14637);
nand U17940 (N_17940,N_14448,N_11568);
nor U17941 (N_17941,N_11560,N_10434);
xor U17942 (N_17942,N_11436,N_12063);
xor U17943 (N_17943,N_14322,N_14469);
and U17944 (N_17944,N_11033,N_13169);
or U17945 (N_17945,N_11413,N_13417);
xor U17946 (N_17946,N_13454,N_11096);
or U17947 (N_17947,N_13851,N_14742);
and U17948 (N_17948,N_14950,N_10519);
nor U17949 (N_17949,N_10199,N_14991);
nand U17950 (N_17950,N_12860,N_12881);
xnor U17951 (N_17951,N_11231,N_13303);
and U17952 (N_17952,N_10632,N_12805);
and U17953 (N_17953,N_13228,N_12768);
and U17954 (N_17954,N_10995,N_10675);
or U17955 (N_17955,N_12692,N_13366);
nand U17956 (N_17956,N_12147,N_10896);
nor U17957 (N_17957,N_14767,N_14707);
xor U17958 (N_17958,N_13654,N_13511);
nand U17959 (N_17959,N_13647,N_13478);
nand U17960 (N_17960,N_11731,N_11346);
or U17961 (N_17961,N_13399,N_13261);
or U17962 (N_17962,N_14453,N_14834);
or U17963 (N_17963,N_10019,N_10265);
or U17964 (N_17964,N_13913,N_13302);
or U17965 (N_17965,N_13656,N_12519);
xor U17966 (N_17966,N_13610,N_11794);
nor U17967 (N_17967,N_14662,N_12508);
and U17968 (N_17968,N_13043,N_12214);
and U17969 (N_17969,N_10296,N_13067);
nor U17970 (N_17970,N_12768,N_14735);
nor U17971 (N_17971,N_11520,N_13067);
xnor U17972 (N_17972,N_14008,N_11583);
and U17973 (N_17973,N_13399,N_14948);
xnor U17974 (N_17974,N_13393,N_14755);
xnor U17975 (N_17975,N_11052,N_10956);
and U17976 (N_17976,N_14251,N_13286);
and U17977 (N_17977,N_12295,N_11956);
and U17978 (N_17978,N_13841,N_14413);
xnor U17979 (N_17979,N_11021,N_14050);
nor U17980 (N_17980,N_13047,N_13785);
nand U17981 (N_17981,N_12153,N_11941);
nor U17982 (N_17982,N_12597,N_13739);
xnor U17983 (N_17983,N_14140,N_10840);
and U17984 (N_17984,N_13834,N_13374);
or U17985 (N_17985,N_13940,N_13626);
or U17986 (N_17986,N_12810,N_11950);
and U17987 (N_17987,N_13439,N_11696);
nor U17988 (N_17988,N_13629,N_10842);
nor U17989 (N_17989,N_11614,N_11362);
and U17990 (N_17990,N_14752,N_13985);
or U17991 (N_17991,N_14107,N_12225);
or U17992 (N_17992,N_12849,N_13002);
or U17993 (N_17993,N_13965,N_14983);
or U17994 (N_17994,N_10273,N_13586);
nor U17995 (N_17995,N_10730,N_14303);
nor U17996 (N_17996,N_11369,N_14719);
nand U17997 (N_17997,N_12458,N_13746);
or U17998 (N_17998,N_13534,N_11241);
nor U17999 (N_17999,N_13430,N_11526);
xnor U18000 (N_18000,N_11789,N_12534);
and U18001 (N_18001,N_12567,N_13795);
and U18002 (N_18002,N_10346,N_12827);
and U18003 (N_18003,N_11522,N_13849);
nand U18004 (N_18004,N_11240,N_14085);
or U18005 (N_18005,N_10081,N_14197);
or U18006 (N_18006,N_10423,N_14605);
nor U18007 (N_18007,N_11850,N_14629);
nor U18008 (N_18008,N_13215,N_12532);
nor U18009 (N_18009,N_14353,N_11547);
or U18010 (N_18010,N_13190,N_10240);
and U18011 (N_18011,N_14479,N_10910);
xor U18012 (N_18012,N_13384,N_13235);
or U18013 (N_18013,N_11206,N_12008);
and U18014 (N_18014,N_14660,N_11791);
xor U18015 (N_18015,N_10668,N_13192);
and U18016 (N_18016,N_14620,N_14008);
xnor U18017 (N_18017,N_13424,N_14163);
nand U18018 (N_18018,N_14584,N_14724);
and U18019 (N_18019,N_13303,N_11695);
or U18020 (N_18020,N_12247,N_11338);
nand U18021 (N_18021,N_10702,N_10033);
or U18022 (N_18022,N_11981,N_14083);
or U18023 (N_18023,N_11913,N_10327);
or U18024 (N_18024,N_14190,N_12226);
nor U18025 (N_18025,N_10356,N_13044);
or U18026 (N_18026,N_13213,N_13641);
and U18027 (N_18027,N_12045,N_13865);
or U18028 (N_18028,N_13621,N_11855);
nand U18029 (N_18029,N_10315,N_11172);
nor U18030 (N_18030,N_10039,N_10343);
and U18031 (N_18031,N_14562,N_11989);
xor U18032 (N_18032,N_11085,N_12339);
nor U18033 (N_18033,N_14069,N_13707);
xor U18034 (N_18034,N_11355,N_11682);
or U18035 (N_18035,N_10298,N_13070);
nor U18036 (N_18036,N_13964,N_11755);
nor U18037 (N_18037,N_11500,N_14359);
nor U18038 (N_18038,N_12896,N_14770);
or U18039 (N_18039,N_11201,N_11651);
xnor U18040 (N_18040,N_13364,N_10556);
or U18041 (N_18041,N_12660,N_12297);
xnor U18042 (N_18042,N_11114,N_13737);
nor U18043 (N_18043,N_12981,N_11969);
xor U18044 (N_18044,N_13626,N_12607);
xnor U18045 (N_18045,N_14691,N_13125);
nand U18046 (N_18046,N_13575,N_13963);
nand U18047 (N_18047,N_10851,N_13558);
nand U18048 (N_18048,N_12607,N_12555);
nand U18049 (N_18049,N_11666,N_10556);
nor U18050 (N_18050,N_13019,N_13403);
nor U18051 (N_18051,N_13663,N_10209);
nor U18052 (N_18052,N_13143,N_14200);
or U18053 (N_18053,N_10912,N_14168);
and U18054 (N_18054,N_12586,N_14610);
nor U18055 (N_18055,N_11338,N_14111);
and U18056 (N_18056,N_10952,N_10426);
xor U18057 (N_18057,N_14424,N_12412);
and U18058 (N_18058,N_10717,N_10947);
or U18059 (N_18059,N_10252,N_14601);
nor U18060 (N_18060,N_14902,N_10210);
nor U18061 (N_18061,N_11299,N_13135);
nor U18062 (N_18062,N_13306,N_13334);
nor U18063 (N_18063,N_10667,N_14218);
nor U18064 (N_18064,N_11037,N_11560);
nor U18065 (N_18065,N_11312,N_10013);
xor U18066 (N_18066,N_12445,N_13627);
nor U18067 (N_18067,N_14789,N_13359);
nand U18068 (N_18068,N_13032,N_12253);
xnor U18069 (N_18069,N_12855,N_11248);
nand U18070 (N_18070,N_11614,N_14657);
or U18071 (N_18071,N_14682,N_10622);
xnor U18072 (N_18072,N_10075,N_13592);
nand U18073 (N_18073,N_12027,N_11298);
nand U18074 (N_18074,N_13081,N_10305);
nand U18075 (N_18075,N_13534,N_11090);
nor U18076 (N_18076,N_12190,N_11840);
xnor U18077 (N_18077,N_14676,N_10046);
nor U18078 (N_18078,N_13447,N_11739);
and U18079 (N_18079,N_10270,N_14409);
nor U18080 (N_18080,N_10694,N_12326);
and U18081 (N_18081,N_10680,N_10894);
and U18082 (N_18082,N_10889,N_14490);
xnor U18083 (N_18083,N_11029,N_13772);
nand U18084 (N_18084,N_10604,N_13108);
nand U18085 (N_18085,N_12382,N_10523);
xnor U18086 (N_18086,N_13301,N_14311);
nor U18087 (N_18087,N_13867,N_12753);
and U18088 (N_18088,N_10018,N_13056);
nor U18089 (N_18089,N_10759,N_13861);
nand U18090 (N_18090,N_14340,N_10344);
nand U18091 (N_18091,N_11240,N_13378);
and U18092 (N_18092,N_11373,N_14653);
nor U18093 (N_18093,N_10392,N_10758);
nand U18094 (N_18094,N_10976,N_10374);
or U18095 (N_18095,N_10710,N_11434);
and U18096 (N_18096,N_14507,N_14564);
nand U18097 (N_18097,N_13922,N_10710);
or U18098 (N_18098,N_10245,N_14131);
and U18099 (N_18099,N_13330,N_14791);
and U18100 (N_18100,N_10555,N_11138);
xnor U18101 (N_18101,N_13634,N_10764);
xor U18102 (N_18102,N_14316,N_14910);
nand U18103 (N_18103,N_12039,N_11613);
or U18104 (N_18104,N_12362,N_13291);
nor U18105 (N_18105,N_11709,N_12332);
and U18106 (N_18106,N_14374,N_13238);
xor U18107 (N_18107,N_12203,N_10530);
xnor U18108 (N_18108,N_10549,N_10054);
xor U18109 (N_18109,N_10443,N_13525);
nand U18110 (N_18110,N_13049,N_14318);
nor U18111 (N_18111,N_13512,N_14578);
nor U18112 (N_18112,N_13562,N_11412);
or U18113 (N_18113,N_12806,N_14480);
xnor U18114 (N_18114,N_13031,N_12926);
nor U18115 (N_18115,N_11819,N_11244);
xnor U18116 (N_18116,N_12844,N_12073);
or U18117 (N_18117,N_12923,N_14231);
nand U18118 (N_18118,N_10234,N_14103);
nor U18119 (N_18119,N_11537,N_11133);
xnor U18120 (N_18120,N_12170,N_12445);
xnor U18121 (N_18121,N_13437,N_14914);
or U18122 (N_18122,N_11609,N_11640);
nor U18123 (N_18123,N_14104,N_10459);
nand U18124 (N_18124,N_12057,N_12707);
and U18125 (N_18125,N_11150,N_14163);
nand U18126 (N_18126,N_10429,N_11986);
nor U18127 (N_18127,N_12599,N_12733);
and U18128 (N_18128,N_14470,N_10324);
nor U18129 (N_18129,N_14540,N_11077);
nand U18130 (N_18130,N_12104,N_12287);
nand U18131 (N_18131,N_11325,N_12437);
xor U18132 (N_18132,N_10766,N_14375);
or U18133 (N_18133,N_14442,N_11442);
nand U18134 (N_18134,N_13596,N_10327);
and U18135 (N_18135,N_14516,N_13795);
nor U18136 (N_18136,N_11532,N_10761);
or U18137 (N_18137,N_14454,N_10777);
nor U18138 (N_18138,N_13323,N_14178);
or U18139 (N_18139,N_11826,N_13963);
xnor U18140 (N_18140,N_14553,N_10909);
xnor U18141 (N_18141,N_12537,N_11226);
and U18142 (N_18142,N_11256,N_14625);
nor U18143 (N_18143,N_10411,N_11333);
or U18144 (N_18144,N_10070,N_14634);
nor U18145 (N_18145,N_14878,N_11297);
or U18146 (N_18146,N_11926,N_13054);
nand U18147 (N_18147,N_12694,N_14495);
nor U18148 (N_18148,N_13053,N_14775);
or U18149 (N_18149,N_11342,N_10357);
or U18150 (N_18150,N_12603,N_12793);
or U18151 (N_18151,N_10517,N_13126);
or U18152 (N_18152,N_13734,N_11031);
and U18153 (N_18153,N_14316,N_10983);
nor U18154 (N_18154,N_11998,N_13464);
or U18155 (N_18155,N_13016,N_13758);
xor U18156 (N_18156,N_10291,N_12596);
and U18157 (N_18157,N_12180,N_13423);
nor U18158 (N_18158,N_13793,N_13812);
nor U18159 (N_18159,N_11818,N_11711);
or U18160 (N_18160,N_11168,N_13304);
xnor U18161 (N_18161,N_14146,N_14811);
nand U18162 (N_18162,N_14914,N_10786);
nand U18163 (N_18163,N_13486,N_14267);
or U18164 (N_18164,N_14935,N_13530);
or U18165 (N_18165,N_12831,N_10199);
xor U18166 (N_18166,N_12321,N_12317);
xnor U18167 (N_18167,N_12819,N_13653);
xnor U18168 (N_18168,N_11456,N_13600);
nor U18169 (N_18169,N_11309,N_10000);
nor U18170 (N_18170,N_14190,N_13677);
and U18171 (N_18171,N_13871,N_11562);
and U18172 (N_18172,N_13889,N_12320);
or U18173 (N_18173,N_10324,N_13898);
nor U18174 (N_18174,N_11372,N_11814);
and U18175 (N_18175,N_12178,N_14975);
nand U18176 (N_18176,N_10325,N_13206);
or U18177 (N_18177,N_13074,N_14646);
nand U18178 (N_18178,N_10757,N_14315);
or U18179 (N_18179,N_14928,N_11331);
and U18180 (N_18180,N_10329,N_13973);
and U18181 (N_18181,N_10103,N_14255);
nor U18182 (N_18182,N_14220,N_10121);
xnor U18183 (N_18183,N_13147,N_12954);
xnor U18184 (N_18184,N_13160,N_13876);
nand U18185 (N_18185,N_14866,N_11097);
and U18186 (N_18186,N_14245,N_14743);
xnor U18187 (N_18187,N_14082,N_12255);
and U18188 (N_18188,N_11902,N_10742);
and U18189 (N_18189,N_14460,N_11318);
or U18190 (N_18190,N_11098,N_13283);
xnor U18191 (N_18191,N_13566,N_14748);
or U18192 (N_18192,N_14002,N_11847);
and U18193 (N_18193,N_14458,N_12737);
and U18194 (N_18194,N_10883,N_12232);
nor U18195 (N_18195,N_14893,N_12516);
nor U18196 (N_18196,N_13967,N_13126);
xor U18197 (N_18197,N_14983,N_13773);
nand U18198 (N_18198,N_13653,N_11276);
or U18199 (N_18199,N_11469,N_12994);
nor U18200 (N_18200,N_13858,N_14988);
or U18201 (N_18201,N_13210,N_12034);
nand U18202 (N_18202,N_14970,N_11895);
or U18203 (N_18203,N_11521,N_10448);
nand U18204 (N_18204,N_10930,N_11408);
xnor U18205 (N_18205,N_12735,N_13330);
nand U18206 (N_18206,N_14750,N_10929);
and U18207 (N_18207,N_12617,N_11894);
or U18208 (N_18208,N_10982,N_14235);
xnor U18209 (N_18209,N_10134,N_10218);
nand U18210 (N_18210,N_10090,N_14950);
and U18211 (N_18211,N_10647,N_11365);
or U18212 (N_18212,N_14877,N_11102);
or U18213 (N_18213,N_12687,N_10221);
nand U18214 (N_18214,N_14988,N_14036);
nand U18215 (N_18215,N_10394,N_13108);
or U18216 (N_18216,N_11003,N_10629);
nand U18217 (N_18217,N_11062,N_14191);
and U18218 (N_18218,N_10916,N_12175);
nor U18219 (N_18219,N_14235,N_14747);
and U18220 (N_18220,N_11625,N_11470);
or U18221 (N_18221,N_14062,N_13739);
xnor U18222 (N_18222,N_13343,N_10631);
and U18223 (N_18223,N_10737,N_12674);
xnor U18224 (N_18224,N_11335,N_10121);
nor U18225 (N_18225,N_12381,N_12798);
xor U18226 (N_18226,N_10768,N_12480);
xnor U18227 (N_18227,N_12970,N_10977);
or U18228 (N_18228,N_12668,N_10561);
nor U18229 (N_18229,N_14962,N_10737);
xnor U18230 (N_18230,N_11639,N_12911);
and U18231 (N_18231,N_13427,N_10329);
xnor U18232 (N_18232,N_13574,N_13096);
and U18233 (N_18233,N_14027,N_13222);
and U18234 (N_18234,N_12955,N_14911);
xor U18235 (N_18235,N_14261,N_11156);
xnor U18236 (N_18236,N_12998,N_10033);
xnor U18237 (N_18237,N_13109,N_12520);
xor U18238 (N_18238,N_10898,N_10673);
or U18239 (N_18239,N_14354,N_13423);
or U18240 (N_18240,N_13483,N_12239);
nor U18241 (N_18241,N_12173,N_10183);
nand U18242 (N_18242,N_14519,N_11454);
nor U18243 (N_18243,N_11248,N_11361);
or U18244 (N_18244,N_11010,N_11479);
nor U18245 (N_18245,N_11077,N_14914);
and U18246 (N_18246,N_12705,N_11766);
or U18247 (N_18247,N_10354,N_10678);
and U18248 (N_18248,N_14168,N_14257);
nand U18249 (N_18249,N_14693,N_14900);
and U18250 (N_18250,N_14181,N_13858);
xnor U18251 (N_18251,N_13635,N_10679);
nand U18252 (N_18252,N_14848,N_11573);
and U18253 (N_18253,N_13886,N_14368);
nand U18254 (N_18254,N_11288,N_13640);
nand U18255 (N_18255,N_14858,N_10619);
xnor U18256 (N_18256,N_13222,N_10528);
xnor U18257 (N_18257,N_12122,N_10942);
and U18258 (N_18258,N_13762,N_13672);
or U18259 (N_18259,N_12906,N_13747);
and U18260 (N_18260,N_11511,N_14094);
and U18261 (N_18261,N_14807,N_14414);
and U18262 (N_18262,N_12388,N_12409);
nand U18263 (N_18263,N_10094,N_13675);
nand U18264 (N_18264,N_12272,N_12102);
xor U18265 (N_18265,N_12671,N_14907);
and U18266 (N_18266,N_13770,N_10704);
nor U18267 (N_18267,N_10674,N_13900);
and U18268 (N_18268,N_10357,N_13611);
nand U18269 (N_18269,N_14739,N_14567);
xnor U18270 (N_18270,N_10762,N_13780);
xor U18271 (N_18271,N_11023,N_10707);
nand U18272 (N_18272,N_14522,N_14692);
nand U18273 (N_18273,N_12362,N_14442);
or U18274 (N_18274,N_14566,N_13247);
xor U18275 (N_18275,N_10665,N_12333);
nor U18276 (N_18276,N_13065,N_11725);
or U18277 (N_18277,N_14877,N_13528);
or U18278 (N_18278,N_11183,N_13654);
nor U18279 (N_18279,N_10669,N_14907);
and U18280 (N_18280,N_14396,N_12966);
nand U18281 (N_18281,N_11103,N_10804);
or U18282 (N_18282,N_13577,N_14092);
nand U18283 (N_18283,N_11822,N_13540);
nand U18284 (N_18284,N_12986,N_12558);
nor U18285 (N_18285,N_13541,N_11087);
nor U18286 (N_18286,N_14378,N_14193);
xnor U18287 (N_18287,N_10410,N_12195);
or U18288 (N_18288,N_10929,N_13996);
nand U18289 (N_18289,N_11023,N_14736);
xnor U18290 (N_18290,N_13075,N_12049);
nand U18291 (N_18291,N_11059,N_12869);
nor U18292 (N_18292,N_14368,N_10341);
or U18293 (N_18293,N_11564,N_12837);
or U18294 (N_18294,N_13171,N_12275);
nand U18295 (N_18295,N_10631,N_10578);
or U18296 (N_18296,N_14102,N_14994);
nand U18297 (N_18297,N_11693,N_11668);
and U18298 (N_18298,N_13408,N_13564);
nor U18299 (N_18299,N_12727,N_11272);
and U18300 (N_18300,N_14453,N_13312);
nor U18301 (N_18301,N_12831,N_14506);
and U18302 (N_18302,N_10275,N_11367);
nor U18303 (N_18303,N_13931,N_10158);
nor U18304 (N_18304,N_14783,N_11116);
and U18305 (N_18305,N_12903,N_11209);
xor U18306 (N_18306,N_12304,N_11600);
xnor U18307 (N_18307,N_14692,N_10984);
xor U18308 (N_18308,N_10879,N_12912);
nand U18309 (N_18309,N_10390,N_11253);
or U18310 (N_18310,N_14761,N_10461);
nand U18311 (N_18311,N_12741,N_14764);
or U18312 (N_18312,N_13801,N_12165);
and U18313 (N_18313,N_13880,N_11672);
nor U18314 (N_18314,N_14723,N_12243);
or U18315 (N_18315,N_12795,N_13205);
nor U18316 (N_18316,N_13733,N_11879);
nor U18317 (N_18317,N_11599,N_13051);
and U18318 (N_18318,N_14582,N_11121);
and U18319 (N_18319,N_11363,N_12868);
nor U18320 (N_18320,N_12079,N_14286);
and U18321 (N_18321,N_11822,N_14095);
xor U18322 (N_18322,N_14645,N_14497);
or U18323 (N_18323,N_12966,N_11096);
or U18324 (N_18324,N_11710,N_11841);
nand U18325 (N_18325,N_11782,N_10274);
nand U18326 (N_18326,N_14281,N_12511);
nand U18327 (N_18327,N_10472,N_13337);
nor U18328 (N_18328,N_13890,N_10011);
and U18329 (N_18329,N_13955,N_10153);
and U18330 (N_18330,N_13000,N_12550);
and U18331 (N_18331,N_10724,N_11906);
or U18332 (N_18332,N_14675,N_14033);
nand U18333 (N_18333,N_13459,N_14517);
nor U18334 (N_18334,N_12671,N_12995);
or U18335 (N_18335,N_14030,N_12699);
and U18336 (N_18336,N_11667,N_13494);
nor U18337 (N_18337,N_11033,N_13971);
xor U18338 (N_18338,N_14618,N_11939);
or U18339 (N_18339,N_12006,N_13666);
or U18340 (N_18340,N_14966,N_13569);
xnor U18341 (N_18341,N_12006,N_13197);
and U18342 (N_18342,N_14457,N_11392);
nand U18343 (N_18343,N_13143,N_13699);
nor U18344 (N_18344,N_14387,N_11320);
xnor U18345 (N_18345,N_10311,N_11992);
nor U18346 (N_18346,N_11453,N_10882);
nand U18347 (N_18347,N_13536,N_13380);
or U18348 (N_18348,N_10878,N_14936);
and U18349 (N_18349,N_12842,N_11521);
nand U18350 (N_18350,N_11208,N_14099);
nor U18351 (N_18351,N_13055,N_12921);
nor U18352 (N_18352,N_13472,N_12307);
xnor U18353 (N_18353,N_12037,N_11846);
or U18354 (N_18354,N_14128,N_12781);
nor U18355 (N_18355,N_13489,N_12519);
nand U18356 (N_18356,N_10826,N_13446);
and U18357 (N_18357,N_10822,N_11549);
and U18358 (N_18358,N_11002,N_11297);
xor U18359 (N_18359,N_13599,N_13198);
nand U18360 (N_18360,N_10428,N_11685);
nand U18361 (N_18361,N_10207,N_14273);
nor U18362 (N_18362,N_14041,N_13881);
xor U18363 (N_18363,N_12361,N_11340);
nand U18364 (N_18364,N_12796,N_13351);
and U18365 (N_18365,N_10688,N_11795);
and U18366 (N_18366,N_14786,N_11583);
nand U18367 (N_18367,N_13891,N_10656);
and U18368 (N_18368,N_13932,N_14206);
nor U18369 (N_18369,N_14495,N_13521);
xnor U18370 (N_18370,N_12021,N_10568);
xnor U18371 (N_18371,N_11748,N_11032);
and U18372 (N_18372,N_10092,N_14062);
nand U18373 (N_18373,N_14077,N_14412);
or U18374 (N_18374,N_12860,N_11403);
xor U18375 (N_18375,N_14857,N_14182);
or U18376 (N_18376,N_11369,N_12050);
nor U18377 (N_18377,N_14181,N_10710);
nor U18378 (N_18378,N_12942,N_12529);
nor U18379 (N_18379,N_10462,N_14869);
nand U18380 (N_18380,N_10957,N_11435);
and U18381 (N_18381,N_11646,N_11942);
and U18382 (N_18382,N_11059,N_10390);
xor U18383 (N_18383,N_12694,N_10595);
xnor U18384 (N_18384,N_10927,N_12279);
xor U18385 (N_18385,N_12349,N_14790);
and U18386 (N_18386,N_10586,N_11115);
nand U18387 (N_18387,N_14362,N_13269);
or U18388 (N_18388,N_10236,N_12464);
nor U18389 (N_18389,N_12309,N_13001);
and U18390 (N_18390,N_14087,N_14171);
nor U18391 (N_18391,N_10693,N_14816);
nand U18392 (N_18392,N_12376,N_11016);
or U18393 (N_18393,N_11815,N_10762);
nand U18394 (N_18394,N_11501,N_14151);
and U18395 (N_18395,N_14015,N_10528);
nand U18396 (N_18396,N_10473,N_11783);
xor U18397 (N_18397,N_12149,N_11970);
xor U18398 (N_18398,N_12518,N_11694);
nand U18399 (N_18399,N_14602,N_10811);
nor U18400 (N_18400,N_12459,N_11586);
or U18401 (N_18401,N_11136,N_12622);
or U18402 (N_18402,N_12355,N_12122);
xor U18403 (N_18403,N_13514,N_14468);
xor U18404 (N_18404,N_12974,N_10705);
xnor U18405 (N_18405,N_14226,N_10090);
and U18406 (N_18406,N_14506,N_11410);
and U18407 (N_18407,N_14747,N_10534);
and U18408 (N_18408,N_12254,N_14346);
or U18409 (N_18409,N_10296,N_10475);
or U18410 (N_18410,N_13636,N_13283);
or U18411 (N_18411,N_11998,N_10589);
and U18412 (N_18412,N_12228,N_11412);
and U18413 (N_18413,N_14275,N_11572);
xnor U18414 (N_18414,N_13694,N_13433);
nor U18415 (N_18415,N_14508,N_10030);
and U18416 (N_18416,N_14541,N_14067);
or U18417 (N_18417,N_13414,N_13193);
and U18418 (N_18418,N_11047,N_14201);
nand U18419 (N_18419,N_12950,N_10016);
nor U18420 (N_18420,N_11342,N_10316);
nand U18421 (N_18421,N_13455,N_14808);
and U18422 (N_18422,N_11875,N_14457);
xor U18423 (N_18423,N_10310,N_14554);
or U18424 (N_18424,N_12639,N_14209);
xnor U18425 (N_18425,N_14065,N_13914);
xor U18426 (N_18426,N_14790,N_14974);
nand U18427 (N_18427,N_11160,N_14813);
nor U18428 (N_18428,N_10721,N_10862);
nand U18429 (N_18429,N_10125,N_11145);
and U18430 (N_18430,N_10582,N_14922);
nor U18431 (N_18431,N_12066,N_10718);
or U18432 (N_18432,N_13033,N_12033);
nor U18433 (N_18433,N_11009,N_12647);
xor U18434 (N_18434,N_12436,N_11656);
or U18435 (N_18435,N_11102,N_13374);
nor U18436 (N_18436,N_11944,N_10958);
or U18437 (N_18437,N_13775,N_11797);
and U18438 (N_18438,N_14097,N_12155);
nor U18439 (N_18439,N_13222,N_13136);
nor U18440 (N_18440,N_10268,N_10987);
and U18441 (N_18441,N_12848,N_14121);
nor U18442 (N_18442,N_14609,N_12461);
nor U18443 (N_18443,N_12154,N_11275);
nor U18444 (N_18444,N_12161,N_14652);
and U18445 (N_18445,N_13485,N_12986);
or U18446 (N_18446,N_12536,N_10950);
nand U18447 (N_18447,N_14516,N_12872);
xor U18448 (N_18448,N_14458,N_11460);
nor U18449 (N_18449,N_11216,N_11272);
nand U18450 (N_18450,N_10657,N_13221);
and U18451 (N_18451,N_10152,N_13793);
or U18452 (N_18452,N_10036,N_10990);
or U18453 (N_18453,N_13895,N_14878);
and U18454 (N_18454,N_12402,N_12461);
nand U18455 (N_18455,N_11984,N_12707);
nor U18456 (N_18456,N_14300,N_12704);
and U18457 (N_18457,N_12641,N_10117);
nor U18458 (N_18458,N_12695,N_10173);
xnor U18459 (N_18459,N_13570,N_12921);
or U18460 (N_18460,N_13752,N_14689);
nor U18461 (N_18461,N_10656,N_11574);
and U18462 (N_18462,N_13425,N_13053);
nand U18463 (N_18463,N_14572,N_12486);
and U18464 (N_18464,N_13520,N_10691);
xnor U18465 (N_18465,N_11430,N_11518);
or U18466 (N_18466,N_14532,N_13138);
nor U18467 (N_18467,N_10545,N_11165);
and U18468 (N_18468,N_13580,N_10355);
nor U18469 (N_18469,N_14990,N_13119);
or U18470 (N_18470,N_11752,N_12360);
nor U18471 (N_18471,N_13649,N_10357);
or U18472 (N_18472,N_11910,N_13671);
and U18473 (N_18473,N_13031,N_12060);
nor U18474 (N_18474,N_12129,N_13627);
xor U18475 (N_18475,N_10186,N_11997);
and U18476 (N_18476,N_13990,N_12678);
or U18477 (N_18477,N_13875,N_11359);
nand U18478 (N_18478,N_14900,N_14608);
nand U18479 (N_18479,N_12822,N_14290);
or U18480 (N_18480,N_13230,N_13694);
and U18481 (N_18481,N_10594,N_11772);
xnor U18482 (N_18482,N_12167,N_13460);
nand U18483 (N_18483,N_11158,N_14175);
or U18484 (N_18484,N_14877,N_14002);
and U18485 (N_18485,N_13604,N_12487);
nand U18486 (N_18486,N_12358,N_12555);
nor U18487 (N_18487,N_12298,N_14696);
and U18488 (N_18488,N_12000,N_10563);
or U18489 (N_18489,N_13568,N_10111);
nand U18490 (N_18490,N_13410,N_14647);
or U18491 (N_18491,N_13453,N_14126);
xnor U18492 (N_18492,N_14893,N_10383);
xnor U18493 (N_18493,N_12176,N_12244);
or U18494 (N_18494,N_13904,N_13820);
nor U18495 (N_18495,N_14396,N_12087);
or U18496 (N_18496,N_10220,N_11930);
and U18497 (N_18497,N_14646,N_12656);
or U18498 (N_18498,N_12278,N_10808);
nor U18499 (N_18499,N_11007,N_13152);
or U18500 (N_18500,N_10265,N_11802);
and U18501 (N_18501,N_10327,N_13244);
and U18502 (N_18502,N_12625,N_13577);
nor U18503 (N_18503,N_14499,N_12600);
or U18504 (N_18504,N_12242,N_14438);
xor U18505 (N_18505,N_10180,N_10764);
xor U18506 (N_18506,N_11730,N_13298);
xor U18507 (N_18507,N_11430,N_13595);
and U18508 (N_18508,N_10183,N_11279);
nor U18509 (N_18509,N_12461,N_11654);
or U18510 (N_18510,N_14823,N_14953);
and U18511 (N_18511,N_11267,N_14753);
and U18512 (N_18512,N_11219,N_12391);
or U18513 (N_18513,N_14007,N_12212);
or U18514 (N_18514,N_11527,N_14107);
nor U18515 (N_18515,N_14489,N_12580);
nor U18516 (N_18516,N_12136,N_14671);
nor U18517 (N_18517,N_14622,N_10466);
or U18518 (N_18518,N_11554,N_13690);
nand U18519 (N_18519,N_12075,N_14674);
nor U18520 (N_18520,N_10883,N_13475);
nand U18521 (N_18521,N_11179,N_12833);
xor U18522 (N_18522,N_14635,N_12029);
xor U18523 (N_18523,N_10002,N_14278);
nand U18524 (N_18524,N_14543,N_10419);
nand U18525 (N_18525,N_13234,N_14262);
and U18526 (N_18526,N_14989,N_14363);
xor U18527 (N_18527,N_12372,N_13359);
and U18528 (N_18528,N_14443,N_11990);
nand U18529 (N_18529,N_11240,N_14385);
and U18530 (N_18530,N_13260,N_14228);
nand U18531 (N_18531,N_14595,N_13781);
xnor U18532 (N_18532,N_13175,N_12735);
nor U18533 (N_18533,N_12758,N_10829);
nor U18534 (N_18534,N_14662,N_12145);
nor U18535 (N_18535,N_13551,N_10096);
and U18536 (N_18536,N_10856,N_11134);
and U18537 (N_18537,N_11135,N_10279);
nand U18538 (N_18538,N_12943,N_11049);
and U18539 (N_18539,N_13046,N_11621);
xnor U18540 (N_18540,N_10969,N_14911);
or U18541 (N_18541,N_13990,N_10157);
nor U18542 (N_18542,N_11325,N_12579);
or U18543 (N_18543,N_12060,N_10464);
xor U18544 (N_18544,N_10495,N_11227);
nor U18545 (N_18545,N_12328,N_13467);
or U18546 (N_18546,N_13600,N_13345);
xnor U18547 (N_18547,N_12990,N_12443);
xnor U18548 (N_18548,N_13883,N_12364);
xnor U18549 (N_18549,N_10576,N_14195);
xor U18550 (N_18550,N_12900,N_10249);
and U18551 (N_18551,N_10005,N_10508);
and U18552 (N_18552,N_11110,N_10233);
nor U18553 (N_18553,N_14888,N_14453);
xnor U18554 (N_18554,N_12005,N_14601);
nor U18555 (N_18555,N_11975,N_14009);
nor U18556 (N_18556,N_14486,N_11406);
and U18557 (N_18557,N_14354,N_12164);
or U18558 (N_18558,N_12842,N_14770);
xnor U18559 (N_18559,N_13748,N_10801);
xor U18560 (N_18560,N_13063,N_12760);
or U18561 (N_18561,N_11249,N_10534);
and U18562 (N_18562,N_11698,N_11118);
or U18563 (N_18563,N_11320,N_14993);
or U18564 (N_18564,N_12128,N_13850);
and U18565 (N_18565,N_11469,N_12552);
nand U18566 (N_18566,N_11454,N_10904);
or U18567 (N_18567,N_10468,N_11185);
or U18568 (N_18568,N_13071,N_13523);
or U18569 (N_18569,N_12581,N_14026);
xnor U18570 (N_18570,N_14799,N_11933);
or U18571 (N_18571,N_12675,N_12300);
nand U18572 (N_18572,N_11355,N_10521);
nor U18573 (N_18573,N_14075,N_14765);
nor U18574 (N_18574,N_12731,N_10198);
nor U18575 (N_18575,N_11667,N_13703);
and U18576 (N_18576,N_10815,N_10597);
and U18577 (N_18577,N_10504,N_13741);
or U18578 (N_18578,N_12860,N_12655);
or U18579 (N_18579,N_12667,N_14776);
and U18580 (N_18580,N_13054,N_13400);
or U18581 (N_18581,N_10883,N_11454);
and U18582 (N_18582,N_11374,N_13280);
and U18583 (N_18583,N_12526,N_11831);
and U18584 (N_18584,N_14048,N_10522);
and U18585 (N_18585,N_11531,N_12909);
nor U18586 (N_18586,N_12966,N_11987);
nand U18587 (N_18587,N_13087,N_11551);
xor U18588 (N_18588,N_12501,N_13815);
nor U18589 (N_18589,N_14167,N_11677);
or U18590 (N_18590,N_11360,N_14648);
or U18591 (N_18591,N_13635,N_13813);
or U18592 (N_18592,N_14273,N_14943);
and U18593 (N_18593,N_12822,N_13241);
nor U18594 (N_18594,N_11369,N_12404);
or U18595 (N_18595,N_14249,N_14576);
xnor U18596 (N_18596,N_11728,N_13323);
or U18597 (N_18597,N_10530,N_10228);
nand U18598 (N_18598,N_13013,N_10096);
nand U18599 (N_18599,N_10388,N_11418);
nor U18600 (N_18600,N_13197,N_11181);
nand U18601 (N_18601,N_10017,N_13710);
xnor U18602 (N_18602,N_11121,N_13857);
and U18603 (N_18603,N_10557,N_14823);
nor U18604 (N_18604,N_11817,N_14291);
xor U18605 (N_18605,N_13841,N_10468);
or U18606 (N_18606,N_12912,N_12503);
and U18607 (N_18607,N_12139,N_14316);
nand U18608 (N_18608,N_14348,N_10613);
nand U18609 (N_18609,N_11046,N_14083);
nand U18610 (N_18610,N_13503,N_11019);
xnor U18611 (N_18611,N_14038,N_12783);
and U18612 (N_18612,N_12120,N_14819);
nor U18613 (N_18613,N_10567,N_10755);
and U18614 (N_18614,N_10727,N_13678);
and U18615 (N_18615,N_10451,N_13907);
and U18616 (N_18616,N_10595,N_14795);
nand U18617 (N_18617,N_14697,N_12155);
xor U18618 (N_18618,N_10671,N_12448);
nand U18619 (N_18619,N_13131,N_10663);
xor U18620 (N_18620,N_12412,N_13707);
and U18621 (N_18621,N_11591,N_14094);
and U18622 (N_18622,N_11593,N_12337);
nor U18623 (N_18623,N_13808,N_14069);
nor U18624 (N_18624,N_14515,N_12696);
and U18625 (N_18625,N_14369,N_11584);
nor U18626 (N_18626,N_14280,N_13188);
xnor U18627 (N_18627,N_12094,N_12688);
nand U18628 (N_18628,N_10854,N_10162);
xnor U18629 (N_18629,N_10382,N_10097);
nor U18630 (N_18630,N_12083,N_11029);
and U18631 (N_18631,N_11511,N_11797);
xor U18632 (N_18632,N_11378,N_14081);
nand U18633 (N_18633,N_12145,N_12306);
nor U18634 (N_18634,N_11760,N_13296);
and U18635 (N_18635,N_11263,N_14982);
nor U18636 (N_18636,N_14499,N_14769);
or U18637 (N_18637,N_10399,N_13593);
xor U18638 (N_18638,N_11022,N_10239);
xnor U18639 (N_18639,N_11263,N_13145);
or U18640 (N_18640,N_10728,N_12500);
nand U18641 (N_18641,N_12804,N_12304);
xor U18642 (N_18642,N_13791,N_10492);
nor U18643 (N_18643,N_13371,N_13480);
xnor U18644 (N_18644,N_14772,N_11278);
or U18645 (N_18645,N_12953,N_10108);
or U18646 (N_18646,N_10310,N_11904);
xnor U18647 (N_18647,N_14415,N_12352);
and U18648 (N_18648,N_12330,N_14739);
or U18649 (N_18649,N_11183,N_14512);
nor U18650 (N_18650,N_11155,N_10337);
nor U18651 (N_18651,N_14350,N_13250);
or U18652 (N_18652,N_12816,N_12335);
xor U18653 (N_18653,N_10462,N_11245);
nand U18654 (N_18654,N_11631,N_13482);
or U18655 (N_18655,N_11030,N_14017);
nor U18656 (N_18656,N_10606,N_14188);
nor U18657 (N_18657,N_14602,N_13248);
nand U18658 (N_18658,N_12850,N_14387);
and U18659 (N_18659,N_12803,N_10108);
xor U18660 (N_18660,N_11264,N_12298);
nand U18661 (N_18661,N_11479,N_10832);
xnor U18662 (N_18662,N_10548,N_11136);
nor U18663 (N_18663,N_11841,N_14880);
nand U18664 (N_18664,N_12087,N_10641);
nor U18665 (N_18665,N_10268,N_14824);
or U18666 (N_18666,N_10399,N_12598);
or U18667 (N_18667,N_10064,N_10923);
and U18668 (N_18668,N_11186,N_12020);
nor U18669 (N_18669,N_13517,N_10953);
nand U18670 (N_18670,N_12596,N_13731);
nand U18671 (N_18671,N_10400,N_11875);
or U18672 (N_18672,N_11715,N_14766);
or U18673 (N_18673,N_14255,N_12027);
or U18674 (N_18674,N_12803,N_12933);
or U18675 (N_18675,N_14834,N_11276);
or U18676 (N_18676,N_13916,N_13432);
or U18677 (N_18677,N_11005,N_11002);
and U18678 (N_18678,N_10607,N_12611);
nand U18679 (N_18679,N_10017,N_14950);
nand U18680 (N_18680,N_14175,N_13811);
nor U18681 (N_18681,N_12616,N_14267);
or U18682 (N_18682,N_10788,N_12547);
nand U18683 (N_18683,N_13029,N_10803);
nor U18684 (N_18684,N_13806,N_12283);
nor U18685 (N_18685,N_10090,N_13259);
xnor U18686 (N_18686,N_10812,N_14487);
nand U18687 (N_18687,N_13360,N_12133);
nor U18688 (N_18688,N_10860,N_11810);
xor U18689 (N_18689,N_11245,N_10925);
xor U18690 (N_18690,N_13124,N_11146);
and U18691 (N_18691,N_12810,N_14169);
nor U18692 (N_18692,N_14607,N_11287);
or U18693 (N_18693,N_11648,N_14561);
nand U18694 (N_18694,N_11159,N_10824);
nor U18695 (N_18695,N_12409,N_14953);
nand U18696 (N_18696,N_14757,N_13683);
xor U18697 (N_18697,N_12730,N_13773);
nor U18698 (N_18698,N_13707,N_14508);
nand U18699 (N_18699,N_11136,N_14365);
nor U18700 (N_18700,N_14262,N_13859);
nor U18701 (N_18701,N_12818,N_11987);
nand U18702 (N_18702,N_12445,N_12242);
nor U18703 (N_18703,N_14031,N_14757);
nand U18704 (N_18704,N_12957,N_14523);
xnor U18705 (N_18705,N_10636,N_12556);
xnor U18706 (N_18706,N_11676,N_10608);
and U18707 (N_18707,N_13095,N_13928);
or U18708 (N_18708,N_14847,N_12809);
and U18709 (N_18709,N_14777,N_13878);
nand U18710 (N_18710,N_11722,N_10848);
xor U18711 (N_18711,N_12470,N_14710);
nor U18712 (N_18712,N_10293,N_10620);
nor U18713 (N_18713,N_12262,N_11394);
or U18714 (N_18714,N_13576,N_10114);
or U18715 (N_18715,N_10773,N_12488);
nor U18716 (N_18716,N_11642,N_10677);
nor U18717 (N_18717,N_11792,N_10867);
or U18718 (N_18718,N_11663,N_12487);
nand U18719 (N_18719,N_11753,N_10187);
and U18720 (N_18720,N_12443,N_10592);
xor U18721 (N_18721,N_14463,N_10723);
nand U18722 (N_18722,N_12430,N_11134);
and U18723 (N_18723,N_14271,N_14107);
or U18724 (N_18724,N_13931,N_14856);
nand U18725 (N_18725,N_13614,N_11061);
xnor U18726 (N_18726,N_11808,N_10015);
nor U18727 (N_18727,N_11857,N_13917);
nand U18728 (N_18728,N_11117,N_12418);
nand U18729 (N_18729,N_13758,N_12443);
xnor U18730 (N_18730,N_11394,N_13578);
nand U18731 (N_18731,N_11045,N_12995);
xnor U18732 (N_18732,N_11776,N_13560);
nor U18733 (N_18733,N_11607,N_12835);
xnor U18734 (N_18734,N_12514,N_14133);
xor U18735 (N_18735,N_11297,N_10665);
nand U18736 (N_18736,N_13935,N_10275);
xor U18737 (N_18737,N_14396,N_12680);
xor U18738 (N_18738,N_11319,N_11798);
and U18739 (N_18739,N_11677,N_14857);
and U18740 (N_18740,N_11613,N_13771);
and U18741 (N_18741,N_10182,N_11121);
nor U18742 (N_18742,N_10395,N_13181);
nand U18743 (N_18743,N_13819,N_12076);
nand U18744 (N_18744,N_11454,N_13076);
xor U18745 (N_18745,N_12772,N_10921);
xor U18746 (N_18746,N_11579,N_10763);
nor U18747 (N_18747,N_12309,N_12990);
nand U18748 (N_18748,N_13383,N_12064);
nand U18749 (N_18749,N_14906,N_11965);
xor U18750 (N_18750,N_13795,N_10318);
and U18751 (N_18751,N_14409,N_10258);
and U18752 (N_18752,N_14150,N_10040);
or U18753 (N_18753,N_10107,N_12465);
or U18754 (N_18754,N_11207,N_14731);
or U18755 (N_18755,N_12646,N_10629);
xnor U18756 (N_18756,N_11804,N_10440);
and U18757 (N_18757,N_11989,N_12196);
xor U18758 (N_18758,N_13357,N_14605);
nor U18759 (N_18759,N_13548,N_11338);
xor U18760 (N_18760,N_13719,N_10234);
nand U18761 (N_18761,N_13702,N_13356);
xnor U18762 (N_18762,N_12141,N_12177);
nor U18763 (N_18763,N_11244,N_12331);
and U18764 (N_18764,N_11893,N_13956);
and U18765 (N_18765,N_10164,N_11612);
nand U18766 (N_18766,N_13178,N_12363);
or U18767 (N_18767,N_14445,N_12138);
and U18768 (N_18768,N_11314,N_10242);
and U18769 (N_18769,N_14113,N_14728);
xnor U18770 (N_18770,N_12288,N_10285);
and U18771 (N_18771,N_10341,N_10928);
and U18772 (N_18772,N_11957,N_14562);
xnor U18773 (N_18773,N_14575,N_12451);
or U18774 (N_18774,N_12882,N_11114);
nor U18775 (N_18775,N_12291,N_10727);
and U18776 (N_18776,N_11832,N_10397);
xor U18777 (N_18777,N_13793,N_11320);
xnor U18778 (N_18778,N_14623,N_14174);
nor U18779 (N_18779,N_10778,N_14935);
or U18780 (N_18780,N_11587,N_11283);
nand U18781 (N_18781,N_13943,N_13345);
xor U18782 (N_18782,N_12825,N_14170);
xor U18783 (N_18783,N_12618,N_13736);
xor U18784 (N_18784,N_10081,N_13214);
and U18785 (N_18785,N_10872,N_14237);
and U18786 (N_18786,N_14986,N_12919);
nor U18787 (N_18787,N_13232,N_12644);
xnor U18788 (N_18788,N_13301,N_10196);
and U18789 (N_18789,N_11922,N_13188);
and U18790 (N_18790,N_11819,N_10020);
or U18791 (N_18791,N_13448,N_14830);
and U18792 (N_18792,N_10438,N_10093);
nand U18793 (N_18793,N_12731,N_14445);
or U18794 (N_18794,N_12838,N_11163);
nor U18795 (N_18795,N_12354,N_14393);
or U18796 (N_18796,N_13189,N_11851);
nor U18797 (N_18797,N_14222,N_12835);
nor U18798 (N_18798,N_12694,N_12842);
or U18799 (N_18799,N_14624,N_12095);
or U18800 (N_18800,N_14980,N_12370);
xnor U18801 (N_18801,N_11384,N_11238);
and U18802 (N_18802,N_11559,N_10782);
xor U18803 (N_18803,N_11839,N_14083);
and U18804 (N_18804,N_11472,N_10774);
nor U18805 (N_18805,N_14841,N_12769);
and U18806 (N_18806,N_12098,N_10994);
and U18807 (N_18807,N_13212,N_10786);
and U18808 (N_18808,N_11518,N_12424);
and U18809 (N_18809,N_14756,N_12454);
xnor U18810 (N_18810,N_14122,N_13052);
or U18811 (N_18811,N_14345,N_10267);
and U18812 (N_18812,N_13166,N_12585);
xor U18813 (N_18813,N_13377,N_14569);
or U18814 (N_18814,N_14621,N_11245);
or U18815 (N_18815,N_12763,N_13428);
or U18816 (N_18816,N_14157,N_10678);
nand U18817 (N_18817,N_13877,N_12024);
or U18818 (N_18818,N_13695,N_14723);
nand U18819 (N_18819,N_12703,N_10217);
and U18820 (N_18820,N_14673,N_10794);
and U18821 (N_18821,N_10714,N_13759);
or U18822 (N_18822,N_12648,N_14211);
xnor U18823 (N_18823,N_12966,N_12145);
and U18824 (N_18824,N_11168,N_14937);
nand U18825 (N_18825,N_13776,N_14040);
nor U18826 (N_18826,N_12703,N_13627);
and U18827 (N_18827,N_10931,N_11454);
or U18828 (N_18828,N_13363,N_10207);
and U18829 (N_18829,N_10781,N_12508);
xnor U18830 (N_18830,N_12696,N_14702);
nand U18831 (N_18831,N_14681,N_14531);
or U18832 (N_18832,N_10851,N_12430);
xnor U18833 (N_18833,N_10179,N_11603);
and U18834 (N_18834,N_14971,N_13459);
nand U18835 (N_18835,N_10425,N_13781);
or U18836 (N_18836,N_13912,N_13387);
and U18837 (N_18837,N_10360,N_11134);
or U18838 (N_18838,N_14228,N_10036);
or U18839 (N_18839,N_11404,N_14046);
xor U18840 (N_18840,N_14314,N_14602);
nor U18841 (N_18841,N_10586,N_13957);
or U18842 (N_18842,N_10633,N_14322);
and U18843 (N_18843,N_11813,N_10547);
nor U18844 (N_18844,N_13120,N_14638);
or U18845 (N_18845,N_12781,N_14939);
nor U18846 (N_18846,N_10016,N_12708);
xor U18847 (N_18847,N_11611,N_10113);
nor U18848 (N_18848,N_14767,N_10125);
nand U18849 (N_18849,N_11743,N_10230);
and U18850 (N_18850,N_10833,N_13718);
nand U18851 (N_18851,N_13702,N_14392);
nor U18852 (N_18852,N_11245,N_10749);
nand U18853 (N_18853,N_14269,N_12678);
nor U18854 (N_18854,N_10399,N_13522);
or U18855 (N_18855,N_10060,N_12391);
nand U18856 (N_18856,N_10493,N_13343);
and U18857 (N_18857,N_10302,N_11918);
nor U18858 (N_18858,N_14677,N_10918);
or U18859 (N_18859,N_13919,N_10784);
nor U18860 (N_18860,N_14487,N_13460);
or U18861 (N_18861,N_11725,N_10650);
or U18862 (N_18862,N_14025,N_12777);
and U18863 (N_18863,N_13329,N_11544);
and U18864 (N_18864,N_11711,N_11359);
nor U18865 (N_18865,N_14674,N_14922);
and U18866 (N_18866,N_10163,N_12641);
or U18867 (N_18867,N_12197,N_10853);
nor U18868 (N_18868,N_10135,N_14558);
xnor U18869 (N_18869,N_12293,N_11468);
nor U18870 (N_18870,N_10284,N_13644);
or U18871 (N_18871,N_13372,N_12643);
and U18872 (N_18872,N_10689,N_14476);
or U18873 (N_18873,N_13513,N_10096);
and U18874 (N_18874,N_13462,N_11761);
or U18875 (N_18875,N_13951,N_10093);
xor U18876 (N_18876,N_12920,N_12203);
xnor U18877 (N_18877,N_14053,N_12223);
nand U18878 (N_18878,N_12543,N_14874);
xor U18879 (N_18879,N_14654,N_12045);
nor U18880 (N_18880,N_10776,N_12009);
nor U18881 (N_18881,N_11112,N_12595);
or U18882 (N_18882,N_11855,N_12722);
xor U18883 (N_18883,N_12605,N_13873);
or U18884 (N_18884,N_12432,N_12373);
and U18885 (N_18885,N_14216,N_13455);
xor U18886 (N_18886,N_11812,N_11135);
nor U18887 (N_18887,N_13085,N_13779);
and U18888 (N_18888,N_11949,N_14897);
or U18889 (N_18889,N_10369,N_13407);
xor U18890 (N_18890,N_10698,N_11332);
nor U18891 (N_18891,N_13739,N_14020);
and U18892 (N_18892,N_14008,N_12387);
or U18893 (N_18893,N_11620,N_13186);
xnor U18894 (N_18894,N_12029,N_12430);
and U18895 (N_18895,N_11020,N_10834);
or U18896 (N_18896,N_14387,N_13414);
and U18897 (N_18897,N_14642,N_14753);
xor U18898 (N_18898,N_10302,N_10493);
xor U18899 (N_18899,N_10907,N_13576);
or U18900 (N_18900,N_13929,N_12609);
xnor U18901 (N_18901,N_12958,N_13569);
xnor U18902 (N_18902,N_13163,N_12913);
xnor U18903 (N_18903,N_12418,N_14115);
or U18904 (N_18904,N_11636,N_14876);
xnor U18905 (N_18905,N_13230,N_11498);
nor U18906 (N_18906,N_11805,N_14965);
and U18907 (N_18907,N_12635,N_13930);
nand U18908 (N_18908,N_12228,N_12477);
or U18909 (N_18909,N_12769,N_12934);
xnor U18910 (N_18910,N_12493,N_11212);
xnor U18911 (N_18911,N_12261,N_11160);
nand U18912 (N_18912,N_14022,N_10251);
nand U18913 (N_18913,N_12181,N_10834);
and U18914 (N_18914,N_11743,N_14504);
xor U18915 (N_18915,N_11721,N_10905);
or U18916 (N_18916,N_14692,N_13161);
xor U18917 (N_18917,N_12957,N_12852);
and U18918 (N_18918,N_13828,N_12725);
and U18919 (N_18919,N_11303,N_10459);
nor U18920 (N_18920,N_11073,N_14650);
nor U18921 (N_18921,N_11556,N_11122);
nand U18922 (N_18922,N_14578,N_11864);
and U18923 (N_18923,N_12197,N_13869);
nor U18924 (N_18924,N_11845,N_12014);
nor U18925 (N_18925,N_14498,N_11806);
xor U18926 (N_18926,N_13756,N_14769);
nor U18927 (N_18927,N_11505,N_13407);
and U18928 (N_18928,N_12481,N_12582);
xnor U18929 (N_18929,N_12763,N_10637);
nand U18930 (N_18930,N_10839,N_14742);
nand U18931 (N_18931,N_13086,N_10732);
and U18932 (N_18932,N_13149,N_12917);
or U18933 (N_18933,N_13246,N_10493);
xnor U18934 (N_18934,N_11418,N_13987);
or U18935 (N_18935,N_10961,N_10105);
xor U18936 (N_18936,N_10629,N_14451);
nand U18937 (N_18937,N_10408,N_13096);
xor U18938 (N_18938,N_13456,N_11931);
nor U18939 (N_18939,N_14871,N_14803);
nand U18940 (N_18940,N_13758,N_11072);
and U18941 (N_18941,N_11934,N_11821);
nor U18942 (N_18942,N_14900,N_11392);
and U18943 (N_18943,N_10655,N_11527);
and U18944 (N_18944,N_12290,N_11332);
xnor U18945 (N_18945,N_13538,N_14192);
nand U18946 (N_18946,N_13139,N_13216);
nand U18947 (N_18947,N_13744,N_10606);
nor U18948 (N_18948,N_11925,N_10518);
nor U18949 (N_18949,N_13445,N_14885);
nand U18950 (N_18950,N_11790,N_11867);
xor U18951 (N_18951,N_10089,N_12871);
xnor U18952 (N_18952,N_14192,N_12150);
and U18953 (N_18953,N_14899,N_10268);
nand U18954 (N_18954,N_12376,N_10450);
xnor U18955 (N_18955,N_11122,N_10065);
nor U18956 (N_18956,N_11065,N_12384);
and U18957 (N_18957,N_14024,N_11519);
or U18958 (N_18958,N_13403,N_14896);
nor U18959 (N_18959,N_12728,N_12729);
and U18960 (N_18960,N_12347,N_10429);
nand U18961 (N_18961,N_11426,N_13496);
or U18962 (N_18962,N_10907,N_10893);
or U18963 (N_18963,N_14617,N_13195);
nand U18964 (N_18964,N_14715,N_11755);
nand U18965 (N_18965,N_10513,N_11427);
nor U18966 (N_18966,N_12262,N_10983);
nand U18967 (N_18967,N_12177,N_13813);
nor U18968 (N_18968,N_10867,N_13165);
xnor U18969 (N_18969,N_13602,N_13775);
nand U18970 (N_18970,N_11000,N_14502);
or U18971 (N_18971,N_13573,N_14163);
nand U18972 (N_18972,N_10749,N_13411);
nor U18973 (N_18973,N_12933,N_14707);
or U18974 (N_18974,N_12757,N_14057);
and U18975 (N_18975,N_10131,N_11208);
nand U18976 (N_18976,N_13039,N_10649);
xor U18977 (N_18977,N_11629,N_13991);
nand U18978 (N_18978,N_11943,N_14569);
nand U18979 (N_18979,N_13056,N_12650);
xnor U18980 (N_18980,N_13739,N_11029);
and U18981 (N_18981,N_13342,N_11010);
nand U18982 (N_18982,N_14008,N_12048);
xnor U18983 (N_18983,N_12670,N_13566);
and U18984 (N_18984,N_10741,N_13250);
and U18985 (N_18985,N_13846,N_10123);
nand U18986 (N_18986,N_13922,N_12822);
nor U18987 (N_18987,N_12421,N_12603);
or U18988 (N_18988,N_10060,N_14584);
xor U18989 (N_18989,N_11332,N_11134);
or U18990 (N_18990,N_10134,N_12993);
or U18991 (N_18991,N_12566,N_11819);
nor U18992 (N_18992,N_13907,N_13921);
xnor U18993 (N_18993,N_11178,N_10563);
nand U18994 (N_18994,N_13121,N_10580);
and U18995 (N_18995,N_10955,N_14891);
xnor U18996 (N_18996,N_14902,N_13400);
or U18997 (N_18997,N_13398,N_10547);
nor U18998 (N_18998,N_13337,N_11143);
nand U18999 (N_18999,N_14499,N_11574);
nor U19000 (N_19000,N_12481,N_13522);
and U19001 (N_19001,N_10310,N_14809);
xor U19002 (N_19002,N_11939,N_11074);
xor U19003 (N_19003,N_12716,N_14505);
or U19004 (N_19004,N_10387,N_12530);
nand U19005 (N_19005,N_12875,N_11938);
nand U19006 (N_19006,N_14425,N_11685);
nor U19007 (N_19007,N_12582,N_10399);
or U19008 (N_19008,N_12150,N_14221);
and U19009 (N_19009,N_10187,N_11172);
xnor U19010 (N_19010,N_14248,N_10140);
or U19011 (N_19011,N_10670,N_14892);
nand U19012 (N_19012,N_14147,N_13410);
nor U19013 (N_19013,N_11032,N_11389);
xor U19014 (N_19014,N_14025,N_11938);
or U19015 (N_19015,N_14392,N_13655);
nor U19016 (N_19016,N_11494,N_10601);
nor U19017 (N_19017,N_14083,N_14793);
xor U19018 (N_19018,N_12163,N_13998);
and U19019 (N_19019,N_14741,N_12881);
nor U19020 (N_19020,N_13253,N_10321);
nor U19021 (N_19021,N_11051,N_11009);
nor U19022 (N_19022,N_12199,N_11717);
nor U19023 (N_19023,N_11337,N_12415);
xor U19024 (N_19024,N_13980,N_10458);
or U19025 (N_19025,N_13935,N_14532);
and U19026 (N_19026,N_11790,N_13731);
and U19027 (N_19027,N_12979,N_10032);
nand U19028 (N_19028,N_12308,N_12413);
xnor U19029 (N_19029,N_14275,N_13440);
or U19030 (N_19030,N_12086,N_12967);
nand U19031 (N_19031,N_14972,N_10417);
or U19032 (N_19032,N_12670,N_14197);
and U19033 (N_19033,N_13680,N_12697);
nor U19034 (N_19034,N_10983,N_10354);
and U19035 (N_19035,N_12699,N_14763);
nand U19036 (N_19036,N_11080,N_11188);
nand U19037 (N_19037,N_13797,N_13877);
or U19038 (N_19038,N_10163,N_14017);
or U19039 (N_19039,N_13216,N_11988);
nand U19040 (N_19040,N_14008,N_11747);
nand U19041 (N_19041,N_10544,N_14435);
nor U19042 (N_19042,N_13545,N_10133);
xor U19043 (N_19043,N_11467,N_13833);
nand U19044 (N_19044,N_12816,N_10358);
or U19045 (N_19045,N_10409,N_12652);
or U19046 (N_19046,N_10810,N_12156);
nand U19047 (N_19047,N_12445,N_14350);
or U19048 (N_19048,N_10601,N_12707);
nand U19049 (N_19049,N_13525,N_12011);
xor U19050 (N_19050,N_13560,N_10221);
xor U19051 (N_19051,N_10827,N_10297);
nor U19052 (N_19052,N_11844,N_11816);
nor U19053 (N_19053,N_14415,N_14148);
and U19054 (N_19054,N_12496,N_12747);
nor U19055 (N_19055,N_10110,N_10015);
nor U19056 (N_19056,N_11339,N_10936);
nor U19057 (N_19057,N_12262,N_13951);
xor U19058 (N_19058,N_14908,N_10928);
nand U19059 (N_19059,N_11097,N_11902);
nor U19060 (N_19060,N_13074,N_14484);
xor U19061 (N_19061,N_13677,N_14011);
nor U19062 (N_19062,N_12157,N_14021);
xor U19063 (N_19063,N_12233,N_10220);
and U19064 (N_19064,N_11434,N_14985);
nand U19065 (N_19065,N_11998,N_13177);
and U19066 (N_19066,N_14791,N_10560);
nand U19067 (N_19067,N_10413,N_11180);
xnor U19068 (N_19068,N_12198,N_12981);
nor U19069 (N_19069,N_10747,N_12690);
nand U19070 (N_19070,N_10338,N_10093);
nand U19071 (N_19071,N_11015,N_11082);
xor U19072 (N_19072,N_13459,N_10184);
and U19073 (N_19073,N_10882,N_11450);
and U19074 (N_19074,N_11510,N_10313);
or U19075 (N_19075,N_12275,N_13403);
xnor U19076 (N_19076,N_10751,N_13496);
xnor U19077 (N_19077,N_10444,N_14895);
nand U19078 (N_19078,N_14711,N_10251);
xnor U19079 (N_19079,N_12618,N_12134);
nor U19080 (N_19080,N_10205,N_14742);
nor U19081 (N_19081,N_12232,N_13925);
xnor U19082 (N_19082,N_10588,N_12660);
or U19083 (N_19083,N_14487,N_12108);
xor U19084 (N_19084,N_10477,N_12906);
and U19085 (N_19085,N_12328,N_10418);
and U19086 (N_19086,N_14089,N_10331);
and U19087 (N_19087,N_12826,N_11861);
nor U19088 (N_19088,N_14707,N_12105);
or U19089 (N_19089,N_12633,N_12640);
xor U19090 (N_19090,N_11373,N_10815);
xnor U19091 (N_19091,N_10486,N_12090);
nor U19092 (N_19092,N_12355,N_10931);
or U19093 (N_19093,N_10085,N_14197);
and U19094 (N_19094,N_14741,N_14826);
or U19095 (N_19095,N_11067,N_10553);
or U19096 (N_19096,N_10958,N_14363);
nand U19097 (N_19097,N_13766,N_10640);
xor U19098 (N_19098,N_10090,N_10222);
xor U19099 (N_19099,N_12571,N_10540);
xor U19100 (N_19100,N_11733,N_12911);
nor U19101 (N_19101,N_11388,N_13729);
and U19102 (N_19102,N_14074,N_14824);
nor U19103 (N_19103,N_14964,N_11391);
xor U19104 (N_19104,N_14432,N_13073);
xor U19105 (N_19105,N_12566,N_14969);
and U19106 (N_19106,N_11667,N_12855);
or U19107 (N_19107,N_13507,N_12832);
and U19108 (N_19108,N_11631,N_13960);
and U19109 (N_19109,N_13220,N_11157);
nand U19110 (N_19110,N_13804,N_11154);
or U19111 (N_19111,N_10025,N_12465);
and U19112 (N_19112,N_11357,N_14225);
nor U19113 (N_19113,N_13957,N_12974);
and U19114 (N_19114,N_14054,N_11398);
nand U19115 (N_19115,N_11024,N_13359);
or U19116 (N_19116,N_12643,N_11228);
xnor U19117 (N_19117,N_10168,N_12049);
nor U19118 (N_19118,N_13414,N_10817);
and U19119 (N_19119,N_13875,N_10806);
nor U19120 (N_19120,N_12119,N_14463);
or U19121 (N_19121,N_14587,N_12806);
and U19122 (N_19122,N_12481,N_13412);
xor U19123 (N_19123,N_14455,N_12342);
nand U19124 (N_19124,N_10469,N_12575);
and U19125 (N_19125,N_11330,N_11646);
xor U19126 (N_19126,N_10833,N_12259);
nor U19127 (N_19127,N_11203,N_13582);
or U19128 (N_19128,N_12485,N_13165);
nand U19129 (N_19129,N_12453,N_14269);
and U19130 (N_19130,N_12242,N_12224);
or U19131 (N_19131,N_10822,N_12404);
or U19132 (N_19132,N_12722,N_12417);
or U19133 (N_19133,N_10488,N_14271);
or U19134 (N_19134,N_10174,N_10040);
nand U19135 (N_19135,N_14603,N_10984);
xnor U19136 (N_19136,N_11092,N_14844);
nor U19137 (N_19137,N_13740,N_12564);
nand U19138 (N_19138,N_13530,N_12054);
xor U19139 (N_19139,N_12729,N_12402);
and U19140 (N_19140,N_11566,N_12766);
and U19141 (N_19141,N_13925,N_14088);
or U19142 (N_19142,N_10714,N_10602);
nor U19143 (N_19143,N_10808,N_11191);
or U19144 (N_19144,N_12932,N_14948);
xnor U19145 (N_19145,N_14271,N_14389);
xnor U19146 (N_19146,N_11603,N_13372);
or U19147 (N_19147,N_11909,N_12044);
nand U19148 (N_19148,N_11937,N_11852);
and U19149 (N_19149,N_12262,N_11418);
xor U19150 (N_19150,N_12883,N_14913);
xor U19151 (N_19151,N_11471,N_13134);
xor U19152 (N_19152,N_13299,N_10886);
or U19153 (N_19153,N_13078,N_12707);
or U19154 (N_19154,N_10526,N_10854);
nor U19155 (N_19155,N_10296,N_11186);
and U19156 (N_19156,N_13765,N_13245);
xor U19157 (N_19157,N_10636,N_12017);
nor U19158 (N_19158,N_14986,N_11993);
and U19159 (N_19159,N_12135,N_10537);
nor U19160 (N_19160,N_10605,N_13169);
or U19161 (N_19161,N_14332,N_10961);
nand U19162 (N_19162,N_13866,N_10573);
and U19163 (N_19163,N_11318,N_10303);
nor U19164 (N_19164,N_13994,N_12983);
or U19165 (N_19165,N_10136,N_14180);
and U19166 (N_19166,N_14042,N_10108);
nor U19167 (N_19167,N_12204,N_14355);
xor U19168 (N_19168,N_10394,N_14412);
nor U19169 (N_19169,N_10730,N_14526);
xnor U19170 (N_19170,N_11804,N_12306);
nor U19171 (N_19171,N_12100,N_11378);
xnor U19172 (N_19172,N_13387,N_13324);
xnor U19173 (N_19173,N_12498,N_11751);
or U19174 (N_19174,N_10038,N_12387);
nor U19175 (N_19175,N_12028,N_12126);
or U19176 (N_19176,N_14920,N_13081);
or U19177 (N_19177,N_13051,N_14176);
xnor U19178 (N_19178,N_12382,N_10258);
xnor U19179 (N_19179,N_12126,N_12419);
and U19180 (N_19180,N_13655,N_13591);
or U19181 (N_19181,N_11135,N_10945);
nor U19182 (N_19182,N_12687,N_13818);
or U19183 (N_19183,N_12053,N_11297);
and U19184 (N_19184,N_11026,N_13967);
or U19185 (N_19185,N_12014,N_14762);
nor U19186 (N_19186,N_13345,N_11485);
nor U19187 (N_19187,N_13906,N_11144);
and U19188 (N_19188,N_11884,N_14578);
or U19189 (N_19189,N_14830,N_13721);
xor U19190 (N_19190,N_12277,N_11919);
nor U19191 (N_19191,N_12302,N_14618);
and U19192 (N_19192,N_11053,N_13673);
and U19193 (N_19193,N_14461,N_10284);
nand U19194 (N_19194,N_14183,N_10939);
and U19195 (N_19195,N_11023,N_11571);
xnor U19196 (N_19196,N_11596,N_14063);
xnor U19197 (N_19197,N_11296,N_12054);
and U19198 (N_19198,N_12766,N_10158);
and U19199 (N_19199,N_13521,N_12291);
or U19200 (N_19200,N_11859,N_12236);
or U19201 (N_19201,N_13002,N_10598);
xor U19202 (N_19202,N_13721,N_12026);
nor U19203 (N_19203,N_13661,N_10019);
or U19204 (N_19204,N_12911,N_11918);
xnor U19205 (N_19205,N_13668,N_10923);
xor U19206 (N_19206,N_10613,N_11849);
and U19207 (N_19207,N_10690,N_13434);
and U19208 (N_19208,N_11250,N_10529);
and U19209 (N_19209,N_11513,N_14222);
and U19210 (N_19210,N_13225,N_10463);
xor U19211 (N_19211,N_12788,N_11299);
or U19212 (N_19212,N_13536,N_14136);
nor U19213 (N_19213,N_11205,N_12680);
xnor U19214 (N_19214,N_10825,N_11234);
or U19215 (N_19215,N_10650,N_10764);
or U19216 (N_19216,N_13190,N_14448);
nor U19217 (N_19217,N_12706,N_11582);
nand U19218 (N_19218,N_13798,N_12409);
or U19219 (N_19219,N_13270,N_11273);
xnor U19220 (N_19220,N_10037,N_13176);
and U19221 (N_19221,N_14850,N_12734);
nand U19222 (N_19222,N_10965,N_10572);
or U19223 (N_19223,N_11877,N_14842);
nand U19224 (N_19224,N_13706,N_12845);
xor U19225 (N_19225,N_11929,N_12601);
nand U19226 (N_19226,N_10545,N_14986);
xor U19227 (N_19227,N_10903,N_12572);
or U19228 (N_19228,N_14189,N_13926);
xor U19229 (N_19229,N_12297,N_10561);
xnor U19230 (N_19230,N_11494,N_14982);
nor U19231 (N_19231,N_13855,N_12259);
and U19232 (N_19232,N_12471,N_10844);
nand U19233 (N_19233,N_10678,N_10395);
nor U19234 (N_19234,N_11294,N_12744);
and U19235 (N_19235,N_13753,N_11833);
nand U19236 (N_19236,N_13780,N_10819);
or U19237 (N_19237,N_10950,N_10086);
nand U19238 (N_19238,N_12256,N_11452);
and U19239 (N_19239,N_12493,N_13073);
nor U19240 (N_19240,N_14642,N_14277);
nor U19241 (N_19241,N_11368,N_11153);
and U19242 (N_19242,N_11165,N_14272);
and U19243 (N_19243,N_14801,N_11073);
nor U19244 (N_19244,N_13165,N_12545);
or U19245 (N_19245,N_14697,N_11628);
and U19246 (N_19246,N_11061,N_12692);
or U19247 (N_19247,N_12597,N_12246);
and U19248 (N_19248,N_11119,N_14369);
nor U19249 (N_19249,N_11716,N_14174);
or U19250 (N_19250,N_13863,N_12443);
nand U19251 (N_19251,N_13575,N_10261);
nor U19252 (N_19252,N_11489,N_12754);
or U19253 (N_19253,N_12261,N_13452);
and U19254 (N_19254,N_12942,N_14649);
nand U19255 (N_19255,N_11925,N_12420);
xor U19256 (N_19256,N_10467,N_11171);
nor U19257 (N_19257,N_13835,N_12938);
and U19258 (N_19258,N_11584,N_11970);
xnor U19259 (N_19259,N_11768,N_13310);
nor U19260 (N_19260,N_11876,N_13801);
nand U19261 (N_19261,N_11302,N_14292);
or U19262 (N_19262,N_10934,N_11876);
xor U19263 (N_19263,N_10348,N_12767);
nor U19264 (N_19264,N_13659,N_13372);
or U19265 (N_19265,N_12377,N_10411);
xnor U19266 (N_19266,N_11820,N_14297);
or U19267 (N_19267,N_12735,N_10859);
and U19268 (N_19268,N_11110,N_12413);
xnor U19269 (N_19269,N_11847,N_14745);
xor U19270 (N_19270,N_12358,N_13573);
and U19271 (N_19271,N_12244,N_13564);
nand U19272 (N_19272,N_11726,N_14692);
or U19273 (N_19273,N_12853,N_14909);
nor U19274 (N_19274,N_13115,N_14815);
or U19275 (N_19275,N_13515,N_14524);
xor U19276 (N_19276,N_10913,N_14628);
xor U19277 (N_19277,N_14554,N_13152);
and U19278 (N_19278,N_12048,N_12467);
nor U19279 (N_19279,N_10017,N_10331);
nand U19280 (N_19280,N_12426,N_13744);
nor U19281 (N_19281,N_14988,N_14887);
or U19282 (N_19282,N_12356,N_11778);
nand U19283 (N_19283,N_11800,N_10064);
nor U19284 (N_19284,N_11579,N_12967);
nor U19285 (N_19285,N_11704,N_10378);
nor U19286 (N_19286,N_12942,N_12356);
and U19287 (N_19287,N_13942,N_11103);
nand U19288 (N_19288,N_14555,N_12631);
or U19289 (N_19289,N_14313,N_10718);
nor U19290 (N_19290,N_10910,N_14768);
nor U19291 (N_19291,N_13635,N_13369);
nor U19292 (N_19292,N_11276,N_10618);
xor U19293 (N_19293,N_14420,N_11048);
and U19294 (N_19294,N_12549,N_14168);
nand U19295 (N_19295,N_12385,N_10987);
and U19296 (N_19296,N_12014,N_12762);
and U19297 (N_19297,N_11832,N_10756);
nand U19298 (N_19298,N_13261,N_14265);
or U19299 (N_19299,N_13576,N_10326);
and U19300 (N_19300,N_12082,N_13190);
nand U19301 (N_19301,N_11022,N_11457);
nand U19302 (N_19302,N_13313,N_11474);
xnor U19303 (N_19303,N_11022,N_14324);
xor U19304 (N_19304,N_14195,N_11586);
or U19305 (N_19305,N_12423,N_11966);
nand U19306 (N_19306,N_10826,N_11781);
or U19307 (N_19307,N_11883,N_13043);
nor U19308 (N_19308,N_13849,N_13761);
nand U19309 (N_19309,N_13160,N_13009);
nand U19310 (N_19310,N_13984,N_10312);
and U19311 (N_19311,N_14699,N_11926);
nor U19312 (N_19312,N_10429,N_10492);
and U19313 (N_19313,N_14240,N_13168);
or U19314 (N_19314,N_12911,N_13681);
nor U19315 (N_19315,N_10229,N_12771);
xor U19316 (N_19316,N_10325,N_14875);
nand U19317 (N_19317,N_13367,N_10628);
nand U19318 (N_19318,N_11573,N_14463);
nand U19319 (N_19319,N_10075,N_10280);
xor U19320 (N_19320,N_11824,N_13118);
nor U19321 (N_19321,N_11460,N_12782);
nand U19322 (N_19322,N_14344,N_13998);
or U19323 (N_19323,N_14417,N_11448);
and U19324 (N_19324,N_13566,N_14044);
xnor U19325 (N_19325,N_10526,N_13609);
nor U19326 (N_19326,N_11441,N_14334);
or U19327 (N_19327,N_12166,N_12659);
or U19328 (N_19328,N_13786,N_12805);
or U19329 (N_19329,N_11499,N_14065);
xor U19330 (N_19330,N_10105,N_12607);
or U19331 (N_19331,N_14252,N_14540);
or U19332 (N_19332,N_13045,N_13705);
and U19333 (N_19333,N_10142,N_10288);
and U19334 (N_19334,N_12476,N_13119);
and U19335 (N_19335,N_10351,N_11230);
or U19336 (N_19336,N_13490,N_13589);
nand U19337 (N_19337,N_10663,N_13170);
and U19338 (N_19338,N_13016,N_10580);
or U19339 (N_19339,N_12787,N_14112);
or U19340 (N_19340,N_13204,N_10522);
nor U19341 (N_19341,N_14972,N_10676);
and U19342 (N_19342,N_13531,N_12310);
nor U19343 (N_19343,N_14386,N_10239);
or U19344 (N_19344,N_10267,N_10953);
or U19345 (N_19345,N_11054,N_13644);
nand U19346 (N_19346,N_10224,N_14249);
nor U19347 (N_19347,N_12430,N_12688);
nor U19348 (N_19348,N_11235,N_10226);
xor U19349 (N_19349,N_13256,N_13694);
and U19350 (N_19350,N_10924,N_12867);
or U19351 (N_19351,N_14286,N_14143);
nand U19352 (N_19352,N_12163,N_10195);
and U19353 (N_19353,N_14403,N_11765);
xor U19354 (N_19354,N_11460,N_14769);
and U19355 (N_19355,N_14757,N_13005);
or U19356 (N_19356,N_11602,N_13011);
nor U19357 (N_19357,N_13903,N_14977);
nor U19358 (N_19358,N_12885,N_12606);
and U19359 (N_19359,N_10259,N_11707);
or U19360 (N_19360,N_10933,N_12702);
nand U19361 (N_19361,N_11002,N_13131);
nor U19362 (N_19362,N_12083,N_13001);
nand U19363 (N_19363,N_12791,N_10037);
nor U19364 (N_19364,N_14649,N_14187);
xor U19365 (N_19365,N_12489,N_13647);
xnor U19366 (N_19366,N_11896,N_10344);
and U19367 (N_19367,N_11807,N_10378);
or U19368 (N_19368,N_13235,N_14216);
xor U19369 (N_19369,N_11187,N_11193);
or U19370 (N_19370,N_11381,N_10177);
and U19371 (N_19371,N_13828,N_11879);
or U19372 (N_19372,N_10380,N_11623);
nand U19373 (N_19373,N_13602,N_10147);
nor U19374 (N_19374,N_11851,N_11516);
and U19375 (N_19375,N_11452,N_13417);
nand U19376 (N_19376,N_12701,N_10988);
and U19377 (N_19377,N_14297,N_11605);
and U19378 (N_19378,N_13422,N_12763);
nor U19379 (N_19379,N_13203,N_14856);
nor U19380 (N_19380,N_10906,N_13402);
nand U19381 (N_19381,N_14493,N_12316);
or U19382 (N_19382,N_13614,N_13480);
nor U19383 (N_19383,N_10489,N_11107);
nor U19384 (N_19384,N_13992,N_10200);
nor U19385 (N_19385,N_12317,N_11438);
or U19386 (N_19386,N_12679,N_12021);
and U19387 (N_19387,N_14370,N_14632);
or U19388 (N_19388,N_13377,N_10481);
xnor U19389 (N_19389,N_10921,N_11592);
and U19390 (N_19390,N_14444,N_11046);
or U19391 (N_19391,N_10566,N_11876);
nand U19392 (N_19392,N_12223,N_11056);
nand U19393 (N_19393,N_11512,N_12818);
nand U19394 (N_19394,N_12835,N_11539);
xor U19395 (N_19395,N_12533,N_12346);
xnor U19396 (N_19396,N_10138,N_12311);
or U19397 (N_19397,N_14837,N_10945);
or U19398 (N_19398,N_11042,N_11241);
or U19399 (N_19399,N_10359,N_14547);
and U19400 (N_19400,N_12818,N_14023);
and U19401 (N_19401,N_13529,N_11298);
and U19402 (N_19402,N_11638,N_14375);
xnor U19403 (N_19403,N_10015,N_14803);
or U19404 (N_19404,N_11349,N_14076);
and U19405 (N_19405,N_14962,N_14890);
or U19406 (N_19406,N_10883,N_14619);
xor U19407 (N_19407,N_11590,N_13906);
or U19408 (N_19408,N_14299,N_14609);
or U19409 (N_19409,N_11635,N_12908);
xor U19410 (N_19410,N_12092,N_11527);
nor U19411 (N_19411,N_13544,N_13914);
nor U19412 (N_19412,N_13241,N_12640);
or U19413 (N_19413,N_14547,N_12828);
xnor U19414 (N_19414,N_12469,N_13572);
nand U19415 (N_19415,N_11824,N_10834);
xor U19416 (N_19416,N_11052,N_13677);
xnor U19417 (N_19417,N_14202,N_10267);
nor U19418 (N_19418,N_10296,N_11064);
and U19419 (N_19419,N_12303,N_11368);
nor U19420 (N_19420,N_14194,N_14164);
and U19421 (N_19421,N_14093,N_14530);
xor U19422 (N_19422,N_13782,N_13062);
nor U19423 (N_19423,N_10493,N_10726);
nor U19424 (N_19424,N_10624,N_11213);
xnor U19425 (N_19425,N_10787,N_11610);
nor U19426 (N_19426,N_12634,N_10298);
or U19427 (N_19427,N_11047,N_13868);
xor U19428 (N_19428,N_10087,N_11141);
nor U19429 (N_19429,N_11842,N_13804);
nand U19430 (N_19430,N_13893,N_14806);
xnor U19431 (N_19431,N_10469,N_11966);
xor U19432 (N_19432,N_13578,N_12955);
and U19433 (N_19433,N_10950,N_10284);
xnor U19434 (N_19434,N_11578,N_11161);
and U19435 (N_19435,N_13566,N_12688);
or U19436 (N_19436,N_12629,N_10979);
nor U19437 (N_19437,N_13356,N_11003);
nor U19438 (N_19438,N_10146,N_13311);
nand U19439 (N_19439,N_10927,N_14690);
nor U19440 (N_19440,N_10624,N_12879);
nor U19441 (N_19441,N_12292,N_10030);
nor U19442 (N_19442,N_10246,N_13432);
nand U19443 (N_19443,N_14060,N_14338);
and U19444 (N_19444,N_11284,N_10811);
nand U19445 (N_19445,N_10444,N_11395);
or U19446 (N_19446,N_13043,N_11760);
nor U19447 (N_19447,N_12007,N_11912);
or U19448 (N_19448,N_14011,N_13035);
nand U19449 (N_19449,N_11385,N_12251);
or U19450 (N_19450,N_12363,N_11566);
or U19451 (N_19451,N_14925,N_11803);
or U19452 (N_19452,N_10200,N_11636);
nand U19453 (N_19453,N_11174,N_12398);
nor U19454 (N_19454,N_10425,N_11283);
xor U19455 (N_19455,N_12459,N_11718);
nor U19456 (N_19456,N_11989,N_14449);
and U19457 (N_19457,N_13705,N_11267);
nor U19458 (N_19458,N_11914,N_14203);
and U19459 (N_19459,N_13495,N_10971);
nand U19460 (N_19460,N_12915,N_10750);
nor U19461 (N_19461,N_10428,N_14940);
and U19462 (N_19462,N_10513,N_11979);
xor U19463 (N_19463,N_12429,N_11991);
nand U19464 (N_19464,N_11781,N_10587);
and U19465 (N_19465,N_11999,N_11777);
and U19466 (N_19466,N_12418,N_13027);
xnor U19467 (N_19467,N_13135,N_13328);
or U19468 (N_19468,N_14261,N_11347);
or U19469 (N_19469,N_13741,N_10436);
or U19470 (N_19470,N_11323,N_14853);
nand U19471 (N_19471,N_12132,N_10882);
or U19472 (N_19472,N_14001,N_13478);
nor U19473 (N_19473,N_13807,N_11514);
and U19474 (N_19474,N_10422,N_10018);
nand U19475 (N_19475,N_10761,N_13394);
and U19476 (N_19476,N_12951,N_13051);
or U19477 (N_19477,N_14359,N_12665);
nand U19478 (N_19478,N_10735,N_10397);
nor U19479 (N_19479,N_10811,N_13052);
or U19480 (N_19480,N_14035,N_13658);
nor U19481 (N_19481,N_11395,N_12103);
xnor U19482 (N_19482,N_10463,N_10040);
nand U19483 (N_19483,N_14910,N_13917);
nor U19484 (N_19484,N_12735,N_13953);
or U19485 (N_19485,N_14699,N_12400);
and U19486 (N_19486,N_12993,N_14302);
xnor U19487 (N_19487,N_11716,N_11574);
nand U19488 (N_19488,N_11305,N_14900);
nor U19489 (N_19489,N_13887,N_14060);
or U19490 (N_19490,N_11737,N_10093);
and U19491 (N_19491,N_13705,N_13179);
and U19492 (N_19492,N_12664,N_13936);
xor U19493 (N_19493,N_12820,N_12199);
nand U19494 (N_19494,N_13630,N_14679);
or U19495 (N_19495,N_11333,N_10566);
nor U19496 (N_19496,N_11691,N_14074);
nor U19497 (N_19497,N_11743,N_11609);
nand U19498 (N_19498,N_13372,N_12578);
and U19499 (N_19499,N_12115,N_12604);
or U19500 (N_19500,N_14643,N_12679);
or U19501 (N_19501,N_12327,N_11333);
or U19502 (N_19502,N_14610,N_13177);
nor U19503 (N_19503,N_12469,N_13672);
nand U19504 (N_19504,N_14202,N_10495);
nand U19505 (N_19505,N_11578,N_14639);
or U19506 (N_19506,N_10136,N_14967);
xnor U19507 (N_19507,N_11361,N_12246);
nand U19508 (N_19508,N_11447,N_12432);
nor U19509 (N_19509,N_14726,N_14702);
nor U19510 (N_19510,N_14538,N_10157);
nand U19511 (N_19511,N_12621,N_10498);
nand U19512 (N_19512,N_13970,N_10920);
xor U19513 (N_19513,N_13453,N_13793);
or U19514 (N_19514,N_14002,N_11008);
nor U19515 (N_19515,N_10743,N_13922);
xor U19516 (N_19516,N_12840,N_13668);
or U19517 (N_19517,N_11748,N_10584);
and U19518 (N_19518,N_12624,N_14682);
nor U19519 (N_19519,N_10259,N_10949);
or U19520 (N_19520,N_10414,N_13987);
and U19521 (N_19521,N_12863,N_13061);
or U19522 (N_19522,N_14677,N_13487);
nand U19523 (N_19523,N_13889,N_11789);
and U19524 (N_19524,N_13870,N_13157);
xor U19525 (N_19525,N_10027,N_12620);
nor U19526 (N_19526,N_14776,N_14789);
nand U19527 (N_19527,N_14757,N_13347);
nand U19528 (N_19528,N_11374,N_10808);
xnor U19529 (N_19529,N_13700,N_13390);
and U19530 (N_19530,N_11422,N_10596);
or U19531 (N_19531,N_11368,N_10246);
xnor U19532 (N_19532,N_13406,N_12505);
and U19533 (N_19533,N_11890,N_13769);
or U19534 (N_19534,N_12661,N_13319);
nand U19535 (N_19535,N_14129,N_11167);
and U19536 (N_19536,N_12338,N_14660);
nand U19537 (N_19537,N_11703,N_11617);
or U19538 (N_19538,N_14545,N_13911);
xor U19539 (N_19539,N_12174,N_11021);
xnor U19540 (N_19540,N_11226,N_13421);
or U19541 (N_19541,N_12900,N_14115);
nor U19542 (N_19542,N_14735,N_14023);
and U19543 (N_19543,N_13646,N_14127);
and U19544 (N_19544,N_12944,N_13437);
nand U19545 (N_19545,N_11614,N_14394);
nor U19546 (N_19546,N_10253,N_10684);
xnor U19547 (N_19547,N_14517,N_14822);
or U19548 (N_19548,N_12080,N_14553);
nand U19549 (N_19549,N_12533,N_10601);
nor U19550 (N_19550,N_10792,N_11100);
xnor U19551 (N_19551,N_13336,N_12389);
nand U19552 (N_19552,N_10946,N_10642);
or U19553 (N_19553,N_13655,N_12432);
or U19554 (N_19554,N_10703,N_10162);
xnor U19555 (N_19555,N_10822,N_14873);
nand U19556 (N_19556,N_13065,N_12062);
xor U19557 (N_19557,N_11180,N_14370);
or U19558 (N_19558,N_12412,N_14664);
or U19559 (N_19559,N_14619,N_14361);
and U19560 (N_19560,N_11298,N_12512);
xnor U19561 (N_19561,N_10947,N_12541);
or U19562 (N_19562,N_14591,N_10087);
nand U19563 (N_19563,N_11200,N_12533);
or U19564 (N_19564,N_14861,N_14958);
xnor U19565 (N_19565,N_12681,N_14462);
nor U19566 (N_19566,N_13684,N_10379);
nor U19567 (N_19567,N_11027,N_10924);
nand U19568 (N_19568,N_13402,N_14608);
nor U19569 (N_19569,N_14781,N_13474);
or U19570 (N_19570,N_11811,N_14752);
nor U19571 (N_19571,N_12039,N_10566);
nand U19572 (N_19572,N_13475,N_13042);
xnor U19573 (N_19573,N_13967,N_11438);
nand U19574 (N_19574,N_14132,N_13015);
or U19575 (N_19575,N_11655,N_11692);
and U19576 (N_19576,N_11517,N_13520);
or U19577 (N_19577,N_11283,N_13182);
and U19578 (N_19578,N_11287,N_12071);
nand U19579 (N_19579,N_10036,N_14813);
and U19580 (N_19580,N_13365,N_10250);
xor U19581 (N_19581,N_11937,N_11601);
and U19582 (N_19582,N_12049,N_14952);
xor U19583 (N_19583,N_13875,N_11234);
nor U19584 (N_19584,N_12776,N_12852);
nand U19585 (N_19585,N_10675,N_12816);
xor U19586 (N_19586,N_13966,N_10368);
xnor U19587 (N_19587,N_12468,N_11035);
or U19588 (N_19588,N_11219,N_13247);
nor U19589 (N_19589,N_12381,N_13269);
and U19590 (N_19590,N_14017,N_12322);
xor U19591 (N_19591,N_11048,N_13716);
and U19592 (N_19592,N_12494,N_12456);
and U19593 (N_19593,N_10629,N_12563);
nor U19594 (N_19594,N_12528,N_11672);
or U19595 (N_19595,N_10385,N_13490);
or U19596 (N_19596,N_12994,N_12614);
nand U19597 (N_19597,N_10604,N_14021);
nor U19598 (N_19598,N_12852,N_12594);
and U19599 (N_19599,N_13846,N_10793);
nand U19600 (N_19600,N_12695,N_12520);
nor U19601 (N_19601,N_10918,N_10624);
and U19602 (N_19602,N_13119,N_13935);
xor U19603 (N_19603,N_10022,N_12138);
and U19604 (N_19604,N_13049,N_14074);
and U19605 (N_19605,N_13239,N_14427);
or U19606 (N_19606,N_13171,N_11295);
nor U19607 (N_19607,N_14960,N_10620);
nor U19608 (N_19608,N_12083,N_13092);
nand U19609 (N_19609,N_12914,N_14930);
nor U19610 (N_19610,N_14179,N_10548);
xnor U19611 (N_19611,N_12327,N_10822);
nand U19612 (N_19612,N_13352,N_14226);
xnor U19613 (N_19613,N_13301,N_12451);
or U19614 (N_19614,N_11617,N_12670);
and U19615 (N_19615,N_10894,N_10473);
or U19616 (N_19616,N_13991,N_14092);
xor U19617 (N_19617,N_14012,N_14639);
or U19618 (N_19618,N_14502,N_11796);
nand U19619 (N_19619,N_14500,N_10770);
or U19620 (N_19620,N_11156,N_13987);
nand U19621 (N_19621,N_12342,N_10556);
nand U19622 (N_19622,N_10854,N_13921);
nand U19623 (N_19623,N_12932,N_13008);
nand U19624 (N_19624,N_11604,N_14798);
xnor U19625 (N_19625,N_11038,N_11259);
and U19626 (N_19626,N_13426,N_12189);
or U19627 (N_19627,N_12490,N_14270);
nor U19628 (N_19628,N_12272,N_14864);
xor U19629 (N_19629,N_12659,N_12480);
or U19630 (N_19630,N_11243,N_13549);
or U19631 (N_19631,N_11150,N_13747);
xnor U19632 (N_19632,N_11698,N_12623);
xor U19633 (N_19633,N_12135,N_11618);
or U19634 (N_19634,N_11550,N_11604);
and U19635 (N_19635,N_14569,N_12670);
nand U19636 (N_19636,N_13654,N_11055);
or U19637 (N_19637,N_11036,N_10836);
and U19638 (N_19638,N_11502,N_10810);
xor U19639 (N_19639,N_13442,N_11967);
or U19640 (N_19640,N_11560,N_14288);
nor U19641 (N_19641,N_10166,N_14031);
or U19642 (N_19642,N_14616,N_10373);
xor U19643 (N_19643,N_11034,N_12736);
nor U19644 (N_19644,N_10812,N_10980);
xor U19645 (N_19645,N_14238,N_13851);
or U19646 (N_19646,N_11837,N_10134);
or U19647 (N_19647,N_11432,N_10602);
xor U19648 (N_19648,N_12678,N_12548);
nor U19649 (N_19649,N_10692,N_12996);
nor U19650 (N_19650,N_11871,N_11175);
and U19651 (N_19651,N_11035,N_11421);
nand U19652 (N_19652,N_13568,N_12235);
and U19653 (N_19653,N_13284,N_11014);
nand U19654 (N_19654,N_14354,N_12592);
nor U19655 (N_19655,N_10377,N_10653);
nor U19656 (N_19656,N_10240,N_14871);
xnor U19657 (N_19657,N_14361,N_13946);
xor U19658 (N_19658,N_12799,N_11887);
or U19659 (N_19659,N_10496,N_11666);
nor U19660 (N_19660,N_10480,N_11390);
and U19661 (N_19661,N_10894,N_12050);
xor U19662 (N_19662,N_10095,N_10763);
or U19663 (N_19663,N_14366,N_12818);
nor U19664 (N_19664,N_14313,N_13505);
or U19665 (N_19665,N_11333,N_14881);
nor U19666 (N_19666,N_12320,N_10427);
and U19667 (N_19667,N_14438,N_13274);
nand U19668 (N_19668,N_12496,N_14982);
xnor U19669 (N_19669,N_11953,N_14671);
or U19670 (N_19670,N_14392,N_13540);
nand U19671 (N_19671,N_14814,N_10029);
and U19672 (N_19672,N_14921,N_10252);
or U19673 (N_19673,N_14080,N_10051);
and U19674 (N_19674,N_13307,N_14249);
and U19675 (N_19675,N_10261,N_13195);
nand U19676 (N_19676,N_11625,N_12570);
or U19677 (N_19677,N_11139,N_10230);
nor U19678 (N_19678,N_14241,N_12460);
nor U19679 (N_19679,N_10989,N_13412);
xor U19680 (N_19680,N_10129,N_13734);
or U19681 (N_19681,N_11354,N_14964);
or U19682 (N_19682,N_11369,N_12250);
nor U19683 (N_19683,N_11234,N_11380);
or U19684 (N_19684,N_12701,N_14015);
xor U19685 (N_19685,N_14217,N_14074);
xor U19686 (N_19686,N_11276,N_10520);
xor U19687 (N_19687,N_10383,N_11211);
nor U19688 (N_19688,N_12135,N_13837);
and U19689 (N_19689,N_13947,N_14411);
nand U19690 (N_19690,N_14292,N_10132);
xor U19691 (N_19691,N_12562,N_13718);
and U19692 (N_19692,N_13883,N_13677);
nor U19693 (N_19693,N_14984,N_10765);
xor U19694 (N_19694,N_10715,N_10785);
and U19695 (N_19695,N_14308,N_10458);
or U19696 (N_19696,N_11557,N_11677);
xnor U19697 (N_19697,N_10130,N_11707);
xnor U19698 (N_19698,N_14668,N_10838);
or U19699 (N_19699,N_10663,N_12865);
nand U19700 (N_19700,N_11065,N_10230);
nor U19701 (N_19701,N_10575,N_10235);
or U19702 (N_19702,N_12056,N_10011);
nand U19703 (N_19703,N_10355,N_10888);
and U19704 (N_19704,N_10448,N_11384);
and U19705 (N_19705,N_14034,N_11888);
xor U19706 (N_19706,N_11519,N_13388);
nor U19707 (N_19707,N_13490,N_12646);
nor U19708 (N_19708,N_14146,N_11548);
nor U19709 (N_19709,N_14070,N_12494);
xnor U19710 (N_19710,N_14989,N_11610);
and U19711 (N_19711,N_13522,N_12637);
nand U19712 (N_19712,N_12194,N_11954);
or U19713 (N_19713,N_12832,N_14646);
nand U19714 (N_19714,N_11633,N_11706);
or U19715 (N_19715,N_10389,N_11789);
and U19716 (N_19716,N_11913,N_11848);
and U19717 (N_19717,N_13047,N_13342);
nand U19718 (N_19718,N_10897,N_13020);
and U19719 (N_19719,N_11470,N_10510);
nand U19720 (N_19720,N_13939,N_12147);
or U19721 (N_19721,N_14046,N_13807);
nand U19722 (N_19722,N_12399,N_13220);
nor U19723 (N_19723,N_13598,N_10391);
or U19724 (N_19724,N_12164,N_12744);
xnor U19725 (N_19725,N_14640,N_14812);
or U19726 (N_19726,N_11236,N_12390);
nand U19727 (N_19727,N_13724,N_14686);
or U19728 (N_19728,N_12833,N_12445);
or U19729 (N_19729,N_11040,N_11582);
nor U19730 (N_19730,N_14351,N_12267);
xor U19731 (N_19731,N_11097,N_13797);
xnor U19732 (N_19732,N_11244,N_14224);
nor U19733 (N_19733,N_10655,N_11946);
and U19734 (N_19734,N_13175,N_11059);
xor U19735 (N_19735,N_12119,N_13030);
or U19736 (N_19736,N_11161,N_13328);
nor U19737 (N_19737,N_14597,N_13803);
and U19738 (N_19738,N_10150,N_13662);
nand U19739 (N_19739,N_13333,N_11613);
xnor U19740 (N_19740,N_12778,N_10135);
or U19741 (N_19741,N_14600,N_14368);
or U19742 (N_19742,N_12018,N_11407);
or U19743 (N_19743,N_11621,N_14985);
nand U19744 (N_19744,N_13476,N_10977);
or U19745 (N_19745,N_10574,N_12529);
nand U19746 (N_19746,N_10444,N_11218);
nor U19747 (N_19747,N_11603,N_13977);
nor U19748 (N_19748,N_13650,N_10966);
or U19749 (N_19749,N_13069,N_10408);
nand U19750 (N_19750,N_13420,N_11043);
or U19751 (N_19751,N_12867,N_11677);
nor U19752 (N_19752,N_10626,N_14349);
xnor U19753 (N_19753,N_10120,N_13461);
or U19754 (N_19754,N_11904,N_12895);
xor U19755 (N_19755,N_10988,N_11528);
or U19756 (N_19756,N_12943,N_11359);
xnor U19757 (N_19757,N_14264,N_14648);
xnor U19758 (N_19758,N_13540,N_13440);
and U19759 (N_19759,N_10337,N_11631);
nand U19760 (N_19760,N_14361,N_14515);
xor U19761 (N_19761,N_12548,N_12358);
or U19762 (N_19762,N_11986,N_12202);
and U19763 (N_19763,N_14363,N_11520);
or U19764 (N_19764,N_13834,N_14555);
or U19765 (N_19765,N_10720,N_14876);
and U19766 (N_19766,N_13367,N_11963);
or U19767 (N_19767,N_10514,N_10671);
xnor U19768 (N_19768,N_10955,N_12157);
xnor U19769 (N_19769,N_11848,N_12893);
or U19770 (N_19770,N_11581,N_11053);
or U19771 (N_19771,N_11671,N_11840);
nor U19772 (N_19772,N_10430,N_12393);
nand U19773 (N_19773,N_12736,N_11914);
xor U19774 (N_19774,N_11294,N_13547);
xor U19775 (N_19775,N_10099,N_14354);
xnor U19776 (N_19776,N_11930,N_12908);
xor U19777 (N_19777,N_13820,N_12156);
and U19778 (N_19778,N_12461,N_13332);
or U19779 (N_19779,N_14529,N_10712);
and U19780 (N_19780,N_12140,N_13426);
nor U19781 (N_19781,N_11285,N_10711);
nand U19782 (N_19782,N_13367,N_12151);
nor U19783 (N_19783,N_11101,N_10701);
xnor U19784 (N_19784,N_14118,N_11173);
and U19785 (N_19785,N_10804,N_13260);
nor U19786 (N_19786,N_13075,N_13738);
and U19787 (N_19787,N_13827,N_11849);
nor U19788 (N_19788,N_12532,N_10355);
nand U19789 (N_19789,N_11310,N_14383);
nor U19790 (N_19790,N_13711,N_10419);
nor U19791 (N_19791,N_11149,N_13596);
nand U19792 (N_19792,N_13876,N_10836);
xnor U19793 (N_19793,N_13497,N_13820);
nor U19794 (N_19794,N_13797,N_14756);
and U19795 (N_19795,N_11375,N_13870);
or U19796 (N_19796,N_13645,N_12794);
xnor U19797 (N_19797,N_10603,N_14839);
nor U19798 (N_19798,N_14733,N_10891);
or U19799 (N_19799,N_11664,N_13161);
and U19800 (N_19800,N_14848,N_10497);
xor U19801 (N_19801,N_11152,N_12547);
nor U19802 (N_19802,N_10750,N_10094);
nor U19803 (N_19803,N_13031,N_13486);
or U19804 (N_19804,N_11152,N_10230);
or U19805 (N_19805,N_11336,N_10201);
nand U19806 (N_19806,N_13176,N_12012);
nor U19807 (N_19807,N_10840,N_10928);
nor U19808 (N_19808,N_11346,N_11018);
xor U19809 (N_19809,N_12671,N_10970);
nand U19810 (N_19810,N_12599,N_11674);
and U19811 (N_19811,N_12333,N_14354);
or U19812 (N_19812,N_13864,N_10644);
or U19813 (N_19813,N_13095,N_13828);
or U19814 (N_19814,N_14940,N_14006);
or U19815 (N_19815,N_14514,N_14457);
xor U19816 (N_19816,N_11811,N_14400);
and U19817 (N_19817,N_10726,N_14012);
xnor U19818 (N_19818,N_13091,N_13621);
or U19819 (N_19819,N_14985,N_14137);
and U19820 (N_19820,N_12543,N_12964);
and U19821 (N_19821,N_10246,N_13610);
and U19822 (N_19822,N_12525,N_11546);
and U19823 (N_19823,N_10251,N_12898);
xor U19824 (N_19824,N_12501,N_10293);
nor U19825 (N_19825,N_10241,N_12805);
or U19826 (N_19826,N_12297,N_14728);
nor U19827 (N_19827,N_14422,N_13580);
or U19828 (N_19828,N_11100,N_10777);
xor U19829 (N_19829,N_14214,N_13012);
xnor U19830 (N_19830,N_10563,N_10245);
nand U19831 (N_19831,N_13773,N_12997);
and U19832 (N_19832,N_13108,N_12676);
nor U19833 (N_19833,N_11284,N_14218);
nand U19834 (N_19834,N_10072,N_13384);
xnor U19835 (N_19835,N_11765,N_10207);
or U19836 (N_19836,N_11891,N_10427);
nand U19837 (N_19837,N_13683,N_12309);
nand U19838 (N_19838,N_12172,N_11374);
xnor U19839 (N_19839,N_13443,N_12658);
nand U19840 (N_19840,N_14586,N_13996);
nor U19841 (N_19841,N_12622,N_12548);
nand U19842 (N_19842,N_10049,N_14415);
xor U19843 (N_19843,N_12615,N_10996);
and U19844 (N_19844,N_11344,N_10129);
xnor U19845 (N_19845,N_12304,N_14611);
or U19846 (N_19846,N_11725,N_11766);
or U19847 (N_19847,N_13192,N_11550);
nand U19848 (N_19848,N_14958,N_10897);
nand U19849 (N_19849,N_14963,N_13881);
nand U19850 (N_19850,N_14876,N_10418);
nand U19851 (N_19851,N_10977,N_12982);
nor U19852 (N_19852,N_14965,N_14576);
nand U19853 (N_19853,N_13475,N_13069);
nand U19854 (N_19854,N_14660,N_13036);
and U19855 (N_19855,N_14311,N_14098);
or U19856 (N_19856,N_10794,N_10860);
or U19857 (N_19857,N_14530,N_12386);
or U19858 (N_19858,N_14912,N_13929);
nand U19859 (N_19859,N_13634,N_10719);
and U19860 (N_19860,N_10483,N_13615);
nor U19861 (N_19861,N_13079,N_11602);
nor U19862 (N_19862,N_10378,N_14307);
xor U19863 (N_19863,N_10316,N_11728);
nor U19864 (N_19864,N_10561,N_10909);
nor U19865 (N_19865,N_12242,N_10922);
and U19866 (N_19866,N_11775,N_12900);
and U19867 (N_19867,N_13932,N_14724);
nor U19868 (N_19868,N_11943,N_11621);
nor U19869 (N_19869,N_13272,N_11825);
or U19870 (N_19870,N_11013,N_11638);
xnor U19871 (N_19871,N_11102,N_13213);
nand U19872 (N_19872,N_11621,N_14603);
and U19873 (N_19873,N_13201,N_10307);
and U19874 (N_19874,N_12886,N_12796);
xnor U19875 (N_19875,N_14705,N_12345);
nand U19876 (N_19876,N_14361,N_13038);
and U19877 (N_19877,N_10424,N_13484);
xor U19878 (N_19878,N_10399,N_14067);
xor U19879 (N_19879,N_14102,N_12038);
nand U19880 (N_19880,N_12979,N_14227);
nor U19881 (N_19881,N_14197,N_13978);
nand U19882 (N_19882,N_13237,N_14820);
and U19883 (N_19883,N_10235,N_11404);
or U19884 (N_19884,N_10623,N_12255);
nor U19885 (N_19885,N_13481,N_12959);
xnor U19886 (N_19886,N_12491,N_13850);
and U19887 (N_19887,N_10812,N_12947);
nor U19888 (N_19888,N_11706,N_11055);
nor U19889 (N_19889,N_11915,N_13999);
or U19890 (N_19890,N_11070,N_12498);
nand U19891 (N_19891,N_12271,N_12729);
and U19892 (N_19892,N_12802,N_10838);
and U19893 (N_19893,N_11625,N_13421);
nor U19894 (N_19894,N_13158,N_12049);
nor U19895 (N_19895,N_14196,N_14250);
xnor U19896 (N_19896,N_11214,N_11712);
and U19897 (N_19897,N_13014,N_12707);
and U19898 (N_19898,N_13012,N_12161);
xnor U19899 (N_19899,N_11254,N_11485);
and U19900 (N_19900,N_13068,N_14677);
xnor U19901 (N_19901,N_10467,N_12750);
xnor U19902 (N_19902,N_13983,N_12760);
nand U19903 (N_19903,N_14178,N_11214);
and U19904 (N_19904,N_10922,N_10949);
nor U19905 (N_19905,N_13259,N_11505);
nand U19906 (N_19906,N_10924,N_14753);
and U19907 (N_19907,N_11874,N_12832);
nand U19908 (N_19908,N_11161,N_11728);
or U19909 (N_19909,N_14894,N_10781);
and U19910 (N_19910,N_12801,N_13421);
and U19911 (N_19911,N_12486,N_14301);
nand U19912 (N_19912,N_14479,N_13821);
or U19913 (N_19913,N_12722,N_12455);
xor U19914 (N_19914,N_10386,N_12381);
or U19915 (N_19915,N_14625,N_10119);
nor U19916 (N_19916,N_13628,N_10399);
xor U19917 (N_19917,N_14785,N_12432);
or U19918 (N_19918,N_13103,N_14523);
nand U19919 (N_19919,N_13617,N_11226);
nor U19920 (N_19920,N_14567,N_13561);
nand U19921 (N_19921,N_10871,N_14606);
and U19922 (N_19922,N_11926,N_10640);
xnor U19923 (N_19923,N_11837,N_11358);
xor U19924 (N_19924,N_12400,N_10420);
xor U19925 (N_19925,N_12235,N_14234);
and U19926 (N_19926,N_12222,N_13455);
or U19927 (N_19927,N_11395,N_10388);
and U19928 (N_19928,N_12656,N_11237);
nor U19929 (N_19929,N_13447,N_12362);
nor U19930 (N_19930,N_11235,N_11537);
and U19931 (N_19931,N_11454,N_12101);
nand U19932 (N_19932,N_12941,N_12283);
or U19933 (N_19933,N_13011,N_11224);
nor U19934 (N_19934,N_13347,N_11723);
xor U19935 (N_19935,N_13728,N_14387);
nand U19936 (N_19936,N_12599,N_10840);
or U19937 (N_19937,N_12225,N_11023);
nor U19938 (N_19938,N_10184,N_10722);
or U19939 (N_19939,N_10801,N_13006);
xnor U19940 (N_19940,N_12153,N_11093);
nor U19941 (N_19941,N_13121,N_14295);
nand U19942 (N_19942,N_12278,N_12154);
xor U19943 (N_19943,N_10750,N_14512);
nand U19944 (N_19944,N_12902,N_12814);
or U19945 (N_19945,N_11124,N_14715);
xnor U19946 (N_19946,N_10118,N_13085);
xnor U19947 (N_19947,N_14616,N_11520);
nor U19948 (N_19948,N_10970,N_11762);
and U19949 (N_19949,N_10181,N_10903);
or U19950 (N_19950,N_12899,N_10307);
and U19951 (N_19951,N_11095,N_12728);
nor U19952 (N_19952,N_13602,N_11865);
and U19953 (N_19953,N_14266,N_10793);
or U19954 (N_19954,N_12135,N_10946);
and U19955 (N_19955,N_11193,N_14321);
nor U19956 (N_19956,N_13483,N_13610);
nand U19957 (N_19957,N_10934,N_10719);
nand U19958 (N_19958,N_13605,N_13227);
or U19959 (N_19959,N_14734,N_14919);
or U19960 (N_19960,N_10176,N_14375);
and U19961 (N_19961,N_14984,N_14135);
nand U19962 (N_19962,N_11105,N_11769);
xnor U19963 (N_19963,N_12466,N_11013);
nand U19964 (N_19964,N_14578,N_11159);
nand U19965 (N_19965,N_14189,N_14991);
and U19966 (N_19966,N_10568,N_14063);
nor U19967 (N_19967,N_12096,N_11093);
nand U19968 (N_19968,N_14885,N_12917);
and U19969 (N_19969,N_12604,N_12712);
and U19970 (N_19970,N_11211,N_14650);
nand U19971 (N_19971,N_13972,N_11063);
xnor U19972 (N_19972,N_10575,N_10106);
and U19973 (N_19973,N_10340,N_12419);
nor U19974 (N_19974,N_13883,N_13391);
nor U19975 (N_19975,N_10354,N_14754);
xnor U19976 (N_19976,N_10082,N_11497);
and U19977 (N_19977,N_13289,N_10025);
nor U19978 (N_19978,N_13767,N_14625);
or U19979 (N_19979,N_14666,N_13144);
nand U19980 (N_19980,N_12015,N_14090);
nor U19981 (N_19981,N_12996,N_12027);
and U19982 (N_19982,N_12841,N_13830);
nor U19983 (N_19983,N_11943,N_12481);
nand U19984 (N_19984,N_14144,N_13245);
or U19985 (N_19985,N_11139,N_14157);
and U19986 (N_19986,N_10166,N_14308);
xor U19987 (N_19987,N_11655,N_11720);
or U19988 (N_19988,N_12472,N_10639);
xnor U19989 (N_19989,N_14182,N_14800);
or U19990 (N_19990,N_10001,N_11827);
or U19991 (N_19991,N_13322,N_11706);
and U19992 (N_19992,N_14065,N_13400);
nand U19993 (N_19993,N_10653,N_11086);
and U19994 (N_19994,N_10163,N_14825);
nor U19995 (N_19995,N_14845,N_10113);
nand U19996 (N_19996,N_13206,N_11244);
xnor U19997 (N_19997,N_14364,N_12804);
nor U19998 (N_19998,N_12223,N_14050);
and U19999 (N_19999,N_12675,N_13127);
xor U20000 (N_20000,N_18181,N_17331);
or U20001 (N_20001,N_19742,N_17200);
or U20002 (N_20002,N_18113,N_15969);
nand U20003 (N_20003,N_18689,N_15511);
nor U20004 (N_20004,N_15922,N_17733);
or U20005 (N_20005,N_16703,N_19895);
nor U20006 (N_20006,N_18497,N_19053);
nand U20007 (N_20007,N_15319,N_18818);
nor U20008 (N_20008,N_15484,N_18754);
and U20009 (N_20009,N_17679,N_15241);
and U20010 (N_20010,N_18981,N_15268);
or U20011 (N_20011,N_18567,N_16636);
or U20012 (N_20012,N_18732,N_18734);
xor U20013 (N_20013,N_15286,N_19884);
and U20014 (N_20014,N_19986,N_19100);
and U20015 (N_20015,N_18819,N_17325);
and U20016 (N_20016,N_17667,N_19382);
xnor U20017 (N_20017,N_18120,N_18790);
nor U20018 (N_20018,N_18810,N_19186);
and U20019 (N_20019,N_16765,N_15690);
xnor U20020 (N_20020,N_19590,N_17997);
and U20021 (N_20021,N_15534,N_19518);
xor U20022 (N_20022,N_18404,N_15614);
and U20023 (N_20023,N_19888,N_16237);
or U20024 (N_20024,N_16799,N_16878);
or U20025 (N_20025,N_15877,N_15738);
xnor U20026 (N_20026,N_16708,N_15388);
and U20027 (N_20027,N_17498,N_15299);
nand U20028 (N_20028,N_17504,N_19304);
or U20029 (N_20029,N_16472,N_19224);
xnor U20030 (N_20030,N_18477,N_16341);
xor U20031 (N_20031,N_16055,N_16084);
xor U20032 (N_20032,N_18329,N_18163);
or U20033 (N_20033,N_17598,N_18806);
and U20034 (N_20034,N_17623,N_16390);
xnor U20035 (N_20035,N_18054,N_17905);
xnor U20036 (N_20036,N_18487,N_19584);
nand U20037 (N_20037,N_19420,N_18066);
nor U20038 (N_20038,N_18999,N_18867);
and U20039 (N_20039,N_16033,N_17246);
or U20040 (N_20040,N_19270,N_15081);
and U20041 (N_20041,N_16506,N_16825);
or U20042 (N_20042,N_19551,N_19052);
or U20043 (N_20043,N_15675,N_18218);
nand U20044 (N_20044,N_18983,N_15125);
or U20045 (N_20045,N_16467,N_18808);
xor U20046 (N_20046,N_18648,N_15636);
and U20047 (N_20047,N_15341,N_19804);
and U20048 (N_20048,N_17659,N_17151);
or U20049 (N_20049,N_16406,N_18401);
nand U20050 (N_20050,N_16279,N_19196);
nand U20051 (N_20051,N_18081,N_17430);
xnor U20052 (N_20052,N_15361,N_16042);
and U20053 (N_20053,N_17277,N_19525);
xor U20054 (N_20054,N_18047,N_17383);
nand U20055 (N_20055,N_18598,N_18811);
nand U20056 (N_20056,N_19801,N_15314);
nor U20057 (N_20057,N_16586,N_17730);
or U20058 (N_20058,N_17778,N_17683);
nand U20059 (N_20059,N_16359,N_16764);
nand U20060 (N_20060,N_15265,N_15973);
and U20061 (N_20061,N_16508,N_19930);
or U20062 (N_20062,N_17066,N_18311);
or U20063 (N_20063,N_19635,N_15474);
and U20064 (N_20064,N_17154,N_19935);
and U20065 (N_20065,N_17042,N_19378);
and U20066 (N_20066,N_17368,N_15448);
or U20067 (N_20067,N_15993,N_18505);
nand U20068 (N_20068,N_16327,N_15896);
xor U20069 (N_20069,N_19540,N_18893);
or U20070 (N_20070,N_17356,N_15050);
and U20071 (N_20071,N_17382,N_15137);
xor U20072 (N_20072,N_18501,N_18566);
xnor U20073 (N_20073,N_15572,N_17283);
nand U20074 (N_20074,N_17907,N_19033);
xor U20075 (N_20075,N_16271,N_18882);
xor U20076 (N_20076,N_17089,N_15186);
and U20077 (N_20077,N_18672,N_19848);
and U20078 (N_20078,N_18801,N_15423);
and U20079 (N_20079,N_19812,N_16668);
or U20080 (N_20080,N_17652,N_19618);
and U20081 (N_20081,N_19690,N_19566);
or U20082 (N_20082,N_18117,N_15902);
nor U20083 (N_20083,N_17039,N_17747);
nor U20084 (N_20084,N_18438,N_19293);
xor U20085 (N_20085,N_18305,N_16274);
and U20086 (N_20086,N_16844,N_15348);
or U20087 (N_20087,N_16035,N_15152);
xnor U20088 (N_20088,N_15952,N_15622);
nand U20089 (N_20089,N_18112,N_15356);
nand U20090 (N_20090,N_17065,N_15401);
and U20091 (N_20091,N_18560,N_19898);
and U20092 (N_20092,N_18408,N_17304);
xor U20093 (N_20093,N_18315,N_16137);
xor U20094 (N_20094,N_17397,N_18718);
xnor U20095 (N_20095,N_16995,N_16788);
nor U20096 (N_20096,N_16565,N_18165);
or U20097 (N_20097,N_17645,N_17990);
nand U20098 (N_20098,N_18359,N_19177);
nand U20099 (N_20099,N_15948,N_17661);
nor U20100 (N_20100,N_15544,N_16038);
or U20101 (N_20101,N_16691,N_18619);
nand U20102 (N_20102,N_19836,N_15099);
or U20103 (N_20103,N_19751,N_19573);
and U20104 (N_20104,N_15478,N_16850);
or U20105 (N_20105,N_19694,N_18606);
nand U20106 (N_20106,N_18929,N_17192);
nor U20107 (N_20107,N_19767,N_18240);
nand U20108 (N_20108,N_18472,N_16929);
nor U20109 (N_20109,N_17298,N_19046);
or U20110 (N_20110,N_19607,N_15640);
nand U20111 (N_20111,N_16308,N_19017);
nor U20112 (N_20112,N_17409,N_16334);
nor U20113 (N_20113,N_17163,N_15878);
nor U20114 (N_20114,N_17193,N_15900);
xnor U20115 (N_20115,N_16845,N_17428);
or U20116 (N_20116,N_19120,N_16031);
or U20117 (N_20117,N_18450,N_19636);
or U20118 (N_20118,N_15890,N_17771);
nand U20119 (N_20119,N_19016,N_17293);
nor U20120 (N_20120,N_18904,N_16437);
or U20121 (N_20121,N_19204,N_17396);
xnor U20122 (N_20122,N_15101,N_18595);
xnor U20123 (N_20123,N_17272,N_16438);
or U20124 (N_20124,N_15626,N_16083);
nand U20125 (N_20125,N_16671,N_16603);
and U20126 (N_20126,N_16613,N_15217);
nand U20127 (N_20127,N_19855,N_19743);
xor U20128 (N_20128,N_18225,N_19413);
or U20129 (N_20129,N_17617,N_18600);
and U20130 (N_20130,N_16588,N_17278);
and U20131 (N_20131,N_18607,N_16921);
xnor U20132 (N_20132,N_15812,N_16178);
and U20133 (N_20133,N_16740,N_18015);
xnor U20134 (N_20134,N_17714,N_18280);
nand U20135 (N_20135,N_18362,N_16258);
xor U20136 (N_20136,N_16087,N_15403);
nor U20137 (N_20137,N_15523,N_15098);
or U20138 (N_20138,N_19035,N_15836);
nor U20139 (N_20139,N_17991,N_18773);
nor U20140 (N_20140,N_16628,N_16937);
nand U20141 (N_20141,N_19259,N_18095);
and U20142 (N_20142,N_16062,N_17943);
nand U20143 (N_20143,N_15672,N_17286);
or U20144 (N_20144,N_18223,N_17202);
or U20145 (N_20145,N_15264,N_17461);
nor U20146 (N_20146,N_17091,N_18104);
and U20147 (N_20147,N_16655,N_17988);
nor U20148 (N_20148,N_16804,N_18296);
nand U20149 (N_20149,N_19104,N_17827);
or U20150 (N_20150,N_16635,N_17388);
xnor U20151 (N_20151,N_16514,N_17243);
and U20152 (N_20152,N_19392,N_15479);
and U20153 (N_20153,N_16839,N_15866);
nor U20154 (N_20154,N_17213,N_16101);
nand U20155 (N_20155,N_19334,N_19332);
or U20156 (N_20156,N_18623,N_15542);
and U20157 (N_20157,N_15277,N_15525);
or U20158 (N_20158,N_15038,N_17096);
nor U20159 (N_20159,N_16906,N_16871);
and U20160 (N_20160,N_17033,N_18881);
nor U20161 (N_20161,N_15129,N_16287);
nor U20162 (N_20162,N_17152,N_16591);
xnor U20163 (N_20163,N_17586,N_15008);
or U20164 (N_20164,N_19122,N_15999);
xor U20165 (N_20165,N_16908,N_17385);
xnor U20166 (N_20166,N_16700,N_15467);
or U20167 (N_20167,N_17289,N_16497);
and U20168 (N_20168,N_15698,N_19933);
and U20169 (N_20169,N_17517,N_17234);
nor U20170 (N_20170,N_16365,N_19832);
nand U20171 (N_20171,N_19005,N_15921);
and U20172 (N_20172,N_18554,N_17155);
and U20173 (N_20173,N_16060,N_16932);
nor U20174 (N_20174,N_19133,N_17266);
nand U20175 (N_20175,N_15420,N_19401);
and U20176 (N_20176,N_16429,N_18274);
nor U20177 (N_20177,N_16539,N_18268);
nand U20178 (N_20178,N_19647,N_15965);
and U20179 (N_20179,N_18093,N_15691);
xnor U20180 (N_20180,N_18306,N_18992);
nand U20181 (N_20181,N_17421,N_16134);
nor U20182 (N_20182,N_18677,N_15055);
xnor U20183 (N_20183,N_15564,N_18187);
nor U20184 (N_20184,N_16532,N_16120);
and U20185 (N_20185,N_19858,N_19187);
nor U20186 (N_20186,N_15901,N_19572);
xor U20187 (N_20187,N_17785,N_18536);
xnor U20188 (N_20188,N_15188,N_17693);
or U20189 (N_20189,N_18580,N_15653);
xnor U20190 (N_20190,N_18633,N_19265);
and U20191 (N_20191,N_19312,N_18034);
or U20192 (N_20192,N_17717,N_19949);
xnor U20193 (N_20193,N_16216,N_19143);
nand U20194 (N_20194,N_17427,N_18544);
or U20195 (N_20195,N_18690,N_15214);
nor U20196 (N_20196,N_16209,N_17027);
or U20197 (N_20197,N_18979,N_18746);
and U20198 (N_20198,N_17539,N_15350);
or U20199 (N_20199,N_19211,N_19622);
or U20200 (N_20200,N_15810,N_19765);
or U20201 (N_20201,N_19687,N_16527);
nor U20202 (N_20202,N_16175,N_18177);
nand U20203 (N_20203,N_15285,N_19605);
xnor U20204 (N_20204,N_19337,N_18457);
and U20205 (N_20205,N_16115,N_17405);
or U20206 (N_20206,N_18609,N_16448);
nand U20207 (N_20207,N_18955,N_19171);
or U20208 (N_20208,N_19168,N_17114);
nor U20209 (N_20209,N_17808,N_19314);
or U20210 (N_20210,N_19106,N_18744);
nor U20211 (N_20211,N_15592,N_17115);
xnor U20212 (N_20212,N_19075,N_19020);
nor U20213 (N_20213,N_17822,N_17431);
xor U20214 (N_20214,N_19873,N_17166);
or U20215 (N_20215,N_19841,N_19464);
or U20216 (N_20216,N_18070,N_15760);
nor U20217 (N_20217,N_17005,N_18786);
nor U20218 (N_20218,N_19633,N_18944);
and U20219 (N_20219,N_15439,N_19927);
nand U20220 (N_20220,N_19952,N_17444);
xnor U20221 (N_20221,N_15167,N_17767);
or U20222 (N_20222,N_16148,N_15642);
nand U20223 (N_20223,N_16164,N_16716);
and U20224 (N_20224,N_17466,N_15708);
or U20225 (N_20225,N_17178,N_16447);
and U20226 (N_20226,N_16598,N_16597);
or U20227 (N_20227,N_16678,N_18183);
and U20228 (N_20228,N_17252,N_16785);
nand U20229 (N_20229,N_18594,N_16957);
and U20230 (N_20230,N_18069,N_19004);
or U20231 (N_20231,N_16142,N_15747);
nand U20232 (N_20232,N_19655,N_17496);
and U20233 (N_20233,N_15774,N_17490);
nor U20234 (N_20234,N_16894,N_15359);
nor U20235 (N_20235,N_19821,N_17462);
xnor U20236 (N_20236,N_16939,N_16984);
nand U20237 (N_20237,N_17825,N_15272);
nor U20238 (N_20238,N_17270,N_18193);
and U20239 (N_20239,N_16174,N_16430);
nor U20240 (N_20240,N_16284,N_18476);
or U20241 (N_20241,N_16583,N_16498);
xnor U20242 (N_20242,N_17754,N_15213);
or U20243 (N_20243,N_17608,N_18937);
xor U20244 (N_20244,N_18182,N_16391);
and U20245 (N_20245,N_19970,N_17622);
or U20246 (N_20246,N_16354,N_15425);
nand U20247 (N_20247,N_16873,N_15279);
or U20248 (N_20248,N_17505,N_15907);
nand U20249 (N_20249,N_17875,N_19712);
or U20250 (N_20250,N_15576,N_16130);
nand U20251 (N_20251,N_18565,N_17326);
nor U20252 (N_20252,N_15502,N_15597);
xor U20253 (N_20253,N_18407,N_19134);
or U20254 (N_20254,N_16749,N_19966);
nand U20255 (N_20255,N_18587,N_15624);
nand U20256 (N_20256,N_19676,N_19044);
nor U20257 (N_20257,N_16195,N_16525);
or U20258 (N_20258,N_18755,N_19803);
and U20259 (N_20259,N_19511,N_18221);
nand U20260 (N_20260,N_15360,N_16074);
or U20261 (N_20261,N_19583,N_17620);
and U20262 (N_20262,N_18976,N_15077);
or U20263 (N_20263,N_19084,N_17782);
nand U20264 (N_20264,N_16676,N_18716);
nor U20265 (N_20265,N_16990,N_18701);
nand U20266 (N_20266,N_15234,N_17751);
and U20267 (N_20267,N_15192,N_17551);
or U20268 (N_20268,N_18332,N_19626);
and U20269 (N_20269,N_17101,N_15225);
nor U20270 (N_20270,N_16857,N_17432);
nand U20271 (N_20271,N_15758,N_18875);
nand U20272 (N_20272,N_18303,N_17222);
and U20273 (N_20273,N_15147,N_16732);
or U20274 (N_20274,N_19995,N_19624);
nand U20275 (N_20275,N_16612,N_19737);
or U20276 (N_20276,N_15826,N_18276);
nor U20277 (N_20277,N_16260,N_18398);
or U20278 (N_20278,N_17439,N_17524);
nand U20279 (N_20279,N_17402,N_15091);
xnor U20280 (N_20280,N_18051,N_16286);
xor U20281 (N_20281,N_18661,N_16088);
nand U20282 (N_20282,N_15911,N_17209);
xor U20283 (N_20283,N_15159,N_15575);
nand U20284 (N_20284,N_19740,N_16604);
xnor U20285 (N_20285,N_17641,N_18764);
and U20286 (N_20286,N_18076,N_17833);
nor U20287 (N_20287,N_15524,N_15571);
or U20288 (N_20288,N_16587,N_18556);
or U20289 (N_20289,N_17352,N_17725);
nand U20290 (N_20290,N_19552,N_15431);
or U20291 (N_20291,N_18074,N_18586);
and U20292 (N_20292,N_17902,N_17982);
or U20293 (N_20293,N_19271,N_16493);
nor U20294 (N_20294,N_19711,N_18502);
nor U20295 (N_20295,N_19015,N_17854);
or U20296 (N_20296,N_19846,N_16288);
or U20297 (N_20297,N_17317,N_19919);
xor U20298 (N_20298,N_18319,N_17791);
nand U20299 (N_20299,N_17210,N_17157);
nand U20300 (N_20300,N_18060,N_17216);
xor U20301 (N_20301,N_16832,N_15685);
and U20302 (N_20302,N_15022,N_17310);
xor U20303 (N_20303,N_16553,N_15813);
xor U20304 (N_20304,N_19307,N_15715);
nand U20305 (N_20305,N_15223,N_17533);
xnor U20306 (N_20306,N_16189,N_15288);
and U20307 (N_20307,N_18155,N_18265);
nand U20308 (N_20308,N_19350,N_17819);
nor U20309 (N_20309,N_16199,N_16435);
and U20310 (N_20310,N_15351,N_15606);
or U20311 (N_20311,N_18876,N_19650);
or U20312 (N_20312,N_15851,N_19277);
xnor U20313 (N_20313,N_18304,N_15113);
xor U20314 (N_20314,N_19643,N_18281);
xor U20315 (N_20315,N_19296,N_16868);
and U20316 (N_20316,N_17554,N_15260);
or U20317 (N_20317,N_15405,N_16206);
xor U20318 (N_20318,N_16469,N_16487);
and U20319 (N_20319,N_18235,N_16580);
and U20320 (N_20320,N_18706,N_17106);
and U20321 (N_20321,N_18919,N_19748);
nand U20322 (N_20322,N_17477,N_15271);
or U20323 (N_20323,N_15396,N_15857);
or U20324 (N_20324,N_15028,N_19623);
and U20325 (N_20325,N_18059,N_15251);
xor U20326 (N_20326,N_18243,N_15389);
xnor U20327 (N_20327,N_15230,N_16556);
nand U20328 (N_20328,N_15003,N_15079);
or U20329 (N_20329,N_15639,N_18026);
and U20330 (N_20330,N_16602,N_16901);
nand U20331 (N_20331,N_18640,N_19485);
or U20332 (N_20332,N_19375,N_15834);
nor U20333 (N_20333,N_18599,N_17781);
or U20334 (N_20334,N_19602,N_15300);
nor U20335 (N_20335,N_18577,N_15700);
or U20336 (N_20336,N_17942,N_15753);
nand U20337 (N_20337,N_16898,N_19907);
xor U20338 (N_20338,N_18572,N_17527);
and U20339 (N_20339,N_15864,N_18325);
xor U20340 (N_20340,N_19967,N_19254);
xor U20341 (N_20341,N_18982,N_19893);
or U20342 (N_20342,N_17214,N_18503);
xnor U20343 (N_20343,N_15619,N_17132);
or U20344 (N_20344,N_19613,N_19400);
nor U20345 (N_20345,N_18793,N_16959);
nor U20346 (N_20346,N_18016,N_18114);
nor U20347 (N_20347,N_16006,N_18234);
nor U20348 (N_20348,N_18172,N_17834);
or U20349 (N_20349,N_19632,N_19428);
nand U20350 (N_20350,N_18190,N_16298);
or U20351 (N_20351,N_15682,N_16106);
and U20352 (N_20352,N_15441,N_15017);
xor U20353 (N_20353,N_19792,N_18727);
xor U20354 (N_20354,N_17333,N_18159);
and U20355 (N_20355,N_17004,N_16723);
or U20356 (N_20356,N_19531,N_17451);
and U20357 (N_20357,N_15990,N_15338);
and U20358 (N_20358,N_17790,N_19147);
and U20359 (N_20359,N_18092,N_19688);
or U20360 (N_20360,N_15703,N_18232);
nand U20361 (N_20361,N_15298,N_16413);
xnor U20362 (N_20362,N_18551,N_19809);
or U20363 (N_20363,N_17876,N_17412);
or U20364 (N_20364,N_17122,N_18423);
or U20365 (N_20365,N_17153,N_17689);
or U20366 (N_20366,N_18984,N_18446);
nor U20367 (N_20367,N_17606,N_16236);
nor U20368 (N_20368,N_19191,N_17219);
and U20369 (N_20369,N_17268,N_18042);
nor U20370 (N_20370,N_17478,N_16849);
xor U20371 (N_20371,N_19331,N_15026);
or U20372 (N_20372,N_17036,N_17002);
nand U20373 (N_20373,N_17958,N_15493);
or U20374 (N_20374,N_17457,N_18330);
nand U20375 (N_20375,N_15858,N_15992);
nor U20376 (N_20376,N_19348,N_18056);
and U20377 (N_20377,N_16177,N_19074);
nor U20378 (N_20378,N_18435,N_16803);
and U20379 (N_20379,N_15780,N_15587);
and U20380 (N_20380,N_16985,N_16645);
or U20381 (N_20381,N_19105,N_18058);
nand U20382 (N_20382,N_19166,N_17257);
nand U20383 (N_20383,N_15889,N_17740);
or U20384 (N_20384,N_18430,N_16141);
or U20385 (N_20385,N_15424,N_18781);
nor U20386 (N_20386,N_19825,N_19423);
xor U20387 (N_20387,N_19497,N_15659);
xnor U20388 (N_20388,N_17897,N_17910);
xor U20389 (N_20389,N_15053,N_15793);
xnor U20390 (N_20390,N_16779,N_15428);
or U20391 (N_20391,N_17715,N_17887);
nand U20392 (N_20392,N_19764,N_18237);
or U20393 (N_20393,N_17404,N_17313);
nand U20394 (N_20394,N_16960,N_15920);
and U20395 (N_20395,N_15604,N_19288);
nor U20396 (N_20396,N_17150,N_19154);
or U20397 (N_20397,N_16481,N_18314);
nand U20398 (N_20398,N_17137,N_18552);
nor U20399 (N_20399,N_15057,N_16372);
or U20400 (N_20400,N_15398,N_15983);
xor U20401 (N_20401,N_16766,N_18602);
or U20402 (N_20402,N_16388,N_16250);
or U20403 (N_20403,N_15074,N_17548);
or U20404 (N_20404,N_17953,N_16996);
nor U20405 (N_20405,N_17063,N_15732);
or U20406 (N_20406,N_17773,N_16097);
nand U20407 (N_20407,N_16717,N_18662);
nand U20408 (N_20408,N_15844,N_17672);
and U20409 (N_20409,N_19414,N_17564);
and U20410 (N_20410,N_17060,N_17815);
nand U20411 (N_20411,N_19125,N_18679);
or U20412 (N_20412,N_15471,N_18465);
and U20413 (N_20413,N_19273,N_18410);
or U20414 (N_20414,N_19911,N_16348);
xnor U20415 (N_20415,N_15168,N_16865);
or U20416 (N_20416,N_16893,N_15962);
or U20417 (N_20417,N_18127,N_17816);
xor U20418 (N_20418,N_15964,N_17393);
and U20419 (N_20419,N_15245,N_18555);
xnor U20420 (N_20420,N_15945,N_17770);
or U20421 (N_20421,N_15496,N_15221);
nand U20422 (N_20422,N_18949,N_17124);
xor U20423 (N_20423,N_16049,N_15292);
nor U20424 (N_20424,N_15713,N_19089);
or U20425 (N_20425,N_17529,N_18885);
and U20426 (N_20426,N_19374,N_16646);
or U20427 (N_20427,N_19776,N_15465);
or U20428 (N_20428,N_17845,N_17454);
xor U20429 (N_20429,N_18135,N_15568);
and U20430 (N_20430,N_15436,N_18212);
and U20431 (N_20431,N_16854,N_19426);
nand U20432 (N_20432,N_17817,N_17225);
xor U20433 (N_20433,N_18205,N_18705);
xor U20434 (N_20434,N_15248,N_18749);
nand U20435 (N_20435,N_18965,N_17379);
and U20436 (N_20436,N_17281,N_16020);
xor U20437 (N_20437,N_16807,N_16463);
and U20438 (N_20438,N_19308,N_17322);
nor U20439 (N_20439,N_17500,N_19508);
or U20440 (N_20440,N_19714,N_16217);
nor U20441 (N_20441,N_18709,N_17165);
xor U20442 (N_20442,N_18115,N_18197);
nand U20443 (N_20443,N_16963,N_17125);
and U20444 (N_20444,N_17207,N_17668);
nor U20445 (N_20445,N_19468,N_17471);
nor U20446 (N_20446,N_16369,N_16358);
nor U20447 (N_20447,N_15744,N_19671);
or U20448 (N_20448,N_18767,N_17468);
xnor U20449 (N_20449,N_18474,N_15114);
nor U20450 (N_20450,N_15048,N_18559);
xnor U20451 (N_20451,N_16529,N_19424);
xnor U20452 (N_20452,N_17479,N_15294);
nand U20453 (N_20453,N_16362,N_19183);
nand U20454 (N_20454,N_16666,N_17301);
nor U20455 (N_20455,N_18722,N_17175);
nor U20456 (N_20456,N_18393,N_18852);
or U20457 (N_20457,N_16086,N_16623);
nor U20458 (N_20458,N_18129,N_16210);
xnor U20459 (N_20459,N_18011,N_17727);
and U20460 (N_20460,N_19363,N_18085);
nor U20461 (N_20461,N_15237,N_15840);
or U20462 (N_20462,N_17158,N_19815);
and U20463 (N_20463,N_17968,N_15058);
and U20464 (N_20464,N_17480,N_17093);
and U20465 (N_20465,N_18336,N_18653);
nor U20466 (N_20466,N_15335,N_16801);
xor U20467 (N_20467,N_16465,N_18691);
nand U20468 (N_20468,N_18291,N_17118);
nand U20469 (N_20469,N_15397,N_15566);
nor U20470 (N_20470,N_16971,N_18029);
nand U20471 (N_20471,N_15862,N_15795);
or U20472 (N_20472,N_19360,N_17811);
or U20473 (N_20473,N_15722,N_17945);
or U20474 (N_20474,N_19438,N_19543);
and U20475 (N_20475,N_19582,N_17327);
and U20476 (N_20476,N_18249,N_15417);
and U20477 (N_20477,N_18721,N_16466);
nand U20478 (N_20478,N_18012,N_15580);
and U20479 (N_20479,N_17674,N_16926);
and U20480 (N_20480,N_17535,N_15290);
or U20481 (N_20481,N_19354,N_16283);
or U20482 (N_20482,N_18805,N_16314);
nand U20483 (N_20483,N_16615,N_15908);
and U20484 (N_20484,N_15897,N_17198);
and U20485 (N_20485,N_17923,N_16294);
or U20486 (N_20486,N_15203,N_18561);
and U20487 (N_20487,N_19189,N_15766);
nand U20488 (N_20488,N_17308,N_16238);
nand U20489 (N_20489,N_16114,N_15071);
or U20490 (N_20490,N_19478,N_18510);
or U20491 (N_20491,N_15714,N_18972);
nand U20492 (N_20492,N_17795,N_16907);
nor U20493 (N_20493,N_17611,N_18657);
or U20494 (N_20494,N_18967,N_15193);
nor U20495 (N_20495,N_15106,N_16977);
xor U20496 (N_20496,N_19981,N_15839);
nor U20497 (N_20497,N_16685,N_19081);
and U20498 (N_20498,N_19739,N_19500);
and U20499 (N_20499,N_18943,N_15224);
nor U20500 (N_20500,N_19404,N_18688);
xor U20501 (N_20501,N_17675,N_18024);
or U20502 (N_20502,N_16127,N_18403);
xnor U20503 (N_20503,N_19221,N_18277);
or U20504 (N_20504,N_19145,N_19940);
or U20505 (N_20505,N_18930,N_16639);
nor U20506 (N_20506,N_18517,N_18581);
nand U20507 (N_20507,N_15958,N_16518);
xor U20508 (N_20508,N_15030,N_16292);
xor U20509 (N_20509,N_19985,N_19498);
and U20510 (N_20510,N_18142,N_15131);
nor U20511 (N_20511,N_19736,N_15546);
xor U20512 (N_20512,N_18643,N_19625);
nor U20513 (N_20513,N_16045,N_15573);
nor U20514 (N_20514,N_16139,N_15173);
nor U20515 (N_20515,N_19609,N_17129);
nor U20516 (N_20516,N_16126,N_18484);
nor U20517 (N_20517,N_16777,N_15943);
nor U20518 (N_20518,N_18666,N_19717);
xnor U20519 (N_20519,N_18951,N_15240);
nand U20520 (N_20520,N_17750,N_19396);
and U20521 (N_20521,N_17419,N_15696);
or U20522 (N_20522,N_19102,N_17460);
and U20523 (N_20523,N_16987,N_15387);
nand U20524 (N_20524,N_19529,N_19509);
nand U20525 (N_20525,N_15815,N_17189);
and U20526 (N_20526,N_17447,N_16669);
nand U20527 (N_20527,N_19849,N_15392);
nor U20528 (N_20528,N_18729,N_19116);
xor U20529 (N_20529,N_16817,N_18974);
or U20530 (N_20530,N_19790,N_16630);
nand U20531 (N_20531,N_15354,N_15799);
xnor U20532 (N_20532,N_19250,N_19032);
and U20533 (N_20533,N_16379,N_19333);
or U20534 (N_20534,N_15201,N_15047);
xnor U20535 (N_20535,N_17957,N_18608);
xnor U20536 (N_20536,N_17938,N_18596);
nor U20537 (N_20537,N_18851,N_18761);
xnor U20538 (N_20538,N_19645,N_18860);
nor U20539 (N_20539,N_16160,N_19246);
or U20540 (N_20540,N_16701,N_19048);
nor U20541 (N_20541,N_17149,N_18367);
xor U20542 (N_20542,N_19963,N_17482);
nand U20543 (N_20543,N_15104,N_18337);
xor U20544 (N_20544,N_17259,N_18444);
and U20545 (N_20545,N_19190,N_19514);
xor U20546 (N_20546,N_17871,N_17459);
nor U20547 (N_20547,N_18158,N_17635);
nand U20548 (N_20548,N_18927,N_17831);
nor U20549 (N_20549,N_15516,N_16861);
nand U20550 (N_20550,N_16780,N_16791);
and U20551 (N_20551,N_19559,N_19408);
nor U20552 (N_20552,N_18879,N_19941);
xor U20553 (N_20553,N_17497,N_18039);
nor U20554 (N_20554,N_18239,N_15731);
and U20555 (N_20555,N_18342,N_17848);
nor U20556 (N_20556,N_18802,N_19701);
xnor U20557 (N_20557,N_16755,N_18286);
or U20558 (N_20558,N_16899,N_17956);
nor U20559 (N_20559,N_15233,N_18655);
or U20560 (N_20560,N_15164,N_18571);
xnor U20561 (N_20561,N_18191,N_17377);
or U20562 (N_20562,N_15333,N_15069);
or U20563 (N_20563,N_19578,N_18381);
xnor U20564 (N_20564,N_16823,N_18222);
nor U20565 (N_20565,N_15560,N_19341);
and U20566 (N_20566,N_16856,N_18160);
nor U20567 (N_20567,N_19193,N_15051);
nand U20568 (N_20568,N_18124,N_16896);
nand U20569 (N_20569,N_19069,N_19245);
or U20570 (N_20570,N_16419,N_19778);
nand U20571 (N_20571,N_19150,N_15199);
and U20572 (N_20572,N_18442,N_18796);
xor U20573 (N_20573,N_15100,N_15043);
or U20574 (N_20574,N_16113,N_17557);
nor U20575 (N_20575,N_19544,N_19611);
nor U20576 (N_20576,N_18647,N_18415);
and U20577 (N_20577,N_16482,N_19109);
or U20578 (N_20578,N_16040,N_16345);
or U20579 (N_20579,N_18002,N_16533);
nor U20580 (N_20580,N_19167,N_16952);
nand U20581 (N_20581,N_18918,N_16917);
or U20582 (N_20582,N_16515,N_19780);
and U20583 (N_20583,N_17360,N_17918);
nand U20584 (N_20584,N_15763,N_17037);
and U20585 (N_20585,N_18171,N_18251);
xnor U20586 (N_20586,N_16054,N_17003);
and U20587 (N_20587,N_19845,N_15469);
or U20588 (N_20588,N_16682,N_19987);
nor U20589 (N_20589,N_17264,N_15324);
and U20590 (N_20590,N_19484,N_18912);
nand U20591 (N_20591,N_15197,N_16150);
and U20592 (N_20592,N_16574,N_19515);
xnor U20593 (N_20593,N_16244,N_16434);
or U20594 (N_20594,N_17768,N_19482);
or U20595 (N_20595,N_16902,N_15504);
nand U20596 (N_20596,N_18125,N_17488);
nand U20597 (N_20597,N_17067,N_17450);
and U20598 (N_20598,N_16999,N_17701);
or U20599 (N_20599,N_18140,N_15916);
xnor U20600 (N_20600,N_15784,N_19228);
and U20601 (N_20601,N_19505,N_15347);
nand U20602 (N_20602,N_18216,N_17842);
nor U20603 (N_20603,N_15779,N_16382);
and U20604 (N_20604,N_16798,N_18473);
nor U20605 (N_20605,N_19915,N_15608);
and U20606 (N_20606,N_16725,N_19659);
nand U20607 (N_20607,N_15453,N_16442);
nand U20608 (N_20608,N_18756,N_15015);
xnor U20609 (N_20609,N_15372,N_19151);
nor U20610 (N_20610,N_18695,N_18150);
or U20611 (N_20611,N_15538,N_15154);
xor U20612 (N_20612,N_16226,N_16910);
nand U20613 (N_20613,N_15412,N_15994);
or U20614 (N_20614,N_18211,N_15667);
or U20615 (N_20615,N_18293,N_19297);
nand U20616 (N_20616,N_17362,N_17328);
nand U20617 (N_20617,N_16642,N_17273);
and U20618 (N_20618,N_19603,N_16767);
nor U20619 (N_20619,N_15312,N_15282);
xnor U20620 (N_20620,N_15177,N_18646);
nand U20621 (N_20621,N_15988,N_17699);
nand U20622 (N_20622,N_15327,N_16312);
and U20623 (N_20623,N_17068,N_15689);
xor U20624 (N_20624,N_17824,N_17977);
and U20625 (N_20625,N_18084,N_16507);
nor U20626 (N_20626,N_15332,N_17525);
nand U20627 (N_20627,N_17182,N_16241);
and U20628 (N_20628,N_16255,N_18372);
xnor U20629 (N_20629,N_17986,N_17226);
nand U20630 (N_20630,N_16027,N_19372);
nor U20631 (N_20631,N_16140,N_17981);
nor U20632 (N_20632,N_19580,N_18317);
nor U20633 (N_20633,N_16546,N_15778);
and U20634 (N_20634,N_15909,N_17334);
xnor U20635 (N_20635,N_18735,N_17676);
nor U20636 (N_20636,N_17545,N_18447);
nand U20637 (N_20637,N_18597,N_16576);
nand U20638 (N_20638,N_18528,N_16278);
nand U20639 (N_20639,N_19258,N_18073);
nand U20640 (N_20640,N_16806,N_19407);
nor U20641 (N_20641,N_15872,N_17306);
and U20642 (N_20642,N_19264,N_18354);
xnor U20643 (N_20643,N_16007,N_19057);
nor U20644 (N_20644,N_15035,N_19144);
nor U20645 (N_20645,N_16230,N_17810);
nor U20646 (N_20646,N_18383,N_16843);
nand U20647 (N_20647,N_16151,N_17761);
nor U20648 (N_20648,N_16268,N_15464);
nor U20649 (N_20649,N_15832,N_18116);
or U20650 (N_20650,N_19194,N_15521);
xor U20651 (N_20651,N_15741,N_17392);
and U20652 (N_20652,N_17995,N_18699);
or U20653 (N_20653,N_17798,N_18063);
nand U20654 (N_20654,N_17448,N_15925);
or U20655 (N_20655,N_18040,N_15369);
nor U20656 (N_20656,N_17851,N_15005);
or U20657 (N_20657,N_15442,N_17410);
nand U20658 (N_20658,N_16225,N_17148);
nand U20659 (N_20659,N_15687,N_16531);
and U20660 (N_20660,N_15884,N_19604);
and U20661 (N_20661,N_16895,N_15623);
xor U20662 (N_20662,N_19799,N_17728);
nand U20663 (N_20663,N_18228,N_19315);
or U20664 (N_20664,N_16024,N_19541);
nand U20665 (N_20665,N_18960,N_16485);
nand U20666 (N_20666,N_16479,N_18564);
nor U20667 (N_20667,N_16138,N_17823);
nand U20668 (N_20668,N_19090,N_15761);
and U20669 (N_20669,N_15583,N_16273);
nor U20670 (N_20670,N_18702,N_17522);
and U20671 (N_20671,N_19899,N_15036);
xor U20672 (N_20672,N_17437,N_19184);
xnor U20673 (N_20673,N_16491,N_19910);
xor U20674 (N_20674,N_15379,N_15646);
nor U20675 (N_20675,N_18605,N_18962);
nor U20676 (N_20676,N_19971,N_17110);
or U20677 (N_20677,N_19630,N_16347);
nand U20678 (N_20678,N_17749,N_18866);
and U20679 (N_20679,N_16110,N_15512);
or U20680 (N_20680,N_15590,N_19345);
nand U20681 (N_20681,N_16403,N_17181);
xor U20682 (N_20682,N_18148,N_19094);
nor U20683 (N_20683,N_17241,N_17349);
nand U20684 (N_20684,N_16395,N_18350);
or U20685 (N_20685,N_15370,N_17176);
and U20686 (N_20686,N_16768,N_16794);
and U20687 (N_20687,N_17010,N_16927);
and U20688 (N_20688,N_16829,N_19008);
nor U20689 (N_20689,N_18080,N_17269);
and U20690 (N_20690,N_18445,N_16909);
or U20691 (N_20691,N_15342,N_18263);
nand U20692 (N_20692,N_19087,N_18352);
xnor U20693 (N_20693,N_16980,N_17543);
xnor U20694 (N_20694,N_16316,N_19527);
and U20695 (N_20695,N_17365,N_19922);
nor U20696 (N_20696,N_16408,N_18247);
and U20697 (N_20697,N_15960,N_16103);
nand U20698 (N_20698,N_16681,N_17828);
or U20699 (N_20699,N_19409,N_19364);
or U20700 (N_20700,N_18738,N_17276);
xnor U20701 (N_20701,N_19066,N_16864);
or U20702 (N_20702,N_19951,N_17994);
xor U20703 (N_20703,N_17926,N_16870);
or U20704 (N_20704,N_16322,N_19195);
nand U20705 (N_20705,N_18297,N_18479);
xor U20706 (N_20706,N_15452,N_15382);
and U20707 (N_20707,N_15674,N_16981);
and U20708 (N_20708,N_18464,N_16925);
nor U20709 (N_20709,N_15016,N_15130);
or U20710 (N_20710,N_16831,N_15120);
xnor U20711 (N_20711,N_17783,N_18774);
and U20712 (N_20712,N_19697,N_19289);
or U20713 (N_20713,N_16228,N_18858);
xnor U20714 (N_20714,N_15284,N_17090);
nor U20715 (N_20715,N_16496,N_16069);
nor U20716 (N_20716,N_16459,N_15616);
xor U20717 (N_20717,N_15283,N_19842);
nor U20718 (N_20718,N_15817,N_18259);
or U20719 (N_20719,N_19906,N_17187);
nand U20720 (N_20720,N_19278,N_19774);
nor U20721 (N_20721,N_16759,N_15818);
nand U20722 (N_20722,N_19904,N_18950);
xnor U20723 (N_20723,N_16090,N_17721);
and U20724 (N_20724,N_15794,N_15419);
xnor U20725 (N_20725,N_19668,N_15171);
xor U20726 (N_20726,N_16008,N_16004);
nor U20727 (N_20727,N_19160,N_15932);
nor U20728 (N_20728,N_15589,N_19076);
and U20729 (N_20729,N_17944,N_18419);
nor U20730 (N_20730,N_16184,N_17078);
xor U20731 (N_20731,N_18521,N_18266);
nor U20732 (N_20732,N_19955,N_15355);
xor U20733 (N_20733,N_17575,N_19488);
or U20734 (N_20734,N_15339,N_17144);
nand U20735 (N_20735,N_18273,N_18534);
and U20736 (N_20736,N_16221,N_18920);
nand U20737 (N_20737,N_16267,N_16559);
or U20738 (N_20738,N_18978,N_19926);
or U20739 (N_20739,N_19431,N_15353);
and U20740 (N_20740,N_16675,N_19136);
or U20741 (N_20741,N_16235,N_15447);
and U20742 (N_20742,N_17436,N_16739);
or U20743 (N_20743,N_15729,N_17562);
and U20744 (N_20744,N_18246,N_15893);
xnor U20745 (N_20745,N_16782,N_19817);
nand U20746 (N_20746,N_17510,N_16842);
xor U20747 (N_20747,N_17640,N_19082);
or U20748 (N_20748,N_19208,N_17571);
nand U20749 (N_20749,N_17336,N_19358);
nand U20750 (N_20750,N_19324,N_16738);
and U20751 (N_20751,N_19567,N_15632);
xnor U20752 (N_20752,N_16727,N_16916);
or U20753 (N_20753,N_18931,N_17932);
xnor U20754 (N_20754,N_19925,N_19859);
or U20755 (N_20755,N_17179,N_15445);
nor U20756 (N_20756,N_15968,N_15457);
or U20757 (N_20757,N_18389,N_17417);
or U20758 (N_20758,N_16205,N_16695);
nand U20759 (N_20759,N_19479,N_17865);
xnor U20760 (N_20760,N_16659,N_15185);
nor U20761 (N_20761,N_17920,N_16824);
nor U20762 (N_20762,N_16724,N_16420);
and U20763 (N_20763,N_18369,N_18686);
nand U20764 (N_20764,N_16077,N_16021);
xor U20765 (N_20765,N_18432,N_17694);
and U20766 (N_20766,N_19735,N_17753);
and U20767 (N_20767,N_17073,N_16185);
xor U20768 (N_20768,N_16841,N_17011);
nor U20769 (N_20769,N_15631,N_19684);
nor U20770 (N_20770,N_17669,N_16263);
and U20771 (N_20771,N_15856,N_16504);
nand U20772 (N_20772,N_18956,N_19554);
and U20773 (N_20773,N_17315,N_19310);
xnor U20774 (N_20774,N_16883,N_17350);
and U20775 (N_20775,N_17057,N_16735);
xor U20776 (N_20776,N_17287,N_17296);
and U20777 (N_20777,N_17970,N_16219);
and U20778 (N_20778,N_16066,N_17655);
or U20779 (N_20779,N_16931,N_19495);
nor U20780 (N_20780,N_18496,N_19418);
nor U20781 (N_20781,N_16774,N_17526);
and U20782 (N_20782,N_15459,N_16125);
xnor U20783 (N_20783,N_16462,N_15023);
nor U20784 (N_20784,N_15450,N_16641);
and U20785 (N_20785,N_16988,N_16962);
nand U20786 (N_20786,N_15141,N_19558);
nor U20787 (N_20787,N_19950,N_15970);
and U20788 (N_20788,N_17514,N_16041);
xnor U20789 (N_20789,N_17980,N_18925);
nand U20790 (N_20790,N_15358,N_15855);
nand U20791 (N_20791,N_19294,N_15311);
xor U20792 (N_20792,N_17523,N_19707);
nor U20793 (N_20793,N_17948,N_19127);
nor U20794 (N_20794,N_19242,N_15561);
xor U20795 (N_20795,N_19954,N_15373);
nand U20796 (N_20796,N_19871,N_15320);
nand U20797 (N_20797,N_19012,N_16704);
nand U20798 (N_20798,N_19990,N_15882);
or U20799 (N_20799,N_19857,N_17614);
and U20800 (N_20800,N_15182,N_18615);
nand U20801 (N_20801,N_19503,N_18388);
xnor U20802 (N_20802,N_18550,N_15937);
nor U20803 (N_20803,N_17185,N_19346);
and U20804 (N_20804,N_15644,N_19338);
and U20805 (N_20805,N_17912,N_17199);
and U20806 (N_20806,N_16193,N_19272);
nor U20807 (N_20807,N_15535,N_17610);
xnor U20808 (N_20808,N_18777,N_18004);
nor U20809 (N_20809,N_17805,N_15977);
or U20810 (N_20810,N_15663,N_17032);
xnor U20811 (N_20811,N_15783,N_17563);
or U20812 (N_20812,N_17565,N_16458);
nor U20813 (N_20813,N_17463,N_15656);
xnor U20814 (N_20814,N_16795,N_17474);
or U20815 (N_20815,N_19979,N_19634);
or U20816 (N_20816,N_16548,N_19397);
or U20817 (N_20817,N_18147,N_15737);
xor U20818 (N_20818,N_17707,N_17638);
nand U20819 (N_20819,N_16421,N_18765);
nand U20820 (N_20820,N_16276,N_15529);
nand U20821 (N_20821,N_17022,N_15328);
and U20822 (N_20822,N_19445,N_19230);
xnor U20823 (N_20823,N_18036,N_18998);
or U20824 (N_20824,N_17691,N_18492);
or U20825 (N_20825,N_18558,N_18531);
nor U20826 (N_20826,N_16384,N_17801);
nor U20827 (N_20827,N_16197,N_17550);
nor U20828 (N_20828,N_16443,N_15635);
nand U20829 (N_20829,N_17489,N_15061);
nor U20830 (N_20830,N_18038,N_18427);
and U20831 (N_20831,N_15915,N_15025);
or U20832 (N_20832,N_19079,N_18631);
and U20833 (N_20833,N_19077,N_17262);
or U20834 (N_20834,N_16170,N_15410);
nor U20835 (N_20835,N_15124,N_19463);
or U20836 (N_20836,N_16688,N_19660);
nand U20837 (N_20837,N_16606,N_18778);
xor U20838 (N_20838,N_19199,N_18894);
nand U20839 (N_20839,N_18753,N_15684);
nand U20840 (N_20840,N_17058,N_15422);
or U20841 (N_20841,N_19641,N_15717);
nand U20842 (N_20842,N_17711,N_15352);
or U20843 (N_20843,N_19597,N_17794);
nand U20844 (N_20844,N_16998,N_18604);
nor U20845 (N_20845,N_19030,N_15991);
xor U20846 (N_20846,N_15460,N_16440);
or U20847 (N_20847,N_19770,N_18539);
or U20848 (N_20848,N_19417,N_16790);
nor U20849 (N_20849,N_15482,N_15989);
and U20850 (N_20850,N_18470,N_18400);
nor U20851 (N_20851,N_15318,N_16319);
and U20852 (N_20852,N_17600,N_15322);
nor U20853 (N_20853,N_15181,N_17001);
nor U20854 (N_20854,N_18098,N_18639);
nor U20855 (N_20855,N_15581,N_15170);
and U20856 (N_20856,N_16808,N_15105);
or U20857 (N_20857,N_17859,N_15247);
xnor U20858 (N_20858,N_18573,N_19388);
xnor U20859 (N_20859,N_16684,N_17906);
nand U20860 (N_20860,N_17338,N_18353);
nor U20861 (N_20861,N_16397,N_16475);
nor U20862 (N_20862,N_17530,N_15681);
nor U20863 (N_20863,N_18285,N_19885);
nor U20864 (N_20864,N_19439,N_15518);
xor U20865 (N_20865,N_16254,N_17244);
nand U20866 (N_20866,N_18578,N_15394);
nand U20867 (N_20867,N_19681,N_16905);
nor U20868 (N_20868,N_17552,N_19138);
xor U20869 (N_20869,N_19223,N_17035);
nand U20870 (N_20870,N_18119,N_19968);
and U20871 (N_20871,N_18111,N_17267);
nand U20872 (N_20872,N_19894,N_17034);
and U20873 (N_20873,N_15068,N_15118);
nor U20874 (N_20874,N_15975,N_19669);
xnor U20875 (N_20875,N_16991,N_18363);
xnor U20876 (N_20876,N_19619,N_15346);
or U20877 (N_20877,N_15250,N_19593);
xor U20878 (N_20878,N_15876,N_19784);
nor U20879 (N_20879,N_18333,N_18954);
xnor U20880 (N_20880,N_16091,N_17389);
nor U20881 (N_20881,N_19241,N_17050);
or U20882 (N_20882,N_15634,N_19467);
and U20883 (N_20883,N_18553,N_19948);
and U20884 (N_20884,N_16809,N_16023);
or U20885 (N_20885,N_16291,N_19416);
xnor U20886 (N_20886,N_17160,N_15151);
xor U20887 (N_20887,N_15531,N_16647);
nand U20888 (N_20888,N_15734,N_17245);
xnor U20889 (N_20889,N_15688,N_17974);
or U20890 (N_20890,N_16599,N_19506);
nand U20891 (N_20891,N_19425,N_16778);
nor U20892 (N_20892,N_18986,N_16922);
or U20893 (N_20893,N_16680,N_19823);
or U20894 (N_20894,N_17829,N_17879);
or U20895 (N_20895,N_18676,N_19236);
or U20896 (N_20896,N_19107,N_15955);
xor U20897 (N_20897,N_16032,N_16065);
nor U20898 (N_20898,N_17950,N_19197);
nor U20899 (N_20899,N_19434,N_16558);
nor U20900 (N_20900,N_15498,N_19461);
and U20901 (N_20901,N_18525,N_18255);
or U20902 (N_20902,N_16775,N_17570);
nor U20903 (N_20903,N_18585,N_15262);
and U20904 (N_20904,N_17323,N_17126);
nor U20905 (N_20905,N_17186,N_15267);
xor U20906 (N_20906,N_17415,N_18491);
nand U20907 (N_20907,N_19021,N_17703);
nor U20908 (N_20908,N_17596,N_16191);
nand U20909 (N_20909,N_15809,N_16464);
nand U20910 (N_20910,N_19728,N_17128);
or U20911 (N_20911,N_16453,N_19343);
or U20912 (N_20912,N_17233,N_18053);
and U20913 (N_20913,N_15142,N_16411);
or U20914 (N_20914,N_18507,N_15638);
and U20915 (N_20915,N_19367,N_17954);
or U20916 (N_20916,N_15461,N_15776);
and U20917 (N_20917,N_18915,N_18196);
nor U20918 (N_20918,N_18514,N_15665);
or U20919 (N_20919,N_16073,N_18993);
and U20920 (N_20920,N_17853,N_18822);
nor U20921 (N_20921,N_18953,N_15076);
or U20922 (N_20922,N_15711,N_19368);
and U20923 (N_20923,N_19549,N_18617);
xnor U20924 (N_20924,N_17593,N_19599);
and U20925 (N_20925,N_19808,N_18728);
nand U20926 (N_20926,N_17735,N_15202);
nor U20927 (N_20927,N_16828,N_19754);
or U20928 (N_20928,N_19526,N_19798);
xor U20929 (N_20929,N_16425,N_19172);
and U20930 (N_20930,N_18455,N_17546);
xor U20931 (N_20931,N_15565,N_15934);
nand U20932 (N_20932,N_19472,N_18654);
nor U20933 (N_20933,N_19692,N_16629);
xor U20934 (N_20934,N_15501,N_18620);
and U20935 (N_20935,N_17070,N_19276);
or U20936 (N_20936,N_17435,N_19565);
and U20937 (N_20937,N_15429,N_15645);
nand U20938 (N_20938,N_16123,N_15102);
and U20939 (N_20939,N_19957,N_17173);
nand U20940 (N_20940,N_18569,N_19755);
nand U20941 (N_20941,N_18526,N_19256);
or U20942 (N_20942,N_18278,N_16712);
nand U20943 (N_20943,N_16473,N_19861);
nor U20944 (N_20944,N_15660,N_18659);
or U20945 (N_20945,N_17709,N_16488);
or U20946 (N_20946,N_19924,N_18831);
and U20947 (N_20947,N_18256,N_19473);
xnor U20948 (N_20948,N_15280,N_17607);
nor U20949 (N_20949,N_17512,N_16215);
or U20950 (N_20950,N_17886,N_18032);
nand U20951 (N_20951,N_17644,N_17009);
and U20952 (N_20952,N_16085,N_19108);
xnor U20953 (N_20953,N_19207,N_15408);
and U20954 (N_20954,N_18934,N_15550);
and U20955 (N_20955,N_18374,N_17577);
nand U20956 (N_20956,N_16570,N_16585);
or U20957 (N_20957,N_17642,N_16119);
and U20958 (N_20958,N_17108,N_19366);
or U20959 (N_20959,N_18799,N_16328);
nand U20960 (N_20960,N_19571,N_17329);
and U20961 (N_20961,N_17578,N_17793);
xnor U20962 (N_20962,N_16836,N_19493);
xnor U20963 (N_20963,N_19721,N_15579);
and U20964 (N_20964,N_15673,N_19275);
or U20965 (N_20965,N_18052,N_16223);
or U20966 (N_20966,N_18832,N_15843);
nand U20967 (N_20967,N_19499,N_19800);
nor U20968 (N_20968,N_17631,N_15395);
nor U20969 (N_20969,N_15825,N_15654);
nand U20970 (N_20970,N_17744,N_15601);
and U20971 (N_20971,N_19945,N_15174);
xor U20972 (N_20972,N_17134,N_18850);
nand U20973 (N_20973,N_19117,N_17657);
xor U20974 (N_20974,N_18189,N_17156);
nand U20975 (N_20975,N_19181,N_19336);
xnor U20976 (N_20976,N_15440,N_16351);
and U20977 (N_20977,N_15953,N_16058);
nand U20978 (N_20978,N_16194,N_15569);
or U20979 (N_20979,N_19934,N_16520);
nand U20980 (N_20980,N_15764,N_15029);
xor U20981 (N_20981,N_15669,N_18009);
and U20982 (N_20982,N_17646,N_18682);
nand U20983 (N_20983,N_19458,N_19286);
nand U20984 (N_20984,N_16679,N_17384);
nand U20985 (N_20985,N_16370,N_18238);
nand U20986 (N_20986,N_16994,N_17706);
xor U20987 (N_20987,N_17984,N_18136);
xor U20988 (N_20988,N_18645,N_18626);
and U20989 (N_20989,N_19164,N_16251);
xnor U20990 (N_20990,N_18751,N_15468);
or U20991 (N_20991,N_16718,N_17321);
and U20992 (N_20992,N_17251,N_16003);
and U20993 (N_20993,N_15966,N_19600);
xor U20994 (N_20994,N_16152,N_16757);
xnor U20995 (N_20995,N_15123,N_18100);
nand U20996 (N_20996,N_18406,N_15725);
or U20997 (N_20997,N_18725,N_17670);
nand U20998 (N_20998,N_18449,N_15533);
xnor U20999 (N_20999,N_18340,N_18195);
or U21000 (N_21000,N_17502,N_16149);
or U21001 (N_21001,N_19932,N_16935);
or U21002 (N_21002,N_17041,N_17898);
nor U21003 (N_21003,N_16711,N_15033);
xnor U21004 (N_21004,N_18180,N_19614);
nand U21005 (N_21005,N_17343,N_15541);
xnor U21006 (N_21006,N_15706,N_19415);
xnor U21007 (N_21007,N_16158,N_19437);
nor U21008 (N_21008,N_19073,N_17588);
xnor U21009 (N_21009,N_18065,N_16059);
or U21010 (N_21010,N_17062,N_15166);
or U21011 (N_21011,N_19262,N_19347);
or U21012 (N_21012,N_18425,N_17615);
and U21013 (N_21013,N_19997,N_19725);
and U21014 (N_21014,N_19210,N_15238);
xnor U21015 (N_21015,N_19570,N_19773);
or U21016 (N_21016,N_19238,N_15887);
nand U21017 (N_21017,N_19746,N_19412);
nor U21018 (N_21018,N_17724,N_18485);
nand U21019 (N_21019,N_16826,N_17737);
nor U21020 (N_21020,N_15679,N_15559);
and U21021 (N_21021,N_15899,N_19349);
nand U21022 (N_21022,N_15821,N_18697);
xnor U21023 (N_21023,N_15310,N_15554);
nand U21024 (N_21024,N_16589,N_18869);
xnor U21025 (N_21025,N_18396,N_17284);
and U21026 (N_21026,N_18973,N_15824);
nand U21027 (N_21027,N_15499,N_16171);
and U21028 (N_21028,N_17511,N_15751);
or U21029 (N_21029,N_18433,N_16063);
nor U21030 (N_21030,N_19112,N_18708);
xnor U21031 (N_21031,N_19225,N_17743);
xor U21032 (N_21032,N_19699,N_17142);
xor U21033 (N_21033,N_15830,N_16601);
and U21034 (N_21034,N_15736,N_17764);
nor U21035 (N_21035,N_16726,N_17632);
and U21036 (N_21036,N_15957,N_17760);
nor U21037 (N_21037,N_16057,N_16557);
or U21038 (N_21038,N_18020,N_15046);
and U21039 (N_21039,N_17297,N_15532);
and U21040 (N_21040,N_15190,N_18185);
nand U21041 (N_21041,N_18624,N_19555);
or U21042 (N_21042,N_16897,N_16815);
xnor U21043 (N_21043,N_17000,N_18493);
xnor U21044 (N_21044,N_19292,N_15750);
and U21045 (N_21045,N_15391,N_16262);
nand U21046 (N_21046,N_15854,N_17784);
or U21047 (N_21047,N_16016,N_19279);
nand U21048 (N_21048,N_15413,N_15938);
xor U21049 (N_21049,N_15072,N_19805);
and U21050 (N_21050,N_19999,N_16309);
and U21051 (N_21051,N_17109,N_16667);
or U21052 (N_21052,N_17802,N_15980);
nand U21053 (N_21053,N_15567,N_17403);
nor U21054 (N_21054,N_19587,N_19038);
and U21055 (N_21055,N_17594,N_15762);
xor U21056 (N_21056,N_17376,N_16182);
and U21057 (N_21057,N_18512,N_19056);
nor U21058 (N_21058,N_18386,N_19903);
nand U21059 (N_21059,N_16445,N_19357);
xnor U21060 (N_21060,N_16933,N_16721);
xnor U21061 (N_21061,N_19383,N_16376);
xnor U21062 (N_21062,N_15528,N_15364);
and U21063 (N_21063,N_15842,N_17311);
nor U21064 (N_21064,N_16644,N_18582);
xnor U21065 (N_21065,N_15011,N_15807);
or U21066 (N_21066,N_15720,N_15483);
nand U21067 (N_21067,N_16207,N_15676);
and U21068 (N_21068,N_15997,N_15904);
nor U21069 (N_21069,N_17885,N_18420);
or U21070 (N_21070,N_16147,N_16840);
nor U21071 (N_21071,N_19023,N_16029);
nand U21072 (N_21072,N_17826,N_15169);
or U21073 (N_21073,N_15599,N_19606);
and U21074 (N_21074,N_17650,N_16634);
and U21075 (N_21075,N_18863,N_15163);
xnor U21076 (N_21076,N_18495,N_17966);
nand U21077 (N_21077,N_19850,N_19598);
nor U21078 (N_21078,N_18906,N_17271);
nor U21079 (N_21079,N_16222,N_19536);
nor U21080 (N_21080,N_15275,N_18365);
nand U21081 (N_21081,N_17391,N_15014);
xor U21082 (N_21082,N_17777,N_17804);
nand U21083 (N_21083,N_19436,N_16503);
or U21084 (N_21084,N_18685,N_16652);
and U21085 (N_21085,N_17258,N_17964);
and U21086 (N_21086,N_15092,N_15831);
or U21087 (N_21087,N_18548,N_15835);
xnor U21088 (N_21088,N_19028,N_19794);
xor U21089 (N_21089,N_18861,N_17619);
nand U21090 (N_21090,N_19019,N_15122);
or U21091 (N_21091,N_18208,N_15797);
nor U21092 (N_21092,N_18091,N_17038);
nor U21093 (N_21093,N_18840,N_18468);
xor U21094 (N_21094,N_16577,N_15767);
and U21095 (N_21095,N_18466,N_15508);
nor U21096 (N_21096,N_15874,N_15615);
nor U21097 (N_21097,N_17342,N_15135);
nor U21098 (N_21098,N_19274,N_15628);
or U21099 (N_21099,N_15928,N_19328);
nand U21100 (N_21100,N_16953,N_18959);
xnor U21101 (N_21101,N_15374,N_19460);
or U21102 (N_21102,N_17026,N_19205);
and U21103 (N_21103,N_18431,N_17892);
and U21104 (N_21104,N_18380,N_15798);
nor U21105 (N_21105,N_15650,N_16881);
nor U21106 (N_21106,N_19085,N_16470);
and U21107 (N_21107,N_18674,N_17878);
and U21108 (N_21108,N_17521,N_15811);
or U21109 (N_21109,N_15386,N_19745);
nor U21110 (N_21110,N_17025,N_16172);
and U21111 (N_21111,N_16517,N_17992);
xnor U21112 (N_21112,N_18877,N_19031);
nand U21113 (N_21113,N_17881,N_18809);
nor U21114 (N_21114,N_17375,N_18170);
xnor U21115 (N_21115,N_16133,N_15340);
and U21116 (N_21116,N_18299,N_16343);
or U21117 (N_21117,N_15709,N_17145);
xor U21118 (N_21118,N_15080,N_19342);
and U21119 (N_21119,N_18768,N_17807);
nor U21120 (N_21120,N_16761,N_18418);
xor U21121 (N_21121,N_19973,N_16281);
xnor U21122 (N_21122,N_16393,N_17852);
nand U21123 (N_21123,N_16109,N_18204);
xnor U21124 (N_21124,N_18339,N_17408);
or U21125 (N_21125,N_17372,N_19929);
nor U21126 (N_21126,N_16272,N_17069);
nand U21127 (N_21127,N_15649,N_19827);
nand U21128 (N_21128,N_15894,N_18292);
xnor U21129 (N_21129,N_18481,N_15009);
or U21130 (N_21130,N_17690,N_16478);
nor U21131 (N_21131,N_19637,N_18892);
nor U21132 (N_21132,N_16104,N_16584);
xor U21133 (N_21133,N_16310,N_17292);
and U21134 (N_21134,N_19537,N_18279);
nand U21135 (N_21135,N_17075,N_17567);
nand U21136 (N_21136,N_17752,N_15556);
xor U21137 (N_21137,N_17092,N_15578);
nand U21138 (N_21138,N_19200,N_18769);
nor U21139 (N_21139,N_17347,N_18188);
and U21140 (N_21140,N_19174,N_15530);
nor U21141 (N_21141,N_19306,N_16247);
nor U21142 (N_21142,N_16364,N_19010);
nand U21143 (N_21143,N_16526,N_15510);
nand U21144 (N_21144,N_17030,N_18975);
and U21145 (N_21145,N_17249,N_19501);
nor U21146 (N_21146,N_18094,N_17449);
nor U21147 (N_21147,N_15462,N_15458);
nand U21148 (N_21148,N_15295,N_18826);
xor U21149 (N_21149,N_19666,N_19532);
nor U21150 (N_21150,N_16683,N_19080);
or U21151 (N_21151,N_18914,N_16888);
nand U21152 (N_21152,N_19475,N_16792);
nand U21153 (N_21153,N_17424,N_17055);
and U21154 (N_21154,N_16014,N_16621);
or U21155 (N_21155,N_19562,N_17102);
nand U21156 (N_21156,N_18207,N_19560);
nor U21157 (N_21157,N_19553,N_16301);
or U21158 (N_21158,N_19528,N_19513);
xor U21159 (N_21159,N_19867,N_19163);
and U21160 (N_21160,N_18272,N_17361);
and U21161 (N_21161,N_18890,N_18102);
and U21162 (N_21162,N_16385,N_17220);
xnor U21163 (N_21163,N_19788,N_15756);
and U21164 (N_21164,N_19700,N_17135);
xnor U21165 (N_21165,N_15610,N_18452);
or U21166 (N_21166,N_15205,N_15180);
nor U21167 (N_21167,N_19469,N_15609);
or U21168 (N_21168,N_19991,N_15263);
and U21169 (N_21169,N_17604,N_15156);
nand U21170 (N_21170,N_15158,N_19756);
nor U21171 (N_21171,N_17671,N_19486);
or U21172 (N_21172,N_17263,N_17792);
and U21173 (N_21173,N_18644,N_17531);
or U21174 (N_21174,N_15985,N_19627);
xnor U21175 (N_21175,N_17351,N_19086);
and U21176 (N_21176,N_15418,N_15526);
or U21177 (N_21177,N_16781,N_17235);
or U21178 (N_21178,N_18813,N_16246);
nor U21179 (N_21179,N_18033,N_17446);
and U21180 (N_21180,N_16415,N_17800);
and U21181 (N_21181,N_17757,N_17049);
and U21182 (N_21182,N_19487,N_19419);
xor U21183 (N_21183,N_18335,N_16900);
and U21184 (N_21184,N_15207,N_17872);
nor U21185 (N_21185,N_19156,N_16938);
and U21186 (N_21186,N_18696,N_18307);
xor U21187 (N_21187,N_17788,N_16446);
nand U21188 (N_21188,N_18334,N_19339);
nor U21189 (N_21189,N_19068,N_17503);
xor U21190 (N_21190,N_19775,N_19235);
nor U21191 (N_21191,N_17017,N_17473);
nor U21192 (N_21192,N_19771,N_16050);
and U21193 (N_21193,N_19115,N_15155);
and U21194 (N_21194,N_17891,N_19642);
xor U21195 (N_21195,N_18910,N_15336);
or U21196 (N_21196,N_15879,N_15870);
or U21197 (N_21197,N_18440,N_17566);
and U21198 (N_21198,N_15266,N_19060);
nand U21199 (N_21199,N_18356,N_16866);
nand U21200 (N_21200,N_19615,N_18634);
nand U21201 (N_21201,N_19872,N_16734);
and U21202 (N_21202,N_16618,N_15175);
and U21203 (N_21203,N_15411,N_19137);
or U21204 (N_21204,N_19132,N_17658);
nor U21205 (N_21205,N_18994,N_18629);
and U21206 (N_21206,N_19704,N_17374);
xnor U21207 (N_21207,N_18483,N_15536);
or U21208 (N_21208,N_18733,N_18836);
xor U21209 (N_21209,N_18146,N_16593);
nor U21210 (N_21210,N_19640,N_16608);
xor U21211 (N_21211,N_18857,N_17904);
nor U21212 (N_21212,N_19435,N_15509);
nor U21213 (N_21213,N_17601,N_17513);
or U21214 (N_21214,N_17054,N_18717);
nor U21215 (N_21215,N_19958,N_18692);
nor U21216 (N_21216,N_19689,N_17341);
and U21217 (N_21217,N_15334,N_15803);
nand U21218 (N_21218,N_16399,N_15426);
or U21219 (N_21219,N_18853,N_18516);
or U21220 (N_21220,N_16923,N_17621);
or U21221 (N_21221,N_19430,N_17908);
nand U21222 (N_21222,N_19365,N_18504);
xnor U21223 (N_21223,N_16853,N_15770);
nand U21224 (N_21224,N_16837,N_15139);
xnor U21225 (N_21225,N_16699,N_17780);
xnor U21226 (N_21226,N_17762,N_15289);
nand U21227 (N_21227,N_17023,N_18067);
nand U21228 (N_21228,N_17584,N_17592);
nor U21229 (N_21229,N_19329,N_18731);
nor U21230 (N_21230,N_16212,N_15838);
nand U21231 (N_21231,N_16431,N_15777);
and U21232 (N_21232,N_17696,N_19870);
or U21233 (N_21233,N_19875,N_17515);
or U21234 (N_21234,N_17401,N_17532);
xor U21235 (N_21235,N_15801,N_15630);
or U21236 (N_21236,N_16737,N_16208);
nor U21237 (N_21237,N_16423,N_16729);
nand U21238 (N_21238,N_15553,N_16318);
xnor U21239 (N_21239,N_16132,N_16919);
xnor U21240 (N_21240,N_19157,N_16722);
and U21241 (N_21241,N_18966,N_19819);
xnor U21242 (N_21242,N_18167,N_19128);
nor U21243 (N_21243,N_15006,N_17212);
nor U21244 (N_21244,N_19013,N_15409);
xnor U21245 (N_21245,N_18166,N_15273);
xnor U21246 (N_21246,N_17630,N_18771);
or U21247 (N_21247,N_17628,N_19716);
or U21248 (N_21248,N_16121,N_18003);
nor U21249 (N_21249,N_18622,N_18770);
xor U21250 (N_21250,N_18152,N_16436);
xnor U21251 (N_21251,N_18068,N_18128);
nand U21252 (N_21252,N_19399,N_19851);
nand U21253 (N_21253,N_17330,N_17914);
or U21254 (N_21254,N_17133,N_17820);
or U21255 (N_21255,N_18698,N_19201);
and U21256 (N_21256,N_16651,N_15259);
or U21257 (N_21257,N_19535,N_18385);
and U21258 (N_21258,N_15950,N_18312);
nor U21259 (N_21259,N_19917,N_15455);
nor U21260 (N_21260,N_17569,N_17609);
nor U21261 (N_21261,N_17370,N_17453);
nor U21262 (N_21262,N_15527,N_16516);
nand U21263 (N_21263,N_17087,N_19249);
and U21264 (N_21264,N_16265,N_18103);
and U21265 (N_21265,N_18945,N_18414);
or U21266 (N_21266,N_18037,N_15466);
or U21267 (N_21267,N_15368,N_19705);
nor U21268 (N_21268,N_18928,N_16180);
and U21269 (N_21269,N_17900,N_16564);
nand U21270 (N_21270,N_17131,N_15219);
and U21271 (N_21271,N_17146,N_15371);
xnor U21272 (N_21272,N_17006,N_15927);
and U21273 (N_21273,N_17194,N_16116);
xor U21274 (N_21274,N_19041,N_16452);
and U21275 (N_21275,N_19305,N_15194);
or U21276 (N_21276,N_16789,N_17279);
and U21277 (N_21277,N_17180,N_17718);
nor U21278 (N_21278,N_17506,N_16227);
nor U21279 (N_21279,N_19050,N_19993);
xor U21280 (N_21280,N_18841,N_16233);
nor U21281 (N_21281,N_15577,N_19285);
or U21282 (N_21282,N_17639,N_16080);
or U21283 (N_21283,N_17028,N_18022);
and U21284 (N_21284,N_19001,N_18652);
and U21285 (N_21285,N_19824,N_17294);
or U21286 (N_21286,N_15303,N_15138);
xor U21287 (N_21287,N_15157,N_15658);
or U21288 (N_21288,N_19153,N_16486);
nor U21289 (N_21289,N_17371,N_16969);
and U21290 (N_21290,N_16968,N_17018);
and U21291 (N_21291,N_16444,N_16401);
or U21292 (N_21292,N_19969,N_19766);
nor U21293 (N_21293,N_18641,N_15078);
nand U21294 (N_21294,N_18942,N_18752);
or U21295 (N_21295,N_15134,N_17996);
nor U21296 (N_21296,N_19440,N_15150);
and U21297 (N_21297,N_19317,N_19398);
and U21298 (N_21298,N_17821,N_19710);
nand U21299 (N_21299,N_18941,N_19760);
nor U21300 (N_21300,N_15432,N_15924);
nand U21301 (N_21301,N_17925,N_15730);
xor U21302 (N_21302,N_18007,N_18282);
nand U21303 (N_21303,N_17863,N_17367);
nand U21304 (N_21304,N_19921,N_16690);
nor U21305 (N_21305,N_19686,N_18309);
nand U21306 (N_21306,N_19101,N_19691);
nand U21307 (N_21307,N_19379,N_19715);
and U21308 (N_21308,N_15042,N_17962);
nor U21309 (N_21309,N_16750,N_18891);
and U21310 (N_21310,N_16595,N_19896);
and U21311 (N_21311,N_18759,N_18715);
nand U21312 (N_21312,N_17359,N_18301);
xor U21313 (N_21313,N_19179,N_16240);
xor U21314 (N_21314,N_16627,N_16363);
nor U21315 (N_21315,N_16920,N_18287);
or U21316 (N_21316,N_17880,N_18740);
nand U21317 (N_21317,N_18628,N_15671);
xnor U21318 (N_21318,N_18603,N_17355);
nor U21319 (N_21319,N_18723,N_18519);
or U21320 (N_21320,N_15742,N_15407);
xor U21321 (N_21321,N_17786,N_19530);
or U21322 (N_21322,N_15034,N_17307);
or U21323 (N_21323,N_19131,N_19129);
and U21324 (N_21324,N_19695,N_18134);
or U21325 (N_21325,N_16500,N_19362);
nand U21326 (N_21326,N_16835,N_18538);
or U21327 (N_21327,N_16967,N_17612);
or U21328 (N_21328,N_17841,N_18090);
and U21329 (N_21329,N_16944,N_17119);
xnor U21330 (N_21330,N_15570,N_18327);
or U21331 (N_21331,N_16089,N_18651);
and U21332 (N_21332,N_16966,N_18957);
and U21333 (N_21333,N_15517,N_17673);
and U21334 (N_21334,N_17702,N_19009);
or U21335 (N_21335,N_18996,N_16410);
or U21336 (N_21336,N_16914,N_19173);
xnor U21337 (N_21337,N_18889,N_18907);
or U21338 (N_21338,N_17253,N_17960);
and U21339 (N_21339,N_18667,N_18590);
nor U21340 (N_21340,N_19284,N_18258);
and U21341 (N_21341,N_16624,N_16860);
or U21342 (N_21342,N_18592,N_17536);
or U21343 (N_21343,N_18347,N_19466);
and U21344 (N_21344,N_16572,N_17103);
and U21345 (N_21345,N_18373,N_18323);
or U21346 (N_21346,N_19061,N_16653);
xnor U21347 (N_21347,N_16820,N_18995);
xor U21348 (N_21348,N_15956,N_18198);
or U21349 (N_21349,N_16375,N_18179);
nand U21350 (N_21350,N_18843,N_19395);
nand U21351 (N_21351,N_19110,N_18422);
nand U21352 (N_21352,N_17366,N_17809);
or U21353 (N_21353,N_15959,N_17884);
nand U21354 (N_21354,N_16934,N_18936);
or U21355 (N_21355,N_18511,N_18290);
nand U21356 (N_21356,N_19470,N_15149);
nor U21357 (N_21357,N_15406,N_16360);
nand U21358 (N_21358,N_18902,N_17765);
and U21359 (N_21359,N_16153,N_17947);
or U21360 (N_21360,N_15513,N_19912);
or U21361 (N_21361,N_19866,N_15585);
nand U21362 (N_21362,N_17951,N_18532);
nand U21363 (N_21363,N_15926,N_18348);
xnor U21364 (N_21364,N_18713,N_16887);
xnor U21365 (N_21365,N_15771,N_18922);
xor U21366 (N_21366,N_15802,N_18673);
or U21367 (N_21367,N_16633,N_16545);
or U21368 (N_21368,N_16071,N_18463);
nor U21369 (N_21369,N_17452,N_15903);
and U21370 (N_21370,N_16554,N_16156);
and U21371 (N_21371,N_15485,N_17171);
and U21372 (N_21372,N_17206,N_15438);
nand U21373 (N_21373,N_16838,N_15885);
nor U21374 (N_21374,N_17159,N_17339);
nand U21375 (N_21375,N_17534,N_17191);
nor U21376 (N_21376,N_16741,N_19787);
and U21377 (N_21377,N_18460,N_19065);
nor U21378 (N_21378,N_17414,N_19718);
and U21379 (N_21379,N_17624,N_17605);
nor U21380 (N_21380,N_17164,N_18543);
or U21381 (N_21381,N_15719,N_15489);
and U21382 (N_21382,N_19456,N_15128);
and U21383 (N_21383,N_19777,N_16818);
nand U21384 (N_21384,N_16745,N_16731);
nand U21385 (N_21385,N_18739,N_15748);
or U21386 (N_21386,N_15430,N_19198);
or U21387 (N_21387,N_18416,N_15781);
nand U21388 (N_21388,N_19733,N_18872);
nand U21389 (N_21389,N_19257,N_18635);
xor U21390 (N_21390,N_15000,N_17172);
xor U21391 (N_21391,N_17169,N_15710);
nand U21392 (N_21392,N_17242,N_19384);
and U21393 (N_21393,N_18454,N_15216);
nand U21394 (N_21394,N_19252,N_15434);
nor U21395 (N_21395,N_18346,N_16324);
and U21396 (N_21396,N_18656,N_15971);
xor U21397 (N_21397,N_19998,N_18006);
xor U21398 (N_21398,N_16075,N_19226);
nor U21399 (N_21399,N_17312,N_16259);
nor U21400 (N_21400,N_19070,N_17295);
nand U21401 (N_21401,N_16694,N_18379);
xnor U21402 (N_21402,N_16361,N_18328);
xor U21403 (N_21403,N_15757,N_17537);
or U21404 (N_21404,N_18854,N_15886);
xor U21405 (N_21405,N_18848,N_16243);
or U21406 (N_21406,N_16936,N_16643);
xor U21407 (N_21407,N_17218,N_16986);
xor U21408 (N_21408,N_17928,N_19083);
or U21409 (N_21409,N_19564,N_19548);
xor U21410 (N_21410,N_15162,N_16128);
or U21411 (N_21411,N_17656,N_17967);
or U21412 (N_21412,N_18121,N_18837);
or U21413 (N_21413,N_16366,N_19111);
xnor U21414 (N_21414,N_15705,N_16592);
nor U21415 (N_21415,N_18616,N_17256);
xor U21416 (N_21416,N_15027,N_16862);
or U21417 (N_21417,N_18169,N_18490);
nor U21418 (N_21418,N_15212,N_17072);
nor U21419 (N_21419,N_17756,N_16079);
or U21420 (N_21420,N_18803,N_19591);
or U21421 (N_21421,N_19255,N_15891);
xor U21422 (N_21422,N_19579,N_17921);
or U21423 (N_21423,N_17850,N_19595);
or U21424 (N_21424,N_19862,N_19045);
xor U21425 (N_21425,N_19693,N_16879);
or U21426 (N_21426,N_15875,N_18313);
nor U21427 (N_21427,N_18413,N_15549);
or U21428 (N_21428,N_18775,N_18233);
nor U21429 (N_21429,N_15850,N_16111);
nand U21430 (N_21430,N_17704,N_15652);
nand U21431 (N_21431,N_17591,N_18939);
and U21432 (N_21432,N_16947,N_18382);
xor U21433 (N_21433,N_17965,N_16285);
nor U21434 (N_21434,N_19303,N_16293);
nor U21435 (N_21435,N_18987,N_16135);
and U21436 (N_21436,N_16970,N_17422);
and U21437 (N_21437,N_15979,N_15325);
or U21438 (N_21438,N_16992,N_17373);
or U21439 (N_21439,N_18824,N_17407);
and U21440 (N_21440,N_19448,N_19203);
xnor U21441 (N_21441,N_18475,N_18412);
or U21442 (N_21442,N_17629,N_16242);
nand U21443 (N_21443,N_16441,N_18903);
or U21444 (N_21444,N_19443,N_19939);
and U21445 (N_21445,N_15378,N_18500);
xnor U21446 (N_21446,N_16800,N_19651);
and U21447 (N_21447,N_15693,N_19731);
xnor U21448 (N_21448,N_16753,N_18870);
or U21449 (N_21449,N_15160,N_18737);
xor U21450 (N_21450,N_16067,N_19049);
nand U21451 (N_21451,N_17061,N_15007);
nor U21452 (N_21452,N_19984,N_19928);
nor U21453 (N_21453,N_18451,N_17915);
xor U21454 (N_21454,N_18779,N_16993);
or U21455 (N_21455,N_17647,N_16915);
or U21456 (N_21456,N_16847,N_16248);
xnor U21457 (N_21457,N_16535,N_15399);
nor U21458 (N_21458,N_19227,N_17662);
or U21459 (N_21459,N_17909,N_15276);
nor U21460 (N_21460,N_17959,N_17738);
nand U21461 (N_21461,N_16451,N_15662);
nand U21462 (N_21462,N_18486,N_17636);
nor U21463 (N_21463,N_16674,N_19188);
and U21464 (N_21464,N_17797,N_19909);
nor U21465 (N_21465,N_18678,N_18880);
nor U21466 (N_21466,N_16687,N_19161);
nor U21467 (N_21467,N_15321,N_16733);
nor U21468 (N_21468,N_18642,N_18439);
nor U21469 (N_21469,N_15548,N_15257);
xor U21470 (N_21470,N_15052,N_17469);
and U21471 (N_21471,N_16528,N_16396);
or U21472 (N_21472,N_18064,N_17470);
xnor U21473 (N_21473,N_15869,N_15986);
or U21474 (N_21474,N_18043,N_19752);
and U21475 (N_21475,N_15345,N_19977);
and U21476 (N_21476,N_16145,N_19569);
and U21477 (N_21477,N_15145,N_15258);
nor U21478 (N_21478,N_15062,N_18900);
and U21479 (N_21479,N_17864,N_16356);
xor U21480 (N_21480,N_16426,N_15552);
xor U21481 (N_21481,N_15215,N_19708);
or U21482 (N_21482,N_19222,N_16159);
or U21483 (N_21483,N_16961,N_17353);
nand U21484 (N_21484,N_18533,N_16975);
xor U21485 (N_21485,N_15488,N_17051);
or U21486 (N_21486,N_19516,N_15301);
and U21487 (N_21487,N_16196,N_18322);
and U21488 (N_21488,N_19309,N_16884);
nand U21489 (N_21489,N_16590,N_19589);
and U21490 (N_21490,N_17769,N_17660);
and U21491 (N_21491,N_17082,N_17929);
nor U21492 (N_21492,N_16736,N_17763);
nand U21493 (N_21493,N_16290,N_16582);
xor U21494 (N_21494,N_15331,N_18820);
or U21495 (N_21495,N_19703,N_16819);
xnor U21496 (N_21496,N_17116,N_15330);
nor U21497 (N_21497,N_17107,N_15868);
nand U21498 (N_21498,N_19876,N_18459);
nand U21499 (N_21499,N_15176,N_15127);
nand U21500 (N_21500,N_19465,N_17059);
nand U21501 (N_21501,N_18245,N_16428);
nor U21502 (N_21502,N_15366,N_16457);
xnor U21503 (N_21503,N_16911,N_15791);
nor U21504 (N_21504,N_17597,N_18508);
xnor U21505 (N_21505,N_15116,N_15733);
or U21506 (N_21506,N_18601,N_18763);
nor U21507 (N_21507,N_18888,N_16336);
and U21508 (N_21508,N_17618,N_15707);
xnor U21509 (N_21509,N_15187,N_15253);
and U21510 (N_21510,N_18664,N_17890);
nor U21511 (N_21511,N_15557,N_16547);
and U21512 (N_21512,N_18467,N_15668);
nand U21513 (N_21513,N_16903,N_17346);
or U21514 (N_21514,N_18684,N_15841);
nand U21515 (N_21515,N_17441,N_15220);
nand U21516 (N_21516,N_15094,N_16013);
nand U21517 (N_21517,N_15065,N_18001);
nand U21518 (N_21518,N_19251,N_18772);
or U21519 (N_21519,N_15670,N_18638);
or U21520 (N_21520,N_18886,N_17560);
nor U21521 (N_21521,N_17088,N_17130);
or U21522 (N_21522,N_17280,N_19762);
and U21523 (N_21523,N_16605,N_19243);
xor U21524 (N_21524,N_15402,N_19268);
and U21525 (N_21525,N_17021,N_16859);
nor U21526 (N_21526,N_19135,N_19547);
or U21527 (N_21527,N_18375,N_15769);
or U21528 (N_21528,N_15978,N_16392);
or U21529 (N_21529,N_15132,N_19916);
or U21530 (N_21530,N_15981,N_17803);
and U21531 (N_21531,N_19834,N_19018);
nand U21532 (N_21532,N_16822,N_16720);
xnor U21533 (N_21533,N_19678,N_19220);
xor U21534 (N_21534,N_16660,N_18849);
and U21535 (N_21535,N_16339,N_18079);
nor U21536 (N_21536,N_18130,N_18441);
nand U21537 (N_21537,N_16404,N_15584);
xnor U21538 (N_21538,N_19502,N_19055);
xnor U21539 (N_21539,N_18417,N_16124);
nor U21540 (N_21540,N_17516,N_17335);
nand U21541 (N_21541,N_16282,N_19034);
or U21542 (N_21542,N_17076,N_18611);
nand U21543 (N_21543,N_16656,N_18961);
nand U21544 (N_21544,N_16983,N_17561);
nor U21545 (N_21545,N_15755,N_17426);
xnor U21546 (N_21546,N_19213,N_15558);
or U21547 (N_21547,N_18295,N_16561);
or U21548 (N_21548,N_19727,N_15735);
and U21549 (N_21549,N_17491,N_16061);
or U21550 (N_21550,N_18078,N_15456);
and U21551 (N_21551,N_15018,N_18905);
or U21552 (N_21552,N_16882,N_16924);
xnor U21553 (N_21553,N_17423,N_16877);
nand U21554 (N_21554,N_19610,N_16631);
and U21555 (N_21555,N_19802,N_16489);
or U21556 (N_21556,N_17275,N_19298);
and U21557 (N_21557,N_15376,N_19064);
or U21558 (N_21558,N_19300,N_17549);
or U21559 (N_21559,N_19785,N_19818);
nor U21560 (N_21560,N_19826,N_16654);
xor U21561 (N_21561,N_16974,N_18411);
xor U21562 (N_21562,N_16954,N_15206);
nand U21563 (N_21563,N_17538,N_18724);
xor U21564 (N_21564,N_17755,N_15433);
or U21565 (N_21565,N_18588,N_19494);
nor U21566 (N_21566,N_16030,N_19421);
nor U21567 (N_21567,N_15507,N_15828);
xor U21568 (N_21568,N_15883,N_18583);
nor U21569 (N_21569,N_18783,N_15414);
nor U21570 (N_21570,N_15090,N_16257);
and U21571 (N_21571,N_16098,N_19880);
xnor U21572 (N_21572,N_19753,N_18707);
xor U21573 (N_21573,N_18887,N_17983);
and U21574 (N_21574,N_18378,N_15249);
xor U21575 (N_21575,N_15063,N_18700);
xor U21576 (N_21576,N_16555,N_17047);
and U21577 (N_21577,N_16797,N_17418);
or U21578 (N_21578,N_18153,N_17400);
and U21579 (N_21579,N_16144,N_17648);
nor U21580 (N_21580,N_15931,N_17637);
and U21581 (N_21581,N_15343,N_18041);
and U21582 (N_21582,N_19675,N_19943);
nand U21583 (N_21583,N_19761,N_18300);
and U21584 (N_21584,N_16092,N_18613);
xnor U21585 (N_21585,N_17084,N_18748);
or U21586 (N_21586,N_19029,N_19854);
nand U21587 (N_21587,N_17856,N_15621);
nor U21588 (N_21588,N_17541,N_19768);
nor U21589 (N_21589,N_18097,N_18878);
or U21590 (N_21590,N_19586,N_15451);
xor U21591 (N_21591,N_18670,N_15256);
xnor U21592 (N_21592,N_18320,N_18390);
nor U21593 (N_21593,N_19002,N_16492);
and U21594 (N_21594,N_19835,N_16082);
or U21595 (N_21595,N_19451,N_19638);
and U21596 (N_21596,N_16772,N_19908);
nor U21597 (N_21597,N_19449,N_19654);
and U21598 (N_21598,N_18694,N_19983);
xnor U21599 (N_21599,N_18760,N_17603);
xor U21600 (N_21600,N_15888,N_17870);
or U21601 (N_21601,N_18089,N_17840);
and U21602 (N_21602,N_19078,N_17542);
nor U21603 (N_21603,N_17074,N_15070);
nand U21604 (N_21604,N_16368,N_18288);
and U21605 (N_21605,N_17205,N_15317);
and U21606 (N_21606,N_17969,N_15316);
and U21607 (N_21607,N_16387,N_15837);
or U21608 (N_21608,N_16039,N_17456);
nor U21609 (N_21609,N_17494,N_15941);
nor U21610 (N_21610,N_19481,N_18625);
nor U21611 (N_21611,N_17846,N_17695);
nor U21612 (N_21612,N_15773,N_17677);
nand U21613 (N_21613,N_19947,N_18794);
nor U21614 (N_21614,N_15463,N_19734);
or U21615 (N_21615,N_19295,N_19674);
and U21616 (N_21616,N_17818,N_15307);
and U21617 (N_21617,N_17553,N_17147);
or U21618 (N_21618,N_17528,N_19545);
nor U21619 (N_21619,N_18541,N_15588);
nand U21620 (N_21620,N_19709,N_17012);
xnor U21621 (N_21621,N_19644,N_16982);
nand U21622 (N_21622,N_15313,N_16161);
nand U21623 (N_21623,N_17779,N_17556);
and U21624 (N_21624,N_17348,N_18807);
and U21625 (N_21625,N_15204,N_18436);
and U21626 (N_21626,N_15495,N_18371);
xnor U21627 (N_21627,N_16707,N_18392);
or U21628 (N_21628,N_19387,N_17585);
and U21629 (N_21629,N_15329,N_17337);
nor U21630 (N_21630,N_17935,N_16552);
or U21631 (N_21631,N_17888,N_18864);
xor U21632 (N_21632,N_19837,N_16373);
and U21633 (N_21633,N_17849,N_19575);
nor U21634 (N_21634,N_15586,N_19620);
and U21635 (N_21635,N_15481,N_16220);
nand U21636 (N_21636,N_15519,N_15380);
and U21637 (N_21637,N_18141,N_15296);
nand U21638 (N_21638,N_17913,N_17540);
and U21639 (N_21639,N_19840,N_15337);
xor U21640 (N_21640,N_17095,N_18913);
nor U21641 (N_21641,N_19113,N_19381);
and U21642 (N_21642,N_16143,N_16181);
or U21643 (N_21643,N_15443,N_18226);
nand U21644 (N_21644,N_19446,N_17250);
xnor U21645 (N_21645,N_19585,N_18839);
nand U21646 (N_21646,N_17056,N_15242);
nand U21647 (N_21647,N_18494,N_18341);
nor U21648 (N_21648,N_18680,N_16418);
and U21649 (N_21649,N_15021,N_19022);
and U21650 (N_21650,N_17573,N_19099);
xor U21651 (N_21651,N_17475,N_19900);
xor U21652 (N_21652,N_15107,N_18421);
or U21653 (N_21653,N_15724,N_17558);
nand U21654 (N_21654,N_16511,N_15505);
nand U21655 (N_21655,N_18658,N_18298);
nor U21656 (N_21656,N_15477,N_15743);
xnor U21657 (N_21657,N_16812,N_17255);
nand U21658 (N_21658,N_19956,N_18082);
and U21659 (N_21659,N_15143,N_16534);
xor U21660 (N_21660,N_17866,N_18244);
nand U21661 (N_21661,N_18896,N_15375);
xnor U21662 (N_21662,N_16313,N_19538);
nor U21663 (N_21663,N_18145,N_19063);
and U21664 (N_21664,N_18660,N_15789);
nor U21665 (N_21665,N_15494,N_17097);
nor U21666 (N_21666,N_16163,N_18529);
nand U21667 (N_21667,N_19039,N_17044);
and U21668 (N_21668,N_17395,N_19964);
or U21669 (N_21669,N_16886,N_18209);
xor U21670 (N_21670,N_19403,N_18911);
or U21671 (N_21671,N_19093,N_16578);
xnor U21672 (N_21672,N_16494,N_18871);
or U21673 (N_21673,N_17924,N_15075);
xor U21674 (N_21674,N_19749,N_17064);
nor U21675 (N_21675,N_19683,N_18669);
nand U21676 (N_21676,N_17053,N_16179);
xor U21677 (N_21677,N_15381,N_15227);
or U21678 (N_21678,N_17007,N_19889);
nor U21679 (N_21679,N_16068,N_15480);
xnor U21680 (N_21680,N_18236,N_18817);
or U21681 (N_21681,N_19959,N_17949);
xnor U21682 (N_21682,N_16229,N_17167);
xnor U21683 (N_21683,N_19682,N_16275);
nor U21684 (N_21684,N_16099,N_17861);
and U21685 (N_21685,N_16304,N_18156);
nand U21686 (N_21686,N_19905,N_17324);
nor U21687 (N_21687,N_19592,N_19828);
or U21688 (N_21688,N_18048,N_16519);
and U21689 (N_21689,N_18830,N_17464);
or U21690 (N_21690,N_16468,N_17882);
nor U21691 (N_21691,N_15183,N_16374);
xnor U21692 (N_21692,N_17580,N_15612);
or U21693 (N_21693,N_16793,N_15880);
nor U21694 (N_21694,N_18122,N_18021);
and U21695 (N_21695,N_18426,N_18370);
or U21696 (N_21696,N_16872,N_17318);
and U21697 (N_21697,N_15723,N_18345);
nor U21698 (N_21698,N_17386,N_15208);
and U21699 (N_21699,N_15647,N_17837);
nor U21700 (N_21700,N_16760,N_18458);
nand U21701 (N_21701,N_16696,N_17999);
nor U21702 (N_21702,N_17434,N_16665);
xor U21703 (N_21703,N_19653,N_15913);
nand U21704 (N_21704,N_17314,N_19394);
or U21705 (N_21705,N_19234,N_17231);
or U21706 (N_21706,N_15133,N_16773);
nand U21707 (N_21707,N_19248,N_15109);
nand U21708 (N_21708,N_19811,N_15198);
and U21709 (N_21709,N_15302,N_17240);
nor U21710 (N_21710,N_15437,N_16405);
nand U21711 (N_21711,N_17663,N_18203);
and U21712 (N_21712,N_16501,N_19237);
or U21713 (N_21713,N_15191,N_18862);
or U21714 (N_21714,N_15084,N_17572);
nand U21715 (N_21715,N_16846,N_19887);
nor U21716 (N_21716,N_16626,N_18570);
and U21717 (N_21717,N_19779,N_19806);
nor U21718 (N_21718,N_15543,N_15637);
and U21719 (N_21719,N_17776,N_18326);
nor U21720 (N_21720,N_17698,N_15792);
nor U21721 (N_21721,N_18077,N_15848);
xor U21722 (N_21722,N_16813,N_15304);
or U21723 (N_21723,N_17708,N_17741);
nand U21724 (N_21724,N_19492,N_17838);
or U21725 (N_21725,N_16025,N_16852);
and U21726 (N_21726,N_18376,N_18958);
nor U21727 (N_21727,N_16948,N_15195);
xnor U21728 (N_21728,N_18088,N_19789);
xnor U21729 (N_21729,N_15782,N_15492);
and U21730 (N_21730,N_19539,N_18261);
and U21731 (N_21731,N_18321,N_17895);
and U21732 (N_21732,N_17196,N_16956);
nor U21733 (N_21733,N_19027,N_15274);
xor U21734 (N_21734,N_16402,N_19169);
nor U21735 (N_21735,N_17100,N_19982);
xor U21736 (N_21736,N_17433,N_19442);
or U21737 (N_21737,N_16756,N_16640);
xnor U21738 (N_21738,N_19574,N_18405);
nor U21739 (N_21739,N_15228,N_17364);
and U21740 (N_21740,N_18443,N_17867);
and U21741 (N_21741,N_17344,N_15097);
nor U21742 (N_21742,N_17501,N_17029);
and U21743 (N_21743,N_18637,N_15270);
and U21744 (N_21744,N_17104,N_17081);
xor U21745 (N_21745,N_17814,N_19390);
nor U21746 (N_21746,N_17170,N_19706);
and U21747 (N_21747,N_17443,N_19098);
or U21748 (N_21748,N_18681,N_15444);
xor U21749 (N_21749,N_17229,N_18387);
and U21750 (N_21750,N_19820,N_19175);
or U21751 (N_21751,N_18649,N_19831);
xor U21752 (N_21752,N_16269,N_19146);
nand U21753 (N_21753,N_16335,N_18815);
xnor U21754 (N_21754,N_17086,N_18524);
and U21755 (N_21755,N_16350,N_17979);
nor U21756 (N_21756,N_17719,N_19319);
nor U21757 (N_21757,N_18758,N_17583);
or U21758 (N_21758,N_18612,N_19918);
or U21759 (N_21759,N_15473,N_18847);
xnor U21760 (N_21760,N_19992,N_15633);
and U21761 (N_21761,N_17162,N_19679);
nor U21762 (N_21762,N_17726,N_16461);
xnor U21763 (N_21763,N_15385,N_16889);
nor U21764 (N_21764,N_17684,N_19797);
nor U21765 (N_21765,N_18845,N_17917);
and U21766 (N_21766,N_17138,N_19432);
or U21767 (N_21767,N_16713,N_18579);
or U21768 (N_21768,N_16536,N_19869);
xnor U21769 (N_21769,N_16477,N_16394);
and U21770 (N_21770,N_15315,N_18932);
xnor U21771 (N_21771,N_15923,N_17369);
xor U21772 (N_21772,N_15112,N_18842);
xnor U21773 (N_21773,N_19829,N_18377);
xnor U21774 (N_21774,N_17939,N_15677);
xor U21775 (N_21775,N_19124,N_17858);
nor U21776 (N_21776,N_16776,N_18123);
or U21777 (N_21777,N_17445,N_15435);
and U21778 (N_21778,N_16239,N_15996);
and U21779 (N_21779,N_16649,N_16011);
xnor U21780 (N_21780,N_16571,N_16747);
xor U21781 (N_21781,N_19290,N_16001);
or U21782 (N_21782,N_19976,N_16958);
or U21783 (N_21783,N_17303,N_16450);
xor U21784 (N_21784,N_16748,N_17625);
nor U21785 (N_21785,N_19490,N_17893);
or U21786 (N_21786,N_17643,N_15765);
or U21787 (N_21787,N_19975,N_17442);
and U21788 (N_21788,N_16022,N_17111);
and U21789 (N_21789,N_19371,N_18219);
nand U21790 (N_21790,N_16107,N_16307);
xnor U21791 (N_21791,N_17961,N_17547);
or U21792 (N_21792,N_15269,N_18014);
nor U21793 (N_21793,N_17946,N_19781);
nand U21794 (N_21794,N_16698,N_16499);
and U21795 (N_21795,N_18991,N_19865);
and U21796 (N_21796,N_19769,N_16005);
and U21797 (N_21797,N_18257,N_17236);
and U21798 (N_21798,N_18186,N_18814);
xnor U21799 (N_21799,N_17518,N_16046);
xnor U21800 (N_21800,N_17602,N_16253);
or U21801 (N_21801,N_19335,N_16400);
nand U21802 (N_21802,N_15814,N_15039);
and U21803 (N_21803,N_15089,N_19299);
nor U21804 (N_21804,N_15759,N_17774);
xor U21805 (N_21805,N_17345,N_17083);
xor U21806 (N_21806,N_18105,N_18308);
nor U21807 (N_21807,N_16524,N_15860);
and U21808 (N_21808,N_15110,N_16855);
nor U21809 (N_21809,N_17221,N_17836);
nor U21810 (N_21810,N_18178,N_19863);
xnor U21811 (N_21811,N_19311,N_18355);
or U21812 (N_21812,N_17113,N_15236);
nor U21813 (N_21813,N_18229,N_16344);
nand U21814 (N_21814,N_19123,N_16018);
and U21815 (N_21815,N_18990,N_16714);
and U21816 (N_21816,N_18428,N_15545);
or U21817 (N_21817,N_19496,N_19556);
nor U21818 (N_21818,N_17161,N_18453);
nand U21819 (N_21819,N_16136,N_18835);
nand U21820 (N_21820,N_16814,N_19217);
and U21821 (N_21821,N_15184,N_15563);
nand U21822 (N_21822,N_15939,N_16600);
and U21823 (N_21823,N_18901,N_16299);
or U21824 (N_21824,N_15929,N_16380);
nor U21825 (N_21825,N_15095,N_19864);
or U21826 (N_21826,N_15144,N_16677);
nor U21827 (N_21827,N_16483,N_19369);
nand U21828 (N_21828,N_16052,N_19510);
and U21829 (N_21829,N_16827,N_15863);
nand U21830 (N_21830,N_19402,N_18784);
and U21831 (N_21831,N_19036,N_18343);
nor U21832 (N_21832,N_16976,N_16204);
xnor U21833 (N_21833,N_18099,N_19663);
nand U21834 (N_21834,N_15121,N_17123);
and U21835 (N_21835,N_15951,N_19962);
nand U21836 (N_21836,N_15726,N_18873);
nor U21837 (N_21837,N_16231,N_17973);
nor U21838 (N_21838,N_15291,N_16203);
and U21839 (N_21839,N_15002,N_18726);
and U21840 (N_21840,N_16117,N_19747);
nor U21841 (N_21841,N_15020,N_16550);
xor U21842 (N_21842,N_18838,N_19883);
nand U21843 (N_21843,N_18086,N_17616);
xnor U21844 (N_21844,N_16015,N_19744);
nand U21845 (N_21845,N_18589,N_19631);
and U21846 (N_21846,N_17544,N_15344);
nor U21847 (N_21847,N_16876,N_15918);
nor U21848 (N_21848,N_16407,N_16544);
nor U21849 (N_21849,N_19281,N_18139);
xnor U21850 (N_21850,N_17877,N_15196);
xor U21851 (N_21851,N_18462,N_18562);
and U21852 (N_21852,N_17485,N_15136);
xor U21853 (N_21853,N_15111,N_16715);
nor U21854 (N_21854,N_16625,N_19877);
or U21855 (N_21855,N_18241,N_15229);
and U21856 (N_21856,N_16673,N_15404);
and U21857 (N_21857,N_15323,N_15775);
nand U21858 (N_21858,N_18576,N_16594);
xnor U21859 (N_21859,N_16609,N_18448);
or U21860 (N_21860,N_19269,N_15255);
and U21861 (N_21861,N_16377,N_16689);
nand U21862 (N_21862,N_17579,N_17729);
xnor U21863 (N_21863,N_15013,N_19680);
nor U21864 (N_21864,N_17394,N_19879);
or U21865 (N_21865,N_19322,N_19427);
xnor U21866 (N_21866,N_16540,N_16616);
nand U21867 (N_21867,N_18429,N_19546);
or U21868 (N_21868,N_18899,N_15704);
nand U21869 (N_21869,N_19059,N_19406);
and U21870 (N_21870,N_17697,N_17941);
xnor U21871 (N_21871,N_17685,N_18971);
and U21872 (N_21872,N_18762,N_15045);
or U21873 (N_21873,N_16076,N_18399);
xor U21874 (N_21874,N_17857,N_15012);
xor U21875 (N_21875,N_17486,N_19719);
nand U21876 (N_21876,N_18437,N_15119);
xor U21877 (N_21877,N_16771,N_17098);
xnor U21878 (N_21878,N_15562,N_15449);
nand U21879 (N_21879,N_16692,N_19429);
and U21880 (N_21880,N_17508,N_16787);
nor U21881 (N_21881,N_17633,N_19359);
and U21882 (N_21882,N_17716,N_19628);
xor U21883 (N_21883,N_16758,N_15984);
nand U21884 (N_21884,N_18220,N_19410);
and U21885 (N_21885,N_15172,N_17581);
nor U21886 (N_21886,N_15627,N_17955);
xnor U21887 (N_21887,N_17832,N_18789);
xor U21888 (N_21888,N_18154,N_15788);
nand U21889 (N_21889,N_16280,N_17705);
and U21890 (N_21890,N_19656,N_19261);
nand U21891 (N_21891,N_15547,N_19247);
nand U21892 (N_21892,N_15293,N_16784);
xor U21893 (N_21893,N_19216,N_15846);
or U21894 (N_21894,N_17031,N_18192);
nor U21895 (N_21895,N_17043,N_19318);
xnor U21896 (N_21896,N_16202,N_17438);
and U21897 (N_21897,N_15049,N_17843);
and U21898 (N_21898,N_19937,N_19994);
and U21899 (N_21899,N_19024,N_17077);
xnor U21900 (N_21900,N_15044,N_19507);
xnor U21901 (N_21901,N_19126,N_18791);
and U21902 (N_21902,N_16657,N_19810);
nand U21903 (N_21903,N_19980,N_19920);
or U21904 (N_21904,N_16751,N_17358);
xnor U21905 (N_21905,N_15239,N_19212);
nor U21906 (N_21906,N_19266,N_18044);
nand U21907 (N_21907,N_16295,N_15472);
nor U21908 (N_21908,N_19853,N_15148);
and U21909 (N_21909,N_19750,N_18535);
nor U21910 (N_21910,N_18360,N_19512);
nor U21911 (N_21911,N_15933,N_18253);
or U21912 (N_21912,N_19088,N_15620);
nand U21913 (N_21913,N_15503,N_18668);
xor U21914 (N_21914,N_19176,N_16562);
and U21915 (N_21915,N_16867,N_19550);
nand U21916 (N_21916,N_18788,N_16100);
or U21917 (N_21917,N_17665,N_17299);
nand U21918 (N_21918,N_15362,N_15593);
xnor U21919 (N_21919,N_19596,N_19326);
xnor U21920 (N_21920,N_18302,N_18316);
and U21921 (N_21921,N_15906,N_18977);
or U21922 (N_21922,N_15522,N_18461);
nand U21923 (N_21923,N_17860,N_18231);
and U21924 (N_21924,N_15987,N_16513);
xor U21925 (N_21925,N_16353,N_15697);
nand U21926 (N_21926,N_19149,N_15790);
xnor U21927 (N_21927,N_19974,N_15287);
and U21928 (N_21928,N_19229,N_18269);
or U21929 (N_21929,N_16638,N_16743);
nand U21930 (N_21930,N_17487,N_17230);
xor U21931 (N_21931,N_19474,N_18935);
nor U21932 (N_21932,N_17873,N_19844);
and U21933 (N_21933,N_17835,N_18144);
or U21934 (N_21934,N_15059,N_18969);
nand U21935 (N_21935,N_18201,N_17261);
nor U21936 (N_21936,N_15859,N_17168);
nor U21937 (N_21937,N_15871,N_18968);
or U21938 (N_21938,N_19673,N_19520);
and U21939 (N_21939,N_16530,N_17143);
nor U21940 (N_21940,N_16928,N_17332);
or U21941 (N_21941,N_15235,N_17399);
or U21942 (N_21942,N_18710,N_19833);
nor U21943 (N_21943,N_18364,N_16796);
or U21944 (N_21944,N_15153,N_17177);
nand U21945 (N_21945,N_15189,N_16424);
nand U21946 (N_21946,N_18126,N_15490);
nand U21947 (N_21947,N_15829,N_19629);
or U21948 (N_21948,N_15140,N_16752);
nor U21949 (N_21949,N_18741,N_15278);
xor U21950 (N_21950,N_17127,N_18730);
or U21951 (N_21951,N_18663,N_19178);
or U21952 (N_21952,N_16048,N_19897);
nor U21953 (N_21953,N_18792,N_18742);
nand U21954 (N_21954,N_17184,N_16017);
and U21955 (N_21955,N_19182,N_18035);
and U21956 (N_21956,N_17894,N_18549);
xor U21957 (N_21957,N_19114,N_15678);
nor U21958 (N_21958,N_19890,N_17722);
nand U21959 (N_21959,N_16256,N_18224);
and U21960 (N_21960,N_19471,N_19047);
nand U21961 (N_21961,N_15252,N_19096);
nand U21962 (N_21962,N_17758,N_19874);
nor U21963 (N_21963,N_17215,N_18161);
nand U21964 (N_21964,N_18834,N_17406);
nor U21965 (N_21965,N_16637,N_18176);
nand U21966 (N_21966,N_15967,N_15093);
nand U21967 (N_21967,N_18248,N_15067);
nor U21968 (N_21968,N_18747,N_15892);
nor U21969 (N_21969,N_15421,N_18101);
or U21970 (N_21970,N_15954,N_19325);
nor U21971 (N_21971,N_15244,N_16211);
or U21972 (N_21972,N_19557,N_19738);
nand U21973 (N_21973,N_18545,N_17626);
nor U21974 (N_21974,N_16989,N_17568);
xor U21975 (N_21975,N_16710,N_16234);
and U21976 (N_21976,N_16697,N_19159);
or U21977 (N_21977,N_18434,N_15363);
nor U21978 (N_21978,N_19450,N_18980);
nand U21979 (N_21979,N_19214,N_17739);
nand U21980 (N_21980,N_18173,N_17472);
nor U21981 (N_21981,N_18057,N_17019);
or U21982 (N_21982,N_19938,N_17936);
xnor U21983 (N_21983,N_15940,N_17223);
or U21984 (N_21984,N_15655,N_19670);
or U21985 (N_21985,N_19621,N_16709);
xor U21986 (N_21986,N_15905,N_15377);
nor U21987 (N_21987,N_17465,N_16805);
nand U21988 (N_21988,N_17916,N_17411);
or U21989 (N_21989,N_17796,N_18610);
or U21990 (N_21990,N_16830,N_16034);
and U21991 (N_21991,N_16078,N_15103);
and U21992 (N_21992,N_19902,N_18916);
xor U21993 (N_21993,N_18780,N_16495);
xnor U21994 (N_21994,N_18711,N_15357);
xnor U21995 (N_21995,N_17682,N_19783);
nand U21996 (N_21996,N_18856,N_17227);
nor U21997 (N_21997,N_17224,N_18650);
nor U21998 (N_21998,N_18109,N_16427);
and U21999 (N_21999,N_16541,N_18215);
xor U22000 (N_22000,N_18358,N_15486);
and U22001 (N_22001,N_19215,N_18736);
or U22002 (N_22002,N_17519,N_15605);
xnor U22003 (N_22003,N_19316,N_18797);
and U22004 (N_22004,N_19698,N_16270);
nor U22005 (N_22005,N_18005,N_16129);
and U22006 (N_22006,N_18614,N_18636);
xor U22007 (N_22007,N_16026,N_19914);
xnor U22008 (N_22008,N_16297,N_16658);
nor U22009 (N_22009,N_17862,N_17987);
nor U22010 (N_22010,N_15942,N_19726);
or U22011 (N_22011,N_18540,N_15539);
and U22012 (N_22012,N_17429,N_18133);
or U22013 (N_22013,N_15728,N_19219);
xor U22014 (N_22014,N_17692,N_18087);
nand U22015 (N_22015,N_16355,N_16549);
and U22016 (N_22016,N_17080,N_19522);
xor U22017 (N_22017,N_16245,N_17723);
nand U22018 (N_22018,N_16449,N_18478);
or U22019 (N_22019,N_16213,N_15073);
nand U22020 (N_22020,N_16455,N_16289);
nor U22021 (N_22021,N_18833,N_16044);
or U22022 (N_22022,N_17190,N_19092);
nand U22023 (N_22023,N_18083,N_15910);
nor U22024 (N_22024,N_16563,N_19452);
xnor U22025 (N_22025,N_16095,N_16333);
nand U22026 (N_22026,N_18546,N_16037);
nand U22027 (N_22027,N_18106,N_16607);
or U22028 (N_22028,N_15001,N_17976);
nor U22029 (N_22029,N_15820,N_15211);
nand U22030 (N_22030,N_18800,N_15010);
nand U22031 (N_22031,N_18110,N_19361);
and U22032 (N_22032,N_15651,N_17787);
nor U22033 (N_22033,N_17248,N_16786);
xnor U22034 (N_22034,N_16072,N_16386);
nor U22035 (N_22035,N_18574,N_18823);
nor U22036 (N_22036,N_16192,N_18242);
and U22037 (N_22037,N_18946,N_18271);
or U22038 (N_22038,N_18499,N_16266);
and U22039 (N_22039,N_15491,N_16326);
and U22040 (N_22040,N_18859,N_17748);
nor U22041 (N_22041,N_17559,N_17855);
nor U22042 (N_22042,N_16096,N_19594);
xnor U22043 (N_22043,N_16306,N_17014);
or U22044 (N_22044,N_19477,N_16187);
nand U22045 (N_22045,N_18402,N_18675);
nand U22046 (N_22046,N_18162,N_15086);
and U22047 (N_22047,N_15087,N_17112);
and U22048 (N_22048,N_19014,N_16456);
and U22049 (N_22049,N_15574,N_18199);
xor U22050 (N_22050,N_16154,N_18394);
xnor U22051 (N_22051,N_19103,N_17413);
and U22052 (N_22052,N_17040,N_16028);
and U22053 (N_22053,N_15873,N_19931);
nand U22054 (N_22054,N_17141,N_16338);
xor U22055 (N_22055,N_18523,N_17309);
nand U22056 (N_22056,N_18621,N_19180);
nor U22057 (N_22057,N_18267,N_17889);
and U22058 (N_22058,N_18874,N_18013);
nor U22059 (N_22059,N_19302,N_15470);
nor U22060 (N_22060,N_19370,N_16596);
nand U22061 (N_22061,N_18310,N_16261);
or U22062 (N_22062,N_19563,N_19988);
or U22063 (N_22063,N_16851,N_16480);
xor U22064 (N_22064,N_16972,N_19648);
nor U22065 (N_22065,N_15261,N_18947);
xnor U22066 (N_22066,N_16510,N_19608);
and U22067 (N_22067,N_18071,N_15126);
or U22068 (N_22068,N_16094,N_16342);
nand U22069 (N_22069,N_17354,N_19356);
and U22070 (N_22070,N_16460,N_15804);
xor U22071 (N_22071,N_16904,N_19447);
nor U22072 (N_22072,N_19839,N_15349);
and U22073 (N_22073,N_18025,N_18884);
xor U22074 (N_22074,N_19140,N_16560);
or U22075 (N_22075,N_15845,N_16810);
or U22076 (N_22076,N_16190,N_15930);
nand U22077 (N_22077,N_16833,N_19062);
and U22078 (N_22078,N_17211,N_15551);
and U22079 (N_22079,N_16043,N_19489);
nor U22080 (N_22080,N_19051,N_15607);
or U22081 (N_22081,N_19601,N_16131);
xor U22082 (N_22082,N_16521,N_16064);
xnor U22083 (N_22083,N_19504,N_16538);
or U22084 (N_22084,N_19672,N_19965);
and U22085 (N_22085,N_17291,N_18812);
and U22086 (N_22086,N_19386,N_18506);
and U22087 (N_22087,N_19206,N_15281);
nor U22088 (N_22088,N_18575,N_16330);
nor U22089 (N_22089,N_19667,N_15367);
and U22090 (N_22090,N_15019,N_18948);
nor U22091 (N_22091,N_19260,N_19878);
and U22092 (N_22092,N_16122,N_19639);
nand U22093 (N_22093,N_18714,N_16502);
xnor U22094 (N_22094,N_17016,N_18264);
and U22095 (N_22095,N_15680,N_17634);
or U22096 (N_22096,N_18630,N_19521);
nand U22097 (N_22097,N_17664,N_16946);
nand U22098 (N_22098,N_19796,N_16010);
or U22099 (N_22099,N_18000,N_17934);
nand U22100 (N_22100,N_16277,N_19658);
nand U22101 (N_22101,N_17813,N_15146);
xnor U22102 (N_22102,N_15768,N_19616);
and U22103 (N_22103,N_17509,N_16012);
and U22104 (N_22104,N_15209,N_15935);
nor U22105 (N_22105,N_19664,N_18804);
nor U22106 (N_22106,N_17493,N_15218);
xor U22107 (N_22107,N_16036,N_17686);
and U22108 (N_22108,N_16706,N_18787);
or U22109 (N_22109,N_17931,N_16439);
and U22110 (N_22110,N_16476,N_18349);
and U22111 (N_22111,N_17666,N_15243);
nand U22112 (N_22112,N_17772,N_19320);
or U22113 (N_22113,N_16169,N_18970);
xor U22114 (N_22114,N_18522,N_19376);
nor U22115 (N_22115,N_16019,N_19732);
nor U22116 (N_22116,N_18391,N_15056);
and U22117 (N_22117,N_17247,N_16165);
and U22118 (N_22118,N_16264,N_17839);
and U22119 (N_22119,N_16389,N_19830);
or U22120 (N_22120,N_16705,N_16537);
nor U22121 (N_22121,N_17204,N_17499);
and U22122 (N_22122,N_16300,N_19772);
nand U22123 (N_22123,N_15800,N_19612);
nand U22124 (N_22124,N_19860,N_18952);
xor U22125 (N_22125,N_17188,N_16000);
nor U22126 (N_22126,N_16610,N_15178);
or U22127 (N_22127,N_18530,N_15032);
xor U22128 (N_22128,N_16769,N_19391);
xnor U22129 (N_22129,N_19816,N_19459);
xnor U22130 (N_22130,N_15847,N_19713);
nand U22131 (N_22131,N_16009,N_15643);
and U22132 (N_22132,N_15972,N_19524);
nand U22133 (N_22133,N_16620,N_15232);
xnor U22134 (N_22134,N_17847,N_16973);
and U22135 (N_22135,N_16945,N_16070);
and U22136 (N_22136,N_18940,N_17390);
nor U22137 (N_22137,N_17587,N_18924);
and U22138 (N_22138,N_18096,N_18055);
and U22139 (N_22139,N_19996,N_15308);
or U22140 (N_22140,N_15108,N_15613);
nor U22141 (N_22141,N_16454,N_17582);
nand U22142 (N_22142,N_15917,N_15976);
nor U22143 (N_22143,N_17239,N_17483);
nand U22144 (N_22144,N_17919,N_15641);
or U22145 (N_22145,N_15695,N_18324);
nand U22146 (N_22146,N_17174,N_19380);
and U22147 (N_22147,N_17458,N_18289);
nand U22148 (N_22148,N_15727,N_15618);
xnor U22149 (N_22149,N_16664,N_17806);
xnor U22150 (N_22150,N_17896,N_15515);
and U22151 (N_22151,N_19067,N_17265);
nand U22152 (N_22152,N_18671,N_16329);
or U22153 (N_22153,N_19856,N_16398);
and U22154 (N_22154,N_18028,N_16551);
and U22155 (N_22155,N_15365,N_17013);
xnor U22156 (N_22156,N_16311,N_19913);
xor U22157 (N_22157,N_17340,N_19454);
or U22158 (N_22158,N_16232,N_18712);
or U22159 (N_22159,N_15179,N_16157);
xnor U22160 (N_22160,N_17020,N_19652);
xnor U22161 (N_22161,N_19040,N_18254);
nor U22162 (N_22162,N_16346,N_15004);
nand U22163 (N_22163,N_18132,N_16118);
xor U22164 (N_22164,N_16579,N_15024);
or U22165 (N_22165,N_18591,N_17589);
or U22166 (N_22166,N_19267,N_19782);
and U22167 (N_22167,N_18227,N_16505);
or U22168 (N_22168,N_19491,N_15520);
nand U22169 (N_22169,N_17476,N_16650);
nor U22170 (N_22170,N_17024,N_16918);
xor U22171 (N_22171,N_18963,N_15692);
or U22172 (N_22172,N_17495,N_18471);
nor U22173 (N_22173,N_16321,N_18252);
nand U22174 (N_22174,N_15721,N_15914);
nor U22175 (N_22175,N_17254,N_16617);
or U22176 (N_22176,N_16573,N_17288);
nor U22177 (N_22177,N_17217,N_15853);
or U22178 (N_22178,N_18844,N_15200);
nor U22179 (N_22179,N_18895,N_19702);
and U22180 (N_22180,N_19377,N_18318);
or U22181 (N_22181,N_18164,N_17302);
nor U22182 (N_22182,N_16325,N_18217);
or U22183 (N_22183,N_16763,N_18683);
xnor U22184 (N_22184,N_18283,N_19373);
nor U22185 (N_22185,N_16471,N_15816);
or U22186 (N_22186,N_17978,N_15254);
or U22187 (N_22187,N_18593,N_16315);
xnor U22188 (N_22188,N_15037,N_15591);
nor U22189 (N_22189,N_15944,N_18338);
and U22190 (N_22190,N_19814,N_15054);
nor U22191 (N_22191,N_17320,N_17120);
and U22192 (N_22192,N_16047,N_16834);
and U22193 (N_22193,N_17590,N_19989);
or U22194 (N_22194,N_19483,N_19301);
nor U22195 (N_22195,N_18149,N_17105);
xor U22196 (N_22196,N_16176,N_19886);
nor U22197 (N_22197,N_17933,N_18868);
xnor U22198 (N_22198,N_15415,N_15787);
nor U22199 (N_22199,N_15514,N_15305);
xnor U22200 (N_22200,N_18270,N_15982);
xor U22201 (N_22201,N_18537,N_16416);
nand U22202 (N_22202,N_17742,N_17972);
or U22203 (N_22203,N_16848,N_18137);
or U22204 (N_22204,N_17094,N_16816);
nor U22205 (N_22205,N_16056,N_18568);
nor U22206 (N_22206,N_19327,N_19455);
nor U22207 (N_22207,N_17993,N_17052);
nand U22208 (N_22208,N_15326,N_15881);
nand U22209 (N_22209,N_19576,N_16951);
nand U22210 (N_22210,N_18745,N_15912);
xnor U22211 (N_22211,N_19677,N_16632);
and U22212 (N_22212,N_18923,N_18250);
nand U22213 (N_22213,N_19649,N_17274);
nand U22214 (N_22214,N_18072,N_19330);
xnor U22215 (N_22215,N_16200,N_18720);
and U22216 (N_22216,N_17228,N_16522);
and U22217 (N_22217,N_18184,N_19462);
nor U22218 (N_22218,N_18557,N_15754);
nor U22219 (N_22219,N_16303,N_18518);
and U22220 (N_22220,N_16950,N_19519);
and U22221 (N_22221,N_19892,N_18018);
xnor U22222 (N_22222,N_19581,N_17712);
nand U22223 (N_22223,N_16523,N_15231);
nand U22224 (N_22224,N_19185,N_17140);
or U22225 (N_22225,N_18361,N_16105);
nand U22226 (N_22226,N_15919,N_19476);
xnor U22227 (N_22227,N_19662,N_18865);
nand U22228 (N_22228,N_16422,N_15974);
nor U22229 (N_22229,N_17195,N_15827);
xor U22230 (N_22230,N_19165,N_18174);
and U22231 (N_22231,N_16162,N_18351);
nand U22232 (N_22232,N_16811,N_18828);
or U22233 (N_22233,N_15222,N_15947);
nor U22234 (N_22234,N_15066,N_17197);
or U22235 (N_22235,N_18017,N_15497);
nor U22236 (N_22236,N_18921,N_18118);
nor U22237 (N_22237,N_18331,N_19868);
nor U22238 (N_22238,N_16053,N_18766);
nor U22239 (N_22239,N_16214,N_16619);
nand U22240 (N_22240,N_17759,N_19720);
and U22241 (N_22241,N_17653,N_18757);
or U22242 (N_22242,N_19847,N_15694);
or U22243 (N_22243,N_17387,N_19961);
nand U22244 (N_22244,N_18275,N_17927);
nor U22245 (N_22245,N_16168,N_17208);
or U22246 (N_22246,N_18498,N_16614);
xor U22247 (N_22247,N_19724,N_19240);
nand U22248 (N_22248,N_17681,N_16186);
and U22249 (N_22249,N_15961,N_19155);
nor U22250 (N_22250,N_16352,N_17319);
xor U22251 (N_22251,N_19287,N_19730);
and U22252 (N_22252,N_17720,N_18200);
nand U22253 (N_22253,N_16432,N_15712);
nor U22254 (N_22254,N_15600,N_17998);
and U22255 (N_22255,N_15476,N_17260);
and U22256 (N_22256,N_16661,N_16930);
or U22257 (N_22257,N_16166,N_16979);
or U22258 (N_22258,N_19453,N_19534);
or U22259 (N_22259,N_16648,N_17305);
or U22260 (N_22260,N_19152,N_19617);
nor U22261 (N_22261,N_16249,N_15390);
and U22262 (N_22262,N_18964,N_17300);
or U22263 (N_22263,N_15096,N_17989);
nand U22264 (N_22264,N_16146,N_19283);
xor U22265 (N_22265,N_15031,N_18210);
nand U22266 (N_22266,N_18542,N_19444);
nor U22267 (N_22267,N_17425,N_17952);
nor U22268 (N_22268,N_17651,N_18908);
xor U22269 (N_22269,N_16323,N_15833);
nor U22270 (N_22270,N_15661,N_17775);
and U22271 (N_22271,N_16296,N_17595);
nand U22272 (N_22272,N_19263,N_19119);
or U22273 (N_22273,N_17380,N_17232);
and U22274 (N_22274,N_19389,N_17844);
or U22275 (N_22275,N_16198,N_18469);
nand U22276 (N_22276,N_18294,N_19233);
nand U22277 (N_22277,N_18816,N_19006);
xnor U22278 (N_22278,N_17484,N_19542);
nand U22279 (N_22279,N_19685,N_17901);
xor U22280 (N_22280,N_16383,N_17121);
nor U22281 (N_22281,N_17903,N_16102);
and U22282 (N_22282,N_15749,N_17237);
xor U22283 (N_22283,N_15699,N_16880);
nor U22284 (N_22284,N_15849,N_19011);
nand U22285 (N_22285,N_19405,N_15595);
nor U22286 (N_22286,N_19759,N_18395);
xor U22287 (N_22287,N_15702,N_16409);
nand U22288 (N_22288,N_19026,N_18061);
and U22289 (N_22289,N_18010,N_18214);
nand U22290 (N_22290,N_16802,N_15805);
xnor U22291 (N_22291,N_15383,N_19433);
nand U22292 (N_22292,N_17117,N_19457);
or U22293 (N_22293,N_16978,N_18821);
xor U22294 (N_22294,N_19253,N_19095);
or U22295 (N_22295,N_15995,N_18509);
nand U22296 (N_22296,N_19141,N_17812);
nand U22297 (N_22297,N_16357,N_15041);
or U22298 (N_22298,N_19942,N_19393);
or U22299 (N_22299,N_16858,N_15064);
nor U22300 (N_22300,N_16183,N_17678);
xor U22301 (N_22301,N_19091,N_18045);
or U22302 (N_22302,N_17830,N_17203);
or U22303 (N_22303,N_18825,N_19665);
and U22304 (N_22304,N_17883,N_18563);
and U22305 (N_22305,N_15629,N_16964);
and U22306 (N_22306,N_17599,N_15085);
nor U22307 (N_22307,N_16566,N_19953);
and U22308 (N_22308,N_19058,N_16331);
nand U22309 (N_22309,N_16378,N_16663);
nand U22310 (N_22310,N_17015,N_16340);
and U22311 (N_22311,N_15416,N_15625);
xnor U22312 (N_22312,N_17736,N_17363);
or U22313 (N_22313,N_19202,N_19758);
nor U22314 (N_22314,N_15115,N_15537);
or U22315 (N_22315,N_16940,N_18260);
nor U22316 (N_22316,N_16770,N_17071);
nor U22317 (N_22317,N_16490,N_18719);
nor U22318 (N_22318,N_18456,N_19344);
nor U22319 (N_22319,N_15686,N_16611);
nor U22320 (N_22320,N_17085,N_16367);
and U22321 (N_22321,N_16002,N_16173);
nor U22322 (N_22322,N_19891,N_18194);
or U22323 (N_22323,N_15648,N_17688);
xnor U22324 (N_22324,N_18988,N_18397);
nor U22325 (N_22325,N_16224,N_17732);
and U22326 (N_22326,N_15226,N_15506);
nor U22327 (N_22327,N_18230,N_19351);
or U22328 (N_22328,N_18030,N_17766);
nor U22329 (N_22329,N_17440,N_17930);
nand U22330 (N_22330,N_18547,N_16337);
or U22331 (N_22331,N_16672,N_16693);
or U22332 (N_22332,N_18703,N_19162);
xor U22333 (N_22333,N_16762,N_15487);
xnor U22334 (N_22334,N_18409,N_18202);
or U22335 (N_22335,N_18827,N_18488);
nor U22336 (N_22336,N_17975,N_18750);
nand U22337 (N_22337,N_17357,N_19568);
xnor U22338 (N_22338,N_16997,N_16381);
nand U22339 (N_22339,N_17874,N_16783);
or U22340 (N_22340,N_16702,N_19960);
and U22341 (N_22341,N_19158,N_19192);
xnor U22342 (N_22342,N_17046,N_17079);
and U22343 (N_22343,N_15772,N_19231);
xnor U22344 (N_22344,N_16719,N_18008);
xor U22345 (N_22345,N_15393,N_18846);
xor U22346 (N_22346,N_19000,N_19121);
xnor U22347 (N_22347,N_19972,N_15895);
nand U22348 (N_22348,N_17507,N_17746);
xnor U22349 (N_22349,N_19239,N_18019);
nand U22350 (N_22350,N_17940,N_17045);
xnor U22351 (N_22351,N_17963,N_18665);
or U22352 (N_22352,N_19795,N_18027);
xor U22353 (N_22353,N_18926,N_19170);
nor U22354 (N_22354,N_17734,N_18357);
or U22355 (N_22355,N_15060,N_19786);
xor U22356 (N_22356,N_19657,N_17869);
or U22357 (N_22357,N_16414,N_17139);
and U22358 (N_22358,N_15819,N_16081);
nand U22359 (N_22359,N_18151,N_18687);
nand U22360 (N_22360,N_19923,N_16302);
or U22361 (N_22361,N_17136,N_19130);
and U22362 (N_22362,N_17420,N_16320);
nand U22363 (N_22363,N_19646,N_17455);
xnor U22364 (N_22364,N_18175,N_16201);
nor U22365 (N_22365,N_16108,N_16412);
nor U22366 (N_22366,N_18075,N_18985);
and U22367 (N_22367,N_17238,N_16662);
and U22368 (N_22368,N_15582,N_19763);
nand U22369 (N_22369,N_15949,N_19881);
xnor U22370 (N_22370,N_17922,N_16622);
and U22371 (N_22371,N_19037,N_17985);
xnor U22372 (N_22372,N_15210,N_15867);
nand U22373 (N_22373,N_17381,N_18938);
or U22374 (N_22374,N_17899,N_19741);
or U22375 (N_22375,N_19729,N_16912);
and U22376 (N_22376,N_17731,N_18344);
nor U22377 (N_22377,N_19043,N_15040);
nor U22378 (N_22378,N_19353,N_19007);
xnor U22379 (N_22379,N_19561,N_18424);
or U22380 (N_22380,N_19003,N_17576);
and U22381 (N_22381,N_16349,N_18482);
xnor U22382 (N_22382,N_17868,N_18489);
nor U22383 (N_22383,N_18131,N_16874);
and U22384 (N_22384,N_16093,N_17574);
nand U22385 (N_22385,N_19517,N_18704);
nand U22386 (N_22386,N_18997,N_17492);
or U22387 (N_22387,N_15088,N_18909);
or U22388 (N_22388,N_18515,N_19313);
nand U22389 (N_22389,N_16542,N_15823);
xor U22390 (N_22390,N_17467,N_15603);
nand U22391 (N_22391,N_18107,N_15852);
nand U22392 (N_22392,N_15808,N_15657);
xnor U22393 (N_22393,N_15611,N_19838);
and U22394 (N_22394,N_18031,N_18138);
xor U22395 (N_22395,N_17649,N_16742);
and U22396 (N_22396,N_15598,N_18829);
and U22397 (N_22397,N_16943,N_18368);
xor U22398 (N_22398,N_15246,N_18632);
nand U22399 (N_22399,N_15785,N_17627);
or U22400 (N_22400,N_17481,N_17285);
and U22401 (N_22401,N_19071,N_18933);
or U22402 (N_22402,N_19944,N_16754);
nand U22403 (N_22403,N_19523,N_16863);
or U22404 (N_22404,N_16167,N_16218);
xor U22405 (N_22405,N_19422,N_15165);
and U22406 (N_22406,N_16686,N_15384);
nor U22407 (N_22407,N_15786,N_18917);
nor U22408 (N_22408,N_15454,N_19882);
nor U22409 (N_22409,N_15716,N_19588);
or U22410 (N_22410,N_19480,N_19852);
or U22411 (N_22411,N_18480,N_15500);
xor U22412 (N_22412,N_17555,N_18384);
nand U22413 (N_22413,N_19025,N_15822);
xor U22414 (N_22414,N_18795,N_16112);
nor U22415 (N_22415,N_17713,N_16433);
or U22416 (N_22416,N_18743,N_17700);
nor U22417 (N_22417,N_17613,N_16746);
and U22418 (N_22418,N_16317,N_18206);
nor U22419 (N_22419,N_17282,N_19807);
or U22420 (N_22420,N_15666,N_17745);
nor U22421 (N_22421,N_19822,N_15427);
nor U22422 (N_22422,N_19661,N_17520);
or U22423 (N_22423,N_16891,N_18855);
nor U22424 (N_22424,N_19291,N_15806);
xnor U22425 (N_22425,N_16913,N_16332);
nor U22426 (N_22426,N_15946,N_16955);
xor U22427 (N_22427,N_16305,N_19722);
nor U22428 (N_22428,N_15664,N_15309);
nand U22429 (N_22429,N_15861,N_19072);
xnor U22430 (N_22430,N_18262,N_16890);
nor U22431 (N_22431,N_19139,N_18213);
xnor U22432 (N_22432,N_15740,N_16892);
nor U22433 (N_22433,N_19577,N_15752);
or U22434 (N_22434,N_17416,N_18284);
nor U22435 (N_22435,N_16821,N_15596);
nand U22436 (N_22436,N_15297,N_16575);
or U22437 (N_22437,N_18627,N_16188);
nand U22438 (N_22438,N_19441,N_19097);
nand U22439 (N_22439,N_19355,N_16051);
nand U22440 (N_22440,N_17680,N_18157);
or U22441 (N_22441,N_16744,N_16484);
xor U22442 (N_22442,N_15745,N_16949);
xnor U22443 (N_22443,N_18143,N_15594);
and U22444 (N_22444,N_19244,N_19533);
nand U22445 (N_22445,N_15161,N_16568);
and U22446 (N_22446,N_15617,N_16567);
nor U22447 (N_22447,N_17398,N_16942);
or U22448 (N_22448,N_19280,N_16155);
xor U22449 (N_22449,N_19946,N_18798);
nor U22450 (N_22450,N_15963,N_18168);
and U22451 (N_22451,N_19323,N_16941);
nor U22452 (N_22452,N_19936,N_19793);
and U22453 (N_22453,N_19696,N_16728);
nand U22454 (N_22454,N_16474,N_15117);
or U22455 (N_22455,N_16509,N_17799);
xor U22456 (N_22456,N_18618,N_17008);
xnor U22457 (N_22457,N_19340,N_18062);
nand U22458 (N_22458,N_18898,N_17378);
nor U22459 (N_22459,N_15998,N_19385);
nor U22460 (N_22460,N_18693,N_17183);
nor U22461 (N_22461,N_15746,N_17048);
xor U22462 (N_22462,N_16512,N_19118);
xor U22463 (N_22463,N_19142,N_18520);
or U22464 (N_22464,N_17687,N_15936);
xnor U22465 (N_22465,N_18527,N_15865);
nand U22466 (N_22466,N_17099,N_16569);
nand U22467 (N_22467,N_15446,N_19843);
nand U22468 (N_22468,N_17937,N_18785);
nand U22469 (N_22469,N_16730,N_18023);
or U22470 (N_22470,N_16371,N_18049);
nor U22471 (N_22471,N_15475,N_15683);
and U22472 (N_22472,N_19209,N_19321);
or U22473 (N_22473,N_17290,N_18782);
xor U22474 (N_22474,N_19978,N_17911);
or U22475 (N_22475,N_19352,N_18050);
nand U22476 (N_22476,N_16869,N_19813);
xnor U22477 (N_22477,N_16670,N_16965);
nor U22478 (N_22478,N_18046,N_19232);
nand U22479 (N_22479,N_15540,N_16875);
nor U22480 (N_22480,N_16417,N_18883);
nand U22481 (N_22481,N_15400,N_17789);
or U22482 (N_22482,N_17710,N_18989);
or U22483 (N_22483,N_16885,N_17316);
nand U22484 (N_22484,N_19757,N_15796);
xnor U22485 (N_22485,N_16252,N_18897);
xor U22486 (N_22486,N_16543,N_15555);
nand U22487 (N_22487,N_18513,N_15306);
and U22488 (N_22488,N_18776,N_19148);
nor U22489 (N_22489,N_18108,N_15083);
and U22490 (N_22490,N_19282,N_19901);
nand U22491 (N_22491,N_15718,N_19042);
nand U22492 (N_22492,N_15602,N_19723);
nor U22493 (N_22493,N_17654,N_19791);
nand U22494 (N_22494,N_18584,N_15898);
nand U22495 (N_22495,N_17201,N_19411);
and U22496 (N_22496,N_16581,N_19218);
and U22497 (N_22497,N_18366,N_15701);
or U22498 (N_22498,N_17971,N_19054);
nand U22499 (N_22499,N_15739,N_15082);
or U22500 (N_22500,N_16900,N_19075);
xor U22501 (N_22501,N_18616,N_18251);
xnor U22502 (N_22502,N_16732,N_15469);
nand U22503 (N_22503,N_18362,N_19267);
and U22504 (N_22504,N_19410,N_17962);
nand U22505 (N_22505,N_18441,N_15252);
or U22506 (N_22506,N_19806,N_15169);
nand U22507 (N_22507,N_15023,N_16134);
nand U22508 (N_22508,N_15215,N_19376);
and U22509 (N_22509,N_19154,N_15137);
and U22510 (N_22510,N_19016,N_19035);
xor U22511 (N_22511,N_15322,N_17754);
and U22512 (N_22512,N_17435,N_16059);
and U22513 (N_22513,N_15162,N_19415);
or U22514 (N_22514,N_15876,N_19391);
and U22515 (N_22515,N_16221,N_16779);
or U22516 (N_22516,N_19710,N_18154);
nand U22517 (N_22517,N_19625,N_15295);
nand U22518 (N_22518,N_18673,N_18436);
xnor U22519 (N_22519,N_16696,N_15183);
and U22520 (N_22520,N_16802,N_15875);
and U22521 (N_22521,N_17779,N_17641);
xor U22522 (N_22522,N_16659,N_15792);
nand U22523 (N_22523,N_18722,N_15407);
and U22524 (N_22524,N_15272,N_15630);
or U22525 (N_22525,N_15981,N_16563);
nand U22526 (N_22526,N_17057,N_15105);
nand U22527 (N_22527,N_18040,N_19500);
nor U22528 (N_22528,N_19755,N_17264);
or U22529 (N_22529,N_18570,N_17470);
and U22530 (N_22530,N_15091,N_17887);
or U22531 (N_22531,N_16401,N_17596);
and U22532 (N_22532,N_16861,N_15251);
xnor U22533 (N_22533,N_17664,N_17830);
xnor U22534 (N_22534,N_15056,N_18246);
and U22535 (N_22535,N_15576,N_17803);
xor U22536 (N_22536,N_15697,N_15372);
xnor U22537 (N_22537,N_16627,N_19813);
nor U22538 (N_22538,N_17014,N_15991);
nor U22539 (N_22539,N_15766,N_18602);
xnor U22540 (N_22540,N_16065,N_19820);
and U22541 (N_22541,N_15516,N_19662);
xor U22542 (N_22542,N_17012,N_17472);
or U22543 (N_22543,N_17137,N_19548);
nor U22544 (N_22544,N_19593,N_18058);
nor U22545 (N_22545,N_18002,N_18438);
or U22546 (N_22546,N_16870,N_18979);
nand U22547 (N_22547,N_17437,N_17648);
nor U22548 (N_22548,N_16594,N_18975);
xor U22549 (N_22549,N_18255,N_17597);
nor U22550 (N_22550,N_17513,N_16914);
and U22551 (N_22551,N_17583,N_15289);
nor U22552 (N_22552,N_15552,N_19689);
nand U22553 (N_22553,N_16324,N_18182);
or U22554 (N_22554,N_19510,N_17972);
xor U22555 (N_22555,N_16500,N_16118);
or U22556 (N_22556,N_15406,N_15947);
or U22557 (N_22557,N_15998,N_17248);
or U22558 (N_22558,N_15442,N_18446);
nor U22559 (N_22559,N_17575,N_15339);
or U22560 (N_22560,N_17994,N_19974);
xor U22561 (N_22561,N_17256,N_16754);
and U22562 (N_22562,N_18184,N_17025);
nor U22563 (N_22563,N_16740,N_19586);
xnor U22564 (N_22564,N_17693,N_15026);
or U22565 (N_22565,N_16171,N_17605);
and U22566 (N_22566,N_17559,N_15910);
nand U22567 (N_22567,N_15779,N_18796);
or U22568 (N_22568,N_15274,N_15842);
and U22569 (N_22569,N_19926,N_18897);
nor U22570 (N_22570,N_19872,N_17757);
and U22571 (N_22571,N_18352,N_17679);
xor U22572 (N_22572,N_15180,N_19073);
or U22573 (N_22573,N_19977,N_19576);
xor U22574 (N_22574,N_16120,N_18161);
xnor U22575 (N_22575,N_18496,N_19320);
xnor U22576 (N_22576,N_16300,N_15537);
nor U22577 (N_22577,N_17164,N_18193);
nor U22578 (N_22578,N_18728,N_17087);
and U22579 (N_22579,N_19598,N_16901);
nor U22580 (N_22580,N_17597,N_16278);
xor U22581 (N_22581,N_18774,N_15674);
or U22582 (N_22582,N_15309,N_18080);
or U22583 (N_22583,N_15768,N_19040);
and U22584 (N_22584,N_19179,N_18254);
and U22585 (N_22585,N_19932,N_15863);
and U22586 (N_22586,N_17115,N_19306);
nand U22587 (N_22587,N_18931,N_18451);
nor U22588 (N_22588,N_17564,N_17554);
or U22589 (N_22589,N_17024,N_15684);
nand U22590 (N_22590,N_15459,N_16788);
and U22591 (N_22591,N_18978,N_16357);
or U22592 (N_22592,N_19696,N_19111);
nand U22593 (N_22593,N_17987,N_17513);
or U22594 (N_22594,N_18440,N_18384);
xor U22595 (N_22595,N_15525,N_19582);
nand U22596 (N_22596,N_19449,N_17787);
or U22597 (N_22597,N_17028,N_18669);
nor U22598 (N_22598,N_18472,N_16664);
xor U22599 (N_22599,N_16138,N_19328);
and U22600 (N_22600,N_17293,N_19435);
nor U22601 (N_22601,N_16262,N_19060);
nand U22602 (N_22602,N_16561,N_16482);
nor U22603 (N_22603,N_18205,N_16494);
and U22604 (N_22604,N_19669,N_15004);
or U22605 (N_22605,N_19241,N_15369);
and U22606 (N_22606,N_19008,N_19879);
or U22607 (N_22607,N_17644,N_17687);
nand U22608 (N_22608,N_18567,N_19099);
or U22609 (N_22609,N_18390,N_18744);
nand U22610 (N_22610,N_18473,N_19983);
nand U22611 (N_22611,N_17982,N_15512);
or U22612 (N_22612,N_17823,N_15382);
or U22613 (N_22613,N_19794,N_16224);
xor U22614 (N_22614,N_17310,N_18266);
nor U22615 (N_22615,N_15026,N_18577);
xnor U22616 (N_22616,N_18187,N_18991);
nor U22617 (N_22617,N_15727,N_19935);
and U22618 (N_22618,N_19674,N_19582);
and U22619 (N_22619,N_17549,N_18354);
xor U22620 (N_22620,N_18015,N_17452);
nor U22621 (N_22621,N_15488,N_17321);
nor U22622 (N_22622,N_17246,N_16190);
and U22623 (N_22623,N_17285,N_19106);
and U22624 (N_22624,N_18813,N_18580);
or U22625 (N_22625,N_19156,N_18324);
or U22626 (N_22626,N_16331,N_16618);
or U22627 (N_22627,N_19513,N_15616);
nand U22628 (N_22628,N_18498,N_19816);
nor U22629 (N_22629,N_15644,N_17149);
and U22630 (N_22630,N_19070,N_17264);
nand U22631 (N_22631,N_17404,N_19427);
nand U22632 (N_22632,N_19579,N_17943);
or U22633 (N_22633,N_15210,N_16594);
nand U22634 (N_22634,N_19498,N_15449);
nand U22635 (N_22635,N_17624,N_16938);
nand U22636 (N_22636,N_16121,N_18490);
or U22637 (N_22637,N_16785,N_18670);
xor U22638 (N_22638,N_16594,N_17635);
xor U22639 (N_22639,N_17130,N_19881);
nand U22640 (N_22640,N_16761,N_18442);
nor U22641 (N_22641,N_16028,N_19440);
xor U22642 (N_22642,N_17577,N_16029);
nor U22643 (N_22643,N_17870,N_18314);
and U22644 (N_22644,N_15373,N_16741);
or U22645 (N_22645,N_16784,N_17400);
nor U22646 (N_22646,N_16065,N_19758);
nor U22647 (N_22647,N_17767,N_17084);
or U22648 (N_22648,N_19934,N_16056);
nand U22649 (N_22649,N_15654,N_17666);
or U22650 (N_22650,N_18226,N_19550);
xor U22651 (N_22651,N_18814,N_19486);
nor U22652 (N_22652,N_18278,N_16809);
nor U22653 (N_22653,N_19201,N_16910);
xnor U22654 (N_22654,N_17911,N_16122);
xor U22655 (N_22655,N_15289,N_15964);
nand U22656 (N_22656,N_17189,N_15401);
or U22657 (N_22657,N_18314,N_15891);
and U22658 (N_22658,N_16832,N_15375);
or U22659 (N_22659,N_19360,N_19667);
or U22660 (N_22660,N_15294,N_16760);
xnor U22661 (N_22661,N_15629,N_16029);
xnor U22662 (N_22662,N_16497,N_19968);
or U22663 (N_22663,N_18674,N_15310);
nor U22664 (N_22664,N_19190,N_16841);
and U22665 (N_22665,N_16339,N_16962);
xor U22666 (N_22666,N_16323,N_18983);
xor U22667 (N_22667,N_16314,N_18774);
xor U22668 (N_22668,N_15260,N_15763);
nor U22669 (N_22669,N_16293,N_19025);
nor U22670 (N_22670,N_18648,N_15271);
nand U22671 (N_22671,N_18272,N_19003);
xor U22672 (N_22672,N_19735,N_18475);
and U22673 (N_22673,N_15583,N_17387);
nand U22674 (N_22674,N_16021,N_15527);
or U22675 (N_22675,N_16184,N_19465);
nand U22676 (N_22676,N_18985,N_18988);
and U22677 (N_22677,N_18986,N_16384);
nor U22678 (N_22678,N_19902,N_17170);
nor U22679 (N_22679,N_19140,N_18294);
or U22680 (N_22680,N_15724,N_19765);
nand U22681 (N_22681,N_19965,N_16325);
and U22682 (N_22682,N_18467,N_19625);
nor U22683 (N_22683,N_15881,N_16411);
and U22684 (N_22684,N_15373,N_17332);
and U22685 (N_22685,N_18510,N_15807);
or U22686 (N_22686,N_17292,N_19882);
or U22687 (N_22687,N_18263,N_19454);
xnor U22688 (N_22688,N_19534,N_17449);
xnor U22689 (N_22689,N_16023,N_15103);
and U22690 (N_22690,N_16531,N_18370);
and U22691 (N_22691,N_17648,N_19525);
nand U22692 (N_22692,N_15454,N_16866);
or U22693 (N_22693,N_15075,N_17507);
or U22694 (N_22694,N_16272,N_19460);
or U22695 (N_22695,N_18342,N_16562);
xnor U22696 (N_22696,N_18249,N_19004);
and U22697 (N_22697,N_17212,N_16459);
and U22698 (N_22698,N_18352,N_16488);
nand U22699 (N_22699,N_19865,N_16325);
and U22700 (N_22700,N_18928,N_18525);
or U22701 (N_22701,N_18265,N_19857);
xor U22702 (N_22702,N_19641,N_15183);
xnor U22703 (N_22703,N_15885,N_15227);
or U22704 (N_22704,N_15720,N_15342);
xnor U22705 (N_22705,N_16606,N_18110);
or U22706 (N_22706,N_19831,N_15359);
or U22707 (N_22707,N_15129,N_18084);
or U22708 (N_22708,N_17274,N_16930);
or U22709 (N_22709,N_15356,N_19650);
xnor U22710 (N_22710,N_16375,N_17951);
nor U22711 (N_22711,N_17148,N_17074);
nand U22712 (N_22712,N_18673,N_16231);
nor U22713 (N_22713,N_15187,N_16016);
or U22714 (N_22714,N_16953,N_15292);
xor U22715 (N_22715,N_19616,N_17617);
nor U22716 (N_22716,N_19258,N_17534);
nand U22717 (N_22717,N_16243,N_17891);
or U22718 (N_22718,N_15460,N_16534);
or U22719 (N_22719,N_15069,N_15245);
or U22720 (N_22720,N_18240,N_17213);
nor U22721 (N_22721,N_16767,N_19324);
and U22722 (N_22722,N_15253,N_18442);
xnor U22723 (N_22723,N_17116,N_19675);
or U22724 (N_22724,N_19108,N_19683);
xor U22725 (N_22725,N_17039,N_18256);
and U22726 (N_22726,N_18295,N_15549);
or U22727 (N_22727,N_16774,N_19176);
nor U22728 (N_22728,N_17329,N_17091);
xnor U22729 (N_22729,N_16254,N_19470);
or U22730 (N_22730,N_15541,N_17918);
or U22731 (N_22731,N_16848,N_15940);
nand U22732 (N_22732,N_16872,N_17729);
xnor U22733 (N_22733,N_16927,N_15905);
or U22734 (N_22734,N_17850,N_19780);
nand U22735 (N_22735,N_16078,N_16152);
xor U22736 (N_22736,N_18100,N_15972);
xnor U22737 (N_22737,N_15716,N_19553);
nand U22738 (N_22738,N_17213,N_19720);
xnor U22739 (N_22739,N_17373,N_18257);
nand U22740 (N_22740,N_16687,N_15795);
or U22741 (N_22741,N_18980,N_17576);
nand U22742 (N_22742,N_17370,N_19670);
or U22743 (N_22743,N_17017,N_16686);
and U22744 (N_22744,N_15758,N_16553);
and U22745 (N_22745,N_18664,N_19186);
nand U22746 (N_22746,N_18825,N_16091);
and U22747 (N_22747,N_15706,N_16027);
xor U22748 (N_22748,N_19280,N_15550);
nand U22749 (N_22749,N_18632,N_19792);
and U22750 (N_22750,N_19082,N_17061);
and U22751 (N_22751,N_17611,N_16300);
nand U22752 (N_22752,N_18930,N_18090);
nor U22753 (N_22753,N_16462,N_16093);
and U22754 (N_22754,N_16542,N_18098);
xnor U22755 (N_22755,N_16243,N_16889);
or U22756 (N_22756,N_15780,N_16513);
or U22757 (N_22757,N_15675,N_19567);
and U22758 (N_22758,N_15490,N_19960);
nand U22759 (N_22759,N_15050,N_18374);
or U22760 (N_22760,N_17203,N_16943);
nor U22761 (N_22761,N_17772,N_19344);
or U22762 (N_22762,N_15446,N_19608);
or U22763 (N_22763,N_18347,N_15877);
or U22764 (N_22764,N_16426,N_17667);
or U22765 (N_22765,N_17827,N_19204);
or U22766 (N_22766,N_17797,N_18018);
nor U22767 (N_22767,N_15634,N_19423);
nor U22768 (N_22768,N_18203,N_16184);
nor U22769 (N_22769,N_15695,N_19056);
nand U22770 (N_22770,N_15581,N_16893);
nand U22771 (N_22771,N_16493,N_15756);
xor U22772 (N_22772,N_16193,N_18355);
nor U22773 (N_22773,N_15035,N_18494);
xnor U22774 (N_22774,N_18676,N_19756);
xor U22775 (N_22775,N_18389,N_15231);
nand U22776 (N_22776,N_15386,N_17298);
or U22777 (N_22777,N_18310,N_19080);
or U22778 (N_22778,N_18306,N_18420);
and U22779 (N_22779,N_15366,N_15516);
nor U22780 (N_22780,N_18952,N_18293);
nand U22781 (N_22781,N_17160,N_17601);
nand U22782 (N_22782,N_16642,N_19593);
nand U22783 (N_22783,N_19611,N_15485);
nor U22784 (N_22784,N_17442,N_18425);
and U22785 (N_22785,N_15590,N_19126);
and U22786 (N_22786,N_17026,N_17686);
and U22787 (N_22787,N_17333,N_16106);
or U22788 (N_22788,N_19867,N_15053);
nand U22789 (N_22789,N_18723,N_18829);
nand U22790 (N_22790,N_18306,N_19763);
or U22791 (N_22791,N_19794,N_18902);
nor U22792 (N_22792,N_17502,N_16360);
and U22793 (N_22793,N_17265,N_17453);
or U22794 (N_22794,N_18910,N_19733);
or U22795 (N_22795,N_15297,N_19001);
xor U22796 (N_22796,N_16630,N_16289);
nand U22797 (N_22797,N_16479,N_17601);
nor U22798 (N_22798,N_17665,N_18181);
nor U22799 (N_22799,N_15020,N_18936);
or U22800 (N_22800,N_16126,N_16568);
nor U22801 (N_22801,N_16351,N_17886);
or U22802 (N_22802,N_16691,N_17595);
and U22803 (N_22803,N_17989,N_17223);
or U22804 (N_22804,N_15681,N_15682);
xnor U22805 (N_22805,N_19875,N_17512);
xnor U22806 (N_22806,N_17009,N_17957);
xnor U22807 (N_22807,N_15429,N_19392);
nor U22808 (N_22808,N_16200,N_19139);
or U22809 (N_22809,N_19859,N_17082);
or U22810 (N_22810,N_16195,N_16102);
nand U22811 (N_22811,N_17628,N_18247);
or U22812 (N_22812,N_16253,N_19144);
or U22813 (N_22813,N_16901,N_19018);
xnor U22814 (N_22814,N_15143,N_16222);
or U22815 (N_22815,N_17512,N_18482);
nor U22816 (N_22816,N_18232,N_16157);
xor U22817 (N_22817,N_15169,N_15768);
or U22818 (N_22818,N_15357,N_16192);
or U22819 (N_22819,N_18807,N_17816);
xnor U22820 (N_22820,N_17725,N_19667);
or U22821 (N_22821,N_15117,N_16717);
nor U22822 (N_22822,N_17443,N_15122);
nor U22823 (N_22823,N_16418,N_16140);
nor U22824 (N_22824,N_18666,N_18034);
nor U22825 (N_22825,N_17650,N_15611);
or U22826 (N_22826,N_15609,N_15097);
nand U22827 (N_22827,N_17298,N_15166);
xnor U22828 (N_22828,N_17399,N_19574);
or U22829 (N_22829,N_16901,N_19103);
nand U22830 (N_22830,N_18392,N_15080);
or U22831 (N_22831,N_18101,N_16576);
xor U22832 (N_22832,N_19706,N_16641);
nor U22833 (N_22833,N_18650,N_18876);
and U22834 (N_22834,N_15275,N_16331);
xor U22835 (N_22835,N_19985,N_15613);
nor U22836 (N_22836,N_17325,N_17491);
xor U22837 (N_22837,N_19721,N_19615);
xnor U22838 (N_22838,N_19105,N_16649);
or U22839 (N_22839,N_16086,N_19368);
and U22840 (N_22840,N_17212,N_18114);
xor U22841 (N_22841,N_16250,N_19585);
and U22842 (N_22842,N_19428,N_15163);
or U22843 (N_22843,N_18805,N_16433);
nor U22844 (N_22844,N_17905,N_17781);
nor U22845 (N_22845,N_15324,N_18319);
xnor U22846 (N_22846,N_18137,N_15788);
and U22847 (N_22847,N_15095,N_19275);
nand U22848 (N_22848,N_16838,N_16099);
xnor U22849 (N_22849,N_15935,N_17832);
xnor U22850 (N_22850,N_15200,N_15401);
xor U22851 (N_22851,N_17555,N_17356);
nor U22852 (N_22852,N_16826,N_16385);
nand U22853 (N_22853,N_19907,N_19281);
xor U22854 (N_22854,N_18483,N_16990);
and U22855 (N_22855,N_17670,N_19362);
and U22856 (N_22856,N_19540,N_18766);
or U22857 (N_22857,N_19615,N_18933);
xor U22858 (N_22858,N_16325,N_17284);
nor U22859 (N_22859,N_15084,N_18865);
and U22860 (N_22860,N_15499,N_19760);
and U22861 (N_22861,N_15079,N_17745);
and U22862 (N_22862,N_15729,N_15747);
and U22863 (N_22863,N_16902,N_15672);
nor U22864 (N_22864,N_16745,N_15615);
and U22865 (N_22865,N_18474,N_15775);
and U22866 (N_22866,N_15570,N_19345);
nand U22867 (N_22867,N_18942,N_15793);
nand U22868 (N_22868,N_16077,N_19053);
or U22869 (N_22869,N_19382,N_16504);
nor U22870 (N_22870,N_15270,N_15394);
or U22871 (N_22871,N_15040,N_19407);
nand U22872 (N_22872,N_15661,N_15351);
nand U22873 (N_22873,N_17969,N_16193);
nor U22874 (N_22874,N_19648,N_17205);
and U22875 (N_22875,N_17317,N_16269);
and U22876 (N_22876,N_17343,N_16514);
xnor U22877 (N_22877,N_18907,N_19174);
and U22878 (N_22878,N_16803,N_19928);
or U22879 (N_22879,N_17496,N_18537);
or U22880 (N_22880,N_19665,N_18694);
nor U22881 (N_22881,N_18180,N_16060);
nand U22882 (N_22882,N_18041,N_18139);
xor U22883 (N_22883,N_16560,N_16933);
and U22884 (N_22884,N_18767,N_16296);
nand U22885 (N_22885,N_19469,N_19101);
xnor U22886 (N_22886,N_18973,N_17519);
or U22887 (N_22887,N_16390,N_18870);
xnor U22888 (N_22888,N_17933,N_15414);
nor U22889 (N_22889,N_18983,N_18391);
and U22890 (N_22890,N_16398,N_17092);
nor U22891 (N_22891,N_15862,N_18089);
and U22892 (N_22892,N_15498,N_16387);
or U22893 (N_22893,N_16134,N_17569);
nor U22894 (N_22894,N_16710,N_15011);
nor U22895 (N_22895,N_17155,N_15094);
or U22896 (N_22896,N_18477,N_18930);
or U22897 (N_22897,N_15844,N_19630);
and U22898 (N_22898,N_17961,N_19521);
nand U22899 (N_22899,N_17597,N_18195);
xnor U22900 (N_22900,N_19451,N_19151);
or U22901 (N_22901,N_19715,N_17390);
xnor U22902 (N_22902,N_17804,N_18364);
nand U22903 (N_22903,N_18045,N_16777);
nor U22904 (N_22904,N_15051,N_15576);
nor U22905 (N_22905,N_16317,N_18151);
xnor U22906 (N_22906,N_16390,N_18190);
and U22907 (N_22907,N_15390,N_16943);
xnor U22908 (N_22908,N_19035,N_15202);
and U22909 (N_22909,N_16634,N_17389);
and U22910 (N_22910,N_19512,N_15272);
nor U22911 (N_22911,N_16901,N_18976);
nand U22912 (N_22912,N_18210,N_19805);
and U22913 (N_22913,N_16283,N_15927);
and U22914 (N_22914,N_17551,N_19269);
xor U22915 (N_22915,N_19177,N_15151);
nor U22916 (N_22916,N_15097,N_18763);
and U22917 (N_22917,N_16402,N_19066);
nand U22918 (N_22918,N_16203,N_18423);
nor U22919 (N_22919,N_15347,N_18993);
and U22920 (N_22920,N_17407,N_18601);
nor U22921 (N_22921,N_18637,N_16276);
nor U22922 (N_22922,N_17066,N_17846);
nor U22923 (N_22923,N_18447,N_16341);
nand U22924 (N_22924,N_16406,N_19016);
or U22925 (N_22925,N_16626,N_18010);
nor U22926 (N_22926,N_16963,N_16154);
nand U22927 (N_22927,N_17636,N_16915);
and U22928 (N_22928,N_19378,N_18097);
nor U22929 (N_22929,N_15354,N_15870);
nand U22930 (N_22930,N_15645,N_18917);
nor U22931 (N_22931,N_18476,N_18465);
xnor U22932 (N_22932,N_15349,N_19431);
and U22933 (N_22933,N_17444,N_17231);
nand U22934 (N_22934,N_19292,N_18674);
and U22935 (N_22935,N_18675,N_16269);
nand U22936 (N_22936,N_16315,N_17850);
xor U22937 (N_22937,N_18473,N_18684);
xor U22938 (N_22938,N_17048,N_19038);
or U22939 (N_22939,N_18049,N_16096);
xor U22940 (N_22940,N_17598,N_19152);
and U22941 (N_22941,N_17083,N_17664);
nor U22942 (N_22942,N_16391,N_16677);
nand U22943 (N_22943,N_17681,N_19819);
nand U22944 (N_22944,N_18200,N_19193);
nand U22945 (N_22945,N_17611,N_19472);
or U22946 (N_22946,N_17596,N_18371);
xnor U22947 (N_22947,N_18032,N_15638);
and U22948 (N_22948,N_15223,N_19745);
xor U22949 (N_22949,N_16684,N_15336);
and U22950 (N_22950,N_17928,N_15232);
and U22951 (N_22951,N_17992,N_18488);
or U22952 (N_22952,N_18215,N_17773);
xnor U22953 (N_22953,N_18724,N_15895);
and U22954 (N_22954,N_18032,N_16064);
nor U22955 (N_22955,N_16965,N_19235);
nor U22956 (N_22956,N_16042,N_16621);
xnor U22957 (N_22957,N_19758,N_16139);
or U22958 (N_22958,N_18703,N_16087);
or U22959 (N_22959,N_15735,N_15622);
nor U22960 (N_22960,N_16326,N_16479);
and U22961 (N_22961,N_17789,N_15396);
xnor U22962 (N_22962,N_16749,N_18002);
or U22963 (N_22963,N_18792,N_19420);
or U22964 (N_22964,N_15024,N_16247);
xnor U22965 (N_22965,N_19473,N_19799);
xnor U22966 (N_22966,N_17782,N_17605);
nor U22967 (N_22967,N_19901,N_17026);
and U22968 (N_22968,N_16967,N_18737);
nor U22969 (N_22969,N_19199,N_19977);
nand U22970 (N_22970,N_18005,N_15803);
xnor U22971 (N_22971,N_16601,N_18818);
and U22972 (N_22972,N_16462,N_16148);
nor U22973 (N_22973,N_16869,N_16285);
and U22974 (N_22974,N_18415,N_17560);
nand U22975 (N_22975,N_17827,N_16368);
nand U22976 (N_22976,N_15183,N_18648);
xor U22977 (N_22977,N_17321,N_19150);
nor U22978 (N_22978,N_19379,N_16353);
nor U22979 (N_22979,N_19652,N_18610);
or U22980 (N_22980,N_16496,N_16807);
xnor U22981 (N_22981,N_19972,N_16323);
xor U22982 (N_22982,N_17926,N_19220);
nor U22983 (N_22983,N_15135,N_15868);
xnor U22984 (N_22984,N_19054,N_18302);
xor U22985 (N_22985,N_18237,N_18137);
and U22986 (N_22986,N_15682,N_15277);
or U22987 (N_22987,N_16547,N_15686);
xnor U22988 (N_22988,N_17349,N_15791);
nand U22989 (N_22989,N_18060,N_18733);
or U22990 (N_22990,N_19345,N_18135);
and U22991 (N_22991,N_16033,N_16883);
nand U22992 (N_22992,N_16043,N_17478);
xor U22993 (N_22993,N_19618,N_16764);
or U22994 (N_22994,N_15242,N_15124);
nor U22995 (N_22995,N_17759,N_15194);
nor U22996 (N_22996,N_19865,N_18295);
and U22997 (N_22997,N_18354,N_15232);
or U22998 (N_22998,N_18340,N_16190);
nand U22999 (N_22999,N_16522,N_16543);
or U23000 (N_23000,N_15748,N_15691);
and U23001 (N_23001,N_19096,N_19226);
or U23002 (N_23002,N_15881,N_15974);
and U23003 (N_23003,N_18492,N_15183);
xor U23004 (N_23004,N_15161,N_17174);
or U23005 (N_23005,N_17769,N_19819);
xor U23006 (N_23006,N_17684,N_17347);
xnor U23007 (N_23007,N_18481,N_15296);
nor U23008 (N_23008,N_16263,N_18156);
xor U23009 (N_23009,N_18585,N_16489);
nand U23010 (N_23010,N_18702,N_15971);
nand U23011 (N_23011,N_18241,N_19404);
nand U23012 (N_23012,N_19161,N_18528);
xor U23013 (N_23013,N_16707,N_17631);
xnor U23014 (N_23014,N_18602,N_19058);
or U23015 (N_23015,N_17132,N_17694);
xor U23016 (N_23016,N_18718,N_16322);
nand U23017 (N_23017,N_16681,N_16810);
and U23018 (N_23018,N_16860,N_18853);
nor U23019 (N_23019,N_19190,N_19474);
xnor U23020 (N_23020,N_18897,N_16584);
and U23021 (N_23021,N_18714,N_17006);
nor U23022 (N_23022,N_19287,N_19243);
nor U23023 (N_23023,N_17926,N_17072);
nor U23024 (N_23024,N_18811,N_19296);
and U23025 (N_23025,N_18242,N_19542);
and U23026 (N_23026,N_18986,N_16147);
xnor U23027 (N_23027,N_18551,N_17666);
and U23028 (N_23028,N_19077,N_19994);
or U23029 (N_23029,N_15643,N_17009);
xor U23030 (N_23030,N_16004,N_16789);
or U23031 (N_23031,N_18314,N_17417);
nor U23032 (N_23032,N_19159,N_18638);
and U23033 (N_23033,N_15476,N_18015);
nand U23034 (N_23034,N_16627,N_18881);
xor U23035 (N_23035,N_16732,N_19996);
xnor U23036 (N_23036,N_17680,N_19731);
nor U23037 (N_23037,N_17474,N_18692);
and U23038 (N_23038,N_15153,N_17735);
nor U23039 (N_23039,N_15160,N_17155);
or U23040 (N_23040,N_15784,N_16491);
or U23041 (N_23041,N_15451,N_16491);
xnor U23042 (N_23042,N_16901,N_17489);
xor U23043 (N_23043,N_17232,N_16088);
nor U23044 (N_23044,N_16989,N_16229);
nand U23045 (N_23045,N_15003,N_16797);
nor U23046 (N_23046,N_19041,N_16324);
and U23047 (N_23047,N_16059,N_18925);
nor U23048 (N_23048,N_17554,N_19908);
nand U23049 (N_23049,N_18374,N_16550);
nand U23050 (N_23050,N_17294,N_17953);
and U23051 (N_23051,N_17176,N_18426);
nor U23052 (N_23052,N_18814,N_17045);
nand U23053 (N_23053,N_15950,N_18842);
or U23054 (N_23054,N_15286,N_15677);
and U23055 (N_23055,N_19696,N_19059);
or U23056 (N_23056,N_16178,N_15409);
nand U23057 (N_23057,N_19394,N_15227);
or U23058 (N_23058,N_18508,N_19577);
or U23059 (N_23059,N_15293,N_17138);
and U23060 (N_23060,N_15138,N_18592);
or U23061 (N_23061,N_17320,N_16039);
nor U23062 (N_23062,N_16063,N_16858);
or U23063 (N_23063,N_15836,N_18788);
or U23064 (N_23064,N_19266,N_16519);
xor U23065 (N_23065,N_19857,N_15933);
nor U23066 (N_23066,N_15111,N_19084);
nor U23067 (N_23067,N_18830,N_18402);
xor U23068 (N_23068,N_16252,N_15533);
xnor U23069 (N_23069,N_16827,N_19387);
and U23070 (N_23070,N_16243,N_18835);
and U23071 (N_23071,N_19488,N_17019);
nor U23072 (N_23072,N_15718,N_16645);
nand U23073 (N_23073,N_18135,N_18613);
nor U23074 (N_23074,N_16782,N_18068);
and U23075 (N_23075,N_18171,N_16833);
nor U23076 (N_23076,N_15284,N_19884);
and U23077 (N_23077,N_19471,N_18639);
xnor U23078 (N_23078,N_17713,N_17508);
nand U23079 (N_23079,N_17426,N_15804);
xor U23080 (N_23080,N_16898,N_16011);
nor U23081 (N_23081,N_15087,N_19840);
or U23082 (N_23082,N_18682,N_15783);
xnor U23083 (N_23083,N_16911,N_18819);
and U23084 (N_23084,N_17009,N_18205);
and U23085 (N_23085,N_19777,N_18985);
nor U23086 (N_23086,N_17116,N_15592);
nor U23087 (N_23087,N_18846,N_19256);
nand U23088 (N_23088,N_16600,N_16101);
nor U23089 (N_23089,N_17397,N_16809);
and U23090 (N_23090,N_19238,N_17686);
or U23091 (N_23091,N_17316,N_15374);
and U23092 (N_23092,N_19121,N_18210);
xnor U23093 (N_23093,N_16482,N_15894);
xor U23094 (N_23094,N_16138,N_17601);
and U23095 (N_23095,N_19062,N_18659);
nor U23096 (N_23096,N_15139,N_17545);
nand U23097 (N_23097,N_16905,N_18318);
or U23098 (N_23098,N_15476,N_17061);
or U23099 (N_23099,N_15366,N_17083);
and U23100 (N_23100,N_18260,N_19966);
and U23101 (N_23101,N_16516,N_19286);
nand U23102 (N_23102,N_15603,N_18341);
nor U23103 (N_23103,N_16718,N_17139);
and U23104 (N_23104,N_19668,N_15075);
nor U23105 (N_23105,N_15260,N_19858);
and U23106 (N_23106,N_19236,N_15931);
and U23107 (N_23107,N_19225,N_19418);
xor U23108 (N_23108,N_17298,N_19639);
and U23109 (N_23109,N_19272,N_18533);
or U23110 (N_23110,N_16781,N_19536);
nor U23111 (N_23111,N_18168,N_17768);
nand U23112 (N_23112,N_18181,N_18615);
nand U23113 (N_23113,N_19862,N_18149);
nor U23114 (N_23114,N_15717,N_16827);
and U23115 (N_23115,N_18552,N_17917);
xor U23116 (N_23116,N_19232,N_17983);
nor U23117 (N_23117,N_19332,N_19036);
and U23118 (N_23118,N_17585,N_17202);
or U23119 (N_23119,N_19704,N_18164);
nor U23120 (N_23120,N_18196,N_18110);
and U23121 (N_23121,N_16853,N_15992);
nor U23122 (N_23122,N_18819,N_18133);
or U23123 (N_23123,N_17419,N_19551);
and U23124 (N_23124,N_19324,N_18965);
and U23125 (N_23125,N_16679,N_16533);
xnor U23126 (N_23126,N_19748,N_18480);
xnor U23127 (N_23127,N_19621,N_17851);
or U23128 (N_23128,N_15727,N_18248);
and U23129 (N_23129,N_16906,N_18385);
nand U23130 (N_23130,N_19365,N_18286);
xnor U23131 (N_23131,N_17410,N_17768);
and U23132 (N_23132,N_15671,N_18832);
or U23133 (N_23133,N_15613,N_16605);
or U23134 (N_23134,N_16540,N_16171);
and U23135 (N_23135,N_19463,N_15399);
or U23136 (N_23136,N_16192,N_19890);
nand U23137 (N_23137,N_16539,N_16852);
xnor U23138 (N_23138,N_17773,N_17805);
xnor U23139 (N_23139,N_17851,N_15409);
or U23140 (N_23140,N_19228,N_19834);
and U23141 (N_23141,N_19550,N_19360);
and U23142 (N_23142,N_15568,N_18842);
nor U23143 (N_23143,N_19509,N_16236);
xor U23144 (N_23144,N_17263,N_15709);
or U23145 (N_23145,N_15038,N_18342);
or U23146 (N_23146,N_17602,N_15158);
or U23147 (N_23147,N_18749,N_19363);
or U23148 (N_23148,N_15432,N_19716);
nor U23149 (N_23149,N_18074,N_19908);
nand U23150 (N_23150,N_15608,N_16103);
or U23151 (N_23151,N_18847,N_19620);
and U23152 (N_23152,N_17569,N_16892);
or U23153 (N_23153,N_17152,N_19194);
and U23154 (N_23154,N_17605,N_19727);
and U23155 (N_23155,N_17484,N_17904);
nor U23156 (N_23156,N_18422,N_16729);
nand U23157 (N_23157,N_19987,N_16655);
or U23158 (N_23158,N_18470,N_16784);
xor U23159 (N_23159,N_18853,N_19346);
or U23160 (N_23160,N_15895,N_18003);
xor U23161 (N_23161,N_17244,N_18757);
and U23162 (N_23162,N_16368,N_17480);
xor U23163 (N_23163,N_16442,N_15323);
nor U23164 (N_23164,N_16436,N_17093);
nand U23165 (N_23165,N_17640,N_17692);
xor U23166 (N_23166,N_15798,N_17433);
nand U23167 (N_23167,N_16210,N_18424);
nand U23168 (N_23168,N_15496,N_16503);
nor U23169 (N_23169,N_17420,N_19175);
and U23170 (N_23170,N_15864,N_16308);
nor U23171 (N_23171,N_15713,N_19328);
or U23172 (N_23172,N_15086,N_18711);
nor U23173 (N_23173,N_17202,N_16042);
xor U23174 (N_23174,N_16238,N_16085);
and U23175 (N_23175,N_17292,N_18282);
or U23176 (N_23176,N_19341,N_15569);
and U23177 (N_23177,N_17679,N_16877);
xor U23178 (N_23178,N_17197,N_18057);
nand U23179 (N_23179,N_19421,N_16855);
or U23180 (N_23180,N_18224,N_19545);
xor U23181 (N_23181,N_19257,N_18313);
nand U23182 (N_23182,N_19285,N_17264);
nand U23183 (N_23183,N_15970,N_18705);
xor U23184 (N_23184,N_19028,N_15906);
xor U23185 (N_23185,N_17193,N_16123);
nand U23186 (N_23186,N_15448,N_16400);
nand U23187 (N_23187,N_18055,N_17442);
nor U23188 (N_23188,N_18848,N_15893);
or U23189 (N_23189,N_17184,N_16871);
xor U23190 (N_23190,N_19442,N_16612);
nand U23191 (N_23191,N_18067,N_16174);
and U23192 (N_23192,N_17976,N_19344);
and U23193 (N_23193,N_16328,N_17467);
nand U23194 (N_23194,N_16918,N_19403);
or U23195 (N_23195,N_16875,N_15968);
or U23196 (N_23196,N_19004,N_15324);
nor U23197 (N_23197,N_15400,N_17557);
nand U23198 (N_23198,N_16437,N_15601);
nor U23199 (N_23199,N_15952,N_18028);
nor U23200 (N_23200,N_15694,N_16618);
nor U23201 (N_23201,N_15946,N_18524);
or U23202 (N_23202,N_15684,N_18786);
and U23203 (N_23203,N_16008,N_17038);
nor U23204 (N_23204,N_19833,N_17799);
xnor U23205 (N_23205,N_19091,N_18269);
and U23206 (N_23206,N_19782,N_16227);
or U23207 (N_23207,N_15603,N_19306);
nand U23208 (N_23208,N_17412,N_17268);
xor U23209 (N_23209,N_15487,N_18322);
and U23210 (N_23210,N_18880,N_18779);
or U23211 (N_23211,N_19237,N_18602);
or U23212 (N_23212,N_15717,N_17006);
xor U23213 (N_23213,N_19243,N_19668);
nand U23214 (N_23214,N_19603,N_15406);
nand U23215 (N_23215,N_17959,N_18684);
nor U23216 (N_23216,N_16275,N_19223);
or U23217 (N_23217,N_17387,N_16765);
xor U23218 (N_23218,N_16461,N_17192);
xnor U23219 (N_23219,N_16942,N_16535);
xnor U23220 (N_23220,N_15272,N_17472);
xor U23221 (N_23221,N_17922,N_15356);
nand U23222 (N_23222,N_18217,N_17693);
and U23223 (N_23223,N_18332,N_15939);
nand U23224 (N_23224,N_19591,N_18544);
or U23225 (N_23225,N_17777,N_18316);
nand U23226 (N_23226,N_15054,N_18064);
or U23227 (N_23227,N_16801,N_16325);
nand U23228 (N_23228,N_15814,N_19881);
xnor U23229 (N_23229,N_18384,N_19108);
or U23230 (N_23230,N_19176,N_15272);
or U23231 (N_23231,N_15756,N_16106);
xnor U23232 (N_23232,N_17263,N_17447);
and U23233 (N_23233,N_16649,N_15220);
or U23234 (N_23234,N_16989,N_15834);
nor U23235 (N_23235,N_18238,N_16815);
nor U23236 (N_23236,N_18517,N_16272);
and U23237 (N_23237,N_17848,N_19817);
xor U23238 (N_23238,N_15165,N_15348);
nand U23239 (N_23239,N_16740,N_18710);
or U23240 (N_23240,N_19578,N_17300);
nor U23241 (N_23241,N_18764,N_16355);
xnor U23242 (N_23242,N_16336,N_15417);
and U23243 (N_23243,N_19990,N_17691);
or U23244 (N_23244,N_17748,N_15373);
nor U23245 (N_23245,N_18651,N_15959);
nand U23246 (N_23246,N_17913,N_19276);
and U23247 (N_23247,N_18063,N_19707);
nor U23248 (N_23248,N_15848,N_15766);
and U23249 (N_23249,N_17142,N_15211);
xnor U23250 (N_23250,N_15418,N_16584);
xnor U23251 (N_23251,N_16148,N_18139);
nor U23252 (N_23252,N_15114,N_17507);
nand U23253 (N_23253,N_18738,N_19454);
nor U23254 (N_23254,N_18440,N_17390);
nor U23255 (N_23255,N_16961,N_19120);
xor U23256 (N_23256,N_18103,N_17451);
nor U23257 (N_23257,N_17293,N_18592);
xor U23258 (N_23258,N_18712,N_19649);
or U23259 (N_23259,N_16001,N_18577);
xnor U23260 (N_23260,N_19184,N_16449);
xnor U23261 (N_23261,N_19370,N_18908);
nand U23262 (N_23262,N_18233,N_17380);
xor U23263 (N_23263,N_18183,N_16828);
or U23264 (N_23264,N_19408,N_16971);
xnor U23265 (N_23265,N_15770,N_15159);
or U23266 (N_23266,N_15894,N_19647);
or U23267 (N_23267,N_16394,N_19668);
and U23268 (N_23268,N_17365,N_18982);
nand U23269 (N_23269,N_18205,N_17897);
nand U23270 (N_23270,N_17942,N_19935);
and U23271 (N_23271,N_18029,N_16735);
nand U23272 (N_23272,N_15397,N_17961);
xor U23273 (N_23273,N_17710,N_16847);
nand U23274 (N_23274,N_17027,N_15735);
and U23275 (N_23275,N_15801,N_19510);
xnor U23276 (N_23276,N_17426,N_17158);
and U23277 (N_23277,N_17032,N_19583);
nor U23278 (N_23278,N_19938,N_15130);
nor U23279 (N_23279,N_17156,N_18118);
and U23280 (N_23280,N_17166,N_15976);
xnor U23281 (N_23281,N_17516,N_18446);
xor U23282 (N_23282,N_17001,N_15280);
xor U23283 (N_23283,N_18339,N_17154);
or U23284 (N_23284,N_17907,N_17702);
nor U23285 (N_23285,N_15115,N_19523);
nor U23286 (N_23286,N_17027,N_15461);
xor U23287 (N_23287,N_15999,N_17759);
xor U23288 (N_23288,N_17854,N_17277);
xor U23289 (N_23289,N_17245,N_15346);
xnor U23290 (N_23290,N_16998,N_17134);
or U23291 (N_23291,N_17606,N_17212);
nor U23292 (N_23292,N_18532,N_19420);
or U23293 (N_23293,N_17003,N_16879);
nand U23294 (N_23294,N_15487,N_17187);
nand U23295 (N_23295,N_15858,N_17191);
xor U23296 (N_23296,N_16914,N_17188);
nand U23297 (N_23297,N_19651,N_16326);
and U23298 (N_23298,N_15072,N_18074);
xnor U23299 (N_23299,N_18465,N_15816);
xnor U23300 (N_23300,N_18063,N_15943);
or U23301 (N_23301,N_17845,N_19674);
nor U23302 (N_23302,N_16448,N_16406);
nor U23303 (N_23303,N_16307,N_16773);
and U23304 (N_23304,N_19881,N_15137);
xor U23305 (N_23305,N_18321,N_17573);
xnor U23306 (N_23306,N_17824,N_16082);
or U23307 (N_23307,N_19586,N_16936);
or U23308 (N_23308,N_15455,N_19543);
nand U23309 (N_23309,N_17681,N_15817);
and U23310 (N_23310,N_18655,N_18773);
or U23311 (N_23311,N_16675,N_15646);
nand U23312 (N_23312,N_15049,N_16296);
xnor U23313 (N_23313,N_19956,N_19927);
nand U23314 (N_23314,N_16623,N_16260);
xnor U23315 (N_23315,N_16886,N_18528);
nand U23316 (N_23316,N_19547,N_19796);
or U23317 (N_23317,N_18803,N_16895);
nand U23318 (N_23318,N_16940,N_19550);
or U23319 (N_23319,N_17818,N_19943);
xor U23320 (N_23320,N_16039,N_19017);
nand U23321 (N_23321,N_17888,N_15937);
nor U23322 (N_23322,N_19281,N_17645);
or U23323 (N_23323,N_19959,N_16982);
xor U23324 (N_23324,N_16806,N_18489);
nor U23325 (N_23325,N_15718,N_15231);
xor U23326 (N_23326,N_15544,N_15091);
nand U23327 (N_23327,N_17483,N_16753);
or U23328 (N_23328,N_18042,N_17305);
and U23329 (N_23329,N_15877,N_17443);
nand U23330 (N_23330,N_18180,N_18514);
nand U23331 (N_23331,N_17898,N_15924);
and U23332 (N_23332,N_18437,N_18371);
nor U23333 (N_23333,N_15160,N_15473);
xnor U23334 (N_23334,N_15987,N_17377);
nor U23335 (N_23335,N_18994,N_16698);
or U23336 (N_23336,N_18527,N_19055);
nand U23337 (N_23337,N_18530,N_16862);
or U23338 (N_23338,N_19679,N_18487);
xor U23339 (N_23339,N_18865,N_15081);
nand U23340 (N_23340,N_17879,N_15356);
or U23341 (N_23341,N_19669,N_15212);
xnor U23342 (N_23342,N_15628,N_15873);
nand U23343 (N_23343,N_15332,N_15709);
nor U23344 (N_23344,N_16265,N_18047);
nor U23345 (N_23345,N_16276,N_18608);
and U23346 (N_23346,N_17874,N_17892);
and U23347 (N_23347,N_19360,N_17659);
nor U23348 (N_23348,N_19740,N_16579);
and U23349 (N_23349,N_19608,N_17370);
nand U23350 (N_23350,N_15519,N_15370);
xor U23351 (N_23351,N_19391,N_19848);
and U23352 (N_23352,N_15750,N_18572);
nand U23353 (N_23353,N_17876,N_16682);
nor U23354 (N_23354,N_16354,N_16938);
and U23355 (N_23355,N_17014,N_17824);
nor U23356 (N_23356,N_18670,N_15021);
xnor U23357 (N_23357,N_17594,N_19822);
and U23358 (N_23358,N_15905,N_17141);
or U23359 (N_23359,N_17748,N_15307);
or U23360 (N_23360,N_17316,N_16020);
or U23361 (N_23361,N_19933,N_15608);
and U23362 (N_23362,N_18197,N_16523);
or U23363 (N_23363,N_16059,N_17868);
nor U23364 (N_23364,N_15542,N_19174);
nand U23365 (N_23365,N_17054,N_19551);
or U23366 (N_23366,N_15637,N_19729);
nand U23367 (N_23367,N_19763,N_19643);
nor U23368 (N_23368,N_19149,N_15571);
nor U23369 (N_23369,N_19045,N_15754);
and U23370 (N_23370,N_16769,N_18612);
and U23371 (N_23371,N_16120,N_18240);
nor U23372 (N_23372,N_18863,N_17444);
and U23373 (N_23373,N_17068,N_16604);
nand U23374 (N_23374,N_17593,N_17075);
nor U23375 (N_23375,N_16363,N_19685);
nor U23376 (N_23376,N_17768,N_17788);
and U23377 (N_23377,N_18609,N_17776);
nand U23378 (N_23378,N_18816,N_15203);
or U23379 (N_23379,N_19153,N_18621);
xnor U23380 (N_23380,N_19611,N_19329);
xor U23381 (N_23381,N_19688,N_17108);
and U23382 (N_23382,N_19803,N_17629);
nor U23383 (N_23383,N_16550,N_15496);
and U23384 (N_23384,N_18463,N_15731);
nor U23385 (N_23385,N_16771,N_15159);
or U23386 (N_23386,N_16226,N_15432);
nand U23387 (N_23387,N_16835,N_15035);
xnor U23388 (N_23388,N_17386,N_19505);
and U23389 (N_23389,N_17711,N_16291);
xnor U23390 (N_23390,N_15496,N_15164);
xor U23391 (N_23391,N_17707,N_17664);
xnor U23392 (N_23392,N_17338,N_17449);
and U23393 (N_23393,N_17236,N_17357);
nand U23394 (N_23394,N_17359,N_16616);
xnor U23395 (N_23395,N_18680,N_15172);
nor U23396 (N_23396,N_16317,N_16605);
xnor U23397 (N_23397,N_19138,N_17462);
nor U23398 (N_23398,N_16045,N_19557);
or U23399 (N_23399,N_15379,N_16349);
or U23400 (N_23400,N_19440,N_19376);
nand U23401 (N_23401,N_18353,N_16127);
and U23402 (N_23402,N_16834,N_17773);
and U23403 (N_23403,N_19197,N_17897);
nand U23404 (N_23404,N_18370,N_19740);
nand U23405 (N_23405,N_16892,N_15083);
nand U23406 (N_23406,N_18532,N_15760);
or U23407 (N_23407,N_17241,N_16076);
and U23408 (N_23408,N_15474,N_18682);
or U23409 (N_23409,N_19611,N_17932);
and U23410 (N_23410,N_17338,N_18200);
xnor U23411 (N_23411,N_19478,N_17893);
and U23412 (N_23412,N_18405,N_15590);
or U23413 (N_23413,N_15625,N_19886);
and U23414 (N_23414,N_18341,N_16992);
nor U23415 (N_23415,N_16719,N_19116);
nand U23416 (N_23416,N_18583,N_17281);
or U23417 (N_23417,N_19745,N_16753);
nor U23418 (N_23418,N_17437,N_19926);
xor U23419 (N_23419,N_19368,N_16692);
or U23420 (N_23420,N_19464,N_15914);
nor U23421 (N_23421,N_19843,N_16915);
xor U23422 (N_23422,N_16058,N_15170);
xor U23423 (N_23423,N_16609,N_17292);
or U23424 (N_23424,N_17330,N_15773);
or U23425 (N_23425,N_19332,N_16487);
nor U23426 (N_23426,N_18301,N_17794);
and U23427 (N_23427,N_15808,N_17301);
nand U23428 (N_23428,N_17174,N_19074);
xnor U23429 (N_23429,N_17768,N_19070);
xnor U23430 (N_23430,N_15507,N_19965);
nor U23431 (N_23431,N_17403,N_18971);
or U23432 (N_23432,N_16792,N_19688);
xnor U23433 (N_23433,N_18972,N_19963);
nand U23434 (N_23434,N_18083,N_19003);
nor U23435 (N_23435,N_15627,N_17583);
and U23436 (N_23436,N_17398,N_17146);
xnor U23437 (N_23437,N_17118,N_16370);
xor U23438 (N_23438,N_18580,N_18433);
nor U23439 (N_23439,N_16104,N_15642);
nand U23440 (N_23440,N_15131,N_16525);
and U23441 (N_23441,N_19584,N_19683);
nand U23442 (N_23442,N_18226,N_17364);
xnor U23443 (N_23443,N_15841,N_17908);
nand U23444 (N_23444,N_16975,N_17397);
and U23445 (N_23445,N_15343,N_15701);
or U23446 (N_23446,N_18308,N_17555);
or U23447 (N_23447,N_17777,N_19791);
nand U23448 (N_23448,N_18953,N_19942);
nor U23449 (N_23449,N_15159,N_19659);
or U23450 (N_23450,N_17993,N_16067);
xor U23451 (N_23451,N_19349,N_17780);
nor U23452 (N_23452,N_17222,N_15038);
and U23453 (N_23453,N_15268,N_19719);
and U23454 (N_23454,N_18478,N_18296);
nor U23455 (N_23455,N_19997,N_17983);
nor U23456 (N_23456,N_18520,N_17549);
nand U23457 (N_23457,N_16869,N_18656);
and U23458 (N_23458,N_18928,N_18145);
nor U23459 (N_23459,N_15476,N_17509);
nand U23460 (N_23460,N_15017,N_17508);
nand U23461 (N_23461,N_19970,N_19133);
xor U23462 (N_23462,N_19937,N_18433);
and U23463 (N_23463,N_16127,N_19980);
nor U23464 (N_23464,N_19195,N_19370);
xnor U23465 (N_23465,N_17036,N_16827);
xnor U23466 (N_23466,N_16293,N_16716);
or U23467 (N_23467,N_18599,N_15054);
and U23468 (N_23468,N_18887,N_18792);
nand U23469 (N_23469,N_18137,N_15160);
xor U23470 (N_23470,N_15543,N_19861);
nand U23471 (N_23471,N_17155,N_19755);
or U23472 (N_23472,N_19066,N_15244);
nor U23473 (N_23473,N_17064,N_15512);
nor U23474 (N_23474,N_16880,N_17959);
and U23475 (N_23475,N_15874,N_15493);
and U23476 (N_23476,N_16679,N_18593);
nand U23477 (N_23477,N_19430,N_19741);
nand U23478 (N_23478,N_17236,N_18109);
nand U23479 (N_23479,N_15578,N_19383);
or U23480 (N_23480,N_19598,N_16162);
and U23481 (N_23481,N_18219,N_17673);
xnor U23482 (N_23482,N_15656,N_18171);
or U23483 (N_23483,N_19470,N_17556);
and U23484 (N_23484,N_17880,N_18428);
xor U23485 (N_23485,N_16169,N_15549);
or U23486 (N_23486,N_16493,N_17108);
or U23487 (N_23487,N_15576,N_17964);
nor U23488 (N_23488,N_19494,N_17022);
nand U23489 (N_23489,N_19111,N_19674);
or U23490 (N_23490,N_16431,N_19272);
nor U23491 (N_23491,N_15036,N_15975);
xnor U23492 (N_23492,N_16803,N_15391);
nor U23493 (N_23493,N_15384,N_15439);
or U23494 (N_23494,N_16646,N_15838);
nor U23495 (N_23495,N_19946,N_18829);
nor U23496 (N_23496,N_19698,N_16475);
xnor U23497 (N_23497,N_19123,N_19542);
nor U23498 (N_23498,N_16014,N_18515);
and U23499 (N_23499,N_16541,N_16974);
xor U23500 (N_23500,N_17276,N_15291);
nand U23501 (N_23501,N_19544,N_16679);
or U23502 (N_23502,N_17401,N_16190);
xnor U23503 (N_23503,N_15668,N_15622);
and U23504 (N_23504,N_15668,N_18641);
xnor U23505 (N_23505,N_16047,N_19616);
nand U23506 (N_23506,N_17964,N_17523);
nand U23507 (N_23507,N_19299,N_19744);
and U23508 (N_23508,N_15514,N_17883);
xor U23509 (N_23509,N_18760,N_15636);
or U23510 (N_23510,N_18043,N_17117);
xnor U23511 (N_23511,N_16513,N_17366);
xnor U23512 (N_23512,N_19552,N_19141);
or U23513 (N_23513,N_16408,N_19640);
or U23514 (N_23514,N_19644,N_16161);
nor U23515 (N_23515,N_19285,N_17103);
or U23516 (N_23516,N_19160,N_15507);
xor U23517 (N_23517,N_18397,N_15918);
xnor U23518 (N_23518,N_17121,N_19953);
xor U23519 (N_23519,N_15066,N_19593);
nand U23520 (N_23520,N_16571,N_15273);
nor U23521 (N_23521,N_18575,N_18710);
or U23522 (N_23522,N_18126,N_19913);
or U23523 (N_23523,N_17211,N_16687);
nor U23524 (N_23524,N_19535,N_17843);
nor U23525 (N_23525,N_15702,N_15914);
and U23526 (N_23526,N_17202,N_18523);
and U23527 (N_23527,N_19317,N_15036);
nand U23528 (N_23528,N_15339,N_16589);
and U23529 (N_23529,N_16100,N_15065);
or U23530 (N_23530,N_16263,N_17401);
xnor U23531 (N_23531,N_18713,N_16539);
xor U23532 (N_23532,N_18417,N_15944);
nand U23533 (N_23533,N_18507,N_17551);
xor U23534 (N_23534,N_17162,N_15212);
or U23535 (N_23535,N_17986,N_18948);
xor U23536 (N_23536,N_18790,N_15541);
nor U23537 (N_23537,N_17773,N_19408);
or U23538 (N_23538,N_19466,N_18857);
nand U23539 (N_23539,N_15324,N_15553);
nand U23540 (N_23540,N_18886,N_17489);
and U23541 (N_23541,N_16317,N_18102);
nor U23542 (N_23542,N_18602,N_18845);
nand U23543 (N_23543,N_15906,N_15903);
nor U23544 (N_23544,N_15704,N_16968);
and U23545 (N_23545,N_15673,N_15905);
nor U23546 (N_23546,N_16192,N_16129);
nor U23547 (N_23547,N_15631,N_17640);
or U23548 (N_23548,N_15283,N_18340);
and U23549 (N_23549,N_15780,N_15673);
and U23550 (N_23550,N_18856,N_18882);
nand U23551 (N_23551,N_16223,N_19938);
or U23552 (N_23552,N_17802,N_16825);
xnor U23553 (N_23553,N_17479,N_17540);
nand U23554 (N_23554,N_17370,N_15113);
and U23555 (N_23555,N_16782,N_15815);
xor U23556 (N_23556,N_17496,N_19668);
xor U23557 (N_23557,N_19970,N_17414);
and U23558 (N_23558,N_18509,N_15367);
or U23559 (N_23559,N_18761,N_18834);
nand U23560 (N_23560,N_19340,N_18234);
nor U23561 (N_23561,N_18923,N_16416);
nor U23562 (N_23562,N_17032,N_16623);
xor U23563 (N_23563,N_18741,N_19745);
xnor U23564 (N_23564,N_17336,N_19294);
or U23565 (N_23565,N_19321,N_18984);
nand U23566 (N_23566,N_18558,N_15689);
xor U23567 (N_23567,N_19274,N_17098);
nor U23568 (N_23568,N_15575,N_17366);
nand U23569 (N_23569,N_16611,N_17309);
xnor U23570 (N_23570,N_15363,N_18692);
nor U23571 (N_23571,N_19600,N_18829);
or U23572 (N_23572,N_16193,N_15736);
xnor U23573 (N_23573,N_18625,N_16359);
nor U23574 (N_23574,N_15665,N_19368);
xnor U23575 (N_23575,N_16451,N_19395);
nand U23576 (N_23576,N_19038,N_15894);
xnor U23577 (N_23577,N_16677,N_19588);
nor U23578 (N_23578,N_15910,N_19922);
and U23579 (N_23579,N_15650,N_16564);
or U23580 (N_23580,N_18073,N_16681);
or U23581 (N_23581,N_18848,N_19700);
nand U23582 (N_23582,N_17821,N_19771);
nor U23583 (N_23583,N_16904,N_17900);
nor U23584 (N_23584,N_17875,N_15512);
nand U23585 (N_23585,N_19614,N_15042);
and U23586 (N_23586,N_18882,N_18924);
nor U23587 (N_23587,N_18370,N_16111);
nor U23588 (N_23588,N_19585,N_19850);
nor U23589 (N_23589,N_16789,N_16505);
or U23590 (N_23590,N_17774,N_16260);
nand U23591 (N_23591,N_15787,N_19937);
xnor U23592 (N_23592,N_18589,N_16771);
or U23593 (N_23593,N_17298,N_17004);
nand U23594 (N_23594,N_17882,N_18147);
and U23595 (N_23595,N_19616,N_16836);
and U23596 (N_23596,N_19225,N_19589);
nor U23597 (N_23597,N_16943,N_18620);
and U23598 (N_23598,N_17257,N_18447);
nand U23599 (N_23599,N_18202,N_15553);
and U23600 (N_23600,N_19331,N_18060);
or U23601 (N_23601,N_17370,N_16528);
nor U23602 (N_23602,N_18426,N_16407);
nor U23603 (N_23603,N_17772,N_19055);
xor U23604 (N_23604,N_19923,N_18373);
nor U23605 (N_23605,N_18460,N_19187);
nor U23606 (N_23606,N_19763,N_15995);
nor U23607 (N_23607,N_16872,N_15895);
and U23608 (N_23608,N_15415,N_16777);
or U23609 (N_23609,N_18296,N_17702);
or U23610 (N_23610,N_17168,N_19447);
nand U23611 (N_23611,N_15137,N_16312);
nand U23612 (N_23612,N_17210,N_16910);
xnor U23613 (N_23613,N_15184,N_19629);
nand U23614 (N_23614,N_18605,N_19808);
nor U23615 (N_23615,N_18160,N_18691);
nand U23616 (N_23616,N_18841,N_15417);
and U23617 (N_23617,N_16406,N_16974);
and U23618 (N_23618,N_15360,N_17444);
and U23619 (N_23619,N_15179,N_17325);
nor U23620 (N_23620,N_19537,N_17220);
nor U23621 (N_23621,N_15183,N_16419);
or U23622 (N_23622,N_17354,N_15683);
or U23623 (N_23623,N_19776,N_16379);
xor U23624 (N_23624,N_15734,N_16063);
nand U23625 (N_23625,N_16407,N_15391);
nand U23626 (N_23626,N_16552,N_18766);
and U23627 (N_23627,N_16098,N_16006);
nor U23628 (N_23628,N_17887,N_19057);
nand U23629 (N_23629,N_16083,N_15611);
nor U23630 (N_23630,N_18628,N_18513);
or U23631 (N_23631,N_15662,N_15561);
or U23632 (N_23632,N_17707,N_15106);
nor U23633 (N_23633,N_19639,N_18519);
nand U23634 (N_23634,N_18295,N_16364);
nor U23635 (N_23635,N_16952,N_18364);
or U23636 (N_23636,N_17395,N_16953);
xnor U23637 (N_23637,N_19790,N_15647);
nand U23638 (N_23638,N_18524,N_19318);
and U23639 (N_23639,N_19813,N_19566);
or U23640 (N_23640,N_15085,N_17320);
and U23641 (N_23641,N_18441,N_17142);
and U23642 (N_23642,N_19538,N_17966);
xnor U23643 (N_23643,N_15698,N_17112);
and U23644 (N_23644,N_15709,N_15877);
xnor U23645 (N_23645,N_18521,N_19749);
xor U23646 (N_23646,N_16655,N_15991);
nor U23647 (N_23647,N_18217,N_19803);
or U23648 (N_23648,N_16822,N_16994);
xnor U23649 (N_23649,N_16993,N_18973);
xnor U23650 (N_23650,N_15314,N_15687);
or U23651 (N_23651,N_16686,N_15089);
or U23652 (N_23652,N_19393,N_18230);
nand U23653 (N_23653,N_15827,N_15359);
nor U23654 (N_23654,N_15458,N_16078);
and U23655 (N_23655,N_17253,N_17742);
or U23656 (N_23656,N_18090,N_15847);
or U23657 (N_23657,N_16783,N_15789);
nor U23658 (N_23658,N_16020,N_18769);
or U23659 (N_23659,N_16255,N_17750);
and U23660 (N_23660,N_19684,N_16239);
nor U23661 (N_23661,N_16046,N_19272);
nand U23662 (N_23662,N_16694,N_18829);
or U23663 (N_23663,N_15416,N_18097);
nor U23664 (N_23664,N_18025,N_15210);
xnor U23665 (N_23665,N_19574,N_15747);
nor U23666 (N_23666,N_15983,N_16928);
or U23667 (N_23667,N_15811,N_15448);
or U23668 (N_23668,N_19129,N_19527);
nor U23669 (N_23669,N_17630,N_15189);
xor U23670 (N_23670,N_19317,N_16686);
or U23671 (N_23671,N_18985,N_15146);
nor U23672 (N_23672,N_17563,N_18566);
nand U23673 (N_23673,N_18360,N_15988);
or U23674 (N_23674,N_18335,N_15211);
and U23675 (N_23675,N_17446,N_16163);
or U23676 (N_23676,N_15938,N_16027);
xor U23677 (N_23677,N_19335,N_15671);
nand U23678 (N_23678,N_16805,N_16866);
or U23679 (N_23679,N_18240,N_19407);
xnor U23680 (N_23680,N_18665,N_15531);
nor U23681 (N_23681,N_17433,N_16626);
or U23682 (N_23682,N_16230,N_19066);
xor U23683 (N_23683,N_18370,N_16424);
nor U23684 (N_23684,N_19399,N_15307);
xnor U23685 (N_23685,N_17243,N_18056);
xor U23686 (N_23686,N_16928,N_19746);
and U23687 (N_23687,N_18072,N_15788);
and U23688 (N_23688,N_15586,N_19841);
nor U23689 (N_23689,N_16016,N_15144);
nand U23690 (N_23690,N_16431,N_18498);
nand U23691 (N_23691,N_19540,N_18760);
nor U23692 (N_23692,N_18783,N_19324);
and U23693 (N_23693,N_16185,N_16385);
nand U23694 (N_23694,N_17514,N_18189);
nand U23695 (N_23695,N_18090,N_16441);
xor U23696 (N_23696,N_18030,N_18523);
and U23697 (N_23697,N_19379,N_18860);
nor U23698 (N_23698,N_16529,N_17211);
or U23699 (N_23699,N_19705,N_15051);
or U23700 (N_23700,N_15177,N_16265);
and U23701 (N_23701,N_17163,N_19373);
xnor U23702 (N_23702,N_17518,N_15239);
or U23703 (N_23703,N_15589,N_18949);
nand U23704 (N_23704,N_18069,N_15579);
nor U23705 (N_23705,N_15743,N_18948);
or U23706 (N_23706,N_16010,N_18532);
nand U23707 (N_23707,N_17257,N_17616);
and U23708 (N_23708,N_15093,N_16666);
or U23709 (N_23709,N_17329,N_15927);
nor U23710 (N_23710,N_18610,N_16053);
nand U23711 (N_23711,N_18026,N_16549);
xnor U23712 (N_23712,N_19167,N_18004);
nand U23713 (N_23713,N_19004,N_16065);
or U23714 (N_23714,N_19385,N_18617);
and U23715 (N_23715,N_16147,N_17249);
and U23716 (N_23716,N_19066,N_17377);
and U23717 (N_23717,N_15234,N_15272);
and U23718 (N_23718,N_18372,N_19769);
and U23719 (N_23719,N_19041,N_19074);
xor U23720 (N_23720,N_19581,N_15154);
nand U23721 (N_23721,N_15843,N_17998);
nand U23722 (N_23722,N_18694,N_15536);
and U23723 (N_23723,N_19977,N_18292);
xor U23724 (N_23724,N_18871,N_18529);
or U23725 (N_23725,N_18703,N_18994);
nand U23726 (N_23726,N_17497,N_17062);
nand U23727 (N_23727,N_19147,N_18669);
nor U23728 (N_23728,N_16735,N_15760);
xor U23729 (N_23729,N_19229,N_15820);
and U23730 (N_23730,N_17715,N_19124);
xnor U23731 (N_23731,N_17085,N_15442);
nor U23732 (N_23732,N_15765,N_17214);
or U23733 (N_23733,N_18546,N_17892);
nor U23734 (N_23734,N_19796,N_17287);
nand U23735 (N_23735,N_18648,N_17799);
and U23736 (N_23736,N_18493,N_19128);
xor U23737 (N_23737,N_18791,N_19768);
xor U23738 (N_23738,N_15566,N_16278);
nand U23739 (N_23739,N_19216,N_18406);
nor U23740 (N_23740,N_17715,N_16863);
or U23741 (N_23741,N_15130,N_18977);
nand U23742 (N_23742,N_15248,N_19488);
and U23743 (N_23743,N_19990,N_17482);
and U23744 (N_23744,N_19961,N_19393);
xnor U23745 (N_23745,N_15718,N_18938);
nor U23746 (N_23746,N_19681,N_15742);
and U23747 (N_23747,N_15733,N_17318);
and U23748 (N_23748,N_16583,N_18196);
nor U23749 (N_23749,N_19253,N_15938);
xor U23750 (N_23750,N_19076,N_15978);
nor U23751 (N_23751,N_18564,N_18150);
and U23752 (N_23752,N_15984,N_15430);
xnor U23753 (N_23753,N_19848,N_19471);
nor U23754 (N_23754,N_17182,N_17780);
and U23755 (N_23755,N_17359,N_17409);
nand U23756 (N_23756,N_19869,N_16949);
and U23757 (N_23757,N_18484,N_16892);
or U23758 (N_23758,N_16402,N_15111);
nor U23759 (N_23759,N_16396,N_17814);
xor U23760 (N_23760,N_16453,N_16030);
and U23761 (N_23761,N_18142,N_16202);
and U23762 (N_23762,N_15217,N_17976);
or U23763 (N_23763,N_18710,N_18626);
xor U23764 (N_23764,N_15389,N_16555);
or U23765 (N_23765,N_16551,N_19210);
or U23766 (N_23766,N_17533,N_16811);
xnor U23767 (N_23767,N_19065,N_19786);
or U23768 (N_23768,N_17063,N_17425);
nand U23769 (N_23769,N_18879,N_17811);
xor U23770 (N_23770,N_16004,N_15655);
xnor U23771 (N_23771,N_15761,N_18644);
nand U23772 (N_23772,N_18127,N_18724);
and U23773 (N_23773,N_18967,N_15530);
or U23774 (N_23774,N_19858,N_19340);
and U23775 (N_23775,N_19928,N_15771);
xnor U23776 (N_23776,N_16235,N_15953);
and U23777 (N_23777,N_15374,N_17088);
nor U23778 (N_23778,N_17122,N_19638);
nor U23779 (N_23779,N_15096,N_16423);
and U23780 (N_23780,N_19914,N_18014);
nor U23781 (N_23781,N_19449,N_17304);
and U23782 (N_23782,N_15664,N_16723);
or U23783 (N_23783,N_16324,N_15817);
and U23784 (N_23784,N_17984,N_17824);
nor U23785 (N_23785,N_17280,N_16368);
nand U23786 (N_23786,N_15772,N_17963);
and U23787 (N_23787,N_17065,N_18333);
and U23788 (N_23788,N_17016,N_18365);
xnor U23789 (N_23789,N_15808,N_17010);
nor U23790 (N_23790,N_18148,N_18509);
nand U23791 (N_23791,N_18927,N_15663);
or U23792 (N_23792,N_18421,N_18743);
xnor U23793 (N_23793,N_15625,N_15788);
xor U23794 (N_23794,N_16898,N_16538);
nor U23795 (N_23795,N_19899,N_17236);
nor U23796 (N_23796,N_18183,N_16774);
or U23797 (N_23797,N_17558,N_15642);
and U23798 (N_23798,N_19617,N_18586);
xor U23799 (N_23799,N_18840,N_17747);
nand U23800 (N_23800,N_19185,N_18889);
or U23801 (N_23801,N_18292,N_18180);
xor U23802 (N_23802,N_17207,N_18127);
and U23803 (N_23803,N_16388,N_19194);
or U23804 (N_23804,N_18649,N_15735);
nand U23805 (N_23805,N_17062,N_18769);
nor U23806 (N_23806,N_18887,N_18598);
or U23807 (N_23807,N_17896,N_19482);
xnor U23808 (N_23808,N_18505,N_17962);
xnor U23809 (N_23809,N_17344,N_15180);
and U23810 (N_23810,N_16620,N_16484);
or U23811 (N_23811,N_18884,N_17151);
xnor U23812 (N_23812,N_18808,N_19541);
xor U23813 (N_23813,N_15837,N_19152);
xor U23814 (N_23814,N_18608,N_19183);
xor U23815 (N_23815,N_19476,N_15729);
nand U23816 (N_23816,N_15365,N_17177);
or U23817 (N_23817,N_16644,N_16342);
and U23818 (N_23818,N_15417,N_18670);
and U23819 (N_23819,N_17406,N_18228);
and U23820 (N_23820,N_19400,N_19809);
nand U23821 (N_23821,N_19594,N_16707);
or U23822 (N_23822,N_15858,N_19126);
or U23823 (N_23823,N_19113,N_17369);
xnor U23824 (N_23824,N_18763,N_19826);
or U23825 (N_23825,N_16000,N_16136);
or U23826 (N_23826,N_15745,N_15581);
nor U23827 (N_23827,N_19364,N_17009);
xnor U23828 (N_23828,N_17677,N_15206);
xor U23829 (N_23829,N_15747,N_19965);
nand U23830 (N_23830,N_15003,N_16054);
nor U23831 (N_23831,N_18994,N_15949);
xnor U23832 (N_23832,N_16828,N_16389);
nor U23833 (N_23833,N_18007,N_18251);
nor U23834 (N_23834,N_17289,N_17875);
or U23835 (N_23835,N_19580,N_18629);
or U23836 (N_23836,N_16325,N_18780);
or U23837 (N_23837,N_19735,N_16011);
or U23838 (N_23838,N_16586,N_17895);
xnor U23839 (N_23839,N_16846,N_15756);
nand U23840 (N_23840,N_19136,N_15571);
or U23841 (N_23841,N_19512,N_17913);
nand U23842 (N_23842,N_15606,N_16079);
nor U23843 (N_23843,N_16719,N_15369);
nand U23844 (N_23844,N_16944,N_18680);
or U23845 (N_23845,N_17042,N_16278);
and U23846 (N_23846,N_17940,N_18342);
nand U23847 (N_23847,N_18131,N_18807);
or U23848 (N_23848,N_19900,N_17760);
nand U23849 (N_23849,N_15065,N_15652);
nor U23850 (N_23850,N_15182,N_18554);
xor U23851 (N_23851,N_19082,N_18348);
xor U23852 (N_23852,N_18867,N_15104);
xor U23853 (N_23853,N_16347,N_15984);
and U23854 (N_23854,N_16346,N_15847);
or U23855 (N_23855,N_16656,N_16974);
and U23856 (N_23856,N_15358,N_18414);
nand U23857 (N_23857,N_15688,N_16733);
nand U23858 (N_23858,N_16261,N_18431);
nor U23859 (N_23859,N_15978,N_18973);
nand U23860 (N_23860,N_18521,N_16999);
or U23861 (N_23861,N_17811,N_15864);
nand U23862 (N_23862,N_17207,N_16239);
and U23863 (N_23863,N_15545,N_18524);
or U23864 (N_23864,N_18991,N_17263);
and U23865 (N_23865,N_15023,N_16540);
and U23866 (N_23866,N_17792,N_19518);
nand U23867 (N_23867,N_16775,N_15533);
and U23868 (N_23868,N_17351,N_15684);
xor U23869 (N_23869,N_17342,N_19827);
xnor U23870 (N_23870,N_18044,N_15770);
xnor U23871 (N_23871,N_16697,N_18242);
xnor U23872 (N_23872,N_18702,N_15660);
nor U23873 (N_23873,N_17990,N_15678);
and U23874 (N_23874,N_17522,N_16083);
and U23875 (N_23875,N_15574,N_17133);
or U23876 (N_23876,N_17318,N_17104);
xnor U23877 (N_23877,N_17505,N_15655);
nand U23878 (N_23878,N_15151,N_19397);
nand U23879 (N_23879,N_17009,N_17137);
xnor U23880 (N_23880,N_15282,N_17785);
nor U23881 (N_23881,N_17483,N_15758);
nor U23882 (N_23882,N_15757,N_18699);
and U23883 (N_23883,N_18766,N_16066);
or U23884 (N_23884,N_18793,N_15278);
and U23885 (N_23885,N_17474,N_15561);
and U23886 (N_23886,N_15743,N_19056);
nor U23887 (N_23887,N_17900,N_16021);
or U23888 (N_23888,N_18471,N_19965);
nand U23889 (N_23889,N_17274,N_17299);
nor U23890 (N_23890,N_15888,N_16288);
xor U23891 (N_23891,N_15849,N_18111);
xnor U23892 (N_23892,N_19088,N_15027);
and U23893 (N_23893,N_18269,N_17968);
or U23894 (N_23894,N_19721,N_19032);
nor U23895 (N_23895,N_18020,N_19010);
nor U23896 (N_23896,N_15380,N_18366);
nor U23897 (N_23897,N_19860,N_16245);
nand U23898 (N_23898,N_16031,N_16754);
and U23899 (N_23899,N_18262,N_19624);
and U23900 (N_23900,N_15592,N_17834);
xnor U23901 (N_23901,N_19423,N_18333);
and U23902 (N_23902,N_17431,N_19270);
and U23903 (N_23903,N_19235,N_16127);
or U23904 (N_23904,N_18028,N_17713);
and U23905 (N_23905,N_17076,N_15136);
and U23906 (N_23906,N_15810,N_16046);
xor U23907 (N_23907,N_19648,N_17708);
and U23908 (N_23908,N_16972,N_17730);
and U23909 (N_23909,N_16179,N_15153);
xor U23910 (N_23910,N_15274,N_19411);
nor U23911 (N_23911,N_19628,N_16984);
or U23912 (N_23912,N_16695,N_19351);
and U23913 (N_23913,N_15763,N_15185);
nand U23914 (N_23914,N_16052,N_18312);
nor U23915 (N_23915,N_19968,N_15611);
nor U23916 (N_23916,N_17592,N_19131);
and U23917 (N_23917,N_17904,N_19890);
xnor U23918 (N_23918,N_19173,N_18717);
xor U23919 (N_23919,N_19889,N_16525);
xnor U23920 (N_23920,N_17384,N_18544);
nand U23921 (N_23921,N_19715,N_19513);
nor U23922 (N_23922,N_15396,N_19701);
nand U23923 (N_23923,N_18746,N_15499);
nand U23924 (N_23924,N_19587,N_18357);
or U23925 (N_23925,N_15482,N_17778);
and U23926 (N_23926,N_16294,N_19374);
nand U23927 (N_23927,N_19857,N_16615);
nand U23928 (N_23928,N_19415,N_15835);
nor U23929 (N_23929,N_18852,N_15596);
nand U23930 (N_23930,N_17214,N_18384);
and U23931 (N_23931,N_19313,N_18282);
and U23932 (N_23932,N_16842,N_18494);
nor U23933 (N_23933,N_17106,N_18793);
nand U23934 (N_23934,N_15127,N_17575);
nor U23935 (N_23935,N_16188,N_18239);
nor U23936 (N_23936,N_19586,N_19555);
and U23937 (N_23937,N_19387,N_16431);
and U23938 (N_23938,N_15466,N_19044);
nand U23939 (N_23939,N_17486,N_18575);
or U23940 (N_23940,N_16336,N_17790);
nor U23941 (N_23941,N_18994,N_18820);
xor U23942 (N_23942,N_17031,N_17223);
and U23943 (N_23943,N_17615,N_18991);
xnor U23944 (N_23944,N_19608,N_15519);
and U23945 (N_23945,N_18700,N_19712);
nor U23946 (N_23946,N_17442,N_17030);
nand U23947 (N_23947,N_16779,N_16301);
or U23948 (N_23948,N_18284,N_18014);
nor U23949 (N_23949,N_19917,N_19541);
and U23950 (N_23950,N_17314,N_18501);
and U23951 (N_23951,N_19673,N_16503);
and U23952 (N_23952,N_18926,N_15739);
or U23953 (N_23953,N_19647,N_18849);
nand U23954 (N_23954,N_19606,N_16262);
nor U23955 (N_23955,N_16492,N_15518);
and U23956 (N_23956,N_17591,N_18796);
nor U23957 (N_23957,N_16010,N_16616);
or U23958 (N_23958,N_15527,N_16545);
or U23959 (N_23959,N_17879,N_15325);
nor U23960 (N_23960,N_18681,N_16314);
nor U23961 (N_23961,N_16872,N_15203);
and U23962 (N_23962,N_16681,N_17166);
or U23963 (N_23963,N_17590,N_18857);
or U23964 (N_23964,N_15115,N_19486);
or U23965 (N_23965,N_18333,N_18615);
or U23966 (N_23966,N_19211,N_19369);
nand U23967 (N_23967,N_15115,N_17892);
nor U23968 (N_23968,N_19676,N_15577);
nor U23969 (N_23969,N_16562,N_16953);
xor U23970 (N_23970,N_17815,N_19312);
and U23971 (N_23971,N_15029,N_16941);
nand U23972 (N_23972,N_16333,N_18614);
or U23973 (N_23973,N_16609,N_16788);
and U23974 (N_23974,N_16183,N_16818);
nor U23975 (N_23975,N_18322,N_17512);
or U23976 (N_23976,N_15789,N_19562);
xor U23977 (N_23977,N_19619,N_19407);
and U23978 (N_23978,N_17945,N_18338);
xnor U23979 (N_23979,N_19198,N_15105);
xor U23980 (N_23980,N_16671,N_19314);
and U23981 (N_23981,N_16789,N_16521);
or U23982 (N_23982,N_15167,N_17795);
nor U23983 (N_23983,N_19332,N_17147);
and U23984 (N_23984,N_15431,N_16971);
xor U23985 (N_23985,N_18486,N_15965);
nor U23986 (N_23986,N_16018,N_17453);
xor U23987 (N_23987,N_19331,N_15761);
or U23988 (N_23988,N_15024,N_17193);
nand U23989 (N_23989,N_19617,N_17821);
or U23990 (N_23990,N_19556,N_15615);
xnor U23991 (N_23991,N_17403,N_19804);
nor U23992 (N_23992,N_18132,N_18255);
and U23993 (N_23993,N_17841,N_15402);
or U23994 (N_23994,N_15820,N_17913);
or U23995 (N_23995,N_17535,N_15321);
xor U23996 (N_23996,N_15947,N_19197);
xnor U23997 (N_23997,N_17175,N_19677);
nand U23998 (N_23998,N_16361,N_15986);
nand U23999 (N_23999,N_17503,N_17883);
xnor U24000 (N_24000,N_18615,N_19249);
or U24001 (N_24001,N_16512,N_15446);
or U24002 (N_24002,N_18386,N_18837);
nand U24003 (N_24003,N_18229,N_16818);
xor U24004 (N_24004,N_16162,N_18520);
nor U24005 (N_24005,N_18938,N_18955);
or U24006 (N_24006,N_15280,N_18692);
nor U24007 (N_24007,N_15893,N_18594);
xor U24008 (N_24008,N_17916,N_16594);
nor U24009 (N_24009,N_18041,N_16547);
nand U24010 (N_24010,N_16563,N_15301);
or U24011 (N_24011,N_19447,N_16125);
nor U24012 (N_24012,N_17537,N_18975);
nand U24013 (N_24013,N_15003,N_15327);
and U24014 (N_24014,N_16209,N_17523);
xnor U24015 (N_24015,N_16765,N_18506);
nor U24016 (N_24016,N_16383,N_18909);
and U24017 (N_24017,N_19484,N_17368);
and U24018 (N_24018,N_15400,N_19191);
xor U24019 (N_24019,N_18979,N_15841);
or U24020 (N_24020,N_18476,N_15780);
and U24021 (N_24021,N_19744,N_15529);
and U24022 (N_24022,N_19040,N_18195);
and U24023 (N_24023,N_16656,N_15108);
and U24024 (N_24024,N_16791,N_18321);
nand U24025 (N_24025,N_16260,N_16239);
nor U24026 (N_24026,N_18308,N_19010);
xnor U24027 (N_24027,N_15607,N_18312);
and U24028 (N_24028,N_15436,N_17875);
and U24029 (N_24029,N_15247,N_18329);
nor U24030 (N_24030,N_19476,N_18566);
nand U24031 (N_24031,N_18752,N_17541);
nor U24032 (N_24032,N_15582,N_18155);
nor U24033 (N_24033,N_15834,N_16969);
xor U24034 (N_24034,N_17178,N_15060);
nand U24035 (N_24035,N_15312,N_16956);
nand U24036 (N_24036,N_18833,N_17250);
or U24037 (N_24037,N_18274,N_16373);
xor U24038 (N_24038,N_16840,N_18210);
or U24039 (N_24039,N_18601,N_17917);
and U24040 (N_24040,N_17208,N_19652);
nor U24041 (N_24041,N_16293,N_15287);
and U24042 (N_24042,N_18561,N_17191);
xnor U24043 (N_24043,N_15738,N_18612);
and U24044 (N_24044,N_18009,N_16642);
or U24045 (N_24045,N_18445,N_16600);
xnor U24046 (N_24046,N_18408,N_15377);
or U24047 (N_24047,N_15798,N_15646);
or U24048 (N_24048,N_15667,N_19040);
nor U24049 (N_24049,N_16838,N_15334);
xor U24050 (N_24050,N_18267,N_18262);
xor U24051 (N_24051,N_18227,N_19920);
nand U24052 (N_24052,N_16529,N_19750);
or U24053 (N_24053,N_15389,N_16160);
xor U24054 (N_24054,N_19204,N_16371);
and U24055 (N_24055,N_16825,N_18897);
nand U24056 (N_24056,N_16311,N_16426);
nand U24057 (N_24057,N_17103,N_15045);
and U24058 (N_24058,N_17548,N_16519);
or U24059 (N_24059,N_17262,N_19288);
nor U24060 (N_24060,N_17823,N_19950);
nand U24061 (N_24061,N_15346,N_19077);
xor U24062 (N_24062,N_18689,N_18813);
xnor U24063 (N_24063,N_17930,N_17217);
xnor U24064 (N_24064,N_16884,N_16869);
xnor U24065 (N_24065,N_19058,N_15512);
or U24066 (N_24066,N_17602,N_19176);
nor U24067 (N_24067,N_15300,N_18372);
xnor U24068 (N_24068,N_15655,N_18494);
and U24069 (N_24069,N_16535,N_16485);
xor U24070 (N_24070,N_19192,N_19420);
xnor U24071 (N_24071,N_16232,N_15675);
xor U24072 (N_24072,N_16960,N_15327);
xnor U24073 (N_24073,N_17240,N_19874);
nand U24074 (N_24074,N_19520,N_17642);
and U24075 (N_24075,N_17539,N_15493);
and U24076 (N_24076,N_16381,N_18319);
nor U24077 (N_24077,N_15113,N_19015);
xnor U24078 (N_24078,N_15148,N_19802);
nand U24079 (N_24079,N_17009,N_18931);
xor U24080 (N_24080,N_19095,N_19242);
or U24081 (N_24081,N_16305,N_15532);
xnor U24082 (N_24082,N_16818,N_17735);
nand U24083 (N_24083,N_17981,N_19035);
xnor U24084 (N_24084,N_19241,N_15757);
or U24085 (N_24085,N_18292,N_19253);
or U24086 (N_24086,N_18973,N_19100);
xor U24087 (N_24087,N_17697,N_16408);
or U24088 (N_24088,N_18576,N_15102);
nand U24089 (N_24089,N_19979,N_19147);
nor U24090 (N_24090,N_16879,N_19645);
and U24091 (N_24091,N_18041,N_18295);
or U24092 (N_24092,N_16161,N_15587);
xnor U24093 (N_24093,N_19275,N_17914);
nor U24094 (N_24094,N_19915,N_15017);
nand U24095 (N_24095,N_18014,N_19569);
and U24096 (N_24096,N_17814,N_19273);
nor U24097 (N_24097,N_16415,N_15401);
xnor U24098 (N_24098,N_18456,N_16916);
nand U24099 (N_24099,N_17044,N_15540);
and U24100 (N_24100,N_16511,N_18750);
and U24101 (N_24101,N_18991,N_19425);
nor U24102 (N_24102,N_16183,N_16947);
xor U24103 (N_24103,N_17436,N_15021);
nand U24104 (N_24104,N_15107,N_18557);
nor U24105 (N_24105,N_17530,N_18728);
nor U24106 (N_24106,N_19487,N_18506);
nor U24107 (N_24107,N_16402,N_15058);
or U24108 (N_24108,N_16222,N_17542);
and U24109 (N_24109,N_16711,N_15200);
nor U24110 (N_24110,N_16405,N_17030);
nand U24111 (N_24111,N_17248,N_19843);
and U24112 (N_24112,N_16302,N_18936);
nand U24113 (N_24113,N_16163,N_17188);
or U24114 (N_24114,N_18339,N_16141);
xnor U24115 (N_24115,N_16661,N_16621);
xnor U24116 (N_24116,N_18780,N_17817);
and U24117 (N_24117,N_15389,N_15157);
and U24118 (N_24118,N_15465,N_15249);
or U24119 (N_24119,N_16887,N_15938);
xor U24120 (N_24120,N_16496,N_16058);
nor U24121 (N_24121,N_15892,N_18372);
xnor U24122 (N_24122,N_18782,N_18009);
xor U24123 (N_24123,N_15044,N_19748);
nand U24124 (N_24124,N_19217,N_18605);
xnor U24125 (N_24125,N_18921,N_19009);
xor U24126 (N_24126,N_15077,N_15020);
xor U24127 (N_24127,N_19914,N_15998);
nand U24128 (N_24128,N_17413,N_19716);
or U24129 (N_24129,N_15325,N_17884);
nand U24130 (N_24130,N_18261,N_15879);
xnor U24131 (N_24131,N_16948,N_19506);
nor U24132 (N_24132,N_19542,N_15319);
nor U24133 (N_24133,N_16087,N_18023);
nor U24134 (N_24134,N_18091,N_17750);
nor U24135 (N_24135,N_16837,N_16525);
nand U24136 (N_24136,N_15969,N_16032);
or U24137 (N_24137,N_18865,N_18564);
nor U24138 (N_24138,N_16004,N_19005);
xor U24139 (N_24139,N_19260,N_16988);
or U24140 (N_24140,N_16181,N_17616);
nand U24141 (N_24141,N_19515,N_19875);
or U24142 (N_24142,N_19050,N_15181);
and U24143 (N_24143,N_18086,N_15043);
or U24144 (N_24144,N_19651,N_19487);
and U24145 (N_24145,N_16659,N_15251);
nor U24146 (N_24146,N_19539,N_18403);
or U24147 (N_24147,N_15684,N_19128);
nand U24148 (N_24148,N_19048,N_15788);
xor U24149 (N_24149,N_19717,N_18857);
nand U24150 (N_24150,N_18857,N_16263);
nor U24151 (N_24151,N_19084,N_19192);
nand U24152 (N_24152,N_19362,N_17226);
xor U24153 (N_24153,N_19092,N_15508);
xor U24154 (N_24154,N_19971,N_18198);
nand U24155 (N_24155,N_15354,N_17009);
and U24156 (N_24156,N_16164,N_16776);
or U24157 (N_24157,N_17472,N_18154);
xor U24158 (N_24158,N_17103,N_18868);
nand U24159 (N_24159,N_15212,N_19768);
and U24160 (N_24160,N_17093,N_15084);
nor U24161 (N_24161,N_19165,N_18299);
nor U24162 (N_24162,N_18259,N_16544);
xnor U24163 (N_24163,N_19975,N_17064);
and U24164 (N_24164,N_16154,N_15048);
nor U24165 (N_24165,N_15196,N_15625);
and U24166 (N_24166,N_18789,N_15193);
xnor U24167 (N_24167,N_19499,N_17159);
nor U24168 (N_24168,N_17894,N_16465);
nor U24169 (N_24169,N_18654,N_19414);
or U24170 (N_24170,N_19829,N_18156);
nand U24171 (N_24171,N_16848,N_18450);
or U24172 (N_24172,N_18338,N_15067);
nor U24173 (N_24173,N_16816,N_15055);
or U24174 (N_24174,N_18925,N_19299);
xor U24175 (N_24175,N_17095,N_15021);
nand U24176 (N_24176,N_19816,N_18773);
xor U24177 (N_24177,N_19761,N_15462);
and U24178 (N_24178,N_17569,N_17521);
and U24179 (N_24179,N_17535,N_18471);
xor U24180 (N_24180,N_16641,N_16463);
nor U24181 (N_24181,N_17967,N_15950);
or U24182 (N_24182,N_16945,N_17497);
or U24183 (N_24183,N_18172,N_19638);
nand U24184 (N_24184,N_19419,N_15497);
nand U24185 (N_24185,N_18476,N_18773);
nor U24186 (N_24186,N_15376,N_15714);
and U24187 (N_24187,N_15817,N_17270);
and U24188 (N_24188,N_15530,N_17197);
nor U24189 (N_24189,N_19945,N_16096);
nor U24190 (N_24190,N_16109,N_18521);
xnor U24191 (N_24191,N_15272,N_17700);
nand U24192 (N_24192,N_16512,N_18254);
nor U24193 (N_24193,N_18300,N_15447);
nor U24194 (N_24194,N_19730,N_18952);
or U24195 (N_24195,N_18641,N_19915);
nor U24196 (N_24196,N_18082,N_18238);
or U24197 (N_24197,N_17584,N_16997);
xor U24198 (N_24198,N_19763,N_17615);
nand U24199 (N_24199,N_17799,N_18421);
or U24200 (N_24200,N_15083,N_18946);
and U24201 (N_24201,N_19139,N_18691);
nor U24202 (N_24202,N_15083,N_18023);
and U24203 (N_24203,N_19627,N_16989);
nor U24204 (N_24204,N_18690,N_17228);
and U24205 (N_24205,N_17108,N_15825);
nand U24206 (N_24206,N_19201,N_17545);
nor U24207 (N_24207,N_17151,N_17095);
nor U24208 (N_24208,N_19258,N_17771);
nor U24209 (N_24209,N_18805,N_15262);
and U24210 (N_24210,N_16698,N_18293);
nor U24211 (N_24211,N_17631,N_18807);
or U24212 (N_24212,N_16395,N_16431);
nor U24213 (N_24213,N_19739,N_19096);
nor U24214 (N_24214,N_17074,N_17784);
and U24215 (N_24215,N_19587,N_16539);
or U24216 (N_24216,N_15952,N_16543);
and U24217 (N_24217,N_18086,N_17492);
nor U24218 (N_24218,N_15092,N_15605);
xnor U24219 (N_24219,N_19624,N_16091);
nand U24220 (N_24220,N_19188,N_19331);
nor U24221 (N_24221,N_15665,N_17534);
nand U24222 (N_24222,N_18933,N_15134);
and U24223 (N_24223,N_19280,N_19616);
nor U24224 (N_24224,N_18005,N_18795);
nand U24225 (N_24225,N_18711,N_18805);
and U24226 (N_24226,N_16973,N_15510);
nor U24227 (N_24227,N_15451,N_17646);
xnor U24228 (N_24228,N_19747,N_18984);
or U24229 (N_24229,N_19447,N_15421);
nand U24230 (N_24230,N_17643,N_17661);
xnor U24231 (N_24231,N_19438,N_18786);
and U24232 (N_24232,N_18214,N_19745);
or U24233 (N_24233,N_17538,N_16397);
and U24234 (N_24234,N_15644,N_18203);
nand U24235 (N_24235,N_19942,N_16608);
or U24236 (N_24236,N_16337,N_15700);
nand U24237 (N_24237,N_15836,N_19015);
or U24238 (N_24238,N_15423,N_18981);
and U24239 (N_24239,N_16435,N_16444);
or U24240 (N_24240,N_17112,N_18790);
and U24241 (N_24241,N_15501,N_16125);
nand U24242 (N_24242,N_17712,N_16882);
or U24243 (N_24243,N_15283,N_19168);
and U24244 (N_24244,N_17014,N_16889);
xor U24245 (N_24245,N_18047,N_18501);
nor U24246 (N_24246,N_17441,N_16315);
nand U24247 (N_24247,N_15143,N_17074);
and U24248 (N_24248,N_18667,N_19757);
xnor U24249 (N_24249,N_15485,N_15287);
xnor U24250 (N_24250,N_18489,N_19794);
xnor U24251 (N_24251,N_19697,N_18230);
or U24252 (N_24252,N_19812,N_15397);
xor U24253 (N_24253,N_19005,N_17459);
and U24254 (N_24254,N_19632,N_16605);
and U24255 (N_24255,N_16128,N_19285);
nand U24256 (N_24256,N_17253,N_16923);
xnor U24257 (N_24257,N_19416,N_15758);
xnor U24258 (N_24258,N_15357,N_16467);
xor U24259 (N_24259,N_17891,N_17273);
xnor U24260 (N_24260,N_18151,N_16177);
or U24261 (N_24261,N_19032,N_16224);
nand U24262 (N_24262,N_18336,N_18573);
nand U24263 (N_24263,N_19717,N_19609);
nor U24264 (N_24264,N_17257,N_19019);
nand U24265 (N_24265,N_15601,N_16470);
nand U24266 (N_24266,N_17524,N_16399);
xnor U24267 (N_24267,N_17359,N_18313);
xor U24268 (N_24268,N_17496,N_18614);
xnor U24269 (N_24269,N_16166,N_17660);
nand U24270 (N_24270,N_16229,N_19063);
nand U24271 (N_24271,N_15500,N_15443);
and U24272 (N_24272,N_16949,N_16569);
xor U24273 (N_24273,N_17182,N_15091);
nor U24274 (N_24274,N_19535,N_19189);
or U24275 (N_24275,N_17976,N_18294);
nor U24276 (N_24276,N_17916,N_17124);
and U24277 (N_24277,N_18834,N_15665);
or U24278 (N_24278,N_17054,N_15830);
and U24279 (N_24279,N_17143,N_15465);
and U24280 (N_24280,N_19968,N_16631);
or U24281 (N_24281,N_16583,N_19352);
xor U24282 (N_24282,N_17958,N_17877);
or U24283 (N_24283,N_19317,N_16897);
nor U24284 (N_24284,N_17540,N_18785);
nand U24285 (N_24285,N_18436,N_19373);
and U24286 (N_24286,N_18541,N_17222);
nor U24287 (N_24287,N_18256,N_17375);
nand U24288 (N_24288,N_19593,N_18752);
nand U24289 (N_24289,N_18402,N_16718);
xor U24290 (N_24290,N_19701,N_18809);
nor U24291 (N_24291,N_18125,N_18917);
nor U24292 (N_24292,N_17889,N_17347);
and U24293 (N_24293,N_19588,N_16071);
nand U24294 (N_24294,N_18050,N_19458);
or U24295 (N_24295,N_18583,N_17752);
nor U24296 (N_24296,N_17058,N_15372);
nor U24297 (N_24297,N_17522,N_15382);
xor U24298 (N_24298,N_19803,N_19020);
or U24299 (N_24299,N_16056,N_15632);
nand U24300 (N_24300,N_18912,N_19807);
and U24301 (N_24301,N_18222,N_18555);
nor U24302 (N_24302,N_18676,N_15202);
nor U24303 (N_24303,N_15136,N_18471);
and U24304 (N_24304,N_16979,N_17075);
xnor U24305 (N_24305,N_16942,N_18655);
and U24306 (N_24306,N_16203,N_17111);
nor U24307 (N_24307,N_18729,N_16885);
and U24308 (N_24308,N_19324,N_17805);
xor U24309 (N_24309,N_17783,N_17535);
and U24310 (N_24310,N_18049,N_18470);
nand U24311 (N_24311,N_16936,N_19443);
or U24312 (N_24312,N_18265,N_19699);
nand U24313 (N_24313,N_15685,N_16378);
and U24314 (N_24314,N_19577,N_16125);
or U24315 (N_24315,N_19717,N_15033);
nand U24316 (N_24316,N_17337,N_19229);
and U24317 (N_24317,N_19394,N_18949);
or U24318 (N_24318,N_19710,N_17070);
nand U24319 (N_24319,N_15545,N_15660);
and U24320 (N_24320,N_17891,N_18801);
or U24321 (N_24321,N_17953,N_18134);
xor U24322 (N_24322,N_18680,N_15309);
nand U24323 (N_24323,N_15566,N_18265);
or U24324 (N_24324,N_19373,N_16071);
xor U24325 (N_24325,N_16238,N_16663);
xnor U24326 (N_24326,N_19854,N_18971);
xnor U24327 (N_24327,N_17140,N_19637);
nor U24328 (N_24328,N_15061,N_18667);
xnor U24329 (N_24329,N_16511,N_16514);
and U24330 (N_24330,N_19553,N_17703);
nand U24331 (N_24331,N_17479,N_16031);
nand U24332 (N_24332,N_15590,N_19783);
nand U24333 (N_24333,N_16343,N_16481);
nand U24334 (N_24334,N_18579,N_16405);
and U24335 (N_24335,N_17480,N_17452);
xor U24336 (N_24336,N_15174,N_17572);
or U24337 (N_24337,N_15197,N_15035);
or U24338 (N_24338,N_16826,N_17491);
and U24339 (N_24339,N_16021,N_17337);
nand U24340 (N_24340,N_16770,N_19097);
or U24341 (N_24341,N_15608,N_16469);
nor U24342 (N_24342,N_16869,N_15163);
xnor U24343 (N_24343,N_16297,N_19383);
xor U24344 (N_24344,N_17460,N_17745);
nor U24345 (N_24345,N_18150,N_16991);
xor U24346 (N_24346,N_16818,N_19312);
nand U24347 (N_24347,N_17403,N_18136);
and U24348 (N_24348,N_19704,N_19192);
nand U24349 (N_24349,N_18948,N_15554);
nor U24350 (N_24350,N_18037,N_18187);
nand U24351 (N_24351,N_15834,N_17161);
nor U24352 (N_24352,N_15855,N_17969);
xor U24353 (N_24353,N_17492,N_15837);
and U24354 (N_24354,N_17467,N_17012);
xor U24355 (N_24355,N_18916,N_17682);
nor U24356 (N_24356,N_18186,N_17028);
and U24357 (N_24357,N_15900,N_18972);
or U24358 (N_24358,N_15859,N_17664);
or U24359 (N_24359,N_17638,N_15479);
or U24360 (N_24360,N_16022,N_18758);
and U24361 (N_24361,N_18060,N_19732);
xor U24362 (N_24362,N_19705,N_15146);
xnor U24363 (N_24363,N_17875,N_15214);
or U24364 (N_24364,N_18218,N_17066);
xnor U24365 (N_24365,N_17831,N_16735);
nor U24366 (N_24366,N_18975,N_19687);
nor U24367 (N_24367,N_15469,N_15696);
xor U24368 (N_24368,N_15478,N_15792);
xor U24369 (N_24369,N_16152,N_17337);
xnor U24370 (N_24370,N_19334,N_17032);
or U24371 (N_24371,N_17339,N_19982);
nand U24372 (N_24372,N_17812,N_18158);
xor U24373 (N_24373,N_15229,N_16062);
nor U24374 (N_24374,N_15968,N_19538);
or U24375 (N_24375,N_16243,N_19870);
nor U24376 (N_24376,N_18354,N_17312);
nand U24377 (N_24377,N_18161,N_19154);
xnor U24378 (N_24378,N_17206,N_17458);
nand U24379 (N_24379,N_19936,N_15341);
xor U24380 (N_24380,N_16499,N_15028);
and U24381 (N_24381,N_16080,N_19839);
nand U24382 (N_24382,N_19776,N_18439);
nand U24383 (N_24383,N_19539,N_19207);
or U24384 (N_24384,N_16404,N_18473);
and U24385 (N_24385,N_17647,N_19994);
and U24386 (N_24386,N_18042,N_16457);
nand U24387 (N_24387,N_19643,N_19488);
xnor U24388 (N_24388,N_19576,N_15808);
nand U24389 (N_24389,N_18284,N_17783);
or U24390 (N_24390,N_17723,N_19906);
and U24391 (N_24391,N_15312,N_17315);
nand U24392 (N_24392,N_16361,N_19996);
xor U24393 (N_24393,N_18093,N_19781);
nor U24394 (N_24394,N_16777,N_15685);
xor U24395 (N_24395,N_16966,N_18864);
or U24396 (N_24396,N_18748,N_18145);
xor U24397 (N_24397,N_15863,N_18685);
and U24398 (N_24398,N_18780,N_15025);
xnor U24399 (N_24399,N_16017,N_15475);
or U24400 (N_24400,N_18436,N_15967);
xnor U24401 (N_24401,N_16702,N_17883);
and U24402 (N_24402,N_19265,N_15108);
or U24403 (N_24403,N_16292,N_19143);
nor U24404 (N_24404,N_19582,N_16992);
nor U24405 (N_24405,N_18158,N_19239);
xor U24406 (N_24406,N_17761,N_15530);
nand U24407 (N_24407,N_16049,N_15016);
and U24408 (N_24408,N_15260,N_15038);
or U24409 (N_24409,N_18224,N_19157);
and U24410 (N_24410,N_16567,N_18876);
or U24411 (N_24411,N_15363,N_18016);
nand U24412 (N_24412,N_15568,N_16056);
nor U24413 (N_24413,N_17368,N_18756);
nand U24414 (N_24414,N_16817,N_15875);
nor U24415 (N_24415,N_15403,N_18114);
nor U24416 (N_24416,N_16107,N_18007);
nor U24417 (N_24417,N_18997,N_16451);
or U24418 (N_24418,N_18575,N_18074);
nand U24419 (N_24419,N_18989,N_18633);
xnor U24420 (N_24420,N_17978,N_15005);
or U24421 (N_24421,N_15115,N_16402);
nand U24422 (N_24422,N_15278,N_16253);
xor U24423 (N_24423,N_17586,N_17788);
nand U24424 (N_24424,N_18072,N_18747);
or U24425 (N_24425,N_16811,N_19152);
xor U24426 (N_24426,N_17131,N_19583);
xor U24427 (N_24427,N_19337,N_18170);
nor U24428 (N_24428,N_19548,N_18612);
or U24429 (N_24429,N_15554,N_15234);
nor U24430 (N_24430,N_15302,N_16072);
or U24431 (N_24431,N_19134,N_19293);
and U24432 (N_24432,N_17441,N_17577);
xor U24433 (N_24433,N_17567,N_16453);
or U24434 (N_24434,N_19046,N_17095);
xor U24435 (N_24435,N_16156,N_15126);
and U24436 (N_24436,N_17400,N_18156);
nand U24437 (N_24437,N_19315,N_19844);
and U24438 (N_24438,N_18587,N_16542);
and U24439 (N_24439,N_19699,N_16669);
nand U24440 (N_24440,N_16387,N_16677);
nor U24441 (N_24441,N_19306,N_17652);
nand U24442 (N_24442,N_18348,N_17731);
and U24443 (N_24443,N_18819,N_18821);
nor U24444 (N_24444,N_15978,N_18197);
and U24445 (N_24445,N_16768,N_16042);
nand U24446 (N_24446,N_18247,N_16660);
nand U24447 (N_24447,N_15945,N_18293);
nor U24448 (N_24448,N_16485,N_19926);
and U24449 (N_24449,N_15745,N_15336);
and U24450 (N_24450,N_15078,N_18821);
or U24451 (N_24451,N_15416,N_19362);
xnor U24452 (N_24452,N_18519,N_19985);
nor U24453 (N_24453,N_16051,N_16046);
and U24454 (N_24454,N_18703,N_19636);
nor U24455 (N_24455,N_16514,N_17019);
nor U24456 (N_24456,N_17537,N_15798);
nor U24457 (N_24457,N_18287,N_18933);
or U24458 (N_24458,N_15579,N_15398);
or U24459 (N_24459,N_16295,N_15456);
xor U24460 (N_24460,N_15664,N_18722);
nor U24461 (N_24461,N_17858,N_15778);
xor U24462 (N_24462,N_18273,N_18139);
or U24463 (N_24463,N_18911,N_18747);
nand U24464 (N_24464,N_16850,N_15767);
and U24465 (N_24465,N_18492,N_19671);
and U24466 (N_24466,N_17512,N_19407);
or U24467 (N_24467,N_18766,N_15400);
xnor U24468 (N_24468,N_18422,N_15153);
or U24469 (N_24469,N_17335,N_16245);
nand U24470 (N_24470,N_18670,N_15328);
nor U24471 (N_24471,N_17586,N_16070);
nand U24472 (N_24472,N_17593,N_19958);
xor U24473 (N_24473,N_16897,N_17247);
and U24474 (N_24474,N_15681,N_19615);
and U24475 (N_24475,N_18832,N_16775);
nor U24476 (N_24476,N_16280,N_19701);
nor U24477 (N_24477,N_18311,N_17519);
xnor U24478 (N_24478,N_18516,N_15224);
nor U24479 (N_24479,N_15821,N_17656);
nor U24480 (N_24480,N_17879,N_18743);
or U24481 (N_24481,N_15024,N_18161);
nor U24482 (N_24482,N_19532,N_15796);
or U24483 (N_24483,N_18159,N_19398);
or U24484 (N_24484,N_18694,N_16835);
and U24485 (N_24485,N_15422,N_19325);
nand U24486 (N_24486,N_18891,N_17727);
or U24487 (N_24487,N_19054,N_15516);
nor U24488 (N_24488,N_17612,N_19812);
nor U24489 (N_24489,N_15918,N_18856);
nand U24490 (N_24490,N_16307,N_17376);
or U24491 (N_24491,N_18480,N_18854);
nand U24492 (N_24492,N_15819,N_17988);
or U24493 (N_24493,N_16687,N_16396);
or U24494 (N_24494,N_16183,N_19000);
and U24495 (N_24495,N_15648,N_19518);
or U24496 (N_24496,N_18217,N_17852);
nor U24497 (N_24497,N_15232,N_18826);
nand U24498 (N_24498,N_16639,N_17476);
xor U24499 (N_24499,N_19486,N_15153);
nor U24500 (N_24500,N_18531,N_19209);
nor U24501 (N_24501,N_19394,N_16146);
nand U24502 (N_24502,N_16793,N_17483);
and U24503 (N_24503,N_16233,N_18806);
xnor U24504 (N_24504,N_19467,N_16721);
xnor U24505 (N_24505,N_19247,N_18614);
and U24506 (N_24506,N_19863,N_18014);
and U24507 (N_24507,N_18646,N_18386);
xor U24508 (N_24508,N_16505,N_16584);
nand U24509 (N_24509,N_18454,N_16988);
or U24510 (N_24510,N_17175,N_16527);
and U24511 (N_24511,N_17978,N_18537);
and U24512 (N_24512,N_19146,N_18815);
or U24513 (N_24513,N_15620,N_15640);
or U24514 (N_24514,N_15582,N_16881);
or U24515 (N_24515,N_16723,N_18819);
or U24516 (N_24516,N_18549,N_18231);
or U24517 (N_24517,N_17833,N_15976);
or U24518 (N_24518,N_17166,N_19335);
or U24519 (N_24519,N_15350,N_18908);
or U24520 (N_24520,N_15840,N_15069);
xor U24521 (N_24521,N_18852,N_16131);
and U24522 (N_24522,N_16241,N_18165);
xnor U24523 (N_24523,N_17072,N_17414);
xnor U24524 (N_24524,N_17386,N_16028);
and U24525 (N_24525,N_15387,N_15152);
nand U24526 (N_24526,N_17065,N_18998);
nor U24527 (N_24527,N_17108,N_19650);
or U24528 (N_24528,N_16638,N_19914);
nand U24529 (N_24529,N_15163,N_15885);
and U24530 (N_24530,N_16845,N_19243);
and U24531 (N_24531,N_19115,N_18053);
xor U24532 (N_24532,N_19844,N_15635);
and U24533 (N_24533,N_18100,N_17702);
xor U24534 (N_24534,N_15344,N_19889);
nand U24535 (N_24535,N_15605,N_16212);
xor U24536 (N_24536,N_16841,N_19263);
and U24537 (N_24537,N_17501,N_18528);
xor U24538 (N_24538,N_16061,N_15981);
or U24539 (N_24539,N_16581,N_15248);
nand U24540 (N_24540,N_19735,N_15721);
nand U24541 (N_24541,N_16160,N_18052);
or U24542 (N_24542,N_18521,N_18877);
nand U24543 (N_24543,N_19643,N_18574);
xnor U24544 (N_24544,N_19324,N_15743);
xnor U24545 (N_24545,N_15389,N_17094);
nor U24546 (N_24546,N_17915,N_15920);
nor U24547 (N_24547,N_17695,N_17991);
xnor U24548 (N_24548,N_17615,N_18909);
nor U24549 (N_24549,N_17468,N_16753);
or U24550 (N_24550,N_19815,N_17027);
or U24551 (N_24551,N_19520,N_15204);
and U24552 (N_24552,N_19992,N_18023);
nand U24553 (N_24553,N_17018,N_15699);
or U24554 (N_24554,N_16480,N_17603);
nor U24555 (N_24555,N_18906,N_19709);
xnor U24556 (N_24556,N_17274,N_16882);
or U24557 (N_24557,N_19703,N_18833);
nor U24558 (N_24558,N_19987,N_15069);
and U24559 (N_24559,N_19771,N_17906);
or U24560 (N_24560,N_18122,N_17649);
nor U24561 (N_24561,N_18366,N_16681);
or U24562 (N_24562,N_17311,N_15917);
nor U24563 (N_24563,N_19087,N_17662);
or U24564 (N_24564,N_15626,N_16438);
or U24565 (N_24565,N_17989,N_18432);
or U24566 (N_24566,N_16081,N_19812);
or U24567 (N_24567,N_15932,N_16502);
and U24568 (N_24568,N_16782,N_16397);
xnor U24569 (N_24569,N_19868,N_19242);
nor U24570 (N_24570,N_18901,N_16799);
xor U24571 (N_24571,N_18046,N_18137);
or U24572 (N_24572,N_15134,N_18210);
nor U24573 (N_24573,N_19073,N_16071);
xor U24574 (N_24574,N_16266,N_18243);
nand U24575 (N_24575,N_16146,N_16077);
xor U24576 (N_24576,N_15482,N_17015);
and U24577 (N_24577,N_18926,N_19928);
nor U24578 (N_24578,N_18882,N_17561);
nor U24579 (N_24579,N_15598,N_15167);
nand U24580 (N_24580,N_19292,N_16410);
or U24581 (N_24581,N_15788,N_16187);
nor U24582 (N_24582,N_15930,N_18801);
xor U24583 (N_24583,N_17066,N_16680);
nor U24584 (N_24584,N_17042,N_19174);
xor U24585 (N_24585,N_15897,N_16840);
and U24586 (N_24586,N_19270,N_19838);
and U24587 (N_24587,N_18229,N_16248);
xnor U24588 (N_24588,N_16932,N_17468);
or U24589 (N_24589,N_16830,N_17261);
and U24590 (N_24590,N_19640,N_16537);
or U24591 (N_24591,N_18203,N_19794);
and U24592 (N_24592,N_15732,N_19663);
nor U24593 (N_24593,N_18977,N_18329);
nor U24594 (N_24594,N_16943,N_17958);
nand U24595 (N_24595,N_16698,N_17653);
or U24596 (N_24596,N_19947,N_19856);
nand U24597 (N_24597,N_18397,N_16325);
nand U24598 (N_24598,N_15148,N_16034);
and U24599 (N_24599,N_19442,N_18823);
xor U24600 (N_24600,N_16381,N_19829);
and U24601 (N_24601,N_19003,N_16283);
nor U24602 (N_24602,N_18908,N_19845);
nor U24603 (N_24603,N_15186,N_18228);
and U24604 (N_24604,N_15230,N_15283);
and U24605 (N_24605,N_18232,N_17125);
nor U24606 (N_24606,N_15162,N_19224);
xnor U24607 (N_24607,N_15630,N_17521);
nor U24608 (N_24608,N_15226,N_17215);
or U24609 (N_24609,N_17351,N_15732);
nand U24610 (N_24610,N_19182,N_19829);
xnor U24611 (N_24611,N_17008,N_16173);
and U24612 (N_24612,N_15289,N_15327);
and U24613 (N_24613,N_19682,N_19480);
and U24614 (N_24614,N_16847,N_18921);
and U24615 (N_24615,N_15319,N_16158);
xor U24616 (N_24616,N_19514,N_18720);
nor U24617 (N_24617,N_19699,N_19045);
or U24618 (N_24618,N_18031,N_18146);
nor U24619 (N_24619,N_17392,N_15182);
nor U24620 (N_24620,N_18288,N_16232);
nor U24621 (N_24621,N_16104,N_15454);
xnor U24622 (N_24622,N_18911,N_17958);
nand U24623 (N_24623,N_19968,N_15646);
or U24624 (N_24624,N_17276,N_16070);
or U24625 (N_24625,N_18286,N_17397);
nand U24626 (N_24626,N_16862,N_15272);
nor U24627 (N_24627,N_19146,N_17240);
nor U24628 (N_24628,N_16264,N_17314);
xor U24629 (N_24629,N_15743,N_16493);
nor U24630 (N_24630,N_16188,N_15183);
nor U24631 (N_24631,N_18476,N_17952);
or U24632 (N_24632,N_16500,N_16201);
or U24633 (N_24633,N_15340,N_15706);
nor U24634 (N_24634,N_18476,N_16917);
xnor U24635 (N_24635,N_18788,N_18355);
nand U24636 (N_24636,N_19080,N_15271);
and U24637 (N_24637,N_16535,N_17815);
and U24638 (N_24638,N_17893,N_16054);
nand U24639 (N_24639,N_17453,N_19643);
or U24640 (N_24640,N_17695,N_18398);
xnor U24641 (N_24641,N_16006,N_16812);
xor U24642 (N_24642,N_19108,N_19786);
nor U24643 (N_24643,N_15242,N_17755);
nand U24644 (N_24644,N_18305,N_15476);
and U24645 (N_24645,N_19099,N_17169);
or U24646 (N_24646,N_19254,N_19340);
nand U24647 (N_24647,N_15661,N_17806);
xor U24648 (N_24648,N_17281,N_16173);
nor U24649 (N_24649,N_17027,N_15339);
or U24650 (N_24650,N_19172,N_19298);
and U24651 (N_24651,N_19188,N_18805);
or U24652 (N_24652,N_16384,N_18869);
xnor U24653 (N_24653,N_16680,N_15766);
and U24654 (N_24654,N_18885,N_16350);
xnor U24655 (N_24655,N_19065,N_16157);
nand U24656 (N_24656,N_17411,N_16854);
nand U24657 (N_24657,N_15847,N_16211);
nor U24658 (N_24658,N_19780,N_15571);
nand U24659 (N_24659,N_18143,N_17653);
or U24660 (N_24660,N_16237,N_15904);
or U24661 (N_24661,N_19708,N_18043);
nor U24662 (N_24662,N_18115,N_19129);
or U24663 (N_24663,N_19923,N_15418);
or U24664 (N_24664,N_17301,N_17089);
xor U24665 (N_24665,N_17931,N_16773);
xor U24666 (N_24666,N_19445,N_19560);
nor U24667 (N_24667,N_17043,N_19650);
nand U24668 (N_24668,N_19331,N_19894);
or U24669 (N_24669,N_18342,N_19350);
and U24670 (N_24670,N_15003,N_17354);
nor U24671 (N_24671,N_17689,N_16149);
or U24672 (N_24672,N_15937,N_15004);
nor U24673 (N_24673,N_16857,N_15058);
nor U24674 (N_24674,N_17067,N_16090);
nand U24675 (N_24675,N_19573,N_15785);
nand U24676 (N_24676,N_15600,N_18061);
or U24677 (N_24677,N_17820,N_19884);
nand U24678 (N_24678,N_15151,N_19847);
xor U24679 (N_24679,N_19878,N_18175);
or U24680 (N_24680,N_19499,N_16424);
or U24681 (N_24681,N_17222,N_15133);
nor U24682 (N_24682,N_18821,N_17181);
nor U24683 (N_24683,N_18193,N_19209);
xor U24684 (N_24684,N_15579,N_18265);
nor U24685 (N_24685,N_15837,N_19555);
xnor U24686 (N_24686,N_16869,N_18861);
or U24687 (N_24687,N_16885,N_17200);
and U24688 (N_24688,N_18648,N_15164);
and U24689 (N_24689,N_17163,N_15477);
xor U24690 (N_24690,N_17905,N_16838);
and U24691 (N_24691,N_15546,N_18184);
and U24692 (N_24692,N_18339,N_17536);
and U24693 (N_24693,N_19494,N_18290);
nor U24694 (N_24694,N_18441,N_19333);
xnor U24695 (N_24695,N_18403,N_17940);
or U24696 (N_24696,N_15403,N_19885);
and U24697 (N_24697,N_17282,N_15253);
xnor U24698 (N_24698,N_18512,N_17282);
and U24699 (N_24699,N_16489,N_16447);
or U24700 (N_24700,N_17545,N_15815);
nor U24701 (N_24701,N_19908,N_16626);
and U24702 (N_24702,N_18319,N_18289);
and U24703 (N_24703,N_15469,N_18244);
xor U24704 (N_24704,N_15772,N_15698);
xnor U24705 (N_24705,N_15430,N_16334);
nor U24706 (N_24706,N_16226,N_18173);
or U24707 (N_24707,N_17856,N_19334);
and U24708 (N_24708,N_17869,N_15688);
nor U24709 (N_24709,N_16451,N_19785);
and U24710 (N_24710,N_19028,N_17438);
nor U24711 (N_24711,N_17769,N_16445);
and U24712 (N_24712,N_15079,N_18228);
xor U24713 (N_24713,N_16504,N_16013);
xnor U24714 (N_24714,N_15367,N_16090);
xnor U24715 (N_24715,N_18456,N_19921);
xnor U24716 (N_24716,N_19345,N_19608);
or U24717 (N_24717,N_16583,N_16300);
nor U24718 (N_24718,N_15035,N_18463);
or U24719 (N_24719,N_19782,N_19450);
or U24720 (N_24720,N_18399,N_19209);
nor U24721 (N_24721,N_17936,N_18143);
xnor U24722 (N_24722,N_15541,N_19001);
nor U24723 (N_24723,N_18475,N_18196);
and U24724 (N_24724,N_19421,N_15967);
nor U24725 (N_24725,N_16291,N_16279);
nor U24726 (N_24726,N_16909,N_17919);
and U24727 (N_24727,N_17271,N_17867);
and U24728 (N_24728,N_19060,N_18033);
or U24729 (N_24729,N_19244,N_16790);
or U24730 (N_24730,N_15872,N_15505);
xor U24731 (N_24731,N_15236,N_16450);
and U24732 (N_24732,N_16335,N_19800);
xor U24733 (N_24733,N_16198,N_18176);
nor U24734 (N_24734,N_18952,N_19554);
nand U24735 (N_24735,N_17554,N_18581);
nor U24736 (N_24736,N_16758,N_18952);
xor U24737 (N_24737,N_17399,N_17836);
nand U24738 (N_24738,N_18285,N_15681);
and U24739 (N_24739,N_19496,N_16772);
nor U24740 (N_24740,N_18585,N_18096);
nand U24741 (N_24741,N_17418,N_15187);
nor U24742 (N_24742,N_15036,N_19526);
nand U24743 (N_24743,N_18382,N_18150);
nor U24744 (N_24744,N_17345,N_18063);
and U24745 (N_24745,N_16188,N_18026);
or U24746 (N_24746,N_15809,N_19700);
nand U24747 (N_24747,N_19211,N_15316);
and U24748 (N_24748,N_16013,N_15141);
xor U24749 (N_24749,N_16610,N_16662);
xnor U24750 (N_24750,N_19134,N_16350);
nand U24751 (N_24751,N_18261,N_17819);
or U24752 (N_24752,N_16008,N_15875);
xnor U24753 (N_24753,N_15252,N_16535);
or U24754 (N_24754,N_19499,N_15455);
or U24755 (N_24755,N_15641,N_17282);
and U24756 (N_24756,N_19464,N_15277);
and U24757 (N_24757,N_18611,N_19518);
nand U24758 (N_24758,N_17664,N_18050);
and U24759 (N_24759,N_15928,N_19392);
nand U24760 (N_24760,N_18991,N_15130);
nand U24761 (N_24761,N_15351,N_19286);
and U24762 (N_24762,N_18938,N_17204);
and U24763 (N_24763,N_17548,N_18248);
nor U24764 (N_24764,N_15621,N_19696);
and U24765 (N_24765,N_19153,N_18050);
and U24766 (N_24766,N_16663,N_17753);
nor U24767 (N_24767,N_18171,N_18708);
nor U24768 (N_24768,N_15072,N_18750);
nand U24769 (N_24769,N_15750,N_17630);
nand U24770 (N_24770,N_16734,N_17885);
or U24771 (N_24771,N_15605,N_15149);
nor U24772 (N_24772,N_18614,N_17880);
or U24773 (N_24773,N_16127,N_16890);
nand U24774 (N_24774,N_18020,N_18801);
nor U24775 (N_24775,N_16814,N_17622);
xnor U24776 (N_24776,N_17754,N_17933);
or U24777 (N_24777,N_15457,N_15308);
and U24778 (N_24778,N_16906,N_18381);
xnor U24779 (N_24779,N_17100,N_15047);
and U24780 (N_24780,N_19504,N_18609);
nor U24781 (N_24781,N_18558,N_15909);
xnor U24782 (N_24782,N_18408,N_17260);
and U24783 (N_24783,N_15490,N_15884);
nor U24784 (N_24784,N_17231,N_15068);
nor U24785 (N_24785,N_15400,N_16072);
xnor U24786 (N_24786,N_15088,N_17830);
and U24787 (N_24787,N_15312,N_18250);
xnor U24788 (N_24788,N_17232,N_17844);
xor U24789 (N_24789,N_19020,N_18574);
and U24790 (N_24790,N_19141,N_15054);
xor U24791 (N_24791,N_18221,N_18296);
and U24792 (N_24792,N_18513,N_16712);
nand U24793 (N_24793,N_19863,N_18676);
or U24794 (N_24794,N_16733,N_18606);
xnor U24795 (N_24795,N_19251,N_15815);
or U24796 (N_24796,N_17820,N_18868);
nor U24797 (N_24797,N_18897,N_15116);
or U24798 (N_24798,N_16667,N_18653);
nor U24799 (N_24799,N_18794,N_16999);
nor U24800 (N_24800,N_19453,N_19193);
nand U24801 (N_24801,N_15553,N_15197);
or U24802 (N_24802,N_17467,N_15711);
and U24803 (N_24803,N_18457,N_18024);
or U24804 (N_24804,N_19657,N_16678);
and U24805 (N_24805,N_15726,N_15796);
or U24806 (N_24806,N_18481,N_18075);
or U24807 (N_24807,N_19084,N_19927);
or U24808 (N_24808,N_17698,N_15735);
and U24809 (N_24809,N_19039,N_18363);
nor U24810 (N_24810,N_19257,N_18305);
nand U24811 (N_24811,N_15244,N_17691);
nand U24812 (N_24812,N_19588,N_19079);
or U24813 (N_24813,N_16664,N_19300);
xnor U24814 (N_24814,N_17312,N_15525);
or U24815 (N_24815,N_15630,N_18248);
xnor U24816 (N_24816,N_16312,N_17307);
or U24817 (N_24817,N_15904,N_19396);
or U24818 (N_24818,N_16264,N_18555);
and U24819 (N_24819,N_15800,N_19710);
xnor U24820 (N_24820,N_15149,N_15055);
or U24821 (N_24821,N_16570,N_19633);
and U24822 (N_24822,N_16514,N_15777);
and U24823 (N_24823,N_18121,N_19765);
and U24824 (N_24824,N_17333,N_17157);
or U24825 (N_24825,N_17531,N_18698);
or U24826 (N_24826,N_17349,N_19074);
nor U24827 (N_24827,N_15715,N_18917);
or U24828 (N_24828,N_17792,N_18804);
xnor U24829 (N_24829,N_19063,N_15624);
nor U24830 (N_24830,N_15270,N_19982);
or U24831 (N_24831,N_19081,N_18034);
xor U24832 (N_24832,N_18145,N_16294);
nor U24833 (N_24833,N_15287,N_19926);
xor U24834 (N_24834,N_18808,N_18124);
nand U24835 (N_24835,N_15575,N_18036);
xor U24836 (N_24836,N_17448,N_15339);
and U24837 (N_24837,N_17891,N_17822);
and U24838 (N_24838,N_15646,N_18955);
or U24839 (N_24839,N_17989,N_17992);
nor U24840 (N_24840,N_19429,N_17466);
nand U24841 (N_24841,N_18278,N_16738);
xor U24842 (N_24842,N_15273,N_15848);
nor U24843 (N_24843,N_16084,N_19698);
or U24844 (N_24844,N_19388,N_19178);
nor U24845 (N_24845,N_16777,N_15410);
or U24846 (N_24846,N_19675,N_17515);
nand U24847 (N_24847,N_17256,N_16429);
xnor U24848 (N_24848,N_17088,N_17405);
or U24849 (N_24849,N_17951,N_15169);
nand U24850 (N_24850,N_18742,N_17451);
xor U24851 (N_24851,N_16845,N_15567);
and U24852 (N_24852,N_19210,N_19079);
xnor U24853 (N_24853,N_16946,N_19128);
and U24854 (N_24854,N_15071,N_16402);
or U24855 (N_24855,N_18731,N_16269);
nor U24856 (N_24856,N_17193,N_19113);
xnor U24857 (N_24857,N_18798,N_16507);
nand U24858 (N_24858,N_15352,N_17649);
nand U24859 (N_24859,N_16239,N_16219);
nand U24860 (N_24860,N_18591,N_17053);
xor U24861 (N_24861,N_17721,N_15836);
or U24862 (N_24862,N_16748,N_17832);
or U24863 (N_24863,N_15419,N_15318);
or U24864 (N_24864,N_19821,N_19100);
or U24865 (N_24865,N_19067,N_19486);
and U24866 (N_24866,N_17366,N_17519);
xor U24867 (N_24867,N_15995,N_18826);
or U24868 (N_24868,N_15918,N_16144);
nand U24869 (N_24869,N_18566,N_17077);
xor U24870 (N_24870,N_19052,N_18641);
xnor U24871 (N_24871,N_17272,N_17424);
xnor U24872 (N_24872,N_15464,N_18337);
xnor U24873 (N_24873,N_19174,N_15000);
nor U24874 (N_24874,N_15999,N_16998);
nor U24875 (N_24875,N_16270,N_18975);
nand U24876 (N_24876,N_17495,N_15475);
or U24877 (N_24877,N_18495,N_18485);
or U24878 (N_24878,N_16739,N_15238);
nand U24879 (N_24879,N_19230,N_15596);
nor U24880 (N_24880,N_18782,N_17463);
xor U24881 (N_24881,N_19188,N_18783);
nand U24882 (N_24882,N_19713,N_15452);
nand U24883 (N_24883,N_17128,N_18630);
and U24884 (N_24884,N_18268,N_15580);
or U24885 (N_24885,N_17534,N_16635);
xor U24886 (N_24886,N_17508,N_19746);
or U24887 (N_24887,N_16060,N_18400);
or U24888 (N_24888,N_19646,N_19569);
xnor U24889 (N_24889,N_16366,N_18967);
xor U24890 (N_24890,N_18103,N_19648);
nand U24891 (N_24891,N_15037,N_17017);
nor U24892 (N_24892,N_15640,N_16442);
or U24893 (N_24893,N_15084,N_19775);
or U24894 (N_24894,N_19548,N_17919);
nor U24895 (N_24895,N_16872,N_19134);
or U24896 (N_24896,N_15204,N_17702);
nor U24897 (N_24897,N_17452,N_17510);
and U24898 (N_24898,N_16604,N_15533);
nand U24899 (N_24899,N_16104,N_18245);
nor U24900 (N_24900,N_19041,N_19619);
xnor U24901 (N_24901,N_19872,N_19102);
xor U24902 (N_24902,N_16446,N_17731);
nand U24903 (N_24903,N_15141,N_16864);
or U24904 (N_24904,N_17387,N_19040);
and U24905 (N_24905,N_16233,N_18722);
and U24906 (N_24906,N_18518,N_16729);
nor U24907 (N_24907,N_16230,N_15538);
or U24908 (N_24908,N_15310,N_18064);
nor U24909 (N_24909,N_19544,N_16674);
and U24910 (N_24910,N_17639,N_15548);
nor U24911 (N_24911,N_15124,N_16527);
nand U24912 (N_24912,N_16914,N_19104);
xnor U24913 (N_24913,N_15913,N_15184);
or U24914 (N_24914,N_16183,N_16927);
xor U24915 (N_24915,N_16375,N_19097);
xor U24916 (N_24916,N_16919,N_16808);
xnor U24917 (N_24917,N_17042,N_15753);
nor U24918 (N_24918,N_15646,N_18191);
nor U24919 (N_24919,N_17745,N_15059);
nand U24920 (N_24920,N_18463,N_18249);
xor U24921 (N_24921,N_17187,N_18558);
and U24922 (N_24922,N_17846,N_16316);
and U24923 (N_24923,N_19700,N_17887);
or U24924 (N_24924,N_18950,N_18110);
nor U24925 (N_24925,N_15481,N_18660);
nand U24926 (N_24926,N_16599,N_19577);
or U24927 (N_24927,N_16420,N_18377);
or U24928 (N_24928,N_17408,N_15615);
nor U24929 (N_24929,N_16427,N_16857);
xor U24930 (N_24930,N_17469,N_17065);
nor U24931 (N_24931,N_19411,N_18370);
nand U24932 (N_24932,N_16756,N_19187);
and U24933 (N_24933,N_17383,N_16083);
and U24934 (N_24934,N_15226,N_15707);
xnor U24935 (N_24935,N_15830,N_18793);
nor U24936 (N_24936,N_16241,N_19720);
or U24937 (N_24937,N_17452,N_17616);
nand U24938 (N_24938,N_15007,N_17622);
nand U24939 (N_24939,N_18141,N_17593);
xor U24940 (N_24940,N_18804,N_16186);
or U24941 (N_24941,N_16441,N_15380);
and U24942 (N_24942,N_16887,N_18152);
xor U24943 (N_24943,N_18037,N_19788);
nand U24944 (N_24944,N_15043,N_18934);
nor U24945 (N_24945,N_19991,N_19320);
and U24946 (N_24946,N_16303,N_19712);
and U24947 (N_24947,N_15546,N_16455);
nand U24948 (N_24948,N_18922,N_18419);
or U24949 (N_24949,N_16214,N_19001);
and U24950 (N_24950,N_17616,N_18181);
nand U24951 (N_24951,N_15632,N_15454);
nand U24952 (N_24952,N_18281,N_16411);
or U24953 (N_24953,N_17396,N_18332);
nor U24954 (N_24954,N_15036,N_19352);
xor U24955 (N_24955,N_15370,N_18626);
nor U24956 (N_24956,N_16885,N_17312);
nor U24957 (N_24957,N_16583,N_16910);
xor U24958 (N_24958,N_17122,N_19389);
nor U24959 (N_24959,N_15604,N_17930);
or U24960 (N_24960,N_16634,N_15408);
or U24961 (N_24961,N_15228,N_16507);
nand U24962 (N_24962,N_15939,N_15674);
and U24963 (N_24963,N_17927,N_16520);
xor U24964 (N_24964,N_19364,N_19045);
xnor U24965 (N_24965,N_16031,N_18694);
or U24966 (N_24966,N_18681,N_16499);
nand U24967 (N_24967,N_17980,N_15888);
nor U24968 (N_24968,N_19329,N_18746);
or U24969 (N_24969,N_16197,N_15363);
and U24970 (N_24970,N_16776,N_17262);
nand U24971 (N_24971,N_17597,N_17400);
and U24972 (N_24972,N_16072,N_19276);
or U24973 (N_24973,N_18962,N_19747);
nand U24974 (N_24974,N_19048,N_19393);
and U24975 (N_24975,N_18497,N_17417);
or U24976 (N_24976,N_19729,N_17893);
nand U24977 (N_24977,N_19550,N_17465);
nand U24978 (N_24978,N_18763,N_17399);
nand U24979 (N_24979,N_15861,N_16141);
or U24980 (N_24980,N_16864,N_17400);
or U24981 (N_24981,N_19125,N_18106);
or U24982 (N_24982,N_16785,N_19756);
and U24983 (N_24983,N_19254,N_16919);
or U24984 (N_24984,N_17509,N_17864);
or U24985 (N_24985,N_16096,N_17572);
and U24986 (N_24986,N_16706,N_18974);
nor U24987 (N_24987,N_19020,N_19963);
nor U24988 (N_24988,N_19635,N_18388);
nand U24989 (N_24989,N_16912,N_18905);
and U24990 (N_24990,N_19435,N_18356);
xnor U24991 (N_24991,N_18005,N_16702);
xor U24992 (N_24992,N_17789,N_15327);
and U24993 (N_24993,N_17920,N_18035);
nand U24994 (N_24994,N_16384,N_16329);
nand U24995 (N_24995,N_16340,N_15630);
nor U24996 (N_24996,N_18596,N_16777);
nor U24997 (N_24997,N_17132,N_18727);
and U24998 (N_24998,N_19743,N_16949);
nor U24999 (N_24999,N_15973,N_16896);
and U25000 (N_25000,N_21648,N_24902);
and U25001 (N_25001,N_21519,N_24452);
nor U25002 (N_25002,N_23420,N_22315);
nor U25003 (N_25003,N_23429,N_20348);
or U25004 (N_25004,N_23956,N_24504);
nor U25005 (N_25005,N_22039,N_22966);
or U25006 (N_25006,N_23725,N_22437);
nand U25007 (N_25007,N_24953,N_20631);
or U25008 (N_25008,N_23339,N_23716);
nor U25009 (N_25009,N_21255,N_22662);
and U25010 (N_25010,N_23142,N_20810);
nand U25011 (N_25011,N_22059,N_23744);
xor U25012 (N_25012,N_22730,N_24270);
or U25013 (N_25013,N_24245,N_22097);
nor U25014 (N_25014,N_20304,N_21957);
and U25015 (N_25015,N_20727,N_22484);
nor U25016 (N_25016,N_22477,N_21724);
and U25017 (N_25017,N_21671,N_21542);
nand U25018 (N_25018,N_24392,N_22717);
or U25019 (N_25019,N_22664,N_22850);
or U25020 (N_25020,N_21545,N_24974);
xnor U25021 (N_25021,N_21295,N_23895);
nand U25022 (N_25022,N_22405,N_24622);
nand U25023 (N_25023,N_20831,N_24123);
or U25024 (N_25024,N_24237,N_22231);
nor U25025 (N_25025,N_22519,N_21514);
and U25026 (N_25026,N_24439,N_21689);
nand U25027 (N_25027,N_21763,N_22585);
or U25028 (N_25028,N_22323,N_20660);
or U25029 (N_25029,N_20201,N_22109);
nor U25030 (N_25030,N_24859,N_24285);
and U25031 (N_25031,N_21057,N_22541);
nand U25032 (N_25032,N_21361,N_22240);
and U25033 (N_25033,N_23731,N_22598);
nand U25034 (N_25034,N_24102,N_20040);
xor U25035 (N_25035,N_22351,N_21024);
and U25036 (N_25036,N_23506,N_21793);
nor U25037 (N_25037,N_21081,N_21868);
nor U25038 (N_25038,N_21014,N_21201);
nor U25039 (N_25039,N_20123,N_23759);
nand U25040 (N_25040,N_22821,N_22225);
nor U25041 (N_25041,N_24627,N_20490);
nor U25042 (N_25042,N_21573,N_20644);
and U25043 (N_25043,N_21936,N_21235);
nor U25044 (N_25044,N_23553,N_21281);
nor U25045 (N_25045,N_21430,N_20986);
xor U25046 (N_25046,N_23213,N_21277);
or U25047 (N_25047,N_21954,N_23319);
xor U25048 (N_25048,N_24070,N_22700);
xnor U25049 (N_25049,N_20022,N_24604);
xor U25050 (N_25050,N_20371,N_20495);
nor U25051 (N_25051,N_20238,N_20415);
xnor U25052 (N_25052,N_20436,N_23712);
xor U25053 (N_25053,N_24143,N_21878);
and U25054 (N_25054,N_22168,N_20989);
nor U25055 (N_25055,N_23289,N_24309);
nand U25056 (N_25056,N_24053,N_24794);
or U25057 (N_25057,N_22252,N_22822);
and U25058 (N_25058,N_21170,N_23826);
nand U25059 (N_25059,N_20517,N_20536);
xor U25060 (N_25060,N_21016,N_24922);
nor U25061 (N_25061,N_21717,N_20772);
nor U25062 (N_25062,N_24958,N_20577);
xor U25063 (N_25063,N_20394,N_20894);
xor U25064 (N_25064,N_21259,N_24126);
nand U25065 (N_25065,N_20560,N_24684);
xnor U25066 (N_25066,N_21258,N_21985);
and U25067 (N_25067,N_23926,N_20332);
nor U25068 (N_25068,N_24323,N_23059);
and U25069 (N_25069,N_22755,N_23878);
or U25070 (N_25070,N_22615,N_24629);
nor U25071 (N_25071,N_22415,N_24857);
and U25072 (N_25072,N_21529,N_23735);
nor U25073 (N_25073,N_24592,N_22212);
xor U25074 (N_25074,N_22741,N_23574);
nor U25075 (N_25075,N_22995,N_21084);
nor U25076 (N_25076,N_24118,N_24286);
nor U25077 (N_25077,N_21756,N_24410);
nor U25078 (N_25078,N_22567,N_23607);
and U25079 (N_25079,N_24432,N_21173);
or U25080 (N_25080,N_22583,N_23804);
and U25081 (N_25081,N_24434,N_24005);
xor U25082 (N_25082,N_23163,N_23002);
and U25083 (N_25083,N_22658,N_21329);
xor U25084 (N_25084,N_24354,N_24775);
xnor U25085 (N_25085,N_24591,N_20964);
and U25086 (N_25086,N_21758,N_22795);
or U25087 (N_25087,N_22434,N_21718);
or U25088 (N_25088,N_21335,N_21458);
nor U25089 (N_25089,N_24056,N_24771);
xnor U25090 (N_25090,N_23853,N_21994);
nor U25091 (N_25091,N_24447,N_22287);
nor U25092 (N_25092,N_20785,N_21433);
xnor U25093 (N_25093,N_23109,N_22262);
and U25094 (N_25094,N_24222,N_20189);
xor U25095 (N_25095,N_23551,N_20512);
nand U25096 (N_25096,N_21002,N_24893);
nand U25097 (N_25097,N_20082,N_22466);
nor U25098 (N_25098,N_20484,N_22106);
and U25099 (N_25099,N_23998,N_23384);
or U25100 (N_25100,N_21674,N_20423);
or U25101 (N_25101,N_22280,N_22306);
xor U25102 (N_25102,N_20655,N_22126);
nor U25103 (N_25103,N_21203,N_23676);
nand U25104 (N_25104,N_20701,N_24666);
nor U25105 (N_25105,N_21309,N_23792);
or U25106 (N_25106,N_20352,N_23388);
or U25107 (N_25107,N_22612,N_22693);
nor U25108 (N_25108,N_24863,N_21455);
xor U25109 (N_25109,N_23577,N_20069);
or U25110 (N_25110,N_24366,N_21585);
xor U25111 (N_25111,N_22659,N_21066);
and U25112 (N_25112,N_21161,N_20883);
nand U25113 (N_25113,N_23819,N_20893);
nand U25114 (N_25114,N_24426,N_22561);
xnor U25115 (N_25115,N_20104,N_21325);
xnor U25116 (N_25116,N_22356,N_20606);
or U25117 (N_25117,N_20830,N_21572);
nand U25118 (N_25118,N_22569,N_23313);
or U25119 (N_25119,N_21218,N_23254);
or U25120 (N_25120,N_20061,N_22878);
nor U25121 (N_25121,N_21918,N_20190);
or U25122 (N_25122,N_22257,N_23406);
xnor U25123 (N_25123,N_22861,N_23994);
xor U25124 (N_25124,N_21979,N_20438);
nor U25125 (N_25125,N_22803,N_22950);
or U25126 (N_25126,N_22925,N_22532);
nand U25127 (N_25127,N_22956,N_23700);
or U25128 (N_25128,N_22364,N_23341);
nor U25129 (N_25129,N_24647,N_21232);
nor U25130 (N_25130,N_22827,N_22191);
nor U25131 (N_25131,N_24746,N_22312);
and U25132 (N_25132,N_24227,N_21986);
nor U25133 (N_25133,N_23809,N_22103);
and U25134 (N_25134,N_23828,N_22762);
nand U25135 (N_25135,N_22326,N_20308);
or U25136 (N_25136,N_21271,N_21209);
nand U25137 (N_25137,N_21677,N_23549);
nor U25138 (N_25138,N_21703,N_24724);
nand U25139 (N_25139,N_21144,N_24177);
nor U25140 (N_25140,N_24188,N_24362);
or U25141 (N_25141,N_23416,N_24568);
nor U25142 (N_25142,N_20728,N_23714);
nor U25143 (N_25143,N_22376,N_23232);
and U25144 (N_25144,N_21822,N_23447);
and U25145 (N_25145,N_22607,N_22119);
nand U25146 (N_25146,N_20945,N_21076);
xnor U25147 (N_25147,N_23252,N_23327);
xnor U25148 (N_25148,N_20668,N_24171);
xor U25149 (N_25149,N_22746,N_20952);
xnor U25150 (N_25150,N_23790,N_22156);
xor U25151 (N_25151,N_24242,N_23207);
or U25152 (N_25152,N_21995,N_22491);
nand U25153 (N_25153,N_23554,N_22147);
xor U25154 (N_25154,N_22165,N_21072);
nand U25155 (N_25155,N_20891,N_23812);
nand U25156 (N_25156,N_23698,N_24534);
nand U25157 (N_25157,N_24569,N_24906);
nor U25158 (N_25158,N_22565,N_23847);
and U25159 (N_25159,N_21090,N_23365);
or U25160 (N_25160,N_23882,N_22898);
or U25161 (N_25161,N_22733,N_21473);
nand U25162 (N_25162,N_20018,N_21095);
and U25163 (N_25163,N_20678,N_20617);
or U25164 (N_25164,N_20155,N_21908);
nor U25165 (N_25165,N_23247,N_21288);
nand U25166 (N_25166,N_21856,N_24764);
nor U25167 (N_25167,N_23413,N_23007);
xor U25168 (N_25168,N_21182,N_23112);
and U25169 (N_25169,N_20912,N_21788);
or U25170 (N_25170,N_22141,N_21842);
xor U25171 (N_25171,N_23322,N_23987);
and U25172 (N_25172,N_23378,N_22518);
or U25173 (N_25173,N_23501,N_20324);
xor U25174 (N_25174,N_24870,N_23872);
nor U25175 (N_25175,N_21527,N_24483);
xor U25176 (N_25176,N_20759,N_20422);
or U25177 (N_25177,N_24643,N_24217);
xor U25178 (N_25178,N_21738,N_24639);
and U25179 (N_25179,N_20089,N_24539);
and U25180 (N_25180,N_21319,N_22043);
or U25181 (N_25181,N_22193,N_23175);
and U25182 (N_25182,N_21278,N_21816);
and U25183 (N_25183,N_21725,N_23911);
nor U25184 (N_25184,N_24869,N_21583);
nand U25185 (N_25185,N_23284,N_23942);
nor U25186 (N_25186,N_21001,N_22457);
nand U25187 (N_25187,N_23898,N_21949);
nor U25188 (N_25188,N_21592,N_24407);
nor U25189 (N_25189,N_21488,N_23131);
or U25190 (N_25190,N_23432,N_22012);
xor U25191 (N_25191,N_24843,N_23904);
nand U25192 (N_25192,N_24801,N_20712);
nand U25193 (N_25193,N_22230,N_24218);
nand U25194 (N_25194,N_20762,N_20683);
and U25195 (N_25195,N_20420,N_24234);
nor U25196 (N_25196,N_20116,N_20081);
or U25197 (N_25197,N_22789,N_22889);
or U25198 (N_25198,N_20113,N_22482);
xor U25199 (N_25199,N_20313,N_23522);
nand U25200 (N_25200,N_20465,N_20887);
and U25201 (N_25201,N_24679,N_22593);
or U25202 (N_25202,N_20710,N_23585);
nand U25203 (N_25203,N_20718,N_24508);
and U25204 (N_25204,N_20847,N_20358);
nand U25205 (N_25205,N_20354,N_20402);
or U25206 (N_25206,N_20890,N_24206);
nor U25207 (N_25207,N_23177,N_20382);
nor U25208 (N_25208,N_21864,N_23859);
nand U25209 (N_25209,N_21600,N_21041);
xor U25210 (N_25210,N_21409,N_21304);
and U25211 (N_25211,N_24336,N_20130);
and U25212 (N_25212,N_21528,N_20350);
nand U25213 (N_25213,N_21417,N_22723);
nor U25214 (N_25214,N_20799,N_24311);
nand U25215 (N_25215,N_24581,N_21781);
xnor U25216 (N_25216,N_24704,N_24946);
or U25217 (N_25217,N_24661,N_24635);
xor U25218 (N_25218,N_22148,N_23866);
xnor U25219 (N_25219,N_24251,N_21681);
xor U25220 (N_25220,N_24589,N_23715);
xor U25221 (N_25221,N_22074,N_24474);
nand U25222 (N_25222,N_24899,N_23139);
and U25223 (N_25223,N_21422,N_21300);
nor U25224 (N_25224,N_21485,N_20879);
or U25225 (N_25225,N_22027,N_24238);
nor U25226 (N_25226,N_24229,N_20167);
xor U25227 (N_25227,N_23548,N_20496);
nor U25228 (N_25228,N_23963,N_24887);
xnor U25229 (N_25229,N_23583,N_24945);
nand U25230 (N_25230,N_23644,N_21462);
nor U25231 (N_25231,N_22807,N_24258);
and U25232 (N_25232,N_20291,N_20895);
nor U25233 (N_25233,N_23249,N_21608);
nor U25234 (N_25234,N_22247,N_22279);
and U25235 (N_25235,N_22556,N_22031);
or U25236 (N_25236,N_24396,N_23945);
nor U25237 (N_25237,N_22887,N_21429);
or U25238 (N_25238,N_24798,N_21675);
and U25239 (N_25239,N_24282,N_24928);
nand U25240 (N_25240,N_22464,N_24516);
nand U25241 (N_25241,N_23974,N_20741);
nand U25242 (N_25242,N_20822,N_24040);
xnor U25243 (N_25243,N_24532,N_21865);
nand U25244 (N_25244,N_21713,N_21357);
or U25245 (N_25245,N_21178,N_24740);
xnor U25246 (N_25246,N_23831,N_22638);
and U25247 (N_25247,N_23996,N_21132);
xnor U25248 (N_25248,N_21928,N_24570);
nor U25249 (N_25249,N_22844,N_21607);
and U25250 (N_25250,N_21479,N_22014);
or U25251 (N_25251,N_21780,N_21769);
or U25252 (N_25252,N_24440,N_23734);
nand U25253 (N_25253,N_23949,N_23978);
nor U25254 (N_25254,N_23865,N_23056);
or U25255 (N_25255,N_20501,N_23458);
nand U25256 (N_25256,N_21375,N_24663);
nor U25257 (N_25257,N_21241,N_20576);
nand U25258 (N_25258,N_24788,N_24435);
nand U25259 (N_25259,N_24192,N_23933);
xnor U25260 (N_25260,N_22837,N_23491);
and U25261 (N_25261,N_20109,N_22618);
nand U25262 (N_25262,N_20108,N_24909);
xnor U25263 (N_25263,N_24892,N_24668);
and U25264 (N_25264,N_21204,N_20387);
nor U25265 (N_25265,N_21340,N_24265);
nand U25266 (N_25266,N_20633,N_24828);
or U25267 (N_25267,N_22330,N_22258);
nand U25268 (N_25268,N_22571,N_23685);
and U25269 (N_25269,N_21687,N_21152);
nor U25270 (N_25270,N_20223,N_21639);
nor U25271 (N_25271,N_20930,N_23452);
and U25272 (N_25272,N_23114,N_21852);
and U25273 (N_25273,N_21586,N_22564);
nand U25274 (N_25274,N_22739,N_23478);
nor U25275 (N_25275,N_21405,N_23581);
nor U25276 (N_25276,N_22135,N_21475);
and U25277 (N_25277,N_22524,N_22291);
xnor U25278 (N_25278,N_23884,N_21809);
and U25279 (N_25279,N_23084,N_20634);
nor U25280 (N_25280,N_21881,N_20249);
or U25281 (N_25281,N_20596,N_22910);
xnor U25282 (N_25282,N_23306,N_22336);
or U25283 (N_25283,N_23100,N_24182);
nand U25284 (N_25284,N_20974,N_20296);
and U25285 (N_25285,N_20829,N_24866);
xnor U25286 (N_25286,N_23299,N_24768);
and U25287 (N_25287,N_20447,N_20679);
or U25288 (N_25288,N_23245,N_20997);
and U25289 (N_25289,N_20446,N_20823);
nor U25290 (N_25290,N_23939,N_21169);
and U25291 (N_25291,N_23308,N_20186);
nand U25292 (N_25292,N_24636,N_24505);
or U25293 (N_25293,N_23349,N_22278);
and U25294 (N_25294,N_23879,N_20157);
and U25295 (N_25295,N_21109,N_20571);
nand U25296 (N_25296,N_22830,N_20052);
and U25297 (N_25297,N_24071,N_22293);
and U25298 (N_25298,N_24756,N_24518);
nor U25299 (N_25299,N_23375,N_23855);
or U25300 (N_25300,N_23854,N_20359);
xnor U25301 (N_25301,N_22398,N_20675);
or U25302 (N_25302,N_23758,N_20042);
nor U25303 (N_25303,N_24538,N_21368);
nor U25304 (N_25304,N_22800,N_22187);
nor U25305 (N_25305,N_22796,N_21359);
or U25306 (N_25306,N_20903,N_20601);
and U25307 (N_25307,N_24809,N_24415);
or U25308 (N_25308,N_24064,N_24927);
xor U25309 (N_25309,N_22757,N_20318);
nand U25310 (N_25310,N_21937,N_21990);
nor U25311 (N_25311,N_23612,N_24279);
xnor U25312 (N_25312,N_22938,N_24152);
xnor U25313 (N_25313,N_20551,N_23350);
and U25314 (N_25314,N_23653,N_21287);
nor U25315 (N_25315,N_20714,N_23677);
nor U25316 (N_25316,N_21135,N_23166);
nor U25317 (N_25317,N_24094,N_20479);
and U25318 (N_25318,N_20552,N_23627);
and U25319 (N_25319,N_21722,N_24512);
xor U25320 (N_25320,N_23399,N_24687);
xor U25321 (N_25321,N_24521,N_20275);
and U25322 (N_25322,N_21384,N_24487);
xnor U25323 (N_25323,N_20444,N_22184);
nor U25324 (N_25324,N_21880,N_23153);
or U25325 (N_25325,N_21376,N_24000);
and U25326 (N_25326,N_22256,N_22282);
or U25327 (N_25327,N_24904,N_22347);
xor U25328 (N_25328,N_23505,N_23414);
nand U25329 (N_25329,N_24161,N_24417);
xor U25330 (N_25330,N_21834,N_22705);
and U25331 (N_25331,N_20696,N_20885);
nor U25332 (N_25332,N_21194,N_23353);
xor U25333 (N_25333,N_23633,N_22574);
xor U25334 (N_25334,N_23675,N_23280);
xnor U25335 (N_25335,N_20487,N_24820);
nor U25336 (N_25336,N_23740,N_20375);
nor U25337 (N_25337,N_21503,N_21156);
xor U25338 (N_25338,N_22377,N_22406);
and U25339 (N_25339,N_24163,N_24644);
or U25340 (N_25340,N_20385,N_23294);
xor U25341 (N_25341,N_24759,N_22173);
or U25342 (N_25342,N_22728,N_24600);
or U25343 (N_25343,N_24762,N_22128);
and U25344 (N_25344,N_23527,N_23916);
nor U25345 (N_25345,N_24667,N_24903);
and U25346 (N_25346,N_22024,N_23717);
and U25347 (N_25347,N_23212,N_22353);
nand U25348 (N_25348,N_20692,N_24967);
xor U25349 (N_25349,N_20846,N_22344);
nor U25350 (N_25350,N_23558,N_22735);
nand U25351 (N_25351,N_21729,N_24347);
nand U25352 (N_25352,N_20605,N_23287);
nand U25353 (N_25353,N_23107,N_23474);
or U25354 (N_25354,N_22670,N_20248);
nand U25355 (N_25355,N_21495,N_24708);
and U25356 (N_25356,N_23237,N_24059);
nor U25357 (N_25357,N_24291,N_22461);
or U25358 (N_25358,N_23863,N_21302);
nand U25359 (N_25359,N_20302,N_23172);
nand U25360 (N_25360,N_22198,N_23087);
nand U25361 (N_25361,N_24226,N_20724);
or U25362 (N_25362,N_20224,N_23370);
nand U25363 (N_25363,N_23451,N_20393);
xnor U25364 (N_25364,N_23446,N_23116);
or U25365 (N_25365,N_23487,N_20742);
nand U25366 (N_25366,N_23444,N_22947);
or U25367 (N_25367,N_24200,N_20043);
or U25368 (N_25368,N_21716,N_23137);
nor U25369 (N_25369,N_22929,N_24533);
and U25370 (N_25370,N_22804,N_23515);
nand U25371 (N_25371,N_24786,N_21110);
or U25372 (N_25372,N_21186,N_21162);
nor U25373 (N_25373,N_23986,N_21197);
xnor U25374 (N_25374,N_23905,N_22710);
or U25375 (N_25375,N_21884,N_20185);
nor U25376 (N_25376,N_20954,N_21883);
nand U25377 (N_25377,N_24824,N_20079);
or U25378 (N_25378,N_24119,N_24613);
nor U25379 (N_25379,N_23624,N_20648);
nor U25380 (N_25380,N_21737,N_23786);
and U25381 (N_25381,N_23157,N_20896);
nand U25382 (N_25382,N_23423,N_21025);
or U25383 (N_25383,N_21602,N_23862);
xor U25384 (N_25384,N_22276,N_21804);
and U25385 (N_25385,N_24509,N_23938);
nor U25386 (N_25386,N_24793,N_22513);
nand U25387 (N_25387,N_22111,N_22605);
and U25388 (N_25388,N_20661,N_21408);
or U25389 (N_25389,N_22460,N_21089);
or U25390 (N_25390,N_24009,N_20671);
xor U25391 (N_25391,N_22288,N_24901);
xor U25392 (N_25392,N_23188,N_20241);
xor U25393 (N_25393,N_24535,N_23046);
or U25394 (N_25394,N_20784,N_23024);
nor U25395 (N_25395,N_23244,N_21610);
or U25396 (N_25396,N_21018,N_23861);
and U25397 (N_25397,N_22686,N_22685);
and U25398 (N_25398,N_21941,N_21964);
nor U25399 (N_25399,N_22697,N_24263);
and U25400 (N_25400,N_22234,N_22576);
xor U25401 (N_25401,N_21661,N_23201);
and U25402 (N_25402,N_23075,N_24593);
nand U25403 (N_25403,N_24770,N_24128);
and U25404 (N_25404,N_22243,N_20744);
and U25405 (N_25405,N_23101,N_21802);
and U25406 (N_25406,N_23635,N_21521);
nand U25407 (N_25407,N_23405,N_21122);
nand U25408 (N_25408,N_21961,N_24033);
nor U25409 (N_25409,N_22269,N_21410);
or U25410 (N_25410,N_20796,N_21205);
xor U25411 (N_25411,N_24024,N_23104);
nor U25412 (N_25412,N_21873,N_20875);
nand U25413 (N_25413,N_23727,N_21701);
and U25414 (N_25414,N_20738,N_22606);
or U25415 (N_25415,N_24310,N_21164);
nor U25416 (N_25416,N_24905,N_23136);
and U25417 (N_25417,N_20086,N_23517);
nand U25418 (N_25418,N_23482,N_21748);
and U25419 (N_25419,N_23571,N_24380);
and U25420 (N_25420,N_23543,N_21020);
nor U25421 (N_25421,N_21457,N_24081);
xor U25422 (N_25422,N_20817,N_20511);
and U25423 (N_25423,N_24475,N_24711);
or U25424 (N_25424,N_22835,N_21188);
and U25425 (N_25425,N_22836,N_21916);
and U25426 (N_25426,N_20202,N_24657);
nand U25427 (N_25427,N_22885,N_22578);
and U25428 (N_25428,N_22747,N_22150);
xor U25429 (N_25429,N_20148,N_20031);
and U25430 (N_25430,N_22913,N_21782);
xnor U25431 (N_25431,N_23981,N_24865);
nand U25432 (N_25432,N_21832,N_23050);
nand U25433 (N_25433,N_23810,N_21009);
and U25434 (N_25434,N_23564,N_24562);
nor U25435 (N_25435,N_20474,N_23315);
nand U25436 (N_25436,N_21866,N_24448);
nor U25437 (N_25437,N_22715,N_21997);
xnor U25438 (N_25438,N_22213,N_24356);
and U25439 (N_25439,N_22627,N_24428);
nand U25440 (N_25440,N_21172,N_24321);
or U25441 (N_25441,N_22092,N_24162);
or U25442 (N_25442,N_20192,N_21721);
nand U25443 (N_25443,N_21662,N_24046);
and U25444 (N_25444,N_24416,N_20378);
and U25445 (N_25445,N_22855,N_22370);
or U25446 (N_25446,N_22897,N_21029);
nor U25447 (N_25447,N_23578,N_20537);
and U25448 (N_25448,N_22766,N_24577);
nand U25449 (N_25449,N_24083,N_22968);
nand U25450 (N_25450,N_21119,N_21520);
or U25451 (N_25451,N_21776,N_23164);
nand U25452 (N_25452,N_23488,N_20351);
xor U25453 (N_25453,N_20388,N_23134);
nand U25454 (N_25454,N_23325,N_24425);
or U25455 (N_25455,N_21138,N_24032);
and U25456 (N_25456,N_23067,N_23504);
or U25457 (N_25457,N_23559,N_24063);
and U25458 (N_25458,N_23952,N_24895);
and U25459 (N_25459,N_20497,N_21171);
and U25460 (N_25460,N_24283,N_24722);
or U25461 (N_25461,N_24027,N_22081);
and U25462 (N_25462,N_23500,N_23749);
nand U25463 (N_25463,N_23495,N_24842);
xor U25464 (N_25464,N_23982,N_23173);
nand U25465 (N_25465,N_24921,N_23250);
nor U25466 (N_25466,N_23783,N_24385);
nand U25467 (N_25467,N_23178,N_21596);
or U25468 (N_25468,N_20207,N_22399);
xor U25469 (N_25469,N_21059,N_22108);
nand U25470 (N_25470,N_23031,N_21851);
nand U25471 (N_25471,N_24209,N_23681);
or U25472 (N_25472,N_21709,N_22432);
nand U25473 (N_25473,N_22508,N_21441);
nand U25474 (N_25474,N_21920,N_20323);
nor U25475 (N_25475,N_23035,N_23947);
nor U25476 (N_25476,N_20535,N_23115);
nand U25477 (N_25477,N_24883,N_22494);
xor U25478 (N_25478,N_20164,N_21068);
nand U25479 (N_25479,N_21619,N_23169);
xor U25480 (N_25480,N_21168,N_21581);
and U25481 (N_25481,N_23813,N_21033);
or U25482 (N_25482,N_21762,N_23264);
or U25483 (N_25483,N_24954,N_24211);
or U25484 (N_25484,N_20960,N_22403);
or U25485 (N_25485,N_21028,N_21260);
nand U25486 (N_25486,N_21914,N_20600);
xnor U25487 (N_25487,N_24552,N_20797);
nand U25488 (N_25488,N_20128,N_24299);
and U25489 (N_25489,N_20409,N_23679);
and U25490 (N_25490,N_21650,N_22690);
nand U25491 (N_25491,N_23605,N_24148);
or U25492 (N_25492,N_23282,N_20991);
or U25493 (N_25493,N_21142,N_24010);
nand U25494 (N_25494,N_23199,N_24779);
and U25495 (N_25495,N_23346,N_23058);
or U25496 (N_25496,N_23300,N_21970);
and U25497 (N_25497,N_21840,N_23436);
and U25498 (N_25498,N_20435,N_23079);
and U25499 (N_25499,N_21565,N_20855);
nand U25500 (N_25500,N_21785,N_22005);
nand U25501 (N_25501,N_22914,N_21272);
xnor U25502 (N_25502,N_20247,N_20482);
and U25503 (N_25503,N_22629,N_23610);
and U25504 (N_25504,N_22321,N_24382);
and U25505 (N_25505,N_21097,N_22653);
or U25506 (N_25506,N_21871,N_24486);
nor U25507 (N_25507,N_21428,N_24139);
nand U25508 (N_25508,N_23897,N_22176);
nor U25509 (N_25509,N_24312,N_21333);
and U25510 (N_25510,N_20595,N_20333);
and U25511 (N_25511,N_24925,N_20413);
xnor U25512 (N_25512,N_22677,N_21885);
and U25513 (N_25513,N_20956,N_22046);
nand U25514 (N_25514,N_20242,N_23216);
xnor U25515 (N_25515,N_21386,N_21926);
and U25516 (N_25516,N_23730,N_22125);
nand U25517 (N_25517,N_20177,N_20234);
xnor U25518 (N_25518,N_20418,N_24982);
nand U25519 (N_25519,N_24154,N_22902);
nand U25520 (N_25520,N_23077,N_24626);
nand U25521 (N_25521,N_23481,N_23430);
or U25522 (N_25522,N_21017,N_20092);
xor U25523 (N_25523,N_24319,N_20786);
nand U25524 (N_25524,N_24257,N_23138);
or U25525 (N_25525,N_22573,N_20637);
and U25526 (N_25526,N_22030,N_20169);
nor U25527 (N_25527,N_22383,N_23708);
nor U25528 (N_25528,N_23320,N_22767);
and U25529 (N_25529,N_22559,N_23752);
xnor U25530 (N_25530,N_21274,N_20368);
nand U25531 (N_25531,N_20101,N_23307);
and U25532 (N_25532,N_23209,N_20126);
or U25533 (N_25533,N_23726,N_23124);
nor U25534 (N_25534,N_23296,N_22355);
nand U25535 (N_25535,N_23555,N_23015);
or U25536 (N_25536,N_21118,N_20459);
nor U25537 (N_25537,N_20950,N_20257);
nand U25538 (N_25538,N_24610,N_22596);
and U25539 (N_25539,N_21372,N_21911);
nand U25540 (N_25540,N_22599,N_20966);
and U25541 (N_25541,N_21652,N_20119);
nand U25542 (N_25542,N_20691,N_21952);
or U25543 (N_25543,N_24689,N_22765);
xnor U25544 (N_25544,N_22497,N_23367);
xnor U25545 (N_25545,N_23724,N_21369);
nand U25546 (N_25546,N_22145,N_21299);
nand U25547 (N_25547,N_24773,N_24873);
xnor U25548 (N_25548,N_23338,N_24975);
nor U25549 (N_25549,N_24726,N_22036);
or U25550 (N_25550,N_20492,N_20639);
or U25551 (N_25551,N_20852,N_21635);
nand U25552 (N_25552,N_20609,N_22942);
nor U25553 (N_25553,N_24939,N_24551);
xor U25554 (N_25554,N_24145,N_21535);
or U25555 (N_25555,N_20065,N_24179);
or U25556 (N_25556,N_22099,N_22853);
and U25557 (N_25557,N_20494,N_20630);
and U25558 (N_25558,N_20972,N_20199);
and U25559 (N_25559,N_20976,N_23083);
and U25560 (N_25560,N_21759,N_20037);
or U25561 (N_25561,N_24989,N_21736);
nor U25562 (N_25562,N_21502,N_24548);
or U25563 (N_25563,N_21256,N_20808);
or U25564 (N_25564,N_24937,N_24498);
and U25565 (N_25565,N_23834,N_24730);
nand U25566 (N_25566,N_22268,N_20319);
xor U25567 (N_25567,N_24745,N_21129);
nand U25568 (N_25568,N_20908,N_24744);
nor U25569 (N_25569,N_24640,N_22577);
nor U25570 (N_25570,N_21546,N_21202);
nor U25571 (N_25571,N_20299,N_21321);
or U25572 (N_25572,N_23868,N_20342);
and U25573 (N_25573,N_23586,N_23967);
or U25574 (N_25574,N_20431,N_24941);
or U25575 (N_25575,N_20091,N_23875);
or U25576 (N_25576,N_22066,N_20931);
or U25577 (N_25577,N_21151,N_20667);
nand U25578 (N_25578,N_22142,N_24885);
or U25579 (N_25579,N_24601,N_22249);
nor U25580 (N_25580,N_21426,N_23223);
and U25581 (N_25581,N_20032,N_20345);
xor U25582 (N_25582,N_23218,N_21243);
nor U25583 (N_25583,N_22254,N_20014);
and U25584 (N_25584,N_22073,N_21536);
nor U25585 (N_25585,N_21266,N_22290);
nor U25586 (N_25586,N_21967,N_24785);
nand U25587 (N_25587,N_20531,N_22391);
and U25588 (N_25588,N_23467,N_23113);
and U25589 (N_25589,N_24802,N_21747);
nor U25590 (N_25590,N_21909,N_22118);
nand U25591 (N_25591,N_22628,N_20426);
xor U25592 (N_25592,N_22971,N_22110);
or U25593 (N_25593,N_23593,N_23669);
nand U25594 (N_25594,N_23108,N_21934);
or U25595 (N_25595,N_20307,N_20745);
xnor U25596 (N_25596,N_23012,N_21554);
or U25597 (N_25597,N_21975,N_20666);
nor U25598 (N_25598,N_23530,N_23027);
xor U25599 (N_25599,N_24597,N_23547);
and U25600 (N_25600,N_22199,N_22676);
xnor U25601 (N_25601,N_23579,N_20665);
or U25602 (N_25602,N_22200,N_22169);
nand U25603 (N_25603,N_23475,N_20886);
nor U25604 (N_25604,N_22397,N_21888);
nand U25605 (N_25605,N_21350,N_21074);
and U25606 (N_25606,N_22222,N_21000);
or U25607 (N_25607,N_20364,N_22064);
or U25608 (N_25608,N_20858,N_20518);
and U25609 (N_25609,N_20500,N_22023);
xor U25610 (N_25610,N_24160,N_22424);
nor U25611 (N_25611,N_21796,N_24678);
and U25612 (N_25612,N_20862,N_22372);
or U25613 (N_25613,N_20096,N_23394);
nand U25614 (N_25614,N_21270,N_23450);
nor U25615 (N_25615,N_21827,N_23215);
nor U25616 (N_25616,N_23318,N_22204);
nor U25617 (N_25617,N_23063,N_21040);
or U25618 (N_25618,N_24026,N_20020);
nand U25619 (N_25619,N_22038,N_23032);
and U25620 (N_25620,N_22792,N_21160);
nor U25621 (N_25621,N_23052,N_22927);
and U25622 (N_25622,N_20047,N_23838);
xor U25623 (N_25623,N_22158,N_21891);
and U25624 (N_25624,N_23972,N_20704);
xnor U25625 (N_25625,N_22623,N_21571);
xor U25626 (N_25626,N_23372,N_21859);
or U25627 (N_25627,N_24080,N_24840);
xor U25628 (N_25628,N_24527,N_24133);
and U25629 (N_25629,N_22305,N_22619);
and U25630 (N_25630,N_20994,N_20196);
nand U25631 (N_25631,N_21923,N_24039);
nand U25632 (N_25632,N_21431,N_23171);
xnor U25633 (N_25633,N_22456,N_20841);
and U25634 (N_25634,N_24420,N_23606);
or U25635 (N_25635,N_24466,N_20503);
and U25636 (N_25636,N_21108,N_22115);
or U25637 (N_25637,N_24727,N_21338);
and U25638 (N_25638,N_21666,N_21393);
nor U25639 (N_25639,N_20265,N_23584);
or U25640 (N_25640,N_21965,N_20756);
nand U25641 (N_25641,N_21087,N_21358);
xor U25642 (N_25642,N_20640,N_22483);
xor U25643 (N_25643,N_24352,N_22934);
nor U25644 (N_25644,N_21073,N_23529);
xnor U25645 (N_25645,N_23788,N_20243);
and U25646 (N_25646,N_24305,N_22597);
or U25647 (N_25647,N_21198,N_23867);
or U25648 (N_25648,N_23049,N_23615);
or U25649 (N_25649,N_20327,N_21191);
nand U25650 (N_25650,N_24950,N_22773);
xnor U25651 (N_25651,N_21378,N_20335);
or U25652 (N_25652,N_22946,N_20499);
and U25653 (N_25653,N_21678,N_23279);
xnor U25654 (N_25654,N_24402,N_22078);
and U25655 (N_25655,N_24110,N_23371);
or U25656 (N_25656,N_20432,N_24813);
nand U25657 (N_25657,N_22226,N_24654);
nand U25658 (N_25658,N_23424,N_21366);
nor U25659 (N_25659,N_24962,N_22825);
xor U25660 (N_25660,N_21398,N_22362);
nor U25661 (N_25661,N_20578,N_23566);
nor U25662 (N_25662,N_22554,N_21027);
nor U25663 (N_25663,N_21220,N_24164);
xnor U25664 (N_25664,N_22941,N_22393);
nor U25665 (N_25665,N_23980,N_24275);
nor U25666 (N_25666,N_23043,N_20763);
xnor U25667 (N_25667,N_23540,N_20463);
or U25668 (N_25668,N_23358,N_21963);
or U25669 (N_25669,N_22587,N_24598);
and U25670 (N_25670,N_20188,N_22998);
xnor U25671 (N_25671,N_23640,N_20506);
and U25672 (N_25672,N_20557,N_23797);
nand U25673 (N_25673,N_24924,N_24774);
nand U25674 (N_25674,N_22032,N_20780);
or U25675 (N_25675,N_24725,N_23140);
nor U25676 (N_25676,N_23628,N_21212);
or U25677 (N_25677,N_20688,N_22845);
nand U25678 (N_25678,N_22161,N_20235);
and U25679 (N_25679,N_23833,N_21945);
nand U25680 (N_25680,N_20262,N_20638);
or U25681 (N_25681,N_23160,N_24278);
xnor U25682 (N_25682,N_24423,N_21726);
xnor U25683 (N_25683,N_22840,N_21070);
and U25684 (N_25684,N_20442,N_24093);
xor U25685 (N_25685,N_21133,N_24455);
or U25686 (N_25686,N_24694,N_20569);
nor U25687 (N_25687,N_22431,N_23846);
or U25688 (N_25688,N_23626,N_20703);
or U25689 (N_25689,N_24215,N_20029);
and U25690 (N_25690,N_21052,N_22886);
nor U25691 (N_25691,N_21649,N_22450);
xor U25692 (N_25692,N_24121,N_24868);
nor U25693 (N_25693,N_23328,N_22764);
nand U25694 (N_25694,N_21676,N_22572);
nor U25695 (N_25695,N_22195,N_22881);
and U25696 (N_25696,N_24030,N_20543);
and U25697 (N_25697,N_21233,N_23014);
and U25698 (N_25698,N_24244,N_22172);
nor U25699 (N_25699,N_22797,N_21377);
xor U25700 (N_25700,N_22149,N_23782);
nor U25701 (N_25701,N_21697,N_23435);
xor U25702 (N_25702,N_23380,N_22553);
nor U25703 (N_25703,N_20755,N_22339);
or U25704 (N_25704,N_21533,N_21695);
nor U25705 (N_25705,N_21245,N_20253);
and U25706 (N_25706,N_22275,N_24706);
nor U25707 (N_25707,N_22244,N_24442);
or U25708 (N_25708,N_23093,N_24343);
nor U25709 (N_25709,N_23448,N_23419);
xnor U25710 (N_25710,N_23565,N_24190);
or U25711 (N_25711,N_23772,N_23620);
nand U25712 (N_25712,N_24876,N_23691);
nand U25713 (N_25713,N_23599,N_20546);
xor U25714 (N_25714,N_20983,N_24743);
and U25715 (N_25715,N_21587,N_20451);
xor U25716 (N_25716,N_22453,N_24308);
and U25717 (N_25717,N_23594,N_23873);
or U25718 (N_25718,N_21181,N_21230);
and U25719 (N_25719,N_22608,N_23351);
and U25720 (N_25720,N_22691,N_23190);
xnor U25721 (N_25721,N_23901,N_23964);
or U25722 (N_25722,N_21214,N_20062);
xnor U25723 (N_25723,N_22642,N_23030);
or U25724 (N_25724,N_21563,N_23796);
nor U25725 (N_25725,N_24993,N_23720);
xnor U25726 (N_25726,N_23842,N_24467);
or U25727 (N_25727,N_20558,N_22643);
xor U25728 (N_25728,N_24734,N_21279);
and U25729 (N_25729,N_23654,N_20166);
and U25730 (N_25730,N_22015,N_21958);
nor U25731 (N_25731,N_23428,N_21844);
or U25732 (N_25732,N_21773,N_22386);
nand U25733 (N_25733,N_20211,N_20574);
xnor U25734 (N_25734,N_21854,N_21910);
nand U25735 (N_25735,N_24973,N_20090);
nor U25736 (N_25736,N_22439,N_22472);
nor U25737 (N_25737,N_24100,N_21276);
xnor U25738 (N_25738,N_23438,N_20857);
and U25739 (N_25739,N_21707,N_22361);
or U25740 (N_25740,N_24044,N_20850);
nand U25741 (N_25741,N_20088,N_22901);
xor U25742 (N_25742,N_24176,N_22235);
and U25743 (N_25743,N_23211,N_24193);
and U25744 (N_25744,N_20411,N_23622);
or U25745 (N_25745,N_21297,N_20821);
and U25746 (N_25746,N_21071,N_22872);
and U25747 (N_25747,N_22444,N_24254);
and U25748 (N_25748,N_23902,N_23957);
or U25749 (N_25749,N_24304,N_23983);
or U25750 (N_25750,N_24208,N_23954);
xor U25751 (N_25751,N_20412,N_22748);
nor U25752 (N_25752,N_22033,N_21486);
nor U25753 (N_25753,N_21591,N_20424);
and U25754 (N_25754,N_21744,N_21806);
nor U25755 (N_25755,N_24716,N_23080);
nand U25756 (N_25756,N_23234,N_22068);
or U25757 (N_25757,N_21614,N_22954);
xnor U25758 (N_25758,N_23422,N_23756);
or U25759 (N_25759,N_24616,N_20532);
nor U25760 (N_25760,N_23130,N_24790);
nor U25761 (N_25761,N_22352,N_22055);
or U25762 (N_25762,N_22000,N_21882);
or U25763 (N_25763,N_20768,N_21549);
or U25764 (N_25764,N_24898,N_23376);
nand U25765 (N_25765,N_23688,N_21578);
or U25766 (N_25766,N_20656,N_21927);
xnor U25767 (N_25767,N_21250,N_23183);
or U25768 (N_25768,N_23999,N_24826);
xnor U25769 (N_25769,N_20138,N_22631);
xnor U25770 (N_25770,N_21886,N_24368);
nor U25771 (N_25771,N_20876,N_20038);
nor U25772 (N_25772,N_21438,N_22819);
nor U25773 (N_25773,N_21054,N_20927);
nor U25774 (N_25774,N_24367,N_20021);
xnor U25775 (N_25775,N_22003,N_20870);
or U25776 (N_25776,N_24112,N_22134);
nand U25777 (N_25777,N_20619,N_21559);
nor U25778 (N_25778,N_22548,N_21765);
nand U25779 (N_25779,N_21705,N_23231);
and U25780 (N_25780,N_20407,N_22862);
and U25781 (N_25781,N_21248,N_22263);
or U25782 (N_25782,N_21490,N_23821);
nand U25783 (N_25783,N_24872,N_20851);
and U25784 (N_25784,N_21050,N_24513);
and U25785 (N_25785,N_21498,N_21869);
or U25786 (N_25786,N_22614,N_22603);
nand U25787 (N_25787,N_22663,N_24077);
or U25788 (N_25788,N_23013,N_23006);
nor U25789 (N_25789,N_21450,N_24894);
or U25790 (N_25790,N_23496,N_21643);
nor U25791 (N_25791,N_20056,N_20674);
or U25792 (N_25792,N_20859,N_23143);
and U25793 (N_25793,N_22301,N_24065);
xor U25794 (N_25794,N_23065,N_24414);
xnor U25795 (N_25795,N_22622,N_23129);
xnor U25796 (N_25796,N_23512,N_20168);
nor U25797 (N_25797,N_23870,N_22098);
or U25798 (N_25798,N_23814,N_21826);
nor U25799 (N_25799,N_23638,N_21222);
or U25800 (N_25800,N_23754,N_24671);
nand U25801 (N_25801,N_24896,N_21080);
nand U25802 (N_25802,N_22217,N_23528);
and U25803 (N_25803,N_24550,N_22381);
and U25804 (N_25804,N_22979,N_20611);
or U25805 (N_25805,N_22939,N_22626);
nand U25806 (N_25806,N_21128,N_21810);
nand U25807 (N_25807,N_20370,N_24970);
and U25808 (N_25808,N_20585,N_24624);
nand U25809 (N_25809,N_23818,N_24986);
nor U25810 (N_25810,N_24130,N_23687);
or U25811 (N_25811,N_22325,N_22345);
nor U25812 (N_25812,N_20798,N_24567);
or U25813 (N_25813,N_24966,N_20549);
xnor U25814 (N_25814,N_22724,N_20920);
xnor U25815 (N_25815,N_20183,N_20080);
nand U25816 (N_25816,N_20100,N_22749);
nor U25817 (N_25817,N_22544,N_20897);
xor U25818 (N_25818,N_21858,N_21951);
nor U25819 (N_25819,N_24912,N_22740);
nand U25820 (N_25820,N_21343,N_23295);
nand U25821 (N_25821,N_20095,N_20854);
nor U25822 (N_25822,N_22320,N_22480);
or U25823 (N_25823,N_24288,N_23368);
and U25824 (N_25824,N_23777,N_20213);
nor U25825 (N_25825,N_23966,N_21634);
nand U25826 (N_25826,N_23989,N_22248);
xor U25827 (N_25827,N_22006,N_20152);
xor U25828 (N_25828,N_21148,N_24069);
nor U25829 (N_25829,N_23892,N_21739);
xnor U25830 (N_25830,N_22408,N_20868);
nor U25831 (N_25831,N_21595,N_22820);
nand U25832 (N_25832,N_20764,N_24555);
and U25833 (N_25833,N_20524,N_22096);
nor U25834 (N_25834,N_24249,N_22937);
xor U25835 (N_25835,N_20131,N_21166);
nor U25836 (N_25836,N_23410,N_22136);
or U25837 (N_25837,N_22049,N_21938);
xnor U25838 (N_25838,N_24342,N_21821);
nand U25839 (N_25839,N_23580,N_20534);
or U25840 (N_25840,N_23243,N_24919);
xnor U25841 (N_25841,N_20973,N_24767);
and U25842 (N_25842,N_23747,N_20137);
nand U25843 (N_25843,N_22333,N_20561);
or U25844 (N_25844,N_24836,N_24106);
xor U25845 (N_25845,N_24563,N_23618);
nand U25846 (N_25846,N_22970,N_21456);
nor U25847 (N_25847,N_24350,N_24231);
and U25848 (N_25848,N_21574,N_21680);
or U25849 (N_25849,N_23266,N_24159);
or U25850 (N_25850,N_22646,N_24041);
and U25851 (N_25851,N_24472,N_21267);
xor U25852 (N_25852,N_23466,N_23914);
xor U25853 (N_25853,N_22775,N_23588);
and U25854 (N_25854,N_21894,N_22534);
or U25855 (N_25855,N_23656,N_21219);
nor U25856 (N_25856,N_21702,N_21293);
xnor U25857 (N_25857,N_20214,N_21682);
xnor U25858 (N_25858,N_22394,N_22799);
nor U25859 (N_25859,N_24651,N_23274);
nor U25860 (N_25860,N_24203,N_22181);
nand U25861 (N_25861,N_20448,N_21123);
xor U25862 (N_25862,N_22936,N_20312);
nand U25863 (N_25863,N_20864,N_24963);
nand U25864 (N_25864,N_24782,N_24138);
nor U25865 (N_25865,N_23141,N_22487);
nand U25866 (N_25866,N_20765,N_23761);
xnor U25867 (N_25867,N_22152,N_21314);
and U25868 (N_25868,N_22458,N_23541);
xnor U25869 (N_25869,N_23508,N_21672);
xor U25870 (N_25870,N_24075,N_23713);
nor U25871 (N_25871,N_24101,N_22153);
or U25872 (N_25872,N_22223,N_24686);
or U25873 (N_25873,N_23061,N_24008);
xor U25874 (N_25874,N_22208,N_22684);
or U25875 (N_25875,N_24653,N_24322);
nor U25876 (N_25876,N_20916,N_20525);
nand U25877 (N_25877,N_24248,N_21190);
xnor U25878 (N_25878,N_22501,N_23745);
or U25879 (N_25879,N_22769,N_22018);
or U25880 (N_25880,N_20336,N_24676);
and U25881 (N_25881,N_24401,N_21657);
or U25882 (N_25882,N_23664,N_24575);
nor U25883 (N_25883,N_22751,N_21541);
xnor U25884 (N_25884,N_20256,N_20274);
or U25885 (N_25885,N_23096,N_20953);
xor U25886 (N_25886,N_23238,N_20658);
xnor U25887 (N_25887,N_21416,N_23489);
nand U25888 (N_25888,N_20636,N_24923);
and U25889 (N_25889,N_20039,N_20686);
nand U25890 (N_25890,N_22459,N_20978);
nor U25891 (N_25891,N_22616,N_23312);
and U25892 (N_25892,N_22101,N_23227);
nand U25893 (N_25893,N_21720,N_23076);
xnor U25894 (N_25894,N_23969,N_22652);
xnor U25895 (N_25895,N_22065,N_23699);
and U25896 (N_25896,N_21508,N_23283);
nor U25897 (N_25897,N_23894,N_22516);
nor U25898 (N_25898,N_20464,N_24109);
and U25899 (N_25899,N_24977,N_23292);
and U25900 (N_25900,N_21402,N_21217);
nand U25901 (N_25901,N_21311,N_22343);
nand U25902 (N_25902,N_20384,N_21930);
xnor U25903 (N_25903,N_22549,N_21030);
xnor U25904 (N_25904,N_20399,N_21828);
nor U25905 (N_25905,N_24098,N_24777);
and U25906 (N_25906,N_24763,N_23655);
xnor U25907 (N_25907,N_24184,N_22084);
or U25908 (N_25908,N_20392,N_23841);
and U25909 (N_25909,N_23337,N_24611);
or U25910 (N_25910,N_23305,N_23582);
or U25911 (N_25911,N_21921,N_20509);
nor U25912 (N_25912,N_24316,N_22695);
xor U25913 (N_25913,N_24720,N_22289);
or U25914 (N_25914,N_22253,N_24675);
nor U25915 (N_25915,N_24655,N_24879);
or U25916 (N_25916,N_22433,N_21553);
xor U25917 (N_25917,N_23099,N_20254);
and U25918 (N_25918,N_20527,N_21224);
nor U25919 (N_25919,N_22177,N_22438);
xnor U25920 (N_25920,N_24462,N_20259);
and U25921 (N_25921,N_24605,N_22194);
or U25922 (N_25922,N_22959,N_24942);
nand U25923 (N_25923,N_21513,N_21861);
or U25924 (N_25924,N_24698,N_23456);
nand U25925 (N_25925,N_20376,N_24223);
nand U25926 (N_25926,N_24594,N_22944);
nand U25927 (N_25927,N_20292,N_24246);
nand U25928 (N_25928,N_21706,N_20616);
nand U25929 (N_25929,N_23222,N_20866);
xor U25930 (N_25930,N_23513,N_22933);
nor U25931 (N_25931,N_24378,N_20730);
xnor U25932 (N_25932,N_24528,N_23364);
or U25933 (N_25933,N_22903,N_23526);
xnor U25934 (N_25934,N_23003,N_22783);
xnor U25935 (N_25935,N_21588,N_20200);
or U25936 (N_25936,N_22373,N_24943);
or U25937 (N_25937,N_23631,N_24015);
and U25938 (N_25938,N_22267,N_24180);
nand U25939 (N_25939,N_20971,N_20699);
xnor U25940 (N_25940,N_21653,N_20405);
and U25941 (N_25941,N_21038,N_21741);
nand U25942 (N_25942,N_22641,N_23029);
or U25943 (N_25943,N_24662,N_21523);
nor U25944 (N_25944,N_21387,N_21154);
xor U25945 (N_25945,N_21093,N_22988);
xnor U25946 (N_25946,N_22535,N_22056);
and U25947 (N_25947,N_22703,N_23297);
or U25948 (N_25948,N_22858,N_22857);
nor U25949 (N_25949,N_21026,N_21406);
nand U25950 (N_25950,N_21252,N_20996);
nor U25951 (N_25951,N_20219,N_20593);
xnor U25952 (N_25952,N_22241,N_20267);
nand U25953 (N_25953,N_23133,N_23692);
or U25954 (N_25954,N_20221,N_23360);
or U25955 (N_25955,N_23017,N_20396);
nor U25956 (N_25956,N_22645,N_22088);
and U25957 (N_25957,N_22720,N_22167);
xnor U25958 (N_25958,N_23673,N_24554);
xnor U25959 (N_25959,N_24247,N_22299);
nor U25960 (N_25960,N_21929,N_21568);
nand U25961 (N_25961,N_24300,N_23816);
nor U25962 (N_25962,N_22219,N_20058);
xor U25963 (N_25963,N_24799,N_22699);
or U25964 (N_25964,N_20329,N_22621);
xor U25965 (N_25965,N_20874,N_23225);
nor U25966 (N_25966,N_23202,N_20641);
or U25967 (N_25967,N_20073,N_24882);
nor U25968 (N_25968,N_22563,N_24099);
and U25969 (N_25969,N_21342,N_23767);
nor U25970 (N_25970,N_24012,N_20145);
and U25971 (N_25971,N_22452,N_23154);
nand U25972 (N_25972,N_24105,N_21628);
nand U25973 (N_25973,N_23118,N_23009);
xor U25974 (N_25974,N_20900,N_22260);
and U25975 (N_25975,N_20708,N_24692);
and U25976 (N_25976,N_21145,N_21446);
or U25977 (N_25977,N_20050,N_21206);
nor U25978 (N_25978,N_20690,N_22923);
and U25979 (N_25979,N_24680,N_20070);
or U25980 (N_25980,N_21499,N_22112);
nand U25981 (N_25981,N_21752,N_21956);
or U25982 (N_25982,N_20162,N_22304);
nand U25983 (N_25983,N_20832,N_21900);
or U25984 (N_25984,N_21835,N_21176);
nand U25985 (N_25985,N_22696,N_24938);
nand U25986 (N_25986,N_24948,N_22197);
or U25987 (N_25987,N_20063,N_24150);
nand U25988 (N_25988,N_20212,N_23248);
nand U25989 (N_25989,N_24038,N_24672);
nand U25990 (N_25990,N_23275,N_23755);
or U25991 (N_25991,N_22546,N_24339);
nand U25992 (N_25992,N_21439,N_24732);
or U25993 (N_25993,N_24645,N_23652);
and U25994 (N_25994,N_22635,N_24817);
or U25995 (N_25995,N_21112,N_22727);
and U25996 (N_25996,N_21745,N_21394);
xnor U25997 (N_25997,N_20899,N_24369);
and U25998 (N_25998,N_24233,N_23604);
nor U25999 (N_25999,N_20709,N_24983);
nand U26000 (N_26000,N_24370,N_24742);
and U26001 (N_26001,N_22911,N_20813);
or U26002 (N_26002,N_20921,N_20258);
and U26003 (N_26003,N_21494,N_24845);
nand U26004 (N_26004,N_23357,N_22838);
and U26005 (N_26005,N_21895,N_21972);
nand U26006 (N_26006,N_21555,N_24837);
nand U26007 (N_26007,N_23903,N_22759);
xor U26008 (N_26008,N_21764,N_20305);
or U26009 (N_26009,N_22271,N_24849);
xor U26010 (N_26010,N_23906,N_20542);
xor U26011 (N_26011,N_22729,N_21771);
nor U26012 (N_26012,N_20677,N_23317);
nor U26013 (N_26013,N_20746,N_24830);
xnor U26014 (N_26014,N_24699,N_21723);
and U26015 (N_26015,N_24978,N_24074);
nor U26016 (N_26016,N_24090,N_20654);
nand U26017 (N_26017,N_22805,N_24731);
xnor U26018 (N_26018,N_20282,N_21413);
and U26019 (N_26019,N_21500,N_20579);
nor U26020 (N_26020,N_24739,N_24296);
or U26021 (N_26021,N_20515,N_24482);
nand U26022 (N_26022,N_24351,N_22545);
xnor U26023 (N_26023,N_20001,N_24652);
or U26024 (N_26024,N_21374,N_20044);
xor U26025 (N_26025,N_22847,N_20657);
xor U26026 (N_26026,N_23857,N_20801);
and U26027 (N_26027,N_22632,N_22486);
nand U26028 (N_26028,N_23941,N_21149);
nand U26029 (N_26029,N_20226,N_24326);
xnor U26030 (N_26030,N_24276,N_23149);
xnor U26031 (N_26031,N_23064,N_22337);
nand U26032 (N_26032,N_24891,N_24549);
nand U26033 (N_26033,N_20610,N_21484);
xnor U26034 (N_26034,N_21395,N_24858);
or U26035 (N_26035,N_24373,N_24082);
nor U26036 (N_26036,N_23680,N_22890);
nand U26037 (N_26037,N_21912,N_23705);
nor U26038 (N_26038,N_24328,N_20700);
or U26039 (N_26039,N_21175,N_24232);
nor U26040 (N_26040,N_24795,N_23682);
xnor U26041 (N_26041,N_21794,N_20584);
and U26042 (N_26042,N_24796,N_23743);
nor U26043 (N_26043,N_22485,N_23463);
nor U26044 (N_26044,N_23710,N_22874);
and U26045 (N_26045,N_23418,N_20072);
xor U26046 (N_26046,N_22196,N_24700);
nand U26047 (N_26047,N_23829,N_20872);
xor U26048 (N_26048,N_21999,N_22308);
and U26049 (N_26049,N_21522,N_23971);
or U26050 (N_26050,N_21823,N_20760);
or U26051 (N_26051,N_20721,N_24846);
and U26052 (N_26052,N_22045,N_20905);
or U26053 (N_26053,N_23385,N_23591);
xnor U26054 (N_26054,N_21575,N_23779);
and U26055 (N_26055,N_24994,N_24712);
or U26056 (N_26056,N_24262,N_24155);
and U26057 (N_26057,N_24197,N_20819);
nor U26058 (N_26058,N_21814,N_24526);
nor U26059 (N_26059,N_24413,N_21290);
nor U26060 (N_26060,N_24113,N_22314);
nand U26061 (N_26061,N_24783,N_21116);
and U26062 (N_26062,N_20747,N_20365);
xor U26063 (N_26063,N_24089,N_23912);
nor U26064 (N_26064,N_23869,N_20740);
xor U26065 (N_26065,N_24838,N_21993);
and U26066 (N_26066,N_20349,N_23089);
nor U26067 (N_26067,N_23085,N_24185);
xor U26068 (N_26068,N_22649,N_21221);
or U26069 (N_26069,N_23127,N_21786);
nor U26070 (N_26070,N_24596,N_22660);
and U26071 (N_26071,N_22107,N_21901);
xor U26072 (N_26072,N_20456,N_22958);
nor U26073 (N_26073,N_23927,N_23521);
nand U26074 (N_26074,N_24068,N_21251);
xor U26075 (N_26075,N_22600,N_20794);
xnor U26076 (N_26076,N_24642,N_23091);
nand U26077 (N_26077,N_24052,N_23286);
and U26078 (N_26078,N_22841,N_20889);
xor U26079 (N_26079,N_22785,N_23820);
xnor U26080 (N_26080,N_22205,N_24463);
nor U26081 (N_26081,N_21187,N_20936);
and U26082 (N_26082,N_21324,N_24207);
xnor U26083 (N_26083,N_21483,N_20570);
xnor U26084 (N_26084,N_24586,N_21935);
nand U26085 (N_26085,N_24446,N_23723);
nor U26086 (N_26086,N_23625,N_23773);
and U26087 (N_26087,N_21373,N_20485);
and U26088 (N_26088,N_23806,N_23343);
and U26089 (N_26089,N_21658,N_23329);
or U26090 (N_26090,N_21510,N_20078);
nor U26091 (N_26091,N_24952,N_24393);
and U26092 (N_26092,N_21157,N_24035);
xor U26093 (N_26093,N_23811,N_23426);
xnor U26094 (N_26094,N_20173,N_24571);
and U26095 (N_26095,N_22020,N_23507);
xnor U26096 (N_26096,N_22283,N_23390);
nand U26097 (N_26097,N_23544,N_20583);
and U26098 (N_26098,N_23764,N_21797);
nand U26099 (N_26099,N_23614,N_21807);
or U26100 (N_26100,N_20132,N_23028);
xnor U26101 (N_26101,N_22489,N_21609);
or U26102 (N_26102,N_22943,N_20103);
nor U26103 (N_26103,N_23589,N_23039);
and U26104 (N_26104,N_20337,N_23995);
or U26105 (N_26105,N_22731,N_21693);
or U26106 (N_26106,N_21955,N_22492);
xor U26107 (N_26107,N_22170,N_21006);
xor U26108 (N_26108,N_24588,N_21032);
xor U26109 (N_26109,N_20628,N_22409);
xnor U26110 (N_26110,N_20961,N_23915);
nand U26111 (N_26111,N_23403,N_21254);
or U26112 (N_26112,N_23005,N_20008);
xor U26113 (N_26113,N_23962,N_23442);
and U26114 (N_26114,N_20161,N_21102);
xnor U26115 (N_26115,N_24236,N_20726);
nand U26116 (N_26116,N_20158,N_24104);
and U26117 (N_26117,N_22552,N_20325);
and U26118 (N_26118,N_23407,N_20277);
nor U26119 (N_26119,N_20907,N_22752);
nor U26120 (N_26120,N_24881,N_22806);
nand U26121 (N_26121,N_24514,N_21509);
nand U26122 (N_26122,N_22522,N_24789);
or U26123 (N_26123,N_23472,N_21061);
nand U26124 (N_26124,N_21213,N_20892);
xnor U26125 (N_26125,N_22852,N_23876);
xnor U26126 (N_26126,N_22782,N_20938);
and U26127 (N_26127,N_21363,N_24997);
nand U26128 (N_26128,N_20877,N_22454);
nor U26129 (N_26129,N_21530,N_23850);
and U26130 (N_26130,N_22104,N_23257);
nand U26131 (N_26131,N_24332,N_22823);
or U26132 (N_26132,N_20932,N_20278);
and U26133 (N_26133,N_20943,N_20000);
and U26134 (N_26134,N_22809,N_21210);
xnor U26135 (N_26135,N_23400,N_20689);
or U26136 (N_26136,N_21688,N_24582);
xnor U26137 (N_26137,N_24465,N_23389);
nand U26138 (N_26138,N_21799,N_23411);
and U26139 (N_26139,N_21636,N_21246);
or U26140 (N_26140,N_22527,N_22448);
and U26141 (N_26141,N_24360,N_22427);
or U26142 (N_26142,N_22867,N_20998);
or U26143 (N_26143,N_21174,N_20510);
nand U26144 (N_26144,N_20647,N_21120);
and U26145 (N_26145,N_23460,N_23877);
xnor U26146 (N_26146,N_24468,N_21576);
xor U26147 (N_26147,N_23803,N_21385);
nor U26148 (N_26148,N_20075,N_22617);
or U26149 (N_26149,N_24957,N_21339);
and U26150 (N_26150,N_22303,N_20414);
xnor U26151 (N_26151,N_22816,N_20838);
nand U26152 (N_26152,N_24524,N_21326);
nor U26153 (N_26153,N_20844,N_21667);
nand U26154 (N_26154,N_20204,N_23182);
and U26155 (N_26155,N_20194,N_22499);
and U26156 (N_26156,N_22215,N_23235);
and U26157 (N_26157,N_20947,N_22114);
and U26158 (N_26158,N_23040,N_22185);
xor U26159 (N_26159,N_21534,N_23449);
or U26160 (N_26160,N_20629,N_22793);
nand U26161 (N_26161,N_21504,N_21558);
and U26162 (N_26162,N_24816,N_22651);
xnor U26163 (N_26163,N_21464,N_21950);
nand U26164 (N_26164,N_22363,N_24747);
or U26165 (N_26165,N_24451,N_23709);
xnor U26166 (N_26166,N_23519,N_22609);
nand U26167 (N_26167,N_23937,N_24935);
nor U26168 (N_26168,N_20030,N_22318);
and U26169 (N_26169,N_21114,N_24166);
or U26170 (N_26170,N_22429,N_23126);
xor U26171 (N_26171,N_21892,N_24481);
xor U26172 (N_26172,N_21981,N_23661);
or U26173 (N_26173,N_23732,N_24375);
xor U26174 (N_26174,N_23168,N_23738);
xnor U26175 (N_26175,N_21803,N_23748);
and U26176 (N_26176,N_23044,N_20587);
or U26177 (N_26177,N_20003,N_22790);
xnor U26178 (N_26178,N_20301,N_24136);
nand U26179 (N_26179,N_21679,N_20702);
or U26180 (N_26180,N_24115,N_20729);
xor U26181 (N_26181,N_22388,N_24062);
and U26182 (N_26182,N_21401,N_21654);
and U26183 (N_26183,N_20645,N_23856);
nand U26184 (N_26184,N_22159,N_21904);
nor U26185 (N_26185,N_22776,N_24290);
nand U26186 (N_26186,N_24028,N_21328);
nand U26187 (N_26187,N_22581,N_24403);
and U26188 (N_26188,N_24985,N_23890);
and U26189 (N_26189,N_20910,N_20568);
or U26190 (N_26190,N_20419,N_24269);
or U26191 (N_26191,N_22949,N_21184);
nand U26192 (N_26192,N_24387,N_22905);
nand U26193 (N_26193,N_22105,N_23155);
nor U26194 (N_26194,N_24807,N_22892);
or U26195 (N_26195,N_22848,N_24134);
and U26196 (N_26196,N_24797,N_20783);
xnor U26197 (N_26197,N_22041,N_24703);
nand U26198 (N_26198,N_21813,N_20809);
or U26199 (N_26199,N_22192,N_20328);
nor U26200 (N_26200,N_21552,N_24878);
and U26201 (N_26201,N_22644,N_20612);
nor U26202 (N_26202,N_24491,N_24556);
nand U26203 (N_26203,N_23047,N_21862);
nor U26204 (N_26204,N_20904,N_23885);
xnor U26205 (N_26205,N_24287,N_21442);
and U26206 (N_26206,N_20627,N_22967);
or U26207 (N_26207,N_20439,N_23462);
nor U26208 (N_26208,N_21757,N_21437);
xnor U26209 (N_26209,N_23194,N_23923);
xnor U26210 (N_26210,N_22238,N_21265);
or U26211 (N_26211,N_21257,N_24971);
nand U26212 (N_26212,N_23953,N_23511);
or U26213 (N_26213,N_23961,N_21984);
xnor U26214 (N_26214,N_22401,N_21512);
or U26215 (N_26215,N_22976,N_20230);
nand U26216 (N_26216,N_21261,N_21860);
nor U26217 (N_26217,N_23929,N_24437);
or U26218 (N_26218,N_20433,N_21282);
and U26219 (N_26219,N_20906,N_24058);
nor U26220 (N_26220,N_24006,N_23233);
nor U26221 (N_26221,N_23665,N_21887);
xor U26222 (N_26222,N_20924,N_20300);
xnor U26223 (N_26223,N_24292,N_23455);
nor U26224 (N_26224,N_23147,N_24913);
nor U26225 (N_26225,N_24981,N_22869);
nor U26226 (N_26226,N_21617,N_22570);
nor U26227 (N_26227,N_24780,N_23480);
and U26228 (N_26228,N_22980,N_21380);
nand U26229 (N_26229,N_22264,N_22907);
nor U26230 (N_26230,N_22610,N_22784);
and U26231 (N_26231,N_20969,N_21371);
nor U26232 (N_26232,N_24835,N_20251);
nand U26233 (N_26233,N_20112,N_21597);
and U26234 (N_26234,N_20670,N_24271);
nand U26235 (N_26235,N_21966,N_23135);
and U26236 (N_26236,N_23671,N_20767);
nand U26237 (N_26237,N_21412,N_23556);
and U26238 (N_26238,N_21472,N_20295);
xnor U26239 (N_26239,N_23184,N_24781);
or U26240 (N_26240,N_22509,N_20860);
or U26241 (N_26241,N_20184,N_23545);
nor U26242 (N_26242,N_24408,N_20923);
xnor U26243 (N_26243,N_21857,N_21127);
nand U26244 (N_26244,N_23355,N_24157);
or U26245 (N_26245,N_20015,N_21476);
nand U26246 (N_26246,N_24295,N_21390);
or U26247 (N_26247,N_22374,N_22022);
or U26248 (N_26248,N_23345,N_22495);
nor U26249 (N_26249,N_22008,N_24674);
nand U26250 (N_26250,N_20594,N_20962);
or U26251 (N_26251,N_22926,N_24501);
or U26252 (N_26252,N_20538,N_22179);
and U26253 (N_26253,N_22137,N_24456);
nor U26254 (N_26254,N_24409,N_21269);
nand U26255 (N_26255,N_21663,N_24353);
and U26256 (N_26256,N_22918,N_24146);
nor U26257 (N_26257,N_20268,N_24216);
nand U26258 (N_26258,N_21043,N_22859);
and U26259 (N_26259,N_23674,N_20098);
and U26260 (N_26260,N_20357,N_24839);
nor U26261 (N_26261,N_23285,N_22261);
xnor U26262 (N_26262,N_22537,N_23268);
nor U26263 (N_26263,N_20353,N_22983);
and U26264 (N_26264,N_24529,N_24202);
nor U26265 (N_26265,N_23246,N_21004);
and U26266 (N_26266,N_21023,N_22340);
nor U26267 (N_26267,N_23667,N_20460);
or U26268 (N_26268,N_22190,N_20149);
or U26269 (N_26269,N_22166,N_20915);
or U26270 (N_26270,N_20232,N_20935);
nand U26271 (N_26271,N_23263,N_20793);
nor U26272 (N_26272,N_22912,N_24002);
xor U26273 (N_26273,N_22536,N_22965);
nand U26274 (N_26274,N_21598,N_23896);
nand U26275 (N_26275,N_21917,N_20306);
or U26276 (N_26276,N_23608,N_23262);
or U26277 (N_26277,N_22744,N_23765);
nor U26278 (N_26278,N_21754,N_21354);
nand U26279 (N_26279,N_21656,N_24537);
and U26280 (N_26280,N_23051,N_22714);
and U26281 (N_26281,N_20735,N_22871);
nor U26282 (N_26282,N_23486,N_24395);
nand U26283 (N_26283,N_21590,N_20416);
or U26284 (N_26284,N_21660,N_20085);
nor U26285 (N_26285,N_22551,N_21969);
or U26286 (N_26286,N_24825,N_20475);
nand U26287 (N_26287,N_24500,N_21849);
or U26288 (N_26288,N_23161,N_24076);
nor U26289 (N_26289,N_21399,N_24506);
nor U26290 (N_26290,N_21336,N_24114);
nand U26291 (N_26291,N_21031,N_22981);
nor U26292 (N_26292,N_21049,N_22991);
nor U26293 (N_26293,N_22817,N_23766);
nand U26294 (N_26294,N_22542,N_20853);
and U26295 (N_26295,N_24129,N_23219);
xor U26296 (N_26296,N_24804,N_24705);
and U26297 (N_26297,N_23471,N_21165);
xor U26298 (N_26298,N_24457,N_21382);
or U26299 (N_26299,N_21420,N_22832);
and U26300 (N_26300,N_23798,N_21155);
or U26301 (N_26301,N_22013,N_23827);
nand U26302 (N_26302,N_21613,N_20122);
or U26303 (N_26303,N_21570,N_23026);
and U26304 (N_26304,N_22704,N_23036);
or U26305 (N_26305,N_23081,N_21491);
nand U26306 (N_26306,N_21231,N_21327);
nand U26307 (N_26307,N_22884,N_21897);
or U26308 (N_26308,N_24167,N_20404);
nor U26309 (N_26309,N_22722,N_23629);
and U26310 (N_26310,N_21481,N_22986);
or U26311 (N_26311,N_21604,N_22171);
nor U26312 (N_26312,N_20753,N_20310);
or U26313 (N_26313,N_22309,N_21150);
xor U26314 (N_26314,N_22580,N_21240);
nand U26315 (N_26315,N_24980,N_20563);
and U26316 (N_26316,N_23010,N_20602);
or U26317 (N_26317,N_20806,N_24313);
xor U26318 (N_26318,N_21117,N_23801);
nor U26319 (N_26319,N_22407,N_21863);
and U26320 (N_26320,N_24436,N_24438);
xnor U26321 (N_26321,N_21242,N_21467);
or U26322 (N_26322,N_22506,N_20303);
xnor U26323 (N_26323,N_24374,N_21121);
and U26324 (N_26324,N_22673,N_21124);
or U26325 (N_26325,N_20814,N_20967);
or U26326 (N_26326,N_21103,N_21146);
xor U26327 (N_26327,N_20369,N_20215);
or U26328 (N_26328,N_24023,N_22977);
and U26329 (N_26329,N_21193,N_20143);
or U26330 (N_26330,N_20009,N_20217);
nor U26331 (N_26331,N_24815,N_23395);
nor U26332 (N_26332,N_21480,N_24572);
or U26333 (N_26333,N_21694,N_21211);
nor U26334 (N_26334,N_24765,N_24625);
or U26335 (N_26335,N_24488,N_21352);
nor U26336 (N_26336,N_24805,N_22987);
or U26337 (N_26337,N_23893,N_21974);
xor U26338 (N_26338,N_22341,N_23062);
xnor U26339 (N_26339,N_21820,N_22441);
nor U26340 (N_26340,N_20284,N_22095);
nand U26341 (N_26341,N_20925,N_20736);
nor U26342 (N_26342,N_23560,N_22883);
nor U26343 (N_26343,N_20286,N_23078);
nand U26344 (N_26344,N_20564,N_21237);
xor U26345 (N_26345,N_21180,N_24717);
or U26346 (N_26346,N_23499,N_23090);
nor U26347 (N_26347,N_21291,N_22786);
or U26348 (N_26348,N_21962,N_23146);
nor U26349 (N_26349,N_24411,N_22113);
nand U26350 (N_26350,N_21825,N_21646);
nor U26351 (N_26351,N_23753,N_23907);
and U26352 (N_26352,N_24803,N_23839);
xor U26353 (N_26353,N_21551,N_21808);
nor U26354 (N_26354,N_21313,N_21454);
or U26355 (N_26355,N_22689,N_24095);
and U26356 (N_26356,N_20279,N_24990);
nor U26357 (N_26357,N_24511,N_22864);
nand U26358 (N_26358,N_23132,N_21465);
or U26359 (N_26359,N_23787,N_23241);
and U26360 (N_26360,N_24810,N_24646);
nand U26361 (N_26361,N_20380,N_21360);
and U26362 (N_26362,N_23693,N_23666);
and U26363 (N_26363,N_23975,N_20663);
nor U26364 (N_26364,N_20664,N_24272);
and U26365 (N_26365,N_22594,N_22425);
nor U26366 (N_26366,N_24718,N_23992);
nor U26367 (N_26367,N_22920,N_23004);
or U26368 (N_26368,N_22380,N_24031);
or U26369 (N_26369,N_22909,N_23925);
nand U26370 (N_26370,N_24930,N_24831);
and U26371 (N_26371,N_22661,N_20059);
or U26372 (N_26372,N_23150,N_23960);
nor U26373 (N_26373,N_21922,N_24832);
xor U26374 (N_26374,N_23802,N_20434);
and U26375 (N_26375,N_24480,N_24381);
and U26376 (N_26376,N_24460,N_21800);
nand U26377 (N_26377,N_20529,N_20381);
and U26378 (N_26378,N_22906,N_20115);
or U26379 (N_26379,N_22750,N_22359);
nand U26380 (N_26380,N_24918,N_24037);
nand U26381 (N_26381,N_22350,N_24741);
xor U26382 (N_26382,N_22395,N_20240);
or U26383 (N_26383,N_22162,N_23598);
xor U26384 (N_26384,N_24995,N_23373);
nor U26385 (N_26385,N_22557,N_22637);
nor U26386 (N_26386,N_20141,N_22029);
nor U26387 (N_26387,N_20575,N_24107);
or U26388 (N_26388,N_21870,N_20263);
and U26389 (N_26389,N_22712,N_24595);
or U26390 (N_26390,N_23968,N_21977);
and U26391 (N_26391,N_20770,N_24201);
nor U26392 (N_26392,N_20624,N_22072);
nand U26393 (N_26393,N_24917,N_24968);
nor U26394 (N_26394,N_20491,N_20842);
nand U26395 (N_26395,N_23795,N_20264);
or U26396 (N_26396,N_20133,N_22931);
or U26397 (N_26397,N_22010,N_21615);
nor U26398 (N_26398,N_24599,N_21381);
nand U26399 (N_26399,N_23069,N_20165);
nor U26400 (N_26400,N_23354,N_20097);
nand U26401 (N_26401,N_24683,N_20250);
nand U26402 (N_26402,N_21011,N_22132);
nor U26403 (N_26403,N_22985,N_20142);
and U26404 (N_26404,N_23415,N_21691);
or U26405 (N_26405,N_21396,N_22462);
xor U26406 (N_26406,N_20731,N_20926);
nand U26407 (N_26407,N_24204,N_23468);
nand U26408 (N_26408,N_20315,N_20618);
xnor U26409 (N_26409,N_21749,N_20087);
nand U26410 (N_26410,N_21787,N_21306);
nand U26411 (N_26411,N_23823,N_21449);
and U26412 (N_26412,N_21331,N_23361);
or U26413 (N_26413,N_21307,N_20163);
or U26414 (N_26414,N_22953,N_20653);
or U26415 (N_26415,N_21341,N_22708);
xnor U26416 (N_26416,N_23278,N_24195);
and U26417 (N_26417,N_22666,N_22588);
and U26418 (N_26418,N_23651,N_21069);
nor U26419 (N_26419,N_20010,N_21692);
nand U26420 (N_26420,N_24690,N_22310);
nor U26421 (N_26421,N_21735,N_23538);
nor U26422 (N_26422,N_20803,N_20951);
nor U26423 (N_26423,N_22478,N_22888);
or U26424 (N_26424,N_22202,N_24228);
xnor U26425 (N_26425,N_22826,N_21708);
and U26426 (N_26426,N_24829,N_23323);
and U26427 (N_26427,N_20553,N_23762);
nor U26428 (N_26428,N_21841,N_21208);
and U26429 (N_26429,N_21655,N_24758);
xor U26430 (N_26430,N_22412,N_23145);
or U26431 (N_26431,N_24390,N_24709);
nor U26432 (N_26432,N_21837,N_24658);
xor U26433 (N_26433,N_20440,N_21633);
nor U26434 (N_26434,N_20347,N_23304);
and U26435 (N_26435,N_24243,N_21022);
nor U26436 (N_26436,N_23729,N_20778);
xnor U26437 (N_26437,N_20425,N_21478);
or U26438 (N_26438,N_24673,N_23793);
and U26439 (N_26439,N_24517,N_24330);
or U26440 (N_26440,N_23490,N_23016);
xor U26441 (N_26441,N_22082,N_20064);
nor U26442 (N_26442,N_24760,N_21622);
or U26443 (N_26443,N_24819,N_23509);
or U26444 (N_26444,N_21647,N_23159);
nor U26445 (N_26445,N_22692,N_22281);
nand U26446 (N_26446,N_24877,N_24833);
or U26447 (N_26447,N_22379,N_24173);
or U26448 (N_26448,N_22770,N_23590);
nand U26449 (N_26449,N_24125,N_20372);
nand U26450 (N_26450,N_24067,N_21346);
or U26451 (N_26451,N_21264,N_23985);
and U26452 (N_26452,N_21423,N_23746);
or U26453 (N_26453,N_22706,N_22378);
and U26454 (N_26454,N_24441,N_24476);
nand U26455 (N_26455,N_21451,N_22738);
or U26456 (N_26456,N_20297,N_20965);
nand U26457 (N_26457,N_20591,N_21310);
or U26458 (N_26458,N_23919,N_21980);
or U26459 (N_26459,N_20635,N_20833);
or U26460 (N_26460,N_20208,N_20450);
and U26461 (N_26461,N_22993,N_22928);
xnor U26462 (N_26462,N_20840,N_22087);
or U26463 (N_26463,N_23683,N_20057);
xor U26464 (N_26464,N_24492,N_20550);
and U26465 (N_26465,N_23979,N_20071);
nor U26466 (N_26466,N_23269,N_20984);
nor U26467 (N_26467,N_20643,N_23060);
xnor U26468 (N_26468,N_21818,N_21403);
nand U26469 (N_26469,N_22763,N_21244);
nand U26470 (N_26470,N_21177,N_24608);
nand U26471 (N_26471,N_24669,N_23922);
or U26472 (N_26472,N_24034,N_24695);
nand U26473 (N_26473,N_23092,N_24137);
nand U26474 (N_26474,N_20672,N_21215);
nor U26475 (N_26475,N_24048,N_24055);
nor U26476 (N_26476,N_24165,N_23186);
or U26477 (N_26477,N_23958,N_21618);
nor U26478 (N_26478,N_20839,N_23479);
or U26479 (N_26479,N_21008,N_21383);
xnor U26480 (N_26480,N_21189,N_23534);
or U26481 (N_26481,N_21104,N_20005);
or U26482 (N_26482,N_20837,N_20871);
and U26483 (N_26483,N_24349,N_22655);
nor U26484 (N_26484,N_20175,N_21010);
nor U26485 (N_26485,N_23068,N_23737);
and U26486 (N_26486,N_22479,N_20266);
xnor U26487 (N_26487,N_23402,N_24298);
nor U26488 (N_26488,N_20707,N_22070);
nor U26489 (N_26489,N_21733,N_24124);
xor U26490 (N_26490,N_20706,N_22533);
nor U26491 (N_26491,N_23535,N_20562);
nand U26492 (N_26492,N_21630,N_20867);
xor U26493 (N_26493,N_21976,N_20455);
nand U26494 (N_26494,N_20792,N_21624);
and U26495 (N_26495,N_23258,N_22054);
nor U26496 (N_26496,N_20386,N_22266);
xnor U26497 (N_26497,N_24051,N_23794);
nand U26498 (N_26498,N_24404,N_23151);
nand U26499 (N_26499,N_24609,N_20060);
or U26500 (N_26500,N_22245,N_24754);
nand U26501 (N_26501,N_21779,N_23045);
or U26502 (N_26502,N_24984,N_21332);
nor U26503 (N_26503,N_23335,N_23592);
and U26504 (N_26504,N_21064,N_22220);
nand U26505 (N_26505,N_22265,N_23632);
nand U26506 (N_26506,N_24723,N_24559);
or U26507 (N_26507,N_21247,N_21163);
or U26508 (N_26508,N_20662,N_20129);
nor U26509 (N_26509,N_24519,N_22560);
or U26510 (N_26510,N_24057,N_22451);
and U26511 (N_26511,N_23769,N_21896);
xnor U26512 (N_26512,N_22389,N_23251);
nand U26513 (N_26513,N_24996,N_22716);
xnor U26514 (N_26514,N_24965,N_20970);
nor U26515 (N_26515,N_24281,N_24696);
xor U26516 (N_26516,N_24017,N_23977);
xnor U26517 (N_26517,N_21526,N_20421);
and U26518 (N_26518,N_21746,N_21115);
or U26519 (N_26519,N_20187,N_20845);
or U26520 (N_26520,N_24345,N_22422);
xor U26521 (N_26521,N_21947,N_21419);
or U26522 (N_26522,N_22052,N_24334);
and U26523 (N_26523,N_21496,N_23845);
xnor U26524 (N_26524,N_22295,N_20942);
nor U26525 (N_26525,N_20937,N_22313);
nand U26526 (N_26526,N_22292,N_24307);
nor U26527 (N_26527,N_20153,N_21925);
and U26528 (N_26528,N_22440,N_22390);
or U26529 (N_26529,N_20244,N_24241);
xnor U26530 (N_26530,N_21829,N_20812);
or U26531 (N_26531,N_23331,N_21195);
nand U26532 (N_26532,N_21569,N_22349);
nand U26533 (N_26533,N_24681,N_21715);
nor U26534 (N_26534,N_20769,N_24787);
nand U26535 (N_26535,N_20955,N_21991);
and U26536 (N_26536,N_22322,N_20990);
and U26537 (N_26537,N_20713,N_24564);
nor U26538 (N_26538,N_23253,N_24677);
xnor U26539 (N_26539,N_21424,N_24628);
nand U26540 (N_26540,N_20825,N_20135);
or U26541 (N_26541,N_21594,N_23473);
nand U26542 (N_26542,N_24280,N_24620);
or U26543 (N_26543,N_24318,N_22873);
and U26544 (N_26544,N_20988,N_20884);
xnor U26545 (N_26545,N_21616,N_20720);
nand U26546 (N_26546,N_23281,N_22250);
or U26547 (N_26547,N_22975,N_22251);
and U26548 (N_26548,N_24848,N_20346);
and U26549 (N_26549,N_22924,N_24391);
xor U26550 (N_26550,N_22687,N_20929);
nor U26551 (N_26551,N_22067,N_22455);
xor U26552 (N_26552,N_20356,N_22589);
or U26553 (N_26553,N_21942,N_20613);
nand U26554 (N_26554,N_24297,N_24016);
or U26555 (N_26555,N_23928,N_22414);
nand U26556 (N_26556,N_23377,N_23120);
and U26557 (N_26557,N_21743,N_21096);
xnor U26558 (N_26558,N_23427,N_21948);
and U26559 (N_26559,N_21511,N_22683);
xor U26560 (N_26560,N_22410,N_21099);
xnor U26561 (N_26561,N_24430,N_21493);
nor U26562 (N_26562,N_21685,N_23048);
or U26563 (N_26563,N_22868,N_23770);
nand U26564 (N_26564,N_23440,N_21037);
xor U26565 (N_26565,N_21474,N_21216);
or U26566 (N_26566,N_21605,N_22849);
nor U26567 (N_26567,N_22229,N_21728);
or U26568 (N_26568,N_23198,N_21750);
and U26569 (N_26569,N_21086,N_23900);
and U26570 (N_26570,N_22206,N_23984);
and U26571 (N_26571,N_24266,N_22334);
and U26572 (N_26572,N_21516,N_22525);
xnor U26573 (N_26573,N_23988,N_20260);
xor U26574 (N_26574,N_21906,N_20363);
and U26575 (N_26575,N_20111,N_22392);
and U26576 (N_26576,N_21063,N_24617);
xnor U26577 (N_26577,N_24174,N_24693);
or U26578 (N_26578,N_24273,N_24618);
nor U26579 (N_26579,N_21443,N_20176);
or U26580 (N_26580,N_21337,N_22421);
xor U26581 (N_26581,N_24910,N_20992);
nand U26582 (N_26582,N_21603,N_21223);
nor U26583 (N_26583,N_22017,N_20231);
nor U26584 (N_26584,N_21348,N_23739);
xor U26585 (N_26585,N_21626,N_23476);
nand U26586 (N_26586,N_20245,N_22815);
xnor U26587 (N_26587,N_22435,N_22592);
nand U26588 (N_26588,N_20599,N_21400);
or U26589 (N_26589,N_22420,N_23650);
or U26590 (N_26590,N_22915,N_22028);
nor U26591 (N_26591,N_22044,N_21819);
or U26592 (N_26592,N_20790,N_23434);
or U26593 (N_26593,N_21434,N_23881);
xor U26594 (N_26594,N_23383,N_24458);
nand U26595 (N_26595,N_21196,N_23074);
nand U26596 (N_26596,N_24738,N_23617);
xor U26597 (N_26597,N_23503,N_23822);
nand U26598 (N_26598,N_23609,N_22493);
or U26599 (N_26599,N_22948,N_23381);
and U26600 (N_26600,N_21772,N_21284);
and U26601 (N_26601,N_21989,N_24748);
or U26602 (N_26602,N_23023,N_23363);
nor U26603 (N_26603,N_20160,N_24333);
nand U26604 (N_26604,N_22511,N_21351);
nor U26605 (N_26605,N_21704,N_20483);
xor U26606 (N_26606,N_20836,N_22002);
and U26607 (N_26607,N_21753,N_20033);
xor U26608 (N_26608,N_24499,N_23704);
xnor U26609 (N_26609,N_24092,N_23537);
nor U26610 (N_26610,N_20461,N_22242);
nor U26611 (N_26611,N_20758,N_22284);
and U26612 (N_26612,N_24969,N_20276);
and U26613 (N_26613,N_24359,N_22633);
xor U26614 (N_26614,N_23616,N_23008);
and U26615 (N_26615,N_23332,N_21875);
nor U26616 (N_26616,N_20271,N_21731);
xnor U26617 (N_26617,N_22026,N_21623);
and U26618 (N_26618,N_22060,N_24823);
or U26619 (N_26619,N_20649,N_23393);
and U26620 (N_26620,N_23097,N_21506);
nor U26621 (N_26621,N_21560,N_22209);
nor U26622 (N_26622,N_23849,N_23662);
or U26623 (N_26623,N_21460,N_22298);
or U26624 (N_26624,N_20283,N_22048);
xnor U26625 (N_26625,N_21548,N_21045);
or U26626 (N_26626,N_20554,N_20389);
and U26627 (N_26627,N_23011,N_24641);
nor U26628 (N_26628,N_20220,N_24880);
xor U26629 (N_26629,N_22473,N_24169);
nor U26630 (N_26630,N_20099,N_23461);
or U26631 (N_26631,N_22919,N_20650);
nand U26632 (N_26632,N_22367,N_22718);
nand U26633 (N_26633,N_23660,N_20555);
and U26634 (N_26634,N_24707,N_21060);
xor U26635 (N_26635,N_24583,N_23603);
xor U26636 (N_26636,N_21389,N_22590);
nand U26637 (N_26637,N_20408,N_21515);
nand U26638 (N_26638,N_20361,N_21487);
nand U26639 (N_26639,N_23639,N_21082);
nand U26640 (N_26640,N_23721,N_20330);
and U26641 (N_26641,N_21482,N_22745);
xor U26642 (N_26642,N_21058,N_22709);
nor U26643 (N_26643,N_24142,N_24449);
and U26644 (N_26644,N_24900,N_22025);
nand U26645 (N_26645,N_21207,N_22719);
and U26646 (N_26646,N_23277,N_23970);
nor U26647 (N_26647,N_21960,N_22357);
or U26648 (N_26648,N_22777,N_24736);
and U26649 (N_26649,N_21627,N_20011);
or U26650 (N_26650,N_23887,N_20614);
nand U26651 (N_26651,N_21055,N_22297);
or U26652 (N_26652,N_20339,N_24947);
nand U26653 (N_26653,N_24751,N_24587);
nor U26654 (N_26654,N_22001,N_21065);
or U26655 (N_26655,N_24198,N_22151);
xnor U26656 (N_26656,N_21407,N_24852);
nand U26657 (N_26657,N_24536,N_22880);
and U26658 (N_26658,N_21843,N_24340);
nand U26659 (N_26659,N_23707,N_22019);
and U26660 (N_26660,N_22648,N_21919);
nor U26661 (N_26661,N_22989,N_23392);
nor U26662 (N_26662,N_21268,N_22829);
xor U26663 (N_26663,N_20124,N_21367);
xnor U26664 (N_26664,N_23848,N_22675);
nor U26665 (N_26665,N_21111,N_23917);
nor U26666 (N_26666,N_21035,N_22007);
nand U26667 (N_26667,N_21285,N_20441);
and U26668 (N_26668,N_22419,N_23959);
nand U26669 (N_26669,N_23784,N_20816);
nor U26670 (N_26670,N_20255,N_24578);
xnor U26671 (N_26671,N_21642,N_23441);
xnor U26672 (N_26672,N_23630,N_24088);
nor U26673 (N_26673,N_22382,N_20580);
and U26674 (N_26674,N_21466,N_22207);
xnor U26675 (N_26675,N_20261,N_20828);
xnor U26676 (N_26676,N_23832,N_24664);
and U26677 (N_26677,N_22601,N_24619);
and U26678 (N_26678,N_23156,N_24256);
nand U26679 (N_26679,N_24079,N_20722);
nor U26680 (N_26680,N_21298,N_24633);
xnor U26681 (N_26681,N_22945,N_21019);
or U26682 (N_26682,N_23706,N_24961);
nor U26683 (N_26683,N_21898,N_20331);
xnor U26684 (N_26684,N_24638,N_20526);
nor U26685 (N_26685,N_24444,N_23431);
xor U26686 (N_26686,N_23170,N_23098);
xor U26687 (N_26687,N_24992,N_20888);
xnor U26688 (N_26688,N_24860,N_22042);
and U26689 (N_26689,N_22051,N_21470);
and U26690 (N_26690,N_22385,N_22384);
or U26691 (N_26691,N_23022,N_22180);
nand U26692 (N_26692,N_24907,N_24043);
xnor U26693 (N_26693,N_21239,N_21136);
nand U26694 (N_26694,N_20680,N_24021);
xnor U26695 (N_26695,N_20498,N_20505);
or U26696 (N_26696,N_24111,N_22726);
or U26697 (N_26697,N_23210,N_22865);
and U26698 (N_26698,N_22595,N_20140);
xnor U26699 (N_26699,N_20026,N_24560);
or U26700 (N_26700,N_22978,N_20469);
xor U26701 (N_26701,N_24778,N_20118);
nor U26702 (N_26702,N_24821,N_22203);
nor U26703 (N_26703,N_23494,N_22737);
xor U26704 (N_26704,N_23265,N_22488);
and U26705 (N_26705,N_22761,N_23465);
xor U26706 (N_26706,N_21850,N_22863);
nor U26707 (N_26707,N_24871,N_21902);
xnor U26708 (N_26708,N_24191,N_24443);
xor U26709 (N_26709,N_23454,N_22430);
and U26710 (N_26710,N_20134,N_22061);
nor U26711 (N_26711,N_24178,N_22736);
nand U26712 (N_26712,N_21959,N_24621);
nor U26713 (N_26713,N_23643,N_20144);
or U26714 (N_26714,N_23542,N_21760);
xor U26715 (N_26715,N_20597,N_24072);
xnor U26716 (N_26716,N_24637,N_23273);
nand U26717 (N_26717,N_22300,N_20734);
or U26718 (N_26718,N_23366,N_21751);
xnor U26719 (N_26719,N_21414,N_21789);
xnor U26720 (N_26720,N_20216,N_23751);
or U26721 (N_26721,N_20150,N_20607);
xnor U26722 (N_26722,N_24960,N_20293);
or U26723 (N_26723,N_22210,N_22311);
xnor U26724 (N_26724,N_23288,N_22650);
and U26725 (N_26725,N_24235,N_21471);
and U26726 (N_26726,N_24461,N_23602);
or U26727 (N_26727,N_20467,N_21640);
nor U26728 (N_26728,N_22917,N_20901);
or U26729 (N_26729,N_21228,N_23843);
nor U26730 (N_26730,N_20410,N_21790);
nor U26731 (N_26731,N_23386,N_24959);
xnor U26732 (N_26732,N_22779,N_20761);
xor U26733 (N_26733,N_22602,N_24510);
xnor U26734 (N_26734,N_20592,N_23437);
and U26735 (N_26735,N_22713,N_23736);
nand U26736 (N_26736,N_21696,N_21740);
xor U26737 (N_26737,N_23781,N_23412);
or U26738 (N_26738,N_21088,N_21003);
xnor U26739 (N_26739,N_23568,N_24289);
and U26740 (N_26740,N_22227,N_24911);
xnor U26741 (N_26741,N_22021,N_22539);
xnor U26742 (N_26742,N_20544,N_22760);
or U26743 (N_26743,N_20341,N_22122);
and U26744 (N_26744,N_24205,N_22854);
or U26745 (N_26745,N_21355,N_20659);
and U26746 (N_26746,N_21344,N_20400);
and U26747 (N_26747,N_23909,N_20233);
or U26748 (N_26748,N_20398,N_24853);
or U26749 (N_26749,N_24450,N_22891);
nor U26750 (N_26750,N_23356,N_22416);
nor U26751 (N_26751,N_20773,N_20445);
nor U26752 (N_26752,N_22348,N_21107);
xnor U26753 (N_26753,N_23789,N_22426);
or U26754 (N_26754,N_20869,N_22449);
nand U26755 (N_26755,N_21320,N_23498);
and U26756 (N_26756,N_21273,N_21877);
nand U26757 (N_26757,N_20541,N_23931);
nor U26758 (N_26758,N_20159,N_23404);
or U26759 (N_26759,N_22547,N_20835);
xor U26760 (N_26760,N_21943,N_23573);
nor U26761 (N_26761,N_23775,N_20697);
nand U26762 (N_26762,N_23719,N_21447);
xnor U26763 (N_26763,N_20222,N_23815);
xnor U26764 (N_26764,N_24855,N_23757);
nor U26765 (N_26765,N_20881,N_21275);
xnor U26766 (N_26766,N_23497,N_22870);
or U26767 (N_26767,N_20795,N_20856);
nand U26768 (N_26768,N_22969,N_21734);
nand U26769 (N_26769,N_21939,N_24096);
nor U26770 (N_26770,N_21668,N_23401);
or U26771 (N_26771,N_20084,N_21584);
nand U26772 (N_26772,N_24784,N_22930);
nand U26773 (N_26773,N_21440,N_22811);
nand U26774 (N_26774,N_23733,N_23379);
and U26775 (N_26775,N_22732,N_20987);
nand U26776 (N_26776,N_22080,N_24187);
nor U26777 (N_26777,N_23206,N_20695);
and U26778 (N_26778,N_21670,N_20125);
nand U26779 (N_26779,N_23936,N_21531);
or U26780 (N_26780,N_20035,N_23935);
nor U26781 (N_26781,N_24818,N_24147);
and U26782 (N_26782,N_20685,N_20403);
and U26783 (N_26783,N_22839,N_21988);
or U26784 (N_26784,N_24520,N_20559);
or U26785 (N_26785,N_20174,N_20646);
and U26786 (N_26786,N_24301,N_21083);
nor U26787 (N_26787,N_23347,N_21730);
and U26788 (N_26788,N_20982,N_23678);
or U26789 (N_26789,N_23310,N_22665);
xor U26790 (N_26790,N_24851,N_23567);
xor U26791 (N_26791,N_21459,N_23672);
and U26792 (N_26792,N_20229,N_24153);
or U26793 (N_26793,N_20598,N_23272);
and U26794 (N_26794,N_20322,N_24103);
nor U26795 (N_26795,N_22555,N_23484);
or U26796 (N_26796,N_22810,N_20136);
and U26797 (N_26797,N_23291,N_22117);
and U26798 (N_26798,N_22639,N_23516);
xnor U26799 (N_26799,N_22604,N_24576);
nor U26800 (N_26800,N_22436,N_22694);
or U26801 (N_26801,N_24020,N_21317);
and U26802 (N_26802,N_22116,N_22698);
nand U26803 (N_26803,N_23038,N_24127);
and U26804 (N_26804,N_23808,N_24433);
nand U26805 (N_26805,N_24268,N_23102);
or U26806 (N_26806,N_23502,N_20272);
nand U26807 (N_26807,N_20589,N_22189);
or U26808 (N_26808,N_23697,N_24753);
nand U26809 (N_26809,N_22960,N_24073);
nor U26810 (N_26810,N_21732,N_20417);
xnor U26811 (N_26811,N_21007,N_23718);
nand U26812 (N_26812,N_20788,N_24255);
and U26813 (N_26813,N_22916,N_20682);
or U26814 (N_26814,N_24400,N_21577);
and U26815 (N_26815,N_24936,N_23229);
nand U26816 (N_26816,N_21625,N_20757);
nand U26817 (N_26817,N_21579,N_23546);
nor U26818 (N_26818,N_22164,N_23825);
xnor U26819 (N_26819,N_20457,N_23561);
and U26820 (N_26820,N_20170,N_23298);
and U26821 (N_26821,N_20114,N_22418);
and U26822 (N_26822,N_24007,N_20237);
or U26823 (N_26823,N_21404,N_24776);
and U26824 (N_26824,N_21547,N_20508);
nor U26825 (N_26825,N_24004,N_23483);
xor U26826 (N_26826,N_20834,N_20615);
or U26827 (N_26827,N_22050,N_20547);
nand U26828 (N_26828,N_23562,N_22224);
nor U26829 (N_26829,N_21953,N_24987);
nand U26830 (N_26830,N_24489,N_23162);
xor U26831 (N_26831,N_24014,N_22680);
xnor U26832 (N_26832,N_23864,N_24557);
nor U26833 (N_26833,N_20023,N_21079);
xor U26834 (N_26834,N_21077,N_20717);
nor U26835 (N_26835,N_21141,N_21855);
or U26836 (N_26836,N_20053,N_22672);
nand U26837 (N_26837,N_23910,N_23111);
xor U26838 (N_26838,N_23106,N_20355);
nand U26839 (N_26839,N_23025,N_21589);
xor U26840 (N_26840,N_23955,N_21659);
nor U26841 (N_26841,N_24013,N_24697);
nor U26842 (N_26842,N_22360,N_24822);
xnor U26843 (N_26843,N_23239,N_24314);
xor U26844 (N_26844,N_21853,N_23342);
or U26845 (N_26845,N_20802,N_20476);
nand U26846 (N_26846,N_22417,N_24988);
xnor U26847 (N_26847,N_22828,N_20181);
and U26848 (N_26848,N_22973,N_23634);
and U26849 (N_26849,N_22335,N_24545);
and U26850 (N_26850,N_23348,N_20326);
nand U26851 (N_26851,N_20340,N_20941);
nand U26852 (N_26852,N_24579,N_24602);
nor U26853 (N_26853,N_24976,N_21078);
and U26854 (N_26854,N_22895,N_21983);
or U26855 (N_26855,N_24710,N_20604);
nor U26856 (N_26856,N_20919,N_21125);
nor U26857 (N_26857,N_22346,N_24940);
or U26858 (N_26858,N_22338,N_24224);
xor U26859 (N_26859,N_23220,N_23359);
nor U26860 (N_26860,N_24565,N_23457);
and U26861 (N_26861,N_23071,N_22327);
xnor U26862 (N_26862,N_23741,N_22842);
nand U26863 (N_26863,N_23445,N_20913);
nor U26864 (N_26864,N_21199,N_20651);
and U26865 (N_26865,N_20946,N_23000);
or U26866 (N_26866,N_24632,N_22354);
nand U26867 (N_26867,N_21690,N_22814);
and U26868 (N_26868,N_22962,N_23271);
nor U26869 (N_26869,N_23443,N_23874);
nand U26870 (N_26870,N_24484,N_23302);
nor U26871 (N_26871,N_21322,N_24324);
nor U26872 (N_26872,N_20344,N_24502);
xor U26873 (N_26873,N_22034,N_20239);
nand U26874 (N_26874,N_21036,N_23144);
and U26875 (N_26875,N_21140,N_22992);
or U26876 (N_26876,N_23940,N_24239);
and U26877 (N_26877,N_23659,N_21427);
xor U26878 (N_26878,N_23181,N_21303);
nand U26879 (N_26879,N_22721,N_21292);
nand U26880 (N_26880,N_20863,N_22562);
nor U26881 (N_26881,N_20107,N_20019);
xor U26882 (N_26882,N_21334,N_23125);
nor U26883 (N_26883,N_20981,N_21931);
and U26884 (N_26884,N_22860,N_21768);
and U26885 (N_26885,N_24149,N_22669);
nor U26886 (N_26886,N_22465,N_21651);
and U26887 (N_26887,N_24338,N_22239);
or U26888 (N_26888,N_21200,N_20944);
nand U26889 (N_26889,N_21944,N_23601);
xnor U26890 (N_26890,N_21249,N_23425);
or U26891 (N_26891,N_20139,N_23204);
nor U26892 (N_26892,N_21540,N_21973);
nor U26893 (N_26893,N_22876,N_24478);
xor U26894 (N_26894,N_20782,N_22531);
xor U26895 (N_26895,N_22974,N_24543);
or U26896 (N_26896,N_20800,N_24084);
nor U26897 (N_26897,N_23623,N_24862);
or U26898 (N_26898,N_20652,N_23187);
nor U26899 (N_26899,N_24590,N_20914);
nand U26900 (N_26900,N_23637,N_21815);
or U26901 (N_26901,N_23576,N_20733);
xnor U26902 (N_26902,N_20311,N_24445);
and U26903 (N_26903,N_22813,N_22259);
and U26904 (N_26904,N_20519,N_21879);
xor U26905 (N_26905,N_20979,N_20811);
and U26906 (N_26906,N_20771,N_21039);
or U26907 (N_26907,N_22302,N_24424);
xnor U26908 (N_26908,N_22218,N_23217);
xnor U26909 (N_26909,N_20366,N_21778);
xor U26910 (N_26910,N_21507,N_21448);
or U26911 (N_26911,N_21130,N_24861);
nor U26912 (N_26912,N_21167,N_21349);
or U26913 (N_26913,N_22144,N_21710);
and U26914 (N_26914,N_24522,N_20977);
nand U26915 (N_26915,N_21316,N_20443);
nor U26916 (N_26916,N_21664,N_22515);
nand U26917 (N_26917,N_23477,N_21391);
or U26918 (N_26918,N_22328,N_20449);
xor U26919 (N_26919,N_23991,N_20480);
xor U26920 (N_26920,N_24284,N_24714);
or U26921 (N_26921,N_22808,N_21876);
nand U26922 (N_26922,N_23311,N_24972);
nand U26923 (N_26923,N_23054,N_23600);
and U26924 (N_26924,N_21067,N_20428);
or U26925 (N_26925,N_24473,N_22774);
or U26926 (N_26926,N_21836,N_24931);
nand U26927 (N_26927,N_21347,N_22538);
or U26928 (N_26928,N_20225,N_20391);
and U26929 (N_26929,N_22086,N_21397);
nand U26930 (N_26930,N_22528,N_24429);
nand U26931 (N_26931,N_24019,N_22972);
xnor U26932 (N_26932,N_23055,N_22834);
or U26933 (N_26933,N_23575,N_24250);
nor U26934 (N_26934,N_22964,N_22365);
nor U26935 (N_26935,N_20246,N_22091);
nand U26936 (N_26936,N_23037,N_22475);
nor U26937 (N_26937,N_22982,N_20288);
or U26938 (N_26938,N_22375,N_23020);
xnor U26939 (N_26939,N_20523,N_22657);
and U26940 (N_26940,N_23711,N_20198);
xor U26941 (N_26941,N_24485,N_22996);
xor U26942 (N_26942,N_21712,N_22178);
xnor U26943 (N_26943,N_21034,N_21134);
xnor U26944 (N_26944,N_24210,N_24108);
or U26945 (N_26945,N_21229,N_24431);
or U26946 (N_26946,N_21629,N_22211);
and U26947 (N_26947,N_24181,N_20007);
and U26948 (N_26948,N_20046,N_20909);
and U26949 (N_26949,N_21620,N_24259);
and U26950 (N_26950,N_21830,N_21890);
and U26951 (N_26951,N_22780,N_22232);
xnor U26952 (N_26952,N_20466,N_20236);
xnor U26953 (N_26953,N_23621,N_21783);
nand U26954 (N_26954,N_24388,N_20074);
or U26955 (N_26955,N_23965,N_22831);
nand U26956 (N_26956,N_21874,N_21774);
or U26957 (N_26957,N_20777,N_21308);
or U26958 (N_26958,N_22678,N_23072);
nand U26959 (N_26959,N_21669,N_24515);
and U26960 (N_26960,N_22702,N_24357);
or U26961 (N_26961,N_20478,N_24606);
xnor U26962 (N_26962,N_24932,N_23776);
or U26963 (N_26963,N_20516,N_20625);
nor U26964 (N_26964,N_20210,N_21665);
and U26965 (N_26965,N_21543,N_22272);
xnor U26966 (N_26966,N_23525,N_23053);
xnor U26967 (N_26967,N_23805,N_22123);
nor U26968 (N_26968,N_22656,N_21544);
xnor U26969 (N_26969,N_22155,N_20775);
xor U26970 (N_26970,N_20195,N_20958);
xnor U26971 (N_26971,N_22120,N_20093);
xor U26972 (N_26972,N_20397,N_24302);
nand U26973 (N_26973,N_24036,N_24603);
nor U26974 (N_26974,N_23158,N_21978);
and U26975 (N_26975,N_23976,N_24331);
or U26976 (N_26976,N_24659,N_22447);
nor U26977 (N_26977,N_24856,N_24186);
and U26978 (N_26978,N_21015,N_24897);
nor U26979 (N_26979,N_22443,N_24277);
nand U26980 (N_26980,N_21131,N_21593);
nand U26981 (N_26981,N_24915,N_24344);
and U26982 (N_26982,N_20566,N_23532);
nor U26983 (N_26983,N_20048,N_22787);
nand U26984 (N_26984,N_24844,N_21345);
and U26985 (N_26985,N_22233,N_24361);
or U26986 (N_26986,N_22102,N_23398);
nand U26987 (N_26987,N_24670,N_20963);
or U26988 (N_26988,N_20367,N_20959);
and U26989 (N_26989,N_21621,N_22504);
and U26990 (N_26990,N_20147,N_24812);
or U26991 (N_26991,N_21489,N_24729);
nand U26992 (N_26992,N_23572,N_20076);
or U26993 (N_26993,N_24022,N_22285);
nand U26994 (N_26994,N_20603,N_21158);
and U26995 (N_26995,N_23791,N_24054);
nor U26996 (N_26996,N_23073,N_22270);
nor U26997 (N_26997,N_23648,N_20377);
xnor U26998 (N_26998,N_23837,N_22725);
xnor U26999 (N_26999,N_22575,N_21497);
nor U27000 (N_27000,N_22957,N_23070);
nor U27001 (N_27001,N_22711,N_20287);
xor U27002 (N_27002,N_23408,N_24542);
nor U27003 (N_27003,N_22671,N_24631);
xor U27004 (N_27004,N_20621,N_24398);
nand U27005 (N_27005,N_21226,N_23179);
xnor U27006 (N_27006,N_24890,N_22182);
or U27007 (N_27007,N_24120,N_23824);
nand U27008 (N_27008,N_22053,N_22402);
nor U27009 (N_27009,N_20034,N_22063);
nor U27010 (N_27010,N_22183,N_20787);
and U27011 (N_27011,N_21425,N_22674);
nor U27012 (N_27012,N_23242,N_20565);
nand U27013 (N_27013,N_24558,N_24086);
xnor U27014 (N_27014,N_20626,N_24214);
nor U27015 (N_27015,N_22990,N_22503);
nor U27016 (N_27016,N_24728,N_22530);
xnor U27017 (N_27017,N_23918,N_20865);
xnor U27018 (N_27018,N_21641,N_23728);
or U27019 (N_27019,N_21766,N_21012);
nor U27020 (N_27020,N_20452,N_20383);
or U27021 (N_27021,N_22316,N_22502);
and U27022 (N_27022,N_21645,N_20739);
xor U27023 (N_27023,N_22558,N_23750);
or U27024 (N_27024,N_24315,N_24341);
nand U27025 (N_27025,N_24850,N_20766);
or U27026 (N_27026,N_23510,N_22620);
nor U27027 (N_27027,N_23840,N_23221);
or U27028 (N_27028,N_24212,N_24566);
or U27029 (N_27029,N_24665,N_23860);
and U27030 (N_27030,N_23226,N_21289);
nor U27031 (N_27031,N_22512,N_23702);
nor U27032 (N_27032,N_24045,N_21113);
nand U27033 (N_27033,N_21370,N_22016);
xor U27034 (N_27034,N_24490,N_24991);
nor U27035 (N_27035,N_23122,N_21719);
nor U27036 (N_27036,N_21812,N_22758);
nand U27037 (N_27037,N_22468,N_23303);
and U27038 (N_27038,N_21262,N_22035);
xnor U27039 (N_27039,N_24220,N_22851);
or U27040 (N_27040,N_22069,N_22090);
or U27041 (N_27041,N_23200,N_21062);
and U27042 (N_27042,N_20013,N_22812);
nor U27043 (N_27043,N_24497,N_20513);
or U27044 (N_27044,N_21518,N_21100);
and U27045 (N_27045,N_20489,N_23374);
nand U27046 (N_27046,N_23951,N_20581);
xor U27047 (N_27047,N_20121,N_22668);
and U27048 (N_27048,N_20209,N_23663);
nand U27049 (N_27049,N_22368,N_24122);
xor U27050 (N_27050,N_22071,N_20789);
xor U27051 (N_27051,N_20083,N_22778);
or U27052 (N_27052,N_24003,N_23524);
or U27053 (N_27053,N_23260,N_21445);
or U27054 (N_27054,N_21538,N_21755);
xor U27055 (N_27055,N_22772,N_21611);
xor U27056 (N_27056,N_23033,N_20298);
nand U27057 (N_27057,N_20016,N_23763);
xor U27058 (N_27058,N_23333,N_24363);
nand U27059 (N_27059,N_23492,N_23316);
nor U27060 (N_27060,N_21356,N_22517);
xor U27061 (N_27061,N_20228,N_24172);
nor U27062 (N_27062,N_24406,N_20182);
xnor U27063 (N_27063,N_22329,N_20294);
xnor U27064 (N_27064,N_24649,N_24384);
and U27065 (N_27065,N_23290,N_24213);
or U27066 (N_27066,N_20818,N_20521);
or U27067 (N_27067,N_22490,N_24469);
and U27068 (N_27068,N_22951,N_22319);
nor U27069 (N_27069,N_22083,N_24761);
xor U27070 (N_27070,N_22476,N_23557);
nand U27071 (N_27071,N_21699,N_24721);
or U27072 (N_27072,N_24735,N_21637);
or U27073 (N_27073,N_23670,N_24531);
or U27074 (N_27074,N_24061,N_22510);
xnor U27075 (N_27075,N_22246,N_23695);
nand U27076 (N_27076,N_23417,N_22824);
xor U27077 (N_27077,N_23470,N_24377);
nand U27078 (N_27078,N_24464,N_20218);
xor U27079 (N_27079,N_20172,N_22077);
xnor U27080 (N_27080,N_23095,N_21940);
and U27081 (N_27081,N_20105,N_24117);
or U27082 (N_27082,N_20077,N_24688);
or U27083 (N_27083,N_20504,N_20669);
nand U27084 (N_27084,N_21392,N_23932);
nor U27085 (N_27085,N_23536,N_23324);
and U27086 (N_27086,N_23613,N_24419);
xor U27087 (N_27087,N_20933,N_21727);
nor U27088 (N_27088,N_24656,N_22636);
xor U27089 (N_27089,N_24889,N_23261);
xor U27090 (N_27090,N_22396,N_21183);
nand U27091 (N_27091,N_24348,N_20582);
or U27092 (N_27092,N_20281,N_21280);
and U27093 (N_27093,N_22818,N_20642);
xnor U27094 (N_27094,N_20289,N_23469);
and U27095 (N_27095,N_24346,N_24196);
and U27096 (N_27096,N_24221,N_22754);
or U27097 (N_27097,N_23701,N_20805);
and U27098 (N_27098,N_22274,N_20458);
or U27099 (N_27099,N_24337,N_21085);
nand U27100 (N_27100,N_23148,N_23817);
or U27101 (N_27101,N_23197,N_21501);
nand U27102 (N_27102,N_23722,N_23082);
xor U27103 (N_27103,N_23344,N_22875);
and U27104 (N_27104,N_22277,N_21432);
or U27105 (N_27105,N_20684,N_21452);
nor U27106 (N_27106,N_24325,N_20470);
nor U27107 (N_27107,N_20917,N_22057);
nand U27108 (N_27108,N_22591,N_20573);
and U27109 (N_27109,N_20102,N_20273);
xor U27110 (N_27110,N_20693,N_24496);
and U27111 (N_27111,N_20179,N_24757);
nand U27112 (N_27112,N_22579,N_24132);
and U27113 (N_27113,N_20827,N_21318);
nor U27114 (N_27114,N_20430,N_23464);
nand U27115 (N_27115,N_22550,N_21056);
nand U27116 (N_27116,N_23858,N_21312);
and U27117 (N_27117,N_24691,N_24574);
xnor U27118 (N_27118,N_21517,N_24358);
xor U27119 (N_27119,N_23774,N_22143);
nor U27120 (N_27120,N_24459,N_23485);
nor U27121 (N_27121,N_24623,N_23387);
or U27122 (N_27122,N_21435,N_24479);
nand U27123 (N_27123,N_24066,N_24170);
or U27124 (N_27124,N_23569,N_22342);
or U27125 (N_27125,N_22900,N_21305);
or U27126 (N_27126,N_21946,N_21315);
and U27127 (N_27127,N_20843,N_23899);
or U27128 (N_27128,N_24806,N_22228);
or U27129 (N_27129,N_20066,N_23913);
and U27130 (N_27130,N_23852,N_22358);
nand U27131 (N_27131,N_20820,N_22743);
nor U27132 (N_27132,N_21833,N_23844);
nor U27133 (N_27133,N_22133,N_22188);
and U27134 (N_27134,N_22984,N_24573);
or U27135 (N_27135,N_20406,N_21091);
xor U27136 (N_27136,N_23189,N_23228);
nand U27137 (N_27137,N_24230,N_23094);
nor U27138 (N_27138,N_21094,N_24018);
or U27139 (N_27139,N_24523,N_20146);
xor U27140 (N_27140,N_23944,N_24546);
nor U27141 (N_27141,N_21323,N_21537);
xnor U27142 (N_27142,N_24194,N_22856);
nor U27143 (N_27143,N_20027,N_23690);
nand U27144 (N_27144,N_21227,N_24719);
nand U27145 (N_27145,N_23696,N_22894);
or U27146 (N_27146,N_20025,N_21838);
nand U27147 (N_27147,N_23196,N_21770);
and U27148 (N_27148,N_24713,N_23174);
or U27149 (N_27149,N_20068,N_24364);
nand U27150 (N_27150,N_23453,N_23883);
nor U27151 (N_27151,N_21044,N_22470);
nor U27152 (N_27152,N_22994,N_23830);
xor U27153 (N_27153,N_24612,N_22568);
xor U27154 (N_27154,N_24888,N_21933);
nor U27155 (N_27155,N_24650,N_20985);
nand U27156 (N_27156,N_23836,N_22011);
and U27157 (N_27157,N_21889,N_20502);
or U27158 (N_27158,N_23205,N_23167);
and U27159 (N_27159,N_23658,N_22688);
nand U27160 (N_27160,N_20486,N_24530);
nand U27161 (N_27161,N_20462,N_24955);
nor U27162 (N_27162,N_21698,N_23034);
or U27163 (N_27163,N_21263,N_22075);
and U27164 (N_27164,N_22582,N_24001);
nor U27165 (N_27165,N_20051,N_20360);
nor U27166 (N_27166,N_20737,N_24964);
nand U27167 (N_27167,N_21784,N_20171);
and U27168 (N_27168,N_23684,N_24933);
xnor U27169 (N_27169,N_24422,N_20548);
nor U27170 (N_27170,N_24405,N_21013);
xor U27171 (N_27171,N_24372,N_20934);
xor U27172 (N_27172,N_23110,N_23563);
nor U27173 (N_27173,N_21913,N_24394);
xnor U27174 (N_27174,N_23018,N_23439);
or U27175 (N_27175,N_22540,N_20343);
nor U27176 (N_27176,N_20120,N_23041);
nand U27177 (N_27177,N_23799,N_22154);
nor U27178 (N_27178,N_20898,N_22387);
nand U27179 (N_27179,N_24140,N_23531);
xnor U27180 (N_27180,N_23396,N_24584);
or U27181 (N_27181,N_24561,N_20533);
or U27182 (N_27182,N_22781,N_22463);
xnor U27183 (N_27183,N_22935,N_20041);
nand U27184 (N_27184,N_21899,N_24047);
xor U27185 (N_27185,N_23550,N_20252);
or U27186 (N_27186,N_20911,N_20752);
xnor U27187 (N_27187,N_20995,N_21798);
nand U27188 (N_27188,N_20918,N_21153);
and U27189 (N_27189,N_24320,N_20620);
xnor U27190 (N_27190,N_22634,N_21379);
xor U27191 (N_27191,N_20321,N_20804);
nand U27192 (N_27192,N_22428,N_20949);
nor U27193 (N_27193,N_23152,N_22201);
xor U27194 (N_27194,N_20957,N_23421);
or U27195 (N_27195,N_20227,N_22679);
nand U27196 (N_27196,N_22294,N_20530);
xor U27197 (N_27197,N_23943,N_22520);
and U27198 (N_27198,N_20694,N_24240);
nor U27199 (N_27199,N_24808,N_21463);
nand U27200 (N_27200,N_24547,N_20401);
nand U27201 (N_27201,N_22175,N_20471);
or U27202 (N_27202,N_20751,N_22474);
nand U27203 (N_27203,N_22400,N_24800);
nand U27204 (N_27204,N_23240,N_24525);
or U27205 (N_27205,N_24875,N_21982);
nand U27206 (N_27206,N_20110,N_22961);
and U27207 (N_27207,N_24934,N_20012);
xor U27208 (N_27208,N_23382,N_22640);
or U27209 (N_27209,N_23619,N_21539);
xor U27210 (N_27210,N_23362,N_23165);
and U27211 (N_27211,N_21143,N_23694);
xor U27212 (N_27212,N_20514,N_21046);
nor U27213 (N_27213,N_22221,N_21714);
xor U27214 (N_27214,N_24585,N_23086);
and U27215 (N_27215,N_21139,N_24791);
and U27216 (N_27216,N_22882,N_24553);
or U27217 (N_27217,N_24151,N_23851);
and U27218 (N_27218,N_24306,N_20429);
nand U27219 (N_27219,N_22893,N_23646);
xor U27220 (N_27220,N_22922,N_20776);
or U27221 (N_27221,N_24029,N_23276);
xnor U27222 (N_27222,N_21700,N_23330);
xor U27223 (N_27223,N_21075,N_24979);
or U27224 (N_27224,N_21364,N_24580);
nand U27225 (N_27225,N_21021,N_23270);
and U27226 (N_27226,N_21792,N_24383);
xor U27227 (N_27227,N_23948,N_23689);
nor U27228 (N_27228,N_20269,N_22771);
xnor U27229 (N_27229,N_24454,N_21192);
nor U27230 (N_27230,N_22788,N_21562);
xor U27231 (N_27231,N_22707,N_21831);
or U27232 (N_27232,N_21042,N_22317);
or U27233 (N_27233,N_22514,N_20815);
nor U27234 (N_27234,N_22163,N_20861);
and U27235 (N_27235,N_20968,N_20156);
nand U27236 (N_27236,N_24261,N_22753);
or U27237 (N_27237,N_24867,N_23523);
or U27238 (N_27238,N_21179,N_21932);
xor U27239 (N_27239,N_22058,N_22442);
nand U27240 (N_27240,N_20024,N_20290);
nand U27241 (N_27241,N_23301,N_20623);
and U27242 (N_27242,N_22500,N_20203);
nor U27243 (N_27243,N_23888,N_20939);
and U27244 (N_27244,N_23871,N_23533);
xnor U27245 (N_27245,N_20362,N_21453);
nor U27246 (N_27246,N_21582,N_24634);
nor U27247 (N_27247,N_24199,N_23119);
and U27248 (N_27248,N_21286,N_21996);
and U27249 (N_27249,N_24376,N_24253);
and U27250 (N_27250,N_23336,N_21492);
and U27251 (N_27251,N_21053,N_21234);
or U27252 (N_27252,N_21848,N_22047);
and U27253 (N_27253,N_22498,N_20873);
or U27254 (N_27254,N_20338,N_24914);
and U27255 (N_27255,N_20725,N_22999);
xor U27256 (N_27256,N_21775,N_21411);
nand U27257 (N_27257,N_23990,N_20488);
nor U27258 (N_27258,N_24956,N_23021);
nand U27259 (N_27259,N_22877,N_24225);
or U27260 (N_27260,N_21388,N_21436);
and U27261 (N_27261,N_21468,N_21867);
or U27262 (N_27262,N_20940,N_20522);
xor U27263 (N_27263,N_21801,N_23611);
xor U27264 (N_27264,N_23208,N_24060);
xnor U27265 (N_27265,N_22286,N_24168);
or U27266 (N_27266,N_21845,N_23321);
nor U27267 (N_27267,N_24874,N_24399);
or U27268 (N_27268,N_21811,N_24951);
nor U27269 (N_27269,N_21296,N_24750);
nor U27270 (N_27270,N_21915,N_24183);
xnor U27271 (N_27271,N_22140,N_23835);
and U27272 (N_27272,N_22505,N_24049);
nor U27273 (N_27273,N_24495,N_24944);
xor U27274 (N_27274,N_20608,N_22273);
nand U27275 (N_27275,N_20824,N_21742);
or U27276 (N_27276,N_24303,N_21777);
or U27277 (N_27277,N_20055,N_20705);
and U27278 (N_27278,N_24175,N_22004);
or U27279 (N_27279,N_22174,N_22681);
xor U27280 (N_27280,N_22611,N_24752);
xor U27281 (N_27281,N_22413,N_21048);
and U27282 (N_27282,N_24386,N_20004);
nand U27283 (N_27283,N_24317,N_20754);
nand U27284 (N_27284,N_20774,N_21631);
nand U27285 (N_27285,N_22186,N_22507);
nand U27286 (N_27286,N_20622,N_22009);
nand U27287 (N_27287,N_21992,N_24920);
nor U27288 (N_27288,N_20280,N_20902);
nand U27289 (N_27289,N_21580,N_22613);
or U27290 (N_27290,N_20049,N_22369);
or U27291 (N_27291,N_20698,N_22742);
and U27292 (N_27292,N_23595,N_20151);
xnor U27293 (N_27293,N_22331,N_24847);
nor U27294 (N_27294,N_24477,N_24607);
xor U27295 (N_27295,N_23214,N_24156);
xor U27296 (N_27296,N_20567,N_22921);
nand U27297 (N_27297,N_22255,N_22130);
xnor U27298 (N_27298,N_20017,N_20320);
nand U27299 (N_27299,N_23103,N_20191);
nand U27300 (N_27300,N_21567,N_23657);
and U27301 (N_27301,N_20545,N_22682);
nor U27302 (N_27302,N_20980,N_22146);
xor U27303 (N_27303,N_22371,N_24042);
and U27304 (N_27304,N_24397,N_22446);
xnor U27305 (N_27305,N_23997,N_23326);
xnor U27306 (N_27306,N_24267,N_22529);
nor U27307 (N_27307,N_21505,N_21477);
nor U27308 (N_27308,N_20481,N_20673);
nand U27309 (N_27309,N_24421,N_24379);
nand U27310 (N_27310,N_22798,N_20178);
or U27311 (N_27311,N_22160,N_22904);
xor U27312 (N_27312,N_20472,N_21444);
or U27313 (N_27313,N_24630,N_23930);
or U27314 (N_27314,N_24389,N_20539);
and U27315 (N_27315,N_24293,N_20878);
and U27316 (N_27316,N_20028,N_24085);
nand U27317 (N_27317,N_21415,N_21684);
and U27318 (N_27318,N_21968,N_20468);
nor U27319 (N_27319,N_23908,N_24503);
nor U27320 (N_27320,N_23921,N_24418);
xnor U27321 (N_27321,N_23369,N_20849);
xnor U27322 (N_27322,N_23518,N_24841);
and U27323 (N_27323,N_22833,N_23309);
or U27324 (N_27324,N_23780,N_21612);
or U27325 (N_27325,N_23267,N_23570);
nand U27326 (N_27326,N_23314,N_24087);
or U27327 (N_27327,N_23391,N_20180);
nand U27328 (N_27328,N_21761,N_24908);
xnor U27329 (N_27329,N_24427,N_22908);
and U27330 (N_27330,N_23934,N_20590);
and U27331 (N_27331,N_20586,N_24470);
nor U27332 (N_27332,N_20528,N_23340);
nor U27333 (N_27333,N_24660,N_21638);
or U27334 (N_27334,N_24614,N_23185);
xor U27335 (N_27335,N_22423,N_21137);
nor U27336 (N_27336,N_21098,N_24219);
xor U27337 (N_27337,N_21601,N_24011);
nor U27338 (N_27338,N_21686,N_23642);
nand U27339 (N_27339,N_20588,N_21905);
or U27340 (N_27340,N_20205,N_24864);
nand U27341 (N_27341,N_20743,N_21106);
and U27342 (N_27342,N_21469,N_23645);
nand U27343 (N_27343,N_23520,N_21365);
nand U27344 (N_27344,N_23191,N_22997);
xor U27345 (N_27345,N_23195,N_22734);
and U27346 (N_27346,N_22138,N_22094);
or U27347 (N_27347,N_23019,N_20948);
or U27348 (N_27348,N_22366,N_20848);
nor U27349 (N_27349,N_20723,N_23768);
or U27350 (N_27350,N_23742,N_21092);
xor U27351 (N_27351,N_23409,N_21418);
xnor U27352 (N_27352,N_23596,N_20427);
nor U27353 (N_27353,N_23924,N_24929);
xor U27354 (N_27354,N_22127,N_23880);
and U27355 (N_27355,N_23946,N_24091);
and U27356 (N_27356,N_20520,N_20395);
or U27357 (N_27357,N_22566,N_20715);
and U27358 (N_27358,N_21893,N_22791);
and U27359 (N_27359,N_24854,N_24507);
nand U27360 (N_27360,N_20379,N_24365);
xnor U27361 (N_27361,N_23641,N_23760);
xnor U27362 (N_27362,N_21987,N_20285);
nor U27363 (N_27363,N_20477,N_24755);
and U27364 (N_27364,N_22332,N_22496);
or U27365 (N_27365,N_21283,N_20334);
and U27366 (N_27366,N_20632,N_23397);
xor U27367 (N_27367,N_20749,N_22129);
nand U27368 (N_27368,N_20540,N_22037);
xnor U27369 (N_27369,N_21846,N_24886);
xnor U27370 (N_27370,N_20880,N_20993);
or U27371 (N_27371,N_23771,N_22157);
nor U27372 (N_27372,N_22236,N_24749);
xor U27373 (N_27373,N_22481,N_24615);
nor U27374 (N_27374,N_23256,N_22131);
or U27375 (N_27375,N_20314,N_23807);
or U27376 (N_27376,N_22526,N_21421);
or U27377 (N_27377,N_23433,N_20975);
and U27378 (N_27378,N_21461,N_20473);
nand U27379 (N_27379,N_20067,N_20791);
or U27380 (N_27380,N_24264,N_22584);
and U27381 (N_27381,N_20493,N_22756);
and U27382 (N_27382,N_24701,N_24371);
nand U27383 (N_27383,N_23993,N_22324);
nor U27384 (N_27384,N_24772,N_20127);
nor U27385 (N_27385,N_24493,N_20826);
or U27386 (N_27386,N_24335,N_21791);
xor U27387 (N_27387,N_20687,N_21353);
or U27388 (N_27388,N_24144,N_23459);
nor U27389 (N_27389,N_21238,N_21005);
or U27390 (N_27390,N_22879,N_21711);
nand U27391 (N_27391,N_24811,N_20437);
xnor U27392 (N_27392,N_23066,N_23203);
or U27393 (N_27393,N_23649,N_21047);
nor U27394 (N_27394,N_21683,N_22040);
nand U27395 (N_27395,N_23352,N_21971);
nor U27396 (N_27396,N_23800,N_23636);
nor U27397 (N_27397,N_23552,N_22214);
nand U27398 (N_27398,N_20094,N_22467);
and U27399 (N_27399,N_22667,N_21805);
and U27400 (N_27400,N_20390,N_22100);
nor U27401 (N_27401,N_24682,N_23597);
or U27402 (N_27402,N_24131,N_22216);
nand U27403 (N_27403,N_20779,N_22093);
and U27404 (N_27404,N_23192,N_20781);
xnor U27405 (N_27405,N_24685,N_23334);
and U27406 (N_27406,N_23057,N_24769);
and U27407 (N_27407,N_21362,N_21564);
and U27408 (N_27408,N_21817,N_22701);
nor U27409 (N_27409,N_20373,N_21673);
and U27410 (N_27410,N_22647,N_23785);
and U27411 (N_27411,N_24050,N_20270);
and U27412 (N_27412,N_20036,N_24294);
nand U27413 (N_27413,N_21550,N_24252);
nor U27414 (N_27414,N_20117,N_24097);
and U27415 (N_27415,N_22445,N_21824);
xnor U27416 (N_27416,N_22899,N_24926);
nor U27417 (N_27417,N_22940,N_22237);
and U27418 (N_27418,N_21185,N_20206);
nand U27419 (N_27419,N_23224,N_22955);
or U27420 (N_27420,N_24189,N_21847);
nor U27421 (N_27421,N_24544,N_23886);
xnor U27422 (N_27422,N_21105,N_23176);
and U27423 (N_27423,N_21225,N_20572);
xor U27424 (N_27424,N_22089,N_20316);
nand U27425 (N_27425,N_21294,N_22121);
or U27426 (N_27426,N_24715,N_22307);
or U27427 (N_27427,N_20374,N_20556);
and U27428 (N_27428,N_24141,N_20197);
nand U27429 (N_27429,N_20454,N_20054);
or U27430 (N_27430,N_21126,N_20711);
or U27431 (N_27431,N_21524,N_22932);
nand U27432 (N_27432,N_22586,N_23668);
nand U27433 (N_27433,N_23105,N_21924);
xnor U27434 (N_27434,N_22801,N_24648);
xor U27435 (N_27435,N_24327,N_24355);
nand U27436 (N_27436,N_24274,N_24834);
nor U27437 (N_27437,N_23647,N_24135);
xnor U27438 (N_27438,N_22768,N_24471);
nand U27439 (N_27439,N_23539,N_21236);
or U27440 (N_27440,N_22471,N_20154);
nor U27441 (N_27441,N_21903,N_23973);
and U27442 (N_27442,N_22625,N_21599);
and U27443 (N_27443,N_22411,N_24078);
or U27444 (N_27444,N_22896,N_22802);
nand U27445 (N_27445,N_23950,N_23703);
nor U27446 (N_27446,N_20732,N_20999);
xor U27447 (N_27447,N_20507,N_22654);
nor U27448 (N_27448,N_22624,N_24025);
xor U27449 (N_27449,N_24827,N_24412);
xor U27450 (N_27450,N_22952,N_22139);
nor U27451 (N_27451,N_20106,N_23180);
nand U27452 (N_27452,N_20748,N_21556);
xnor U27453 (N_27453,N_23128,N_24814);
nor U27454 (N_27454,N_23686,N_24766);
and U27455 (N_27455,N_20882,N_22543);
nor U27456 (N_27456,N_20719,N_21051);
nand U27457 (N_27457,N_20002,N_23293);
nand U27458 (N_27458,N_21907,N_21330);
or U27459 (N_27459,N_20681,N_21566);
xnor U27460 (N_27460,N_24541,N_22846);
xnor U27461 (N_27461,N_21872,N_20317);
xnor U27462 (N_27462,N_23891,N_24116);
nor U27463 (N_27463,N_20309,N_20750);
or U27464 (N_27464,N_22124,N_24792);
nand U27465 (N_27465,N_21767,N_21532);
nand U27466 (N_27466,N_23121,N_20807);
nand U27467 (N_27467,N_21561,N_24998);
nand U27468 (N_27468,N_21644,N_24702);
and U27469 (N_27469,N_20045,N_20453);
nor U27470 (N_27470,N_23193,N_24453);
and U27471 (N_27471,N_24999,N_24540);
xnor U27472 (N_27472,N_20006,N_23514);
and U27473 (N_27473,N_21998,N_22630);
and U27474 (N_27474,N_23587,N_21839);
xnor U27475 (N_27475,N_20716,N_22085);
xor U27476 (N_27476,N_22062,N_21632);
and U27477 (N_27477,N_20928,N_24494);
nor U27478 (N_27478,N_23230,N_21557);
nor U27479 (N_27479,N_20193,N_21253);
xnor U27480 (N_27480,N_23117,N_22523);
nand U27481 (N_27481,N_21525,N_22866);
and U27482 (N_27482,N_22076,N_23778);
nor U27483 (N_27483,N_24884,N_22404);
nor U27484 (N_27484,N_22469,N_23920);
or U27485 (N_27485,N_23042,N_21101);
and U27486 (N_27486,N_24733,N_24949);
and U27487 (N_27487,N_21301,N_23493);
nor U27488 (N_27488,N_22963,N_23001);
or U27489 (N_27489,N_22079,N_21795);
or U27490 (N_27490,N_24329,N_22794);
and U27491 (N_27491,N_23889,N_21159);
nor U27492 (N_27492,N_21606,N_23236);
and U27493 (N_27493,N_24158,N_23088);
nor U27494 (N_27494,N_24916,N_24737);
or U27495 (N_27495,N_22843,N_22521);
xor U27496 (N_27496,N_21147,N_20922);
xor U27497 (N_27497,N_20676,N_22296);
nand U27498 (N_27498,N_23259,N_23255);
or U27499 (N_27499,N_23123,N_24260);
or U27500 (N_27500,N_21689,N_24166);
xor U27501 (N_27501,N_21382,N_23846);
or U27502 (N_27502,N_21598,N_22141);
nor U27503 (N_27503,N_23272,N_22794);
and U27504 (N_27504,N_23842,N_24198);
xnor U27505 (N_27505,N_23489,N_21812);
and U27506 (N_27506,N_22350,N_24004);
and U27507 (N_27507,N_22308,N_20047);
nand U27508 (N_27508,N_23906,N_23998);
or U27509 (N_27509,N_22153,N_22626);
nand U27510 (N_27510,N_24163,N_22647);
or U27511 (N_27511,N_22398,N_22025);
nand U27512 (N_27512,N_22969,N_22011);
and U27513 (N_27513,N_23828,N_22076);
and U27514 (N_27514,N_21083,N_23296);
nand U27515 (N_27515,N_22045,N_22238);
and U27516 (N_27516,N_21776,N_21720);
nand U27517 (N_27517,N_22544,N_21279);
and U27518 (N_27518,N_23660,N_21556);
or U27519 (N_27519,N_23139,N_22878);
or U27520 (N_27520,N_22416,N_24895);
nand U27521 (N_27521,N_20913,N_20660);
or U27522 (N_27522,N_21644,N_23656);
xor U27523 (N_27523,N_21998,N_22067);
and U27524 (N_27524,N_20853,N_24928);
nor U27525 (N_27525,N_24735,N_24319);
nand U27526 (N_27526,N_21560,N_22809);
or U27527 (N_27527,N_24677,N_21190);
and U27528 (N_27528,N_23657,N_23187);
and U27529 (N_27529,N_21600,N_24003);
xor U27530 (N_27530,N_23761,N_21826);
or U27531 (N_27531,N_22227,N_20500);
and U27532 (N_27532,N_21828,N_21706);
nor U27533 (N_27533,N_21100,N_20493);
xor U27534 (N_27534,N_24847,N_20963);
and U27535 (N_27535,N_24481,N_20129);
nand U27536 (N_27536,N_21916,N_20378);
or U27537 (N_27537,N_21806,N_21952);
or U27538 (N_27538,N_20683,N_21792);
and U27539 (N_27539,N_21243,N_21361);
or U27540 (N_27540,N_20962,N_20818);
xor U27541 (N_27541,N_22720,N_21306);
nor U27542 (N_27542,N_24683,N_23040);
xor U27543 (N_27543,N_22426,N_22261);
and U27544 (N_27544,N_20137,N_21603);
and U27545 (N_27545,N_22786,N_24077);
or U27546 (N_27546,N_23483,N_22054);
nand U27547 (N_27547,N_24157,N_22714);
or U27548 (N_27548,N_21019,N_21052);
nor U27549 (N_27549,N_21875,N_22534);
nand U27550 (N_27550,N_21151,N_22308);
or U27551 (N_27551,N_20448,N_20815);
or U27552 (N_27552,N_20517,N_21584);
or U27553 (N_27553,N_21390,N_20495);
and U27554 (N_27554,N_23952,N_22847);
nor U27555 (N_27555,N_24551,N_23379);
or U27556 (N_27556,N_24928,N_24816);
nor U27557 (N_27557,N_23336,N_21582);
nand U27558 (N_27558,N_24820,N_24116);
and U27559 (N_27559,N_21512,N_23170);
or U27560 (N_27560,N_20018,N_22284);
xor U27561 (N_27561,N_24581,N_22388);
xor U27562 (N_27562,N_24584,N_24938);
and U27563 (N_27563,N_21289,N_22897);
or U27564 (N_27564,N_20095,N_21327);
or U27565 (N_27565,N_20264,N_23555);
or U27566 (N_27566,N_22817,N_24946);
or U27567 (N_27567,N_23983,N_22326);
and U27568 (N_27568,N_21061,N_21728);
nand U27569 (N_27569,N_22927,N_23432);
and U27570 (N_27570,N_20320,N_22237);
or U27571 (N_27571,N_23056,N_23284);
nand U27572 (N_27572,N_21463,N_24986);
or U27573 (N_27573,N_21642,N_22877);
and U27574 (N_27574,N_23111,N_22397);
xnor U27575 (N_27575,N_21330,N_20179);
and U27576 (N_27576,N_23226,N_21066);
nand U27577 (N_27577,N_20006,N_21419);
xnor U27578 (N_27578,N_20725,N_24801);
and U27579 (N_27579,N_24602,N_20005);
and U27580 (N_27580,N_24945,N_20173);
or U27581 (N_27581,N_22504,N_21987);
nor U27582 (N_27582,N_22471,N_21169);
and U27583 (N_27583,N_23367,N_21366);
and U27584 (N_27584,N_20831,N_21014);
xnor U27585 (N_27585,N_20160,N_20135);
and U27586 (N_27586,N_22195,N_22809);
and U27587 (N_27587,N_21197,N_22522);
nor U27588 (N_27588,N_24759,N_21459);
and U27589 (N_27589,N_21284,N_24128);
and U27590 (N_27590,N_24293,N_20813);
nor U27591 (N_27591,N_21264,N_24156);
nand U27592 (N_27592,N_21067,N_22481);
nor U27593 (N_27593,N_23668,N_24418);
or U27594 (N_27594,N_21717,N_24026);
xor U27595 (N_27595,N_24072,N_20661);
and U27596 (N_27596,N_20665,N_23306);
and U27597 (N_27597,N_24708,N_20981);
nand U27598 (N_27598,N_23335,N_21758);
nand U27599 (N_27599,N_24560,N_24095);
nand U27600 (N_27600,N_23524,N_24932);
nand U27601 (N_27601,N_20776,N_20204);
and U27602 (N_27602,N_22356,N_20788);
xnor U27603 (N_27603,N_22817,N_24084);
xnor U27604 (N_27604,N_23042,N_22003);
and U27605 (N_27605,N_23841,N_22737);
xor U27606 (N_27606,N_24706,N_22015);
nor U27607 (N_27607,N_22720,N_20046);
nand U27608 (N_27608,N_24737,N_20616);
xor U27609 (N_27609,N_20136,N_24525);
nand U27610 (N_27610,N_24755,N_23464);
and U27611 (N_27611,N_22674,N_22794);
nand U27612 (N_27612,N_20059,N_24910);
xnor U27613 (N_27613,N_22802,N_20253);
nand U27614 (N_27614,N_22650,N_22547);
nor U27615 (N_27615,N_24057,N_23044);
xor U27616 (N_27616,N_21203,N_24598);
xor U27617 (N_27617,N_20572,N_21345);
nand U27618 (N_27618,N_24554,N_23645);
and U27619 (N_27619,N_21652,N_24083);
nor U27620 (N_27620,N_22479,N_20306);
or U27621 (N_27621,N_22013,N_24027);
xor U27622 (N_27622,N_22566,N_20762);
or U27623 (N_27623,N_21974,N_24507);
nand U27624 (N_27624,N_22112,N_20969);
nor U27625 (N_27625,N_20000,N_22321);
xnor U27626 (N_27626,N_23001,N_23618);
xor U27627 (N_27627,N_21811,N_23725);
nor U27628 (N_27628,N_23128,N_24161);
xnor U27629 (N_27629,N_22278,N_24782);
nor U27630 (N_27630,N_20374,N_24187);
or U27631 (N_27631,N_20499,N_21080);
or U27632 (N_27632,N_20840,N_20884);
and U27633 (N_27633,N_21170,N_20987);
and U27634 (N_27634,N_23295,N_20816);
xor U27635 (N_27635,N_20903,N_23688);
and U27636 (N_27636,N_24423,N_21291);
and U27637 (N_27637,N_24111,N_23276);
nor U27638 (N_27638,N_20215,N_20204);
nor U27639 (N_27639,N_21590,N_23842);
nand U27640 (N_27640,N_23955,N_20136);
nor U27641 (N_27641,N_23423,N_20336);
and U27642 (N_27642,N_20297,N_20430);
xnor U27643 (N_27643,N_20436,N_22685);
and U27644 (N_27644,N_21406,N_21793);
xor U27645 (N_27645,N_21896,N_21878);
xnor U27646 (N_27646,N_21332,N_24909);
and U27647 (N_27647,N_20741,N_23224);
and U27648 (N_27648,N_22636,N_23965);
or U27649 (N_27649,N_24571,N_20480);
and U27650 (N_27650,N_22802,N_21952);
xor U27651 (N_27651,N_22761,N_22377);
or U27652 (N_27652,N_20688,N_21386);
xnor U27653 (N_27653,N_21259,N_21012);
nand U27654 (N_27654,N_20156,N_24915);
and U27655 (N_27655,N_23711,N_21068);
nor U27656 (N_27656,N_20422,N_20180);
nand U27657 (N_27657,N_21475,N_24787);
xnor U27658 (N_27658,N_22921,N_22933);
nand U27659 (N_27659,N_23023,N_24721);
and U27660 (N_27660,N_23856,N_21692);
xnor U27661 (N_27661,N_24314,N_21154);
and U27662 (N_27662,N_23299,N_21183);
xnor U27663 (N_27663,N_20063,N_24524);
or U27664 (N_27664,N_21665,N_22791);
and U27665 (N_27665,N_20288,N_23703);
and U27666 (N_27666,N_20127,N_21418);
nor U27667 (N_27667,N_24584,N_24114);
nand U27668 (N_27668,N_22539,N_23239);
nor U27669 (N_27669,N_22928,N_24610);
or U27670 (N_27670,N_24962,N_24698);
or U27671 (N_27671,N_24688,N_22586);
and U27672 (N_27672,N_23161,N_21649);
xnor U27673 (N_27673,N_24680,N_23222);
xnor U27674 (N_27674,N_22791,N_23614);
nor U27675 (N_27675,N_20613,N_20423);
nor U27676 (N_27676,N_22724,N_20425);
and U27677 (N_27677,N_21333,N_21919);
nand U27678 (N_27678,N_20922,N_23726);
or U27679 (N_27679,N_23981,N_22058);
and U27680 (N_27680,N_20149,N_24272);
nor U27681 (N_27681,N_21136,N_20855);
nor U27682 (N_27682,N_20704,N_23501);
nor U27683 (N_27683,N_24491,N_23878);
xnor U27684 (N_27684,N_24787,N_24136);
and U27685 (N_27685,N_24627,N_22172);
nand U27686 (N_27686,N_21434,N_21998);
nor U27687 (N_27687,N_21370,N_24346);
nor U27688 (N_27688,N_22953,N_21725);
xor U27689 (N_27689,N_22994,N_20842);
or U27690 (N_27690,N_22056,N_20000);
or U27691 (N_27691,N_22337,N_21225);
and U27692 (N_27692,N_20929,N_20369);
nor U27693 (N_27693,N_20706,N_21961);
or U27694 (N_27694,N_22911,N_24618);
xor U27695 (N_27695,N_20151,N_20112);
nand U27696 (N_27696,N_24160,N_21037);
or U27697 (N_27697,N_24961,N_22653);
or U27698 (N_27698,N_23997,N_23858);
nand U27699 (N_27699,N_22501,N_23364);
or U27700 (N_27700,N_21131,N_20818);
nand U27701 (N_27701,N_24162,N_23611);
xor U27702 (N_27702,N_21542,N_23615);
and U27703 (N_27703,N_24290,N_22383);
nor U27704 (N_27704,N_21187,N_20460);
xnor U27705 (N_27705,N_22985,N_24456);
nor U27706 (N_27706,N_21412,N_24451);
xor U27707 (N_27707,N_23355,N_24377);
nand U27708 (N_27708,N_22367,N_20004);
nand U27709 (N_27709,N_22846,N_21622);
nor U27710 (N_27710,N_23634,N_20609);
xor U27711 (N_27711,N_20754,N_24696);
and U27712 (N_27712,N_22053,N_22822);
and U27713 (N_27713,N_24225,N_20904);
nand U27714 (N_27714,N_24842,N_22325);
xnor U27715 (N_27715,N_21291,N_22176);
nand U27716 (N_27716,N_24768,N_20558);
xor U27717 (N_27717,N_24884,N_24370);
and U27718 (N_27718,N_23117,N_20386);
xnor U27719 (N_27719,N_23034,N_21618);
nor U27720 (N_27720,N_20078,N_20733);
or U27721 (N_27721,N_22182,N_21251);
nor U27722 (N_27722,N_21663,N_22872);
nand U27723 (N_27723,N_23413,N_21635);
nor U27724 (N_27724,N_23988,N_24338);
xor U27725 (N_27725,N_22008,N_24902);
or U27726 (N_27726,N_23880,N_23527);
nand U27727 (N_27727,N_23283,N_22176);
and U27728 (N_27728,N_24830,N_23517);
or U27729 (N_27729,N_24298,N_21985);
nand U27730 (N_27730,N_21732,N_22710);
xor U27731 (N_27731,N_21581,N_24202);
xor U27732 (N_27732,N_24668,N_23240);
nor U27733 (N_27733,N_20402,N_23833);
nand U27734 (N_27734,N_23480,N_24431);
nand U27735 (N_27735,N_21043,N_22240);
nor U27736 (N_27736,N_23608,N_22254);
nor U27737 (N_27737,N_20334,N_21717);
or U27738 (N_27738,N_21642,N_20653);
or U27739 (N_27739,N_20745,N_20709);
xor U27740 (N_27740,N_23350,N_20397);
nor U27741 (N_27741,N_24646,N_20890);
and U27742 (N_27742,N_22859,N_20042);
nand U27743 (N_27743,N_22276,N_22361);
or U27744 (N_27744,N_20904,N_20687);
xor U27745 (N_27745,N_20225,N_21166);
xor U27746 (N_27746,N_24158,N_20518);
nor U27747 (N_27747,N_21541,N_24574);
and U27748 (N_27748,N_20980,N_20822);
nand U27749 (N_27749,N_22665,N_22430);
and U27750 (N_27750,N_21121,N_21923);
nand U27751 (N_27751,N_21114,N_22041);
or U27752 (N_27752,N_21694,N_20352);
nand U27753 (N_27753,N_22689,N_22911);
or U27754 (N_27754,N_24233,N_24068);
and U27755 (N_27755,N_22502,N_24952);
xnor U27756 (N_27756,N_22421,N_23117);
or U27757 (N_27757,N_22318,N_20350);
nor U27758 (N_27758,N_22571,N_20663);
xor U27759 (N_27759,N_24198,N_22579);
xnor U27760 (N_27760,N_22181,N_24994);
xnor U27761 (N_27761,N_22141,N_24199);
or U27762 (N_27762,N_20290,N_20152);
and U27763 (N_27763,N_23901,N_21642);
nor U27764 (N_27764,N_22967,N_21993);
and U27765 (N_27765,N_21380,N_21571);
and U27766 (N_27766,N_22832,N_22719);
xnor U27767 (N_27767,N_21485,N_20179);
and U27768 (N_27768,N_22409,N_22039);
and U27769 (N_27769,N_21678,N_23727);
and U27770 (N_27770,N_24404,N_22192);
xnor U27771 (N_27771,N_24863,N_21257);
xnor U27772 (N_27772,N_21752,N_24232);
nand U27773 (N_27773,N_24810,N_23090);
nor U27774 (N_27774,N_21193,N_24658);
and U27775 (N_27775,N_20961,N_20862);
nor U27776 (N_27776,N_22275,N_20880);
nor U27777 (N_27777,N_20478,N_23046);
nand U27778 (N_27778,N_23043,N_20529);
or U27779 (N_27779,N_23742,N_23757);
nand U27780 (N_27780,N_22919,N_23128);
or U27781 (N_27781,N_24547,N_22616);
nand U27782 (N_27782,N_23962,N_20311);
nand U27783 (N_27783,N_22031,N_23337);
nand U27784 (N_27784,N_24409,N_20281);
and U27785 (N_27785,N_23392,N_24874);
nand U27786 (N_27786,N_23110,N_23726);
and U27787 (N_27787,N_23234,N_24157);
and U27788 (N_27788,N_20501,N_23963);
or U27789 (N_27789,N_24209,N_21321);
and U27790 (N_27790,N_24357,N_20089);
xnor U27791 (N_27791,N_20452,N_23336);
xnor U27792 (N_27792,N_24895,N_24827);
and U27793 (N_27793,N_22521,N_24324);
nor U27794 (N_27794,N_21421,N_20588);
xnor U27795 (N_27795,N_20409,N_24036);
xor U27796 (N_27796,N_21996,N_22606);
xnor U27797 (N_27797,N_24474,N_21818);
or U27798 (N_27798,N_20019,N_23361);
nor U27799 (N_27799,N_23490,N_23412);
xor U27800 (N_27800,N_20224,N_21335);
xnor U27801 (N_27801,N_24237,N_24315);
xnor U27802 (N_27802,N_22313,N_22647);
nand U27803 (N_27803,N_20582,N_21236);
nor U27804 (N_27804,N_24936,N_22011);
xor U27805 (N_27805,N_21387,N_23402);
and U27806 (N_27806,N_20636,N_23412);
xnor U27807 (N_27807,N_23455,N_23277);
and U27808 (N_27808,N_24251,N_21979);
and U27809 (N_27809,N_20998,N_23587);
nor U27810 (N_27810,N_22425,N_22160);
or U27811 (N_27811,N_24702,N_21495);
nand U27812 (N_27812,N_24732,N_24245);
nand U27813 (N_27813,N_24139,N_20962);
nand U27814 (N_27814,N_20551,N_22760);
xnor U27815 (N_27815,N_20129,N_21801);
nand U27816 (N_27816,N_24230,N_21498);
nand U27817 (N_27817,N_24844,N_24087);
xnor U27818 (N_27818,N_23232,N_24895);
or U27819 (N_27819,N_20591,N_21186);
xnor U27820 (N_27820,N_20511,N_23068);
or U27821 (N_27821,N_20409,N_20814);
and U27822 (N_27822,N_22543,N_23729);
xnor U27823 (N_27823,N_20722,N_22050);
and U27824 (N_27824,N_22226,N_24727);
xor U27825 (N_27825,N_22204,N_24625);
or U27826 (N_27826,N_23272,N_24590);
nand U27827 (N_27827,N_21759,N_20773);
xnor U27828 (N_27828,N_22536,N_21905);
or U27829 (N_27829,N_24760,N_20843);
nor U27830 (N_27830,N_23649,N_23628);
xnor U27831 (N_27831,N_22314,N_24938);
or U27832 (N_27832,N_21780,N_24639);
and U27833 (N_27833,N_23101,N_23295);
and U27834 (N_27834,N_22764,N_24193);
and U27835 (N_27835,N_22101,N_24651);
xnor U27836 (N_27836,N_24877,N_22325);
nand U27837 (N_27837,N_20118,N_22787);
xor U27838 (N_27838,N_22390,N_20855);
and U27839 (N_27839,N_24286,N_22214);
and U27840 (N_27840,N_24278,N_20352);
nand U27841 (N_27841,N_20120,N_21088);
xor U27842 (N_27842,N_24038,N_24929);
or U27843 (N_27843,N_21744,N_24374);
or U27844 (N_27844,N_21278,N_22847);
nor U27845 (N_27845,N_24134,N_23542);
nor U27846 (N_27846,N_22126,N_22243);
and U27847 (N_27847,N_23887,N_20351);
nor U27848 (N_27848,N_24775,N_22295);
and U27849 (N_27849,N_20327,N_20565);
nor U27850 (N_27850,N_20991,N_23245);
xnor U27851 (N_27851,N_23806,N_23715);
or U27852 (N_27852,N_20413,N_20349);
nor U27853 (N_27853,N_24112,N_20885);
or U27854 (N_27854,N_24113,N_22142);
and U27855 (N_27855,N_24393,N_23322);
and U27856 (N_27856,N_23899,N_22785);
xnor U27857 (N_27857,N_24129,N_21172);
xnor U27858 (N_27858,N_21560,N_24107);
xor U27859 (N_27859,N_24601,N_20402);
nand U27860 (N_27860,N_22271,N_23661);
nor U27861 (N_27861,N_23903,N_21287);
nor U27862 (N_27862,N_20731,N_22396);
and U27863 (N_27863,N_21532,N_22002);
nor U27864 (N_27864,N_22507,N_22317);
and U27865 (N_27865,N_24324,N_21602);
and U27866 (N_27866,N_24969,N_20463);
and U27867 (N_27867,N_23036,N_22177);
or U27868 (N_27868,N_23163,N_23436);
and U27869 (N_27869,N_24191,N_20234);
nor U27870 (N_27870,N_24240,N_24794);
nand U27871 (N_27871,N_24672,N_22353);
or U27872 (N_27872,N_23840,N_22847);
or U27873 (N_27873,N_22492,N_23317);
xnor U27874 (N_27874,N_24523,N_20870);
and U27875 (N_27875,N_21442,N_23469);
nor U27876 (N_27876,N_22465,N_23128);
nand U27877 (N_27877,N_22937,N_20054);
nand U27878 (N_27878,N_20225,N_20939);
xnor U27879 (N_27879,N_22214,N_23704);
and U27880 (N_27880,N_20094,N_23985);
nand U27881 (N_27881,N_23303,N_23014);
or U27882 (N_27882,N_20420,N_24403);
and U27883 (N_27883,N_23708,N_24338);
nor U27884 (N_27884,N_22233,N_23310);
nor U27885 (N_27885,N_21120,N_22155);
xnor U27886 (N_27886,N_24602,N_24929);
or U27887 (N_27887,N_21049,N_20517);
xor U27888 (N_27888,N_23961,N_23299);
xor U27889 (N_27889,N_22968,N_23396);
nor U27890 (N_27890,N_22345,N_20430);
and U27891 (N_27891,N_23966,N_23306);
xor U27892 (N_27892,N_23895,N_22535);
or U27893 (N_27893,N_21694,N_23140);
and U27894 (N_27894,N_23896,N_24728);
xor U27895 (N_27895,N_22735,N_20133);
or U27896 (N_27896,N_23711,N_21593);
and U27897 (N_27897,N_21827,N_20006);
xnor U27898 (N_27898,N_23332,N_20941);
xnor U27899 (N_27899,N_20602,N_24723);
nand U27900 (N_27900,N_23461,N_20028);
nor U27901 (N_27901,N_24633,N_21131);
nor U27902 (N_27902,N_24540,N_24712);
or U27903 (N_27903,N_24421,N_23884);
or U27904 (N_27904,N_21237,N_24006);
or U27905 (N_27905,N_21729,N_22520);
nand U27906 (N_27906,N_23431,N_23867);
nand U27907 (N_27907,N_23758,N_24674);
nand U27908 (N_27908,N_23641,N_21879);
or U27909 (N_27909,N_21757,N_23834);
and U27910 (N_27910,N_21063,N_20553);
or U27911 (N_27911,N_23473,N_22030);
nor U27912 (N_27912,N_23537,N_22024);
nor U27913 (N_27913,N_23264,N_23160);
nand U27914 (N_27914,N_22036,N_24503);
and U27915 (N_27915,N_22481,N_22643);
nand U27916 (N_27916,N_21823,N_24115);
nand U27917 (N_27917,N_21472,N_24749);
nand U27918 (N_27918,N_22095,N_22691);
or U27919 (N_27919,N_24782,N_22559);
nand U27920 (N_27920,N_20277,N_23513);
or U27921 (N_27921,N_20253,N_22303);
and U27922 (N_27922,N_22551,N_23802);
or U27923 (N_27923,N_23959,N_21421);
xor U27924 (N_27924,N_24021,N_24416);
or U27925 (N_27925,N_21772,N_23306);
and U27926 (N_27926,N_21981,N_20245);
nor U27927 (N_27927,N_22339,N_21615);
xnor U27928 (N_27928,N_24221,N_21191);
nand U27929 (N_27929,N_23237,N_20782);
xor U27930 (N_27930,N_22599,N_21560);
nand U27931 (N_27931,N_21592,N_20927);
or U27932 (N_27932,N_21860,N_20369);
and U27933 (N_27933,N_23656,N_23356);
and U27934 (N_27934,N_23701,N_21847);
xor U27935 (N_27935,N_23082,N_24257);
nor U27936 (N_27936,N_24235,N_21247);
and U27937 (N_27937,N_24521,N_21681);
nor U27938 (N_27938,N_24099,N_23072);
nand U27939 (N_27939,N_24208,N_20928);
nand U27940 (N_27940,N_22269,N_21727);
nand U27941 (N_27941,N_20691,N_22883);
and U27942 (N_27942,N_22257,N_21662);
nand U27943 (N_27943,N_22322,N_21977);
nand U27944 (N_27944,N_20943,N_23262);
or U27945 (N_27945,N_24865,N_24126);
xnor U27946 (N_27946,N_24749,N_22990);
or U27947 (N_27947,N_22228,N_23279);
nor U27948 (N_27948,N_24627,N_23836);
xor U27949 (N_27949,N_21079,N_24283);
and U27950 (N_27950,N_23605,N_23309);
and U27951 (N_27951,N_22977,N_22303);
nor U27952 (N_27952,N_20757,N_20990);
nor U27953 (N_27953,N_24178,N_22956);
nor U27954 (N_27954,N_23547,N_24310);
nand U27955 (N_27955,N_22380,N_24853);
xnor U27956 (N_27956,N_20404,N_20739);
nand U27957 (N_27957,N_21473,N_24145);
nor U27958 (N_27958,N_21093,N_22370);
nor U27959 (N_27959,N_22783,N_21438);
xor U27960 (N_27960,N_24991,N_24548);
nand U27961 (N_27961,N_21207,N_23277);
nand U27962 (N_27962,N_24693,N_23221);
or U27963 (N_27963,N_23207,N_20784);
nand U27964 (N_27964,N_22529,N_20659);
nand U27965 (N_27965,N_22225,N_22435);
and U27966 (N_27966,N_24171,N_23387);
nor U27967 (N_27967,N_21846,N_22659);
or U27968 (N_27968,N_20929,N_22263);
xnor U27969 (N_27969,N_22388,N_20718);
nor U27970 (N_27970,N_21141,N_24530);
xnor U27971 (N_27971,N_23683,N_22781);
nor U27972 (N_27972,N_22135,N_23696);
or U27973 (N_27973,N_21527,N_21329);
or U27974 (N_27974,N_24368,N_24609);
xor U27975 (N_27975,N_23008,N_20434);
or U27976 (N_27976,N_23985,N_24581);
and U27977 (N_27977,N_21288,N_23381);
and U27978 (N_27978,N_20136,N_21181);
xnor U27979 (N_27979,N_20396,N_23775);
nor U27980 (N_27980,N_23075,N_24480);
and U27981 (N_27981,N_20808,N_21532);
nor U27982 (N_27982,N_23354,N_23467);
nand U27983 (N_27983,N_21238,N_24763);
or U27984 (N_27984,N_22485,N_20665);
nand U27985 (N_27985,N_20262,N_20459);
nor U27986 (N_27986,N_21693,N_24022);
or U27987 (N_27987,N_24230,N_23921);
or U27988 (N_27988,N_21328,N_24019);
xnor U27989 (N_27989,N_20135,N_21171);
nor U27990 (N_27990,N_23822,N_20720);
nand U27991 (N_27991,N_21413,N_24585);
or U27992 (N_27992,N_20567,N_23271);
xnor U27993 (N_27993,N_22314,N_23956);
nand U27994 (N_27994,N_24601,N_24887);
nor U27995 (N_27995,N_20772,N_23827);
nand U27996 (N_27996,N_21419,N_22147);
xor U27997 (N_27997,N_23228,N_22848);
nand U27998 (N_27998,N_23377,N_21554);
nor U27999 (N_27999,N_23700,N_22773);
nand U28000 (N_28000,N_22374,N_23243);
nand U28001 (N_28001,N_21677,N_20422);
nand U28002 (N_28002,N_24183,N_23034);
and U28003 (N_28003,N_21966,N_21708);
xor U28004 (N_28004,N_22447,N_24263);
nor U28005 (N_28005,N_22450,N_22546);
and U28006 (N_28006,N_22276,N_22681);
or U28007 (N_28007,N_20817,N_20318);
nor U28008 (N_28008,N_21871,N_22903);
and U28009 (N_28009,N_24683,N_20578);
nor U28010 (N_28010,N_23946,N_21878);
and U28011 (N_28011,N_23041,N_22769);
nor U28012 (N_28012,N_22108,N_20837);
and U28013 (N_28013,N_24352,N_24693);
nand U28014 (N_28014,N_20602,N_21710);
or U28015 (N_28015,N_23520,N_24693);
or U28016 (N_28016,N_22436,N_24499);
nand U28017 (N_28017,N_20677,N_20979);
nor U28018 (N_28018,N_20985,N_21003);
or U28019 (N_28019,N_21417,N_24608);
and U28020 (N_28020,N_21303,N_23767);
nor U28021 (N_28021,N_23663,N_23956);
and U28022 (N_28022,N_23644,N_20196);
nor U28023 (N_28023,N_22056,N_21193);
xor U28024 (N_28024,N_24755,N_22710);
and U28025 (N_28025,N_23641,N_22109);
xor U28026 (N_28026,N_22562,N_24780);
nand U28027 (N_28027,N_20428,N_24406);
nor U28028 (N_28028,N_24291,N_21488);
nand U28029 (N_28029,N_20271,N_20508);
or U28030 (N_28030,N_21832,N_24821);
or U28031 (N_28031,N_20409,N_21696);
nand U28032 (N_28032,N_23866,N_23578);
nor U28033 (N_28033,N_24306,N_24010);
and U28034 (N_28034,N_22950,N_24433);
and U28035 (N_28035,N_23666,N_21392);
nor U28036 (N_28036,N_21142,N_21674);
nand U28037 (N_28037,N_22568,N_21858);
nand U28038 (N_28038,N_24285,N_20280);
nor U28039 (N_28039,N_24631,N_24890);
or U28040 (N_28040,N_21595,N_24042);
or U28041 (N_28041,N_20844,N_24166);
nor U28042 (N_28042,N_23675,N_23843);
nor U28043 (N_28043,N_24838,N_21425);
nor U28044 (N_28044,N_24133,N_20747);
nor U28045 (N_28045,N_20998,N_23684);
nor U28046 (N_28046,N_23756,N_21746);
or U28047 (N_28047,N_20004,N_21965);
and U28048 (N_28048,N_20508,N_24952);
xnor U28049 (N_28049,N_23066,N_23111);
or U28050 (N_28050,N_24015,N_21124);
xor U28051 (N_28051,N_24773,N_22460);
or U28052 (N_28052,N_23877,N_20782);
and U28053 (N_28053,N_20752,N_23669);
and U28054 (N_28054,N_23671,N_20198);
xor U28055 (N_28055,N_24059,N_21882);
and U28056 (N_28056,N_24865,N_22635);
and U28057 (N_28057,N_20679,N_24572);
or U28058 (N_28058,N_20725,N_23705);
xnor U28059 (N_28059,N_24171,N_23072);
xor U28060 (N_28060,N_23347,N_22102);
and U28061 (N_28061,N_20353,N_23237);
nand U28062 (N_28062,N_24735,N_22668);
xor U28063 (N_28063,N_20438,N_21112);
xnor U28064 (N_28064,N_23814,N_20723);
nand U28065 (N_28065,N_23498,N_24557);
xnor U28066 (N_28066,N_20813,N_21235);
nor U28067 (N_28067,N_22061,N_24226);
nor U28068 (N_28068,N_21849,N_22254);
and U28069 (N_28069,N_24929,N_24142);
or U28070 (N_28070,N_22132,N_20726);
and U28071 (N_28071,N_23593,N_24712);
nor U28072 (N_28072,N_23181,N_23245);
nor U28073 (N_28073,N_24060,N_20482);
and U28074 (N_28074,N_20301,N_20299);
nor U28075 (N_28075,N_21522,N_22076);
or U28076 (N_28076,N_20808,N_21114);
xor U28077 (N_28077,N_22844,N_23353);
nand U28078 (N_28078,N_24266,N_20050);
or U28079 (N_28079,N_20812,N_23831);
xor U28080 (N_28080,N_22878,N_21318);
xor U28081 (N_28081,N_23217,N_22885);
nand U28082 (N_28082,N_23531,N_21854);
xor U28083 (N_28083,N_23240,N_22896);
or U28084 (N_28084,N_22981,N_23780);
or U28085 (N_28085,N_23781,N_22314);
or U28086 (N_28086,N_24967,N_23834);
or U28087 (N_28087,N_20558,N_21222);
xor U28088 (N_28088,N_20712,N_20477);
xor U28089 (N_28089,N_21453,N_22822);
or U28090 (N_28090,N_21786,N_22910);
xor U28091 (N_28091,N_21453,N_22639);
or U28092 (N_28092,N_22550,N_22598);
xor U28093 (N_28093,N_24335,N_22000);
nand U28094 (N_28094,N_22570,N_22126);
or U28095 (N_28095,N_20670,N_24653);
nor U28096 (N_28096,N_24841,N_21624);
or U28097 (N_28097,N_20036,N_22081);
or U28098 (N_28098,N_24707,N_21045);
and U28099 (N_28099,N_22443,N_24833);
nor U28100 (N_28100,N_20722,N_21666);
nand U28101 (N_28101,N_22918,N_20267);
xor U28102 (N_28102,N_20625,N_20631);
xor U28103 (N_28103,N_24834,N_23575);
xor U28104 (N_28104,N_21903,N_23170);
xor U28105 (N_28105,N_23738,N_23667);
nor U28106 (N_28106,N_20486,N_21229);
xnor U28107 (N_28107,N_22878,N_21405);
xor U28108 (N_28108,N_21257,N_23648);
xor U28109 (N_28109,N_21162,N_23716);
nor U28110 (N_28110,N_22311,N_22992);
nand U28111 (N_28111,N_23329,N_21676);
or U28112 (N_28112,N_20125,N_21565);
xnor U28113 (N_28113,N_21344,N_21273);
and U28114 (N_28114,N_24972,N_24655);
and U28115 (N_28115,N_21157,N_22880);
and U28116 (N_28116,N_24706,N_24664);
xor U28117 (N_28117,N_22243,N_22805);
nand U28118 (N_28118,N_21559,N_23088);
nand U28119 (N_28119,N_20708,N_20020);
nand U28120 (N_28120,N_22384,N_24051);
and U28121 (N_28121,N_24918,N_23748);
or U28122 (N_28122,N_24323,N_20423);
nor U28123 (N_28123,N_22060,N_21213);
xnor U28124 (N_28124,N_23072,N_21214);
and U28125 (N_28125,N_24676,N_24662);
xnor U28126 (N_28126,N_22647,N_24690);
xnor U28127 (N_28127,N_23284,N_21700);
nand U28128 (N_28128,N_24075,N_21957);
nand U28129 (N_28129,N_23858,N_20205);
and U28130 (N_28130,N_20486,N_21244);
or U28131 (N_28131,N_21870,N_20405);
nand U28132 (N_28132,N_21592,N_21741);
nand U28133 (N_28133,N_20244,N_22264);
or U28134 (N_28134,N_20302,N_20673);
nor U28135 (N_28135,N_22253,N_22004);
and U28136 (N_28136,N_21151,N_24940);
or U28137 (N_28137,N_22241,N_21479);
nand U28138 (N_28138,N_22198,N_22243);
or U28139 (N_28139,N_20123,N_21211);
or U28140 (N_28140,N_20899,N_20378);
nand U28141 (N_28141,N_21671,N_20481);
or U28142 (N_28142,N_21548,N_21275);
nand U28143 (N_28143,N_22227,N_23681);
or U28144 (N_28144,N_21701,N_24599);
xnor U28145 (N_28145,N_22731,N_24998);
or U28146 (N_28146,N_23672,N_20666);
nand U28147 (N_28147,N_22791,N_22495);
nor U28148 (N_28148,N_20919,N_20762);
or U28149 (N_28149,N_21614,N_22097);
nand U28150 (N_28150,N_20282,N_20351);
nand U28151 (N_28151,N_23458,N_22921);
and U28152 (N_28152,N_20891,N_24702);
nor U28153 (N_28153,N_24966,N_23901);
nand U28154 (N_28154,N_24423,N_21811);
nor U28155 (N_28155,N_21935,N_24477);
nand U28156 (N_28156,N_24810,N_23878);
nor U28157 (N_28157,N_22814,N_24127);
and U28158 (N_28158,N_24018,N_22192);
and U28159 (N_28159,N_22044,N_20226);
nor U28160 (N_28160,N_20988,N_22419);
nand U28161 (N_28161,N_24849,N_21822);
nand U28162 (N_28162,N_20349,N_24369);
nor U28163 (N_28163,N_21544,N_21296);
or U28164 (N_28164,N_21888,N_24409);
and U28165 (N_28165,N_21494,N_20262);
nor U28166 (N_28166,N_20506,N_24597);
xnor U28167 (N_28167,N_24721,N_22984);
nor U28168 (N_28168,N_20608,N_20430);
xnor U28169 (N_28169,N_22000,N_22076);
or U28170 (N_28170,N_24887,N_21840);
or U28171 (N_28171,N_24145,N_23432);
xor U28172 (N_28172,N_23551,N_21558);
nand U28173 (N_28173,N_23409,N_23312);
or U28174 (N_28174,N_21407,N_22136);
and U28175 (N_28175,N_22264,N_23832);
nand U28176 (N_28176,N_21131,N_21213);
nand U28177 (N_28177,N_24349,N_21228);
or U28178 (N_28178,N_23434,N_20599);
xnor U28179 (N_28179,N_24854,N_21811);
or U28180 (N_28180,N_24467,N_23156);
and U28181 (N_28181,N_20900,N_22556);
or U28182 (N_28182,N_23372,N_24291);
and U28183 (N_28183,N_23639,N_22976);
nand U28184 (N_28184,N_23357,N_24008);
or U28185 (N_28185,N_22818,N_21167);
xor U28186 (N_28186,N_21957,N_23091);
or U28187 (N_28187,N_22182,N_21771);
nand U28188 (N_28188,N_24981,N_22442);
or U28189 (N_28189,N_21397,N_22625);
nor U28190 (N_28190,N_21398,N_20465);
nand U28191 (N_28191,N_22728,N_21420);
and U28192 (N_28192,N_22734,N_24314);
nand U28193 (N_28193,N_22779,N_22927);
or U28194 (N_28194,N_21961,N_24709);
or U28195 (N_28195,N_24946,N_24213);
nand U28196 (N_28196,N_24299,N_24164);
nor U28197 (N_28197,N_21634,N_22099);
nor U28198 (N_28198,N_23434,N_20572);
nand U28199 (N_28199,N_24050,N_21235);
xnor U28200 (N_28200,N_22795,N_24504);
nor U28201 (N_28201,N_23916,N_24483);
and U28202 (N_28202,N_20436,N_20471);
nand U28203 (N_28203,N_22790,N_23678);
nor U28204 (N_28204,N_22636,N_21625);
xor U28205 (N_28205,N_20188,N_21779);
nor U28206 (N_28206,N_21442,N_21203);
xnor U28207 (N_28207,N_21187,N_20646);
and U28208 (N_28208,N_21555,N_21347);
and U28209 (N_28209,N_22259,N_21550);
xnor U28210 (N_28210,N_21024,N_20333);
xor U28211 (N_28211,N_24737,N_23834);
or U28212 (N_28212,N_22881,N_20532);
nor U28213 (N_28213,N_23637,N_20433);
or U28214 (N_28214,N_22710,N_20765);
nor U28215 (N_28215,N_24160,N_21177);
xor U28216 (N_28216,N_21710,N_24596);
and U28217 (N_28217,N_20880,N_22360);
nand U28218 (N_28218,N_23736,N_21620);
nor U28219 (N_28219,N_22150,N_23366);
or U28220 (N_28220,N_21051,N_22143);
nor U28221 (N_28221,N_22363,N_22938);
nand U28222 (N_28222,N_22636,N_21565);
and U28223 (N_28223,N_23984,N_22184);
xor U28224 (N_28224,N_23121,N_20448);
or U28225 (N_28225,N_22954,N_22993);
and U28226 (N_28226,N_22110,N_23576);
and U28227 (N_28227,N_24603,N_22755);
nand U28228 (N_28228,N_23509,N_20071);
nor U28229 (N_28229,N_24851,N_22694);
and U28230 (N_28230,N_24754,N_22308);
nor U28231 (N_28231,N_23401,N_20912);
nand U28232 (N_28232,N_21871,N_24669);
or U28233 (N_28233,N_22109,N_24320);
and U28234 (N_28234,N_22461,N_22801);
xnor U28235 (N_28235,N_22361,N_21243);
nand U28236 (N_28236,N_23790,N_22541);
or U28237 (N_28237,N_20498,N_22672);
xor U28238 (N_28238,N_20701,N_21535);
and U28239 (N_28239,N_22143,N_24095);
nand U28240 (N_28240,N_23802,N_20062);
or U28241 (N_28241,N_22564,N_21778);
xor U28242 (N_28242,N_21898,N_24152);
nand U28243 (N_28243,N_23969,N_20761);
and U28244 (N_28244,N_22300,N_22607);
and U28245 (N_28245,N_21619,N_22041);
and U28246 (N_28246,N_24247,N_21896);
nor U28247 (N_28247,N_22902,N_22877);
and U28248 (N_28248,N_24933,N_24134);
and U28249 (N_28249,N_20033,N_22837);
or U28250 (N_28250,N_23870,N_20776);
or U28251 (N_28251,N_24340,N_22116);
nor U28252 (N_28252,N_22770,N_20478);
nand U28253 (N_28253,N_24191,N_24741);
nor U28254 (N_28254,N_24418,N_21525);
or U28255 (N_28255,N_22460,N_21420);
nand U28256 (N_28256,N_23731,N_21770);
nor U28257 (N_28257,N_20466,N_21599);
or U28258 (N_28258,N_24307,N_24762);
xnor U28259 (N_28259,N_21253,N_22634);
xnor U28260 (N_28260,N_22441,N_21847);
and U28261 (N_28261,N_23139,N_23123);
nand U28262 (N_28262,N_20739,N_22738);
nand U28263 (N_28263,N_22975,N_22616);
and U28264 (N_28264,N_21950,N_23358);
xor U28265 (N_28265,N_20648,N_20736);
nand U28266 (N_28266,N_20124,N_21614);
or U28267 (N_28267,N_24873,N_20453);
and U28268 (N_28268,N_24992,N_23503);
and U28269 (N_28269,N_22688,N_21104);
and U28270 (N_28270,N_20340,N_20208);
or U28271 (N_28271,N_22509,N_22125);
xor U28272 (N_28272,N_24942,N_22013);
and U28273 (N_28273,N_23658,N_20998);
xor U28274 (N_28274,N_20005,N_22193);
nor U28275 (N_28275,N_21381,N_24517);
xor U28276 (N_28276,N_21566,N_22223);
or U28277 (N_28277,N_22826,N_21230);
nand U28278 (N_28278,N_23967,N_20336);
xor U28279 (N_28279,N_22294,N_23009);
nand U28280 (N_28280,N_20044,N_22304);
nand U28281 (N_28281,N_24489,N_21621);
xnor U28282 (N_28282,N_22243,N_21008);
nor U28283 (N_28283,N_21143,N_20714);
or U28284 (N_28284,N_22283,N_24588);
and U28285 (N_28285,N_21945,N_21120);
and U28286 (N_28286,N_24107,N_24893);
xor U28287 (N_28287,N_23836,N_20376);
nor U28288 (N_28288,N_23914,N_24314);
and U28289 (N_28289,N_22849,N_22342);
nand U28290 (N_28290,N_23683,N_20032);
and U28291 (N_28291,N_22013,N_22021);
xnor U28292 (N_28292,N_24487,N_20236);
xor U28293 (N_28293,N_22239,N_23980);
xor U28294 (N_28294,N_24414,N_24148);
or U28295 (N_28295,N_24318,N_20950);
and U28296 (N_28296,N_21273,N_23031);
and U28297 (N_28297,N_23744,N_22870);
nor U28298 (N_28298,N_23558,N_22020);
xnor U28299 (N_28299,N_20849,N_24329);
and U28300 (N_28300,N_22316,N_21507);
nand U28301 (N_28301,N_23416,N_23878);
nand U28302 (N_28302,N_21477,N_23854);
nor U28303 (N_28303,N_21854,N_22355);
and U28304 (N_28304,N_22444,N_20376);
xor U28305 (N_28305,N_24562,N_24254);
and U28306 (N_28306,N_24035,N_23562);
nand U28307 (N_28307,N_22298,N_20024);
nand U28308 (N_28308,N_24264,N_24790);
or U28309 (N_28309,N_23231,N_23462);
nor U28310 (N_28310,N_24537,N_24199);
or U28311 (N_28311,N_23823,N_23936);
and U28312 (N_28312,N_24809,N_21123);
or U28313 (N_28313,N_23745,N_22700);
and U28314 (N_28314,N_21591,N_24197);
and U28315 (N_28315,N_21447,N_22672);
and U28316 (N_28316,N_22274,N_22902);
and U28317 (N_28317,N_23744,N_21068);
or U28318 (N_28318,N_20183,N_24589);
nand U28319 (N_28319,N_22717,N_21326);
nand U28320 (N_28320,N_20046,N_21426);
and U28321 (N_28321,N_20788,N_21730);
nor U28322 (N_28322,N_22413,N_20847);
xor U28323 (N_28323,N_21672,N_23055);
and U28324 (N_28324,N_23675,N_22642);
nand U28325 (N_28325,N_23772,N_21427);
nand U28326 (N_28326,N_21010,N_22344);
nor U28327 (N_28327,N_23174,N_20455);
nor U28328 (N_28328,N_20466,N_21833);
nor U28329 (N_28329,N_20667,N_22252);
nand U28330 (N_28330,N_21681,N_21723);
nand U28331 (N_28331,N_24900,N_24006);
xor U28332 (N_28332,N_20796,N_23738);
nand U28333 (N_28333,N_24897,N_22457);
or U28334 (N_28334,N_20945,N_21881);
nand U28335 (N_28335,N_21415,N_22414);
nor U28336 (N_28336,N_21575,N_23282);
xor U28337 (N_28337,N_21342,N_22282);
nor U28338 (N_28338,N_20457,N_20393);
or U28339 (N_28339,N_23697,N_22756);
and U28340 (N_28340,N_21828,N_21205);
xnor U28341 (N_28341,N_22927,N_22055);
and U28342 (N_28342,N_24680,N_22563);
and U28343 (N_28343,N_22537,N_23865);
or U28344 (N_28344,N_20272,N_23898);
xnor U28345 (N_28345,N_21740,N_20516);
xnor U28346 (N_28346,N_22259,N_23974);
nor U28347 (N_28347,N_22212,N_20607);
or U28348 (N_28348,N_20302,N_22909);
nor U28349 (N_28349,N_21710,N_20249);
or U28350 (N_28350,N_21322,N_23053);
and U28351 (N_28351,N_21069,N_20619);
and U28352 (N_28352,N_21486,N_24155);
nor U28353 (N_28353,N_22004,N_20354);
or U28354 (N_28354,N_23041,N_24493);
xnor U28355 (N_28355,N_20268,N_21540);
nand U28356 (N_28356,N_20755,N_24577);
and U28357 (N_28357,N_24897,N_20526);
or U28358 (N_28358,N_24601,N_22089);
or U28359 (N_28359,N_20462,N_22811);
and U28360 (N_28360,N_23041,N_20215);
nor U28361 (N_28361,N_20820,N_24948);
xor U28362 (N_28362,N_23243,N_22670);
xnor U28363 (N_28363,N_20296,N_20074);
nand U28364 (N_28364,N_21410,N_21459);
xor U28365 (N_28365,N_23297,N_20191);
or U28366 (N_28366,N_24330,N_24253);
nor U28367 (N_28367,N_20955,N_23304);
nor U28368 (N_28368,N_20822,N_23032);
or U28369 (N_28369,N_23328,N_24197);
and U28370 (N_28370,N_21876,N_24184);
xnor U28371 (N_28371,N_23506,N_23992);
nand U28372 (N_28372,N_22694,N_23498);
xor U28373 (N_28373,N_20203,N_21921);
or U28374 (N_28374,N_23392,N_23994);
or U28375 (N_28375,N_22925,N_23326);
xor U28376 (N_28376,N_24416,N_20911);
xnor U28377 (N_28377,N_22940,N_21098);
xor U28378 (N_28378,N_24910,N_20125);
nand U28379 (N_28379,N_22319,N_23875);
or U28380 (N_28380,N_24311,N_24739);
nand U28381 (N_28381,N_20629,N_22745);
nand U28382 (N_28382,N_23518,N_23244);
or U28383 (N_28383,N_23429,N_22326);
or U28384 (N_28384,N_23350,N_22989);
nor U28385 (N_28385,N_23555,N_22976);
nand U28386 (N_28386,N_24508,N_23338);
nor U28387 (N_28387,N_23116,N_24101);
nor U28388 (N_28388,N_21525,N_22493);
xnor U28389 (N_28389,N_24952,N_21908);
and U28390 (N_28390,N_21261,N_23828);
nand U28391 (N_28391,N_22478,N_24677);
and U28392 (N_28392,N_23340,N_24549);
xnor U28393 (N_28393,N_23966,N_20062);
nor U28394 (N_28394,N_20626,N_24350);
nor U28395 (N_28395,N_20960,N_21853);
nor U28396 (N_28396,N_22911,N_23448);
nor U28397 (N_28397,N_24187,N_22293);
xor U28398 (N_28398,N_21599,N_20025);
or U28399 (N_28399,N_21666,N_24348);
nor U28400 (N_28400,N_21391,N_22787);
nand U28401 (N_28401,N_22774,N_20776);
nor U28402 (N_28402,N_22258,N_20439);
nand U28403 (N_28403,N_23940,N_24194);
nand U28404 (N_28404,N_21205,N_22713);
and U28405 (N_28405,N_22939,N_22663);
nand U28406 (N_28406,N_23696,N_20806);
xnor U28407 (N_28407,N_21830,N_22112);
nand U28408 (N_28408,N_21902,N_24050);
nand U28409 (N_28409,N_20763,N_20711);
nor U28410 (N_28410,N_24607,N_24791);
and U28411 (N_28411,N_21813,N_21676);
nor U28412 (N_28412,N_22722,N_21783);
or U28413 (N_28413,N_20256,N_24424);
xnor U28414 (N_28414,N_21048,N_24665);
or U28415 (N_28415,N_22186,N_23567);
and U28416 (N_28416,N_20423,N_23281);
nor U28417 (N_28417,N_24196,N_21243);
xnor U28418 (N_28418,N_22924,N_21175);
nor U28419 (N_28419,N_22834,N_21476);
xor U28420 (N_28420,N_24411,N_22501);
and U28421 (N_28421,N_23884,N_23841);
or U28422 (N_28422,N_21527,N_23167);
nand U28423 (N_28423,N_20543,N_24917);
nand U28424 (N_28424,N_22482,N_22288);
xnor U28425 (N_28425,N_24653,N_24717);
nand U28426 (N_28426,N_24862,N_20890);
xor U28427 (N_28427,N_22579,N_23901);
or U28428 (N_28428,N_24437,N_23862);
and U28429 (N_28429,N_24466,N_21721);
nand U28430 (N_28430,N_24836,N_24167);
and U28431 (N_28431,N_24314,N_20145);
and U28432 (N_28432,N_22197,N_22559);
or U28433 (N_28433,N_20893,N_24357);
nand U28434 (N_28434,N_22451,N_22503);
and U28435 (N_28435,N_21046,N_23019);
or U28436 (N_28436,N_24298,N_23087);
or U28437 (N_28437,N_23028,N_20225);
xnor U28438 (N_28438,N_21763,N_24981);
nand U28439 (N_28439,N_22169,N_24835);
nand U28440 (N_28440,N_23250,N_20107);
or U28441 (N_28441,N_21239,N_22023);
nand U28442 (N_28442,N_20412,N_22832);
xor U28443 (N_28443,N_23137,N_22067);
and U28444 (N_28444,N_22484,N_20668);
xnor U28445 (N_28445,N_23194,N_24824);
xnor U28446 (N_28446,N_24702,N_23115);
nor U28447 (N_28447,N_23413,N_20644);
and U28448 (N_28448,N_21889,N_23733);
and U28449 (N_28449,N_22827,N_23284);
nand U28450 (N_28450,N_20681,N_23861);
nand U28451 (N_28451,N_21791,N_20869);
nand U28452 (N_28452,N_21695,N_20095);
or U28453 (N_28453,N_21351,N_22930);
xnor U28454 (N_28454,N_24099,N_23483);
nor U28455 (N_28455,N_22245,N_24706);
or U28456 (N_28456,N_22256,N_22842);
xnor U28457 (N_28457,N_22420,N_22328);
nor U28458 (N_28458,N_21803,N_24593);
or U28459 (N_28459,N_20004,N_20454);
nand U28460 (N_28460,N_23116,N_23610);
xor U28461 (N_28461,N_21679,N_24889);
and U28462 (N_28462,N_21090,N_22435);
or U28463 (N_28463,N_24040,N_23976);
nand U28464 (N_28464,N_20084,N_20857);
nor U28465 (N_28465,N_21738,N_23091);
and U28466 (N_28466,N_20886,N_24961);
or U28467 (N_28467,N_23461,N_22308);
nor U28468 (N_28468,N_22607,N_22932);
nor U28469 (N_28469,N_23486,N_22529);
and U28470 (N_28470,N_20386,N_21649);
xor U28471 (N_28471,N_24330,N_24168);
nand U28472 (N_28472,N_23487,N_22944);
nand U28473 (N_28473,N_24891,N_20245);
nand U28474 (N_28474,N_24241,N_24036);
and U28475 (N_28475,N_22280,N_23411);
nor U28476 (N_28476,N_20636,N_23780);
or U28477 (N_28477,N_23361,N_20095);
and U28478 (N_28478,N_20197,N_24796);
or U28479 (N_28479,N_24677,N_21919);
nand U28480 (N_28480,N_20082,N_22675);
or U28481 (N_28481,N_20198,N_21839);
xnor U28482 (N_28482,N_22761,N_21182);
nand U28483 (N_28483,N_20173,N_24530);
or U28484 (N_28484,N_22969,N_20865);
or U28485 (N_28485,N_21718,N_21628);
nor U28486 (N_28486,N_24866,N_22876);
or U28487 (N_28487,N_24279,N_24789);
nor U28488 (N_28488,N_20628,N_21247);
xnor U28489 (N_28489,N_20635,N_21229);
or U28490 (N_28490,N_22073,N_20140);
or U28491 (N_28491,N_23015,N_21144);
xor U28492 (N_28492,N_21793,N_20750);
xnor U28493 (N_28493,N_24104,N_22184);
nand U28494 (N_28494,N_20637,N_21740);
nand U28495 (N_28495,N_22868,N_21868);
and U28496 (N_28496,N_24306,N_20098);
nor U28497 (N_28497,N_21004,N_20510);
nor U28498 (N_28498,N_24193,N_23089);
nand U28499 (N_28499,N_21886,N_23570);
xor U28500 (N_28500,N_20507,N_23431);
and U28501 (N_28501,N_20111,N_20550);
and U28502 (N_28502,N_22735,N_21982);
xnor U28503 (N_28503,N_23490,N_24120);
nand U28504 (N_28504,N_22025,N_22311);
nor U28505 (N_28505,N_21514,N_21102);
and U28506 (N_28506,N_24920,N_23059);
nor U28507 (N_28507,N_21133,N_24605);
and U28508 (N_28508,N_23719,N_21104);
xor U28509 (N_28509,N_23211,N_23367);
and U28510 (N_28510,N_20187,N_23663);
and U28511 (N_28511,N_23648,N_23312);
xnor U28512 (N_28512,N_23213,N_21343);
and U28513 (N_28513,N_20026,N_23909);
and U28514 (N_28514,N_24697,N_24216);
nand U28515 (N_28515,N_23842,N_24221);
nand U28516 (N_28516,N_24075,N_23627);
nand U28517 (N_28517,N_21975,N_24118);
xor U28518 (N_28518,N_21533,N_22360);
xnor U28519 (N_28519,N_23874,N_21745);
xor U28520 (N_28520,N_22164,N_24068);
nand U28521 (N_28521,N_22149,N_21344);
nor U28522 (N_28522,N_20379,N_20972);
xor U28523 (N_28523,N_21328,N_24506);
nand U28524 (N_28524,N_23241,N_22640);
nor U28525 (N_28525,N_23549,N_22850);
and U28526 (N_28526,N_21527,N_20169);
and U28527 (N_28527,N_22139,N_21194);
nand U28528 (N_28528,N_20798,N_23134);
nand U28529 (N_28529,N_24546,N_22481);
nor U28530 (N_28530,N_22349,N_21316);
and U28531 (N_28531,N_24596,N_20284);
xnor U28532 (N_28532,N_23561,N_20476);
nand U28533 (N_28533,N_23729,N_23681);
nor U28534 (N_28534,N_22346,N_23863);
nor U28535 (N_28535,N_24256,N_20062);
nor U28536 (N_28536,N_22017,N_23681);
nand U28537 (N_28537,N_23888,N_23492);
or U28538 (N_28538,N_20948,N_21997);
xnor U28539 (N_28539,N_20086,N_22046);
xnor U28540 (N_28540,N_22137,N_24211);
nand U28541 (N_28541,N_24742,N_22922);
or U28542 (N_28542,N_22669,N_23008);
or U28543 (N_28543,N_21750,N_24979);
nand U28544 (N_28544,N_21089,N_23196);
and U28545 (N_28545,N_24106,N_23969);
or U28546 (N_28546,N_20539,N_20752);
nand U28547 (N_28547,N_23316,N_21416);
or U28548 (N_28548,N_21723,N_20496);
nand U28549 (N_28549,N_21141,N_23706);
nor U28550 (N_28550,N_24347,N_24700);
xor U28551 (N_28551,N_21656,N_24094);
or U28552 (N_28552,N_20583,N_20332);
nor U28553 (N_28553,N_20741,N_21736);
nand U28554 (N_28554,N_22092,N_20949);
xor U28555 (N_28555,N_23252,N_22946);
xor U28556 (N_28556,N_21740,N_20657);
or U28557 (N_28557,N_22367,N_24485);
xnor U28558 (N_28558,N_22115,N_22812);
and U28559 (N_28559,N_20023,N_23413);
nand U28560 (N_28560,N_21863,N_21630);
nor U28561 (N_28561,N_20886,N_22516);
and U28562 (N_28562,N_24672,N_22682);
nand U28563 (N_28563,N_23272,N_24149);
or U28564 (N_28564,N_20606,N_23356);
and U28565 (N_28565,N_20553,N_23942);
and U28566 (N_28566,N_20616,N_23799);
nor U28567 (N_28567,N_22420,N_24275);
nand U28568 (N_28568,N_22031,N_20159);
xor U28569 (N_28569,N_20903,N_21602);
xnor U28570 (N_28570,N_24053,N_21435);
and U28571 (N_28571,N_24855,N_20758);
and U28572 (N_28572,N_24261,N_20052);
or U28573 (N_28573,N_20207,N_22611);
nor U28574 (N_28574,N_24535,N_24953);
nor U28575 (N_28575,N_20824,N_23819);
or U28576 (N_28576,N_22968,N_20678);
nor U28577 (N_28577,N_22335,N_22249);
xor U28578 (N_28578,N_24078,N_20224);
or U28579 (N_28579,N_24539,N_21492);
and U28580 (N_28580,N_22292,N_20931);
xor U28581 (N_28581,N_22345,N_21226);
or U28582 (N_28582,N_22027,N_22323);
xnor U28583 (N_28583,N_22798,N_22144);
or U28584 (N_28584,N_20647,N_24656);
nand U28585 (N_28585,N_22362,N_24808);
and U28586 (N_28586,N_22605,N_24705);
or U28587 (N_28587,N_24159,N_24808);
or U28588 (N_28588,N_21183,N_23623);
nor U28589 (N_28589,N_23314,N_20305);
xor U28590 (N_28590,N_20528,N_23532);
and U28591 (N_28591,N_20007,N_20295);
nand U28592 (N_28592,N_20027,N_23503);
or U28593 (N_28593,N_22125,N_20454);
nand U28594 (N_28594,N_20396,N_24161);
nand U28595 (N_28595,N_21914,N_23326);
or U28596 (N_28596,N_20774,N_23670);
nor U28597 (N_28597,N_23075,N_24101);
xor U28598 (N_28598,N_22728,N_20053);
nor U28599 (N_28599,N_23100,N_22773);
nor U28600 (N_28600,N_20902,N_23048);
nand U28601 (N_28601,N_21343,N_22872);
and U28602 (N_28602,N_24463,N_22121);
nand U28603 (N_28603,N_22056,N_21392);
xnor U28604 (N_28604,N_23616,N_20353);
nor U28605 (N_28605,N_24337,N_20052);
and U28606 (N_28606,N_24416,N_20945);
nand U28607 (N_28607,N_24449,N_23208);
nor U28608 (N_28608,N_23405,N_21615);
nor U28609 (N_28609,N_21718,N_21844);
or U28610 (N_28610,N_24528,N_23814);
xor U28611 (N_28611,N_22931,N_24122);
or U28612 (N_28612,N_20045,N_22226);
or U28613 (N_28613,N_21264,N_23894);
xor U28614 (N_28614,N_20785,N_21912);
and U28615 (N_28615,N_22675,N_21033);
nand U28616 (N_28616,N_21036,N_22889);
nand U28617 (N_28617,N_20377,N_21682);
or U28618 (N_28618,N_21451,N_22212);
nand U28619 (N_28619,N_23339,N_22639);
nand U28620 (N_28620,N_24300,N_20442);
and U28621 (N_28621,N_22337,N_24117);
xnor U28622 (N_28622,N_20465,N_24272);
nor U28623 (N_28623,N_21480,N_24730);
nand U28624 (N_28624,N_20102,N_23064);
or U28625 (N_28625,N_21452,N_24242);
nor U28626 (N_28626,N_21612,N_20260);
or U28627 (N_28627,N_20773,N_23780);
nand U28628 (N_28628,N_23247,N_22815);
xnor U28629 (N_28629,N_23133,N_24384);
xnor U28630 (N_28630,N_23592,N_23297);
and U28631 (N_28631,N_23580,N_20856);
or U28632 (N_28632,N_22777,N_23240);
xor U28633 (N_28633,N_23318,N_21481);
or U28634 (N_28634,N_20833,N_22336);
nand U28635 (N_28635,N_23392,N_21124);
nand U28636 (N_28636,N_21772,N_21720);
nor U28637 (N_28637,N_21676,N_21513);
xnor U28638 (N_28638,N_21420,N_20609);
or U28639 (N_28639,N_21008,N_23211);
or U28640 (N_28640,N_22129,N_22337);
xnor U28641 (N_28641,N_22544,N_24196);
or U28642 (N_28642,N_24971,N_20417);
or U28643 (N_28643,N_23074,N_23130);
nand U28644 (N_28644,N_21555,N_20847);
nand U28645 (N_28645,N_24833,N_21290);
or U28646 (N_28646,N_20497,N_22794);
and U28647 (N_28647,N_20489,N_23761);
or U28648 (N_28648,N_24662,N_20056);
and U28649 (N_28649,N_22958,N_20814);
or U28650 (N_28650,N_22138,N_22404);
nand U28651 (N_28651,N_24314,N_20835);
nand U28652 (N_28652,N_23539,N_22701);
xnor U28653 (N_28653,N_21052,N_24326);
or U28654 (N_28654,N_22919,N_24782);
nor U28655 (N_28655,N_22920,N_24704);
nand U28656 (N_28656,N_23195,N_22997);
and U28657 (N_28657,N_22246,N_20281);
nand U28658 (N_28658,N_24195,N_22166);
or U28659 (N_28659,N_21106,N_21677);
and U28660 (N_28660,N_23137,N_23062);
nand U28661 (N_28661,N_22542,N_23988);
nand U28662 (N_28662,N_24711,N_24255);
and U28663 (N_28663,N_24221,N_24925);
nor U28664 (N_28664,N_20340,N_22048);
xnor U28665 (N_28665,N_23795,N_22991);
nor U28666 (N_28666,N_24902,N_23118);
xnor U28667 (N_28667,N_23214,N_22456);
or U28668 (N_28668,N_22734,N_23987);
or U28669 (N_28669,N_22180,N_22996);
xor U28670 (N_28670,N_23018,N_20960);
nor U28671 (N_28671,N_21299,N_23385);
nand U28672 (N_28672,N_20483,N_24717);
xnor U28673 (N_28673,N_22895,N_22024);
nor U28674 (N_28674,N_22764,N_24649);
or U28675 (N_28675,N_21944,N_22153);
or U28676 (N_28676,N_24039,N_22822);
xor U28677 (N_28677,N_22084,N_23653);
nor U28678 (N_28678,N_22269,N_22171);
and U28679 (N_28679,N_21671,N_20728);
nor U28680 (N_28680,N_22024,N_20551);
or U28681 (N_28681,N_22498,N_20555);
nor U28682 (N_28682,N_22871,N_23036);
or U28683 (N_28683,N_24915,N_22051);
or U28684 (N_28684,N_24293,N_24031);
nand U28685 (N_28685,N_21122,N_22996);
nor U28686 (N_28686,N_22484,N_22246);
xor U28687 (N_28687,N_24230,N_22661);
xnor U28688 (N_28688,N_24729,N_24023);
or U28689 (N_28689,N_24706,N_21333);
or U28690 (N_28690,N_21275,N_20927);
nor U28691 (N_28691,N_20749,N_20213);
or U28692 (N_28692,N_22928,N_21732);
nand U28693 (N_28693,N_24573,N_21881);
or U28694 (N_28694,N_24001,N_22107);
nor U28695 (N_28695,N_21036,N_20288);
or U28696 (N_28696,N_23604,N_21985);
and U28697 (N_28697,N_20157,N_20271);
or U28698 (N_28698,N_21205,N_22364);
nand U28699 (N_28699,N_21858,N_22038);
nand U28700 (N_28700,N_20661,N_23562);
nand U28701 (N_28701,N_20146,N_20192);
nand U28702 (N_28702,N_23579,N_22255);
nand U28703 (N_28703,N_20221,N_24337);
xor U28704 (N_28704,N_22641,N_21682);
or U28705 (N_28705,N_22800,N_20457);
or U28706 (N_28706,N_20812,N_21099);
nand U28707 (N_28707,N_21714,N_22133);
nor U28708 (N_28708,N_20789,N_23929);
or U28709 (N_28709,N_21326,N_21911);
nand U28710 (N_28710,N_22399,N_21338);
xor U28711 (N_28711,N_23398,N_24109);
nand U28712 (N_28712,N_20548,N_24387);
nand U28713 (N_28713,N_22460,N_21962);
and U28714 (N_28714,N_23576,N_24603);
nor U28715 (N_28715,N_23342,N_23062);
xnor U28716 (N_28716,N_23507,N_23561);
and U28717 (N_28717,N_24897,N_21183);
xnor U28718 (N_28718,N_24553,N_23283);
nand U28719 (N_28719,N_24743,N_22318);
nor U28720 (N_28720,N_24587,N_21064);
xnor U28721 (N_28721,N_20816,N_21308);
and U28722 (N_28722,N_20450,N_23505);
nor U28723 (N_28723,N_23128,N_20318);
and U28724 (N_28724,N_24089,N_23975);
or U28725 (N_28725,N_24336,N_20182);
xor U28726 (N_28726,N_24471,N_23421);
or U28727 (N_28727,N_22151,N_21210);
xnor U28728 (N_28728,N_23622,N_24723);
or U28729 (N_28729,N_21566,N_21635);
nand U28730 (N_28730,N_23764,N_20695);
and U28731 (N_28731,N_24586,N_20298);
nand U28732 (N_28732,N_24684,N_24084);
nor U28733 (N_28733,N_20438,N_21081);
or U28734 (N_28734,N_20145,N_22596);
and U28735 (N_28735,N_22721,N_20331);
nand U28736 (N_28736,N_20116,N_23976);
and U28737 (N_28737,N_20226,N_24487);
nand U28738 (N_28738,N_24013,N_20800);
and U28739 (N_28739,N_21515,N_22343);
nor U28740 (N_28740,N_20149,N_22908);
and U28741 (N_28741,N_20450,N_20397);
nand U28742 (N_28742,N_23104,N_21392);
or U28743 (N_28743,N_21278,N_20945);
and U28744 (N_28744,N_20838,N_24171);
xor U28745 (N_28745,N_20782,N_23626);
and U28746 (N_28746,N_21397,N_22913);
and U28747 (N_28747,N_24860,N_21634);
xnor U28748 (N_28748,N_21794,N_23083);
nand U28749 (N_28749,N_20536,N_24754);
nand U28750 (N_28750,N_21351,N_20551);
nand U28751 (N_28751,N_20255,N_23652);
or U28752 (N_28752,N_21874,N_24042);
and U28753 (N_28753,N_21858,N_23451);
xnor U28754 (N_28754,N_21408,N_22631);
and U28755 (N_28755,N_20878,N_21471);
and U28756 (N_28756,N_21778,N_22570);
nand U28757 (N_28757,N_24031,N_22418);
and U28758 (N_28758,N_23382,N_22721);
and U28759 (N_28759,N_24091,N_24336);
or U28760 (N_28760,N_24329,N_23547);
and U28761 (N_28761,N_20910,N_24610);
nor U28762 (N_28762,N_24802,N_23010);
nor U28763 (N_28763,N_23137,N_23095);
xnor U28764 (N_28764,N_20558,N_20208);
nand U28765 (N_28765,N_22666,N_23357);
and U28766 (N_28766,N_20150,N_22493);
nand U28767 (N_28767,N_20568,N_21684);
and U28768 (N_28768,N_21733,N_22309);
xor U28769 (N_28769,N_24322,N_21325);
nand U28770 (N_28770,N_20729,N_24234);
or U28771 (N_28771,N_21858,N_20861);
xor U28772 (N_28772,N_23510,N_23453);
nand U28773 (N_28773,N_22597,N_21320);
and U28774 (N_28774,N_24342,N_22087);
xor U28775 (N_28775,N_21188,N_20106);
and U28776 (N_28776,N_20877,N_24565);
nand U28777 (N_28777,N_24065,N_24014);
xnor U28778 (N_28778,N_22951,N_22208);
nor U28779 (N_28779,N_20683,N_22533);
nand U28780 (N_28780,N_23635,N_23801);
or U28781 (N_28781,N_22993,N_23305);
or U28782 (N_28782,N_20719,N_20744);
nor U28783 (N_28783,N_23798,N_23627);
and U28784 (N_28784,N_21665,N_24890);
or U28785 (N_28785,N_20127,N_21623);
nor U28786 (N_28786,N_20212,N_21586);
nor U28787 (N_28787,N_24353,N_23257);
or U28788 (N_28788,N_23136,N_21284);
and U28789 (N_28789,N_20977,N_22699);
nor U28790 (N_28790,N_20991,N_22393);
nor U28791 (N_28791,N_22982,N_22482);
or U28792 (N_28792,N_23931,N_24684);
nor U28793 (N_28793,N_21477,N_24854);
and U28794 (N_28794,N_20745,N_22661);
nor U28795 (N_28795,N_24651,N_21539);
or U28796 (N_28796,N_22780,N_24620);
xor U28797 (N_28797,N_22464,N_22488);
or U28798 (N_28798,N_21679,N_24884);
xor U28799 (N_28799,N_23536,N_23391);
nand U28800 (N_28800,N_23086,N_21581);
nand U28801 (N_28801,N_22571,N_22708);
nand U28802 (N_28802,N_20139,N_23957);
nand U28803 (N_28803,N_22990,N_22861);
nand U28804 (N_28804,N_22447,N_20060);
nor U28805 (N_28805,N_23637,N_24902);
xnor U28806 (N_28806,N_22847,N_20572);
nand U28807 (N_28807,N_20646,N_22637);
nor U28808 (N_28808,N_24798,N_23208);
nor U28809 (N_28809,N_21154,N_22371);
nand U28810 (N_28810,N_21013,N_21960);
or U28811 (N_28811,N_24369,N_20488);
nor U28812 (N_28812,N_20040,N_20123);
and U28813 (N_28813,N_22788,N_23197);
xor U28814 (N_28814,N_20249,N_24019);
nand U28815 (N_28815,N_22847,N_23721);
and U28816 (N_28816,N_22503,N_23508);
or U28817 (N_28817,N_20596,N_23534);
and U28818 (N_28818,N_23789,N_24218);
and U28819 (N_28819,N_24647,N_20263);
nor U28820 (N_28820,N_24665,N_24406);
nor U28821 (N_28821,N_22830,N_20321);
nor U28822 (N_28822,N_24570,N_24664);
or U28823 (N_28823,N_21074,N_23411);
xnor U28824 (N_28824,N_21537,N_23061);
and U28825 (N_28825,N_21021,N_20383);
xnor U28826 (N_28826,N_24475,N_23368);
xor U28827 (N_28827,N_21999,N_20814);
nor U28828 (N_28828,N_20956,N_24068);
nand U28829 (N_28829,N_24632,N_23529);
nand U28830 (N_28830,N_23248,N_21464);
nor U28831 (N_28831,N_24817,N_20808);
and U28832 (N_28832,N_23293,N_24364);
nor U28833 (N_28833,N_23926,N_24664);
or U28834 (N_28834,N_23042,N_24685);
xnor U28835 (N_28835,N_20115,N_20920);
or U28836 (N_28836,N_24198,N_20851);
or U28837 (N_28837,N_24007,N_23706);
nor U28838 (N_28838,N_23023,N_23732);
nor U28839 (N_28839,N_20184,N_22736);
xor U28840 (N_28840,N_24659,N_23252);
nor U28841 (N_28841,N_20665,N_24127);
nand U28842 (N_28842,N_22228,N_20526);
xnor U28843 (N_28843,N_21236,N_20735);
xnor U28844 (N_28844,N_20658,N_23520);
nor U28845 (N_28845,N_20558,N_21184);
or U28846 (N_28846,N_24084,N_20740);
or U28847 (N_28847,N_23420,N_22337);
nand U28848 (N_28848,N_22826,N_20041);
xor U28849 (N_28849,N_23592,N_22367);
and U28850 (N_28850,N_24634,N_24165);
nor U28851 (N_28851,N_21504,N_24275);
and U28852 (N_28852,N_20204,N_21758);
nor U28853 (N_28853,N_20367,N_21447);
and U28854 (N_28854,N_22334,N_21409);
xor U28855 (N_28855,N_24385,N_21913);
nand U28856 (N_28856,N_24162,N_22731);
and U28857 (N_28857,N_23904,N_21621);
nor U28858 (N_28858,N_22259,N_22894);
nor U28859 (N_28859,N_21181,N_23964);
and U28860 (N_28860,N_24982,N_20145);
and U28861 (N_28861,N_21324,N_22548);
xor U28862 (N_28862,N_20541,N_20125);
nand U28863 (N_28863,N_24286,N_22752);
nor U28864 (N_28864,N_21522,N_21619);
nor U28865 (N_28865,N_21236,N_20973);
nor U28866 (N_28866,N_20738,N_21968);
or U28867 (N_28867,N_23873,N_21590);
xor U28868 (N_28868,N_21018,N_20348);
xor U28869 (N_28869,N_24346,N_22484);
or U28870 (N_28870,N_24242,N_24831);
xnor U28871 (N_28871,N_24777,N_23444);
nor U28872 (N_28872,N_20880,N_22522);
xnor U28873 (N_28873,N_23035,N_24422);
and U28874 (N_28874,N_24885,N_22060);
xor U28875 (N_28875,N_20452,N_22812);
xnor U28876 (N_28876,N_24567,N_22904);
nor U28877 (N_28877,N_20541,N_20108);
and U28878 (N_28878,N_22422,N_23024);
nor U28879 (N_28879,N_21635,N_20442);
xnor U28880 (N_28880,N_24294,N_21330);
and U28881 (N_28881,N_21732,N_21581);
xnor U28882 (N_28882,N_24395,N_23870);
nand U28883 (N_28883,N_24778,N_21223);
xor U28884 (N_28884,N_24465,N_21078);
nor U28885 (N_28885,N_20880,N_24489);
and U28886 (N_28886,N_22080,N_20606);
and U28887 (N_28887,N_21296,N_22111);
nand U28888 (N_28888,N_22015,N_24219);
xnor U28889 (N_28889,N_20141,N_22963);
xor U28890 (N_28890,N_24801,N_20079);
nand U28891 (N_28891,N_22698,N_20130);
nand U28892 (N_28892,N_23823,N_22703);
xor U28893 (N_28893,N_24070,N_21420);
and U28894 (N_28894,N_22705,N_20782);
nor U28895 (N_28895,N_23233,N_24250);
or U28896 (N_28896,N_21567,N_23993);
nand U28897 (N_28897,N_20040,N_22305);
and U28898 (N_28898,N_20878,N_24250);
and U28899 (N_28899,N_21174,N_22430);
nand U28900 (N_28900,N_21835,N_22121);
xor U28901 (N_28901,N_20853,N_24181);
and U28902 (N_28902,N_23490,N_22951);
xor U28903 (N_28903,N_22730,N_24627);
nor U28904 (N_28904,N_24441,N_20341);
and U28905 (N_28905,N_24606,N_22476);
xnor U28906 (N_28906,N_20260,N_22592);
xnor U28907 (N_28907,N_21884,N_22274);
and U28908 (N_28908,N_20304,N_21445);
nand U28909 (N_28909,N_20428,N_22237);
and U28910 (N_28910,N_24172,N_21076);
and U28911 (N_28911,N_24486,N_20655);
and U28912 (N_28912,N_21274,N_22263);
or U28913 (N_28913,N_24005,N_24822);
xnor U28914 (N_28914,N_20425,N_20150);
xnor U28915 (N_28915,N_22044,N_20756);
nor U28916 (N_28916,N_22183,N_24081);
and U28917 (N_28917,N_21565,N_21784);
or U28918 (N_28918,N_22409,N_23444);
xnor U28919 (N_28919,N_20757,N_24902);
nor U28920 (N_28920,N_24785,N_21826);
or U28921 (N_28921,N_21389,N_24795);
and U28922 (N_28922,N_21857,N_21548);
xor U28923 (N_28923,N_23327,N_23868);
nand U28924 (N_28924,N_21652,N_21662);
nor U28925 (N_28925,N_23745,N_23295);
xnor U28926 (N_28926,N_20197,N_20526);
nand U28927 (N_28927,N_22584,N_20499);
xor U28928 (N_28928,N_21015,N_21048);
xnor U28929 (N_28929,N_20715,N_22172);
or U28930 (N_28930,N_22560,N_24773);
nand U28931 (N_28931,N_20722,N_22772);
nand U28932 (N_28932,N_24680,N_21848);
nand U28933 (N_28933,N_22326,N_24209);
and U28934 (N_28934,N_22413,N_21781);
and U28935 (N_28935,N_24054,N_24961);
or U28936 (N_28936,N_24667,N_21269);
xnor U28937 (N_28937,N_24561,N_21695);
nor U28938 (N_28938,N_22442,N_21590);
and U28939 (N_28939,N_24567,N_22858);
or U28940 (N_28940,N_23339,N_24025);
nor U28941 (N_28941,N_21861,N_20964);
and U28942 (N_28942,N_23030,N_22370);
nor U28943 (N_28943,N_20895,N_23774);
or U28944 (N_28944,N_24799,N_24838);
and U28945 (N_28945,N_23441,N_20491);
nand U28946 (N_28946,N_23127,N_20953);
xor U28947 (N_28947,N_23096,N_20772);
xnor U28948 (N_28948,N_23299,N_23489);
xor U28949 (N_28949,N_22846,N_20513);
nand U28950 (N_28950,N_23646,N_22685);
or U28951 (N_28951,N_20057,N_22241);
nor U28952 (N_28952,N_20031,N_23164);
or U28953 (N_28953,N_20020,N_23392);
and U28954 (N_28954,N_24552,N_24633);
or U28955 (N_28955,N_24795,N_20129);
xor U28956 (N_28956,N_20896,N_23342);
xnor U28957 (N_28957,N_20654,N_20610);
nor U28958 (N_28958,N_20234,N_21890);
nand U28959 (N_28959,N_23401,N_21445);
nand U28960 (N_28960,N_21983,N_23477);
and U28961 (N_28961,N_22318,N_21079);
nand U28962 (N_28962,N_21674,N_20962);
xnor U28963 (N_28963,N_20016,N_22508);
xor U28964 (N_28964,N_20000,N_22592);
and U28965 (N_28965,N_24612,N_20202);
nor U28966 (N_28966,N_20965,N_23131);
nand U28967 (N_28967,N_22150,N_24154);
nand U28968 (N_28968,N_21470,N_20050);
nand U28969 (N_28969,N_24644,N_22981);
xnor U28970 (N_28970,N_20702,N_23573);
or U28971 (N_28971,N_20612,N_22911);
nor U28972 (N_28972,N_24408,N_20409);
nand U28973 (N_28973,N_21079,N_21371);
or U28974 (N_28974,N_22511,N_21202);
or U28975 (N_28975,N_23351,N_23257);
and U28976 (N_28976,N_21531,N_20172);
and U28977 (N_28977,N_22342,N_20276);
nand U28978 (N_28978,N_24626,N_21929);
and U28979 (N_28979,N_22341,N_23361);
nor U28980 (N_28980,N_23462,N_22362);
nor U28981 (N_28981,N_21902,N_24618);
xnor U28982 (N_28982,N_24190,N_22094);
or U28983 (N_28983,N_24481,N_24606);
nor U28984 (N_28984,N_22273,N_20400);
nor U28985 (N_28985,N_21985,N_23797);
or U28986 (N_28986,N_20418,N_24788);
or U28987 (N_28987,N_21307,N_22315);
or U28988 (N_28988,N_20874,N_21239);
nor U28989 (N_28989,N_24103,N_20458);
or U28990 (N_28990,N_24480,N_22823);
nor U28991 (N_28991,N_24619,N_22424);
nand U28992 (N_28992,N_23924,N_23446);
nand U28993 (N_28993,N_20578,N_20405);
nor U28994 (N_28994,N_21054,N_22732);
and U28995 (N_28995,N_21540,N_20508);
nor U28996 (N_28996,N_21921,N_21846);
xnor U28997 (N_28997,N_22373,N_20933);
nor U28998 (N_28998,N_24633,N_23786);
and U28999 (N_28999,N_20780,N_24328);
or U29000 (N_29000,N_22649,N_24409);
and U29001 (N_29001,N_24227,N_23695);
and U29002 (N_29002,N_21803,N_21509);
or U29003 (N_29003,N_24805,N_21302);
xnor U29004 (N_29004,N_23521,N_21042);
nand U29005 (N_29005,N_23398,N_20305);
nor U29006 (N_29006,N_22893,N_20712);
and U29007 (N_29007,N_23339,N_22229);
nor U29008 (N_29008,N_22007,N_21811);
nor U29009 (N_29009,N_22857,N_20455);
or U29010 (N_29010,N_23466,N_23866);
or U29011 (N_29011,N_21434,N_22176);
or U29012 (N_29012,N_20014,N_20588);
nand U29013 (N_29013,N_23563,N_22863);
nor U29014 (N_29014,N_22899,N_24426);
xor U29015 (N_29015,N_22426,N_21111);
or U29016 (N_29016,N_23378,N_23747);
nand U29017 (N_29017,N_21198,N_24534);
or U29018 (N_29018,N_20286,N_24040);
and U29019 (N_29019,N_23117,N_23832);
xor U29020 (N_29020,N_22585,N_23229);
nor U29021 (N_29021,N_22825,N_24107);
xnor U29022 (N_29022,N_20620,N_23820);
nor U29023 (N_29023,N_21856,N_22329);
or U29024 (N_29024,N_23139,N_21429);
nor U29025 (N_29025,N_24760,N_22951);
nand U29026 (N_29026,N_23020,N_23309);
and U29027 (N_29027,N_22532,N_22458);
and U29028 (N_29028,N_20679,N_20180);
or U29029 (N_29029,N_20593,N_23885);
or U29030 (N_29030,N_23990,N_22276);
nor U29031 (N_29031,N_23379,N_21513);
and U29032 (N_29032,N_20492,N_23054);
and U29033 (N_29033,N_23909,N_24458);
and U29034 (N_29034,N_23675,N_23268);
nor U29035 (N_29035,N_21733,N_20917);
xnor U29036 (N_29036,N_20397,N_23781);
nor U29037 (N_29037,N_20814,N_23595);
or U29038 (N_29038,N_24410,N_23106);
or U29039 (N_29039,N_21807,N_24728);
and U29040 (N_29040,N_24241,N_24274);
or U29041 (N_29041,N_22507,N_24840);
or U29042 (N_29042,N_21701,N_22672);
and U29043 (N_29043,N_21505,N_24707);
nand U29044 (N_29044,N_22962,N_20301);
or U29045 (N_29045,N_23847,N_24222);
nor U29046 (N_29046,N_23079,N_24152);
nor U29047 (N_29047,N_21965,N_23743);
or U29048 (N_29048,N_21575,N_21016);
or U29049 (N_29049,N_24962,N_22627);
and U29050 (N_29050,N_22581,N_20370);
or U29051 (N_29051,N_20623,N_21743);
nand U29052 (N_29052,N_23101,N_20160);
nand U29053 (N_29053,N_21148,N_23500);
nor U29054 (N_29054,N_21808,N_21292);
and U29055 (N_29055,N_23737,N_22918);
nand U29056 (N_29056,N_23971,N_20086);
nor U29057 (N_29057,N_24046,N_24978);
and U29058 (N_29058,N_24250,N_22411);
nor U29059 (N_29059,N_21184,N_23258);
nand U29060 (N_29060,N_24202,N_21298);
and U29061 (N_29061,N_20367,N_23759);
xor U29062 (N_29062,N_24690,N_20823);
or U29063 (N_29063,N_21789,N_20474);
xor U29064 (N_29064,N_22187,N_23288);
or U29065 (N_29065,N_24896,N_22805);
or U29066 (N_29066,N_23074,N_23638);
nor U29067 (N_29067,N_22274,N_21910);
xor U29068 (N_29068,N_20966,N_23348);
or U29069 (N_29069,N_20304,N_22437);
nor U29070 (N_29070,N_24705,N_21015);
nand U29071 (N_29071,N_20321,N_23396);
and U29072 (N_29072,N_22742,N_22844);
or U29073 (N_29073,N_20263,N_20682);
or U29074 (N_29074,N_22455,N_23889);
xor U29075 (N_29075,N_23001,N_23069);
or U29076 (N_29076,N_20509,N_24585);
and U29077 (N_29077,N_24971,N_21602);
and U29078 (N_29078,N_23645,N_24736);
or U29079 (N_29079,N_21682,N_22305);
xnor U29080 (N_29080,N_24387,N_22869);
nand U29081 (N_29081,N_24967,N_22226);
nand U29082 (N_29082,N_20747,N_20341);
xnor U29083 (N_29083,N_23036,N_22118);
nand U29084 (N_29084,N_20299,N_20626);
or U29085 (N_29085,N_21000,N_21661);
or U29086 (N_29086,N_21556,N_22020);
nand U29087 (N_29087,N_20874,N_22111);
nor U29088 (N_29088,N_20300,N_20196);
nor U29089 (N_29089,N_22062,N_21383);
xor U29090 (N_29090,N_22511,N_24768);
or U29091 (N_29091,N_22707,N_20721);
xnor U29092 (N_29092,N_23070,N_22974);
nand U29093 (N_29093,N_24494,N_21952);
nor U29094 (N_29094,N_23720,N_22357);
nor U29095 (N_29095,N_20963,N_22748);
and U29096 (N_29096,N_22755,N_21627);
nor U29097 (N_29097,N_24827,N_22209);
or U29098 (N_29098,N_21007,N_21474);
nand U29099 (N_29099,N_22805,N_21057);
xor U29100 (N_29100,N_24325,N_24387);
nor U29101 (N_29101,N_20784,N_24522);
nand U29102 (N_29102,N_21254,N_21290);
and U29103 (N_29103,N_22455,N_23660);
nand U29104 (N_29104,N_20985,N_20276);
or U29105 (N_29105,N_24229,N_20653);
nor U29106 (N_29106,N_24239,N_21110);
or U29107 (N_29107,N_21362,N_20429);
or U29108 (N_29108,N_21413,N_21054);
or U29109 (N_29109,N_24645,N_21556);
and U29110 (N_29110,N_22581,N_24679);
or U29111 (N_29111,N_24623,N_20477);
nor U29112 (N_29112,N_21458,N_24435);
and U29113 (N_29113,N_24163,N_22140);
xor U29114 (N_29114,N_20977,N_23552);
nor U29115 (N_29115,N_22382,N_22408);
xnor U29116 (N_29116,N_20183,N_20344);
xor U29117 (N_29117,N_23603,N_20458);
nor U29118 (N_29118,N_21033,N_21234);
nand U29119 (N_29119,N_23212,N_22850);
nor U29120 (N_29120,N_22718,N_24339);
nor U29121 (N_29121,N_23916,N_23679);
and U29122 (N_29122,N_23129,N_22200);
nor U29123 (N_29123,N_23934,N_21158);
and U29124 (N_29124,N_21949,N_23606);
nand U29125 (N_29125,N_21835,N_20600);
and U29126 (N_29126,N_20639,N_20823);
xnor U29127 (N_29127,N_22505,N_23825);
xor U29128 (N_29128,N_21216,N_24091);
nand U29129 (N_29129,N_23986,N_23414);
xor U29130 (N_29130,N_23404,N_20683);
nand U29131 (N_29131,N_20913,N_21627);
xnor U29132 (N_29132,N_24825,N_20299);
nor U29133 (N_29133,N_20493,N_24556);
nor U29134 (N_29134,N_24359,N_21900);
and U29135 (N_29135,N_23991,N_24088);
nand U29136 (N_29136,N_22076,N_21355);
xor U29137 (N_29137,N_23060,N_21007);
and U29138 (N_29138,N_21145,N_20282);
and U29139 (N_29139,N_22158,N_23285);
nor U29140 (N_29140,N_21722,N_22236);
nand U29141 (N_29141,N_24131,N_21785);
nand U29142 (N_29142,N_23622,N_20156);
or U29143 (N_29143,N_21263,N_20019);
or U29144 (N_29144,N_20864,N_21993);
xnor U29145 (N_29145,N_20718,N_21811);
and U29146 (N_29146,N_21031,N_20758);
and U29147 (N_29147,N_21303,N_23077);
nand U29148 (N_29148,N_22135,N_23252);
nand U29149 (N_29149,N_20773,N_23074);
and U29150 (N_29150,N_24380,N_22462);
nand U29151 (N_29151,N_20684,N_21929);
nand U29152 (N_29152,N_23314,N_21478);
and U29153 (N_29153,N_22967,N_24977);
nand U29154 (N_29154,N_22341,N_23231);
nand U29155 (N_29155,N_21112,N_24151);
or U29156 (N_29156,N_22008,N_21293);
and U29157 (N_29157,N_23553,N_24896);
nor U29158 (N_29158,N_24640,N_22980);
xor U29159 (N_29159,N_22065,N_21512);
nor U29160 (N_29160,N_22439,N_20707);
or U29161 (N_29161,N_20507,N_24881);
nand U29162 (N_29162,N_20735,N_23295);
nor U29163 (N_29163,N_23455,N_20277);
nand U29164 (N_29164,N_24658,N_23066);
nor U29165 (N_29165,N_24155,N_24002);
nand U29166 (N_29166,N_23744,N_24227);
or U29167 (N_29167,N_20113,N_22224);
xnor U29168 (N_29168,N_20840,N_20448);
and U29169 (N_29169,N_23452,N_22090);
nor U29170 (N_29170,N_24550,N_20937);
nand U29171 (N_29171,N_20899,N_23213);
or U29172 (N_29172,N_22929,N_20073);
nor U29173 (N_29173,N_24570,N_24082);
xor U29174 (N_29174,N_24541,N_24251);
or U29175 (N_29175,N_20024,N_22364);
xnor U29176 (N_29176,N_24005,N_21010);
nand U29177 (N_29177,N_23505,N_21053);
nor U29178 (N_29178,N_24196,N_21238);
nor U29179 (N_29179,N_20235,N_24729);
nor U29180 (N_29180,N_20578,N_22013);
xnor U29181 (N_29181,N_21524,N_21245);
xor U29182 (N_29182,N_24067,N_22623);
or U29183 (N_29183,N_23389,N_22974);
xor U29184 (N_29184,N_21117,N_20471);
or U29185 (N_29185,N_22820,N_21747);
xnor U29186 (N_29186,N_23764,N_22510);
nand U29187 (N_29187,N_21231,N_21485);
xor U29188 (N_29188,N_22922,N_24916);
or U29189 (N_29189,N_22843,N_24188);
nand U29190 (N_29190,N_23623,N_22629);
nor U29191 (N_29191,N_23137,N_21189);
xnor U29192 (N_29192,N_24754,N_21134);
xnor U29193 (N_29193,N_20661,N_20687);
and U29194 (N_29194,N_22087,N_23341);
and U29195 (N_29195,N_23609,N_23697);
and U29196 (N_29196,N_23262,N_24604);
nand U29197 (N_29197,N_22577,N_22763);
nor U29198 (N_29198,N_20103,N_23098);
and U29199 (N_29199,N_21154,N_24595);
or U29200 (N_29200,N_23374,N_21477);
nand U29201 (N_29201,N_20945,N_20215);
xor U29202 (N_29202,N_24591,N_22962);
nor U29203 (N_29203,N_21836,N_24135);
nor U29204 (N_29204,N_21018,N_21600);
and U29205 (N_29205,N_20726,N_22502);
and U29206 (N_29206,N_22601,N_22755);
nor U29207 (N_29207,N_23948,N_23433);
or U29208 (N_29208,N_21813,N_23374);
xnor U29209 (N_29209,N_20571,N_24946);
xnor U29210 (N_29210,N_24696,N_21407);
nor U29211 (N_29211,N_23812,N_24575);
xnor U29212 (N_29212,N_21243,N_24281);
nand U29213 (N_29213,N_23206,N_24598);
or U29214 (N_29214,N_24592,N_21136);
nand U29215 (N_29215,N_24189,N_24245);
xnor U29216 (N_29216,N_24464,N_24617);
nand U29217 (N_29217,N_21081,N_24157);
xnor U29218 (N_29218,N_24253,N_21716);
nor U29219 (N_29219,N_21936,N_23750);
nor U29220 (N_29220,N_21854,N_24685);
xor U29221 (N_29221,N_21985,N_20239);
nor U29222 (N_29222,N_21518,N_22177);
nor U29223 (N_29223,N_24731,N_21351);
xnor U29224 (N_29224,N_22645,N_23572);
xnor U29225 (N_29225,N_24819,N_24364);
and U29226 (N_29226,N_21695,N_22367);
and U29227 (N_29227,N_21411,N_22456);
and U29228 (N_29228,N_22448,N_22895);
or U29229 (N_29229,N_24559,N_23681);
or U29230 (N_29230,N_20800,N_22788);
and U29231 (N_29231,N_24177,N_24537);
or U29232 (N_29232,N_24561,N_20581);
or U29233 (N_29233,N_22214,N_23012);
or U29234 (N_29234,N_22589,N_20071);
nand U29235 (N_29235,N_22972,N_20958);
xnor U29236 (N_29236,N_22680,N_23545);
nand U29237 (N_29237,N_20625,N_23979);
nor U29238 (N_29238,N_21563,N_24899);
xnor U29239 (N_29239,N_21093,N_24073);
nand U29240 (N_29240,N_24572,N_22955);
nand U29241 (N_29241,N_22529,N_20191);
xor U29242 (N_29242,N_22975,N_20434);
or U29243 (N_29243,N_20635,N_23928);
xnor U29244 (N_29244,N_22818,N_21960);
xnor U29245 (N_29245,N_24403,N_23184);
nand U29246 (N_29246,N_20480,N_21380);
and U29247 (N_29247,N_24829,N_20446);
and U29248 (N_29248,N_21733,N_20845);
nor U29249 (N_29249,N_23416,N_20077);
xnor U29250 (N_29250,N_23376,N_22437);
nor U29251 (N_29251,N_24589,N_22295);
or U29252 (N_29252,N_20035,N_22761);
xnor U29253 (N_29253,N_21548,N_22224);
nand U29254 (N_29254,N_22514,N_24123);
or U29255 (N_29255,N_22442,N_20163);
and U29256 (N_29256,N_22750,N_24245);
nand U29257 (N_29257,N_24981,N_24409);
xor U29258 (N_29258,N_21619,N_22915);
nor U29259 (N_29259,N_24118,N_22338);
and U29260 (N_29260,N_20112,N_24619);
and U29261 (N_29261,N_24717,N_24892);
xor U29262 (N_29262,N_23799,N_23391);
nand U29263 (N_29263,N_22786,N_20855);
nor U29264 (N_29264,N_23108,N_23051);
and U29265 (N_29265,N_23950,N_24117);
nand U29266 (N_29266,N_21903,N_22660);
nand U29267 (N_29267,N_23194,N_22911);
xnor U29268 (N_29268,N_22426,N_23418);
and U29269 (N_29269,N_23073,N_21080);
xor U29270 (N_29270,N_24188,N_24126);
and U29271 (N_29271,N_24286,N_24723);
xor U29272 (N_29272,N_24243,N_23371);
or U29273 (N_29273,N_23831,N_20670);
xnor U29274 (N_29274,N_21958,N_23526);
and U29275 (N_29275,N_21829,N_20902);
nand U29276 (N_29276,N_22864,N_20579);
xor U29277 (N_29277,N_20454,N_22757);
or U29278 (N_29278,N_23674,N_24625);
or U29279 (N_29279,N_24233,N_20342);
nand U29280 (N_29280,N_23135,N_20531);
and U29281 (N_29281,N_21675,N_21926);
or U29282 (N_29282,N_21379,N_23388);
and U29283 (N_29283,N_20880,N_21515);
nor U29284 (N_29284,N_21685,N_23287);
nand U29285 (N_29285,N_20391,N_24165);
xnor U29286 (N_29286,N_21895,N_22949);
nand U29287 (N_29287,N_23815,N_23776);
or U29288 (N_29288,N_21161,N_23489);
or U29289 (N_29289,N_22260,N_24547);
nand U29290 (N_29290,N_22561,N_23055);
and U29291 (N_29291,N_24222,N_23615);
nor U29292 (N_29292,N_20695,N_22384);
nand U29293 (N_29293,N_23977,N_22398);
nand U29294 (N_29294,N_23115,N_22487);
or U29295 (N_29295,N_24731,N_22625);
nor U29296 (N_29296,N_23640,N_22291);
nor U29297 (N_29297,N_22705,N_20317);
xor U29298 (N_29298,N_20660,N_21434);
or U29299 (N_29299,N_24937,N_21793);
xor U29300 (N_29300,N_23684,N_21701);
nand U29301 (N_29301,N_24479,N_22008);
nor U29302 (N_29302,N_24987,N_22307);
xor U29303 (N_29303,N_21010,N_22028);
and U29304 (N_29304,N_22809,N_22374);
nand U29305 (N_29305,N_23249,N_23455);
and U29306 (N_29306,N_22035,N_21634);
nor U29307 (N_29307,N_20578,N_24136);
nand U29308 (N_29308,N_22232,N_24227);
or U29309 (N_29309,N_21155,N_20765);
and U29310 (N_29310,N_20450,N_20605);
xor U29311 (N_29311,N_21189,N_20097);
and U29312 (N_29312,N_20950,N_21190);
xor U29313 (N_29313,N_23491,N_20038);
and U29314 (N_29314,N_24433,N_23950);
and U29315 (N_29315,N_22826,N_23588);
or U29316 (N_29316,N_23059,N_20473);
xnor U29317 (N_29317,N_23916,N_20494);
xor U29318 (N_29318,N_21434,N_21197);
and U29319 (N_29319,N_21868,N_23203);
nor U29320 (N_29320,N_23197,N_24206);
or U29321 (N_29321,N_20052,N_20013);
xor U29322 (N_29322,N_22412,N_23197);
nand U29323 (N_29323,N_21798,N_20153);
nor U29324 (N_29324,N_23933,N_22925);
xnor U29325 (N_29325,N_21106,N_20399);
xnor U29326 (N_29326,N_21456,N_22133);
or U29327 (N_29327,N_23820,N_23293);
xor U29328 (N_29328,N_22578,N_22295);
nand U29329 (N_29329,N_23239,N_23573);
nor U29330 (N_29330,N_20667,N_24453);
nor U29331 (N_29331,N_24878,N_24314);
nand U29332 (N_29332,N_23593,N_22753);
or U29333 (N_29333,N_23699,N_23905);
nand U29334 (N_29334,N_24818,N_24931);
or U29335 (N_29335,N_23464,N_24389);
nor U29336 (N_29336,N_23357,N_22663);
nand U29337 (N_29337,N_22711,N_22977);
or U29338 (N_29338,N_23785,N_20700);
nand U29339 (N_29339,N_23379,N_20057);
xor U29340 (N_29340,N_21926,N_24435);
and U29341 (N_29341,N_21329,N_20174);
and U29342 (N_29342,N_24976,N_24864);
nand U29343 (N_29343,N_24497,N_22598);
nor U29344 (N_29344,N_21917,N_24002);
xnor U29345 (N_29345,N_21795,N_24406);
and U29346 (N_29346,N_23518,N_20180);
nor U29347 (N_29347,N_23173,N_24599);
and U29348 (N_29348,N_24232,N_21193);
nand U29349 (N_29349,N_22065,N_20840);
nand U29350 (N_29350,N_22103,N_24948);
xnor U29351 (N_29351,N_21352,N_20045);
xnor U29352 (N_29352,N_23519,N_22356);
nor U29353 (N_29353,N_23723,N_22576);
nor U29354 (N_29354,N_20582,N_24409);
xor U29355 (N_29355,N_22482,N_22337);
nand U29356 (N_29356,N_23941,N_23506);
nand U29357 (N_29357,N_22766,N_21235);
xor U29358 (N_29358,N_20785,N_21887);
or U29359 (N_29359,N_21416,N_21721);
nand U29360 (N_29360,N_22491,N_22599);
or U29361 (N_29361,N_24462,N_20761);
nor U29362 (N_29362,N_24060,N_24248);
xor U29363 (N_29363,N_24873,N_20258);
nor U29364 (N_29364,N_20576,N_22277);
nor U29365 (N_29365,N_20634,N_21805);
xnor U29366 (N_29366,N_23455,N_22525);
nor U29367 (N_29367,N_24470,N_21289);
or U29368 (N_29368,N_21576,N_20920);
nor U29369 (N_29369,N_24552,N_21821);
and U29370 (N_29370,N_22948,N_21333);
nor U29371 (N_29371,N_23131,N_22145);
xnor U29372 (N_29372,N_23104,N_22117);
or U29373 (N_29373,N_21622,N_22291);
nand U29374 (N_29374,N_24244,N_24729);
xor U29375 (N_29375,N_23258,N_24268);
or U29376 (N_29376,N_20585,N_23251);
xor U29377 (N_29377,N_24427,N_21175);
and U29378 (N_29378,N_24843,N_24690);
nor U29379 (N_29379,N_24940,N_23954);
nor U29380 (N_29380,N_23776,N_20589);
or U29381 (N_29381,N_21081,N_20055);
and U29382 (N_29382,N_20456,N_23892);
xnor U29383 (N_29383,N_24674,N_24432);
or U29384 (N_29384,N_22212,N_23986);
or U29385 (N_29385,N_20396,N_24514);
and U29386 (N_29386,N_23192,N_24722);
xor U29387 (N_29387,N_21557,N_22620);
nand U29388 (N_29388,N_20286,N_24090);
nand U29389 (N_29389,N_20645,N_20392);
and U29390 (N_29390,N_22096,N_21469);
xor U29391 (N_29391,N_20319,N_21755);
and U29392 (N_29392,N_20924,N_22836);
or U29393 (N_29393,N_23515,N_23103);
nand U29394 (N_29394,N_21682,N_20604);
nand U29395 (N_29395,N_24012,N_21622);
nor U29396 (N_29396,N_23466,N_23744);
nor U29397 (N_29397,N_22665,N_20755);
and U29398 (N_29398,N_24837,N_21075);
and U29399 (N_29399,N_24399,N_21374);
nor U29400 (N_29400,N_21791,N_22959);
or U29401 (N_29401,N_20601,N_23300);
xnor U29402 (N_29402,N_22930,N_20265);
nand U29403 (N_29403,N_23236,N_22662);
nor U29404 (N_29404,N_20602,N_23514);
xor U29405 (N_29405,N_22579,N_21624);
xor U29406 (N_29406,N_22557,N_22580);
or U29407 (N_29407,N_20697,N_23736);
xnor U29408 (N_29408,N_23043,N_24556);
or U29409 (N_29409,N_20433,N_20822);
xor U29410 (N_29410,N_23213,N_21228);
or U29411 (N_29411,N_20789,N_24732);
nor U29412 (N_29412,N_23618,N_22061);
nand U29413 (N_29413,N_23093,N_20809);
and U29414 (N_29414,N_23220,N_23470);
and U29415 (N_29415,N_24758,N_20850);
or U29416 (N_29416,N_22479,N_20149);
nor U29417 (N_29417,N_22244,N_23317);
nor U29418 (N_29418,N_24628,N_24235);
xnor U29419 (N_29419,N_22014,N_23712);
or U29420 (N_29420,N_24363,N_23186);
xnor U29421 (N_29421,N_20977,N_23865);
xor U29422 (N_29422,N_22323,N_24016);
or U29423 (N_29423,N_21863,N_23534);
nor U29424 (N_29424,N_23261,N_24515);
nor U29425 (N_29425,N_22739,N_24503);
or U29426 (N_29426,N_23086,N_20262);
and U29427 (N_29427,N_24711,N_22328);
or U29428 (N_29428,N_22053,N_23024);
xnor U29429 (N_29429,N_23120,N_22632);
nand U29430 (N_29430,N_23745,N_23036);
or U29431 (N_29431,N_21222,N_22268);
nor U29432 (N_29432,N_20313,N_24488);
and U29433 (N_29433,N_22164,N_23710);
nor U29434 (N_29434,N_24847,N_20692);
nand U29435 (N_29435,N_24704,N_22025);
or U29436 (N_29436,N_23373,N_21002);
nor U29437 (N_29437,N_21910,N_23150);
nand U29438 (N_29438,N_20839,N_21268);
and U29439 (N_29439,N_23388,N_24274);
nand U29440 (N_29440,N_24191,N_24950);
and U29441 (N_29441,N_21878,N_22690);
nor U29442 (N_29442,N_24631,N_20721);
and U29443 (N_29443,N_21136,N_22654);
and U29444 (N_29444,N_21734,N_20677);
and U29445 (N_29445,N_22903,N_22863);
nor U29446 (N_29446,N_23093,N_23427);
xor U29447 (N_29447,N_20215,N_20950);
or U29448 (N_29448,N_22072,N_24454);
or U29449 (N_29449,N_22494,N_24928);
xor U29450 (N_29450,N_24887,N_24798);
and U29451 (N_29451,N_23656,N_20102);
nor U29452 (N_29452,N_21132,N_23729);
and U29453 (N_29453,N_24962,N_24924);
or U29454 (N_29454,N_23343,N_24254);
and U29455 (N_29455,N_20158,N_21183);
nand U29456 (N_29456,N_22366,N_23470);
xnor U29457 (N_29457,N_24550,N_21117);
xnor U29458 (N_29458,N_21009,N_23415);
or U29459 (N_29459,N_22100,N_20479);
and U29460 (N_29460,N_24088,N_22532);
nor U29461 (N_29461,N_24041,N_20783);
nand U29462 (N_29462,N_22087,N_22890);
nor U29463 (N_29463,N_20695,N_22491);
nor U29464 (N_29464,N_21687,N_23107);
and U29465 (N_29465,N_23445,N_23338);
and U29466 (N_29466,N_24564,N_24995);
nand U29467 (N_29467,N_22006,N_24793);
or U29468 (N_29468,N_20752,N_22436);
nand U29469 (N_29469,N_24228,N_24704);
and U29470 (N_29470,N_24892,N_24598);
nor U29471 (N_29471,N_24637,N_22034);
nand U29472 (N_29472,N_22848,N_23847);
xor U29473 (N_29473,N_23486,N_22185);
nand U29474 (N_29474,N_22527,N_22773);
nor U29475 (N_29475,N_20899,N_22947);
nor U29476 (N_29476,N_22303,N_20453);
or U29477 (N_29477,N_20723,N_24974);
nand U29478 (N_29478,N_22510,N_24808);
and U29479 (N_29479,N_21264,N_24152);
or U29480 (N_29480,N_21942,N_22291);
xor U29481 (N_29481,N_21783,N_23782);
or U29482 (N_29482,N_24143,N_22978);
and U29483 (N_29483,N_23578,N_21756);
xor U29484 (N_29484,N_23344,N_20117);
and U29485 (N_29485,N_24965,N_24859);
nor U29486 (N_29486,N_23606,N_23621);
or U29487 (N_29487,N_20061,N_21619);
nand U29488 (N_29488,N_24316,N_21466);
nor U29489 (N_29489,N_24000,N_23390);
or U29490 (N_29490,N_21562,N_21420);
and U29491 (N_29491,N_23914,N_21964);
and U29492 (N_29492,N_23916,N_23508);
xor U29493 (N_29493,N_24467,N_22755);
xor U29494 (N_29494,N_23107,N_24511);
nor U29495 (N_29495,N_21464,N_22452);
nand U29496 (N_29496,N_21304,N_21114);
and U29497 (N_29497,N_22191,N_23072);
nand U29498 (N_29498,N_21985,N_23018);
nor U29499 (N_29499,N_20905,N_23120);
nand U29500 (N_29500,N_24174,N_24401);
or U29501 (N_29501,N_20524,N_24502);
nor U29502 (N_29502,N_24153,N_21300);
and U29503 (N_29503,N_20541,N_24711);
nor U29504 (N_29504,N_20108,N_22499);
or U29505 (N_29505,N_23021,N_23677);
nand U29506 (N_29506,N_20900,N_20454);
xnor U29507 (N_29507,N_23891,N_23807);
or U29508 (N_29508,N_21833,N_22756);
or U29509 (N_29509,N_21830,N_21037);
and U29510 (N_29510,N_20480,N_20077);
nand U29511 (N_29511,N_21386,N_23004);
xnor U29512 (N_29512,N_24093,N_22048);
and U29513 (N_29513,N_20652,N_23940);
nand U29514 (N_29514,N_24627,N_20150);
xnor U29515 (N_29515,N_22772,N_24470);
nand U29516 (N_29516,N_20359,N_24538);
nand U29517 (N_29517,N_20625,N_23171);
and U29518 (N_29518,N_22833,N_24014);
xor U29519 (N_29519,N_20851,N_20300);
and U29520 (N_29520,N_21280,N_23098);
nand U29521 (N_29521,N_20345,N_22178);
and U29522 (N_29522,N_22294,N_21824);
nand U29523 (N_29523,N_20014,N_23599);
and U29524 (N_29524,N_23166,N_20861);
and U29525 (N_29525,N_22580,N_21914);
nand U29526 (N_29526,N_21599,N_23825);
nand U29527 (N_29527,N_24716,N_20742);
nand U29528 (N_29528,N_24250,N_22065);
and U29529 (N_29529,N_20259,N_24042);
nor U29530 (N_29530,N_20304,N_23234);
nor U29531 (N_29531,N_21488,N_21979);
or U29532 (N_29532,N_20231,N_22552);
nand U29533 (N_29533,N_20270,N_21010);
nand U29534 (N_29534,N_21976,N_24263);
or U29535 (N_29535,N_24249,N_20956);
and U29536 (N_29536,N_24961,N_20585);
or U29537 (N_29537,N_22794,N_20786);
xor U29538 (N_29538,N_20788,N_22955);
or U29539 (N_29539,N_22586,N_24989);
or U29540 (N_29540,N_20222,N_21591);
xnor U29541 (N_29541,N_22202,N_20275);
and U29542 (N_29542,N_23627,N_22343);
or U29543 (N_29543,N_24273,N_20206);
xnor U29544 (N_29544,N_20861,N_24545);
and U29545 (N_29545,N_23242,N_23753);
xnor U29546 (N_29546,N_24663,N_21700);
xnor U29547 (N_29547,N_23529,N_22706);
nand U29548 (N_29548,N_22980,N_20228);
or U29549 (N_29549,N_23540,N_22059);
nor U29550 (N_29550,N_23139,N_20117);
nor U29551 (N_29551,N_23440,N_20974);
xor U29552 (N_29552,N_24641,N_20138);
nor U29553 (N_29553,N_23934,N_20886);
nand U29554 (N_29554,N_22508,N_22003);
xor U29555 (N_29555,N_21923,N_23802);
xor U29556 (N_29556,N_23386,N_21815);
or U29557 (N_29557,N_21666,N_24691);
or U29558 (N_29558,N_20893,N_21712);
nor U29559 (N_29559,N_20178,N_21756);
nor U29560 (N_29560,N_24125,N_24477);
or U29561 (N_29561,N_22489,N_23436);
or U29562 (N_29562,N_20734,N_21308);
and U29563 (N_29563,N_22329,N_24111);
nand U29564 (N_29564,N_21093,N_23363);
or U29565 (N_29565,N_23880,N_20265);
and U29566 (N_29566,N_21278,N_22736);
nor U29567 (N_29567,N_21930,N_24595);
nand U29568 (N_29568,N_21594,N_22279);
and U29569 (N_29569,N_22299,N_24370);
nor U29570 (N_29570,N_23007,N_22244);
nand U29571 (N_29571,N_22257,N_22712);
nor U29572 (N_29572,N_21627,N_23823);
nor U29573 (N_29573,N_24524,N_23607);
xnor U29574 (N_29574,N_24791,N_22513);
nand U29575 (N_29575,N_22128,N_24556);
nand U29576 (N_29576,N_20704,N_21110);
or U29577 (N_29577,N_20985,N_21865);
or U29578 (N_29578,N_23403,N_20530);
or U29579 (N_29579,N_21123,N_21618);
or U29580 (N_29580,N_21538,N_22763);
nor U29581 (N_29581,N_23807,N_23887);
xnor U29582 (N_29582,N_22279,N_24625);
or U29583 (N_29583,N_22090,N_20179);
xnor U29584 (N_29584,N_20251,N_24018);
and U29585 (N_29585,N_21345,N_24795);
nor U29586 (N_29586,N_20081,N_20642);
or U29587 (N_29587,N_23462,N_23629);
nand U29588 (N_29588,N_22787,N_23926);
xnor U29589 (N_29589,N_20681,N_23547);
and U29590 (N_29590,N_22227,N_20337);
or U29591 (N_29591,N_20616,N_22781);
nor U29592 (N_29592,N_21525,N_20104);
xor U29593 (N_29593,N_21481,N_20551);
nor U29594 (N_29594,N_24802,N_21936);
or U29595 (N_29595,N_23676,N_23117);
xor U29596 (N_29596,N_20972,N_22614);
or U29597 (N_29597,N_21000,N_22759);
or U29598 (N_29598,N_24667,N_22980);
and U29599 (N_29599,N_24258,N_20315);
nor U29600 (N_29600,N_21508,N_24401);
nand U29601 (N_29601,N_24518,N_22852);
nor U29602 (N_29602,N_23346,N_20054);
xor U29603 (N_29603,N_24075,N_23355);
nor U29604 (N_29604,N_21632,N_23261);
or U29605 (N_29605,N_20090,N_23817);
and U29606 (N_29606,N_20973,N_20991);
xor U29607 (N_29607,N_22110,N_21029);
nor U29608 (N_29608,N_22566,N_21528);
nand U29609 (N_29609,N_24031,N_22008);
and U29610 (N_29610,N_23007,N_23760);
and U29611 (N_29611,N_20299,N_23316);
or U29612 (N_29612,N_22934,N_22788);
and U29613 (N_29613,N_23550,N_22760);
or U29614 (N_29614,N_23978,N_21778);
nand U29615 (N_29615,N_24215,N_22492);
or U29616 (N_29616,N_24070,N_21418);
nor U29617 (N_29617,N_21535,N_20812);
or U29618 (N_29618,N_20965,N_21549);
xnor U29619 (N_29619,N_21701,N_21315);
xnor U29620 (N_29620,N_22750,N_21845);
and U29621 (N_29621,N_23705,N_21961);
or U29622 (N_29622,N_24110,N_21538);
nand U29623 (N_29623,N_21703,N_24125);
nand U29624 (N_29624,N_24859,N_21781);
and U29625 (N_29625,N_23247,N_23538);
xor U29626 (N_29626,N_21181,N_22139);
and U29627 (N_29627,N_24906,N_21157);
xor U29628 (N_29628,N_23916,N_21287);
or U29629 (N_29629,N_22961,N_24839);
nand U29630 (N_29630,N_21092,N_20907);
xnor U29631 (N_29631,N_20547,N_23796);
or U29632 (N_29632,N_21325,N_21442);
or U29633 (N_29633,N_21571,N_23024);
nand U29634 (N_29634,N_23774,N_22051);
nand U29635 (N_29635,N_21147,N_23129);
xor U29636 (N_29636,N_20409,N_22891);
or U29637 (N_29637,N_20951,N_22279);
or U29638 (N_29638,N_21812,N_21920);
and U29639 (N_29639,N_23636,N_20559);
and U29640 (N_29640,N_24887,N_24608);
or U29641 (N_29641,N_21585,N_20549);
xnor U29642 (N_29642,N_22699,N_21265);
or U29643 (N_29643,N_21546,N_24423);
nand U29644 (N_29644,N_21402,N_22676);
nand U29645 (N_29645,N_21273,N_24346);
xnor U29646 (N_29646,N_23414,N_22629);
nor U29647 (N_29647,N_20795,N_24965);
nand U29648 (N_29648,N_21521,N_24458);
xor U29649 (N_29649,N_20803,N_24326);
or U29650 (N_29650,N_23428,N_20137);
nand U29651 (N_29651,N_21021,N_20476);
or U29652 (N_29652,N_24824,N_22660);
nand U29653 (N_29653,N_24172,N_21995);
xor U29654 (N_29654,N_20917,N_24892);
nor U29655 (N_29655,N_23813,N_22437);
nand U29656 (N_29656,N_24056,N_22520);
nor U29657 (N_29657,N_23207,N_22540);
xnor U29658 (N_29658,N_22742,N_24472);
and U29659 (N_29659,N_20739,N_23686);
and U29660 (N_29660,N_23363,N_24729);
or U29661 (N_29661,N_22747,N_22724);
xor U29662 (N_29662,N_23622,N_20532);
or U29663 (N_29663,N_23963,N_23437);
xor U29664 (N_29664,N_20249,N_20616);
nor U29665 (N_29665,N_23959,N_23512);
nor U29666 (N_29666,N_21907,N_22159);
nor U29667 (N_29667,N_21931,N_24688);
nand U29668 (N_29668,N_20917,N_21940);
xor U29669 (N_29669,N_21412,N_24881);
xor U29670 (N_29670,N_20557,N_22963);
nor U29671 (N_29671,N_24784,N_21461);
nor U29672 (N_29672,N_21991,N_20142);
nor U29673 (N_29673,N_23220,N_20232);
nand U29674 (N_29674,N_21579,N_21821);
nand U29675 (N_29675,N_21721,N_24549);
nor U29676 (N_29676,N_22428,N_23939);
nor U29677 (N_29677,N_24027,N_22305);
nand U29678 (N_29678,N_22864,N_20094);
or U29679 (N_29679,N_23881,N_20637);
and U29680 (N_29680,N_24487,N_20366);
and U29681 (N_29681,N_20911,N_24310);
nor U29682 (N_29682,N_21162,N_21712);
nand U29683 (N_29683,N_23826,N_21710);
or U29684 (N_29684,N_22223,N_21160);
nand U29685 (N_29685,N_24470,N_23938);
nand U29686 (N_29686,N_24724,N_21707);
nand U29687 (N_29687,N_23554,N_20781);
and U29688 (N_29688,N_22898,N_24469);
xor U29689 (N_29689,N_24659,N_20531);
nor U29690 (N_29690,N_22194,N_21439);
xor U29691 (N_29691,N_21591,N_23632);
nor U29692 (N_29692,N_22700,N_21660);
nand U29693 (N_29693,N_21441,N_20892);
or U29694 (N_29694,N_20049,N_21624);
nor U29695 (N_29695,N_23347,N_22834);
and U29696 (N_29696,N_20971,N_24610);
and U29697 (N_29697,N_23030,N_23831);
and U29698 (N_29698,N_21343,N_21902);
xor U29699 (N_29699,N_24510,N_23863);
nor U29700 (N_29700,N_20016,N_23834);
nor U29701 (N_29701,N_21094,N_23517);
and U29702 (N_29702,N_22827,N_21525);
and U29703 (N_29703,N_23789,N_21245);
nand U29704 (N_29704,N_23026,N_24287);
xnor U29705 (N_29705,N_22808,N_20181);
nand U29706 (N_29706,N_20244,N_20800);
or U29707 (N_29707,N_22453,N_23822);
and U29708 (N_29708,N_22835,N_20315);
nand U29709 (N_29709,N_21482,N_20813);
nand U29710 (N_29710,N_21655,N_24482);
nor U29711 (N_29711,N_22885,N_21437);
nor U29712 (N_29712,N_21934,N_23498);
xnor U29713 (N_29713,N_23672,N_20149);
nor U29714 (N_29714,N_22872,N_20490);
or U29715 (N_29715,N_20862,N_23614);
and U29716 (N_29716,N_22807,N_23192);
or U29717 (N_29717,N_24784,N_20702);
or U29718 (N_29718,N_21744,N_24995);
nand U29719 (N_29719,N_21892,N_21879);
nor U29720 (N_29720,N_23195,N_21923);
or U29721 (N_29721,N_22497,N_22708);
xor U29722 (N_29722,N_22809,N_22822);
and U29723 (N_29723,N_24327,N_23631);
or U29724 (N_29724,N_22037,N_21087);
nor U29725 (N_29725,N_23937,N_21842);
nand U29726 (N_29726,N_23715,N_23423);
and U29727 (N_29727,N_21983,N_22655);
or U29728 (N_29728,N_20835,N_24084);
xor U29729 (N_29729,N_22806,N_20334);
nor U29730 (N_29730,N_22188,N_22838);
or U29731 (N_29731,N_20734,N_23700);
nor U29732 (N_29732,N_23569,N_21413);
and U29733 (N_29733,N_24536,N_22803);
or U29734 (N_29734,N_22094,N_20730);
xnor U29735 (N_29735,N_22367,N_20389);
or U29736 (N_29736,N_23673,N_21925);
nand U29737 (N_29737,N_20635,N_22187);
and U29738 (N_29738,N_24610,N_22771);
and U29739 (N_29739,N_22381,N_21179);
xor U29740 (N_29740,N_21712,N_22768);
nor U29741 (N_29741,N_21478,N_21740);
nor U29742 (N_29742,N_21663,N_20990);
xnor U29743 (N_29743,N_20469,N_22653);
or U29744 (N_29744,N_24302,N_21281);
or U29745 (N_29745,N_23931,N_20689);
or U29746 (N_29746,N_20820,N_24636);
xor U29747 (N_29747,N_24799,N_20481);
xnor U29748 (N_29748,N_21294,N_22497);
nor U29749 (N_29749,N_20703,N_21738);
xnor U29750 (N_29750,N_22881,N_23924);
nor U29751 (N_29751,N_20692,N_21374);
xnor U29752 (N_29752,N_21471,N_21082);
and U29753 (N_29753,N_24496,N_24270);
xnor U29754 (N_29754,N_22448,N_24850);
or U29755 (N_29755,N_23082,N_21139);
and U29756 (N_29756,N_22744,N_20795);
xnor U29757 (N_29757,N_24166,N_23249);
or U29758 (N_29758,N_24549,N_21719);
nand U29759 (N_29759,N_24175,N_20038);
and U29760 (N_29760,N_24699,N_22880);
xor U29761 (N_29761,N_23318,N_24887);
and U29762 (N_29762,N_22461,N_20192);
xor U29763 (N_29763,N_20835,N_20459);
or U29764 (N_29764,N_20748,N_22184);
xnor U29765 (N_29765,N_23186,N_23658);
xor U29766 (N_29766,N_24853,N_23867);
and U29767 (N_29767,N_22890,N_22299);
or U29768 (N_29768,N_21946,N_21893);
nor U29769 (N_29769,N_21850,N_22689);
xnor U29770 (N_29770,N_22334,N_24318);
or U29771 (N_29771,N_23866,N_23062);
xor U29772 (N_29772,N_22860,N_21516);
or U29773 (N_29773,N_23327,N_21711);
and U29774 (N_29774,N_21877,N_24279);
nor U29775 (N_29775,N_24057,N_23666);
or U29776 (N_29776,N_22881,N_24556);
xnor U29777 (N_29777,N_24243,N_20123);
nor U29778 (N_29778,N_23243,N_22730);
nor U29779 (N_29779,N_23685,N_21640);
or U29780 (N_29780,N_23177,N_22386);
nand U29781 (N_29781,N_22326,N_21671);
or U29782 (N_29782,N_22667,N_22767);
xnor U29783 (N_29783,N_21541,N_24546);
or U29784 (N_29784,N_24761,N_23802);
nor U29785 (N_29785,N_20104,N_22788);
nand U29786 (N_29786,N_22637,N_21652);
nor U29787 (N_29787,N_20685,N_23477);
or U29788 (N_29788,N_23616,N_20442);
and U29789 (N_29789,N_24602,N_23058);
xor U29790 (N_29790,N_23591,N_20582);
nand U29791 (N_29791,N_20025,N_21060);
and U29792 (N_29792,N_20756,N_20642);
nor U29793 (N_29793,N_23834,N_20642);
or U29794 (N_29794,N_21823,N_24381);
or U29795 (N_29795,N_21746,N_24955);
nor U29796 (N_29796,N_22992,N_22235);
nand U29797 (N_29797,N_24602,N_24773);
nor U29798 (N_29798,N_21461,N_23528);
nand U29799 (N_29799,N_22776,N_23958);
nand U29800 (N_29800,N_21543,N_23771);
nand U29801 (N_29801,N_22370,N_23351);
xor U29802 (N_29802,N_22558,N_21859);
nand U29803 (N_29803,N_20263,N_24071);
xor U29804 (N_29804,N_23858,N_22881);
nor U29805 (N_29805,N_24139,N_21790);
nor U29806 (N_29806,N_24510,N_23139);
or U29807 (N_29807,N_20177,N_23415);
xor U29808 (N_29808,N_24044,N_21668);
and U29809 (N_29809,N_23863,N_22990);
and U29810 (N_29810,N_21701,N_24720);
or U29811 (N_29811,N_22445,N_21182);
and U29812 (N_29812,N_21630,N_24571);
and U29813 (N_29813,N_22939,N_22309);
nor U29814 (N_29814,N_23231,N_22731);
or U29815 (N_29815,N_23855,N_23520);
and U29816 (N_29816,N_23992,N_23896);
nand U29817 (N_29817,N_23089,N_21283);
nand U29818 (N_29818,N_24167,N_22592);
and U29819 (N_29819,N_22220,N_21667);
and U29820 (N_29820,N_22627,N_21087);
or U29821 (N_29821,N_24390,N_22245);
nor U29822 (N_29822,N_24332,N_22463);
nand U29823 (N_29823,N_20151,N_20489);
xor U29824 (N_29824,N_21486,N_20278);
xor U29825 (N_29825,N_22702,N_22307);
or U29826 (N_29826,N_22095,N_21862);
or U29827 (N_29827,N_23745,N_24844);
xnor U29828 (N_29828,N_22059,N_21714);
or U29829 (N_29829,N_23427,N_24112);
xnor U29830 (N_29830,N_22432,N_22832);
and U29831 (N_29831,N_20591,N_22181);
or U29832 (N_29832,N_23955,N_24162);
nor U29833 (N_29833,N_24490,N_20309);
or U29834 (N_29834,N_20703,N_22569);
or U29835 (N_29835,N_21316,N_23893);
nor U29836 (N_29836,N_22142,N_24587);
or U29837 (N_29837,N_21631,N_24823);
nand U29838 (N_29838,N_21437,N_22526);
nand U29839 (N_29839,N_22953,N_21744);
or U29840 (N_29840,N_23425,N_23202);
nand U29841 (N_29841,N_21155,N_22753);
xnor U29842 (N_29842,N_22282,N_22767);
nand U29843 (N_29843,N_23569,N_21634);
or U29844 (N_29844,N_20577,N_21731);
xor U29845 (N_29845,N_23965,N_21241);
nor U29846 (N_29846,N_21639,N_24231);
and U29847 (N_29847,N_23242,N_21517);
or U29848 (N_29848,N_20521,N_22884);
nor U29849 (N_29849,N_20783,N_22595);
and U29850 (N_29850,N_21478,N_21258);
xor U29851 (N_29851,N_24006,N_23066);
nand U29852 (N_29852,N_21306,N_24286);
nor U29853 (N_29853,N_24420,N_23131);
nor U29854 (N_29854,N_20966,N_24134);
and U29855 (N_29855,N_24490,N_22858);
nor U29856 (N_29856,N_24489,N_24682);
nand U29857 (N_29857,N_24057,N_22856);
nand U29858 (N_29858,N_20582,N_22075);
nand U29859 (N_29859,N_20454,N_20872);
or U29860 (N_29860,N_24008,N_23056);
nand U29861 (N_29861,N_24187,N_22485);
and U29862 (N_29862,N_21537,N_23127);
and U29863 (N_29863,N_20094,N_22385);
nand U29864 (N_29864,N_24643,N_24939);
and U29865 (N_29865,N_22932,N_20022);
nand U29866 (N_29866,N_24410,N_23132);
nor U29867 (N_29867,N_24808,N_24475);
nand U29868 (N_29868,N_21154,N_22583);
nor U29869 (N_29869,N_24457,N_24638);
or U29870 (N_29870,N_20711,N_24952);
xnor U29871 (N_29871,N_23903,N_24710);
xnor U29872 (N_29872,N_21052,N_24415);
or U29873 (N_29873,N_22032,N_21465);
nor U29874 (N_29874,N_20143,N_20703);
or U29875 (N_29875,N_22895,N_21795);
nor U29876 (N_29876,N_20939,N_24863);
nor U29877 (N_29877,N_24247,N_21357);
and U29878 (N_29878,N_22574,N_20448);
and U29879 (N_29879,N_21217,N_20168);
or U29880 (N_29880,N_23210,N_24144);
nand U29881 (N_29881,N_22083,N_21556);
or U29882 (N_29882,N_21086,N_21460);
nand U29883 (N_29883,N_21377,N_20587);
nand U29884 (N_29884,N_20502,N_24537);
xnor U29885 (N_29885,N_23670,N_20747);
or U29886 (N_29886,N_23168,N_22633);
and U29887 (N_29887,N_23417,N_23583);
and U29888 (N_29888,N_23281,N_21841);
or U29889 (N_29889,N_21449,N_22715);
nor U29890 (N_29890,N_21071,N_24322);
nor U29891 (N_29891,N_23853,N_24190);
or U29892 (N_29892,N_23340,N_21917);
xor U29893 (N_29893,N_20675,N_23802);
or U29894 (N_29894,N_23905,N_22203);
nor U29895 (N_29895,N_21285,N_21793);
xnor U29896 (N_29896,N_21863,N_23051);
and U29897 (N_29897,N_20197,N_24130);
xor U29898 (N_29898,N_21475,N_22518);
or U29899 (N_29899,N_21110,N_21585);
and U29900 (N_29900,N_20060,N_22302);
nand U29901 (N_29901,N_21597,N_20992);
nand U29902 (N_29902,N_20942,N_21844);
and U29903 (N_29903,N_22694,N_22403);
xor U29904 (N_29904,N_22522,N_22246);
or U29905 (N_29905,N_24534,N_20319);
or U29906 (N_29906,N_24551,N_20932);
or U29907 (N_29907,N_22507,N_22635);
xor U29908 (N_29908,N_20101,N_21945);
xor U29909 (N_29909,N_23646,N_20121);
xor U29910 (N_29910,N_24021,N_21697);
nand U29911 (N_29911,N_21890,N_22382);
nand U29912 (N_29912,N_22901,N_20315);
and U29913 (N_29913,N_20535,N_22002);
nand U29914 (N_29914,N_20498,N_20172);
or U29915 (N_29915,N_24381,N_23079);
or U29916 (N_29916,N_22318,N_22111);
nor U29917 (N_29917,N_20969,N_20595);
xnor U29918 (N_29918,N_23064,N_24438);
nand U29919 (N_29919,N_24979,N_20997);
nor U29920 (N_29920,N_22742,N_23894);
nor U29921 (N_29921,N_21499,N_20879);
xor U29922 (N_29922,N_21917,N_21476);
and U29923 (N_29923,N_20201,N_24449);
and U29924 (N_29924,N_21014,N_20188);
nand U29925 (N_29925,N_20266,N_21004);
and U29926 (N_29926,N_24766,N_21753);
nand U29927 (N_29927,N_22620,N_22281);
nor U29928 (N_29928,N_24197,N_24960);
or U29929 (N_29929,N_21675,N_22649);
xnor U29930 (N_29930,N_23722,N_21934);
nor U29931 (N_29931,N_22532,N_24123);
and U29932 (N_29932,N_24634,N_21798);
nor U29933 (N_29933,N_20461,N_22492);
or U29934 (N_29934,N_23947,N_21360);
and U29935 (N_29935,N_22282,N_21336);
and U29936 (N_29936,N_21940,N_23509);
or U29937 (N_29937,N_23665,N_23622);
xnor U29938 (N_29938,N_23679,N_21398);
or U29939 (N_29939,N_24197,N_22708);
and U29940 (N_29940,N_20023,N_20773);
and U29941 (N_29941,N_21001,N_20412);
nand U29942 (N_29942,N_20294,N_23580);
xor U29943 (N_29943,N_21253,N_20508);
or U29944 (N_29944,N_20354,N_22749);
xor U29945 (N_29945,N_21587,N_23674);
nor U29946 (N_29946,N_20488,N_23953);
nand U29947 (N_29947,N_24742,N_24432);
xnor U29948 (N_29948,N_22651,N_21386);
and U29949 (N_29949,N_23075,N_23554);
xor U29950 (N_29950,N_22643,N_22144);
xnor U29951 (N_29951,N_23543,N_20673);
nor U29952 (N_29952,N_20834,N_22346);
nor U29953 (N_29953,N_21425,N_24647);
nor U29954 (N_29954,N_20795,N_23876);
xnor U29955 (N_29955,N_20406,N_21719);
or U29956 (N_29956,N_23480,N_22443);
or U29957 (N_29957,N_23298,N_21275);
nand U29958 (N_29958,N_21623,N_22231);
or U29959 (N_29959,N_21814,N_22500);
or U29960 (N_29960,N_21597,N_21218);
nand U29961 (N_29961,N_24792,N_22490);
or U29962 (N_29962,N_24522,N_22445);
xor U29963 (N_29963,N_21180,N_20553);
nand U29964 (N_29964,N_22622,N_20188);
nor U29965 (N_29965,N_21152,N_20616);
nand U29966 (N_29966,N_20370,N_23018);
and U29967 (N_29967,N_22052,N_22722);
or U29968 (N_29968,N_21606,N_24469);
nand U29969 (N_29969,N_20438,N_21727);
xnor U29970 (N_29970,N_21778,N_22839);
nor U29971 (N_29971,N_24832,N_20162);
nand U29972 (N_29972,N_23541,N_21873);
and U29973 (N_29973,N_21379,N_20666);
and U29974 (N_29974,N_24721,N_23225);
and U29975 (N_29975,N_21269,N_20496);
and U29976 (N_29976,N_23357,N_23100);
xor U29977 (N_29977,N_20368,N_22550);
nor U29978 (N_29978,N_23646,N_24321);
or U29979 (N_29979,N_23357,N_20010);
and U29980 (N_29980,N_21458,N_24980);
nor U29981 (N_29981,N_20213,N_23700);
or U29982 (N_29982,N_20734,N_22637);
nor U29983 (N_29983,N_21227,N_20353);
or U29984 (N_29984,N_20481,N_20154);
and U29985 (N_29985,N_23572,N_23739);
nor U29986 (N_29986,N_24050,N_21203);
xnor U29987 (N_29987,N_24623,N_24359);
nand U29988 (N_29988,N_22287,N_24940);
xor U29989 (N_29989,N_24937,N_23517);
or U29990 (N_29990,N_23832,N_23821);
or U29991 (N_29991,N_23693,N_22030);
nor U29992 (N_29992,N_24747,N_22053);
and U29993 (N_29993,N_20129,N_21895);
and U29994 (N_29994,N_20359,N_23719);
and U29995 (N_29995,N_20529,N_23623);
and U29996 (N_29996,N_20086,N_21414);
nor U29997 (N_29997,N_23267,N_20251);
nor U29998 (N_29998,N_22329,N_24447);
or U29999 (N_29999,N_21380,N_22664);
and U30000 (N_30000,N_28329,N_27607);
xnor U30001 (N_30001,N_28897,N_25851);
or U30002 (N_30002,N_29332,N_27022);
nor U30003 (N_30003,N_29930,N_25921);
xnor U30004 (N_30004,N_27576,N_29000);
nor U30005 (N_30005,N_25421,N_25539);
xor U30006 (N_30006,N_29391,N_29133);
nand U30007 (N_30007,N_29182,N_28709);
and U30008 (N_30008,N_25487,N_29272);
or U30009 (N_30009,N_26588,N_25123);
and U30010 (N_30010,N_29890,N_29501);
and U30011 (N_30011,N_25357,N_25246);
nor U30012 (N_30012,N_26900,N_25391);
nand U30013 (N_30013,N_25644,N_27541);
xnor U30014 (N_30014,N_29657,N_27561);
nand U30015 (N_30015,N_29028,N_27106);
xor U30016 (N_30016,N_26997,N_27830);
and U30017 (N_30017,N_29454,N_25871);
and U30018 (N_30018,N_26769,N_27744);
and U30019 (N_30019,N_28664,N_26504);
and U30020 (N_30020,N_25397,N_28227);
or U30021 (N_30021,N_25564,N_25738);
or U30022 (N_30022,N_25625,N_25124);
nor U30023 (N_30023,N_25173,N_29975);
nand U30024 (N_30024,N_28778,N_25719);
xnor U30025 (N_30025,N_29956,N_25418);
nor U30026 (N_30026,N_28049,N_29648);
xor U30027 (N_30027,N_28938,N_25776);
or U30028 (N_30028,N_25009,N_25960);
nor U30029 (N_30029,N_26058,N_29686);
nor U30030 (N_30030,N_29100,N_29216);
xnor U30031 (N_30031,N_26061,N_29345);
nand U30032 (N_30032,N_28679,N_29872);
nor U30033 (N_30033,N_28443,N_28280);
nor U30034 (N_30034,N_28427,N_28405);
nor U30035 (N_30035,N_27874,N_26305);
nor U30036 (N_30036,N_27581,N_29246);
nor U30037 (N_30037,N_28321,N_26816);
nand U30038 (N_30038,N_28170,N_25076);
xnor U30039 (N_30039,N_26282,N_28113);
and U30040 (N_30040,N_26913,N_27345);
or U30041 (N_30041,N_27493,N_27883);
nand U30042 (N_30042,N_25066,N_26520);
nand U30043 (N_30043,N_26136,N_27146);
or U30044 (N_30044,N_28590,N_29409);
nor U30045 (N_30045,N_28392,N_27461);
and U30046 (N_30046,N_26181,N_26856);
xor U30047 (N_30047,N_29072,N_25255);
nor U30048 (N_30048,N_25297,N_28437);
nor U30049 (N_30049,N_25126,N_27954);
nand U30050 (N_30050,N_26435,N_27509);
nor U30051 (N_30051,N_25556,N_28480);
nor U30052 (N_30052,N_27013,N_29421);
and U30053 (N_30053,N_26398,N_26076);
or U30054 (N_30054,N_26985,N_29469);
and U30055 (N_30055,N_28573,N_27439);
xnor U30056 (N_30056,N_27431,N_27846);
or U30057 (N_30057,N_25178,N_29435);
nor U30058 (N_30058,N_26096,N_27807);
or U30059 (N_30059,N_29557,N_26278);
nand U30060 (N_30060,N_25611,N_27520);
nor U30061 (N_30061,N_26855,N_27787);
and U30062 (N_30062,N_25285,N_28109);
nand U30063 (N_30063,N_28757,N_25417);
nor U30064 (N_30064,N_27501,N_28220);
nor U30065 (N_30065,N_27735,N_29467);
nor U30066 (N_30066,N_29418,N_29088);
nor U30067 (N_30067,N_25197,N_29462);
and U30068 (N_30068,N_29154,N_26047);
nand U30069 (N_30069,N_27843,N_28067);
nor U30070 (N_30070,N_28345,N_27546);
xnor U30071 (N_30071,N_25508,N_29430);
xor U30072 (N_30072,N_27241,N_28805);
and U30073 (N_30073,N_27024,N_26902);
or U30074 (N_30074,N_25745,N_27690);
nor U30075 (N_30075,N_29884,N_26568);
nand U30076 (N_30076,N_26409,N_29719);
and U30077 (N_30077,N_29665,N_28568);
nor U30078 (N_30078,N_29453,N_28207);
nand U30079 (N_30079,N_29006,N_28536);
nand U30080 (N_30080,N_28663,N_29024);
or U30081 (N_30081,N_28990,N_27422);
nor U30082 (N_30082,N_26625,N_27869);
and U30083 (N_30083,N_27988,N_27417);
and U30084 (N_30084,N_28712,N_27266);
nor U30085 (N_30085,N_29188,N_26438);
or U30086 (N_30086,N_25732,N_27770);
or U30087 (N_30087,N_27038,N_27108);
and U30088 (N_30088,N_27623,N_26102);
or U30089 (N_30089,N_27223,N_27965);
nor U30090 (N_30090,N_28639,N_26138);
or U30091 (N_30091,N_29228,N_25182);
and U30092 (N_30092,N_29653,N_28434);
nand U30093 (N_30093,N_26035,N_29911);
or U30094 (N_30094,N_29475,N_25744);
nor U30095 (N_30095,N_27238,N_29639);
xnor U30096 (N_30096,N_28241,N_26935);
xnor U30097 (N_30097,N_29477,N_26089);
nor U30098 (N_30098,N_26145,N_27386);
or U30099 (N_30099,N_29023,N_29539);
xnor U30100 (N_30100,N_27357,N_26280);
or U30101 (N_30101,N_25021,N_29715);
xor U30102 (N_30102,N_28159,N_26784);
nor U30103 (N_30103,N_27762,N_27505);
or U30104 (N_30104,N_29160,N_26279);
nor U30105 (N_30105,N_28933,N_26942);
or U30106 (N_30106,N_25504,N_28237);
and U30107 (N_30107,N_29481,N_28126);
or U30108 (N_30108,N_28307,N_25779);
and U30109 (N_30109,N_26992,N_28319);
xnor U30110 (N_30110,N_25687,N_29830);
nor U30111 (N_30111,N_29752,N_27193);
nand U30112 (N_30112,N_27259,N_28470);
xnor U30113 (N_30113,N_25057,N_28406);
nor U30114 (N_30114,N_27851,N_25427);
nor U30115 (N_30115,N_28727,N_26761);
xnor U30116 (N_30116,N_25631,N_28014);
or U30117 (N_30117,N_28649,N_27496);
or U30118 (N_30118,N_28693,N_26502);
xnor U30119 (N_30119,N_28796,N_26969);
nand U30120 (N_30120,N_29874,N_29230);
or U30121 (N_30121,N_28950,N_27902);
and U30122 (N_30122,N_29910,N_25794);
or U30123 (N_30123,N_25437,N_27174);
nand U30124 (N_30124,N_27910,N_29928);
and U30125 (N_30125,N_26898,N_27061);
nor U30126 (N_30126,N_27283,N_25050);
nor U30127 (N_30127,N_28694,N_28128);
or U30128 (N_30128,N_25848,N_27708);
xnor U30129 (N_30129,N_26051,N_25395);
nor U30130 (N_30130,N_29105,N_27254);
and U30131 (N_30131,N_28094,N_26238);
and U30132 (N_30132,N_28048,N_27306);
and U30133 (N_30133,N_26612,N_26890);
and U30134 (N_30134,N_28129,N_26150);
nand U30135 (N_30135,N_27127,N_28070);
xnor U30136 (N_30136,N_29480,N_27327);
nand U30137 (N_30137,N_29732,N_28251);
or U30138 (N_30138,N_26328,N_26283);
nor U30139 (N_30139,N_26836,N_27556);
xor U30140 (N_30140,N_25747,N_28783);
nor U30141 (N_30141,N_26513,N_29035);
nand U30142 (N_30142,N_27229,N_29735);
xnor U30143 (N_30143,N_29738,N_27453);
and U30144 (N_30144,N_26249,N_27483);
or U30145 (N_30145,N_28707,N_29651);
or U30146 (N_30146,N_26731,N_27391);
and U30147 (N_30147,N_27582,N_29399);
xnor U30148 (N_30148,N_25812,N_25345);
xnor U30149 (N_30149,N_29450,N_29753);
nor U30150 (N_30150,N_29168,N_27522);
nor U30151 (N_30151,N_29823,N_27781);
or U30152 (N_30152,N_28389,N_29840);
nor U30153 (N_30153,N_28855,N_28672);
xor U30154 (N_30154,N_25046,N_27957);
xor U30155 (N_30155,N_27815,N_26754);
and U30156 (N_30156,N_27725,N_25193);
nand U30157 (N_30157,N_26814,N_26812);
nand U30158 (N_30158,N_26930,N_28817);
nor U30159 (N_30159,N_28540,N_28487);
or U30160 (N_30160,N_25840,N_25630);
xnor U30161 (N_30161,N_27497,N_26643);
or U30162 (N_30162,N_27432,N_28968);
nor U30163 (N_30163,N_29256,N_26804);
and U30164 (N_30164,N_27868,N_29093);
nand U30165 (N_30165,N_28118,N_26851);
or U30166 (N_30166,N_27151,N_25167);
or U30167 (N_30167,N_28650,N_25484);
nand U30168 (N_30168,N_29565,N_26323);
or U30169 (N_30169,N_27875,N_27399);
or U30170 (N_30170,N_27655,N_26811);
nor U30171 (N_30171,N_26962,N_29184);
xor U30172 (N_30172,N_25331,N_25424);
or U30173 (N_30173,N_26826,N_25927);
xor U30174 (N_30174,N_25224,N_27312);
xnor U30175 (N_30175,N_27699,N_27118);
and U30176 (N_30176,N_25805,N_26426);
and U30177 (N_30177,N_25730,N_26265);
nand U30178 (N_30178,N_28042,N_28833);
or U30179 (N_30179,N_26469,N_26009);
xnor U30180 (N_30180,N_27540,N_29192);
nor U30181 (N_30181,N_28583,N_25992);
xnor U30182 (N_30182,N_25514,N_28815);
xnor U30183 (N_30183,N_25010,N_26715);
or U30184 (N_30184,N_27436,N_29270);
xor U30185 (N_30185,N_25834,N_27754);
or U30186 (N_30186,N_26878,N_29658);
nor U30187 (N_30187,N_28646,N_25324);
xnor U30188 (N_30188,N_29961,N_28748);
or U30189 (N_30189,N_27612,N_25983);
or U30190 (N_30190,N_28006,N_27333);
or U30191 (N_30191,N_28408,N_27308);
nor U30192 (N_30192,N_29948,N_29425);
and U30193 (N_30193,N_28099,N_26941);
nand U30194 (N_30194,N_25451,N_25233);
nand U30195 (N_30195,N_28024,N_25517);
xor U30196 (N_30196,N_28054,N_28386);
nand U30197 (N_30197,N_25646,N_27156);
or U30198 (N_30198,N_29718,N_28019);
and U30199 (N_30199,N_25172,N_27646);
nand U30200 (N_30200,N_25202,N_28597);
or U30201 (N_30201,N_29624,N_25392);
or U30202 (N_30202,N_28073,N_27299);
nand U30203 (N_30203,N_26146,N_29115);
nand U30204 (N_30204,N_26778,N_27008);
and U30205 (N_30205,N_25410,N_27304);
nand U30206 (N_30206,N_28290,N_25238);
nor U30207 (N_30207,N_25617,N_25802);
and U30208 (N_30208,N_28465,N_28656);
and U30209 (N_30209,N_25523,N_28965);
nor U30210 (N_30210,N_29233,N_26362);
xnor U30211 (N_30211,N_29553,N_27588);
and U30212 (N_30212,N_26001,N_28236);
nand U30213 (N_30213,N_25847,N_26149);
xnor U30214 (N_30214,N_26561,N_28840);
nor U30215 (N_30215,N_28885,N_27023);
xnor U30216 (N_30216,N_25203,N_25213);
nor U30217 (N_30217,N_25234,N_25362);
xnor U30218 (N_30218,N_29295,N_25225);
nand U30219 (N_30219,N_29011,N_29380);
nor U30220 (N_30220,N_29713,N_25998);
nor U30221 (N_30221,N_25917,N_25654);
nor U30222 (N_30222,N_25852,N_26662);
or U30223 (N_30223,N_29424,N_25121);
or U30224 (N_30224,N_25304,N_25069);
and U30225 (N_30225,N_28491,N_27185);
nand U30226 (N_30226,N_29936,N_25994);
nand U30227 (N_30227,N_29045,N_29969);
xnor U30228 (N_30228,N_27506,N_26949);
or U30229 (N_30229,N_26335,N_29893);
xor U30230 (N_30230,N_27705,N_25622);
nor U30231 (N_30231,N_28934,N_25912);
nand U30232 (N_30232,N_25715,N_25170);
xnor U30233 (N_30233,N_25416,N_28410);
or U30234 (N_30234,N_25758,N_25907);
or U30235 (N_30235,N_29222,N_28746);
and U30236 (N_30236,N_26522,N_26459);
and U30237 (N_30237,N_29509,N_27911);
xor U30238 (N_30238,N_25598,N_28056);
and U30239 (N_30239,N_26166,N_26555);
nor U30240 (N_30240,N_29009,N_26592);
nand U30241 (N_30241,N_25742,N_29330);
xnor U30242 (N_30242,N_29277,N_26532);
nor U30243 (N_30243,N_25816,N_26195);
and U30244 (N_30244,N_28636,N_29204);
nand U30245 (N_30245,N_27889,N_28806);
nor U30246 (N_30246,N_29153,N_29241);
xor U30247 (N_30247,N_26691,N_29121);
nand U30248 (N_30248,N_28501,N_26671);
and U30249 (N_30249,N_27792,N_29536);
or U30250 (N_30250,N_29073,N_28452);
and U30251 (N_30251,N_27611,N_26611);
xor U30252 (N_30252,N_26553,N_29212);
nor U30253 (N_30253,N_28530,N_25107);
nor U30254 (N_30254,N_25720,N_29808);
xor U30255 (N_30255,N_25181,N_25322);
nand U30256 (N_30256,N_29452,N_29774);
or U30257 (N_30257,N_25078,N_28257);
xnor U30258 (N_30258,N_29263,N_29328);
or U30259 (N_30259,N_28017,N_29704);
xor U30260 (N_30260,N_27726,N_25534);
or U30261 (N_30261,N_29499,N_28412);
or U30262 (N_30262,N_26641,N_29125);
and U30263 (N_30263,N_26547,N_25343);
nor U30264 (N_30264,N_27321,N_26636);
nor U30265 (N_30265,N_29485,N_26460);
and U30266 (N_30266,N_25649,N_27950);
or U30267 (N_30267,N_26037,N_29642);
and U30268 (N_30268,N_26334,N_28433);
xor U30269 (N_30269,N_28710,N_28359);
or U30270 (N_30270,N_27437,N_26098);
xnor U30271 (N_30271,N_27580,N_25810);
nand U30272 (N_30272,N_27504,N_29800);
nand U30273 (N_30273,N_26714,N_29322);
nor U30274 (N_30274,N_25929,N_26099);
and U30275 (N_30275,N_28670,N_29532);
and U30276 (N_30276,N_29787,N_29419);
or U30277 (N_30277,N_28228,N_28326);
or U30278 (N_30278,N_25228,N_28528);
and U30279 (N_30279,N_28479,N_27180);
and U30280 (N_30280,N_26415,N_28913);
xnor U30281 (N_30281,N_25084,N_29525);
nor U30282 (N_30282,N_28552,N_27122);
nor U30283 (N_30283,N_25925,N_29381);
nand U30284 (N_30284,N_27375,N_27753);
xor U30285 (N_30285,N_25281,N_28988);
nor U30286 (N_30286,N_26331,N_25363);
or U30287 (N_30287,N_28874,N_26767);
or U30288 (N_30288,N_26235,N_28620);
nand U30289 (N_30289,N_26780,N_29312);
or U30290 (N_30290,N_29124,N_28596);
nor U30291 (N_30291,N_27277,N_26683);
or U30292 (N_30292,N_28854,N_28174);
or U30293 (N_30293,N_26228,N_25976);
xnor U30294 (N_30294,N_27228,N_25133);
or U30295 (N_30295,N_27877,N_25465);
and U30296 (N_30296,N_27416,N_26340);
xnor U30297 (N_30297,N_29831,N_26926);
nor U30298 (N_30298,N_26017,N_26198);
xnor U30299 (N_30299,N_25559,N_28811);
or U30300 (N_30300,N_29794,N_29937);
or U30301 (N_30301,N_27101,N_27313);
nor U30302 (N_30302,N_28134,N_29822);
xnor U30303 (N_30303,N_28202,N_25067);
nor U30304 (N_30304,N_25950,N_25866);
and U30305 (N_30305,N_26940,N_29051);
xnor U30306 (N_30306,N_27756,N_29321);
xnor U30307 (N_30307,N_28436,N_29194);
and U30308 (N_30308,N_25278,N_29346);
nor U30309 (N_30309,N_25970,N_28751);
or U30310 (N_30310,N_25361,N_29074);
xnor U30311 (N_30311,N_26674,N_27855);
xnor U30312 (N_30312,N_29206,N_28363);
xor U30313 (N_30313,N_25058,N_27609);
xor U30314 (N_30314,N_26736,N_25853);
nor U30315 (N_30315,N_27727,N_25910);
nor U30316 (N_30316,N_28377,N_25911);
and U30317 (N_30317,N_28844,N_29492);
nor U30318 (N_30318,N_29638,N_26085);
nor U30319 (N_30319,N_26159,N_29520);
or U30320 (N_30320,N_27641,N_28585);
xnor U30321 (N_30321,N_27925,N_26933);
or U30322 (N_30322,N_28496,N_27964);
xor U30323 (N_30323,N_27824,N_25938);
nand U30324 (N_30324,N_25746,N_26680);
nor U30325 (N_30325,N_25889,N_28269);
nand U30326 (N_30326,N_27892,N_25651);
nor U30327 (N_30327,N_26798,N_26312);
or U30328 (N_30328,N_27643,N_29636);
nor U30329 (N_30329,N_28763,N_26893);
xnor U30330 (N_30330,N_26946,N_26425);
xor U30331 (N_30331,N_27656,N_29057);
or U30332 (N_30332,N_25501,N_28275);
or U30333 (N_30333,N_27361,N_29298);
xor U30334 (N_30334,N_29145,N_27105);
xnor U30335 (N_30335,N_27595,N_28162);
and U30336 (N_30336,N_26496,N_27909);
nand U30337 (N_30337,N_28801,N_28420);
nand U30338 (N_30338,N_29482,N_29913);
nor U30339 (N_30339,N_27730,N_28995);
xor U30340 (N_30340,N_28047,N_27667);
nor U30341 (N_30341,N_25899,N_25967);
or U30342 (N_30342,N_27788,N_26807);
and U30343 (N_30343,N_25118,N_29143);
nand U30344 (N_30344,N_28268,N_26071);
and U30345 (N_30345,N_25731,N_26869);
nor U30346 (N_30346,N_27207,N_26886);
nand U30347 (N_30347,N_29142,N_27132);
or U30348 (N_30348,N_27376,N_28400);
or U30349 (N_30349,N_26706,N_27535);
and U30350 (N_30350,N_26923,N_25982);
nand U30351 (N_30351,N_27503,N_26395);
or U30352 (N_30352,N_25433,N_27281);
and U30353 (N_30353,N_26704,N_28419);
nor U30354 (N_30354,N_28695,N_26201);
nand U30355 (N_30355,N_25261,N_28058);
nor U30356 (N_30356,N_27847,N_27090);
nor U30357 (N_30357,N_29628,N_26506);
or U30358 (N_30358,N_29369,N_29020);
nor U30359 (N_30359,N_27343,N_25165);
nand U30360 (N_30360,N_25192,N_28050);
nor U30361 (N_30361,N_25521,N_29221);
or U30362 (N_30362,N_28028,N_26556);
and U30363 (N_30363,N_26212,N_29554);
and U30364 (N_30364,N_25896,N_27394);
or U30365 (N_30365,N_28474,N_26377);
nor U30366 (N_30366,N_26669,N_29140);
nand U30367 (N_30367,N_27462,N_25364);
and U30368 (N_30368,N_26422,N_29629);
nand U30369 (N_30369,N_26824,N_26260);
xnor U30370 (N_30370,N_28401,N_29848);
or U30371 (N_30371,N_27931,N_27470);
and U30372 (N_30372,N_26021,N_29404);
nor U30373 (N_30373,N_27459,N_27069);
and U30374 (N_30374,N_29052,N_26183);
and U30375 (N_30375,N_25216,N_26066);
or U30376 (N_30376,N_28473,N_28715);
nand U30377 (N_30377,N_27669,N_25830);
and U30378 (N_30378,N_25700,N_27665);
or U30379 (N_30379,N_27408,N_28285);
xor U30380 (N_30380,N_26549,N_25702);
nand U30381 (N_30381,N_27691,N_26000);
nor U30382 (N_30382,N_28218,N_25485);
nor U30383 (N_30383,N_29799,N_27679);
xnor U30384 (N_30384,N_26289,N_25495);
nand U30385 (N_30385,N_26818,N_29616);
and U30386 (N_30386,N_25372,N_29083);
or U30387 (N_30387,N_27401,N_29875);
or U30388 (N_30388,N_26874,N_29313);
or U30389 (N_30389,N_27620,N_27508);
and U30390 (N_30390,N_25340,N_25301);
nor U30391 (N_30391,N_29873,N_28538);
nor U30392 (N_30392,N_25140,N_29862);
and U30393 (N_30393,N_27164,N_27117);
and U30394 (N_30394,N_27237,N_29640);
nand U30395 (N_30395,N_25270,N_29511);
and U30396 (N_30396,N_28399,N_27256);
xor U30397 (N_30397,N_26803,N_26120);
xor U30398 (N_30398,N_27760,N_26026);
or U30399 (N_30399,N_27553,N_26450);
nand U30400 (N_30400,N_27252,N_25052);
or U30401 (N_30401,N_25125,N_29250);
nand U30402 (N_30402,N_27110,N_28151);
nor U30403 (N_30403,N_28522,N_29156);
nand U30404 (N_30404,N_29227,N_28212);
xnor U30405 (N_30405,N_29667,N_27196);
or U30406 (N_30406,N_27668,N_26483);
or U30407 (N_30407,N_29089,N_27739);
and U30408 (N_30408,N_25577,N_26288);
xor U30409 (N_30409,N_27919,N_27269);
or U30410 (N_30410,N_29441,N_26112);
or U30411 (N_30411,N_26924,N_28276);
nand U30412 (N_30412,N_26581,N_26226);
xor U30413 (N_30413,N_25130,N_26330);
xnor U30414 (N_30414,N_26954,N_29497);
nand U30415 (N_30415,N_28441,N_28816);
and U30416 (N_30416,N_28618,N_27428);
nor U30417 (N_30417,N_25457,N_27373);
nor U30418 (N_30418,N_28572,N_25690);
nor U30419 (N_30419,N_29048,N_27949);
or U30420 (N_30420,N_29560,N_28026);
nand U30421 (N_30421,N_29285,N_26567);
xor U30422 (N_30422,N_28061,N_27542);
and U30423 (N_30423,N_26478,N_29754);
xor U30424 (N_30424,N_27692,N_26388);
or U30425 (N_30425,N_28426,N_26995);
or U30426 (N_30426,N_26870,N_26859);
or U30427 (N_30427,N_27568,N_28372);
nor U30428 (N_30428,N_26336,N_26106);
xor U30429 (N_30429,N_29084,N_25722);
nand U30430 (N_30430,N_27005,N_28700);
xor U30431 (N_30431,N_27440,N_29682);
nor U30432 (N_30432,N_25979,N_27050);
and U30433 (N_30433,N_27091,N_27075);
or U30434 (N_30434,N_27625,N_29484);
or U30435 (N_30435,N_28983,N_27029);
or U30436 (N_30436,N_26861,N_27732);
xor U30437 (N_30437,N_25455,N_29879);
nand U30438 (N_30438,N_27275,N_26487);
or U30439 (N_30439,N_25112,N_28547);
xor U30440 (N_30440,N_26854,N_26215);
nor U30441 (N_30441,N_27034,N_25920);
nor U30442 (N_30442,N_26782,N_26417);
xnor U30443 (N_30443,N_29097,N_28834);
or U30444 (N_30444,N_29589,N_26494);
xor U30445 (N_30445,N_25775,N_26243);
xnor U30446 (N_30446,N_27642,N_27743);
nand U30447 (N_30447,N_29559,N_26871);
or U30448 (N_30448,N_28052,N_29921);
xnor U30449 (N_30449,N_27396,N_28772);
xnor U30450 (N_30450,N_28098,N_27201);
nand U30451 (N_30451,N_29350,N_28110);
xnor U30452 (N_30452,N_25520,N_25342);
or U30453 (N_30453,N_26927,N_25116);
or U30454 (N_30454,N_26116,N_26405);
nand U30455 (N_30455,N_26653,N_28245);
nor U30456 (N_30456,N_25439,N_29098);
nand U30457 (N_30457,N_27162,N_25034);
and U30458 (N_30458,N_26967,N_27188);
xnor U30459 (N_30459,N_26578,N_29371);
and U30460 (N_30460,N_25619,N_29155);
xor U30461 (N_30461,N_26648,N_28843);
xnor U30462 (N_30462,N_29551,N_28402);
xnor U30463 (N_30463,N_29694,N_26781);
nor U30464 (N_30464,N_27823,N_28367);
and U30465 (N_30465,N_29306,N_25669);
or U30466 (N_30466,N_25932,N_27064);
nand U30467 (N_30467,N_27413,N_29780);
xnor U30468 (N_30468,N_28430,N_28252);
nor U30469 (N_30469,N_25043,N_29195);
xor U30470 (N_30470,N_27000,N_27340);
or U30471 (N_30471,N_28297,N_29232);
nand U30472 (N_30472,N_25373,N_29027);
or U30473 (N_30473,N_28232,N_29515);
and U30474 (N_30474,N_25529,N_29608);
nand U30475 (N_30475,N_29615,N_29683);
and U30476 (N_30476,N_28502,N_25632);
xor U30477 (N_30477,N_27358,N_28503);
xnor U30478 (N_30478,N_27472,N_26844);
or U30479 (N_30479,N_26348,N_27487);
and U30480 (N_30480,N_29326,N_25110);
and U30481 (N_30481,N_27996,N_25657);
nand U30482 (N_30482,N_25119,N_29953);
nand U30483 (N_30483,N_26253,N_25263);
and U30484 (N_30484,N_29386,N_25254);
nor U30485 (N_30485,N_28658,N_26701);
or U30486 (N_30486,N_28160,N_27992);
nand U30487 (N_30487,N_29144,N_27866);
nor U30488 (N_30488,N_28553,N_28066);
nor U30489 (N_30489,N_28594,N_29957);
nand U30490 (N_30490,N_26117,N_29336);
nor U30491 (N_30491,N_27115,N_27498);
or U30492 (N_30492,N_29411,N_27764);
nor U30493 (N_30493,N_25243,N_29113);
or U30494 (N_30494,N_29550,N_25264);
xnor U30495 (N_30495,N_27537,N_26374);
xnor U30496 (N_30496,N_28645,N_28859);
nand U30497 (N_30497,N_25764,N_26274);
and U30498 (N_30498,N_27516,N_25567);
xor U30499 (N_30499,N_26843,N_27079);
and U30500 (N_30500,N_25381,N_26188);
nand U30501 (N_30501,N_25902,N_26928);
and U30502 (N_30502,N_26901,N_27589);
and U30503 (N_30503,N_27818,N_29561);
and U30504 (N_30504,N_29941,N_25576);
nand U30505 (N_30505,N_26621,N_25241);
nand U30506 (N_30506,N_29149,N_26564);
and U30507 (N_30507,N_29672,N_28025);
or U30508 (N_30508,N_28595,N_28787);
xnor U30509 (N_30509,N_27930,N_29824);
and U30510 (N_30510,N_28475,N_26719);
nand U30511 (N_30511,N_29979,N_29367);
xnor U30512 (N_30512,N_25865,N_26703);
or U30513 (N_30513,N_26794,N_25205);
or U30514 (N_30514,N_28023,N_29058);
or U30515 (N_30515,N_26449,N_28177);
nand U30516 (N_30516,N_25668,N_28320);
nand U30517 (N_30517,N_29586,N_28599);
nor U30518 (N_30518,N_28705,N_29169);
xnor U30519 (N_30519,N_29977,N_29798);
or U30520 (N_30520,N_28004,N_25175);
and U30521 (N_30521,N_27037,N_28685);
and U30522 (N_30522,N_28413,N_29131);
and U30523 (N_30523,N_25122,N_28878);
or U30524 (N_30524,N_28515,N_28814);
nand U30525 (N_30525,N_27558,N_26702);
xor U30526 (N_30526,N_29157,N_26268);
nor U30527 (N_30527,N_26054,N_27002);
nand U30528 (N_30528,N_28891,N_25763);
nor U30529 (N_30529,N_25411,N_26064);
and U30530 (N_30530,N_27555,N_28225);
nor U30531 (N_30531,N_26984,N_27584);
xor U30532 (N_30532,N_25442,N_25699);
nor U30533 (N_30533,N_25931,N_29400);
and U30534 (N_30534,N_28975,N_25120);
nor U30535 (N_30535,N_29374,N_29078);
and U30536 (N_30536,N_26231,N_28924);
nor U30537 (N_30537,N_29700,N_29340);
nor U30538 (N_30538,N_27712,N_29993);
or U30539 (N_30539,N_26975,N_29292);
or U30540 (N_30540,N_25818,N_27322);
nand U30541 (N_30541,N_29293,N_27402);
xor U30542 (N_30542,N_27485,N_27678);
and U30543 (N_30543,N_28623,N_28575);
or U30544 (N_30544,N_28082,N_27009);
nor U30545 (N_30545,N_29687,N_26062);
or U30546 (N_30546,N_26888,N_25100);
and U30547 (N_30547,N_29461,N_29833);
nand U30548 (N_30548,N_26451,N_28365);
or U30549 (N_30549,N_28264,N_29388);
nor U30550 (N_30550,N_29578,N_28346);
or U30551 (N_30551,N_27368,N_26891);
xnor U30552 (N_30552,N_27897,N_25869);
or U30553 (N_30553,N_25060,N_25835);
xnor U30554 (N_30554,N_25494,N_26809);
nand U30555 (N_30555,N_29670,N_27385);
nand U30556 (N_30556,N_28385,N_25924);
or U30557 (N_30557,N_27438,N_25900);
and U30558 (N_30558,N_28929,N_27779);
nand U30559 (N_30559,N_27249,N_27246);
nor U30560 (N_30560,N_28549,N_27325);
nor U30561 (N_30561,N_25180,N_25939);
or U30562 (N_30562,N_25903,N_25694);
and U30563 (N_30563,N_25952,N_26887);
and U30564 (N_30564,N_29231,N_26213);
nand U30565 (N_30565,N_28488,N_27100);
xnor U30566 (N_30566,N_29067,N_25326);
nor U30567 (N_30567,N_26293,N_29934);
or U30568 (N_30568,N_27626,N_25603);
and U30569 (N_30569,N_26810,N_28578);
nand U30570 (N_30570,N_25565,N_27077);
and U30571 (N_30571,N_28369,N_26980);
nor U30572 (N_30572,N_29444,N_26637);
xnor U30573 (N_30573,N_25291,N_25015);
xnor U30574 (N_30574,N_26276,N_27452);
and U30575 (N_30575,N_27415,N_28652);
xnor U30576 (N_30576,N_28261,N_25637);
or U30577 (N_30577,N_25695,N_29455);
and U30578 (N_30578,N_25605,N_26392);
nor U30579 (N_30579,N_27466,N_29076);
nand U30580 (N_30580,N_29107,N_28088);
nor U30581 (N_30581,N_28880,N_26203);
xnor U30582 (N_30582,N_27849,N_25020);
nor U30583 (N_30583,N_27200,N_26295);
nor U30584 (N_30584,N_27884,N_26486);
nor U30585 (N_30585,N_29165,N_29432);
nand U30586 (N_30586,N_29773,N_28898);
nand U30587 (N_30587,N_27020,N_26936);
nand U30588 (N_30588,N_25280,N_26971);
nand U30589 (N_30589,N_26088,N_27819);
and U30590 (N_30590,N_25473,N_26402);
xnor U30591 (N_30591,N_28836,N_27710);
or U30592 (N_30592,N_29855,N_29967);
xnor U30593 (N_30593,N_28725,N_29917);
xnor U30594 (N_30594,N_27016,N_26059);
or U30595 (N_30595,N_28714,N_29591);
nand U30596 (N_30596,N_27015,N_28906);
xnor U30597 (N_30597,N_27011,N_27857);
nor U30598 (N_30598,N_25204,N_27941);
xnor U30599 (N_30599,N_28062,N_26760);
or U30600 (N_30600,N_29239,N_25890);
and U30601 (N_30601,N_26317,N_26056);
or U30602 (N_30602,N_26663,N_26616);
and U30603 (N_30603,N_26762,N_27551);
xnor U30604 (N_30604,N_28166,N_28970);
and U30605 (N_30605,N_27586,N_27421);
and U30606 (N_30606,N_27123,N_26858);
or U30607 (N_30607,N_25025,N_27251);
or U30608 (N_30608,N_25393,N_27374);
nand U30609 (N_30609,N_25708,N_28462);
nor U30610 (N_30610,N_25837,N_25492);
nand U30611 (N_30611,N_26829,N_25648);
xnor U30612 (N_30612,N_27515,N_27046);
nor U30613 (N_30613,N_26287,N_28262);
nand U30614 (N_30614,N_25901,N_25832);
xor U30615 (N_30615,N_28895,N_25143);
and U30616 (N_30616,N_26877,N_25538);
or U30617 (N_30617,N_28655,N_27209);
and U30618 (N_30618,N_27799,N_25554);
nand U30619 (N_30619,N_28295,N_25171);
nand U30620 (N_30620,N_28096,N_25895);
nor U30621 (N_30621,N_27088,N_26303);
xnor U30622 (N_30622,N_29618,N_28500);
or U30623 (N_30623,N_26294,N_27419);
and U30624 (N_30624,N_25436,N_28856);
and U30625 (N_30625,N_25660,N_28072);
and U30626 (N_30626,N_29673,N_26633);
and U30627 (N_30627,N_27587,N_26004);
or U30628 (N_30628,N_25949,N_29201);
or U30629 (N_30629,N_29579,N_25621);
nor U30630 (N_30630,N_26477,N_28451);
or U30631 (N_30631,N_25582,N_29111);
or U30632 (N_30632,N_26991,N_27882);
nand U30633 (N_30633,N_27226,N_27733);
nand U30634 (N_30634,N_26597,N_26675);
and U30635 (N_30635,N_26508,N_29723);
and U30636 (N_30636,N_26756,N_27724);
nand U30637 (N_30637,N_26127,N_25139);
xnor U30638 (N_30638,N_26593,N_28195);
nor U30639 (N_30639,N_25445,N_26434);
nor U30640 (N_30640,N_29054,N_28292);
nor U30641 (N_30641,N_25456,N_29796);
or U30642 (N_30642,N_27554,N_27471);
xor U30643 (N_30643,N_28069,N_28366);
nand U30644 (N_30644,N_29759,N_26712);
or U30645 (N_30645,N_26727,N_29849);
nand U30646 (N_30646,N_29207,N_25131);
xnor U30647 (N_30647,N_27006,N_27356);
or U30648 (N_30648,N_28689,N_26952);
and U30649 (N_30649,N_26515,N_27280);
nor U30650 (N_30650,N_26920,N_26979);
and U30651 (N_30651,N_25461,N_28724);
nor U30652 (N_30652,N_28223,N_28135);
xor U30653 (N_30653,N_28481,N_27121);
nor U30654 (N_30654,N_25815,N_25467);
nand U30655 (N_30655,N_29254,N_26423);
xor U30656 (N_30656,N_26599,N_25793);
nand U30657 (N_30657,N_28394,N_25022);
nor U30658 (N_30658,N_27731,N_25675);
nor U30659 (N_30659,N_27190,N_27605);
nand U30660 (N_30660,N_27221,N_28318);
and U30661 (N_30661,N_25258,N_27684);
and U30662 (N_30662,N_29746,N_28560);
and U30663 (N_30663,N_29697,N_28512);
xor U30664 (N_30664,N_28669,N_29433);
or U30665 (N_30665,N_26257,N_27972);
nand U30666 (N_30666,N_25985,N_27255);
xnor U30667 (N_30667,N_27570,N_26177);
nand U30668 (N_30668,N_29770,N_27932);
or U30669 (N_30669,N_28642,N_28121);
xor U30670 (N_30670,N_27946,N_27053);
xnor U30671 (N_30671,N_26729,N_27397);
nand U30672 (N_30672,N_28704,N_25044);
or U30673 (N_30673,N_29662,N_25849);
xnor U30674 (N_30674,N_25218,N_28603);
nor U30675 (N_30675,N_26443,N_26505);
or U30676 (N_30676,N_29428,N_28581);
xor U30677 (N_30677,N_25403,N_25102);
and U30678 (N_30678,N_28145,N_27746);
or U30679 (N_30679,N_26453,N_26694);
or U30680 (N_30680,N_26692,N_28742);
nor U30681 (N_30681,N_28953,N_28463);
or U30682 (N_30682,N_27740,N_26668);
nor U30683 (N_30683,N_27295,N_25018);
or U30684 (N_30684,N_28130,N_26628);
nor U30685 (N_30685,N_26677,N_25188);
nor U30686 (N_30686,N_29013,N_25993);
nor U30687 (N_30687,N_28472,N_29032);
xnor U30688 (N_30688,N_27552,N_27456);
xor U30689 (N_30689,N_25366,N_26529);
or U30690 (N_30690,N_25592,N_26391);
xor U30691 (N_30691,N_27337,N_27645);
nor U30692 (N_30692,N_25916,N_27359);
and U30693 (N_30693,N_25024,N_28119);
nor U30694 (N_30694,N_27126,N_27955);
or U30695 (N_30695,N_26531,N_28222);
or U30696 (N_30696,N_28404,N_26455);
nor U30697 (N_30697,N_28137,N_27181);
or U30698 (N_30698,N_27870,N_28409);
or U30699 (N_30699,N_27194,N_26291);
or U30700 (N_30700,N_26216,N_26918);
nor U30701 (N_30701,N_26830,N_25946);
xor U30702 (N_30702,N_28739,N_27795);
nand U30703 (N_30703,N_26619,N_25771);
xor U30704 (N_30704,N_28306,N_28272);
nand U30705 (N_30705,N_29614,N_25293);
nor U30706 (N_30706,N_29126,N_28776);
nand U30707 (N_30707,N_26618,N_25097);
xor U30708 (N_30708,N_25666,N_27003);
and U30709 (N_30709,N_29997,N_26292);
nand U30710 (N_30710,N_25803,N_27927);
xnor U30711 (N_30711,N_28390,N_27247);
nand U30712 (N_30712,N_29300,N_26446);
nor U30713 (N_30713,N_26551,N_29264);
xnor U30714 (N_30714,N_27817,N_26247);
nand U30715 (N_30715,N_28154,N_29650);
nor U30716 (N_30716,N_26376,N_28764);
xor U30717 (N_30717,N_25858,N_29114);
or U30718 (N_30718,N_26430,N_29693);
xor U30719 (N_30719,N_26896,N_28798);
or U30720 (N_30720,N_27474,N_27619);
xor U30721 (N_30721,N_28910,N_26604);
and U30722 (N_30722,N_25283,N_25251);
or U30723 (N_30723,N_28055,N_27030);
xnor U30724 (N_30724,N_25796,N_25141);
and U30725 (N_30725,N_25295,N_28974);
nor U30726 (N_30726,N_27518,N_28612);
nand U30727 (N_30727,N_27311,N_27709);
nand U30728 (N_30728,N_29516,N_25714);
nand U30729 (N_30729,N_26214,N_27894);
nand U30730 (N_30730,N_28782,N_27478);
xor U30731 (N_30731,N_29413,N_27007);
nor U30732 (N_30732,N_26421,N_26302);
and U30733 (N_30733,N_29584,N_29838);
nand U30734 (N_30734,N_27986,N_29376);
or U30735 (N_30735,N_26755,N_25149);
and U30736 (N_30736,N_26246,N_25490);
and U30737 (N_30737,N_25158,N_29804);
nor U30738 (N_30738,N_28767,N_26850);
nand U30739 (N_30739,N_29783,N_29172);
or U30740 (N_30740,N_25596,N_25402);
xor U30741 (N_30741,N_29880,N_25750);
xnor U30742 (N_30742,N_25684,N_26501);
or U30743 (N_30743,N_27059,N_27912);
nor U30744 (N_30744,N_26350,N_25031);
nand U30745 (N_30745,N_27435,N_27107);
nor U30746 (N_30746,N_27152,N_27670);
xor U30747 (N_30747,N_25341,N_29033);
and U30748 (N_30748,N_25332,N_26823);
or U30749 (N_30749,N_26732,N_26038);
nor U30750 (N_30750,N_26759,N_29716);
nand U30751 (N_30751,N_29427,N_29276);
and U30752 (N_30752,N_26559,N_25498);
or U30753 (N_30753,N_25820,N_25479);
nor U30754 (N_30754,N_28283,N_27157);
nor U30755 (N_30755,N_28187,N_27481);
and U30756 (N_30756,N_25502,N_28471);
nor U30757 (N_30757,N_27039,N_27323);
xnor U30758 (N_30758,N_28358,N_29106);
nand U30759 (N_30759,N_26074,N_29731);
xnor U30760 (N_30760,N_28887,N_26457);
and U30761 (N_30761,N_28498,N_25047);
nor U30762 (N_30762,N_29183,N_25049);
xor U30763 (N_30763,N_26649,N_27550);
xnor U30764 (N_30764,N_28976,N_27082);
and U30765 (N_30765,N_29664,N_25358);
xor U30766 (N_30766,N_27213,N_29205);
and U30767 (N_30767,N_28935,N_27838);
or U30768 (N_30768,N_26063,N_27720);
or U30769 (N_30769,N_29705,N_25151);
nor U30770 (N_30770,N_25590,N_25634);
nand U30771 (N_30771,N_29310,N_29029);
nor U30772 (N_30772,N_29181,N_28155);
xor U30773 (N_30773,N_27736,N_26086);
or U30774 (N_30774,N_26899,N_27342);
xor U30775 (N_30775,N_28514,N_27657);
xor U30776 (N_30776,N_27494,N_25313);
or U30777 (N_30777,N_27549,N_29856);
and U30778 (N_30778,N_29217,N_27898);
or U30779 (N_30779,N_29070,N_28735);
nand U30780 (N_30780,N_26640,N_27043);
nor U30781 (N_30781,N_25989,N_26366);
nand U30782 (N_30782,N_28830,N_27652);
nor U30783 (N_30783,N_29304,N_29050);
nor U30784 (N_30784,N_25999,N_26406);
nor U30785 (N_30785,N_29069,N_29085);
and U30786 (N_30786,N_29789,N_27261);
or U30787 (N_30787,N_25256,N_29595);
nand U30788 (N_30788,N_27879,N_25200);
nand U30789 (N_30789,N_27074,N_28698);
nand U30790 (N_30790,N_27761,N_25365);
nand U30791 (N_30791,N_28532,N_26825);
nor U30792 (N_30792,N_25923,N_25222);
or U30793 (N_30793,N_28138,N_29778);
xor U30794 (N_30794,N_28270,N_27800);
nor U30795 (N_30795,N_29337,N_25476);
nor U30796 (N_30796,N_27203,N_29902);
nand U30797 (N_30797,N_29825,N_27216);
nor U30798 (N_30798,N_29980,N_28007);
nand U30799 (N_30799,N_28510,N_29502);
nor U30800 (N_30800,N_28075,N_29179);
nor U30801 (N_30801,N_28312,N_25400);
nor U30802 (N_30802,N_29582,N_29747);
and U30803 (N_30803,N_25981,N_27718);
nor U30804 (N_30804,N_29991,N_26978);
or U30805 (N_30805,N_26084,N_25017);
xnor U30806 (N_30806,N_28005,N_28435);
nand U30807 (N_30807,N_25080,N_27728);
and U30808 (N_30808,N_28982,N_26452);
xor U30809 (N_30809,N_27786,N_27463);
xnor U30810 (N_30810,N_26594,N_29030);
nand U30811 (N_30811,N_29174,N_26557);
or U30812 (N_30812,N_26341,N_29066);
or U30813 (N_30813,N_29535,N_28826);
or U30814 (N_30814,N_26262,N_26134);
xor U30815 (N_30815,N_25555,N_25547);
nor U30816 (N_30816,N_27398,N_25333);
xnor U30817 (N_30817,N_26034,N_25825);
xor U30818 (N_30818,N_28468,N_29417);
and U30819 (N_30819,N_27148,N_29707);
or U30820 (N_30820,N_26454,N_27896);
nor U30821 (N_30821,N_25897,N_26309);
and U30822 (N_30822,N_28820,N_25551);
nand U30823 (N_30823,N_25432,N_29517);
or U30824 (N_30824,N_27137,N_26516);
xnor U30825 (N_30825,N_25829,N_27636);
nand U30826 (N_30826,N_25370,N_25886);
nand U30827 (N_30827,N_25645,N_26783);
nor U30828 (N_30828,N_29710,N_28453);
xor U30829 (N_30829,N_27853,N_29909);
xnor U30830 (N_30830,N_28476,N_27414);
or U30831 (N_30831,N_28686,N_25103);
xnor U30832 (N_30832,N_29549,N_27087);
or U30833 (N_30833,N_25536,N_25870);
and U30834 (N_30834,N_26414,N_28823);
or U30835 (N_30835,N_25497,N_28615);
nor U30836 (N_30836,N_28955,N_26768);
nor U30837 (N_30837,N_29307,N_27716);
xor U30838 (N_30838,N_28980,N_29200);
or U30839 (N_30839,N_27388,N_27763);
nand U30840 (N_30840,N_28657,N_27887);
nor U30841 (N_30841,N_28901,N_27135);
and U30842 (N_30842,N_28635,N_29191);
nand U30843 (N_30843,N_26480,N_26381);
xor U30844 (N_30844,N_28550,N_28758);
nor U30845 (N_30845,N_28238,N_27242);
or U30846 (N_30846,N_27693,N_28165);
xor U30847 (N_30847,N_27328,N_28964);
nor U30848 (N_30848,N_25459,N_29692);
or U30849 (N_30849,N_29922,N_25063);
xnor U30850 (N_30850,N_28752,N_25795);
and U30851 (N_30851,N_26242,N_25821);
and U30852 (N_30852,N_28180,N_26013);
nor U30853 (N_30853,N_27512,N_28095);
nand U30854 (N_30854,N_26290,N_27686);
nand U30855 (N_30855,N_29898,N_28477);
and U30856 (N_30856,N_29829,N_27747);
and U30857 (N_30857,N_25132,N_29575);
nor U30858 (N_30858,N_25438,N_26343);
and U30859 (N_30859,N_25503,N_25670);
xnor U30860 (N_30860,N_28508,N_25040);
and U30861 (N_30861,N_27395,N_26407);
and U30862 (N_30862,N_26573,N_25549);
or U30863 (N_30863,N_26642,N_25138);
xor U30864 (N_30864,N_29574,N_27338);
or U30865 (N_30865,N_29213,N_29924);
xor U30866 (N_30866,N_28604,N_27715);
nor U30867 (N_30867,N_28083,N_27507);
or U30868 (N_30868,N_29809,N_25723);
xor U30869 (N_30869,N_27199,N_28644);
and U30870 (N_30870,N_25686,N_29580);
and U30871 (N_30871,N_27968,N_29806);
nor U30872 (N_30872,N_26046,N_27310);
or U30873 (N_30873,N_26681,N_29319);
nand U30874 (N_30874,N_29378,N_27314);
nor U30875 (N_30875,N_28022,N_29382);
nand U30876 (N_30876,N_29699,N_27890);
nor U30877 (N_30877,N_27169,N_28115);
or U30878 (N_30878,N_27975,N_25360);
or U30879 (N_30879,N_29305,N_27409);
nand U30880 (N_30880,N_26224,N_26277);
xor U30881 (N_30881,N_27521,N_28215);
nor U30882 (N_30882,N_27995,N_28517);
xor U30883 (N_30883,N_26442,N_28230);
nand U30884 (N_30884,N_27780,N_28125);
or U30885 (N_30885,N_28789,N_29514);
and U30886 (N_30886,N_26587,N_26646);
nand U30887 (N_30887,N_26707,N_25059);
and U30888 (N_30888,N_28324,N_29904);
nor U30889 (N_30889,N_27172,N_27168);
and U30890 (N_30890,N_25936,N_25153);
nor U30891 (N_30891,N_27274,N_26266);
xnor U30892 (N_30892,N_25734,N_28884);
nor U30893 (N_30893,N_29563,N_25836);
nor U30894 (N_30894,N_26543,N_28233);
nor U30895 (N_30895,N_25077,N_29585);
or U30896 (N_30896,N_27316,N_25481);
xor U30897 (N_30897,N_28467,N_27202);
or U30898 (N_30898,N_27973,N_26300);
xor U30899 (N_30899,N_29632,N_27465);
and U30900 (N_30900,N_29741,N_25591);
or U30901 (N_30901,N_28265,N_25328);
or U30902 (N_30902,N_26327,N_26223);
or U30903 (N_30903,N_27532,N_26148);
or U30904 (N_30904,N_27791,N_29814);
nor U30905 (N_30905,N_28922,N_28396);
or U30906 (N_30906,N_27351,N_25085);
or U30907 (N_30907,N_28041,N_27806);
or U30908 (N_30908,N_28986,N_27287);
nand U30909 (N_30909,N_26281,N_25334);
or U30910 (N_30910,N_29620,N_26499);
nor U30911 (N_30911,N_27035,N_25862);
nand U30912 (N_30912,N_27723,N_25541);
xor U30913 (N_30913,N_25081,N_28785);
and U30914 (N_30914,N_28956,N_29861);
or U30915 (N_30915,N_29858,N_29761);
nor U30916 (N_30916,N_29465,N_25867);
nor U30917 (N_30917,N_26128,N_26225);
nand U30918 (N_30918,N_29422,N_28065);
nor U30919 (N_30919,N_26069,N_27993);
xnor U30920 (N_30920,N_26542,N_28876);
nor U30921 (N_30921,N_27575,N_26774);
or U30922 (N_30922,N_28384,N_28565);
or U30923 (N_30923,N_26318,N_28337);
and U30924 (N_30924,N_29137,N_25537);
or U30925 (N_30925,N_25926,N_29262);
nand U30926 (N_30926,N_27592,N_27051);
nand U30927 (N_30927,N_28011,N_28093);
nand U30928 (N_30928,N_27054,N_29403);
nand U30929 (N_30929,N_28168,N_26191);
xnor U30930 (N_30930,N_27412,N_25874);
nor U30931 (N_30931,N_26286,N_27630);
nor U30932 (N_30932,N_29109,N_25681);
or U30933 (N_30933,N_29981,N_26082);
and U30934 (N_30934,N_26524,N_27382);
and U30935 (N_30935,N_28726,N_29540);
and U30936 (N_30936,N_29416,N_25610);
nor U30937 (N_30937,N_26672,N_26320);
and U30938 (N_30938,N_25389,N_25159);
and U30939 (N_30939,N_27565,N_25808);
or U30940 (N_30940,N_29966,N_25799);
xor U30941 (N_30941,N_27070,N_26070);
and U30942 (N_30942,N_25562,N_25868);
and U30943 (N_30943,N_28478,N_25491);
nand U30944 (N_30944,N_28667,N_25876);
and U30945 (N_30945,N_27205,N_28322);
or U30946 (N_30946,N_29352,N_28544);
or U30947 (N_30947,N_27618,N_29479);
xnor U30948 (N_30948,N_25428,N_27197);
or U30949 (N_30949,N_28893,N_29588);
and U30950 (N_30950,N_27405,N_27469);
nor U30951 (N_30951,N_28484,N_29817);
or U30952 (N_30952,N_25941,N_27856);
nand U30953 (N_30953,N_27563,N_26563);
xnor U30954 (N_30954,N_29963,N_28696);
or U30955 (N_30955,N_27638,N_28605);
or U30956 (N_30956,N_29587,N_28266);
nor U30957 (N_30957,N_28981,N_27057);
xor U30958 (N_30958,N_26245,N_28060);
xor U30959 (N_30959,N_28450,N_25226);
or U30960 (N_30960,N_26721,N_28221);
and U30961 (N_30961,N_27966,N_29721);
and U30962 (N_30962,N_26171,N_27782);
and U30963 (N_30963,N_29764,N_29448);
or U30964 (N_30964,N_26109,N_26411);
and U30965 (N_30965,N_29603,N_29860);
or U30966 (N_30966,N_26155,N_29583);
or U30967 (N_30967,N_26527,N_28203);
xnor U30968 (N_30968,N_28448,N_28106);
and U30969 (N_30969,N_28659,N_28941);
nor U30970 (N_30970,N_25781,N_25323);
and U30971 (N_30971,N_28625,N_28716);
nor U30972 (N_30972,N_26831,N_28647);
and U30973 (N_30973,N_25493,N_27591);
and U30974 (N_30974,N_28352,N_27517);
and U30975 (N_30975,N_25161,N_26699);
or U30976 (N_30976,N_26306,N_29989);
xnor U30977 (N_30977,N_28756,N_25398);
xnor U30978 (N_30978,N_27350,N_26605);
xnor U30979 (N_30979,N_25462,N_28087);
or U30980 (N_30980,N_26550,N_25996);
or U30981 (N_30981,N_27093,N_26202);
xor U30982 (N_30982,N_28079,N_25545);
nor U30983 (N_30983,N_27529,N_26817);
xnor U30984 (N_30984,N_26753,N_29274);
and U30985 (N_30985,N_28189,N_28835);
nand U30986 (N_30986,N_25737,N_25553);
or U30987 (N_30987,N_26833,N_27141);
or U30988 (N_30988,N_29148,N_29370);
or U30989 (N_30989,N_28818,N_26751);
nor U30990 (N_30990,N_25065,N_25894);
xor U30991 (N_30991,N_26473,N_29865);
and U30992 (N_30992,N_29494,N_26802);
nor U30993 (N_30993,N_26271,N_25797);
and U30994 (N_30994,N_25505,N_29970);
nand U30995 (N_30995,N_28178,N_28851);
and U30996 (N_30996,N_25933,N_28633);
xnor U30997 (N_30997,N_27562,N_28688);
nor U30998 (N_30998,N_26582,N_25838);
or U30999 (N_30999,N_25969,N_26010);
xor U31000 (N_31000,N_25072,N_29742);
nand U31001 (N_31001,N_29164,N_27253);
xnor U31002 (N_31002,N_28872,N_28912);
nor U31003 (N_31003,N_26456,N_26534);
and U31004 (N_31004,N_26372,N_25918);
and U31005 (N_31005,N_26645,N_25288);
nand U31006 (N_31006,N_27027,N_26947);
nand U31007 (N_31007,N_28579,N_29138);
or U31008 (N_31008,N_29299,N_28444);
xor U31009 (N_31009,N_27426,N_28792);
nand U31010 (N_31010,N_29189,N_25613);
nor U31011 (N_31011,N_29832,N_25447);
nand U31012 (N_31012,N_25658,N_28235);
or U31013 (N_31013,N_26269,N_26418);
or U31014 (N_31014,N_28971,N_26700);
nand U31015 (N_31015,N_29266,N_27915);
and U31016 (N_31016,N_28786,N_29135);
xnor U31017 (N_31017,N_26733,N_26044);
and U31018 (N_31018,N_27697,N_29807);
or U31019 (N_31019,N_28860,N_25013);
xnor U31020 (N_31020,N_26015,N_25284);
nor U31021 (N_31021,N_28574,N_26169);
nor U31022 (N_31022,N_29901,N_27793);
nor U31023 (N_31023,N_25273,N_26382);
nor U31024 (N_31024,N_25055,N_26726);
and U31025 (N_31025,N_25955,N_28628);
nand U31026 (N_31026,N_28832,N_29478);
nor U31027 (N_31027,N_29437,N_27944);
nand U31028 (N_31028,N_26027,N_25995);
and U31029 (N_31029,N_29625,N_26813);
or U31030 (N_31030,N_29275,N_27928);
nand U31031 (N_31031,N_28589,N_28888);
nor U31032 (N_31032,N_26765,N_28043);
or U31033 (N_31033,N_28584,N_28181);
nor U31034 (N_31034,N_27400,N_27564);
nor U31035 (N_31035,N_25157,N_27878);
xnor U31036 (N_31036,N_25189,N_25195);
nor U31037 (N_31037,N_29488,N_29512);
nand U31038 (N_31038,N_25905,N_25425);
or U31039 (N_31039,N_26848,N_26141);
or U31040 (N_31040,N_26012,N_25252);
or U31041 (N_31041,N_26590,N_29982);
and U31042 (N_31042,N_29351,N_25176);
nand U31043 (N_31043,N_28214,N_29987);
nand U31044 (N_31044,N_29363,N_25543);
and U31045 (N_31045,N_29593,N_29090);
nor U31046 (N_31046,N_27755,N_26301);
nor U31047 (N_31047,N_26519,N_26390);
nor U31048 (N_31048,N_29522,N_25512);
xnor U31049 (N_31049,N_28493,N_26772);
or U31050 (N_31050,N_29447,N_25227);
nand U31051 (N_31051,N_28209,N_25682);
and U31052 (N_31052,N_27648,N_26296);
or U31053 (N_31053,N_25399,N_27264);
xnor U31054 (N_31054,N_25000,N_26852);
and U31055 (N_31055,N_27947,N_27873);
nand U31056 (N_31056,N_28064,N_26790);
or U31057 (N_31057,N_27816,N_27784);
or U31058 (N_31058,N_27904,N_27384);
or U31059 (N_31059,N_25208,N_27293);
nand U31060 (N_31060,N_27130,N_26839);
and U31061 (N_31061,N_27839,N_29049);
xor U31062 (N_31062,N_29257,N_29839);
xnor U31063 (N_31063,N_28879,N_25388);
xnor U31064 (N_31064,N_27622,N_27033);
nor U31065 (N_31065,N_28703,N_25877);
nor U31066 (N_31066,N_26419,N_26591);
or U31067 (N_31067,N_25962,N_26747);
nor U31068 (N_31068,N_29592,N_26250);
or U31069 (N_31069,N_28734,N_25136);
nor U31070 (N_31070,N_28142,N_26526);
xor U31071 (N_31071,N_26077,N_25800);
nor U31072 (N_31072,N_27921,N_28442);
or U31073 (N_31073,N_29243,N_27309);
xor U31074 (N_31074,N_28662,N_28520);
nand U31075 (N_31075,N_26110,N_26598);
nor U31076 (N_31076,N_26763,N_25299);
or U31077 (N_31077,N_26170,N_28951);
nand U31078 (N_31078,N_29990,N_27425);
or U31079 (N_31079,N_27102,N_27086);
or U31080 (N_31080,N_29354,N_28486);
and U31081 (N_31081,N_28164,N_27372);
nand U31082 (N_31082,N_27010,N_26298);
and U31083 (N_31083,N_28849,N_25602);
xor U31084 (N_31084,N_27833,N_28799);
and U31085 (N_31085,N_29353,N_29343);
nand U31086 (N_31086,N_25267,N_28606);
nor U31087 (N_31087,N_28684,N_27773);
nand U31088 (N_31088,N_28925,N_26353);
or U31089 (N_31089,N_25987,N_28750);
or U31090 (N_31090,N_29785,N_26710);
or U31091 (N_31091,N_29954,N_29951);
nand U31092 (N_31092,N_25396,N_26622);
and U31093 (N_31093,N_25780,N_25676);
nor U31094 (N_31094,N_26693,N_26894);
nand U31095 (N_31095,N_27189,N_27796);
or U31096 (N_31096,N_26864,N_29680);
xnor U31097 (N_31097,N_28626,N_29442);
nor U31098 (N_31098,N_26822,N_29226);
and U31099 (N_31099,N_26773,N_25348);
nor U31100 (N_31100,N_25783,N_25525);
xor U31101 (N_31101,N_25579,N_26689);
nor U31102 (N_31102,N_29590,N_26081);
and U31103 (N_31103,N_28918,N_25948);
or U31104 (N_31104,N_28395,N_28499);
or U31105 (N_31105,N_26832,N_28624);
nor U31106 (N_31106,N_28205,N_26631);
and U31107 (N_31107,N_28894,N_29309);
nand U31108 (N_31108,N_28291,N_28349);
nor U31109 (N_31109,N_25856,N_25701);
nand U31110 (N_31110,N_25578,N_25071);
and U31111 (N_31111,N_26006,N_26471);
nand U31112 (N_31112,N_25231,N_26221);
nand U31113 (N_31113,N_25443,N_25826);
xor U31114 (N_31114,N_26094,N_26917);
or U31115 (N_31115,N_25721,N_25953);
nand U31116 (N_31116,N_28845,N_28561);
or U31117 (N_31117,N_27076,N_29562);
nand U31118 (N_31118,N_26718,N_29283);
or U31119 (N_31119,N_27676,N_29637);
nand U31120 (N_31120,N_25873,N_29871);
xor U31121 (N_31121,N_25471,N_28759);
nor U31122 (N_31122,N_27834,N_25094);
nor U31123 (N_31123,N_29470,N_25450);
xnor U31124 (N_31124,N_28422,N_28002);
nand U31125 (N_31125,N_26654,N_26915);
xnor U31126 (N_31126,N_25516,N_27608);
and U31127 (N_31127,N_27173,N_29679);
nor U31128 (N_31128,N_25513,N_25434);
nor U31129 (N_31129,N_27539,N_27906);
or U31130 (N_31130,N_26873,N_25991);
xnor U31131 (N_31131,N_27214,N_29249);
and U31132 (N_31132,N_26771,N_27078);
or U31133 (N_31133,N_25609,N_26022);
and U31134 (N_31134,N_26867,N_26895);
nor U31135 (N_31135,N_25679,N_26355);
xor U31136 (N_31136,N_26990,N_26698);
nand U31137 (N_31137,N_26371,N_29613);
and U31138 (N_31138,N_26196,N_26491);
nor U31139 (N_31139,N_26678,N_27585);
or U31140 (N_31140,N_25390,N_26209);
nor U31141 (N_31141,N_27195,N_26129);
xnor U31142 (N_31142,N_25884,N_25185);
nor U31143 (N_31143,N_27683,N_29555);
or U31144 (N_31144,N_26999,N_29964);
nand U31145 (N_31145,N_27530,N_27381);
nor U31146 (N_31146,N_28611,N_27632);
nand U31147 (N_31147,N_27797,N_28749);
or U31148 (N_31148,N_27433,N_27689);
nand U31149 (N_31149,N_28998,N_26157);
and U31150 (N_31150,N_28718,N_28828);
xnor U31151 (N_31151,N_29394,N_27854);
nor U31152 (N_31152,N_25573,N_28428);
nand U31153 (N_31153,N_26068,N_29493);
and U31154 (N_31154,N_25374,N_27206);
nand U31155 (N_31155,N_25790,N_27766);
and U31156 (N_31156,N_25789,N_25581);
nand U31157 (N_31157,N_25035,N_26842);
or U31158 (N_31158,N_27706,N_28107);
or U31159 (N_31159,N_28947,N_29038);
nand U31160 (N_31160,N_28928,N_28454);
and U31161 (N_31161,N_28063,N_29092);
nor U31162 (N_31162,N_27159,N_28010);
or U31163 (N_31163,N_26458,N_27476);
nor U31164 (N_31164,N_26151,N_28984);
xor U31165 (N_31165,N_28614,N_26562);
and U31166 (N_31166,N_25235,N_25356);
xnor U31167 (N_31167,N_27829,N_27095);
xor U31168 (N_31168,N_25697,N_25768);
and U31169 (N_31169,N_26795,N_26717);
nor U31170 (N_31170,N_28665,N_29323);
xnor U31171 (N_31171,N_29717,N_27065);
and U31172 (N_31172,N_28952,N_26664);
and U31173 (N_31173,N_26730,N_27017);
and U31174 (N_31174,N_26126,N_29128);
and U31175 (N_31175,N_27774,N_27406);
and U31176 (N_31176,N_28960,N_29530);
and U31177 (N_31177,N_28996,N_29342);
or U31178 (N_31178,N_27777,N_25219);
xnor U31179 (N_31179,N_28091,N_29797);
nand U31180 (N_31180,N_26186,N_29701);
nor U31181 (N_31181,N_28519,N_27933);
nand U31182 (N_31182,N_27794,N_29041);
and U31183 (N_31183,N_25506,N_26687);
or U31184 (N_31184,N_27072,N_27484);
nand U31185 (N_31185,N_28361,N_26711);
and U31186 (N_31186,N_26552,N_26445);
and U31187 (N_31187,N_26114,N_27279);
nand U31188 (N_31188,N_28545,N_27475);
xnor U31189 (N_31189,N_25570,N_29572);
and U31190 (N_31190,N_25638,N_25317);
xor U31191 (N_31191,N_27977,N_26108);
nand U31192 (N_31192,N_28198,N_27032);
and U31193 (N_31193,N_26218,N_26845);
nor U31194 (N_31194,N_26510,N_26972);
nand U31195 (N_31195,N_28284,N_25751);
nor U31196 (N_31196,N_28917,N_25906);
nor U31197 (N_31197,N_26132,N_26060);
or U31198 (N_31198,N_25041,N_26586);
or U31199 (N_31199,N_29681,N_28892);
nor U31200 (N_31200,N_27778,N_28108);
and U31201 (N_31201,N_27543,N_28846);
xor U31202 (N_31202,N_27895,N_27347);
and U31203 (N_31203,N_25488,N_26741);
xnor U31204 (N_31204,N_25005,N_28877);
xor U31205 (N_31205,N_27765,N_27499);
or U31206 (N_31206,N_28954,N_27672);
xnor U31207 (N_31207,N_26354,N_27989);
xnor U31208 (N_31208,N_26101,N_28423);
nor U31209 (N_31209,N_26614,N_28161);
or U31210 (N_31210,N_25464,N_27814);
or U31211 (N_31211,N_25664,N_27835);
or U31212 (N_31212,N_25718,N_26875);
nor U31213 (N_31213,N_25306,N_28039);
nand U31214 (N_31214,N_28021,N_28886);
and U31215 (N_31215,N_26241,N_28966);
or U31216 (N_31216,N_26053,N_28666);
xor U31217 (N_31217,N_28190,N_27116);
nand U31218 (N_31218,N_29025,N_26661);
nand U31219 (N_31219,N_25279,N_27084);
or U31220 (N_31220,N_28857,N_29545);
xnor U31221 (N_31221,N_27232,N_26897);
and U31222 (N_31222,N_28882,N_28147);
xor U31223 (N_31223,N_25320,N_25470);
and U31224 (N_31224,N_26955,N_28341);
nand U31225 (N_31225,N_28397,N_28059);
nor U31226 (N_31226,N_28457,N_27886);
nand U31227 (N_31227,N_27662,N_25683);
xor U31228 (N_31228,N_29962,N_26036);
xor U31229 (N_31229,N_25368,N_27446);
nand U31230 (N_31230,N_28774,N_29606);
and U31231 (N_31231,N_26575,N_27260);
xor U31232 (N_31232,N_29766,N_26745);
or U31233 (N_31233,N_28483,N_26651);
or U31234 (N_31234,N_25229,N_26356);
xnor U31235 (N_31235,N_26488,N_29971);
and U31236 (N_31236,N_29724,N_26394);
or U31237 (N_31237,N_26624,N_29668);
nand U31238 (N_31238,N_25446,N_26708);
or U31239 (N_31239,N_25419,N_25217);
nor U31240 (N_31240,N_28156,N_26067);
xnor U31241 (N_31241,N_28921,N_28548);
nand U31242 (N_31242,N_29537,N_27841);
or U31243 (N_31243,N_27571,N_27745);
and U31244 (N_31244,N_26509,N_26118);
and U31245 (N_31245,N_25083,N_26912);
or U31246 (N_31246,N_25893,N_28761);
nand U31247 (N_31247,N_25308,N_27048);
or U31248 (N_31248,N_29842,N_25841);
nor U31249 (N_31249,N_28020,N_29745);
nand U31250 (N_31250,N_25431,N_26479);
or U31251 (N_31251,N_26050,N_25532);
or U31252 (N_31252,N_28949,N_25262);
or U31253 (N_31253,N_29605,N_27063);
nor U31254 (N_31254,N_29542,N_29630);
nor U31255 (N_31255,N_29412,N_25560);
nor U31256 (N_31256,N_27651,N_29473);
xor U31257 (N_31257,N_25351,N_26609);
nor U31258 (N_31258,N_27951,N_26299);
xnor U31259 (N_31259,N_26503,N_26304);
nor U31260 (N_31260,N_27998,N_27248);
and U31261 (N_31261,N_29158,N_25452);
xor U31262 (N_31262,N_28100,N_29214);
and U31263 (N_31263,N_27025,N_25641);
xor U31264 (N_31264,N_28809,N_26908);
and U31265 (N_31265,N_27278,N_26834);
xor U31266 (N_31266,N_26160,N_29258);
nand U31267 (N_31267,N_26865,N_28870);
xnor U31268 (N_31268,N_29870,N_29460);
nand U31269 (N_31269,N_29518,N_26474);
or U31270 (N_31270,N_25209,N_25716);
and U31271 (N_31271,N_25274,N_25961);
and U31272 (N_31272,N_26174,N_29756);
xnor U31273 (N_31273,N_27990,N_28505);
nor U31274 (N_31274,N_25627,N_29360);
xor U31275 (N_31275,N_25748,N_27236);
and U31276 (N_31276,N_26507,N_29958);
and U31277 (N_31277,N_28900,N_29123);
nand U31278 (N_31278,N_27629,N_27089);
nand U31279 (N_31279,N_25135,N_25008);
or U31280 (N_31280,N_28883,N_27907);
xor U31281 (N_31281,N_26073,N_26180);
xnor U31282 (N_31282,N_27624,N_25934);
nor U31283 (N_31283,N_28302,N_26133);
nor U31284 (N_31284,N_27407,N_28033);
or U31285 (N_31285,N_27741,N_25885);
nand U31286 (N_31286,N_27534,N_25002);
nor U31287 (N_31287,N_29919,N_27852);
xnor U31288 (N_31288,N_25845,N_28172);
or U31289 (N_31289,N_27544,N_26437);
nand U31290 (N_31290,N_29570,N_25665);
nand U31291 (N_31291,N_25177,N_28057);
and U31292 (N_31292,N_26248,N_29468);
xor U31293 (N_31293,N_29757,N_25230);
xor U31294 (N_31294,N_25872,N_27559);
and U31295 (N_31295,N_28588,N_28850);
nor U31296 (N_31296,N_27031,N_26029);
nand U31297 (N_31297,N_29224,N_28987);
nor U31298 (N_31298,N_26385,N_25292);
nand U31299 (N_31299,N_29273,N_25959);
nor U31300 (N_31300,N_28101,N_29379);
and U31301 (N_31301,N_29932,N_29423);
or U31302 (N_31302,N_27899,N_27828);
nand U31303 (N_31303,N_29122,N_28899);
nor U31304 (N_31304,N_26523,N_29837);
or U31305 (N_31305,N_28046,N_29776);
xor U31306 (N_31306,N_26685,N_28909);
xor U31307 (N_31307,N_25453,N_28077);
nor U31308 (N_31308,N_28271,N_29631);
nand U31309 (N_31309,N_25011,N_27377);
and U31310 (N_31310,N_25325,N_25422);
nor U31311 (N_31311,N_26931,N_29034);
and U31312 (N_31312,N_25327,N_28728);
and U31313 (N_31313,N_28013,N_28289);
or U31314 (N_31314,N_25844,N_29660);
nand U31315 (N_31315,N_29359,N_26359);
or U31316 (N_31316,N_26123,N_28580);
or U31317 (N_31317,N_28852,N_27449);
or U31318 (N_31318,N_25164,N_25168);
nor U31319 (N_31319,N_27859,N_28112);
nand U31320 (N_31320,N_26684,N_29026);
nand U31321 (N_31321,N_26165,N_27598);
nand U31322 (N_31322,N_28616,N_25864);
xnor U31323 (N_31323,N_29251,N_29740);
nand U31324 (N_31324,N_29510,N_25940);
and U31325 (N_31325,N_27477,N_25335);
nor U31326 (N_31326,N_27523,N_25792);
nor U31327 (N_31327,N_26639,N_26236);
and U31328 (N_31328,N_25099,N_27707);
nor U31329 (N_31329,N_25801,N_26974);
and U31330 (N_31330,N_29779,N_29490);
or U31331 (N_31331,N_27671,N_28296);
or U31332 (N_31332,N_28730,N_27663);
xnor U31333 (N_31333,N_27257,N_26929);
nand U31334 (N_31334,N_25997,N_29247);
nand U31335 (N_31335,N_29244,N_27334);
nor U31336 (N_31336,N_29889,N_27429);
nor U31337 (N_31337,N_25607,N_26600);
and U31338 (N_31338,N_29202,N_29327);
xor U31339 (N_31339,N_25713,N_26267);
nand U31340 (N_31340,N_28371,N_28537);
nor U31341 (N_31341,N_27702,N_28314);
nor U31342 (N_31342,N_29220,N_28777);
and U31343 (N_31343,N_25033,N_29946);
nand U31344 (N_31344,N_28425,N_25111);
nor U31345 (N_31345,N_25773,N_25965);
xor U31346 (N_31346,N_29944,N_27913);
and U31347 (N_31347,N_27486,N_26880);
or U31348 (N_31348,N_25386,N_26321);
nand U31349 (N_31349,N_29895,N_25672);
nor U31350 (N_31350,N_28294,N_28199);
nand U31351 (N_31351,N_29062,N_26725);
nand U31352 (N_31352,N_28864,N_27871);
and U31353 (N_31353,N_26776,N_29392);
and U31354 (N_31354,N_28081,N_26011);
nor U31355 (N_31355,N_29471,N_25369);
xor U31356 (N_31356,N_26998,N_25148);
nor U31357 (N_31357,N_27861,N_25661);
nand U31358 (N_31358,N_26989,N_27131);
and U31359 (N_31359,N_25287,N_25248);
or U31360 (N_31360,N_27635,N_27370);
nand U31361 (N_31361,N_28382,N_27424);
or U31362 (N_31362,N_29375,N_26837);
and U31363 (N_31363,N_25653,N_28263);
nand U31364 (N_31364,N_28398,N_28668);
and U31365 (N_31365,N_27445,N_25007);
and U31366 (N_31366,N_27704,N_29821);
and U31367 (N_31367,N_26951,N_25460);
nor U31368 (N_31368,N_28380,N_29324);
nor U31369 (N_31369,N_27457,N_29811);
xnor U31370 (N_31370,N_28169,N_29573);
nor U31371 (N_31371,N_27099,N_27826);
nor U31372 (N_31372,N_29659,N_27916);
nor U31373 (N_31373,N_29698,N_29358);
nand U31374 (N_31374,N_25974,N_29750);
or U31375 (N_31375,N_27365,N_28741);
and U31376 (N_31376,N_27547,N_27315);
xnor U31377 (N_31377,N_28258,N_28464);
or U31378 (N_31378,N_28038,N_25518);
nand U31379 (N_31379,N_28338,N_28555);
nor U31380 (N_31380,N_26750,N_29110);
or U31381 (N_31381,N_29543,N_25642);
nor U31382 (N_31382,N_28506,N_25966);
or U31383 (N_31383,N_26777,N_27939);
nand U31384 (N_31384,N_27160,N_26210);
xnor U31385 (N_31385,N_26533,N_26546);
nor U31386 (N_31386,N_28335,N_28226);
nor U31387 (N_31387,N_29383,N_27473);
nor U31388 (N_31388,N_29920,N_29663);
and U31389 (N_31389,N_25029,N_28961);
nand U31390 (N_31390,N_29942,N_26968);
xnor U31391 (N_31391,N_25575,N_28866);
nand U31392 (N_31392,N_25823,N_25833);
nand U31393 (N_31393,N_28414,N_25947);
nor U31394 (N_31394,N_25557,N_26797);
xnor U31395 (N_31395,N_25978,N_27812);
or U31396 (N_31396,N_25733,N_27262);
nor U31397 (N_31397,N_28201,N_26647);
or U31398 (N_31398,N_26650,N_26554);
and U31399 (N_31399,N_28328,N_28300);
or U31400 (N_31400,N_28770,N_25584);
xor U31401 (N_31401,N_28936,N_25774);
nand U31402 (N_31402,N_29847,N_26275);
nand U31403 (N_31403,N_27296,N_29900);
nand U31404 (N_31404,N_26577,N_28000);
nor U31405 (N_31405,N_26369,N_29318);
or U31406 (N_31406,N_27355,N_27569);
xnor U31407 (N_31407,N_25788,N_26113);
and U31408 (N_31408,N_26259,N_29255);
nor U31409 (N_31409,N_27092,N_29851);
nand U31410 (N_31410,N_25215,N_27339);
or U31411 (N_31411,N_26482,N_26876);
or U31412 (N_31412,N_28641,N_29408);
and U31413 (N_31413,N_25647,N_28163);
and U31414 (N_31414,N_29674,N_26996);
nor U31415 (N_31415,N_29506,N_27383);
nand U31416 (N_31416,N_27867,N_27335);
nor U31417 (N_31417,N_26976,N_25240);
and U31418 (N_31418,N_29019,N_29385);
xor U31419 (N_31419,N_27803,N_28871);
nor U31420 (N_31420,N_29329,N_29706);
or U31421 (N_31421,N_26465,N_25975);
and U31422 (N_31422,N_27984,N_29387);
nand U31423 (N_31423,N_29344,N_29278);
or U31424 (N_31424,N_26403,N_29015);
nand U31425 (N_31425,N_27062,N_25310);
nand U31426 (N_31426,N_25186,N_25423);
or U31427 (N_31427,N_26799,N_26862);
and U31428 (N_31428,N_27052,N_26273);
xnor U31429 (N_31429,N_27666,N_26705);
and U31430 (N_31430,N_27096,N_29777);
nor U31431 (N_31431,N_29791,N_28492);
xnor U31432 (N_31432,N_28432,N_28788);
or U31433 (N_31433,N_28114,N_27566);
or U31434 (N_31434,N_29690,N_29016);
xor U31435 (N_31435,N_25888,N_26217);
and U31436 (N_31436,N_27354,N_28923);
nand U31437 (N_31437,N_28743,N_26948);
xnor U31438 (N_31438,N_25271,N_26254);
xnor U31439 (N_31439,N_26497,N_27292);
xnor U31440 (N_31440,N_25696,N_25674);
xor U31441 (N_31441,N_25190,N_26737);
nor U31442 (N_31442,N_28074,N_28171);
and U31443 (N_31443,N_27183,N_29063);
nand U31444 (N_31444,N_27154,N_29643);
nand U31445 (N_31445,N_25724,N_27790);
nor U31446 (N_31446,N_27526,N_29297);
or U31447 (N_31447,N_27769,N_26828);
nor U31448 (N_31448,N_29644,N_28865);
nor U31449 (N_31449,N_29193,N_27982);
or U31450 (N_31450,N_26087,N_25318);
or U31451 (N_31451,N_28908,N_27067);
or U31452 (N_31452,N_27443,N_29666);
and U31453 (N_31453,N_29599,N_28243);
xnor U31454 (N_31454,N_26589,N_29521);
nor U31455 (N_31455,N_26179,N_25698);
xnor U31456 (N_31456,N_27548,N_29739);
and U31457 (N_31457,N_29671,N_25891);
and U31458 (N_31458,N_29002,N_25064);
nand U31459 (N_31459,N_27211,N_27171);
nand U31460 (N_31460,N_29429,N_27245);
or U31461 (N_31461,N_28391,N_29906);
nor U31462 (N_31462,N_25692,N_25359);
or U31463 (N_31463,N_26316,N_29600);
xnor U31464 (N_31464,N_25415,N_26481);
and U31465 (N_31465,N_25070,N_26907);
and U31466 (N_31466,N_28638,N_29236);
nor U31467 (N_31467,N_27970,N_26879);
xor U31468 (N_31468,N_29402,N_28001);
nor U31469 (N_31469,N_28355,N_27808);
nand U31470 (N_31470,N_28340,N_25354);
and U31471 (N_31471,N_26838,N_27974);
nand U31472 (N_31472,N_28969,N_29998);
nand U31473 (N_31473,N_29938,N_29347);
nor U31474 (N_31474,N_27514,N_28288);
nor U31475 (N_31475,N_27600,N_29491);
and U31476 (N_31476,N_29623,N_25898);
or U31477 (N_31477,N_27848,N_26525);
xnor U31478 (N_31478,N_29781,N_29864);
xor U31479 (N_31479,N_25237,N_27888);
nand U31480 (N_31480,N_27677,N_26764);
nand U31481 (N_31481,N_27420,N_29410);
nor U31482 (N_31482,N_28640,N_27634);
or U31483 (N_31483,N_25530,N_25882);
xnor U31484 (N_31484,N_26904,N_28158);
nor U31485 (N_31485,N_26024,N_27482);
nor U31486 (N_31486,N_28504,N_27610);
or U31487 (N_31487,N_28674,N_25006);
xor U31488 (N_31488,N_28570,N_25860);
nor U31489 (N_31489,N_26429,N_29317);
and U31490 (N_31490,N_25785,N_29737);
nor U31491 (N_31491,N_28810,N_28327);
xor U31492 (N_31492,N_27742,N_26779);
or U31493 (N_31493,N_27997,N_26357);
nor U31494 (N_31494,N_27557,N_29405);
nor U31495 (N_31495,N_27133,N_27698);
nand U31496 (N_31496,N_29259,N_26801);
nand U31497 (N_31497,N_27827,N_27410);
or U31498 (N_31498,N_28242,N_25770);
nor U31499 (N_31499,N_25298,N_27060);
xor U31500 (N_31500,N_27273,N_28627);
and U31501 (N_31501,N_27184,N_28287);
nand U31502 (N_31502,N_26052,N_29548);
nor U31503 (N_31503,N_29810,N_28080);
nor U31504 (N_31504,N_29036,N_29676);
nor U31505 (N_31505,N_27811,N_25212);
xnor U31506 (N_31506,N_25150,N_26007);
nand U31507 (N_31507,N_26805,N_27695);
nand U31508 (N_31508,N_29064,N_26911);
nor U31509 (N_31509,N_25588,N_29134);
nor U31510 (N_31510,N_26461,N_25639);
or U31511 (N_31511,N_25384,N_29112);
or U31512 (N_31512,N_28518,N_28313);
nand U31513 (N_31513,N_27876,N_29722);
or U31514 (N_31514,N_25239,N_28930);
nor U31515 (N_31515,N_25032,N_25244);
xor U31516 (N_31516,N_26560,N_25524);
or U31517 (N_31517,N_26956,N_29280);
xor U31518 (N_31518,N_25757,N_26667);
nand U31519 (N_31519,N_27574,N_25964);
and U31520 (N_31520,N_27577,N_28839);
and U31521 (N_31521,N_28812,N_26676);
and U31522 (N_31522,N_28717,N_29547);
nor U31523 (N_31523,N_27979,N_27300);
nor U31524 (N_31524,N_25663,N_28308);
and U31525 (N_31525,N_27653,N_28356);
or U31526 (N_31526,N_29355,N_28336);
nand U31527 (N_31527,N_25257,N_25709);
nand U31528 (N_31528,N_25378,N_26462);
and U31529 (N_31529,N_26872,N_27352);
or U31530 (N_31530,N_29844,N_29362);
or U31531 (N_31531,N_26881,N_26748);
nand U31532 (N_31532,N_29260,N_29908);
and U31533 (N_31533,N_27348,N_29568);
or U31534 (N_31534,N_27045,N_28111);
and U31535 (N_31535,N_26743,N_27270);
xnor U31536 (N_31536,N_29208,N_29845);
or U31537 (N_31537,N_28562,N_26466);
xor U31538 (N_31538,N_28092,N_28902);
nand U31539 (N_31539,N_28619,N_28030);
or U31540 (N_31540,N_25863,N_26690);
or U31541 (N_31541,N_29912,N_29459);
xor U31542 (N_31542,N_25813,N_26796);
nand U31543 (N_31543,N_27492,N_26005);
or U31544 (N_31544,N_26576,N_26744);
and U31545 (N_31545,N_29556,N_28303);
and U31546 (N_31546,N_27004,N_28701);
or U31547 (N_31547,N_25382,N_28213);
nor U31548 (N_31548,N_26463,N_28144);
or U31549 (N_31549,N_25113,N_26416);
or U31550 (N_31550,N_29972,N_26207);
nand U31551 (N_31551,N_28661,N_26695);
xnor U31552 (N_31552,N_27138,N_26135);
nor U31553 (N_31553,N_25943,N_25134);
or U31554 (N_31554,N_29440,N_25615);
xnor U31555 (N_31555,N_25739,N_26270);
nor U31556 (N_31556,N_26168,N_26673);
xor U31557 (N_31557,N_26970,N_26023);
xor U31558 (N_31558,N_29758,N_29238);
xor U31559 (N_31559,N_27371,N_27567);
nor U31560 (N_31560,N_25145,N_25915);
nand U31561 (N_31561,N_29271,N_27963);
or U31562 (N_31562,N_28018,N_26606);
nand U31563 (N_31563,N_26793,N_29876);
and U31564 (N_31564,N_28957,N_25753);
xor U31565 (N_31565,N_29198,N_28723);
or U31566 (N_31566,N_26042,N_26018);
nor U31567 (N_31567,N_29768,N_28896);
nor U31568 (N_31568,N_25194,N_26347);
xor U31569 (N_31569,N_25626,N_25206);
or U31570 (N_31570,N_26339,N_28342);
xor U31571 (N_31571,N_27945,N_25586);
nand U31572 (N_31572,N_26163,N_29727);
nand U31573 (N_31573,N_28084,N_28629);
or U31574 (N_31574,N_25412,N_27495);
xnor U31575 (N_31575,N_25472,N_25956);
or U31576 (N_31576,N_29366,N_28334);
and U31577 (N_31577,N_27014,N_27616);
and U31578 (N_31578,N_28706,N_29826);
nand U31579 (N_31579,N_25566,N_28489);
nand U31580 (N_31580,N_26987,N_26623);
or U31581 (N_31581,N_29751,N_27664);
or U31582 (N_31582,N_27862,N_26397);
nor U31583 (N_31583,N_25680,N_27186);
nor U31584 (N_31584,N_25535,N_28388);
and U31585 (N_31585,N_26709,N_28609);
or U31586 (N_31586,N_28122,N_29296);
nor U31587 (N_31587,N_26827,N_28992);
xor U31588 (N_31588,N_27301,N_27593);
nand U31589 (N_31589,N_26957,N_28415);
xor U31590 (N_31590,N_29649,N_29899);
nor U31591 (N_31591,N_26324,N_26882);
nor U31592 (N_31592,N_25819,N_27073);
nor U31593 (N_31593,N_26384,N_29767);
nand U31594 (N_31594,N_26313,N_27403);
and U31595 (N_31595,N_25268,N_29496);
nor U31596 (N_31596,N_29617,N_27136);
xor U31597 (N_31597,N_26724,N_25735);
and U31598 (N_31598,N_27080,N_29281);
xnor U31599 (N_31599,N_29820,N_27243);
and U31600 (N_31600,N_27192,N_28943);
or U31601 (N_31601,N_27937,N_29611);
and U31602 (N_31602,N_25809,N_25859);
xor U31603 (N_31603,N_25430,N_27681);
and U31604 (N_31604,N_29685,N_27533);
nor U31605 (N_31605,N_28136,N_25522);
xnor U31606 (N_31606,N_26185,N_26841);
and U31607 (N_31607,N_28133,N_28847);
nor U31608 (N_31608,N_26048,N_26517);
xor U31609 (N_31609,N_28123,N_25624);
and U31610 (N_31610,N_29237,N_27140);
or U31611 (N_31611,N_29196,N_29267);
or U31612 (N_31612,N_26632,N_26003);
and U31613 (N_31613,N_28255,N_29734);
xor U31614 (N_31614,N_28034,N_28543);
and U31615 (N_31615,N_27929,N_29314);
or U31616 (N_31616,N_29014,N_26432);
or U31617 (N_31617,N_26285,N_28978);
and U31618 (N_31618,N_28979,N_29161);
nand U31619 (N_31619,N_28920,N_28239);
nor U31620 (N_31620,N_25827,N_26072);
nand U31621 (N_31621,N_29438,N_29130);
or U31622 (N_31622,N_27602,N_29933);
and U31623 (N_31623,N_25290,N_25887);
or U31624 (N_31624,N_28085,N_27893);
or U31625 (N_31625,N_29117,N_26176);
nand U31626 (N_31626,N_25883,N_29714);
nand U31627 (N_31627,N_26993,N_26815);
xor U31628 (N_31628,N_28557,N_27392);
or U31629 (N_31629,N_28738,N_26124);
nor U31630 (N_31630,N_26239,N_28677);
and U31631 (N_31631,N_29486,N_27331);
nand U31632 (N_31632,N_28692,N_26107);
and U31633 (N_31633,N_28800,N_27510);
nand U31634 (N_31634,N_26615,N_25957);
nor U31635 (N_31635,N_25875,N_29684);
and U31636 (N_31636,N_27748,N_27985);
and U31637 (N_31637,N_26866,N_26538);
nor U31638 (N_31638,N_26670,N_29635);
or U31639 (N_31639,N_25383,N_28985);
and U31640 (N_31640,N_28779,N_25276);
xor U31641 (N_31641,N_29983,N_25091);
nand U31642 (N_31642,N_26361,N_28354);
nor U31643 (N_31643,N_29489,N_26630);
and U31644 (N_31644,N_27272,N_29736);
nand U31645 (N_31645,N_25593,N_26256);
or U31646 (N_31646,N_28298,N_29364);
or U31647 (N_31647,N_27288,N_29725);
nor U31648 (N_31648,N_29331,N_26092);
xor U31649 (N_31649,N_28323,N_26139);
xor U31650 (N_31650,N_26986,N_27500);
xnor U31651 (N_31651,N_27379,N_27881);
xor U31652 (N_31652,N_25449,N_25908);
and U31653 (N_31653,N_28274,N_27324);
nor U31654 (N_31654,N_28097,N_26156);
xor U31655 (N_31655,N_25704,N_25677);
nor U31656 (N_31656,N_28775,N_25319);
nand U31657 (N_31657,N_29472,N_28044);
or U31658 (N_31658,N_25951,N_25174);
xnor U31659 (N_31659,N_29420,N_25016);
nor U31660 (N_31660,N_26184,N_25850);
or U31661 (N_31661,N_25249,N_28858);
nand U31662 (N_31662,N_26569,N_26652);
nand U31663 (N_31663,N_25260,N_27991);
nand U31664 (N_31664,N_29476,N_25154);
nor U31665 (N_31665,N_29308,N_28148);
xor U31666 (N_31666,N_29225,N_25115);
and U31667 (N_31667,N_29645,N_27717);
xor U31668 (N_31668,N_29819,N_25401);
xnor U31669 (N_31669,N_27750,N_25688);
xnor U31670 (N_31670,N_28566,N_29190);
xnor U31671 (N_31671,N_25477,N_25275);
and U31672 (N_31672,N_28076,N_26227);
xor U31673 (N_31673,N_25385,N_26448);
nand U31674 (N_31674,N_29999,N_28868);
or U31675 (N_31675,N_29056,N_25636);
nand U31676 (N_31676,N_28569,N_26122);
or U31677 (N_31677,N_28914,N_27837);
nor U31678 (N_31678,N_27525,N_25300);
or U31679 (N_31679,N_28032,N_29655);
nor U31680 (N_31680,N_28533,N_25643);
and U31681 (N_31681,N_25778,N_26365);
and U31682 (N_31682,N_28373,N_27673);
nand U31683 (N_31683,N_25707,N_27125);
or U31684 (N_31684,N_26596,N_27330);
xnor U31685 (N_31685,N_28374,N_29678);
and U31686 (N_31686,N_27969,N_27167);
xor U31687 (N_31687,N_29108,N_28634);
nand U31688 (N_31688,N_28140,N_26333);
and U31689 (N_31689,N_27150,N_27914);
nor U31690 (N_31690,N_25056,N_26545);
and U31691 (N_31691,N_25604,N_29457);
nor U31692 (N_31692,N_26020,N_26131);
and U31693 (N_31693,N_28120,N_25073);
nand U31694 (N_31694,N_29652,N_26696);
or U31695 (N_31695,N_27967,N_26206);
xnor U31696 (N_31696,N_26757,N_29389);
or U31697 (N_31697,N_27938,N_29377);
xnor U31698 (N_31698,N_27230,N_25620);
xor U31699 (N_31699,N_25376,N_28523);
or U31700 (N_31700,N_28036,N_25089);
nand U31701 (N_31701,N_28325,N_28370);
nand U31702 (N_31702,N_29315,N_28873);
or U31703 (N_31703,N_28339,N_28051);
nand U31704 (N_31704,N_26857,N_28012);
or U31705 (N_31705,N_25307,N_29523);
nor U31706 (N_31706,N_26439,N_25023);
or U31707 (N_31707,N_25413,N_25349);
xnor U31708 (N_31708,N_28529,N_27714);
and U31709 (N_31709,N_25594,N_26792);
or U31710 (N_31710,N_28485,N_29602);
xor U31711 (N_31711,N_28711,N_28630);
xor U31712 (N_31712,N_26758,N_25762);
xnor U31713 (N_31713,N_26938,N_28526);
or U31714 (N_31714,N_29836,N_26973);
and U31715 (N_31715,N_29534,N_28753);
nor U31716 (N_31716,N_25977,N_25727);
or U31717 (N_31717,N_29883,N_27479);
nor U31718 (N_31718,N_28153,N_25036);
and U31719 (N_31719,N_28586,N_26716);
and U31720 (N_31720,N_27128,N_25429);
or U31721 (N_31721,N_27427,N_29119);
or U31722 (N_31722,N_28009,N_29564);
nor U31723 (N_31723,N_26558,N_29772);
or U31724 (N_31724,N_28278,N_26161);
and U31725 (N_31725,N_26518,N_27464);
xnor U31726 (N_31726,N_27844,N_29607);
and U31727 (N_31727,N_29891,N_26187);
xnor U31728 (N_31728,N_26821,N_27621);
or U31729 (N_31729,N_28632,N_26511);
nand U31730 (N_31730,N_29445,N_25191);
or U31731 (N_31731,N_29669,N_25109);
xor U31732 (N_31732,N_27850,N_26352);
or U31733 (N_31733,N_28907,N_26585);
and U31734 (N_31734,N_28702,N_25662);
nor U31735 (N_31735,N_29677,N_25092);
xnor U31736 (N_31736,N_26713,N_28248);
nand U31737 (N_31737,N_25972,N_26953);
nand U31738 (N_31738,N_29627,N_26906);
and U31739 (N_31739,N_26958,N_26498);
and U31740 (N_31740,N_27071,N_28186);
xor U31741 (N_31741,N_26660,N_28387);
xnor U31742 (N_31742,N_25540,N_25769);
nor U31743 (N_31743,N_25027,N_28691);
nor U31744 (N_31744,N_25984,N_26922);
or U31745 (N_31745,N_27149,N_29464);
or U31746 (N_31746,N_28494,N_29749);
nor U31747 (N_31747,N_26785,N_29646);
nand U31748 (N_31748,N_26090,N_25303);
or U31749 (N_31749,N_28803,N_25265);
xor U31750 (N_31750,N_25652,N_25093);
xnor U31751 (N_31751,N_25469,N_28682);
nand U31752 (N_31752,N_26412,N_27298);
and U31753 (N_31753,N_29612,N_27390);
and U31754 (N_31754,N_25944,N_26193);
and U31755 (N_31755,N_28766,N_25223);
xor U31756 (N_31756,N_25531,N_26766);
or U31757 (N_31757,N_25798,N_27948);
or U31758 (N_31758,N_29708,N_25406);
nand U31759 (N_31759,N_27083,N_25408);
and U31760 (N_31760,N_26079,N_27163);
and U31761 (N_31761,N_28781,N_26571);
nor U31762 (N_31762,N_29769,N_25904);
nor U31763 (N_31763,N_25068,N_27810);
xnor U31764 (N_31764,N_29888,N_27617);
nand U31765 (N_31765,N_29104,N_26988);
and U31766 (N_31766,N_27468,N_29656);
or U31767 (N_31767,N_28944,N_26147);
and U31768 (N_31768,N_29373,N_28447);
or U31769 (N_31769,N_26629,N_29567);
nand U31770 (N_31770,N_29771,N_29974);
nand U31771 (N_31771,N_25404,N_28680);
and U31772 (N_31772,N_28721,N_25377);
or U31773 (N_31773,N_29235,N_29728);
xor U31774 (N_31774,N_28368,N_29571);
xnor U31775 (N_31775,N_25220,N_27719);
nand U31776 (N_31776,N_25272,N_27222);
or U31777 (N_31777,N_26584,N_27289);
nor U31778 (N_31778,N_26028,N_29439);
nand U31779 (N_31779,N_26208,N_25533);
nand U31780 (N_31780,N_25693,N_28438);
nand U31781 (N_31781,N_29702,N_28127);
or U31782 (N_31782,N_28150,N_29075);
nand U31783 (N_31783,N_29042,N_26885);
nand U31784 (N_31784,N_27224,N_27660);
nor U31785 (N_31785,N_25051,N_26916);
nor U31786 (N_31786,N_25546,N_26847);
nand U31787 (N_31787,N_28516,N_28259);
nand U31788 (N_31788,N_28554,N_28771);
or U31789 (N_31789,N_27749,N_25963);
nor U31790 (N_31790,N_26521,N_28293);
and U31791 (N_31791,N_27258,N_25919);
xor U31792 (N_31792,N_26620,N_28736);
nor U31793 (N_31793,N_29059,N_29022);
xor U31794 (N_31794,N_27511,N_27244);
and U31795 (N_31795,N_29597,N_25061);
nor U31796 (N_31796,N_28286,N_28197);
nand U31797 (N_31797,N_25786,N_29334);
xnor U31798 (N_31798,N_28769,N_25426);
and U31799 (N_31799,N_27318,N_27363);
xnor U31800 (N_31800,N_29099,N_26919);
or U31801 (N_31801,N_29955,N_29415);
nand U31802 (N_31802,N_26065,N_28317);
nand U31803 (N_31803,N_29040,N_28755);
nand U31804 (N_31804,N_28600,N_29905);
nand U31805 (N_31805,N_25314,N_27820);
xor U31806 (N_31806,N_25760,N_27654);
and U31807 (N_31807,N_26427,N_27649);
nand U31808 (N_31808,N_28103,N_29529);
xor U31809 (N_31809,N_27647,N_27772);
nor U31810 (N_31810,N_26607,N_25635);
nand U31811 (N_31811,N_28535,N_28822);
or U31812 (N_31812,N_26514,N_27239);
nand U31813 (N_31813,N_28673,N_27802);
nand U31814 (N_31814,N_29086,N_28086);
nor U31815 (N_31815,N_28497,N_27176);
nand U31816 (N_31816,N_25930,N_27366);
xnor U31817 (N_31817,N_25854,N_26389);
and U31818 (N_31818,N_28745,N_25014);
xor U31819 (N_31819,N_26008,N_25019);
xor U31820 (N_31820,N_26808,N_29348);
and U31821 (N_31821,N_26040,N_26396);
nand U31822 (N_31822,N_28247,N_26634);
and U31823 (N_31823,N_26775,N_25496);
or U31824 (N_31824,N_25210,N_28343);
nand U31825 (N_31825,N_28838,N_25026);
xor U31826 (N_31826,N_28919,N_28016);
and U31827 (N_31827,N_28973,N_29598);
nand U31828 (N_31828,N_25346,N_29763);
or U31829 (N_31829,N_28564,N_27276);
xor U31830 (N_31830,N_28362,N_27659);
and U31831 (N_31831,N_29524,N_26379);
nor U31832 (N_31832,N_25824,N_29215);
nor U31833 (N_31833,N_27068,N_27836);
and U31834 (N_31834,N_27158,N_27983);
nor U31835 (N_31835,N_25105,N_28521);
nand U31836 (N_31836,N_25321,N_27329);
or U31837 (N_31837,N_29170,N_27145);
nor U31838 (N_31838,N_29211,N_27326);
and U31839 (N_31839,N_27783,N_27282);
and U31840 (N_31840,N_26495,N_29827);
xnor U31841 (N_31841,N_29795,N_26530);
and U31842 (N_31842,N_29449,N_28417);
or U31843 (N_31843,N_29007,N_25117);
nand U31844 (N_31844,N_29995,N_28378);
and U31845 (N_31845,N_28146,N_27924);
nor U31846 (N_31846,N_29801,N_28139);
nor U31847 (N_31847,N_27134,N_26820);
nor U31848 (N_31848,N_27344,N_26686);
nor U31849 (N_31849,N_27001,N_28994);
nand U31850 (N_31850,N_25563,N_28015);
nor U31851 (N_31851,N_28143,N_27842);
and U31852 (N_31852,N_26934,N_26178);
xor U31853 (N_31853,N_29709,N_27572);
or U31854 (N_31854,N_28141,N_28525);
nand U31855 (N_31855,N_27042,N_27179);
or U31856 (N_31856,N_26441,N_26603);
or U31857 (N_31857,N_28260,N_29897);
nand U31858 (N_31858,N_27109,N_27804);
and U31859 (N_31859,N_29361,N_27775);
or U31860 (N_31860,N_29641,N_25945);
or U31861 (N_31861,N_26332,N_29601);
nand U31862 (N_31862,N_26580,N_29021);
xor U31863 (N_31863,N_26791,N_27606);
and U31864 (N_31864,N_25550,N_29828);
xnor U31865 (N_31865,N_29245,N_29047);
nand U31866 (N_31866,N_26189,N_26739);
and U31867 (N_31867,N_26078,N_26994);
nor U31868 (N_31868,N_29176,N_27923);
nand U31869 (N_31869,N_28513,N_27290);
nor U31870 (N_31870,N_26853,N_26787);
nand U31871 (N_31871,N_27055,N_25527);
nand U31872 (N_31872,N_28461,N_29129);
or U31873 (N_31873,N_25088,N_29436);
nor U31874 (N_31874,N_25942,N_26031);
and U31875 (N_31875,N_29010,N_28008);
nor U31876 (N_31876,N_27231,N_26222);
and U31877 (N_31877,N_26540,N_27813);
or U31878 (N_31878,N_25759,N_26666);
and U31879 (N_31879,N_28315,N_25179);
xor U31880 (N_31880,N_28459,N_25142);
nand U31881 (N_31881,N_26375,N_27832);
or U31882 (N_31882,N_29116,N_29177);
nand U31883 (N_31883,N_25305,N_29907);
nor U31884 (N_31884,N_25441,N_28551);
nor U31885 (N_31885,N_27644,N_26635);
nor U31886 (N_31886,N_29286,N_28183);
nand U31887 (N_31887,N_27943,N_26230);
nor U31888 (N_31888,N_26788,N_29039);
or U31889 (N_31889,N_26682,N_25277);
or U31890 (N_31890,N_28807,N_28591);
xnor U31891 (N_31891,N_26945,N_29765);
nor U31892 (N_31892,N_29269,N_29894);
nand U31893 (N_31893,N_27303,N_29151);
nor U31894 (N_31894,N_29311,N_25608);
xor U31895 (N_31895,N_29755,N_27721);
or U31896 (N_31896,N_27144,N_25717);
or U31897 (N_31897,N_25913,N_25096);
xor U31898 (N_31898,N_29818,N_26905);
and U31899 (N_31899,N_28211,N_25221);
nor U31900 (N_31900,N_27885,N_29284);
and U31901 (N_31901,N_29929,N_29793);
nand U31902 (N_31902,N_27346,N_27175);
xor U31903 (N_31903,N_28760,N_29604);
xor U31904 (N_31904,N_26002,N_25104);
xnor U31905 (N_31905,N_25160,N_26039);
and U31906 (N_31906,N_26143,N_29290);
and U31907 (N_31907,N_27026,N_28418);
xnor U31908 (N_31908,N_26153,N_25814);
xor U31909 (N_31909,N_28439,N_26903);
xor U31910 (N_31910,N_29302,N_27081);
or U31911 (N_31911,N_29786,N_29458);
or U31912 (N_31912,N_28571,N_29903);
or U31913 (N_31913,N_27976,N_29495);
nand U31914 (N_31914,N_28179,N_27711);
or U31915 (N_31915,N_28124,N_29843);
xnor U31916 (N_31916,N_26137,N_26346);
xor U31917 (N_31917,N_25169,N_26665);
nor U31918 (N_31918,N_28311,N_27738);
nor U31919 (N_31919,N_29973,N_29853);
nand U31920 (N_31920,N_25375,N_27341);
nor U31921 (N_31921,N_28813,N_29519);
nand U31922 (N_31922,N_27177,N_28791);
and U31923 (N_31923,N_29178,N_25302);
nor U31924 (N_31924,N_25380,N_27418);
nor U31925 (N_31925,N_29918,N_27597);
and U31926 (N_31926,N_28729,N_26057);
or U31927 (N_31927,N_27353,N_28862);
nor U31928 (N_31928,N_26251,N_28608);
or U31929 (N_31929,N_28376,N_29407);
or U31930 (N_31930,N_27536,N_29301);
and U31931 (N_31931,N_26570,N_29654);
and U31932 (N_31932,N_27737,N_25509);
xor U31933 (N_31933,N_27019,N_28890);
or U31934 (N_31934,N_27294,N_25614);
or U31935 (N_31935,N_25628,N_29915);
nor U31936 (N_31936,N_27389,N_25673);
xor U31937 (N_31937,N_27560,N_28456);
nor U31938 (N_31938,N_28316,N_27604);
nor U31939 (N_31939,N_26016,N_26447);
nand U31940 (N_31940,N_25574,N_26800);
nor U31941 (N_31941,N_28105,N_28889);
nand U31942 (N_31942,N_29852,N_26030);
xor U31943 (N_31943,N_26536,N_26400);
or U31944 (N_31944,N_28254,N_27111);
and U31945 (N_31945,N_29622,N_29866);
and U31946 (N_31946,N_25146,N_28867);
nand U31947 (N_31947,N_28613,N_25468);
and U31948 (N_31948,N_25811,N_25108);
nor U31949 (N_31949,N_26152,N_28747);
and U31950 (N_31950,N_25528,N_27178);
nand U31951 (N_31951,N_28653,N_25166);
nand U31952 (N_31952,N_29610,N_27590);
and U31953 (N_31953,N_27573,N_28277);
xnor U31954 (N_31954,N_27809,N_25526);
xor U31955 (N_31955,N_26091,N_26656);
and U31956 (N_31956,N_25004,N_29037);
or U31957 (N_31957,N_25766,N_28224);
and U31958 (N_31958,N_25042,N_27959);
and U31959 (N_31959,N_25474,N_27722);
nand U31960 (N_31960,N_27114,N_25655);
xnor U31961 (N_31961,N_28279,N_27926);
nor U31962 (N_31962,N_27961,N_25755);
xor U31963 (N_31963,N_29141,N_29368);
and U31964 (N_31964,N_25352,N_26537);
xor U31965 (N_31965,N_25752,N_29081);
xor U31966 (N_31966,N_25347,N_29527);
nand U31967 (N_31967,N_25245,N_28946);
and U31968 (N_31968,N_27940,N_26572);
or U31969 (N_31969,N_28676,N_26378);
xor U31970 (N_31970,N_29703,N_28559);
and U31971 (N_31971,N_27012,N_29743);
or U31972 (N_31972,N_28249,N_29261);
or U31973 (N_31973,N_25286,N_25706);
nand U31974 (N_31974,N_27235,N_25127);
and U31975 (N_31975,N_26489,N_28853);
and U31976 (N_31976,N_27182,N_26158);
and U31977 (N_31977,N_29118,N_28333);
nor U31978 (N_31978,N_28740,N_26175);
or U31979 (N_31979,N_28660,N_27627);
and U31980 (N_31980,N_29349,N_26914);
nor U31981 (N_31981,N_25253,N_28848);
xnor U31982 (N_31982,N_28206,N_28131);
xor U31983 (N_31983,N_26849,N_28754);
and U31984 (N_31984,N_29095,N_27467);
nor U31985 (N_31985,N_26045,N_27491);
nand U31986 (N_31986,N_28310,N_26601);
xor U31987 (N_31987,N_27864,N_29729);
and U31988 (N_31988,N_27952,N_25973);
and U31989 (N_31989,N_29434,N_26965);
nor U31990 (N_31990,N_28963,N_26229);
nand U31991 (N_31991,N_28989,N_26464);
or U31992 (N_31992,N_26164,N_28959);
and U31993 (N_31993,N_27215,N_25640);
xnor U31994 (N_31994,N_28357,N_26909);
nor U31995 (N_31995,N_28071,N_28732);
or U31996 (N_31996,N_25294,N_29988);
or U31997 (N_31997,N_29147,N_28188);
xnor U31998 (N_31998,N_25048,N_25315);
xor U31999 (N_31999,N_25350,N_29994);
and U32000 (N_32000,N_26493,N_29885);
nand U32001 (N_32001,N_27332,N_28132);
or U32002 (N_32002,N_25667,N_25074);
xor U32003 (N_32003,N_28089,N_27210);
nand U32004 (N_32004,N_26205,N_26742);
and U32005 (N_32005,N_27028,N_27901);
nand U32006 (N_32006,N_27872,N_28622);
and U32007 (N_32007,N_27268,N_26167);
or U32008 (N_32008,N_28267,N_27981);
xnor U32009 (N_32009,N_29935,N_26162);
and U32010 (N_32010,N_25339,N_26200);
xor U32011 (N_32011,N_26237,N_25782);
xnor U32012 (N_32012,N_25880,N_27112);
nand U32013 (N_32013,N_27143,N_27688);
and U32014 (N_32014,N_29939,N_28229);
and U32015 (N_32015,N_27822,N_27920);
nor U32016 (N_32016,N_27165,N_25054);
or U32017 (N_32017,N_26528,N_25791);
and U32018 (N_32018,N_25114,N_27021);
and U32019 (N_32019,N_26368,N_26199);
or U32020 (N_32020,N_28250,N_28842);
and U32021 (N_32021,N_25980,N_26370);
xor U32022 (N_32022,N_25510,N_27284);
nand U32023 (N_32023,N_27640,N_28191);
or U32024 (N_32024,N_27538,N_25367);
nor U32025 (N_32025,N_28045,N_27958);
and U32026 (N_32026,N_25726,N_28744);
and U32027 (N_32027,N_25689,N_25095);
or U32028 (N_32028,N_28937,N_26345);
nand U32029 (N_32029,N_29396,N_28546);
and U32030 (N_32030,N_29456,N_26121);
or U32031 (N_32031,N_26192,N_26373);
xnor U32032 (N_32032,N_25571,N_27953);
nor U32033 (N_32033,N_25846,N_27674);
xnor U32034 (N_32034,N_29209,N_25337);
nand U32035 (N_32035,N_28993,N_26658);
nor U32036 (N_32036,N_26746,N_27661);
or U32037 (N_32037,N_26364,N_25703);
nand U32038 (N_32038,N_25152,N_28802);
and U32039 (N_32039,N_27825,N_26314);
nor U32040 (N_32040,N_29968,N_25106);
or U32041 (N_32041,N_26033,N_27129);
nor U32042 (N_32042,N_28511,N_27450);
or U32043 (N_32043,N_25729,N_27319);
and U32044 (N_32044,N_26408,N_25822);
nand U32045 (N_32045,N_29507,N_25914);
nor U32046 (N_32046,N_29406,N_28731);
and U32047 (N_32047,N_26548,N_29834);
nand U32048 (N_32048,N_25879,N_26233);
nor U32049 (N_32049,N_27219,N_29474);
xor U32050 (N_32050,N_27444,N_27918);
xnor U32051 (N_32051,N_25062,N_25098);
nand U32052 (N_32052,N_26100,N_28903);
and U32053 (N_32053,N_25458,N_25269);
or U32054 (N_32054,N_27234,N_25353);
xor U32055 (N_32055,N_27900,N_26424);
nor U32056 (N_32056,N_29483,N_29265);
nand U32057 (N_32057,N_28507,N_27170);
xnor U32058 (N_32058,N_26014,N_26360);
nor U32059 (N_32059,N_28331,N_29812);
nor U32060 (N_32060,N_26720,N_29782);
nor U32061 (N_32061,N_29923,N_29139);
and U32062 (N_32062,N_25037,N_29146);
nor U32063 (N_32063,N_28610,N_27291);
nand U32064 (N_32064,N_29150,N_28593);
nand U32065 (N_32065,N_26284,N_29120);
nor U32066 (N_32066,N_29882,N_28793);
nor U32067 (N_32067,N_28773,N_28364);
and U32068 (N_32068,N_26204,N_27685);
nand U32069 (N_32069,N_28332,N_27801);
or U32070 (N_32070,N_26840,N_29869);
or U32071 (N_32071,N_28244,N_29792);
nor U32072 (N_32072,N_25309,N_25922);
nand U32073 (N_32073,N_26436,N_28697);
nor U32074 (N_32074,N_29487,N_29163);
and U32075 (N_32075,N_25743,N_29775);
nor U32076 (N_32076,N_29320,N_29949);
nor U32077 (N_32077,N_29925,N_25710);
nor U32078 (N_32078,N_29541,N_25338);
nand U32079 (N_32079,N_29609,N_25861);
and U32080 (N_32080,N_27233,N_28577);
and U32081 (N_32081,N_27650,N_28246);
nand U32082 (N_32082,N_25784,N_28948);
nor U32083 (N_32083,N_26032,N_28421);
nand U32084 (N_32084,N_25475,N_28795);
nor U32085 (N_32085,N_28445,N_28231);
nand U32086 (N_32086,N_27935,N_28029);
nand U32087 (N_32087,N_27047,N_26387);
and U32088 (N_32088,N_28827,N_27579);
nor U32089 (N_32089,N_25435,N_29279);
xnor U32090 (N_32090,N_28824,N_28780);
nor U32091 (N_32091,N_27066,N_25128);
and U32092 (N_32092,N_29080,N_25754);
xor U32093 (N_32093,N_27393,N_28563);
xnor U32094 (N_32094,N_26119,N_29068);
or U32095 (N_32095,N_29633,N_28681);
or U32096 (N_32096,N_29210,N_25129);
nand U32097 (N_32097,N_29841,N_27166);
nor U32098 (N_32098,N_29132,N_25144);
xnor U32099 (N_32099,N_27204,N_27489);
nor U32100 (N_32100,N_26740,N_25448);
nand U32101 (N_32101,N_25282,N_28737);
nor U32102 (N_32102,N_29531,N_26565);
and U32103 (N_32103,N_25935,N_29916);
nor U32104 (N_32104,N_28208,N_29945);
nor U32105 (N_32105,N_26219,N_28804);
and U32106 (N_32106,N_29943,N_25618);
nand U32107 (N_32107,N_28719,N_29082);
or U32108 (N_32108,N_25777,N_26485);
xnor U32109 (N_32109,N_28416,N_25685);
nor U32110 (N_32110,N_26943,N_26566);
nand U32111 (N_32111,N_27805,N_26734);
and U32112 (N_32112,N_28102,N_26351);
xor U32113 (N_32113,N_29186,N_26932);
nor U32114 (N_32114,N_29947,N_26983);
and U32115 (N_32115,N_25909,N_28196);
nor U32116 (N_32116,N_28643,N_25650);
nand U32117 (N_32117,N_29384,N_28927);
nand U32118 (N_32118,N_26910,N_25201);
nor U32119 (N_32119,N_29395,N_29252);
nor U32120 (N_32120,N_27603,N_26326);
nand U32121 (N_32121,N_29316,N_25355);
and U32122 (N_32122,N_25289,N_28455);
and U32123 (N_32123,N_26194,N_29505);
or U32124 (N_32124,N_29846,N_29508);
nor U32125 (N_32125,N_29952,N_27891);
and U32126 (N_32126,N_29626,N_26921);
nor U32127 (N_32127,N_28940,N_25463);
or U32128 (N_32128,N_29528,N_25568);
and U32129 (N_32129,N_29008,N_28539);
nand U32130 (N_32130,N_29730,N_27840);
and U32131 (N_32131,N_28299,N_27978);
nor U32132 (N_32132,N_29253,N_28527);
and U32133 (N_32133,N_27378,N_29071);
nand U32134 (N_32134,N_29696,N_26657);
or U32135 (N_32135,N_25606,N_26083);
nor U32136 (N_32136,N_29857,N_27628);
xnor U32137 (N_32137,N_25311,N_29733);
and U32138 (N_32138,N_25183,N_29762);
or U32139 (N_32139,N_29001,N_25086);
or U32140 (N_32140,N_25542,N_29234);
nand U32141 (N_32141,N_27757,N_28304);
nand U32142 (N_32142,N_29060,N_25156);
xor U32143 (N_32143,N_28301,N_26358);
or U32144 (N_32144,N_28869,N_29356);
nor U32145 (N_32145,N_28204,N_25756);
or U32146 (N_32146,N_25211,N_28942);
nor U32147 (N_32147,N_25187,N_26386);
or U32148 (N_32148,N_25379,N_25155);
nor U32149 (N_32149,N_25039,N_29504);
xnor U32150 (N_32150,N_29712,N_28192);
xnor U32151 (N_32151,N_27220,N_27513);
or U32152 (N_32152,N_25741,N_26142);
nor U32153 (N_32153,N_29748,N_27208);
xnor U32154 (N_32154,N_27124,N_26541);
nand U32155 (N_32155,N_27094,N_27734);
nand U32156 (N_32156,N_27225,N_25807);
and U32157 (N_32157,N_26363,N_25968);
xnor U32158 (N_32158,N_27490,N_26093);
or U32159 (N_32159,N_29341,N_26103);
and U32160 (N_32160,N_26595,N_27187);
or U32161 (N_32161,N_25740,N_25659);
or U32162 (N_32162,N_27267,N_25817);
and U32163 (N_32163,N_27633,N_27682);
or U32164 (N_32164,N_28429,N_29596);
nand U32165 (N_32165,N_28531,N_25988);
xor U32166 (N_32166,N_29867,N_26608);
nor U32167 (N_32167,N_27404,N_28648);
nand U32168 (N_32168,N_25580,N_29959);
and U32169 (N_32169,N_29594,N_26602);
and U32170 (N_32170,N_29094,N_25387);
nor U32171 (N_32171,N_25214,N_27018);
or U32172 (N_32172,N_25162,N_27768);
nor U32173 (N_32173,N_27454,N_27583);
or U32174 (N_32174,N_27615,N_25394);
or U32175 (N_32175,N_26444,N_29187);
and U32176 (N_32176,N_27905,N_25831);
and U32177 (N_32177,N_25597,N_29077);
or U32178 (N_32178,N_25344,N_29914);
or U32179 (N_32179,N_25828,N_25767);
and U32180 (N_32180,N_27447,N_25711);
nand U32181 (N_32181,N_25336,N_25583);
nand U32182 (N_32182,N_29242,N_28592);
nand U32183 (N_32183,N_28117,N_28078);
nand U32184 (N_32184,N_29815,N_25629);
or U32185 (N_32185,N_26467,N_27198);
and U32186 (N_32186,N_26728,N_26638);
and U32187 (N_32187,N_29503,N_26043);
and U32188 (N_32188,N_27860,N_29288);
xor U32189 (N_32189,N_28273,N_26105);
nand U32190 (N_32190,N_28939,N_29558);
and U32191 (N_32191,N_28819,N_29868);
or U32192 (N_32192,N_28053,N_26627);
nor U32193 (N_32193,N_26307,N_25454);
nand U32194 (N_32194,N_27098,N_28602);
nand U32195 (N_32195,N_28379,N_28524);
nand U32196 (N_32196,N_25499,N_27441);
nor U32197 (N_32197,N_26115,N_27594);
and U32198 (N_32198,N_25247,N_28654);
nand U32199 (N_32199,N_26297,N_28733);
nand U32200 (N_32200,N_25937,N_25316);
or U32201 (N_32201,N_29960,N_28482);
and U32202 (N_32202,N_29863,N_25407);
and U32203 (N_32203,N_28393,N_26490);
nor U32204 (N_32204,N_26735,N_25414);
nor U32205 (N_32205,N_25558,N_25878);
or U32206 (N_32206,N_26172,N_29398);
and U32207 (N_32207,N_26981,N_25236);
nand U32208 (N_32208,N_26095,N_25207);
nor U32209 (N_32209,N_27758,N_25045);
xnor U32210 (N_32210,N_27631,N_29173);
nand U32211 (N_32211,N_25986,N_28831);
xnor U32212 (N_32212,N_26173,N_29805);
and U32213 (N_32213,N_27307,N_29577);
xnor U32214 (N_32214,N_29004,N_26470);
nand U32215 (N_32215,N_29291,N_27858);
or U32216 (N_32216,N_25971,N_29065);
and U32217 (N_32217,N_27058,N_27713);
xor U32218 (N_32218,N_25420,N_25371);
and U32219 (N_32219,N_25725,N_26959);
and U32220 (N_32220,N_29197,N_29289);
xnor U32221 (N_32221,N_27980,N_26019);
or U32222 (N_32222,N_26190,N_29985);
or U32223 (N_32223,N_29689,N_27942);
nor U32224 (N_32224,N_29466,N_28282);
nand U32225 (N_32225,N_28360,N_27103);
xor U32226 (N_32226,N_29357,N_26319);
nor U32227 (N_32227,N_29726,N_27380);
or U32228 (N_32228,N_25843,N_27120);
xor U32229 (N_32229,N_29546,N_29003);
xnor U32230 (N_32230,N_25656,N_25196);
xor U32231 (N_32231,N_26512,N_26892);
or U32232 (N_32232,N_28353,N_29218);
and U32233 (N_32233,N_29223,N_29802);
and U32234 (N_32234,N_28037,N_27917);
and U32235 (N_32235,N_26367,N_29619);
nor U32236 (N_32236,N_28687,N_29996);
nor U32237 (N_32237,N_29881,N_25772);
nand U32238 (N_32238,N_27637,N_26789);
nor U32239 (N_32239,N_26863,N_28157);
nor U32240 (N_32240,N_28932,N_27263);
and U32241 (N_32241,N_27364,N_28152);
and U32242 (N_32242,N_25242,N_28837);
nand U32243 (N_32243,N_25552,N_25147);
or U32244 (N_32244,N_27845,N_29675);
or U32245 (N_32245,N_25101,N_27367);
and U32246 (N_32246,N_26626,N_27218);
and U32247 (N_32247,N_26322,N_28194);
nand U32248 (N_32248,N_27297,N_27217);
or U32249 (N_32249,N_27789,N_25312);
nand U32250 (N_32250,N_26960,N_29103);
xnor U32251 (N_32251,N_28861,N_29498);
xor U32252 (N_32252,N_27191,N_25892);
and U32253 (N_32253,N_26475,N_25572);
xnor U32254 (N_32254,N_29835,N_29414);
nand U32255 (N_32255,N_25633,N_26329);
nand U32256 (N_32256,N_27729,N_26574);
xor U32257 (N_32257,N_29159,N_26393);
or U32258 (N_32258,N_27639,N_28460);
nor U32259 (N_32259,N_27041,N_25329);
nor U32260 (N_32260,N_28375,N_25857);
and U32261 (N_32261,N_29372,N_27044);
xor U32262 (N_32262,N_26738,N_29185);
nand U32263 (N_32263,N_28407,N_27703);
and U32264 (N_32264,N_28576,N_26428);
or U32265 (N_32265,N_27265,N_25082);
and U32266 (N_32266,N_27999,N_29647);
and U32267 (N_32267,N_26819,N_28466);
nor U32268 (N_32268,N_29931,N_26111);
and U32269 (N_32269,N_26579,N_27776);
and U32270 (N_32270,N_25199,N_26786);
or U32271 (N_32271,N_28808,N_25728);
nand U32272 (N_32272,N_26610,N_29533);
or U32273 (N_32273,N_29171,N_28958);
and U32274 (N_32274,N_27286,N_29325);
or U32275 (N_32275,N_25712,N_26963);
xnor U32276 (N_32276,N_27880,N_29282);
nand U32277 (N_32277,N_25761,N_29287);
xor U32278 (N_32278,N_29986,N_26342);
nand U32279 (N_32279,N_28541,N_29538);
nand U32280 (N_32280,N_28175,N_27908);
nor U32281 (N_32281,N_25330,N_27362);
nor U32282 (N_32282,N_26337,N_26232);
xor U32283 (N_32283,N_25616,N_29926);
xnor U32284 (N_32284,N_26255,N_28253);
nand U32285 (N_32285,N_26140,N_25053);
or U32286 (N_32286,N_28234,N_29788);
and U32287 (N_32287,N_29790,N_26264);
and U32288 (N_32288,N_26950,N_29877);
or U32289 (N_32289,N_27865,N_28219);
nor U32290 (N_32290,N_26679,N_26404);
nand U32291 (N_32291,N_29859,N_28167);
nand U32292 (N_32292,N_25612,N_28675);
and U32293 (N_32293,N_28469,N_26272);
nand U32294 (N_32294,N_29965,N_25787);
nor U32295 (N_32295,N_29569,N_25137);
nand U32296 (N_32296,N_28825,N_27701);
nor U32297 (N_32297,N_25483,N_28582);
and U32298 (N_32298,N_26075,N_27411);
or U32299 (N_32299,N_28962,N_25804);
nand U32300 (N_32300,N_25079,N_28309);
nand U32301 (N_32301,N_28182,N_28350);
xor U32302 (N_32302,N_27250,N_26125);
nor U32303 (N_32303,N_29992,N_27922);
nor U32304 (N_32304,N_27771,N_29166);
xnor U32305 (N_32305,N_28637,N_29365);
xnor U32306 (N_32306,N_26868,N_28035);
or U32307 (N_32307,N_25184,N_25671);
nand U32308 (N_32308,N_29031,N_29744);
and U32309 (N_32309,N_26835,N_29526);
and U32310 (N_32310,N_25409,N_28911);
or U32311 (N_32311,N_26433,N_28040);
xnor U32312 (N_32312,N_27161,N_28090);
nor U32313 (N_32313,N_25003,N_27369);
or U32314 (N_32314,N_28598,N_25090);
or U32315 (N_32315,N_29294,N_25705);
and U32316 (N_32316,N_26049,N_25561);
nand U32317 (N_32317,N_28330,N_25250);
nand U32318 (N_32318,N_27613,N_25198);
nor U32319 (N_32319,N_28068,N_29127);
nor U32320 (N_32320,N_25990,N_25296);
nor U32321 (N_32321,N_29091,N_29451);
and U32322 (N_32322,N_25600,N_26688);
and U32323 (N_32323,N_26383,N_25544);
nand U32324 (N_32324,N_28762,N_25030);
nand U32325 (N_32325,N_28587,N_28678);
and U32326 (N_32326,N_26749,N_28915);
and U32327 (N_32327,N_26697,N_28176);
and U32328 (N_32328,N_29463,N_26041);
and U32329 (N_32329,N_27936,N_28281);
nand U32330 (N_32330,N_26258,N_29813);
xor U32331 (N_32331,N_25839,N_29044);
or U32332 (N_32332,N_26468,N_29335);
xor U32333 (N_32333,N_28631,N_29621);
nand U32334 (N_32334,N_29338,N_28794);
nor U32335 (N_32335,N_26539,N_27227);
and U32336 (N_32336,N_29012,N_28411);
nand U32337 (N_32337,N_28617,N_27545);
xor U32338 (N_32338,N_29333,N_29061);
xor U32339 (N_32339,N_28905,N_29393);
and U32340 (N_32340,N_25480,N_29390);
nor U32341 (N_32341,N_25585,N_27962);
xor U32342 (N_32342,N_28621,N_27448);
nand U32343 (N_32343,N_26263,N_28790);
nand U32344 (N_32344,N_27285,N_26055);
or U32345 (N_32345,N_27153,N_28347);
xor U32346 (N_32346,N_26401,N_27387);
nor U32347 (N_32347,N_27903,N_25405);
nor U32348 (N_32348,N_25444,N_27759);
or U32349 (N_32349,N_26939,N_26104);
and U32350 (N_32350,N_25765,N_27528);
nor U32351 (N_32351,N_27752,N_27821);
nor U32352 (N_32352,N_28863,N_28690);
and U32353 (N_32353,N_27036,N_27480);
nand U32354 (N_32354,N_25736,N_27142);
xnor U32355 (N_32355,N_28031,N_26966);
nor U32356 (N_32356,N_29339,N_28003);
xor U32357 (N_32357,N_26964,N_27271);
nand U32358 (N_32358,N_26220,N_29443);
nor U32359 (N_32359,N_26944,N_27360);
nand U32360 (N_32360,N_26846,N_27460);
or U32361 (N_32361,N_29219,N_25881);
nand U32362 (N_32362,N_28193,N_26244);
and U32363 (N_32363,N_27700,N_25478);
nand U32364 (N_32364,N_27785,N_27155);
and U32365 (N_32365,N_28671,N_25001);
and U32366 (N_32366,N_29431,N_25623);
nor U32367 (N_32367,N_28841,N_29513);
and U32368 (N_32368,N_25087,N_27614);
xor U32369 (N_32369,N_29691,N_27113);
xor U32370 (N_32370,N_28784,N_27519);
xor U32371 (N_32371,N_28184,N_26431);
nand U32372 (N_32372,N_25440,N_29167);
nor U32373 (N_32373,N_29711,N_25678);
and U32374 (N_32374,N_29878,N_27694);
nand U32375 (N_32375,N_26261,N_27531);
and U32376 (N_32376,N_28713,N_28821);
nor U32377 (N_32377,N_29896,N_29268);
nor U32378 (N_32378,N_27451,N_25466);
nor U32379 (N_32379,N_28200,N_29544);
nand U32380 (N_32380,N_28383,N_25958);
nor U32381 (N_32381,N_26889,N_29854);
or U32382 (N_32382,N_27675,N_29927);
nand U32383 (N_32383,N_28997,N_27317);
nor U32384 (N_32384,N_28556,N_28495);
or U32385 (N_32385,N_26380,N_26440);
nor U32386 (N_32386,N_28344,N_25163);
xor U32387 (N_32387,N_27049,N_26025);
xor U32388 (N_32388,N_27596,N_29892);
nor U32389 (N_32389,N_29203,N_27578);
nor U32390 (N_32390,N_28351,N_25954);
and U32391 (N_32391,N_25515,N_27956);
nand U32392 (N_32392,N_26182,N_25548);
or U32393 (N_32393,N_26806,N_25028);
or U32394 (N_32394,N_26977,N_27442);
and U32395 (N_32395,N_27599,N_29017);
or U32396 (N_32396,N_25855,N_29046);
and U32397 (N_32397,N_27305,N_27524);
and U32398 (N_32398,N_29940,N_29087);
or U32399 (N_32399,N_28217,N_25587);
xnor U32400 (N_32400,N_26252,N_26937);
nor U32401 (N_32401,N_27119,N_29886);
nor U32402 (N_32402,N_27863,N_25569);
and U32403 (N_32403,N_28977,N_28999);
or U32404 (N_32404,N_29162,N_29101);
xnor U32405 (N_32405,N_26310,N_29576);
xnor U32406 (N_32406,N_28534,N_29816);
and U32407 (N_32407,N_29053,N_26234);
xnor U32408 (N_32408,N_26860,N_29199);
or U32409 (N_32409,N_27423,N_29096);
xnor U32410 (N_32410,N_26613,N_25266);
nand U32411 (N_32411,N_28722,N_26325);
and U32412 (N_32412,N_29079,N_26399);
and U32413 (N_32413,N_28424,N_25599);
xnor U32414 (N_32414,N_27527,N_29978);
nor U32415 (N_32415,N_25589,N_27601);
xnor U32416 (N_32416,N_26752,N_29180);
and U32417 (N_32417,N_29303,N_29976);
and U32418 (N_32418,N_29152,N_25595);
or U32419 (N_32419,N_29688,N_25806);
nor U32420 (N_32420,N_25507,N_27085);
xnor U32421 (N_32421,N_28116,N_29175);
xnor U32422 (N_32422,N_28904,N_28651);
or U32423 (N_32423,N_27147,N_29950);
xor U32424 (N_32424,N_28881,N_29634);
nand U32425 (N_32425,N_29401,N_28446);
and U32426 (N_32426,N_25259,N_27104);
nand U32427 (N_32427,N_26476,N_27212);
nand U32428 (N_32428,N_25749,N_27751);
nor U32429 (N_32429,N_26315,N_26583);
xor U32430 (N_32430,N_29446,N_27040);
xor U32431 (N_32431,N_26144,N_25012);
nor U32432 (N_32432,N_29018,N_28683);
and U32433 (N_32433,N_28381,N_26338);
nand U32434 (N_32434,N_28458,N_25482);
nor U32435 (N_32435,N_26472,N_27056);
xnor U32436 (N_32436,N_25842,N_26130);
or U32437 (N_32437,N_25511,N_28256);
xor U32438 (N_32438,N_26154,N_25232);
xor U32439 (N_32439,N_28558,N_27097);
and U32440 (N_32440,N_26492,N_26349);
and U32441 (N_32441,N_25038,N_28708);
nand U32442 (N_32442,N_28916,N_27658);
and U32443 (N_32443,N_27488,N_25519);
nor U32444 (N_32444,N_26723,N_25601);
nor U32445 (N_32445,N_26308,N_25486);
nand U32446 (N_32446,N_28567,N_28875);
and U32447 (N_32447,N_26344,N_25489);
xnor U32448 (N_32448,N_29803,N_28720);
and U32449 (N_32449,N_26197,N_29581);
or U32450 (N_32450,N_29552,N_29248);
xor U32451 (N_32451,N_28972,N_28765);
xnor U32452 (N_32452,N_28991,N_27934);
and U32453 (N_32453,N_28768,N_26925);
and U32454 (N_32454,N_28240,N_26770);
xnor U32455 (N_32455,N_26644,N_28440);
nand U32456 (N_32456,N_26211,N_27458);
and U32457 (N_32457,N_28542,N_28431);
nor U32458 (N_32458,N_27696,N_27687);
or U32459 (N_32459,N_28607,N_27349);
or U32460 (N_32460,N_28601,N_27240);
or U32461 (N_32461,N_28027,N_27430);
and U32462 (N_32462,N_29984,N_26500);
or U32463 (N_32463,N_26544,N_26080);
or U32464 (N_32464,N_26883,N_28699);
nand U32465 (N_32465,N_27767,N_29500);
xor U32466 (N_32466,N_27434,N_26420);
and U32467 (N_32467,N_27987,N_26659);
and U32468 (N_32468,N_27302,N_29850);
and U32469 (N_32469,N_29229,N_29005);
nor U32470 (N_32470,N_25075,N_28926);
nand U32471 (N_32471,N_29240,N_27798);
xor U32472 (N_32472,N_26410,N_25691);
or U32473 (N_32473,N_28348,N_29043);
nor U32474 (N_32474,N_28490,N_28173);
nand U32475 (N_32475,N_26240,N_26655);
xor U32476 (N_32476,N_29566,N_27320);
nor U32477 (N_32477,N_29720,N_26884);
nor U32478 (N_32478,N_29055,N_26617);
nand U32479 (N_32479,N_29661,N_26311);
xnor U32480 (N_32480,N_26982,N_28509);
or U32481 (N_32481,N_29784,N_27455);
and U32482 (N_32482,N_28829,N_29102);
and U32483 (N_32483,N_27971,N_27139);
or U32484 (N_32484,N_25928,N_27502);
or U32485 (N_32485,N_26961,N_28967);
xor U32486 (N_32486,N_28149,N_28185);
xor U32487 (N_32487,N_26535,N_26097);
nor U32488 (N_32488,N_26484,N_28797);
xor U32489 (N_32489,N_28945,N_27831);
xor U32490 (N_32490,N_29887,N_28305);
xor U32491 (N_32491,N_29760,N_27680);
xor U32492 (N_32492,N_29397,N_27336);
and U32493 (N_32493,N_29136,N_28210);
nand U32494 (N_32494,N_27960,N_26722);
xnor U32495 (N_32495,N_29695,N_28931);
or U32496 (N_32496,N_28216,N_28104);
nor U32497 (N_32497,N_29426,N_28403);
and U32498 (N_32498,N_28449,N_26413);
and U32499 (N_32499,N_25500,N_27994);
nand U32500 (N_32500,N_29472,N_25941);
nor U32501 (N_32501,N_29396,N_27362);
or U32502 (N_32502,N_26523,N_26962);
nand U32503 (N_32503,N_29713,N_27466);
xor U32504 (N_32504,N_26213,N_26185);
xnor U32505 (N_32505,N_25554,N_25830);
nor U32506 (N_32506,N_28900,N_26415);
nand U32507 (N_32507,N_26237,N_29350);
xnor U32508 (N_32508,N_25923,N_27567);
and U32509 (N_32509,N_25389,N_29975);
xor U32510 (N_32510,N_26202,N_29931);
or U32511 (N_32511,N_27324,N_27658);
nand U32512 (N_32512,N_26836,N_26445);
xor U32513 (N_32513,N_28287,N_26725);
nor U32514 (N_32514,N_28334,N_28875);
or U32515 (N_32515,N_26364,N_27630);
or U32516 (N_32516,N_25960,N_28183);
nand U32517 (N_32517,N_29126,N_26106);
or U32518 (N_32518,N_29588,N_25309);
xnor U32519 (N_32519,N_28345,N_27331);
or U32520 (N_32520,N_26559,N_26683);
xnor U32521 (N_32521,N_28295,N_29093);
nand U32522 (N_32522,N_28077,N_27417);
or U32523 (N_32523,N_26102,N_25931);
xor U32524 (N_32524,N_25537,N_26192);
or U32525 (N_32525,N_27458,N_27387);
and U32526 (N_32526,N_26009,N_27650);
or U32527 (N_32527,N_27264,N_26491);
xor U32528 (N_32528,N_27227,N_28362);
nand U32529 (N_32529,N_25089,N_27947);
and U32530 (N_32530,N_27663,N_28862);
nor U32531 (N_32531,N_29660,N_28389);
or U32532 (N_32532,N_29028,N_25950);
xor U32533 (N_32533,N_26403,N_28028);
or U32534 (N_32534,N_26402,N_25908);
or U32535 (N_32535,N_26827,N_29911);
or U32536 (N_32536,N_27534,N_29241);
nor U32537 (N_32537,N_25198,N_25411);
and U32538 (N_32538,N_27203,N_28671);
nand U32539 (N_32539,N_28622,N_26829);
and U32540 (N_32540,N_28609,N_25293);
and U32541 (N_32541,N_26142,N_29717);
xor U32542 (N_32542,N_27378,N_26140);
and U32543 (N_32543,N_26326,N_29375);
or U32544 (N_32544,N_28463,N_26541);
and U32545 (N_32545,N_27373,N_29610);
and U32546 (N_32546,N_28989,N_25310);
nor U32547 (N_32547,N_28991,N_29111);
nor U32548 (N_32548,N_28150,N_28702);
and U32549 (N_32549,N_28805,N_29864);
xnor U32550 (N_32550,N_28475,N_27275);
nand U32551 (N_32551,N_28820,N_28849);
or U32552 (N_32552,N_26897,N_28228);
nor U32553 (N_32553,N_27597,N_25711);
and U32554 (N_32554,N_27566,N_28747);
and U32555 (N_32555,N_29799,N_29636);
nand U32556 (N_32556,N_27138,N_29363);
and U32557 (N_32557,N_26872,N_27445);
or U32558 (N_32558,N_25388,N_27702);
or U32559 (N_32559,N_27383,N_27654);
xor U32560 (N_32560,N_25437,N_28552);
or U32561 (N_32561,N_26864,N_26541);
and U32562 (N_32562,N_27714,N_27308);
nand U32563 (N_32563,N_25451,N_26040);
nor U32564 (N_32564,N_26756,N_28571);
xor U32565 (N_32565,N_25502,N_28691);
and U32566 (N_32566,N_27286,N_25605);
nand U32567 (N_32567,N_27901,N_26662);
nand U32568 (N_32568,N_29601,N_25942);
nand U32569 (N_32569,N_26940,N_28253);
xor U32570 (N_32570,N_29616,N_27025);
xnor U32571 (N_32571,N_27925,N_26647);
or U32572 (N_32572,N_29310,N_28730);
xnor U32573 (N_32573,N_25066,N_28884);
xor U32574 (N_32574,N_26571,N_26584);
nand U32575 (N_32575,N_29784,N_29255);
and U32576 (N_32576,N_29693,N_29362);
nand U32577 (N_32577,N_28725,N_28534);
xnor U32578 (N_32578,N_27209,N_26851);
and U32579 (N_32579,N_25467,N_25607);
and U32580 (N_32580,N_28705,N_27290);
nor U32581 (N_32581,N_25128,N_27037);
nor U32582 (N_32582,N_25124,N_29564);
and U32583 (N_32583,N_26543,N_28662);
xor U32584 (N_32584,N_26905,N_29711);
and U32585 (N_32585,N_26741,N_29000);
xor U32586 (N_32586,N_28395,N_25463);
or U32587 (N_32587,N_28395,N_26792);
and U32588 (N_32588,N_26255,N_28443);
xor U32589 (N_32589,N_25405,N_26608);
nand U32590 (N_32590,N_29110,N_28744);
and U32591 (N_32591,N_27659,N_28277);
nor U32592 (N_32592,N_27267,N_27608);
xnor U32593 (N_32593,N_26763,N_28795);
or U32594 (N_32594,N_29606,N_27604);
nor U32595 (N_32595,N_26380,N_26949);
xnor U32596 (N_32596,N_29726,N_26594);
and U32597 (N_32597,N_26547,N_29742);
and U32598 (N_32598,N_29646,N_28423);
and U32599 (N_32599,N_27941,N_26693);
and U32600 (N_32600,N_27439,N_26345);
and U32601 (N_32601,N_26950,N_27244);
and U32602 (N_32602,N_25123,N_27470);
nor U32603 (N_32603,N_29279,N_26156);
xnor U32604 (N_32604,N_28006,N_25345);
or U32605 (N_32605,N_29159,N_25365);
nand U32606 (N_32606,N_25493,N_26245);
and U32607 (N_32607,N_27013,N_25891);
nand U32608 (N_32608,N_27322,N_28713);
and U32609 (N_32609,N_25927,N_29189);
nand U32610 (N_32610,N_27602,N_29469);
nor U32611 (N_32611,N_28611,N_28069);
nor U32612 (N_32612,N_25808,N_28594);
nand U32613 (N_32613,N_26890,N_25450);
xnor U32614 (N_32614,N_29452,N_28635);
and U32615 (N_32615,N_28051,N_27881);
and U32616 (N_32616,N_25323,N_27011);
nand U32617 (N_32617,N_26828,N_26171);
nand U32618 (N_32618,N_25710,N_25911);
nor U32619 (N_32619,N_28601,N_27456);
xnor U32620 (N_32620,N_25235,N_26768);
nor U32621 (N_32621,N_29033,N_28490);
nor U32622 (N_32622,N_29166,N_26824);
nor U32623 (N_32623,N_26165,N_29466);
or U32624 (N_32624,N_27215,N_27845);
xor U32625 (N_32625,N_26499,N_25592);
xnor U32626 (N_32626,N_25239,N_27818);
nor U32627 (N_32627,N_26602,N_27194);
nand U32628 (N_32628,N_25334,N_29366);
nand U32629 (N_32629,N_28989,N_25299);
and U32630 (N_32630,N_27659,N_29772);
nand U32631 (N_32631,N_27384,N_26475);
nand U32632 (N_32632,N_26367,N_28147);
nand U32633 (N_32633,N_29884,N_27757);
nand U32634 (N_32634,N_27557,N_28555);
or U32635 (N_32635,N_29916,N_25822);
or U32636 (N_32636,N_25049,N_25595);
nor U32637 (N_32637,N_27258,N_29738);
and U32638 (N_32638,N_27663,N_26180);
nor U32639 (N_32639,N_29861,N_26158);
nor U32640 (N_32640,N_27772,N_28381);
nand U32641 (N_32641,N_25660,N_26009);
and U32642 (N_32642,N_26371,N_27458);
nand U32643 (N_32643,N_27157,N_25206);
and U32644 (N_32644,N_25878,N_25360);
and U32645 (N_32645,N_26704,N_27686);
or U32646 (N_32646,N_25363,N_25941);
xor U32647 (N_32647,N_26848,N_28507);
and U32648 (N_32648,N_29338,N_28023);
and U32649 (N_32649,N_25349,N_27499);
nor U32650 (N_32650,N_25159,N_28839);
and U32651 (N_32651,N_27360,N_25079);
or U32652 (N_32652,N_28908,N_25654);
or U32653 (N_32653,N_25265,N_28113);
nand U32654 (N_32654,N_25983,N_27063);
xnor U32655 (N_32655,N_27509,N_25706);
nor U32656 (N_32656,N_29743,N_25158);
and U32657 (N_32657,N_26190,N_28117);
nand U32658 (N_32658,N_25709,N_25629);
xor U32659 (N_32659,N_25227,N_29998);
or U32660 (N_32660,N_25889,N_28470);
nand U32661 (N_32661,N_25318,N_29651);
and U32662 (N_32662,N_26736,N_25445);
or U32663 (N_32663,N_26374,N_27690);
and U32664 (N_32664,N_25498,N_25998);
nor U32665 (N_32665,N_29602,N_26754);
xor U32666 (N_32666,N_25096,N_27890);
xor U32667 (N_32667,N_28361,N_27453);
xnor U32668 (N_32668,N_28022,N_25017);
nand U32669 (N_32669,N_25690,N_28802);
and U32670 (N_32670,N_26424,N_25448);
xor U32671 (N_32671,N_27746,N_25562);
xnor U32672 (N_32672,N_25079,N_27259);
nand U32673 (N_32673,N_28471,N_26032);
and U32674 (N_32674,N_25552,N_25930);
nand U32675 (N_32675,N_26099,N_29124);
or U32676 (N_32676,N_27451,N_25409);
and U32677 (N_32677,N_29575,N_29554);
nor U32678 (N_32678,N_27159,N_27930);
or U32679 (N_32679,N_28029,N_25785);
and U32680 (N_32680,N_25756,N_26189);
or U32681 (N_32681,N_27287,N_25030);
and U32682 (N_32682,N_25155,N_29296);
or U32683 (N_32683,N_26890,N_26668);
nor U32684 (N_32684,N_28145,N_26182);
or U32685 (N_32685,N_28718,N_29102);
xnor U32686 (N_32686,N_27908,N_26878);
nand U32687 (N_32687,N_26362,N_27136);
nor U32688 (N_32688,N_26067,N_28532);
nor U32689 (N_32689,N_26236,N_29900);
or U32690 (N_32690,N_26922,N_26299);
nand U32691 (N_32691,N_29990,N_28589);
nor U32692 (N_32692,N_29869,N_28597);
or U32693 (N_32693,N_26923,N_26862);
or U32694 (N_32694,N_28745,N_29923);
nand U32695 (N_32695,N_26612,N_29934);
nor U32696 (N_32696,N_28535,N_28143);
nor U32697 (N_32697,N_28317,N_25278);
xnor U32698 (N_32698,N_28972,N_29156);
and U32699 (N_32699,N_27781,N_26668);
nand U32700 (N_32700,N_27508,N_25125);
xor U32701 (N_32701,N_25224,N_28930);
nand U32702 (N_32702,N_26449,N_25116);
xor U32703 (N_32703,N_28130,N_29091);
or U32704 (N_32704,N_27224,N_27980);
xor U32705 (N_32705,N_28279,N_26296);
nor U32706 (N_32706,N_25670,N_26979);
or U32707 (N_32707,N_27954,N_25037);
and U32708 (N_32708,N_27569,N_28543);
xnor U32709 (N_32709,N_27963,N_28271);
nor U32710 (N_32710,N_28941,N_26692);
or U32711 (N_32711,N_25231,N_29866);
nor U32712 (N_32712,N_28976,N_29850);
or U32713 (N_32713,N_26302,N_25156);
or U32714 (N_32714,N_26692,N_26880);
nand U32715 (N_32715,N_29436,N_28994);
xor U32716 (N_32716,N_29603,N_27314);
and U32717 (N_32717,N_25308,N_26465);
or U32718 (N_32718,N_26133,N_27959);
nand U32719 (N_32719,N_28821,N_26531);
nor U32720 (N_32720,N_28903,N_27586);
nor U32721 (N_32721,N_28239,N_25680);
nor U32722 (N_32722,N_25605,N_27929);
or U32723 (N_32723,N_28532,N_25071);
nor U32724 (N_32724,N_27126,N_25550);
nand U32725 (N_32725,N_27238,N_26776);
nand U32726 (N_32726,N_28849,N_26900);
or U32727 (N_32727,N_28139,N_25929);
and U32728 (N_32728,N_25930,N_29512);
and U32729 (N_32729,N_25640,N_27097);
nor U32730 (N_32730,N_29095,N_26561);
and U32731 (N_32731,N_26532,N_29689);
nand U32732 (N_32732,N_28743,N_28559);
nand U32733 (N_32733,N_25875,N_27192);
nor U32734 (N_32734,N_27649,N_25734);
and U32735 (N_32735,N_28342,N_28147);
xor U32736 (N_32736,N_29081,N_27073);
or U32737 (N_32737,N_27486,N_29039);
or U32738 (N_32738,N_25389,N_27157);
and U32739 (N_32739,N_26900,N_27102);
nor U32740 (N_32740,N_29784,N_29706);
xnor U32741 (N_32741,N_29272,N_29635);
xnor U32742 (N_32742,N_27575,N_29615);
xnor U32743 (N_32743,N_27036,N_29396);
or U32744 (N_32744,N_25032,N_25390);
and U32745 (N_32745,N_29312,N_26304);
and U32746 (N_32746,N_25088,N_27443);
xnor U32747 (N_32747,N_29873,N_27769);
xnor U32748 (N_32748,N_29578,N_28083);
or U32749 (N_32749,N_27378,N_28432);
or U32750 (N_32750,N_27481,N_26746);
xnor U32751 (N_32751,N_29616,N_27635);
nand U32752 (N_32752,N_25943,N_25613);
xnor U32753 (N_32753,N_26066,N_28344);
xnor U32754 (N_32754,N_25517,N_28279);
nand U32755 (N_32755,N_28048,N_29663);
nand U32756 (N_32756,N_25736,N_28834);
xnor U32757 (N_32757,N_26582,N_28062);
nand U32758 (N_32758,N_27068,N_28777);
or U32759 (N_32759,N_28070,N_27912);
xor U32760 (N_32760,N_27430,N_25164);
nor U32761 (N_32761,N_27339,N_29539);
nand U32762 (N_32762,N_29999,N_25790);
nor U32763 (N_32763,N_29885,N_28873);
nand U32764 (N_32764,N_29494,N_26727);
or U32765 (N_32765,N_25318,N_28023);
nor U32766 (N_32766,N_25867,N_26799);
xor U32767 (N_32767,N_25886,N_25503);
and U32768 (N_32768,N_26701,N_28455);
xor U32769 (N_32769,N_27860,N_29347);
xor U32770 (N_32770,N_27683,N_29352);
and U32771 (N_32771,N_28999,N_28328);
nor U32772 (N_32772,N_25028,N_29206);
nand U32773 (N_32773,N_28641,N_26280);
nand U32774 (N_32774,N_26348,N_26309);
and U32775 (N_32775,N_28042,N_28716);
or U32776 (N_32776,N_25003,N_25912);
or U32777 (N_32777,N_27618,N_26619);
xor U32778 (N_32778,N_26512,N_27175);
xnor U32779 (N_32779,N_26909,N_25017);
xnor U32780 (N_32780,N_29357,N_25534);
or U32781 (N_32781,N_29795,N_26630);
or U32782 (N_32782,N_27260,N_28347);
nor U32783 (N_32783,N_27172,N_27818);
nand U32784 (N_32784,N_28764,N_28198);
or U32785 (N_32785,N_26543,N_25755);
or U32786 (N_32786,N_28740,N_29479);
and U32787 (N_32787,N_26218,N_29898);
xnor U32788 (N_32788,N_25628,N_27252);
nor U32789 (N_32789,N_29558,N_25299);
or U32790 (N_32790,N_29129,N_25019);
or U32791 (N_32791,N_27873,N_28858);
nor U32792 (N_32792,N_28089,N_26235);
xor U32793 (N_32793,N_28929,N_28412);
nor U32794 (N_32794,N_27490,N_26798);
or U32795 (N_32795,N_25420,N_25526);
and U32796 (N_32796,N_26730,N_29719);
xor U32797 (N_32797,N_25482,N_26151);
and U32798 (N_32798,N_28744,N_25162);
xnor U32799 (N_32799,N_25869,N_25423);
or U32800 (N_32800,N_27631,N_29795);
xor U32801 (N_32801,N_29102,N_29291);
nor U32802 (N_32802,N_27608,N_25059);
xnor U32803 (N_32803,N_29784,N_25035);
xnor U32804 (N_32804,N_28685,N_28815);
nor U32805 (N_32805,N_27428,N_26598);
and U32806 (N_32806,N_28046,N_29931);
nor U32807 (N_32807,N_27976,N_26847);
and U32808 (N_32808,N_29286,N_29722);
or U32809 (N_32809,N_25220,N_28369);
or U32810 (N_32810,N_28529,N_27853);
or U32811 (N_32811,N_27410,N_26331);
xnor U32812 (N_32812,N_28729,N_25518);
nor U32813 (N_32813,N_28936,N_25091);
xor U32814 (N_32814,N_27773,N_25447);
nand U32815 (N_32815,N_26942,N_28084);
xor U32816 (N_32816,N_29606,N_27401);
nor U32817 (N_32817,N_28366,N_27923);
or U32818 (N_32818,N_27210,N_25109);
nand U32819 (N_32819,N_26511,N_29139);
nor U32820 (N_32820,N_26283,N_26040);
nor U32821 (N_32821,N_26536,N_26157);
nor U32822 (N_32822,N_29608,N_27469);
xnor U32823 (N_32823,N_27970,N_25704);
or U32824 (N_32824,N_25110,N_27771);
and U32825 (N_32825,N_27962,N_25191);
nor U32826 (N_32826,N_26960,N_26377);
xor U32827 (N_32827,N_29231,N_25542);
nand U32828 (N_32828,N_26550,N_28538);
nor U32829 (N_32829,N_26358,N_25455);
nor U32830 (N_32830,N_28132,N_28782);
nor U32831 (N_32831,N_29282,N_25222);
xnor U32832 (N_32832,N_27169,N_27562);
xnor U32833 (N_32833,N_29738,N_29763);
nor U32834 (N_32834,N_25125,N_27601);
and U32835 (N_32835,N_25626,N_29807);
xor U32836 (N_32836,N_26639,N_26699);
or U32837 (N_32837,N_29698,N_27553);
xor U32838 (N_32838,N_28769,N_25566);
nor U32839 (N_32839,N_26967,N_25502);
or U32840 (N_32840,N_27089,N_25486);
nand U32841 (N_32841,N_25398,N_27676);
or U32842 (N_32842,N_29894,N_28330);
xor U32843 (N_32843,N_27349,N_28687);
nor U32844 (N_32844,N_27526,N_27167);
xor U32845 (N_32845,N_29176,N_27678);
nor U32846 (N_32846,N_28754,N_25299);
or U32847 (N_32847,N_27800,N_25521);
nand U32848 (N_32848,N_26278,N_28081);
or U32849 (N_32849,N_29682,N_25212);
nor U32850 (N_32850,N_25759,N_27350);
and U32851 (N_32851,N_27760,N_27485);
and U32852 (N_32852,N_27505,N_29541);
nor U32853 (N_32853,N_29111,N_26198);
xor U32854 (N_32854,N_27191,N_27702);
xor U32855 (N_32855,N_26407,N_25922);
or U32856 (N_32856,N_26346,N_26246);
and U32857 (N_32857,N_25739,N_29797);
and U32858 (N_32858,N_28866,N_28120);
nor U32859 (N_32859,N_28875,N_29927);
nand U32860 (N_32860,N_28059,N_26494);
nor U32861 (N_32861,N_28742,N_29225);
or U32862 (N_32862,N_28987,N_28936);
or U32863 (N_32863,N_29558,N_28454);
and U32864 (N_32864,N_28280,N_28402);
nand U32865 (N_32865,N_27105,N_26806);
nor U32866 (N_32866,N_27970,N_29923);
nand U32867 (N_32867,N_27596,N_25023);
xor U32868 (N_32868,N_27157,N_27492);
xor U32869 (N_32869,N_25005,N_28459);
and U32870 (N_32870,N_25081,N_29295);
nand U32871 (N_32871,N_29905,N_27671);
and U32872 (N_32872,N_26916,N_25180);
and U32873 (N_32873,N_25989,N_25286);
xor U32874 (N_32874,N_29685,N_28610);
nand U32875 (N_32875,N_25670,N_27733);
nor U32876 (N_32876,N_25655,N_27958);
nand U32877 (N_32877,N_28816,N_27189);
and U32878 (N_32878,N_25527,N_27880);
nand U32879 (N_32879,N_26049,N_29722);
and U32880 (N_32880,N_26302,N_27215);
or U32881 (N_32881,N_28094,N_26336);
nand U32882 (N_32882,N_29873,N_27778);
and U32883 (N_32883,N_26038,N_26937);
and U32884 (N_32884,N_28426,N_25884);
and U32885 (N_32885,N_29224,N_25545);
nand U32886 (N_32886,N_29238,N_25941);
nor U32887 (N_32887,N_26974,N_25677);
nand U32888 (N_32888,N_29087,N_27551);
or U32889 (N_32889,N_25451,N_26402);
and U32890 (N_32890,N_28595,N_28437);
and U32891 (N_32891,N_29453,N_25385);
nand U32892 (N_32892,N_27586,N_28836);
xor U32893 (N_32893,N_28645,N_25563);
nand U32894 (N_32894,N_26112,N_28564);
and U32895 (N_32895,N_29736,N_28111);
or U32896 (N_32896,N_25396,N_25390);
and U32897 (N_32897,N_28302,N_25989);
nor U32898 (N_32898,N_25240,N_29178);
xor U32899 (N_32899,N_27182,N_28638);
or U32900 (N_32900,N_28853,N_29060);
nand U32901 (N_32901,N_26644,N_27946);
nor U32902 (N_32902,N_27893,N_28448);
nor U32903 (N_32903,N_28747,N_27862);
or U32904 (N_32904,N_27041,N_26071);
and U32905 (N_32905,N_26150,N_27258);
and U32906 (N_32906,N_25020,N_25796);
nor U32907 (N_32907,N_25169,N_28633);
and U32908 (N_32908,N_26473,N_29425);
nand U32909 (N_32909,N_25212,N_27026);
and U32910 (N_32910,N_29190,N_28991);
or U32911 (N_32911,N_29043,N_28330);
nor U32912 (N_32912,N_26582,N_27343);
nand U32913 (N_32913,N_28929,N_27417);
nor U32914 (N_32914,N_27424,N_29968);
nor U32915 (N_32915,N_26039,N_28278);
nand U32916 (N_32916,N_27954,N_25801);
and U32917 (N_32917,N_25707,N_28679);
nor U32918 (N_32918,N_26589,N_26790);
xnor U32919 (N_32919,N_26630,N_27938);
and U32920 (N_32920,N_27998,N_28772);
or U32921 (N_32921,N_28349,N_25238);
xnor U32922 (N_32922,N_28176,N_27094);
nor U32923 (N_32923,N_26664,N_28720);
xor U32924 (N_32924,N_26181,N_26222);
xnor U32925 (N_32925,N_27026,N_27238);
xor U32926 (N_32926,N_25143,N_29386);
or U32927 (N_32927,N_28351,N_26310);
nor U32928 (N_32928,N_25863,N_28515);
nor U32929 (N_32929,N_29322,N_28960);
xor U32930 (N_32930,N_27215,N_25424);
nand U32931 (N_32931,N_25741,N_26754);
nor U32932 (N_32932,N_25506,N_25913);
or U32933 (N_32933,N_28407,N_27363);
nor U32934 (N_32934,N_28090,N_27758);
nand U32935 (N_32935,N_25931,N_27254);
nand U32936 (N_32936,N_26641,N_29584);
xnor U32937 (N_32937,N_29565,N_25027);
nor U32938 (N_32938,N_29043,N_29959);
or U32939 (N_32939,N_25492,N_29356);
or U32940 (N_32940,N_29259,N_25503);
xnor U32941 (N_32941,N_25971,N_29288);
nand U32942 (N_32942,N_27498,N_25867);
xor U32943 (N_32943,N_25009,N_26619);
or U32944 (N_32944,N_28960,N_26650);
xnor U32945 (N_32945,N_29959,N_26000);
nand U32946 (N_32946,N_28315,N_26112);
or U32947 (N_32947,N_26358,N_27203);
or U32948 (N_32948,N_28949,N_29560);
xor U32949 (N_32949,N_29375,N_25590);
xnor U32950 (N_32950,N_29195,N_29160);
xnor U32951 (N_32951,N_28697,N_29325);
and U32952 (N_32952,N_26138,N_27413);
or U32953 (N_32953,N_27417,N_26267);
or U32954 (N_32954,N_29352,N_28451);
xnor U32955 (N_32955,N_27333,N_25993);
nor U32956 (N_32956,N_28224,N_25809);
nand U32957 (N_32957,N_26283,N_26108);
xnor U32958 (N_32958,N_26175,N_29093);
and U32959 (N_32959,N_28130,N_27858);
nand U32960 (N_32960,N_29242,N_26014);
or U32961 (N_32961,N_26652,N_27425);
xor U32962 (N_32962,N_28861,N_25830);
and U32963 (N_32963,N_29000,N_29389);
nand U32964 (N_32964,N_26172,N_26847);
xor U32965 (N_32965,N_28630,N_25321);
xor U32966 (N_32966,N_27832,N_29572);
nor U32967 (N_32967,N_26647,N_26686);
nand U32968 (N_32968,N_26125,N_28503);
nand U32969 (N_32969,N_27662,N_26454);
and U32970 (N_32970,N_28866,N_29374);
or U32971 (N_32971,N_25382,N_25621);
nor U32972 (N_32972,N_28237,N_27706);
nor U32973 (N_32973,N_28581,N_25271);
xor U32974 (N_32974,N_28721,N_26857);
or U32975 (N_32975,N_27689,N_26026);
nand U32976 (N_32976,N_26389,N_26714);
xor U32977 (N_32977,N_26961,N_28984);
nor U32978 (N_32978,N_26404,N_29120);
nand U32979 (N_32979,N_27248,N_25782);
or U32980 (N_32980,N_25880,N_26894);
and U32981 (N_32981,N_25809,N_26097);
nor U32982 (N_32982,N_28336,N_27213);
or U32983 (N_32983,N_26896,N_25085);
xor U32984 (N_32984,N_27794,N_27341);
xnor U32985 (N_32985,N_29554,N_25129);
nand U32986 (N_32986,N_28880,N_29360);
xnor U32987 (N_32987,N_29613,N_26752);
or U32988 (N_32988,N_26796,N_25053);
xor U32989 (N_32989,N_27868,N_27160);
nand U32990 (N_32990,N_27206,N_27575);
nor U32991 (N_32991,N_28634,N_28620);
or U32992 (N_32992,N_26828,N_29364);
or U32993 (N_32993,N_25010,N_27140);
nand U32994 (N_32994,N_27140,N_26913);
nor U32995 (N_32995,N_26413,N_25283);
or U32996 (N_32996,N_28983,N_28922);
and U32997 (N_32997,N_27206,N_29055);
nor U32998 (N_32998,N_27858,N_29859);
nor U32999 (N_32999,N_25485,N_25958);
and U33000 (N_33000,N_26244,N_28910);
nor U33001 (N_33001,N_28291,N_26207);
xor U33002 (N_33002,N_28191,N_29449);
or U33003 (N_33003,N_26179,N_27353);
xor U33004 (N_33004,N_28911,N_25654);
and U33005 (N_33005,N_28585,N_27356);
and U33006 (N_33006,N_28664,N_28672);
or U33007 (N_33007,N_27001,N_26500);
and U33008 (N_33008,N_26300,N_27232);
xnor U33009 (N_33009,N_26927,N_29729);
or U33010 (N_33010,N_29823,N_26699);
xnor U33011 (N_33011,N_27672,N_29151);
nor U33012 (N_33012,N_27117,N_27488);
nor U33013 (N_33013,N_29449,N_25664);
xnor U33014 (N_33014,N_26196,N_27382);
xor U33015 (N_33015,N_29648,N_28967);
nor U33016 (N_33016,N_27527,N_29133);
or U33017 (N_33017,N_29196,N_28380);
xor U33018 (N_33018,N_28422,N_27960);
or U33019 (N_33019,N_28949,N_29905);
and U33020 (N_33020,N_28021,N_26710);
nor U33021 (N_33021,N_29560,N_25224);
xnor U33022 (N_33022,N_28412,N_26460);
and U33023 (N_33023,N_26734,N_27405);
nand U33024 (N_33024,N_29148,N_28987);
nor U33025 (N_33025,N_27674,N_25164);
nor U33026 (N_33026,N_28627,N_27837);
or U33027 (N_33027,N_29005,N_29441);
xnor U33028 (N_33028,N_26982,N_27315);
and U33029 (N_33029,N_26086,N_25889);
nor U33030 (N_33030,N_29379,N_25258);
or U33031 (N_33031,N_29615,N_27100);
nand U33032 (N_33032,N_25433,N_28303);
nor U33033 (N_33033,N_25622,N_27432);
nor U33034 (N_33034,N_29170,N_26993);
or U33035 (N_33035,N_26021,N_29586);
nand U33036 (N_33036,N_27457,N_28917);
and U33037 (N_33037,N_29102,N_26820);
xor U33038 (N_33038,N_27315,N_28793);
or U33039 (N_33039,N_26691,N_25898);
nor U33040 (N_33040,N_26520,N_26470);
xnor U33041 (N_33041,N_29662,N_28709);
xor U33042 (N_33042,N_29009,N_25999);
and U33043 (N_33043,N_25880,N_28954);
nand U33044 (N_33044,N_25679,N_27775);
and U33045 (N_33045,N_26402,N_28594);
or U33046 (N_33046,N_29695,N_26305);
xor U33047 (N_33047,N_25593,N_28085);
or U33048 (N_33048,N_29398,N_26759);
nor U33049 (N_33049,N_28449,N_28107);
xor U33050 (N_33050,N_27533,N_28954);
and U33051 (N_33051,N_25901,N_26158);
nand U33052 (N_33052,N_26203,N_29555);
nor U33053 (N_33053,N_28748,N_26932);
and U33054 (N_33054,N_28780,N_28931);
or U33055 (N_33055,N_28470,N_28052);
or U33056 (N_33056,N_27988,N_25939);
xnor U33057 (N_33057,N_27457,N_27245);
xor U33058 (N_33058,N_28121,N_28806);
nor U33059 (N_33059,N_29458,N_25050);
or U33060 (N_33060,N_28848,N_25990);
and U33061 (N_33061,N_29523,N_27708);
nand U33062 (N_33062,N_29634,N_25961);
nor U33063 (N_33063,N_27726,N_25796);
or U33064 (N_33064,N_29960,N_25346);
nor U33065 (N_33065,N_29678,N_25869);
or U33066 (N_33066,N_27273,N_26194);
nor U33067 (N_33067,N_27603,N_29883);
or U33068 (N_33068,N_27003,N_26612);
nand U33069 (N_33069,N_27523,N_27945);
nor U33070 (N_33070,N_26900,N_27076);
and U33071 (N_33071,N_25011,N_27840);
xnor U33072 (N_33072,N_28496,N_26717);
and U33073 (N_33073,N_27392,N_26278);
xnor U33074 (N_33074,N_29135,N_28027);
xor U33075 (N_33075,N_28618,N_29886);
and U33076 (N_33076,N_26039,N_28358);
xnor U33077 (N_33077,N_28244,N_29906);
nor U33078 (N_33078,N_26374,N_27808);
or U33079 (N_33079,N_29946,N_29845);
or U33080 (N_33080,N_29569,N_29046);
xnor U33081 (N_33081,N_26219,N_28784);
nor U33082 (N_33082,N_29463,N_27494);
nor U33083 (N_33083,N_29210,N_29066);
xnor U33084 (N_33084,N_26071,N_27408);
nand U33085 (N_33085,N_26522,N_29693);
nand U33086 (N_33086,N_28944,N_27820);
and U33087 (N_33087,N_25373,N_27619);
nor U33088 (N_33088,N_29848,N_26769);
nor U33089 (N_33089,N_28151,N_26779);
nor U33090 (N_33090,N_27638,N_27636);
xor U33091 (N_33091,N_25874,N_28220);
nand U33092 (N_33092,N_27429,N_27356);
xor U33093 (N_33093,N_27750,N_27211);
nand U33094 (N_33094,N_29716,N_28919);
and U33095 (N_33095,N_26717,N_25146);
nor U33096 (N_33096,N_26048,N_26143);
nand U33097 (N_33097,N_28075,N_26620);
nand U33098 (N_33098,N_25636,N_27976);
nor U33099 (N_33099,N_29763,N_26837);
xor U33100 (N_33100,N_28182,N_29199);
nand U33101 (N_33101,N_27767,N_27682);
nand U33102 (N_33102,N_28320,N_26078);
nand U33103 (N_33103,N_27445,N_27683);
or U33104 (N_33104,N_28144,N_29848);
nor U33105 (N_33105,N_25292,N_26396);
nand U33106 (N_33106,N_29620,N_25134);
nand U33107 (N_33107,N_28176,N_29857);
nor U33108 (N_33108,N_29005,N_25341);
nand U33109 (N_33109,N_27850,N_28315);
xor U33110 (N_33110,N_28564,N_29200);
xnor U33111 (N_33111,N_29425,N_25853);
nor U33112 (N_33112,N_28577,N_27172);
nand U33113 (N_33113,N_27994,N_26936);
xnor U33114 (N_33114,N_27618,N_27152);
nor U33115 (N_33115,N_25016,N_29043);
nand U33116 (N_33116,N_25763,N_27300);
and U33117 (N_33117,N_27117,N_25631);
xor U33118 (N_33118,N_28017,N_26918);
nand U33119 (N_33119,N_27105,N_29603);
or U33120 (N_33120,N_28533,N_26261);
or U33121 (N_33121,N_28763,N_27479);
xor U33122 (N_33122,N_27257,N_29297);
nand U33123 (N_33123,N_28744,N_25994);
nand U33124 (N_33124,N_29529,N_25937);
nand U33125 (N_33125,N_27060,N_28714);
xor U33126 (N_33126,N_27719,N_27492);
or U33127 (N_33127,N_27096,N_29456);
nor U33128 (N_33128,N_28544,N_27118);
and U33129 (N_33129,N_27468,N_28219);
or U33130 (N_33130,N_26149,N_29205);
and U33131 (N_33131,N_26486,N_27207);
and U33132 (N_33132,N_25644,N_29743);
and U33133 (N_33133,N_28848,N_25205);
and U33134 (N_33134,N_28167,N_27945);
and U33135 (N_33135,N_29452,N_29684);
xnor U33136 (N_33136,N_29381,N_29996);
nand U33137 (N_33137,N_27228,N_28938);
nor U33138 (N_33138,N_29088,N_26777);
and U33139 (N_33139,N_28947,N_27193);
nand U33140 (N_33140,N_29377,N_28829);
nand U33141 (N_33141,N_27923,N_27645);
or U33142 (N_33142,N_28850,N_27134);
nor U33143 (N_33143,N_27154,N_28538);
or U33144 (N_33144,N_25021,N_29533);
or U33145 (N_33145,N_25960,N_27621);
nand U33146 (N_33146,N_25234,N_28493);
nand U33147 (N_33147,N_28327,N_25621);
nor U33148 (N_33148,N_27170,N_29328);
nor U33149 (N_33149,N_28848,N_28302);
nand U33150 (N_33150,N_25059,N_28771);
nand U33151 (N_33151,N_27687,N_29827);
nand U33152 (N_33152,N_26673,N_26520);
and U33153 (N_33153,N_26227,N_29614);
and U33154 (N_33154,N_25454,N_29439);
nor U33155 (N_33155,N_29750,N_29302);
nand U33156 (N_33156,N_29803,N_28326);
xnor U33157 (N_33157,N_28613,N_25703);
and U33158 (N_33158,N_28400,N_29051);
and U33159 (N_33159,N_27465,N_28584);
and U33160 (N_33160,N_29846,N_28416);
nand U33161 (N_33161,N_25533,N_25526);
nor U33162 (N_33162,N_27227,N_28168);
and U33163 (N_33163,N_26566,N_28039);
or U33164 (N_33164,N_29033,N_26736);
and U33165 (N_33165,N_25663,N_26423);
xnor U33166 (N_33166,N_25029,N_26933);
xor U33167 (N_33167,N_26855,N_26478);
nor U33168 (N_33168,N_29117,N_25838);
nand U33169 (N_33169,N_28735,N_26259);
nor U33170 (N_33170,N_28133,N_28627);
and U33171 (N_33171,N_27065,N_29278);
and U33172 (N_33172,N_28447,N_26715);
nor U33173 (N_33173,N_28706,N_28545);
nor U33174 (N_33174,N_28064,N_29387);
nand U33175 (N_33175,N_26415,N_26308);
nor U33176 (N_33176,N_26867,N_28364);
xnor U33177 (N_33177,N_26088,N_28715);
nand U33178 (N_33178,N_25916,N_29231);
or U33179 (N_33179,N_29434,N_25387);
or U33180 (N_33180,N_28304,N_25876);
and U33181 (N_33181,N_28742,N_28769);
nor U33182 (N_33182,N_29346,N_25342);
xnor U33183 (N_33183,N_29720,N_28714);
and U33184 (N_33184,N_26480,N_26420);
and U33185 (N_33185,N_27823,N_26617);
or U33186 (N_33186,N_29114,N_26402);
nor U33187 (N_33187,N_25719,N_29160);
nand U33188 (N_33188,N_29347,N_29716);
and U33189 (N_33189,N_25721,N_28183);
nor U33190 (N_33190,N_28984,N_25067);
xnor U33191 (N_33191,N_26225,N_27097);
or U33192 (N_33192,N_28814,N_28991);
and U33193 (N_33193,N_26590,N_28353);
or U33194 (N_33194,N_27391,N_25020);
and U33195 (N_33195,N_28820,N_29278);
nor U33196 (N_33196,N_26017,N_29298);
nand U33197 (N_33197,N_25702,N_26220);
nand U33198 (N_33198,N_25350,N_27501);
or U33199 (N_33199,N_25343,N_27253);
nand U33200 (N_33200,N_25881,N_29901);
or U33201 (N_33201,N_25963,N_28896);
xnor U33202 (N_33202,N_26206,N_27224);
nand U33203 (N_33203,N_25391,N_25997);
and U33204 (N_33204,N_27353,N_27100);
or U33205 (N_33205,N_27324,N_25120);
nand U33206 (N_33206,N_29965,N_25491);
nor U33207 (N_33207,N_26135,N_27063);
or U33208 (N_33208,N_28778,N_29569);
nand U33209 (N_33209,N_27080,N_28907);
nand U33210 (N_33210,N_27944,N_29304);
nand U33211 (N_33211,N_26709,N_29966);
or U33212 (N_33212,N_26184,N_27360);
nor U33213 (N_33213,N_25927,N_28584);
nor U33214 (N_33214,N_29264,N_26613);
and U33215 (N_33215,N_28472,N_27381);
nand U33216 (N_33216,N_29581,N_29742);
nand U33217 (N_33217,N_26103,N_26755);
xnor U33218 (N_33218,N_29294,N_26139);
nor U33219 (N_33219,N_25829,N_26779);
nand U33220 (N_33220,N_28593,N_28621);
nand U33221 (N_33221,N_28120,N_25642);
or U33222 (N_33222,N_29007,N_27356);
nand U33223 (N_33223,N_29483,N_26775);
nor U33224 (N_33224,N_29841,N_29732);
and U33225 (N_33225,N_26923,N_27604);
and U33226 (N_33226,N_25042,N_27505);
and U33227 (N_33227,N_27230,N_26594);
nand U33228 (N_33228,N_27826,N_29343);
or U33229 (N_33229,N_26711,N_29501);
nor U33230 (N_33230,N_27037,N_25584);
nor U33231 (N_33231,N_26060,N_27583);
nand U33232 (N_33232,N_29376,N_25580);
and U33233 (N_33233,N_28638,N_25217);
and U33234 (N_33234,N_27024,N_25587);
xor U33235 (N_33235,N_27480,N_28836);
xnor U33236 (N_33236,N_26822,N_28185);
xnor U33237 (N_33237,N_29206,N_28434);
or U33238 (N_33238,N_25787,N_27120);
xnor U33239 (N_33239,N_25851,N_26028);
and U33240 (N_33240,N_28823,N_28300);
xor U33241 (N_33241,N_25895,N_29087);
or U33242 (N_33242,N_25602,N_27246);
nand U33243 (N_33243,N_25237,N_27923);
or U33244 (N_33244,N_26474,N_27272);
nand U33245 (N_33245,N_28481,N_29360);
and U33246 (N_33246,N_29065,N_26679);
nand U33247 (N_33247,N_29891,N_28449);
or U33248 (N_33248,N_27073,N_27928);
or U33249 (N_33249,N_26878,N_26480);
xnor U33250 (N_33250,N_29843,N_29088);
xnor U33251 (N_33251,N_26273,N_27436);
xor U33252 (N_33252,N_27075,N_25612);
or U33253 (N_33253,N_28608,N_29335);
nor U33254 (N_33254,N_28639,N_25206);
or U33255 (N_33255,N_27105,N_25200);
nand U33256 (N_33256,N_29670,N_27802);
nand U33257 (N_33257,N_25682,N_26985);
and U33258 (N_33258,N_28650,N_27865);
nor U33259 (N_33259,N_25275,N_25951);
and U33260 (N_33260,N_29572,N_25247);
or U33261 (N_33261,N_25430,N_25646);
and U33262 (N_33262,N_27346,N_27390);
or U33263 (N_33263,N_26338,N_28618);
or U33264 (N_33264,N_26434,N_28691);
nor U33265 (N_33265,N_29655,N_29742);
xnor U33266 (N_33266,N_25210,N_29959);
xnor U33267 (N_33267,N_26532,N_29215);
nand U33268 (N_33268,N_29193,N_25814);
and U33269 (N_33269,N_25834,N_29684);
nand U33270 (N_33270,N_27618,N_28790);
nand U33271 (N_33271,N_27169,N_25109);
xor U33272 (N_33272,N_27632,N_29588);
nand U33273 (N_33273,N_27189,N_29757);
nand U33274 (N_33274,N_29645,N_28160);
xor U33275 (N_33275,N_26310,N_28368);
or U33276 (N_33276,N_28774,N_26176);
nand U33277 (N_33277,N_25150,N_28379);
or U33278 (N_33278,N_28634,N_28222);
and U33279 (N_33279,N_25384,N_26913);
nor U33280 (N_33280,N_25932,N_29145);
nand U33281 (N_33281,N_26200,N_29128);
nand U33282 (N_33282,N_29735,N_26885);
nor U33283 (N_33283,N_28391,N_25307);
xnor U33284 (N_33284,N_27784,N_29345);
or U33285 (N_33285,N_29158,N_27679);
or U33286 (N_33286,N_29344,N_26841);
nor U33287 (N_33287,N_29304,N_29174);
nand U33288 (N_33288,N_27367,N_29391);
xnor U33289 (N_33289,N_26427,N_28777);
nor U33290 (N_33290,N_26056,N_26730);
nor U33291 (N_33291,N_29039,N_27996);
or U33292 (N_33292,N_29778,N_27059);
nand U33293 (N_33293,N_26857,N_26718);
and U33294 (N_33294,N_29729,N_26271);
or U33295 (N_33295,N_25710,N_29949);
nor U33296 (N_33296,N_25808,N_26184);
xor U33297 (N_33297,N_28202,N_26755);
nor U33298 (N_33298,N_28658,N_25645);
xor U33299 (N_33299,N_26757,N_26427);
nand U33300 (N_33300,N_27182,N_26608);
and U33301 (N_33301,N_26171,N_25048);
or U33302 (N_33302,N_29833,N_28696);
nor U33303 (N_33303,N_28817,N_25007);
nand U33304 (N_33304,N_26863,N_29235);
nor U33305 (N_33305,N_25382,N_27635);
nand U33306 (N_33306,N_26806,N_26539);
and U33307 (N_33307,N_26175,N_29189);
xor U33308 (N_33308,N_25621,N_29013);
nor U33309 (N_33309,N_29765,N_26211);
and U33310 (N_33310,N_26210,N_26831);
and U33311 (N_33311,N_25291,N_26077);
xor U33312 (N_33312,N_25997,N_25689);
nor U33313 (N_33313,N_25961,N_27127);
nand U33314 (N_33314,N_28761,N_26823);
or U33315 (N_33315,N_29280,N_25677);
xnor U33316 (N_33316,N_28633,N_28372);
nor U33317 (N_33317,N_27396,N_25601);
or U33318 (N_33318,N_26812,N_26843);
nand U33319 (N_33319,N_26963,N_26553);
xor U33320 (N_33320,N_27801,N_25703);
nand U33321 (N_33321,N_28693,N_28019);
or U33322 (N_33322,N_29226,N_26776);
nand U33323 (N_33323,N_28987,N_29860);
nand U33324 (N_33324,N_25769,N_28327);
nor U33325 (N_33325,N_29930,N_27455);
or U33326 (N_33326,N_28847,N_29336);
nor U33327 (N_33327,N_27687,N_29633);
nand U33328 (N_33328,N_26681,N_26695);
nand U33329 (N_33329,N_29414,N_26440);
xnor U33330 (N_33330,N_29804,N_26326);
or U33331 (N_33331,N_28949,N_25850);
nor U33332 (N_33332,N_27785,N_25517);
and U33333 (N_33333,N_29707,N_27184);
xor U33334 (N_33334,N_28872,N_27638);
xor U33335 (N_33335,N_29435,N_29944);
nor U33336 (N_33336,N_25365,N_25994);
xor U33337 (N_33337,N_29246,N_29972);
nand U33338 (N_33338,N_29762,N_25515);
or U33339 (N_33339,N_26992,N_26759);
and U33340 (N_33340,N_26266,N_26287);
and U33341 (N_33341,N_29890,N_27159);
nor U33342 (N_33342,N_25042,N_26383);
nand U33343 (N_33343,N_25442,N_25366);
xnor U33344 (N_33344,N_29880,N_27063);
xnor U33345 (N_33345,N_26564,N_28690);
nand U33346 (N_33346,N_27390,N_26636);
and U33347 (N_33347,N_29695,N_25869);
nor U33348 (N_33348,N_27182,N_29762);
nand U33349 (N_33349,N_26417,N_25788);
nand U33350 (N_33350,N_26475,N_25002);
and U33351 (N_33351,N_29538,N_28955);
or U33352 (N_33352,N_27608,N_27078);
or U33353 (N_33353,N_26557,N_29021);
or U33354 (N_33354,N_27294,N_29709);
or U33355 (N_33355,N_28545,N_28539);
and U33356 (N_33356,N_26939,N_25961);
xor U33357 (N_33357,N_28190,N_26184);
nand U33358 (N_33358,N_27555,N_29314);
nor U33359 (N_33359,N_26772,N_29486);
nand U33360 (N_33360,N_28367,N_25780);
or U33361 (N_33361,N_29763,N_25738);
nor U33362 (N_33362,N_29468,N_29876);
xnor U33363 (N_33363,N_25123,N_26082);
and U33364 (N_33364,N_27012,N_25142);
nand U33365 (N_33365,N_27160,N_28766);
xnor U33366 (N_33366,N_25186,N_29917);
nand U33367 (N_33367,N_25993,N_26626);
or U33368 (N_33368,N_29124,N_25588);
nor U33369 (N_33369,N_29351,N_28529);
and U33370 (N_33370,N_27241,N_29819);
nor U33371 (N_33371,N_27009,N_28635);
and U33372 (N_33372,N_26275,N_25823);
nor U33373 (N_33373,N_28029,N_29081);
nand U33374 (N_33374,N_29335,N_28133);
nand U33375 (N_33375,N_27648,N_26663);
nor U33376 (N_33376,N_28123,N_25605);
nand U33377 (N_33377,N_27822,N_28207);
and U33378 (N_33378,N_29618,N_27862);
xnor U33379 (N_33379,N_28896,N_26001);
nor U33380 (N_33380,N_25155,N_25929);
nor U33381 (N_33381,N_27063,N_28982);
nand U33382 (N_33382,N_25605,N_27101);
and U33383 (N_33383,N_29485,N_25325);
nand U33384 (N_33384,N_28679,N_25658);
or U33385 (N_33385,N_27672,N_27920);
or U33386 (N_33386,N_27017,N_26840);
xor U33387 (N_33387,N_28312,N_27134);
or U33388 (N_33388,N_29011,N_28846);
or U33389 (N_33389,N_27628,N_26905);
nand U33390 (N_33390,N_25650,N_28988);
nand U33391 (N_33391,N_26028,N_25610);
nor U33392 (N_33392,N_25283,N_27639);
xor U33393 (N_33393,N_26700,N_29245);
nor U33394 (N_33394,N_29343,N_26067);
nand U33395 (N_33395,N_25358,N_27738);
nor U33396 (N_33396,N_25677,N_28534);
nand U33397 (N_33397,N_25286,N_29146);
nand U33398 (N_33398,N_25203,N_29087);
nand U33399 (N_33399,N_27080,N_29111);
nand U33400 (N_33400,N_25157,N_28282);
xor U33401 (N_33401,N_26412,N_25597);
or U33402 (N_33402,N_28473,N_27213);
nor U33403 (N_33403,N_26627,N_29623);
nand U33404 (N_33404,N_25793,N_27816);
nor U33405 (N_33405,N_26862,N_27201);
or U33406 (N_33406,N_28801,N_27285);
nand U33407 (N_33407,N_25583,N_27661);
nor U33408 (N_33408,N_28678,N_28204);
nor U33409 (N_33409,N_27563,N_29527);
xor U33410 (N_33410,N_28842,N_28925);
and U33411 (N_33411,N_28224,N_27767);
nand U33412 (N_33412,N_25339,N_29079);
xnor U33413 (N_33413,N_29195,N_29805);
and U33414 (N_33414,N_29916,N_28443);
or U33415 (N_33415,N_28539,N_28770);
nor U33416 (N_33416,N_27853,N_25708);
nor U33417 (N_33417,N_28646,N_29926);
nor U33418 (N_33418,N_27528,N_29237);
nand U33419 (N_33419,N_29400,N_28698);
nand U33420 (N_33420,N_28772,N_25871);
nor U33421 (N_33421,N_27888,N_25672);
nand U33422 (N_33422,N_27447,N_25415);
nor U33423 (N_33423,N_27007,N_29985);
xnor U33424 (N_33424,N_26141,N_26627);
nor U33425 (N_33425,N_26671,N_25186);
xnor U33426 (N_33426,N_27168,N_26169);
xnor U33427 (N_33427,N_25700,N_26592);
nor U33428 (N_33428,N_28951,N_28580);
and U33429 (N_33429,N_27723,N_28638);
and U33430 (N_33430,N_29975,N_26966);
nand U33431 (N_33431,N_29472,N_29527);
nand U33432 (N_33432,N_25476,N_26285);
nand U33433 (N_33433,N_25681,N_27376);
and U33434 (N_33434,N_26158,N_27948);
nor U33435 (N_33435,N_26179,N_27169);
nor U33436 (N_33436,N_27518,N_28503);
xor U33437 (N_33437,N_26642,N_27728);
nand U33438 (N_33438,N_29417,N_29915);
nor U33439 (N_33439,N_26726,N_27751);
nand U33440 (N_33440,N_25088,N_25075);
nand U33441 (N_33441,N_25479,N_26188);
and U33442 (N_33442,N_26653,N_26796);
or U33443 (N_33443,N_25792,N_25703);
or U33444 (N_33444,N_26937,N_28472);
or U33445 (N_33445,N_27838,N_25629);
xor U33446 (N_33446,N_25786,N_27003);
nand U33447 (N_33447,N_27203,N_29917);
nor U33448 (N_33448,N_29712,N_27308);
nand U33449 (N_33449,N_28425,N_26468);
xnor U33450 (N_33450,N_29047,N_25636);
and U33451 (N_33451,N_28914,N_26127);
or U33452 (N_33452,N_26186,N_26796);
and U33453 (N_33453,N_28105,N_29029);
nand U33454 (N_33454,N_27252,N_29056);
and U33455 (N_33455,N_26807,N_25791);
nor U33456 (N_33456,N_29746,N_26891);
nand U33457 (N_33457,N_29601,N_25876);
and U33458 (N_33458,N_29123,N_26774);
and U33459 (N_33459,N_29256,N_26246);
nand U33460 (N_33460,N_28640,N_26251);
nor U33461 (N_33461,N_25333,N_26601);
or U33462 (N_33462,N_29341,N_29862);
xor U33463 (N_33463,N_29242,N_28411);
nand U33464 (N_33464,N_27798,N_29473);
nor U33465 (N_33465,N_27578,N_27390);
nor U33466 (N_33466,N_25049,N_25042);
nand U33467 (N_33467,N_26044,N_25943);
or U33468 (N_33468,N_26567,N_29956);
nand U33469 (N_33469,N_28530,N_27422);
and U33470 (N_33470,N_26858,N_26892);
or U33471 (N_33471,N_29374,N_27392);
xnor U33472 (N_33472,N_29729,N_26379);
nor U33473 (N_33473,N_25683,N_29185);
or U33474 (N_33474,N_26440,N_26267);
or U33475 (N_33475,N_29658,N_26597);
nor U33476 (N_33476,N_26702,N_27969);
or U33477 (N_33477,N_26293,N_26899);
and U33478 (N_33478,N_28370,N_29007);
nand U33479 (N_33479,N_26856,N_27932);
nand U33480 (N_33480,N_26488,N_27358);
and U33481 (N_33481,N_29228,N_27866);
or U33482 (N_33482,N_28747,N_29341);
or U33483 (N_33483,N_29118,N_25283);
and U33484 (N_33484,N_27738,N_28817);
nor U33485 (N_33485,N_28939,N_28172);
xor U33486 (N_33486,N_29808,N_29455);
nor U33487 (N_33487,N_25104,N_26557);
nand U33488 (N_33488,N_27773,N_28365);
and U33489 (N_33489,N_28918,N_27806);
xnor U33490 (N_33490,N_25832,N_26088);
nand U33491 (N_33491,N_26297,N_27400);
xnor U33492 (N_33492,N_27548,N_26822);
nand U33493 (N_33493,N_26318,N_25090);
nor U33494 (N_33494,N_28422,N_26813);
and U33495 (N_33495,N_27293,N_26259);
nand U33496 (N_33496,N_27035,N_25160);
nor U33497 (N_33497,N_28886,N_29283);
nand U33498 (N_33498,N_26448,N_29661);
nor U33499 (N_33499,N_25173,N_26391);
nor U33500 (N_33500,N_29730,N_26421);
and U33501 (N_33501,N_29114,N_29421);
xor U33502 (N_33502,N_25338,N_28308);
nand U33503 (N_33503,N_27300,N_26793);
or U33504 (N_33504,N_26597,N_28945);
xnor U33505 (N_33505,N_29330,N_25212);
or U33506 (N_33506,N_25698,N_27681);
and U33507 (N_33507,N_28740,N_25995);
xor U33508 (N_33508,N_28392,N_28659);
and U33509 (N_33509,N_28190,N_25306);
nand U33510 (N_33510,N_25914,N_26352);
or U33511 (N_33511,N_28585,N_26830);
nand U33512 (N_33512,N_27740,N_27419);
nand U33513 (N_33513,N_25611,N_26478);
and U33514 (N_33514,N_29045,N_28190);
nor U33515 (N_33515,N_27580,N_26076);
or U33516 (N_33516,N_29042,N_26628);
nand U33517 (N_33517,N_27679,N_26728);
and U33518 (N_33518,N_27228,N_29226);
or U33519 (N_33519,N_29822,N_29791);
xor U33520 (N_33520,N_29990,N_28482);
nor U33521 (N_33521,N_26426,N_27675);
nand U33522 (N_33522,N_29198,N_26563);
nand U33523 (N_33523,N_29438,N_28066);
or U33524 (N_33524,N_27936,N_25565);
or U33525 (N_33525,N_25834,N_25739);
and U33526 (N_33526,N_29295,N_29261);
or U33527 (N_33527,N_29818,N_27003);
nor U33528 (N_33528,N_28272,N_26778);
xor U33529 (N_33529,N_28600,N_27228);
nand U33530 (N_33530,N_26426,N_29006);
nand U33531 (N_33531,N_29657,N_28043);
xnor U33532 (N_33532,N_29373,N_25812);
xnor U33533 (N_33533,N_26691,N_25184);
nand U33534 (N_33534,N_29968,N_28575);
and U33535 (N_33535,N_28320,N_27044);
and U33536 (N_33536,N_26403,N_27972);
xor U33537 (N_33537,N_25523,N_27571);
nor U33538 (N_33538,N_29411,N_28166);
xor U33539 (N_33539,N_28628,N_29118);
or U33540 (N_33540,N_29045,N_25462);
and U33541 (N_33541,N_26424,N_26420);
nand U33542 (N_33542,N_26949,N_25126);
or U33543 (N_33543,N_28435,N_26034);
and U33544 (N_33544,N_26815,N_27187);
or U33545 (N_33545,N_26817,N_25495);
nor U33546 (N_33546,N_28385,N_27145);
xor U33547 (N_33547,N_27609,N_29793);
xor U33548 (N_33548,N_29057,N_27936);
nor U33549 (N_33549,N_25190,N_26391);
nor U33550 (N_33550,N_28370,N_27849);
or U33551 (N_33551,N_26669,N_25643);
or U33552 (N_33552,N_28922,N_29015);
and U33553 (N_33553,N_28755,N_26303);
and U33554 (N_33554,N_27502,N_29370);
xor U33555 (N_33555,N_26018,N_28954);
or U33556 (N_33556,N_29163,N_27365);
nor U33557 (N_33557,N_27169,N_26441);
nor U33558 (N_33558,N_29061,N_27302);
nand U33559 (N_33559,N_28400,N_27544);
or U33560 (N_33560,N_26996,N_29434);
or U33561 (N_33561,N_26945,N_25288);
and U33562 (N_33562,N_27059,N_25328);
nand U33563 (N_33563,N_29859,N_27853);
and U33564 (N_33564,N_27858,N_25593);
xor U33565 (N_33565,N_27901,N_25003);
or U33566 (N_33566,N_26882,N_29566);
xnor U33567 (N_33567,N_26219,N_26839);
and U33568 (N_33568,N_28012,N_26255);
xnor U33569 (N_33569,N_29511,N_28987);
nor U33570 (N_33570,N_29262,N_29320);
or U33571 (N_33571,N_29363,N_25837);
or U33572 (N_33572,N_28644,N_29221);
or U33573 (N_33573,N_27976,N_28315);
and U33574 (N_33574,N_29803,N_27094);
xnor U33575 (N_33575,N_26386,N_26092);
nor U33576 (N_33576,N_25129,N_28451);
and U33577 (N_33577,N_28819,N_28905);
or U33578 (N_33578,N_25118,N_28445);
nand U33579 (N_33579,N_29868,N_27088);
and U33580 (N_33580,N_25240,N_25218);
nand U33581 (N_33581,N_29863,N_25957);
nor U33582 (N_33582,N_26014,N_28202);
or U33583 (N_33583,N_26123,N_26347);
nand U33584 (N_33584,N_29840,N_29101);
nor U33585 (N_33585,N_26330,N_29099);
nand U33586 (N_33586,N_26074,N_25183);
nand U33587 (N_33587,N_26758,N_29202);
xnor U33588 (N_33588,N_26426,N_25677);
or U33589 (N_33589,N_29705,N_25396);
or U33590 (N_33590,N_27433,N_25755);
nand U33591 (N_33591,N_26150,N_27260);
nand U33592 (N_33592,N_29074,N_28287);
and U33593 (N_33593,N_28960,N_25739);
or U33594 (N_33594,N_25522,N_27892);
or U33595 (N_33595,N_28245,N_25542);
and U33596 (N_33596,N_26721,N_27542);
and U33597 (N_33597,N_27572,N_28090);
and U33598 (N_33598,N_28504,N_28598);
or U33599 (N_33599,N_27394,N_27950);
or U33600 (N_33600,N_27442,N_25804);
nor U33601 (N_33601,N_26690,N_26774);
and U33602 (N_33602,N_25768,N_25053);
or U33603 (N_33603,N_26428,N_25311);
xnor U33604 (N_33604,N_25882,N_27967);
nor U33605 (N_33605,N_27015,N_27113);
nor U33606 (N_33606,N_29442,N_25355);
nor U33607 (N_33607,N_27782,N_26991);
and U33608 (N_33608,N_29975,N_25709);
nor U33609 (N_33609,N_28756,N_25695);
nand U33610 (N_33610,N_28120,N_25566);
xor U33611 (N_33611,N_25842,N_26097);
and U33612 (N_33612,N_26053,N_25645);
or U33613 (N_33613,N_26925,N_25954);
nor U33614 (N_33614,N_26375,N_25473);
nand U33615 (N_33615,N_27836,N_28778);
xnor U33616 (N_33616,N_28664,N_27362);
nor U33617 (N_33617,N_28693,N_26500);
nor U33618 (N_33618,N_29106,N_29292);
nor U33619 (N_33619,N_29845,N_25248);
or U33620 (N_33620,N_25358,N_28409);
nor U33621 (N_33621,N_27043,N_27831);
and U33622 (N_33622,N_25693,N_28126);
or U33623 (N_33623,N_25223,N_26404);
nand U33624 (N_33624,N_29933,N_29050);
or U33625 (N_33625,N_26741,N_28921);
and U33626 (N_33626,N_29845,N_29370);
xnor U33627 (N_33627,N_29836,N_27557);
and U33628 (N_33628,N_27170,N_25282);
and U33629 (N_33629,N_27682,N_26734);
and U33630 (N_33630,N_28046,N_27710);
xnor U33631 (N_33631,N_27205,N_27153);
and U33632 (N_33632,N_27084,N_27968);
and U33633 (N_33633,N_29047,N_29459);
xnor U33634 (N_33634,N_25609,N_25990);
or U33635 (N_33635,N_25904,N_27597);
nor U33636 (N_33636,N_27113,N_27937);
nand U33637 (N_33637,N_29892,N_27717);
or U33638 (N_33638,N_26700,N_25388);
xnor U33639 (N_33639,N_27123,N_26954);
or U33640 (N_33640,N_28628,N_28398);
xor U33641 (N_33641,N_26291,N_25717);
nor U33642 (N_33642,N_25071,N_26810);
and U33643 (N_33643,N_27048,N_25324);
xnor U33644 (N_33644,N_26113,N_25932);
xor U33645 (N_33645,N_28224,N_29401);
and U33646 (N_33646,N_25013,N_27970);
and U33647 (N_33647,N_27509,N_27475);
nand U33648 (N_33648,N_27157,N_27373);
nor U33649 (N_33649,N_28896,N_25848);
and U33650 (N_33650,N_28345,N_25534);
and U33651 (N_33651,N_27667,N_28034);
and U33652 (N_33652,N_26187,N_25268);
nand U33653 (N_33653,N_25654,N_27757);
xor U33654 (N_33654,N_28034,N_29870);
xnor U33655 (N_33655,N_28395,N_28962);
nand U33656 (N_33656,N_26232,N_27476);
or U33657 (N_33657,N_29669,N_25287);
xnor U33658 (N_33658,N_29102,N_28721);
and U33659 (N_33659,N_26878,N_27161);
nor U33660 (N_33660,N_26381,N_28379);
nand U33661 (N_33661,N_29766,N_29538);
or U33662 (N_33662,N_27203,N_25642);
or U33663 (N_33663,N_27444,N_26303);
xor U33664 (N_33664,N_26453,N_26136);
nor U33665 (N_33665,N_27382,N_25717);
xnor U33666 (N_33666,N_29469,N_28940);
and U33667 (N_33667,N_27951,N_28527);
xnor U33668 (N_33668,N_25625,N_25075);
xor U33669 (N_33669,N_29021,N_28659);
and U33670 (N_33670,N_25433,N_26541);
nand U33671 (N_33671,N_28012,N_25279);
xor U33672 (N_33672,N_28379,N_28204);
or U33673 (N_33673,N_28791,N_25987);
or U33674 (N_33674,N_27237,N_26124);
nand U33675 (N_33675,N_26158,N_25048);
and U33676 (N_33676,N_26111,N_29081);
xor U33677 (N_33677,N_28844,N_25326);
nand U33678 (N_33678,N_29594,N_28350);
xor U33679 (N_33679,N_26481,N_29202);
and U33680 (N_33680,N_25269,N_29997);
and U33681 (N_33681,N_26235,N_27652);
nand U33682 (N_33682,N_27265,N_25797);
nand U33683 (N_33683,N_25194,N_27567);
nor U33684 (N_33684,N_26073,N_29646);
xnor U33685 (N_33685,N_27702,N_25443);
xor U33686 (N_33686,N_28426,N_27376);
and U33687 (N_33687,N_29372,N_26150);
and U33688 (N_33688,N_27790,N_26131);
or U33689 (N_33689,N_27745,N_26823);
and U33690 (N_33690,N_25126,N_28622);
xor U33691 (N_33691,N_28896,N_28631);
xnor U33692 (N_33692,N_25148,N_29492);
nor U33693 (N_33693,N_28648,N_26752);
and U33694 (N_33694,N_29740,N_27536);
nor U33695 (N_33695,N_26481,N_26418);
xnor U33696 (N_33696,N_26427,N_28827);
and U33697 (N_33697,N_27740,N_28600);
xnor U33698 (N_33698,N_29803,N_26893);
and U33699 (N_33699,N_27861,N_28126);
xnor U33700 (N_33700,N_26054,N_26981);
or U33701 (N_33701,N_27483,N_26338);
or U33702 (N_33702,N_29825,N_25401);
nor U33703 (N_33703,N_25637,N_25717);
and U33704 (N_33704,N_25241,N_29019);
or U33705 (N_33705,N_28339,N_25534);
nor U33706 (N_33706,N_29561,N_26775);
nor U33707 (N_33707,N_29843,N_29273);
nor U33708 (N_33708,N_28673,N_26270);
and U33709 (N_33709,N_27130,N_25651);
xor U33710 (N_33710,N_26891,N_25755);
or U33711 (N_33711,N_27491,N_29489);
nand U33712 (N_33712,N_27213,N_26682);
and U33713 (N_33713,N_27506,N_25021);
xnor U33714 (N_33714,N_26928,N_26429);
or U33715 (N_33715,N_28227,N_27554);
and U33716 (N_33716,N_29706,N_28806);
xnor U33717 (N_33717,N_27280,N_26255);
or U33718 (N_33718,N_29187,N_29366);
xnor U33719 (N_33719,N_27675,N_26978);
nor U33720 (N_33720,N_25880,N_29630);
nand U33721 (N_33721,N_26275,N_28298);
nand U33722 (N_33722,N_27170,N_26527);
or U33723 (N_33723,N_29580,N_26411);
or U33724 (N_33724,N_27163,N_25794);
xnor U33725 (N_33725,N_26751,N_29515);
nand U33726 (N_33726,N_26559,N_28560);
or U33727 (N_33727,N_26024,N_27564);
and U33728 (N_33728,N_29560,N_25575);
xor U33729 (N_33729,N_25169,N_25679);
nor U33730 (N_33730,N_26713,N_29440);
nor U33731 (N_33731,N_28837,N_26656);
nor U33732 (N_33732,N_28346,N_26070);
nor U33733 (N_33733,N_25473,N_26374);
nand U33734 (N_33734,N_28420,N_28815);
nor U33735 (N_33735,N_26035,N_29747);
and U33736 (N_33736,N_29132,N_29211);
and U33737 (N_33737,N_26912,N_29964);
or U33738 (N_33738,N_25440,N_27455);
nand U33739 (N_33739,N_28251,N_27352);
or U33740 (N_33740,N_25306,N_27346);
and U33741 (N_33741,N_28325,N_27533);
xnor U33742 (N_33742,N_25801,N_29801);
and U33743 (N_33743,N_26731,N_26517);
and U33744 (N_33744,N_25491,N_29685);
nor U33745 (N_33745,N_26166,N_26848);
nor U33746 (N_33746,N_27361,N_25072);
or U33747 (N_33747,N_29448,N_29877);
nor U33748 (N_33748,N_28373,N_26681);
or U33749 (N_33749,N_26223,N_28756);
or U33750 (N_33750,N_28604,N_27702);
nand U33751 (N_33751,N_26560,N_29918);
nand U33752 (N_33752,N_28482,N_25710);
or U33753 (N_33753,N_26770,N_25313);
nand U33754 (N_33754,N_25241,N_27186);
nand U33755 (N_33755,N_25435,N_29934);
or U33756 (N_33756,N_27813,N_25300);
xnor U33757 (N_33757,N_27586,N_29509);
or U33758 (N_33758,N_26442,N_27242);
nor U33759 (N_33759,N_27874,N_28456);
nor U33760 (N_33760,N_28893,N_28815);
nor U33761 (N_33761,N_27685,N_25299);
xor U33762 (N_33762,N_28206,N_25204);
nand U33763 (N_33763,N_29115,N_28292);
nand U33764 (N_33764,N_25676,N_25686);
and U33765 (N_33765,N_29968,N_28931);
xor U33766 (N_33766,N_29562,N_29041);
nand U33767 (N_33767,N_25601,N_29197);
xor U33768 (N_33768,N_26662,N_28571);
nand U33769 (N_33769,N_25066,N_25826);
and U33770 (N_33770,N_28081,N_28845);
nor U33771 (N_33771,N_25111,N_28338);
and U33772 (N_33772,N_28522,N_25758);
or U33773 (N_33773,N_29019,N_27422);
nand U33774 (N_33774,N_28181,N_28211);
and U33775 (N_33775,N_25368,N_26322);
and U33776 (N_33776,N_25193,N_26678);
xnor U33777 (N_33777,N_26833,N_28200);
nor U33778 (N_33778,N_25886,N_29904);
or U33779 (N_33779,N_28319,N_28042);
and U33780 (N_33780,N_28875,N_29332);
or U33781 (N_33781,N_26358,N_25701);
or U33782 (N_33782,N_27011,N_27370);
nor U33783 (N_33783,N_26694,N_29094);
and U33784 (N_33784,N_27258,N_29595);
nor U33785 (N_33785,N_29208,N_28820);
xor U33786 (N_33786,N_29472,N_26442);
or U33787 (N_33787,N_25299,N_28229);
xor U33788 (N_33788,N_26748,N_26828);
or U33789 (N_33789,N_28438,N_26239);
and U33790 (N_33790,N_26823,N_28948);
xnor U33791 (N_33791,N_28757,N_26516);
xor U33792 (N_33792,N_29387,N_29272);
nand U33793 (N_33793,N_27615,N_25895);
nand U33794 (N_33794,N_27223,N_28037);
and U33795 (N_33795,N_25198,N_26553);
nand U33796 (N_33796,N_29884,N_27367);
nand U33797 (N_33797,N_25914,N_26934);
nand U33798 (N_33798,N_27188,N_28343);
and U33799 (N_33799,N_26260,N_26833);
and U33800 (N_33800,N_27813,N_26135);
or U33801 (N_33801,N_29379,N_29823);
and U33802 (N_33802,N_28545,N_27500);
nor U33803 (N_33803,N_26152,N_27093);
or U33804 (N_33804,N_29202,N_26262);
nand U33805 (N_33805,N_26976,N_26506);
or U33806 (N_33806,N_26951,N_29561);
nand U33807 (N_33807,N_27543,N_29657);
and U33808 (N_33808,N_25347,N_27232);
xnor U33809 (N_33809,N_27261,N_27812);
nor U33810 (N_33810,N_27896,N_25658);
nor U33811 (N_33811,N_27852,N_29997);
nor U33812 (N_33812,N_26250,N_26075);
and U33813 (N_33813,N_28361,N_28581);
or U33814 (N_33814,N_28796,N_28334);
nand U33815 (N_33815,N_27507,N_26323);
nor U33816 (N_33816,N_26981,N_28402);
nand U33817 (N_33817,N_29451,N_28519);
xor U33818 (N_33818,N_28194,N_29285);
nor U33819 (N_33819,N_26728,N_27029);
nor U33820 (N_33820,N_27101,N_28732);
and U33821 (N_33821,N_25692,N_28229);
xor U33822 (N_33822,N_26608,N_25046);
and U33823 (N_33823,N_29728,N_26049);
xor U33824 (N_33824,N_28054,N_28609);
and U33825 (N_33825,N_25673,N_25692);
xnor U33826 (N_33826,N_26949,N_26315);
nor U33827 (N_33827,N_26118,N_27844);
nand U33828 (N_33828,N_25986,N_26797);
xor U33829 (N_33829,N_28135,N_26864);
and U33830 (N_33830,N_29252,N_25284);
or U33831 (N_33831,N_28138,N_29995);
and U33832 (N_33832,N_27487,N_27982);
nand U33833 (N_33833,N_27989,N_26968);
xor U33834 (N_33834,N_28870,N_28276);
or U33835 (N_33835,N_29190,N_27282);
and U33836 (N_33836,N_29404,N_26646);
nor U33837 (N_33837,N_27099,N_26400);
or U33838 (N_33838,N_29978,N_28966);
or U33839 (N_33839,N_29273,N_26618);
and U33840 (N_33840,N_28279,N_26353);
or U33841 (N_33841,N_27380,N_29663);
nand U33842 (N_33842,N_26125,N_25277);
xnor U33843 (N_33843,N_27045,N_27900);
and U33844 (N_33844,N_29419,N_28532);
xor U33845 (N_33845,N_25226,N_26434);
nand U33846 (N_33846,N_29748,N_29889);
nand U33847 (N_33847,N_27284,N_26677);
and U33848 (N_33848,N_25699,N_28223);
nand U33849 (N_33849,N_26957,N_29950);
nand U33850 (N_33850,N_26441,N_26623);
and U33851 (N_33851,N_27901,N_25345);
nand U33852 (N_33852,N_27213,N_27728);
xnor U33853 (N_33853,N_28705,N_28336);
or U33854 (N_33854,N_25116,N_29461);
and U33855 (N_33855,N_28477,N_26900);
xnor U33856 (N_33856,N_26515,N_28653);
xor U33857 (N_33857,N_25454,N_28179);
nor U33858 (N_33858,N_29712,N_26297);
nand U33859 (N_33859,N_28758,N_29903);
nor U33860 (N_33860,N_29870,N_29999);
nor U33861 (N_33861,N_28782,N_28404);
nand U33862 (N_33862,N_26022,N_27332);
nor U33863 (N_33863,N_26649,N_28507);
and U33864 (N_33864,N_28096,N_27125);
nand U33865 (N_33865,N_29672,N_27169);
or U33866 (N_33866,N_25536,N_26861);
nand U33867 (N_33867,N_29547,N_29222);
and U33868 (N_33868,N_27160,N_27824);
or U33869 (N_33869,N_29244,N_25067);
nand U33870 (N_33870,N_25847,N_25780);
or U33871 (N_33871,N_27082,N_26581);
or U33872 (N_33872,N_27153,N_29580);
nor U33873 (N_33873,N_28574,N_28746);
xor U33874 (N_33874,N_28581,N_25489);
and U33875 (N_33875,N_26551,N_29192);
nor U33876 (N_33876,N_27765,N_28752);
nand U33877 (N_33877,N_27939,N_28881);
nand U33878 (N_33878,N_28187,N_26568);
and U33879 (N_33879,N_29189,N_28007);
and U33880 (N_33880,N_26747,N_29762);
nor U33881 (N_33881,N_29999,N_29754);
nor U33882 (N_33882,N_26868,N_28947);
xnor U33883 (N_33883,N_27633,N_26171);
nor U33884 (N_33884,N_26461,N_29777);
nor U33885 (N_33885,N_28937,N_29626);
and U33886 (N_33886,N_29945,N_25617);
and U33887 (N_33887,N_27150,N_29519);
nor U33888 (N_33888,N_27283,N_27567);
nor U33889 (N_33889,N_25472,N_25695);
nand U33890 (N_33890,N_29972,N_28756);
or U33891 (N_33891,N_25000,N_27493);
and U33892 (N_33892,N_27230,N_28452);
or U33893 (N_33893,N_28068,N_28060);
nor U33894 (N_33894,N_26824,N_27400);
nor U33895 (N_33895,N_26255,N_26746);
xnor U33896 (N_33896,N_26152,N_29970);
xor U33897 (N_33897,N_29766,N_27032);
and U33898 (N_33898,N_25545,N_25336);
and U33899 (N_33899,N_27260,N_28864);
or U33900 (N_33900,N_25925,N_26972);
nor U33901 (N_33901,N_25476,N_28698);
or U33902 (N_33902,N_28921,N_25995);
or U33903 (N_33903,N_29019,N_27031);
nor U33904 (N_33904,N_28691,N_25572);
nand U33905 (N_33905,N_25936,N_29756);
and U33906 (N_33906,N_25416,N_27774);
nor U33907 (N_33907,N_26701,N_25545);
nor U33908 (N_33908,N_27185,N_29304);
xor U33909 (N_33909,N_28539,N_28050);
and U33910 (N_33910,N_25228,N_25525);
or U33911 (N_33911,N_26783,N_25424);
and U33912 (N_33912,N_29642,N_27586);
xnor U33913 (N_33913,N_25361,N_27481);
nand U33914 (N_33914,N_26347,N_29467);
or U33915 (N_33915,N_28597,N_29349);
nand U33916 (N_33916,N_26092,N_25817);
and U33917 (N_33917,N_28537,N_28493);
xor U33918 (N_33918,N_28239,N_27551);
xnor U33919 (N_33919,N_26966,N_28958);
xor U33920 (N_33920,N_26102,N_27493);
or U33921 (N_33921,N_25771,N_26830);
xor U33922 (N_33922,N_28966,N_25939);
nand U33923 (N_33923,N_26743,N_25564);
nand U33924 (N_33924,N_27878,N_26354);
nor U33925 (N_33925,N_28121,N_25127);
and U33926 (N_33926,N_27154,N_27773);
or U33927 (N_33927,N_25092,N_29979);
nand U33928 (N_33928,N_25468,N_28452);
and U33929 (N_33929,N_27220,N_25361);
xor U33930 (N_33930,N_27222,N_29828);
or U33931 (N_33931,N_28633,N_29226);
or U33932 (N_33932,N_28426,N_26382);
xnor U33933 (N_33933,N_28818,N_26784);
and U33934 (N_33934,N_28251,N_29846);
or U33935 (N_33935,N_29750,N_29246);
or U33936 (N_33936,N_27482,N_25138);
nor U33937 (N_33937,N_25651,N_26279);
nand U33938 (N_33938,N_27182,N_28954);
nand U33939 (N_33939,N_27664,N_25322);
xnor U33940 (N_33940,N_28767,N_27155);
nor U33941 (N_33941,N_25179,N_26539);
xor U33942 (N_33942,N_25586,N_28309);
nand U33943 (N_33943,N_28299,N_26128);
nor U33944 (N_33944,N_29284,N_27385);
and U33945 (N_33945,N_26273,N_27725);
nand U33946 (N_33946,N_28859,N_25537);
xnor U33947 (N_33947,N_27133,N_28374);
xor U33948 (N_33948,N_25788,N_28169);
and U33949 (N_33949,N_28945,N_26734);
xnor U33950 (N_33950,N_27654,N_28730);
and U33951 (N_33951,N_25125,N_25020);
nand U33952 (N_33952,N_26741,N_25058);
and U33953 (N_33953,N_29288,N_26243);
nand U33954 (N_33954,N_27882,N_29640);
or U33955 (N_33955,N_26163,N_28763);
nor U33956 (N_33956,N_25180,N_28561);
xor U33957 (N_33957,N_26070,N_25848);
xor U33958 (N_33958,N_27051,N_26399);
and U33959 (N_33959,N_29054,N_29867);
xnor U33960 (N_33960,N_28202,N_27142);
nand U33961 (N_33961,N_28408,N_27962);
nor U33962 (N_33962,N_29246,N_27089);
nor U33963 (N_33963,N_25450,N_27947);
nand U33964 (N_33964,N_25215,N_28199);
and U33965 (N_33965,N_26349,N_29117);
xnor U33966 (N_33966,N_27520,N_29634);
and U33967 (N_33967,N_28095,N_25890);
or U33968 (N_33968,N_26036,N_29694);
nor U33969 (N_33969,N_26935,N_25017);
nor U33970 (N_33970,N_29239,N_28973);
nand U33971 (N_33971,N_26049,N_27455);
xnor U33972 (N_33972,N_25803,N_28802);
xor U33973 (N_33973,N_26582,N_26808);
xor U33974 (N_33974,N_28546,N_29668);
xor U33975 (N_33975,N_25495,N_25767);
xnor U33976 (N_33976,N_26603,N_25598);
and U33977 (N_33977,N_27074,N_27453);
nor U33978 (N_33978,N_26179,N_25447);
nor U33979 (N_33979,N_25920,N_27633);
nand U33980 (N_33980,N_29094,N_26068);
or U33981 (N_33981,N_27466,N_28919);
or U33982 (N_33982,N_28136,N_25511);
nand U33983 (N_33983,N_28453,N_28724);
nor U33984 (N_33984,N_28109,N_27360);
or U33985 (N_33985,N_28254,N_27600);
nor U33986 (N_33986,N_29807,N_29611);
and U33987 (N_33987,N_25984,N_29564);
xnor U33988 (N_33988,N_25630,N_26343);
and U33989 (N_33989,N_29109,N_26691);
or U33990 (N_33990,N_25509,N_28996);
nand U33991 (N_33991,N_25488,N_25540);
nor U33992 (N_33992,N_28977,N_29858);
or U33993 (N_33993,N_25548,N_29111);
nand U33994 (N_33994,N_27719,N_29106);
or U33995 (N_33995,N_27541,N_25940);
or U33996 (N_33996,N_25092,N_28508);
or U33997 (N_33997,N_26259,N_29875);
nor U33998 (N_33998,N_29827,N_25972);
nand U33999 (N_33999,N_25673,N_28989);
and U34000 (N_34000,N_26392,N_27654);
or U34001 (N_34001,N_25681,N_25908);
nand U34002 (N_34002,N_26097,N_26361);
or U34003 (N_34003,N_26408,N_26612);
and U34004 (N_34004,N_25640,N_26643);
nor U34005 (N_34005,N_29293,N_29732);
and U34006 (N_34006,N_28183,N_27628);
or U34007 (N_34007,N_26894,N_27098);
or U34008 (N_34008,N_28590,N_27844);
or U34009 (N_34009,N_28256,N_25374);
or U34010 (N_34010,N_28992,N_29099);
xor U34011 (N_34011,N_29329,N_25359);
nor U34012 (N_34012,N_28124,N_25292);
and U34013 (N_34013,N_25959,N_27956);
or U34014 (N_34014,N_26024,N_25098);
and U34015 (N_34015,N_26008,N_27946);
or U34016 (N_34016,N_26550,N_27845);
nand U34017 (N_34017,N_28100,N_25616);
or U34018 (N_34018,N_27803,N_27216);
xnor U34019 (N_34019,N_28164,N_28945);
or U34020 (N_34020,N_28141,N_25770);
nand U34021 (N_34021,N_29615,N_26704);
xor U34022 (N_34022,N_26131,N_25742);
or U34023 (N_34023,N_28779,N_27242);
and U34024 (N_34024,N_26531,N_28390);
or U34025 (N_34025,N_26465,N_26546);
nor U34026 (N_34026,N_26260,N_28785);
xnor U34027 (N_34027,N_25314,N_27662);
nand U34028 (N_34028,N_28480,N_27918);
nor U34029 (N_34029,N_28372,N_29298);
or U34030 (N_34030,N_28090,N_26284);
nand U34031 (N_34031,N_26355,N_25599);
or U34032 (N_34032,N_26532,N_25879);
xnor U34033 (N_34033,N_28722,N_25970);
or U34034 (N_34034,N_26119,N_25888);
and U34035 (N_34035,N_26735,N_26524);
nand U34036 (N_34036,N_27549,N_25523);
nor U34037 (N_34037,N_26517,N_29273);
xor U34038 (N_34038,N_25935,N_27489);
or U34039 (N_34039,N_28604,N_27995);
nor U34040 (N_34040,N_25403,N_29590);
nor U34041 (N_34041,N_28937,N_27845);
or U34042 (N_34042,N_25859,N_27144);
nor U34043 (N_34043,N_28102,N_25087);
nor U34044 (N_34044,N_25420,N_25933);
nor U34045 (N_34045,N_28566,N_25195);
nor U34046 (N_34046,N_29864,N_28081);
and U34047 (N_34047,N_26539,N_25257);
and U34048 (N_34048,N_27175,N_25000);
or U34049 (N_34049,N_27832,N_29433);
or U34050 (N_34050,N_26108,N_26219);
nor U34051 (N_34051,N_26935,N_25825);
xnor U34052 (N_34052,N_26765,N_29817);
nor U34053 (N_34053,N_25228,N_27564);
and U34054 (N_34054,N_27530,N_25614);
nor U34055 (N_34055,N_25337,N_28314);
and U34056 (N_34056,N_28254,N_28252);
nor U34057 (N_34057,N_25618,N_29365);
and U34058 (N_34058,N_26581,N_28670);
and U34059 (N_34059,N_28997,N_27901);
xor U34060 (N_34060,N_26102,N_27756);
and U34061 (N_34061,N_26558,N_25258);
or U34062 (N_34062,N_26880,N_29878);
xnor U34063 (N_34063,N_29009,N_28652);
nand U34064 (N_34064,N_27581,N_29827);
and U34065 (N_34065,N_26926,N_29969);
xnor U34066 (N_34066,N_28065,N_26277);
nor U34067 (N_34067,N_27173,N_26753);
xnor U34068 (N_34068,N_25821,N_25627);
xnor U34069 (N_34069,N_26114,N_27771);
nor U34070 (N_34070,N_25681,N_26689);
xor U34071 (N_34071,N_27417,N_28628);
nor U34072 (N_34072,N_25386,N_28780);
and U34073 (N_34073,N_29035,N_26720);
and U34074 (N_34074,N_27493,N_27562);
xnor U34075 (N_34075,N_29086,N_28549);
nand U34076 (N_34076,N_28937,N_28405);
nor U34077 (N_34077,N_26712,N_25521);
nand U34078 (N_34078,N_27777,N_25717);
or U34079 (N_34079,N_25979,N_26660);
nand U34080 (N_34080,N_29727,N_27118);
xnor U34081 (N_34081,N_29433,N_29934);
nor U34082 (N_34082,N_25262,N_29208);
or U34083 (N_34083,N_25328,N_26918);
nor U34084 (N_34084,N_26149,N_25486);
nor U34085 (N_34085,N_29047,N_27722);
or U34086 (N_34086,N_25075,N_25602);
nor U34087 (N_34087,N_29657,N_29343);
or U34088 (N_34088,N_26760,N_26548);
and U34089 (N_34089,N_27297,N_27773);
or U34090 (N_34090,N_27091,N_26524);
nor U34091 (N_34091,N_27334,N_26790);
nor U34092 (N_34092,N_26245,N_28682);
or U34093 (N_34093,N_28947,N_29864);
nor U34094 (N_34094,N_26249,N_27267);
xor U34095 (N_34095,N_29314,N_27399);
or U34096 (N_34096,N_25270,N_26221);
nor U34097 (N_34097,N_28794,N_29532);
nand U34098 (N_34098,N_29478,N_28910);
nand U34099 (N_34099,N_25697,N_28816);
nor U34100 (N_34100,N_27561,N_29103);
or U34101 (N_34101,N_26943,N_29394);
and U34102 (N_34102,N_27660,N_25105);
and U34103 (N_34103,N_27976,N_25743);
nand U34104 (N_34104,N_26587,N_26584);
xor U34105 (N_34105,N_26956,N_26023);
xnor U34106 (N_34106,N_29202,N_27893);
nor U34107 (N_34107,N_27948,N_29673);
nand U34108 (N_34108,N_26034,N_29160);
nand U34109 (N_34109,N_25673,N_28371);
and U34110 (N_34110,N_29252,N_26700);
nor U34111 (N_34111,N_25278,N_29207);
and U34112 (N_34112,N_25019,N_26842);
nand U34113 (N_34113,N_27392,N_25310);
xor U34114 (N_34114,N_26757,N_26445);
nand U34115 (N_34115,N_27189,N_28001);
xor U34116 (N_34116,N_27242,N_28827);
nor U34117 (N_34117,N_28348,N_25075);
xor U34118 (N_34118,N_28867,N_29180);
nor U34119 (N_34119,N_26279,N_25501);
nand U34120 (N_34120,N_29140,N_27837);
nand U34121 (N_34121,N_29354,N_27989);
nor U34122 (N_34122,N_27269,N_28056);
nand U34123 (N_34123,N_27916,N_25190);
nor U34124 (N_34124,N_25188,N_28556);
nor U34125 (N_34125,N_29499,N_28695);
nand U34126 (N_34126,N_28679,N_28674);
xnor U34127 (N_34127,N_28216,N_25423);
nor U34128 (N_34128,N_28654,N_26151);
nand U34129 (N_34129,N_27101,N_25132);
nand U34130 (N_34130,N_27137,N_28628);
and U34131 (N_34131,N_26045,N_29409);
or U34132 (N_34132,N_26394,N_29861);
and U34133 (N_34133,N_28440,N_25648);
or U34134 (N_34134,N_28042,N_28585);
xor U34135 (N_34135,N_25136,N_28233);
xor U34136 (N_34136,N_28037,N_29605);
nor U34137 (N_34137,N_26717,N_28577);
or U34138 (N_34138,N_28259,N_29923);
nor U34139 (N_34139,N_28670,N_25879);
or U34140 (N_34140,N_25547,N_28794);
nor U34141 (N_34141,N_26131,N_27826);
nor U34142 (N_34142,N_28053,N_26677);
or U34143 (N_34143,N_29396,N_25920);
or U34144 (N_34144,N_26449,N_26060);
xnor U34145 (N_34145,N_25759,N_29980);
xor U34146 (N_34146,N_26895,N_28739);
or U34147 (N_34147,N_27845,N_28550);
or U34148 (N_34148,N_25485,N_27058);
nand U34149 (N_34149,N_25913,N_28083);
nand U34150 (N_34150,N_25484,N_26158);
or U34151 (N_34151,N_25031,N_27175);
and U34152 (N_34152,N_27704,N_28769);
nor U34153 (N_34153,N_28310,N_25700);
xnor U34154 (N_34154,N_29236,N_29115);
or U34155 (N_34155,N_28323,N_25588);
or U34156 (N_34156,N_27522,N_26784);
nor U34157 (N_34157,N_25547,N_26639);
xnor U34158 (N_34158,N_25593,N_27130);
nor U34159 (N_34159,N_29568,N_29583);
xnor U34160 (N_34160,N_25979,N_27793);
xor U34161 (N_34161,N_27564,N_28345);
nor U34162 (N_34162,N_27833,N_27801);
xor U34163 (N_34163,N_28477,N_27800);
or U34164 (N_34164,N_27199,N_26592);
or U34165 (N_34165,N_25835,N_28938);
or U34166 (N_34166,N_26736,N_27638);
nor U34167 (N_34167,N_28805,N_27100);
nor U34168 (N_34168,N_29683,N_27573);
and U34169 (N_34169,N_28732,N_26743);
and U34170 (N_34170,N_26171,N_25180);
xor U34171 (N_34171,N_26104,N_25400);
xor U34172 (N_34172,N_29623,N_25173);
nand U34173 (N_34173,N_27805,N_26692);
or U34174 (N_34174,N_26384,N_29210);
nand U34175 (N_34175,N_28110,N_27731);
xor U34176 (N_34176,N_29392,N_26231);
and U34177 (N_34177,N_25945,N_27290);
xnor U34178 (N_34178,N_25302,N_29646);
xnor U34179 (N_34179,N_27235,N_28934);
nand U34180 (N_34180,N_25553,N_28224);
nor U34181 (N_34181,N_27626,N_25202);
or U34182 (N_34182,N_28681,N_26777);
nor U34183 (N_34183,N_25706,N_27887);
or U34184 (N_34184,N_25720,N_28990);
nand U34185 (N_34185,N_28142,N_26371);
nand U34186 (N_34186,N_26562,N_28520);
xnor U34187 (N_34187,N_28252,N_27098);
nand U34188 (N_34188,N_26513,N_29381);
nor U34189 (N_34189,N_27508,N_29127);
and U34190 (N_34190,N_27223,N_28087);
nand U34191 (N_34191,N_26803,N_26360);
or U34192 (N_34192,N_27752,N_27453);
nor U34193 (N_34193,N_26806,N_29820);
nor U34194 (N_34194,N_25020,N_29130);
and U34195 (N_34195,N_26790,N_26288);
nand U34196 (N_34196,N_26464,N_25850);
nor U34197 (N_34197,N_29085,N_25439);
and U34198 (N_34198,N_25062,N_26829);
nor U34199 (N_34199,N_29508,N_27666);
nand U34200 (N_34200,N_27421,N_25103);
nand U34201 (N_34201,N_27348,N_27842);
or U34202 (N_34202,N_25273,N_27406);
xnor U34203 (N_34203,N_28564,N_25106);
nor U34204 (N_34204,N_27455,N_29992);
or U34205 (N_34205,N_27645,N_27849);
or U34206 (N_34206,N_26500,N_26773);
and U34207 (N_34207,N_29127,N_27159);
and U34208 (N_34208,N_25088,N_29886);
nand U34209 (N_34209,N_26155,N_28540);
nand U34210 (N_34210,N_27223,N_29696);
nor U34211 (N_34211,N_26763,N_27536);
xnor U34212 (N_34212,N_26406,N_25469);
and U34213 (N_34213,N_28064,N_29111);
xnor U34214 (N_34214,N_25967,N_26559);
or U34215 (N_34215,N_25758,N_25033);
nor U34216 (N_34216,N_27763,N_26040);
xor U34217 (N_34217,N_28494,N_28744);
nand U34218 (N_34218,N_29562,N_25025);
nor U34219 (N_34219,N_27812,N_27862);
xor U34220 (N_34220,N_29507,N_26247);
xnor U34221 (N_34221,N_26634,N_25458);
or U34222 (N_34222,N_27584,N_28246);
or U34223 (N_34223,N_25120,N_25301);
xnor U34224 (N_34224,N_29298,N_27257);
or U34225 (N_34225,N_29161,N_25818);
nor U34226 (N_34226,N_25173,N_29059);
or U34227 (N_34227,N_25235,N_27231);
and U34228 (N_34228,N_25893,N_28489);
or U34229 (N_34229,N_29438,N_29554);
and U34230 (N_34230,N_28519,N_26538);
and U34231 (N_34231,N_26450,N_28581);
or U34232 (N_34232,N_28935,N_25233);
and U34233 (N_34233,N_29558,N_28558);
xor U34234 (N_34234,N_29748,N_27112);
xnor U34235 (N_34235,N_27558,N_27814);
nor U34236 (N_34236,N_26815,N_27827);
nand U34237 (N_34237,N_27590,N_25642);
and U34238 (N_34238,N_27000,N_25682);
xnor U34239 (N_34239,N_27853,N_27803);
and U34240 (N_34240,N_29933,N_26719);
nor U34241 (N_34241,N_28139,N_28038);
nand U34242 (N_34242,N_29907,N_29823);
xor U34243 (N_34243,N_28552,N_25525);
nand U34244 (N_34244,N_28493,N_28765);
or U34245 (N_34245,N_28033,N_25307);
nor U34246 (N_34246,N_29278,N_29246);
or U34247 (N_34247,N_29836,N_29802);
nor U34248 (N_34248,N_25343,N_25624);
and U34249 (N_34249,N_26530,N_27716);
nor U34250 (N_34250,N_25581,N_26323);
or U34251 (N_34251,N_26761,N_26214);
xnor U34252 (N_34252,N_26120,N_27759);
or U34253 (N_34253,N_29140,N_27154);
or U34254 (N_34254,N_29942,N_27717);
or U34255 (N_34255,N_28690,N_28589);
or U34256 (N_34256,N_27155,N_28064);
xor U34257 (N_34257,N_28643,N_27470);
and U34258 (N_34258,N_27285,N_29236);
nand U34259 (N_34259,N_25426,N_25261);
nor U34260 (N_34260,N_25606,N_25229);
and U34261 (N_34261,N_26084,N_28922);
or U34262 (N_34262,N_28279,N_26248);
or U34263 (N_34263,N_27366,N_27097);
xnor U34264 (N_34264,N_29286,N_26752);
xnor U34265 (N_34265,N_28248,N_25352);
or U34266 (N_34266,N_26402,N_28343);
nor U34267 (N_34267,N_28131,N_26620);
nor U34268 (N_34268,N_26759,N_28983);
xor U34269 (N_34269,N_27905,N_29487);
nand U34270 (N_34270,N_27433,N_28718);
nand U34271 (N_34271,N_29216,N_28649);
xnor U34272 (N_34272,N_26346,N_25846);
xnor U34273 (N_34273,N_26099,N_27310);
nor U34274 (N_34274,N_28890,N_26808);
nand U34275 (N_34275,N_29361,N_27961);
nor U34276 (N_34276,N_25465,N_25737);
and U34277 (N_34277,N_29033,N_26759);
and U34278 (N_34278,N_28158,N_28304);
xor U34279 (N_34279,N_26166,N_26287);
and U34280 (N_34280,N_25711,N_29118);
xor U34281 (N_34281,N_28054,N_25963);
or U34282 (N_34282,N_26391,N_28784);
or U34283 (N_34283,N_26037,N_25097);
nand U34284 (N_34284,N_29137,N_29506);
nor U34285 (N_34285,N_29027,N_27434);
nor U34286 (N_34286,N_28279,N_25567);
xor U34287 (N_34287,N_25526,N_26830);
nand U34288 (N_34288,N_28064,N_28840);
nand U34289 (N_34289,N_28598,N_28148);
nor U34290 (N_34290,N_26415,N_26267);
or U34291 (N_34291,N_27017,N_28252);
nor U34292 (N_34292,N_28592,N_27741);
nor U34293 (N_34293,N_28127,N_28802);
or U34294 (N_34294,N_28306,N_29082);
or U34295 (N_34295,N_29734,N_26567);
or U34296 (N_34296,N_26220,N_29533);
and U34297 (N_34297,N_25208,N_28335);
and U34298 (N_34298,N_27306,N_29844);
nand U34299 (N_34299,N_26351,N_29460);
or U34300 (N_34300,N_28696,N_26156);
nor U34301 (N_34301,N_28909,N_27097);
or U34302 (N_34302,N_29371,N_26051);
or U34303 (N_34303,N_25234,N_26824);
and U34304 (N_34304,N_26602,N_29919);
or U34305 (N_34305,N_26367,N_29926);
nand U34306 (N_34306,N_26116,N_29646);
and U34307 (N_34307,N_25324,N_26391);
or U34308 (N_34308,N_25180,N_25223);
nor U34309 (N_34309,N_26461,N_29195);
nand U34310 (N_34310,N_29128,N_29186);
or U34311 (N_34311,N_26400,N_29077);
and U34312 (N_34312,N_28913,N_29559);
nand U34313 (N_34313,N_27569,N_27222);
and U34314 (N_34314,N_26591,N_26471);
nand U34315 (N_34315,N_29893,N_25057);
and U34316 (N_34316,N_28442,N_25778);
or U34317 (N_34317,N_28521,N_25155);
nor U34318 (N_34318,N_27416,N_29514);
xor U34319 (N_34319,N_29425,N_28100);
nor U34320 (N_34320,N_28492,N_27205);
or U34321 (N_34321,N_28088,N_25074);
xnor U34322 (N_34322,N_28234,N_26463);
nor U34323 (N_34323,N_29143,N_28512);
xnor U34324 (N_34324,N_27789,N_29303);
nor U34325 (N_34325,N_27858,N_29631);
and U34326 (N_34326,N_25011,N_25361);
and U34327 (N_34327,N_25787,N_25357);
xnor U34328 (N_34328,N_25318,N_28565);
nand U34329 (N_34329,N_26807,N_28285);
nand U34330 (N_34330,N_27414,N_25491);
and U34331 (N_34331,N_29517,N_25945);
nand U34332 (N_34332,N_29820,N_27722);
nor U34333 (N_34333,N_25104,N_25033);
xnor U34334 (N_34334,N_26850,N_28987);
or U34335 (N_34335,N_28764,N_28376);
nor U34336 (N_34336,N_29359,N_27157);
or U34337 (N_34337,N_27395,N_28322);
nor U34338 (N_34338,N_28647,N_25778);
xor U34339 (N_34339,N_25164,N_29564);
or U34340 (N_34340,N_28295,N_28036);
and U34341 (N_34341,N_29228,N_27109);
or U34342 (N_34342,N_26542,N_26635);
xnor U34343 (N_34343,N_29340,N_28610);
xnor U34344 (N_34344,N_29456,N_27379);
nand U34345 (N_34345,N_25192,N_26165);
nand U34346 (N_34346,N_28458,N_27486);
xnor U34347 (N_34347,N_29580,N_25203);
and U34348 (N_34348,N_25966,N_28851);
or U34349 (N_34349,N_25848,N_25062);
xor U34350 (N_34350,N_26740,N_28671);
and U34351 (N_34351,N_26835,N_28313);
and U34352 (N_34352,N_25732,N_27548);
or U34353 (N_34353,N_26901,N_26322);
and U34354 (N_34354,N_26752,N_29248);
and U34355 (N_34355,N_27682,N_28529);
nand U34356 (N_34356,N_26939,N_26913);
or U34357 (N_34357,N_28692,N_25440);
xor U34358 (N_34358,N_26580,N_26601);
xor U34359 (N_34359,N_25055,N_27653);
nand U34360 (N_34360,N_25331,N_27592);
or U34361 (N_34361,N_25731,N_29182);
nand U34362 (N_34362,N_25509,N_28846);
nand U34363 (N_34363,N_26184,N_28468);
nor U34364 (N_34364,N_29271,N_27512);
nand U34365 (N_34365,N_25064,N_25939);
and U34366 (N_34366,N_27008,N_25382);
xnor U34367 (N_34367,N_27310,N_26258);
nand U34368 (N_34368,N_25893,N_27358);
and U34369 (N_34369,N_26587,N_29363);
and U34370 (N_34370,N_28290,N_26261);
nand U34371 (N_34371,N_25083,N_26967);
nand U34372 (N_34372,N_27097,N_28027);
or U34373 (N_34373,N_27862,N_25137);
nand U34374 (N_34374,N_25159,N_26447);
and U34375 (N_34375,N_27965,N_27997);
and U34376 (N_34376,N_25415,N_29291);
xor U34377 (N_34377,N_29059,N_27790);
or U34378 (N_34378,N_25277,N_27817);
and U34379 (N_34379,N_25408,N_26608);
nor U34380 (N_34380,N_28737,N_29872);
nand U34381 (N_34381,N_28229,N_28635);
nand U34382 (N_34382,N_25405,N_26630);
nor U34383 (N_34383,N_27381,N_29975);
or U34384 (N_34384,N_27293,N_27007);
xor U34385 (N_34385,N_25520,N_29790);
or U34386 (N_34386,N_25371,N_27185);
nor U34387 (N_34387,N_28111,N_29475);
nand U34388 (N_34388,N_25799,N_26362);
and U34389 (N_34389,N_27007,N_29632);
nand U34390 (N_34390,N_27609,N_27907);
xor U34391 (N_34391,N_29114,N_28833);
nand U34392 (N_34392,N_25230,N_27481);
or U34393 (N_34393,N_28323,N_29509);
and U34394 (N_34394,N_25634,N_29144);
xor U34395 (N_34395,N_26255,N_27995);
xnor U34396 (N_34396,N_26899,N_26025);
or U34397 (N_34397,N_25963,N_28033);
nand U34398 (N_34398,N_25977,N_26657);
or U34399 (N_34399,N_26945,N_28227);
and U34400 (N_34400,N_25607,N_25296);
nor U34401 (N_34401,N_25430,N_29113);
nand U34402 (N_34402,N_27815,N_27844);
nand U34403 (N_34403,N_26698,N_25219);
or U34404 (N_34404,N_29357,N_27074);
nor U34405 (N_34405,N_29348,N_28527);
and U34406 (N_34406,N_25727,N_29256);
nor U34407 (N_34407,N_28154,N_26993);
or U34408 (N_34408,N_29530,N_26890);
xor U34409 (N_34409,N_28696,N_25331);
or U34410 (N_34410,N_25588,N_29195);
or U34411 (N_34411,N_26580,N_26300);
xnor U34412 (N_34412,N_26972,N_28960);
nor U34413 (N_34413,N_26865,N_26670);
nand U34414 (N_34414,N_26641,N_26886);
xnor U34415 (N_34415,N_26589,N_28507);
nand U34416 (N_34416,N_27107,N_26262);
and U34417 (N_34417,N_28090,N_26925);
nor U34418 (N_34418,N_26570,N_29771);
or U34419 (N_34419,N_29619,N_27347);
nand U34420 (N_34420,N_29934,N_27116);
nor U34421 (N_34421,N_28614,N_29497);
nor U34422 (N_34422,N_25167,N_28135);
and U34423 (N_34423,N_27016,N_26680);
nand U34424 (N_34424,N_25857,N_27748);
nor U34425 (N_34425,N_28786,N_26807);
nand U34426 (N_34426,N_29630,N_28108);
xnor U34427 (N_34427,N_28199,N_26993);
xnor U34428 (N_34428,N_25937,N_29610);
xor U34429 (N_34429,N_25081,N_27032);
xnor U34430 (N_34430,N_26063,N_29984);
nor U34431 (N_34431,N_25200,N_25844);
nand U34432 (N_34432,N_27205,N_28886);
nand U34433 (N_34433,N_25773,N_26782);
nand U34434 (N_34434,N_26735,N_27020);
nor U34435 (N_34435,N_25960,N_26532);
nand U34436 (N_34436,N_27844,N_26773);
xnor U34437 (N_34437,N_28218,N_29598);
nand U34438 (N_34438,N_29880,N_29239);
nand U34439 (N_34439,N_27382,N_26926);
xor U34440 (N_34440,N_26795,N_27488);
and U34441 (N_34441,N_26252,N_28236);
or U34442 (N_34442,N_25045,N_29659);
xnor U34443 (N_34443,N_28773,N_28022);
and U34444 (N_34444,N_25044,N_27931);
or U34445 (N_34445,N_25877,N_29919);
and U34446 (N_34446,N_29057,N_26811);
xor U34447 (N_34447,N_25117,N_27417);
nor U34448 (N_34448,N_26296,N_27602);
or U34449 (N_34449,N_27903,N_26881);
and U34450 (N_34450,N_29425,N_25089);
nand U34451 (N_34451,N_29580,N_28465);
nor U34452 (N_34452,N_25835,N_28117);
nor U34453 (N_34453,N_25630,N_27017);
or U34454 (N_34454,N_28287,N_27256);
nand U34455 (N_34455,N_27805,N_28976);
and U34456 (N_34456,N_29758,N_29770);
nand U34457 (N_34457,N_27847,N_25588);
or U34458 (N_34458,N_27041,N_25600);
or U34459 (N_34459,N_28026,N_29998);
or U34460 (N_34460,N_25942,N_27554);
xnor U34461 (N_34461,N_25702,N_29241);
xor U34462 (N_34462,N_25061,N_29218);
nor U34463 (N_34463,N_28654,N_26897);
or U34464 (N_34464,N_26162,N_28783);
xnor U34465 (N_34465,N_29378,N_29490);
xor U34466 (N_34466,N_25550,N_27879);
nand U34467 (N_34467,N_28886,N_28474);
and U34468 (N_34468,N_27743,N_28405);
nor U34469 (N_34469,N_28335,N_29099);
xor U34470 (N_34470,N_25718,N_27866);
and U34471 (N_34471,N_26359,N_28825);
nor U34472 (N_34472,N_29967,N_26666);
or U34473 (N_34473,N_26345,N_27730);
xnor U34474 (N_34474,N_28748,N_28988);
xnor U34475 (N_34475,N_25783,N_29642);
or U34476 (N_34476,N_26148,N_29392);
and U34477 (N_34477,N_25588,N_29291);
and U34478 (N_34478,N_28739,N_25292);
nand U34479 (N_34479,N_28303,N_26992);
nor U34480 (N_34480,N_29580,N_25702);
nand U34481 (N_34481,N_29427,N_27282);
xnor U34482 (N_34482,N_28843,N_29130);
xnor U34483 (N_34483,N_26516,N_26558);
or U34484 (N_34484,N_28876,N_25809);
and U34485 (N_34485,N_27652,N_26206);
nand U34486 (N_34486,N_27599,N_29713);
or U34487 (N_34487,N_25962,N_26684);
or U34488 (N_34488,N_27981,N_27809);
nor U34489 (N_34489,N_26775,N_28496);
xor U34490 (N_34490,N_25566,N_27742);
nand U34491 (N_34491,N_26907,N_27113);
nand U34492 (N_34492,N_27576,N_29267);
nand U34493 (N_34493,N_26937,N_26012);
nor U34494 (N_34494,N_29688,N_29610);
nand U34495 (N_34495,N_27587,N_27237);
nor U34496 (N_34496,N_28001,N_25850);
or U34497 (N_34497,N_29199,N_25770);
and U34498 (N_34498,N_29506,N_29492);
and U34499 (N_34499,N_27617,N_26336);
nand U34500 (N_34500,N_26735,N_29760);
or U34501 (N_34501,N_27539,N_26095);
nor U34502 (N_34502,N_28034,N_27566);
xor U34503 (N_34503,N_26688,N_27221);
or U34504 (N_34504,N_27038,N_29540);
nor U34505 (N_34505,N_26472,N_25494);
xnor U34506 (N_34506,N_28896,N_29885);
xnor U34507 (N_34507,N_27066,N_27454);
nand U34508 (N_34508,N_27315,N_28285);
and U34509 (N_34509,N_26081,N_25550);
xnor U34510 (N_34510,N_28968,N_26767);
or U34511 (N_34511,N_28884,N_28251);
and U34512 (N_34512,N_26760,N_26623);
nor U34513 (N_34513,N_26767,N_26036);
or U34514 (N_34514,N_26426,N_29614);
nand U34515 (N_34515,N_27935,N_25653);
and U34516 (N_34516,N_27134,N_25131);
nand U34517 (N_34517,N_27333,N_26454);
xor U34518 (N_34518,N_25657,N_29653);
xor U34519 (N_34519,N_25570,N_28773);
and U34520 (N_34520,N_27637,N_26128);
and U34521 (N_34521,N_25703,N_27520);
nand U34522 (N_34522,N_29404,N_27631);
and U34523 (N_34523,N_28786,N_26289);
nand U34524 (N_34524,N_27871,N_26630);
and U34525 (N_34525,N_25033,N_27785);
xor U34526 (N_34526,N_29693,N_26772);
or U34527 (N_34527,N_29300,N_25144);
nor U34528 (N_34528,N_25570,N_25775);
xnor U34529 (N_34529,N_26607,N_29826);
nand U34530 (N_34530,N_25943,N_25031);
and U34531 (N_34531,N_28958,N_28158);
xnor U34532 (N_34532,N_29614,N_28250);
and U34533 (N_34533,N_27406,N_26972);
nand U34534 (N_34534,N_26894,N_27708);
nand U34535 (N_34535,N_29385,N_27382);
or U34536 (N_34536,N_26441,N_27068);
nand U34537 (N_34537,N_26868,N_26256);
xnor U34538 (N_34538,N_27890,N_26578);
and U34539 (N_34539,N_25004,N_28606);
or U34540 (N_34540,N_27084,N_27967);
or U34541 (N_34541,N_28966,N_27732);
nand U34542 (N_34542,N_26369,N_25462);
nor U34543 (N_34543,N_26094,N_29808);
and U34544 (N_34544,N_26451,N_26988);
or U34545 (N_34545,N_29115,N_28423);
or U34546 (N_34546,N_27578,N_28248);
nand U34547 (N_34547,N_29200,N_26190);
nor U34548 (N_34548,N_29571,N_27922);
xor U34549 (N_34549,N_27863,N_26731);
and U34550 (N_34550,N_26948,N_28527);
xnor U34551 (N_34551,N_26650,N_25002);
nand U34552 (N_34552,N_29197,N_25152);
nand U34553 (N_34553,N_25467,N_28348);
or U34554 (N_34554,N_25914,N_28590);
xnor U34555 (N_34555,N_25316,N_26836);
and U34556 (N_34556,N_26370,N_29725);
or U34557 (N_34557,N_27199,N_25202);
nor U34558 (N_34558,N_29422,N_25184);
nor U34559 (N_34559,N_28584,N_29848);
or U34560 (N_34560,N_27784,N_26749);
nand U34561 (N_34561,N_26002,N_29298);
xor U34562 (N_34562,N_29022,N_27292);
nor U34563 (N_34563,N_26754,N_28715);
nand U34564 (N_34564,N_25395,N_28916);
and U34565 (N_34565,N_26784,N_26740);
xor U34566 (N_34566,N_29632,N_25511);
or U34567 (N_34567,N_29270,N_29975);
and U34568 (N_34568,N_28899,N_25851);
xor U34569 (N_34569,N_25598,N_28897);
xor U34570 (N_34570,N_25586,N_26621);
or U34571 (N_34571,N_27378,N_28719);
xnor U34572 (N_34572,N_25580,N_26418);
or U34573 (N_34573,N_27303,N_28711);
nor U34574 (N_34574,N_25897,N_28586);
or U34575 (N_34575,N_29952,N_29738);
xor U34576 (N_34576,N_28611,N_28573);
or U34577 (N_34577,N_29271,N_28688);
and U34578 (N_34578,N_28850,N_29350);
or U34579 (N_34579,N_29065,N_26956);
xnor U34580 (N_34580,N_25248,N_28488);
and U34581 (N_34581,N_28121,N_28983);
or U34582 (N_34582,N_28263,N_25137);
or U34583 (N_34583,N_25089,N_26391);
nor U34584 (N_34584,N_29398,N_25283);
nor U34585 (N_34585,N_27878,N_27394);
and U34586 (N_34586,N_25613,N_28498);
nand U34587 (N_34587,N_26457,N_26433);
xor U34588 (N_34588,N_26501,N_26744);
nor U34589 (N_34589,N_25764,N_25705);
xnor U34590 (N_34590,N_27281,N_29338);
nor U34591 (N_34591,N_27175,N_28732);
nor U34592 (N_34592,N_26515,N_26347);
or U34593 (N_34593,N_29689,N_25075);
or U34594 (N_34594,N_27979,N_27156);
or U34595 (N_34595,N_26644,N_26212);
nor U34596 (N_34596,N_28317,N_29757);
xor U34597 (N_34597,N_28862,N_26810);
nand U34598 (N_34598,N_28674,N_28093);
nor U34599 (N_34599,N_28724,N_29130);
and U34600 (N_34600,N_26103,N_29223);
and U34601 (N_34601,N_28148,N_29605);
or U34602 (N_34602,N_25034,N_26948);
xor U34603 (N_34603,N_26358,N_29325);
xnor U34604 (N_34604,N_28156,N_26949);
xor U34605 (N_34605,N_28882,N_26777);
nand U34606 (N_34606,N_29623,N_26296);
or U34607 (N_34607,N_29110,N_25326);
xnor U34608 (N_34608,N_27415,N_27087);
or U34609 (N_34609,N_28176,N_29432);
nor U34610 (N_34610,N_25253,N_26105);
nand U34611 (N_34611,N_29598,N_29007);
or U34612 (N_34612,N_28766,N_28421);
and U34613 (N_34613,N_27031,N_27510);
nand U34614 (N_34614,N_25020,N_29572);
or U34615 (N_34615,N_28577,N_29682);
nand U34616 (N_34616,N_27427,N_28331);
nor U34617 (N_34617,N_25302,N_26525);
nor U34618 (N_34618,N_28689,N_27093);
and U34619 (N_34619,N_26882,N_27422);
nor U34620 (N_34620,N_26160,N_28833);
xor U34621 (N_34621,N_25738,N_27874);
nand U34622 (N_34622,N_27264,N_28198);
or U34623 (N_34623,N_25942,N_27755);
or U34624 (N_34624,N_29818,N_29931);
xnor U34625 (N_34625,N_26970,N_29673);
xor U34626 (N_34626,N_29793,N_29632);
nand U34627 (N_34627,N_25781,N_25282);
nor U34628 (N_34628,N_27775,N_29720);
xnor U34629 (N_34629,N_29009,N_27510);
nand U34630 (N_34630,N_26985,N_25696);
nor U34631 (N_34631,N_27992,N_28105);
or U34632 (N_34632,N_25405,N_27673);
nand U34633 (N_34633,N_27887,N_27432);
or U34634 (N_34634,N_28064,N_27268);
xnor U34635 (N_34635,N_28975,N_27746);
or U34636 (N_34636,N_25714,N_29149);
nand U34637 (N_34637,N_27885,N_28904);
xnor U34638 (N_34638,N_26489,N_29157);
or U34639 (N_34639,N_29268,N_25680);
nand U34640 (N_34640,N_27590,N_28816);
nand U34641 (N_34641,N_27998,N_25796);
or U34642 (N_34642,N_28570,N_25500);
nand U34643 (N_34643,N_28594,N_28183);
nand U34644 (N_34644,N_25568,N_26802);
nor U34645 (N_34645,N_27900,N_28850);
nand U34646 (N_34646,N_29634,N_28838);
xnor U34647 (N_34647,N_27536,N_27361);
nor U34648 (N_34648,N_25779,N_27543);
and U34649 (N_34649,N_29801,N_27155);
xnor U34650 (N_34650,N_29684,N_25889);
nand U34651 (N_34651,N_27900,N_27535);
or U34652 (N_34652,N_25377,N_25026);
xor U34653 (N_34653,N_25861,N_25647);
nand U34654 (N_34654,N_28685,N_25487);
or U34655 (N_34655,N_26835,N_25598);
nand U34656 (N_34656,N_29903,N_25448);
or U34657 (N_34657,N_29084,N_25973);
nor U34658 (N_34658,N_26288,N_26970);
and U34659 (N_34659,N_25623,N_27683);
nand U34660 (N_34660,N_26235,N_28973);
or U34661 (N_34661,N_29875,N_26211);
nand U34662 (N_34662,N_28703,N_28185);
nor U34663 (N_34663,N_29385,N_26223);
nand U34664 (N_34664,N_28961,N_26130);
and U34665 (N_34665,N_29315,N_26139);
nor U34666 (N_34666,N_28822,N_25440);
nand U34667 (N_34667,N_28815,N_26351);
xor U34668 (N_34668,N_28432,N_26404);
or U34669 (N_34669,N_26698,N_25280);
nand U34670 (N_34670,N_25411,N_25719);
and U34671 (N_34671,N_28159,N_28396);
and U34672 (N_34672,N_29894,N_28563);
nor U34673 (N_34673,N_26260,N_26708);
or U34674 (N_34674,N_26537,N_26242);
nand U34675 (N_34675,N_25241,N_25527);
nand U34676 (N_34676,N_26253,N_29850);
or U34677 (N_34677,N_26374,N_27257);
nand U34678 (N_34678,N_28751,N_27321);
xnor U34679 (N_34679,N_27532,N_28185);
and U34680 (N_34680,N_27210,N_28214);
nand U34681 (N_34681,N_27953,N_26451);
nand U34682 (N_34682,N_28825,N_25331);
nor U34683 (N_34683,N_26326,N_25407);
or U34684 (N_34684,N_26277,N_25835);
nor U34685 (N_34685,N_29971,N_26611);
nor U34686 (N_34686,N_29563,N_27606);
or U34687 (N_34687,N_28733,N_27381);
or U34688 (N_34688,N_26459,N_25718);
nand U34689 (N_34689,N_28833,N_27425);
nor U34690 (N_34690,N_27158,N_28882);
xor U34691 (N_34691,N_26549,N_25500);
nand U34692 (N_34692,N_29178,N_27236);
nor U34693 (N_34693,N_28257,N_25480);
or U34694 (N_34694,N_25601,N_27718);
xor U34695 (N_34695,N_26391,N_29483);
and U34696 (N_34696,N_28390,N_26347);
or U34697 (N_34697,N_27001,N_29948);
xnor U34698 (N_34698,N_27221,N_27055);
nand U34699 (N_34699,N_26027,N_27273);
and U34700 (N_34700,N_25769,N_28616);
or U34701 (N_34701,N_29712,N_27136);
or U34702 (N_34702,N_27507,N_28889);
and U34703 (N_34703,N_25299,N_27323);
nand U34704 (N_34704,N_25978,N_29078);
xor U34705 (N_34705,N_26432,N_26533);
or U34706 (N_34706,N_26319,N_28948);
nor U34707 (N_34707,N_29420,N_25292);
nand U34708 (N_34708,N_28740,N_28085);
xor U34709 (N_34709,N_28302,N_26965);
xor U34710 (N_34710,N_26763,N_26180);
nor U34711 (N_34711,N_28273,N_26459);
or U34712 (N_34712,N_29338,N_25709);
or U34713 (N_34713,N_27501,N_27533);
and U34714 (N_34714,N_28403,N_26590);
and U34715 (N_34715,N_25052,N_29451);
xor U34716 (N_34716,N_29278,N_29842);
nand U34717 (N_34717,N_29547,N_27830);
or U34718 (N_34718,N_27604,N_26419);
nand U34719 (N_34719,N_29133,N_29435);
xnor U34720 (N_34720,N_25195,N_27491);
and U34721 (N_34721,N_27412,N_26654);
nor U34722 (N_34722,N_25951,N_29197);
nor U34723 (N_34723,N_25785,N_26131);
or U34724 (N_34724,N_27569,N_27733);
nor U34725 (N_34725,N_28085,N_26112);
nor U34726 (N_34726,N_28712,N_27582);
or U34727 (N_34727,N_29503,N_27756);
nand U34728 (N_34728,N_29315,N_29903);
nor U34729 (N_34729,N_28848,N_29118);
and U34730 (N_34730,N_25248,N_26843);
nor U34731 (N_34731,N_29759,N_25921);
nand U34732 (N_34732,N_28730,N_28701);
xor U34733 (N_34733,N_29764,N_25264);
nor U34734 (N_34734,N_29383,N_26986);
or U34735 (N_34735,N_29666,N_27424);
or U34736 (N_34736,N_27464,N_25443);
nor U34737 (N_34737,N_28472,N_29645);
nor U34738 (N_34738,N_28293,N_28883);
or U34739 (N_34739,N_28302,N_25513);
nor U34740 (N_34740,N_26728,N_29421);
or U34741 (N_34741,N_25080,N_25016);
nand U34742 (N_34742,N_29918,N_27931);
xor U34743 (N_34743,N_25605,N_25283);
and U34744 (N_34744,N_26917,N_25368);
and U34745 (N_34745,N_25983,N_28061);
and U34746 (N_34746,N_26760,N_25100);
and U34747 (N_34747,N_28091,N_27131);
nor U34748 (N_34748,N_25927,N_27812);
and U34749 (N_34749,N_28922,N_28752);
nor U34750 (N_34750,N_26925,N_25926);
and U34751 (N_34751,N_28858,N_25143);
nor U34752 (N_34752,N_25056,N_27588);
xnor U34753 (N_34753,N_26296,N_29962);
or U34754 (N_34754,N_29801,N_26468);
xor U34755 (N_34755,N_29226,N_25803);
nand U34756 (N_34756,N_26920,N_27957);
or U34757 (N_34757,N_26198,N_25506);
xnor U34758 (N_34758,N_25048,N_25629);
nor U34759 (N_34759,N_26506,N_27739);
nand U34760 (N_34760,N_25551,N_29107);
or U34761 (N_34761,N_29830,N_28785);
nand U34762 (N_34762,N_25911,N_28869);
or U34763 (N_34763,N_28704,N_27117);
xnor U34764 (N_34764,N_27578,N_29536);
or U34765 (N_34765,N_28140,N_28705);
or U34766 (N_34766,N_27938,N_25332);
xor U34767 (N_34767,N_28562,N_28273);
nand U34768 (N_34768,N_29280,N_28051);
nand U34769 (N_34769,N_28754,N_29489);
nor U34770 (N_34770,N_28568,N_28597);
xor U34771 (N_34771,N_25122,N_25809);
nand U34772 (N_34772,N_25243,N_28230);
and U34773 (N_34773,N_28327,N_25643);
xor U34774 (N_34774,N_28605,N_28968);
or U34775 (N_34775,N_25440,N_25088);
xor U34776 (N_34776,N_27478,N_26647);
xnor U34777 (N_34777,N_28147,N_26006);
or U34778 (N_34778,N_26886,N_27544);
nor U34779 (N_34779,N_28524,N_27533);
nor U34780 (N_34780,N_29656,N_27197);
or U34781 (N_34781,N_28944,N_26755);
nor U34782 (N_34782,N_27258,N_27887);
nand U34783 (N_34783,N_27096,N_25701);
xnor U34784 (N_34784,N_25271,N_29930);
xnor U34785 (N_34785,N_25811,N_25976);
nand U34786 (N_34786,N_25111,N_25138);
nor U34787 (N_34787,N_28755,N_27683);
nor U34788 (N_34788,N_27759,N_25818);
xor U34789 (N_34789,N_29175,N_26543);
and U34790 (N_34790,N_25173,N_27015);
nor U34791 (N_34791,N_27721,N_28661);
xnor U34792 (N_34792,N_29047,N_28372);
nor U34793 (N_34793,N_26127,N_25597);
and U34794 (N_34794,N_29055,N_28214);
xnor U34795 (N_34795,N_29694,N_29456);
nor U34796 (N_34796,N_25268,N_27556);
or U34797 (N_34797,N_27819,N_25854);
nor U34798 (N_34798,N_25275,N_25388);
and U34799 (N_34799,N_26166,N_27525);
or U34800 (N_34800,N_27982,N_27102);
xor U34801 (N_34801,N_27942,N_25332);
nor U34802 (N_34802,N_28867,N_29849);
nor U34803 (N_34803,N_26319,N_29418);
xor U34804 (N_34804,N_27660,N_28536);
nor U34805 (N_34805,N_27238,N_28418);
and U34806 (N_34806,N_27125,N_25174);
and U34807 (N_34807,N_26578,N_27688);
or U34808 (N_34808,N_29819,N_29778);
xnor U34809 (N_34809,N_27378,N_26269);
nand U34810 (N_34810,N_27304,N_26027);
or U34811 (N_34811,N_26784,N_29413);
or U34812 (N_34812,N_26310,N_29484);
or U34813 (N_34813,N_29774,N_29825);
and U34814 (N_34814,N_27915,N_26262);
nor U34815 (N_34815,N_26985,N_25443);
nor U34816 (N_34816,N_28227,N_28577);
xor U34817 (N_34817,N_25465,N_26201);
and U34818 (N_34818,N_28073,N_26524);
or U34819 (N_34819,N_27822,N_27279);
xor U34820 (N_34820,N_29896,N_27326);
xnor U34821 (N_34821,N_28612,N_26978);
and U34822 (N_34822,N_26510,N_29702);
and U34823 (N_34823,N_25017,N_28185);
nor U34824 (N_34824,N_25569,N_25983);
xor U34825 (N_34825,N_27321,N_29304);
and U34826 (N_34826,N_28257,N_27666);
xor U34827 (N_34827,N_26778,N_26580);
nor U34828 (N_34828,N_27990,N_27455);
nor U34829 (N_34829,N_26185,N_27241);
and U34830 (N_34830,N_26834,N_27737);
nand U34831 (N_34831,N_25199,N_28101);
nor U34832 (N_34832,N_27399,N_26472);
xnor U34833 (N_34833,N_29907,N_26166);
nand U34834 (N_34834,N_27908,N_28746);
nand U34835 (N_34835,N_27361,N_28500);
nor U34836 (N_34836,N_26747,N_28107);
or U34837 (N_34837,N_29210,N_25870);
nand U34838 (N_34838,N_26215,N_26944);
and U34839 (N_34839,N_28267,N_26321);
xnor U34840 (N_34840,N_25329,N_27296);
or U34841 (N_34841,N_25810,N_26149);
nor U34842 (N_34842,N_26849,N_29957);
xnor U34843 (N_34843,N_25868,N_28393);
nand U34844 (N_34844,N_27764,N_29827);
xnor U34845 (N_34845,N_26695,N_25781);
xnor U34846 (N_34846,N_29917,N_27902);
xor U34847 (N_34847,N_25172,N_25121);
and U34848 (N_34848,N_28249,N_27595);
xor U34849 (N_34849,N_29747,N_27139);
nor U34850 (N_34850,N_27154,N_25573);
xnor U34851 (N_34851,N_29527,N_27696);
nor U34852 (N_34852,N_28386,N_29402);
nor U34853 (N_34853,N_27025,N_28039);
or U34854 (N_34854,N_29858,N_26058);
or U34855 (N_34855,N_29987,N_29306);
xnor U34856 (N_34856,N_25174,N_28286);
or U34857 (N_34857,N_29803,N_28749);
nand U34858 (N_34858,N_28675,N_29014);
or U34859 (N_34859,N_25521,N_27117);
nor U34860 (N_34860,N_25577,N_28232);
nand U34861 (N_34861,N_25685,N_28375);
or U34862 (N_34862,N_27435,N_25676);
or U34863 (N_34863,N_25194,N_29799);
xor U34864 (N_34864,N_25740,N_25136);
and U34865 (N_34865,N_25744,N_27370);
nor U34866 (N_34866,N_28849,N_27019);
and U34867 (N_34867,N_27410,N_27707);
xor U34868 (N_34868,N_29862,N_28579);
nand U34869 (N_34869,N_28470,N_25473);
nor U34870 (N_34870,N_26944,N_29115);
nand U34871 (N_34871,N_27986,N_27909);
nand U34872 (N_34872,N_27705,N_28076);
or U34873 (N_34873,N_29663,N_29020);
or U34874 (N_34874,N_26930,N_27639);
nand U34875 (N_34875,N_28145,N_27511);
and U34876 (N_34876,N_25929,N_27971);
nor U34877 (N_34877,N_25618,N_27680);
and U34878 (N_34878,N_29983,N_29964);
xnor U34879 (N_34879,N_28585,N_25568);
xnor U34880 (N_34880,N_27604,N_28801);
nor U34881 (N_34881,N_28003,N_28047);
or U34882 (N_34882,N_29209,N_28287);
or U34883 (N_34883,N_29074,N_29056);
nand U34884 (N_34884,N_25307,N_29779);
or U34885 (N_34885,N_26153,N_27516);
nand U34886 (N_34886,N_29565,N_28259);
or U34887 (N_34887,N_29337,N_29096);
nor U34888 (N_34888,N_27617,N_29010);
nand U34889 (N_34889,N_25572,N_25896);
nor U34890 (N_34890,N_25837,N_29596);
nor U34891 (N_34891,N_27225,N_25369);
and U34892 (N_34892,N_27163,N_26763);
and U34893 (N_34893,N_27783,N_26013);
and U34894 (N_34894,N_27290,N_29461);
or U34895 (N_34895,N_25324,N_27320);
or U34896 (N_34896,N_25207,N_29528);
xnor U34897 (N_34897,N_26829,N_29536);
and U34898 (N_34898,N_27177,N_27407);
or U34899 (N_34899,N_25503,N_25140);
and U34900 (N_34900,N_26715,N_27646);
and U34901 (N_34901,N_27625,N_29299);
nand U34902 (N_34902,N_27178,N_27221);
nand U34903 (N_34903,N_29894,N_28048);
nand U34904 (N_34904,N_26609,N_27393);
nand U34905 (N_34905,N_26516,N_26607);
or U34906 (N_34906,N_28240,N_26065);
xor U34907 (N_34907,N_26469,N_26754);
xnor U34908 (N_34908,N_26538,N_25080);
nand U34909 (N_34909,N_25895,N_28675);
xnor U34910 (N_34910,N_29281,N_27910);
and U34911 (N_34911,N_25614,N_29755);
nand U34912 (N_34912,N_26364,N_26263);
nand U34913 (N_34913,N_25070,N_25307);
xnor U34914 (N_34914,N_28147,N_25510);
xor U34915 (N_34915,N_25500,N_28321);
or U34916 (N_34916,N_25838,N_26845);
xnor U34917 (N_34917,N_25508,N_26504);
xor U34918 (N_34918,N_29820,N_26943);
nor U34919 (N_34919,N_29373,N_28938);
or U34920 (N_34920,N_28590,N_28920);
or U34921 (N_34921,N_26105,N_25586);
and U34922 (N_34922,N_28900,N_28802);
xnor U34923 (N_34923,N_27523,N_29289);
nor U34924 (N_34924,N_28455,N_25244);
and U34925 (N_34925,N_28006,N_27927);
nand U34926 (N_34926,N_28432,N_26041);
and U34927 (N_34927,N_27178,N_25433);
nand U34928 (N_34928,N_27900,N_28476);
and U34929 (N_34929,N_28398,N_25461);
xor U34930 (N_34930,N_29563,N_28321);
or U34931 (N_34931,N_26921,N_28406);
nor U34932 (N_34932,N_27550,N_28987);
xnor U34933 (N_34933,N_25923,N_25710);
and U34934 (N_34934,N_27459,N_25079);
nor U34935 (N_34935,N_28707,N_26804);
nor U34936 (N_34936,N_28325,N_25053);
or U34937 (N_34937,N_25470,N_26065);
nor U34938 (N_34938,N_26917,N_28857);
or U34939 (N_34939,N_26935,N_29578);
and U34940 (N_34940,N_29206,N_27316);
nor U34941 (N_34941,N_26163,N_29807);
nand U34942 (N_34942,N_29639,N_25120);
xor U34943 (N_34943,N_25070,N_27217);
xnor U34944 (N_34944,N_29991,N_26420);
or U34945 (N_34945,N_27866,N_27123);
nand U34946 (N_34946,N_28540,N_28005);
xor U34947 (N_34947,N_28265,N_28721);
nor U34948 (N_34948,N_26018,N_29481);
xor U34949 (N_34949,N_29521,N_27802);
nor U34950 (N_34950,N_28132,N_27410);
xnor U34951 (N_34951,N_28545,N_26040);
and U34952 (N_34952,N_25218,N_29231);
and U34953 (N_34953,N_27734,N_29055);
and U34954 (N_34954,N_29713,N_25040);
or U34955 (N_34955,N_26956,N_26333);
and U34956 (N_34956,N_28830,N_28324);
nor U34957 (N_34957,N_25838,N_25486);
xnor U34958 (N_34958,N_27394,N_26540);
nor U34959 (N_34959,N_26345,N_29684);
nor U34960 (N_34960,N_25697,N_25040);
nor U34961 (N_34961,N_27508,N_27373);
or U34962 (N_34962,N_27719,N_28399);
nand U34963 (N_34963,N_26142,N_29725);
xor U34964 (N_34964,N_26242,N_25284);
or U34965 (N_34965,N_29447,N_26299);
nand U34966 (N_34966,N_27670,N_28277);
and U34967 (N_34967,N_25044,N_29977);
or U34968 (N_34968,N_25189,N_25592);
xnor U34969 (N_34969,N_25331,N_27480);
nand U34970 (N_34970,N_25466,N_26351);
nor U34971 (N_34971,N_27202,N_26453);
and U34972 (N_34972,N_26625,N_25504);
or U34973 (N_34973,N_29466,N_27877);
nand U34974 (N_34974,N_28801,N_28365);
or U34975 (N_34975,N_27982,N_25048);
or U34976 (N_34976,N_28091,N_28395);
nor U34977 (N_34977,N_28327,N_26621);
nand U34978 (N_34978,N_29627,N_26528);
xor U34979 (N_34979,N_27701,N_26156);
or U34980 (N_34980,N_25339,N_28210);
and U34981 (N_34981,N_27375,N_26025);
or U34982 (N_34982,N_29858,N_25228);
or U34983 (N_34983,N_27587,N_26524);
or U34984 (N_34984,N_26650,N_28476);
and U34985 (N_34985,N_28248,N_27591);
nand U34986 (N_34986,N_26953,N_28064);
or U34987 (N_34987,N_27212,N_28859);
nand U34988 (N_34988,N_28348,N_29104);
and U34989 (N_34989,N_26582,N_27660);
and U34990 (N_34990,N_29665,N_28692);
nand U34991 (N_34991,N_26421,N_26033);
or U34992 (N_34992,N_25552,N_26480);
or U34993 (N_34993,N_29401,N_26017);
nand U34994 (N_34994,N_25614,N_26624);
or U34995 (N_34995,N_27653,N_29157);
nor U34996 (N_34996,N_27718,N_29109);
nand U34997 (N_34997,N_26164,N_25759);
nand U34998 (N_34998,N_25578,N_27448);
nor U34999 (N_34999,N_25041,N_27643);
or U35000 (N_35000,N_34420,N_31316);
xnor U35001 (N_35001,N_33660,N_34870);
and U35002 (N_35002,N_30363,N_30646);
xnor U35003 (N_35003,N_33281,N_32498);
or U35004 (N_35004,N_34254,N_30305);
xor U35005 (N_35005,N_30522,N_31368);
nand U35006 (N_35006,N_34680,N_32708);
nor U35007 (N_35007,N_32354,N_31643);
and U35008 (N_35008,N_34506,N_30189);
xnor U35009 (N_35009,N_33226,N_32213);
nand U35010 (N_35010,N_34096,N_34628);
nor U35011 (N_35011,N_34522,N_33587);
or U35012 (N_35012,N_33804,N_33408);
or U35013 (N_35013,N_33740,N_31600);
nand U35014 (N_35014,N_31513,N_33510);
and U35015 (N_35015,N_32110,N_34659);
or U35016 (N_35016,N_30162,N_33410);
and U35017 (N_35017,N_33308,N_33617);
nand U35018 (N_35018,N_30784,N_30501);
xor U35019 (N_35019,N_30534,N_30215);
xnor U35020 (N_35020,N_34166,N_33359);
nor U35021 (N_35021,N_31649,N_32374);
or U35022 (N_35022,N_33870,N_33053);
nor U35023 (N_35023,N_30214,N_31914);
and U35024 (N_35024,N_31081,N_33060);
and U35025 (N_35025,N_30406,N_30995);
nand U35026 (N_35026,N_32794,N_34981);
nor U35027 (N_35027,N_34798,N_30874);
nor U35028 (N_35028,N_30124,N_34128);
xnor U35029 (N_35029,N_31650,N_34822);
nor U35030 (N_35030,N_32693,N_32990);
xor U35031 (N_35031,N_34307,N_31349);
and U35032 (N_35032,N_31337,N_33974);
and U35033 (N_35033,N_33718,N_32411);
or U35034 (N_35034,N_30936,N_32297);
or U35035 (N_35035,N_31446,N_32654);
nor U35036 (N_35036,N_33110,N_33954);
and U35037 (N_35037,N_30795,N_33078);
nand U35038 (N_35038,N_31925,N_30659);
nand U35039 (N_35039,N_32049,N_34066);
xor U35040 (N_35040,N_33861,N_30167);
xor U35041 (N_35041,N_34726,N_30509);
nor U35042 (N_35042,N_34860,N_32903);
and U35043 (N_35043,N_34531,N_30365);
and U35044 (N_35044,N_33691,N_34613);
nand U35045 (N_35045,N_33020,N_31669);
nor U35046 (N_35046,N_31211,N_34298);
or U35047 (N_35047,N_33825,N_31308);
or U35048 (N_35048,N_30230,N_30966);
nor U35049 (N_35049,N_30751,N_31348);
nand U35050 (N_35050,N_34791,N_34040);
nor U35051 (N_35051,N_32561,N_30578);
or U35052 (N_35052,N_31978,N_33620);
nand U35053 (N_35053,N_34683,N_32077);
and U35054 (N_35054,N_32384,N_34190);
or U35055 (N_35055,N_32955,N_31634);
or U35056 (N_35056,N_32657,N_33838);
or U35057 (N_35057,N_31757,N_32059);
nor U35058 (N_35058,N_30396,N_34521);
and U35059 (N_35059,N_31760,N_34963);
xor U35060 (N_35060,N_34421,N_34891);
or U35061 (N_35061,N_34487,N_31416);
or U35062 (N_35062,N_34734,N_30634);
and U35063 (N_35063,N_31226,N_30841);
and U35064 (N_35064,N_31155,N_33739);
and U35065 (N_35065,N_31780,N_31539);
nor U35066 (N_35066,N_34856,N_30604);
and U35067 (N_35067,N_34766,N_32375);
nand U35068 (N_35068,N_30603,N_33575);
nor U35069 (N_35069,N_32564,N_30750);
nand U35070 (N_35070,N_30173,N_34476);
and U35071 (N_35071,N_30451,N_31772);
nor U35072 (N_35072,N_33148,N_34896);
nor U35073 (N_35073,N_31454,N_33649);
xnor U35074 (N_35074,N_33550,N_32499);
nor U35075 (N_35075,N_32451,N_32505);
nand U35076 (N_35076,N_31241,N_32702);
and U35077 (N_35077,N_31924,N_33172);
nor U35078 (N_35078,N_32018,N_34480);
and U35079 (N_35079,N_30388,N_33700);
and U35080 (N_35080,N_31351,N_32777);
nand U35081 (N_35081,N_30954,N_34507);
xnor U35082 (N_35082,N_33049,N_32218);
xnor U35083 (N_35083,N_34888,N_30746);
or U35084 (N_35084,N_33250,N_34238);
nor U35085 (N_35085,N_30158,N_30419);
nand U35086 (N_35086,N_33480,N_31755);
xor U35087 (N_35087,N_33367,N_32134);
xnor U35088 (N_35088,N_32754,N_34611);
nand U35089 (N_35089,N_32229,N_33675);
xor U35090 (N_35090,N_33054,N_33569);
xor U35091 (N_35091,N_33249,N_33387);
or U35092 (N_35092,N_34403,N_34099);
and U35093 (N_35093,N_32423,N_32874);
and U35094 (N_35094,N_33628,N_32562);
nor U35095 (N_35095,N_33328,N_30007);
and U35096 (N_35096,N_32947,N_32207);
or U35097 (N_35097,N_32361,N_34219);
and U35098 (N_35098,N_33186,N_34829);
nor U35099 (N_35099,N_30071,N_33541);
xor U35100 (N_35100,N_31277,N_33361);
and U35101 (N_35101,N_31741,N_31897);
nor U35102 (N_35102,N_34097,N_33067);
xor U35103 (N_35103,N_31698,N_31611);
xor U35104 (N_35104,N_30211,N_33109);
and U35105 (N_35105,N_32902,N_31704);
or U35106 (N_35106,N_30528,N_32265);
nand U35107 (N_35107,N_31140,N_31710);
nand U35108 (N_35108,N_31342,N_31778);
or U35109 (N_35109,N_33439,N_32695);
nor U35110 (N_35110,N_32236,N_30182);
or U35111 (N_35111,N_34652,N_33576);
xnor U35112 (N_35112,N_30933,N_30793);
nor U35113 (N_35113,N_33158,N_32452);
and U35114 (N_35114,N_34795,N_33313);
nor U35115 (N_35115,N_30667,N_34644);
nor U35116 (N_35116,N_32492,N_34033);
and U35117 (N_35117,N_33670,N_33114);
or U35118 (N_35118,N_34707,N_33131);
nand U35119 (N_35119,N_32401,N_34002);
or U35120 (N_35120,N_34547,N_32344);
xnor U35121 (N_35121,N_31879,N_33748);
nor U35122 (N_35122,N_32295,N_31522);
nand U35123 (N_35123,N_32853,N_30823);
or U35124 (N_35124,N_30853,N_30693);
or U35125 (N_35125,N_34902,N_31633);
and U35126 (N_35126,N_33830,N_33210);
nand U35127 (N_35127,N_33205,N_32762);
or U35128 (N_35128,N_30168,N_33933);
or U35129 (N_35129,N_30135,N_33925);
nand U35130 (N_35130,N_34903,N_33556);
nor U35131 (N_35131,N_33236,N_34154);
nor U35132 (N_35132,N_33028,N_32007);
nand U35133 (N_35133,N_34148,N_33380);
xor U35134 (N_35134,N_32112,N_31125);
or U35135 (N_35135,N_34398,N_30160);
nand U35136 (N_35136,N_33837,N_32275);
and U35137 (N_35137,N_32830,N_31519);
xor U35138 (N_35138,N_31654,N_34253);
and U35139 (N_35139,N_32216,N_34647);
nor U35140 (N_35140,N_33859,N_31224);
or U35141 (N_35141,N_34520,N_31494);
nor U35142 (N_35142,N_32556,N_34075);
nand U35143 (N_35143,N_30974,N_34625);
xor U35144 (N_35144,N_34880,N_33521);
or U35145 (N_35145,N_31893,N_32628);
and U35146 (N_35146,N_33988,N_34646);
and U35147 (N_35147,N_34882,N_30371);
or U35148 (N_35148,N_34350,N_31439);
or U35149 (N_35149,N_33376,N_31196);
nand U35150 (N_35150,N_34354,N_33461);
or U35151 (N_35151,N_31253,N_32416);
or U35152 (N_35152,N_30929,N_34925);
nor U35153 (N_35153,N_32130,N_33713);
nand U35154 (N_35154,N_31657,N_30502);
nor U35155 (N_35155,N_31737,N_30343);
and U35156 (N_35156,N_34598,N_31424);
or U35157 (N_35157,N_32633,N_32997);
nand U35158 (N_35158,N_31338,N_33287);
or U35159 (N_35159,N_34965,N_34740);
nand U35160 (N_35160,N_34270,N_31181);
xor U35161 (N_35161,N_33145,N_31734);
nand U35162 (N_35162,N_31838,N_32826);
nor U35163 (N_35163,N_33143,N_30236);
nand U35164 (N_35164,N_33737,N_33621);
and U35165 (N_35165,N_32938,N_30468);
or U35166 (N_35166,N_30674,N_31303);
nor U35167 (N_35167,N_33991,N_34678);
xnor U35168 (N_35168,N_34784,N_34782);
or U35169 (N_35169,N_33447,N_30193);
nand U35170 (N_35170,N_34814,N_30309);
xor U35171 (N_35171,N_31302,N_30708);
xnor U35172 (N_35172,N_30876,N_30898);
nand U35173 (N_35173,N_30021,N_31688);
or U35174 (N_35174,N_32076,N_33432);
and U35175 (N_35175,N_30422,N_32811);
and U35176 (N_35176,N_30270,N_32696);
nor U35177 (N_35177,N_30505,N_30955);
nor U35178 (N_35178,N_32943,N_34679);
nor U35179 (N_35179,N_32648,N_33522);
nand U35180 (N_35180,N_31322,N_34473);
nand U35181 (N_35181,N_31639,N_33260);
and U35182 (N_35182,N_30152,N_32138);
and U35183 (N_35183,N_31222,N_31240);
nor U35184 (N_35184,N_31190,N_32540);
nor U35185 (N_35185,N_34789,N_31079);
nand U35186 (N_35186,N_34596,N_34376);
nor U35187 (N_35187,N_30572,N_32527);
nor U35188 (N_35188,N_30884,N_32873);
xor U35189 (N_35189,N_31333,N_34206);
and U35190 (N_35190,N_32918,N_31524);
and U35191 (N_35191,N_34702,N_33563);
and U35192 (N_35192,N_30112,N_34332);
nand U35193 (N_35193,N_32815,N_34998);
and U35194 (N_35194,N_33894,N_31373);
xnor U35195 (N_35195,N_33768,N_33581);
and U35196 (N_35196,N_31840,N_30552);
nand U35197 (N_35197,N_30932,N_34525);
xnor U35198 (N_35198,N_31483,N_33136);
nand U35199 (N_35199,N_33422,N_33906);
nor U35200 (N_35200,N_31213,N_30979);
or U35201 (N_35201,N_32132,N_32688);
xnor U35202 (N_35202,N_31395,N_30553);
nand U35203 (N_35203,N_34992,N_30353);
nor U35204 (N_35204,N_33775,N_33546);
xnor U35205 (N_35205,N_34145,N_34313);
nor U35206 (N_35206,N_30079,N_34057);
xnor U35207 (N_35207,N_31271,N_33070);
nor U35208 (N_35208,N_32140,N_30560);
or U35209 (N_35209,N_33772,N_32158);
nor U35210 (N_35210,N_33398,N_33914);
nor U35211 (N_35211,N_32175,N_32738);
and U35212 (N_35212,N_30299,N_34947);
and U35213 (N_35213,N_34936,N_31481);
xnor U35214 (N_35214,N_30130,N_33736);
nor U35215 (N_35215,N_33732,N_32093);
nor U35216 (N_35216,N_30510,N_33702);
nand U35217 (N_35217,N_30594,N_31580);
xnor U35218 (N_35218,N_32214,N_31396);
xor U35219 (N_35219,N_34738,N_32030);
or U35220 (N_35220,N_30777,N_34560);
nor U35221 (N_35221,N_32432,N_32820);
and U35222 (N_35222,N_33340,N_30986);
nand U35223 (N_35223,N_32987,N_33827);
and U35224 (N_35224,N_34899,N_33125);
or U35225 (N_35225,N_32792,N_33333);
nor U35226 (N_35226,N_34379,N_33468);
nor U35227 (N_35227,N_30856,N_32937);
xnor U35228 (N_35228,N_32819,N_31256);
nor U35229 (N_35229,N_30507,N_33626);
xor U35230 (N_35230,N_34732,N_33252);
nor U35231 (N_35231,N_31503,N_34442);
or U35232 (N_35232,N_32523,N_33195);
and U35233 (N_35233,N_31703,N_30450);
and U35234 (N_35234,N_30174,N_34811);
xnor U35235 (N_35235,N_34243,N_30592);
and U35236 (N_35236,N_31971,N_32259);
or U35237 (N_35237,N_31811,N_31281);
and U35238 (N_35238,N_32181,N_31629);
xor U35239 (N_35239,N_32424,N_31482);
xor U35240 (N_35240,N_32597,N_30383);
or U35241 (N_35241,N_32307,N_32317);
nor U35242 (N_35242,N_33448,N_33600);
or U35243 (N_35243,N_32033,N_32724);
xor U35244 (N_35244,N_33945,N_33265);
nand U35245 (N_35245,N_31341,N_31595);
or U35246 (N_35246,N_30110,N_33685);
or U35247 (N_35247,N_32889,N_30402);
xnor U35248 (N_35248,N_30779,N_31560);
or U35249 (N_35249,N_33355,N_34823);
or U35250 (N_35250,N_34052,N_34858);
xor U35251 (N_35251,N_34861,N_32258);
nor U35252 (N_35252,N_34172,N_31680);
or U35253 (N_35253,N_34278,N_32946);
nor U35254 (N_35254,N_34572,N_31844);
nor U35255 (N_35255,N_31788,N_30577);
nand U35256 (N_35256,N_34482,N_32274);
xor U35257 (N_35257,N_33593,N_31872);
nor U35258 (N_35258,N_34940,N_30725);
and U35259 (N_35259,N_30163,N_30889);
and U35260 (N_35260,N_31013,N_30350);
nand U35261 (N_35261,N_34935,N_32723);
xnor U35262 (N_35262,N_32553,N_30920);
or U35263 (N_35263,N_33025,N_31350);
and U35264 (N_35264,N_30097,N_34720);
nand U35265 (N_35265,N_32612,N_34109);
or U35266 (N_35266,N_32729,N_31541);
and U35267 (N_35267,N_31869,N_31896);
nand U35268 (N_35268,N_34750,N_31051);
or U35269 (N_35269,N_30220,N_30729);
nand U35270 (N_35270,N_33405,N_32766);
xor U35271 (N_35271,N_30653,N_34460);
xor U35272 (N_35272,N_33719,N_31974);
nor U35273 (N_35273,N_33013,N_30487);
and U35274 (N_35274,N_30797,N_31182);
nor U35275 (N_35275,N_33173,N_31983);
nor U35276 (N_35276,N_32653,N_34767);
and U35277 (N_35277,N_31045,N_32056);
and U35278 (N_35278,N_31770,N_31730);
nor U35279 (N_35279,N_33286,N_31834);
and U35280 (N_35280,N_32992,N_33790);
and U35281 (N_35281,N_34471,N_30761);
or U35282 (N_35282,N_33507,N_32771);
xor U35283 (N_35283,N_30030,N_32254);
xnor U35284 (N_35284,N_31156,N_34843);
or U35285 (N_35285,N_30680,N_33757);
nor U35286 (N_35286,N_34068,N_33377);
and U35287 (N_35287,N_30027,N_30748);
nor U35288 (N_35288,N_34853,N_34105);
nand U35289 (N_35289,N_34315,N_30626);
nand U35290 (N_35290,N_31374,N_32448);
or U35291 (N_35291,N_30831,N_30416);
nand U35292 (N_35292,N_33073,N_33912);
nand U35293 (N_35293,N_30414,N_32211);
nor U35294 (N_35294,N_34357,N_30232);
and U35295 (N_35295,N_32340,N_31769);
or U35296 (N_35296,N_33648,N_34859);
xnor U35297 (N_35297,N_33524,N_31832);
nor U35298 (N_35298,N_30605,N_32410);
or U35299 (N_35299,N_33969,N_33033);
or U35300 (N_35300,N_33977,N_30696);
nor U35301 (N_35301,N_33821,N_34526);
nor U35302 (N_35302,N_33088,N_34265);
and U35303 (N_35303,N_31484,N_32541);
and U35304 (N_35304,N_30666,N_31227);
and U35305 (N_35305,N_31728,N_30208);
xor U35306 (N_35306,N_31628,N_30311);
nor U35307 (N_35307,N_33623,N_33035);
nand U35308 (N_35308,N_31866,N_32781);
or U35309 (N_35309,N_31534,N_34378);
and U35310 (N_35310,N_31290,N_32196);
nor U35311 (N_35311,N_30991,N_33389);
xor U35312 (N_35312,N_33966,N_30905);
nor U35313 (N_35313,N_30833,N_31906);
xor U35314 (N_35314,N_33858,N_33193);
or U35315 (N_35315,N_31080,N_32663);
and U35316 (N_35316,N_31310,N_30316);
or U35317 (N_35317,N_30953,N_31176);
nand U35318 (N_35318,N_30170,N_33501);
nor U35319 (N_35319,N_33288,N_33463);
and U35320 (N_35320,N_30896,N_33533);
and U35321 (N_35321,N_31382,N_34592);
and U35322 (N_35322,N_33003,N_34504);
or U35323 (N_35323,N_34677,N_32146);
xnor U35324 (N_35324,N_30420,N_32098);
and U35325 (N_35325,N_34387,N_32571);
xor U35326 (N_35326,N_34836,N_33356);
nor U35327 (N_35327,N_30390,N_31535);
xnor U35328 (N_35328,N_32286,N_30977);
nor U35329 (N_35329,N_33095,N_30520);
or U35330 (N_35330,N_32253,N_34897);
or U35331 (N_35331,N_33061,N_33930);
xor U35332 (N_35332,N_31835,N_33674);
or U35333 (N_35333,N_33490,N_30873);
nand U35334 (N_35334,N_33818,N_32184);
or U35335 (N_35335,N_32817,N_32780);
xnor U35336 (N_35336,N_32062,N_33065);
xor U35337 (N_35337,N_30231,N_33893);
xnor U35338 (N_35338,N_31905,N_32460);
and U35339 (N_35339,N_32339,N_33416);
and U35340 (N_35340,N_33727,N_32271);
nand U35341 (N_35341,N_30964,N_31254);
nor U35342 (N_35342,N_33267,N_31544);
xor U35343 (N_35343,N_33393,N_32143);
xor U35344 (N_35344,N_32201,N_30591);
and U35345 (N_35345,N_30593,N_31588);
nor U35346 (N_35346,N_32659,N_31171);
nor U35347 (N_35347,N_31453,N_32441);
and U35348 (N_35348,N_32881,N_30957);
nor U35349 (N_35349,N_33197,N_31386);
nor U35350 (N_35350,N_34719,N_32869);
or U35351 (N_35351,N_32710,N_33781);
and U35352 (N_35352,N_34092,N_30678);
and U35353 (N_35353,N_33270,N_31391);
xor U35354 (N_35354,N_30331,N_30068);
or U35355 (N_35355,N_33348,N_30969);
nand U35356 (N_35356,N_32300,N_33424);
and U35357 (N_35357,N_32960,N_33445);
xnor U35358 (N_35358,N_30518,N_34001);
xor U35359 (N_35359,N_30769,N_31764);
nand U35360 (N_35360,N_33223,N_34612);
nor U35361 (N_35361,N_30772,N_31022);
xnor U35362 (N_35362,N_31257,N_34689);
nand U35363 (N_35363,N_31486,N_33697);
nor U35364 (N_35364,N_31773,N_34225);
nor U35365 (N_35365,N_32409,N_32249);
nor U35366 (N_35366,N_30151,N_31555);
and U35367 (N_35367,N_30890,N_33624);
nand U35368 (N_35368,N_33666,N_33519);
xnor U35369 (N_35369,N_33374,N_31317);
or U35370 (N_35370,N_34290,N_30098);
nand U35371 (N_35371,N_34517,N_30720);
or U35372 (N_35372,N_31742,N_30171);
and U35373 (N_35373,N_32769,N_32020);
or U35374 (N_35374,N_33758,N_34353);
and U35375 (N_35375,N_32831,N_34153);
and U35376 (N_35376,N_34907,N_32682);
or U35377 (N_35377,N_34283,N_30766);
xor U35378 (N_35378,N_32833,N_33705);
and U35379 (N_35379,N_34110,N_30651);
xor U35380 (N_35380,N_30218,N_32525);
and U35381 (N_35381,N_34852,N_30868);
nand U35382 (N_35382,N_33819,N_30559);
and U35383 (N_35383,N_32719,N_30527);
xnor U35384 (N_35384,N_34498,N_30357);
nor U35385 (N_35385,N_31060,N_32939);
nor U35386 (N_35386,N_34247,N_32805);
nand U35387 (N_35387,N_31249,N_30184);
nand U35388 (N_35388,N_33322,N_32978);
nor U35389 (N_35389,N_30845,N_33080);
or U35390 (N_35390,N_31236,N_32846);
nor U35391 (N_35391,N_34181,N_34863);
xor U35392 (N_35392,N_33651,N_34306);
xnor U35393 (N_35393,N_33560,N_31533);
and U35394 (N_35394,N_34175,N_30973);
and U35395 (N_35395,N_31419,N_34189);
or U35396 (N_35396,N_32728,N_31331);
and U35397 (N_35397,N_31738,N_30844);
nor U35398 (N_35398,N_31444,N_30556);
and U35399 (N_35399,N_33514,N_31507);
and U35400 (N_35400,N_30291,N_31845);
nor U35401 (N_35401,N_31426,N_31752);
nand U35402 (N_35402,N_32208,N_31987);
nor U35403 (N_35403,N_30069,N_34367);
or U35404 (N_35404,N_33085,N_30380);
and U35405 (N_35405,N_33745,N_34410);
xnor U35406 (N_35406,N_33037,N_34669);
nand U35407 (N_35407,N_34709,N_33509);
nand U35408 (N_35408,N_34342,N_32367);
xor U35409 (N_35409,N_34900,N_33228);
or U35410 (N_35410,N_31197,N_33315);
or U35411 (N_35411,N_33590,N_30899);
nand U35412 (N_35412,N_30425,N_31179);
xnor U35413 (N_35413,N_33245,N_30336);
nand U35414 (N_35414,N_31431,N_31665);
nand U35415 (N_35415,N_34366,N_31057);
xor U35416 (N_35416,N_31002,N_33665);
xor U35417 (N_35417,N_33400,N_30429);
nand U35418 (N_35418,N_32630,N_31745);
or U35419 (N_35419,N_32963,N_34042);
and U35420 (N_35420,N_34245,N_34848);
nor U35421 (N_35421,N_31242,N_34281);
or U35422 (N_35422,N_31946,N_30695);
nor U35423 (N_35423,N_31246,N_34733);
or U35424 (N_35424,N_31927,N_30012);
nor U35425 (N_35425,N_33905,N_31707);
xnor U35426 (N_35426,N_33454,N_33518);
or U35427 (N_35427,N_30632,N_33659);
or U35428 (N_35428,N_31420,N_34626);
or U35429 (N_35429,N_31286,N_32390);
xnor U35430 (N_35430,N_30878,N_34444);
nand U35431 (N_35431,N_33981,N_31550);
nor U35432 (N_35432,N_33471,N_34916);
nand U35433 (N_35433,N_31736,N_33196);
nand U35434 (N_35434,N_31437,N_32602);
nor U35435 (N_35435,N_32878,N_34515);
or U35436 (N_35436,N_33795,N_33201);
xnor U35437 (N_35437,N_30226,N_32369);
nor U35438 (N_35438,N_34323,N_34185);
and U35439 (N_35439,N_34474,N_30325);
and U35440 (N_35440,N_32879,N_32611);
nand U35441 (N_35441,N_30424,N_31149);
and U35442 (N_35442,N_30132,N_32035);
nand U35443 (N_35443,N_32109,N_33848);
or U35444 (N_35444,N_34781,N_33744);
nor U35445 (N_35445,N_33544,N_30004);
and U35446 (N_35446,N_33783,N_34402);
xor U35447 (N_35447,N_31212,N_32025);
nand U35448 (N_35448,N_31399,N_34587);
and U35449 (N_35449,N_30804,N_34890);
xnor U35450 (N_35450,N_33127,N_31393);
nor U35451 (N_35451,N_31123,N_31352);
xnor U35452 (N_35452,N_30972,N_34875);
and U35453 (N_35453,N_31911,N_30272);
or U35454 (N_35454,N_32117,N_31314);
nand U35455 (N_35455,N_33126,N_33999);
xnor U35456 (N_35456,N_30948,N_32776);
or U35457 (N_35457,N_30885,N_33268);
nand U35458 (N_35458,N_33618,N_32282);
xnor U35459 (N_35459,N_30257,N_31750);
or U35460 (N_35460,N_30564,N_30665);
or U35461 (N_35461,N_31418,N_32882);
nor U35462 (N_35462,N_32005,N_33984);
or U35463 (N_35463,N_32296,N_30032);
nor U35464 (N_35464,N_32187,N_30176);
or U35465 (N_35465,N_33135,N_31434);
nor U35466 (N_35466,N_31518,N_30718);
xor U35467 (N_35467,N_30862,N_30445);
or U35468 (N_35468,N_31229,N_30565);
nor U35469 (N_35469,N_31116,N_34168);
or U35470 (N_35470,N_32345,N_31613);
nand U35471 (N_35471,N_30723,N_34333);
nor U35472 (N_35472,N_34731,N_33742);
nor U35473 (N_35473,N_31711,N_30356);
nand U35474 (N_35474,N_34151,N_31756);
nand U35475 (N_35475,N_33259,N_30376);
xnor U35476 (N_35476,N_32660,N_34464);
nand U35477 (N_35477,N_32028,N_32359);
nor U35478 (N_35478,N_31111,N_34640);
nand U35479 (N_35479,N_32563,N_32980);
nor U35480 (N_35480,N_33489,N_34475);
or U35481 (N_35481,N_32590,N_32467);
nor U35482 (N_35482,N_34954,N_34501);
nand U35483 (N_35483,N_34576,N_30894);
nand U35484 (N_35484,N_34541,N_30865);
or U35485 (N_35485,N_33474,N_32970);
nand U35486 (N_35486,N_30842,N_32365);
xnor U35487 (N_35487,N_31546,N_33635);
and U35488 (N_35488,N_34761,N_33246);
and U35489 (N_35489,N_33189,N_31159);
xnor U35490 (N_35490,N_33849,N_30724);
nor U35491 (N_35491,N_32048,N_34113);
xor U35492 (N_35492,N_33256,N_32251);
and U35493 (N_35493,N_32012,N_32144);
and U35494 (N_35494,N_30512,N_32545);
nor U35495 (N_35495,N_34548,N_34991);
xnor U35496 (N_35496,N_32924,N_33929);
or U35497 (N_35497,N_31949,N_33238);
nor U35498 (N_35498,N_32736,N_32839);
xor U35499 (N_35499,N_34816,N_31120);
nand U35500 (N_35500,N_33892,N_34447);
nor U35501 (N_35501,N_31531,N_31394);
and U35502 (N_35502,N_33968,N_34840);
or U35503 (N_35503,N_32969,N_30105);
and U35504 (N_35504,N_34165,N_34282);
xnor U35505 (N_35505,N_32161,N_33435);
nor U35506 (N_35506,N_31950,N_30526);
and U35507 (N_35507,N_32320,N_31790);
nor U35508 (N_35508,N_32129,N_31076);
and U35509 (N_35509,N_33225,N_33199);
nand U35510 (N_35510,N_30664,N_34446);
nor U35511 (N_35511,N_32081,N_32362);
nand U35512 (N_35512,N_32044,N_33498);
nor U35513 (N_35513,N_33247,N_31712);
nor U35514 (N_35514,N_34005,N_32412);
and U35515 (N_35515,N_33478,N_30368);
xor U35516 (N_35516,N_31083,N_32318);
and U35517 (N_35517,N_34700,N_34018);
and U35518 (N_35518,N_31873,N_30233);
nand U35519 (N_35519,N_33050,N_33482);
xnor U35520 (N_35520,N_30337,N_30463);
and U35521 (N_35521,N_30555,N_32476);
or U35522 (N_35522,N_33891,N_33342);
nor U35523 (N_35523,N_31774,N_34682);
and U35524 (N_35524,N_31506,N_30539);
xnor U35525 (N_35525,N_32289,N_30655);
nand U35526 (N_35526,N_33952,N_30209);
and U35527 (N_35527,N_33975,N_31876);
and U35528 (N_35528,N_34104,N_34385);
and U35529 (N_35529,N_34792,N_31005);
and U35530 (N_35530,N_31427,N_33588);
and U35531 (N_35531,N_33133,N_31233);
or U35532 (N_35532,N_34242,N_33992);
or U35533 (N_35533,N_33167,N_31377);
nand U35534 (N_35534,N_30148,N_32616);
nor U35535 (N_35535,N_32192,N_32706);
nor U35536 (N_35536,N_34549,N_34509);
xnor U35537 (N_35537,N_31653,N_32000);
nor U35538 (N_35538,N_30827,N_31401);
nor U35539 (N_35539,N_33332,N_33351);
xor U35540 (N_35540,N_33995,N_33683);
nor U35541 (N_35541,N_31597,N_34374);
or U35542 (N_35542,N_31006,N_34911);
and U35543 (N_35543,N_34777,N_30775);
nor U35544 (N_35544,N_31685,N_30610);
nand U35545 (N_35545,N_33916,N_34915);
nand U35546 (N_35546,N_30558,N_33940);
and U35547 (N_35547,N_32971,N_33202);
or U35548 (N_35548,N_30490,N_33711);
and U35549 (N_35549,N_32417,N_33395);
nand U35550 (N_35550,N_33637,N_30541);
nand U35551 (N_35551,N_33753,N_31014);
nor U35552 (N_35552,N_30947,N_30949);
nor U35553 (N_35553,N_33960,N_32419);
and U35554 (N_35554,N_33536,N_32537);
nor U35555 (N_35555,N_33822,N_31509);
and U35556 (N_35556,N_30671,N_34953);
nor U35557 (N_35557,N_34770,N_32246);
nand U35558 (N_35558,N_31450,N_33093);
nand U35559 (N_35559,N_32691,N_30755);
and U35560 (N_35560,N_34978,N_30101);
xor U35561 (N_35561,N_32068,N_31158);
xor U35562 (N_35562,N_33484,N_31104);
xor U35563 (N_35563,N_30574,N_30597);
xor U35564 (N_35564,N_30378,N_31576);
and U35565 (N_35565,N_34204,N_30435);
nor U35566 (N_35566,N_31538,N_33399);
and U35567 (N_35567,N_31623,N_33475);
nor U35568 (N_35568,N_31883,N_30109);
and U35569 (N_35569,N_31325,N_31392);
and U35570 (N_35570,N_31473,N_33039);
nor U35571 (N_35571,N_31210,N_33077);
xnor U35572 (N_35572,N_33301,N_31478);
and U35573 (N_35573,N_33633,N_32999);
or U35574 (N_35574,N_33150,N_30658);
xor U35575 (N_35575,N_30990,N_33586);
xnor U35576 (N_35576,N_32336,N_31019);
and U35577 (N_35577,N_32245,N_32016);
or U35578 (N_35578,N_34755,N_32334);
xnor U35579 (N_35579,N_33881,N_33774);
and U35580 (N_35580,N_32647,N_30499);
and U35581 (N_35581,N_34215,N_33056);
and U35582 (N_35582,N_32935,N_34699);
or U35583 (N_35583,N_30752,N_32205);
nand U35584 (N_35584,N_31296,N_34466);
xor U35585 (N_35585,N_33561,N_33869);
or U35586 (N_35586,N_32023,N_31732);
nand U35587 (N_35587,N_32685,N_34090);
and U35588 (N_35588,N_34049,N_30458);
or U35589 (N_35589,N_34196,N_33803);
nor U35590 (N_35590,N_30840,N_30570);
or U35591 (N_35591,N_31789,N_33862);
nand U35592 (N_35592,N_33455,N_30460);
nor U35593 (N_35593,N_30201,N_32930);
xnor U35594 (N_35594,N_33696,N_31842);
and U35595 (N_35595,N_30623,N_30307);
nor U35596 (N_35596,N_33704,N_30010);
and U35597 (N_35597,N_34372,N_34050);
and U35598 (N_35598,N_34686,N_32588);
nand U35599 (N_35599,N_32893,N_33987);
xor U35600 (N_35600,N_32153,N_31063);
nor U35601 (N_35601,N_30320,N_32321);
or U35602 (N_35602,N_34081,N_31651);
nand U35603 (N_35603,N_32827,N_34234);
and U35604 (N_35604,N_33782,N_33850);
and U35605 (N_35605,N_34663,N_30319);
nor U35606 (N_35606,N_30237,N_31794);
nand U35607 (N_35607,N_34550,N_31345);
and U35608 (N_35608,N_34966,N_32917);
nand U35609 (N_35609,N_34842,N_32119);
or U35610 (N_35610,N_32669,N_34674);
nand U35611 (N_35611,N_33750,N_33609);
nand U35612 (N_35612,N_33627,N_33923);
xnor U35613 (N_35613,N_31828,N_30473);
nand U35614 (N_35614,N_31312,N_33187);
or U35615 (N_35615,N_31364,N_34544);
nor U35616 (N_35616,N_34664,N_30730);
nand U35617 (N_35617,N_33865,N_32619);
or U35618 (N_35618,N_33129,N_32420);
nand U35619 (N_35619,N_31365,N_33024);
nor U35620 (N_35620,N_30400,N_34538);
or U35621 (N_35621,N_32548,N_33951);
nand U35622 (N_35622,N_30489,N_30817);
xor U35623 (N_35623,N_31304,N_34924);
or U35624 (N_35624,N_34794,N_34573);
and U35625 (N_35625,N_31274,N_33253);
or U35626 (N_35626,N_34236,N_34457);
and U35627 (N_35627,N_30206,N_31846);
and U35628 (N_35628,N_31809,N_30087);
or U35629 (N_35629,N_33502,N_34467);
nand U35630 (N_35630,N_31954,N_34881);
or U35631 (N_35631,N_31008,N_32962);
nand U35632 (N_35632,N_31195,N_30581);
or U35633 (N_35633,N_30164,N_34650);
and U35634 (N_35634,N_34303,N_33773);
nand U35635 (N_35635,N_31178,N_34627);
nand U35636 (N_35636,N_31201,N_30428);
nor U35637 (N_35637,N_31353,N_30126);
nor U35638 (N_35638,N_33227,N_32209);
xor U35639 (N_35639,N_34006,N_30017);
or U35640 (N_35640,N_30029,N_30826);
nor U35641 (N_35641,N_31235,N_32624);
or U35642 (N_35642,N_34901,N_33345);
nor U35643 (N_35643,N_34443,N_31822);
and U35644 (N_35644,N_33528,N_31479);
or U35645 (N_35645,N_32454,N_34392);
and U35646 (N_35646,N_33883,N_30447);
xnor U35647 (N_35647,N_31678,N_31723);
nand U35648 (N_35648,N_32637,N_34519);
xnor U35649 (N_35649,N_34400,N_30641);
nor U35650 (N_35650,N_30219,N_30609);
and U35651 (N_35651,N_32155,N_30348);
and U35652 (N_35652,N_34894,N_32105);
or U35653 (N_35653,N_32646,N_34346);
nor U35654 (N_35654,N_32847,N_31232);
and U35655 (N_35655,N_33318,N_33098);
xor U35656 (N_35656,N_33993,N_34721);
nand U35657 (N_35657,N_32974,N_31763);
or U35658 (N_35658,N_33928,N_33128);
nor U35659 (N_35659,N_30346,N_33216);
or U35660 (N_35660,N_34273,N_34300);
xor U35661 (N_35661,N_31165,N_34763);
xor U35662 (N_35662,N_32793,N_32721);
and U35663 (N_35663,N_33299,N_32174);
nand U35664 (N_35664,N_34157,N_34182);
or U35665 (N_35665,N_31072,N_33362);
xnor U35666 (N_35666,N_34029,N_32075);
or U35667 (N_35667,N_31880,N_34162);
or U35668 (N_35668,N_32994,N_34232);
nand U35669 (N_35669,N_30614,N_34158);
or U35670 (N_35670,N_33787,N_31264);
xnor U35671 (N_35671,N_30516,N_32667);
and U35672 (N_35672,N_34320,N_34994);
nand U35673 (N_35673,N_31683,N_33169);
nand U35674 (N_35674,N_31850,N_32765);
and U35675 (N_35675,N_32171,N_33907);
xor U35676 (N_35676,N_34465,N_32844);
and U35677 (N_35677,N_33152,N_32818);
and U35678 (N_35678,N_33801,N_34778);
and U35679 (N_35679,N_31471,N_33272);
xnor U35680 (N_35680,N_34412,N_31169);
or U35681 (N_35681,N_31221,N_32024);
nor U35682 (N_35682,N_34432,N_33446);
and U35683 (N_35683,N_32915,N_34252);
nand U35684 (N_35684,N_30938,N_31340);
nor U35685 (N_35685,N_32579,N_31889);
xor U35686 (N_35686,N_30789,N_31656);
or U35687 (N_35687,N_34494,N_34437);
or U35688 (N_35688,N_33555,N_32399);
or U35689 (N_35689,N_32524,N_31278);
and U35690 (N_35690,N_32923,N_34383);
nor U35691 (N_35691,N_30524,N_30519);
nor U35692 (N_35692,N_32147,N_33284);
nor U35693 (N_35693,N_33203,N_34768);
xnor U35694 (N_35694,N_31442,N_31152);
xor U35695 (N_35695,N_33506,N_33373);
and U35696 (N_35696,N_34551,N_34931);
nor U35697 (N_35697,N_32623,N_30116);
or U35698 (N_35698,N_32900,N_31916);
xor U35699 (N_35699,N_34582,N_34174);
and U35700 (N_35700,N_30903,N_34964);
nor U35701 (N_35701,N_32601,N_33105);
nand U35702 (N_35702,N_32220,N_34929);
or U35703 (N_35703,N_30085,N_33994);
or U35704 (N_35704,N_33494,N_33450);
or U35705 (N_35705,N_34065,N_33092);
and U35706 (N_35706,N_31359,N_30888);
nor U35707 (N_35707,N_31843,N_30656);
nand U35708 (N_35708,N_30417,N_32787);
and U35709 (N_35709,N_32264,N_31529);
nand U35710 (N_35710,N_34136,N_32314);
or U35711 (N_35711,N_34046,N_32250);
and U35712 (N_35712,N_32639,N_31787);
xor U35713 (N_35713,N_31720,N_30550);
or U35714 (N_35714,N_31784,N_31376);
nand U35715 (N_35715,N_31430,N_34079);
nand U35716 (N_35716,N_34380,N_32233);
nor U35717 (N_35717,N_30985,N_30472);
or U35718 (N_35718,N_33321,N_30382);
xnor U35719 (N_35719,N_31570,N_33406);
nor U35720 (N_35720,N_33534,N_32989);
and U35721 (N_35721,N_30200,N_32223);
xnor U35722 (N_35722,N_32341,N_30533);
and U35723 (N_35723,N_34589,N_30044);
xnor U35724 (N_35724,N_31530,N_34553);
and U35725 (N_35725,N_33419,N_33008);
or U35726 (N_35726,N_30054,N_32488);
and U35727 (N_35727,N_30347,N_31614);
or U35728 (N_35728,N_30585,N_34552);
nand U35729 (N_35729,N_30877,N_34570);
xnor U35730 (N_35730,N_34448,N_31875);
nor U35731 (N_35731,N_34711,N_31958);
nand U35732 (N_35732,N_30916,N_30997);
nor U35733 (N_35733,N_34661,N_31715);
nand U35734 (N_35734,N_34008,N_30323);
xor U35735 (N_35735,N_33791,N_34343);
nand U35736 (N_35736,N_30293,N_31996);
and U35737 (N_35737,N_31184,N_32225);
or U35738 (N_35738,N_30015,N_34293);
nand U35739 (N_35739,N_34908,N_33611);
xnor U35740 (N_35740,N_31231,N_34645);
nand U35741 (N_35741,N_32876,N_32356);
xor U35742 (N_35742,N_34974,N_32584);
and U35743 (N_35743,N_31500,N_31260);
xor U35744 (N_35744,N_34280,N_33784);
nor U35745 (N_35745,N_30493,N_30308);
nand U35746 (N_35746,N_30704,N_30286);
xor U35747 (N_35747,N_33834,N_31956);
nand U35748 (N_35748,N_30009,N_32206);
xor U35749 (N_35749,N_31275,N_31370);
nand U35750 (N_35750,N_34462,N_32908);
or U35751 (N_35751,N_33271,N_31878);
or U35752 (N_35752,N_30271,N_34948);
and U35753 (N_35753,N_31099,N_34051);
nand U35754 (N_35754,N_32325,N_31170);
nand U35755 (N_35755,N_30248,N_31306);
xnor U35756 (N_35756,N_32311,N_32617);
xnor U35757 (N_35757,N_30557,N_30476);
and U35758 (N_35758,N_32949,N_33062);
nor U35759 (N_35759,N_32606,N_34969);
and U35760 (N_35760,N_30113,N_31920);
nor U35761 (N_35761,N_30367,N_33168);
or U35762 (N_35762,N_31262,N_34286);
and U35763 (N_35763,N_33604,N_30544);
or U35764 (N_35764,N_32269,N_31818);
nand U35765 (N_35765,N_33571,N_33241);
nand U35766 (N_35766,N_32471,N_31344);
or U35767 (N_35767,N_33817,N_33656);
xor U35768 (N_35768,N_30019,N_31777);
or U35769 (N_35769,N_33273,N_33014);
nor U35770 (N_35770,N_32092,N_31098);
nand U35771 (N_35771,N_32235,N_31646);
nor U35772 (N_35772,N_32408,N_31932);
or U35773 (N_35773,N_31825,N_30229);
or U35774 (N_35774,N_31164,N_32756);
nand U35775 (N_35775,N_32137,N_32227);
nor U35776 (N_35776,N_33155,N_33030);
xor U35777 (N_35777,N_32182,N_31380);
and U35778 (N_35778,N_31874,N_30301);
nand U35779 (N_35779,N_32901,N_34807);
xnor U35780 (N_35780,N_30895,N_30586);
xnor U35781 (N_35781,N_32594,N_33477);
or U35782 (N_35782,N_33512,N_32003);
and U35783 (N_35783,N_33597,N_33767);
nor U35784 (N_35784,N_34797,N_32718);
nor U35785 (N_35785,N_34694,N_31953);
nor U35786 (N_35786,N_31034,N_31462);
nand U35787 (N_35787,N_30542,N_31526);
or U35788 (N_35788,N_31388,N_31269);
xnor U35789 (N_35789,N_30759,N_31801);
nand U35790 (N_35790,N_33113,N_34648);
or U35791 (N_35791,N_31283,N_31892);
or U35792 (N_35792,N_32897,N_31785);
or U35793 (N_35793,N_32570,N_30048);
nor U35794 (N_35794,N_30692,N_34728);
and U35795 (N_35795,N_34369,N_33486);
nand U35796 (N_35796,N_30602,N_30764);
nor U35797 (N_35797,N_31990,N_30956);
and U35798 (N_35798,N_30511,N_30742);
or U35799 (N_35799,N_32324,N_33305);
xnor U35800 (N_35800,N_34806,N_30285);
nand U35801 (N_35801,N_32539,N_33926);
nor U35802 (N_35802,N_34451,N_33672);
nand U35803 (N_35803,N_31870,N_30339);
nor U35804 (N_35804,N_34317,N_30314);
xnor U35805 (N_35805,N_31599,N_30418);
nand U35806 (N_35806,N_32768,N_31065);
and U35807 (N_35807,N_31601,N_34671);
or U35808 (N_35808,N_34425,N_34240);
or U35809 (N_35809,N_32069,N_34787);
and U35810 (N_35810,N_33629,N_30401);
or U35811 (N_35811,N_32114,N_34932);
or U35812 (N_35812,N_33715,N_32124);
or U35813 (N_35813,N_31520,N_32198);
xor U35814 (N_35814,N_30262,N_30663);
nand U35815 (N_35815,N_34291,N_31860);
xor U35816 (N_35816,N_34803,N_32322);
and U35817 (N_35817,N_31686,N_34904);
or U35818 (N_35818,N_34656,N_32305);
and U35819 (N_35819,N_31107,N_33505);
xnor U35820 (N_35820,N_31970,N_34419);
xor U35821 (N_35821,N_30847,N_30508);
or U35822 (N_35822,N_30274,N_30062);
or U35823 (N_35823,N_30807,N_30922);
xor U35824 (N_35824,N_30901,N_31487);
and U35825 (N_35825,N_32516,N_32052);
nor U35826 (N_35826,N_33323,N_31795);
nand U35827 (N_35827,N_30255,N_30801);
or U35828 (N_35828,N_33956,N_30387);
xnor U35829 (N_35829,N_32529,N_32121);
xor U35830 (N_35830,N_31321,N_34438);
or U35831 (N_35831,N_33565,N_30675);
and U35832 (N_35832,N_30821,N_31863);
or U35833 (N_35833,N_34167,N_31583);
xnor U35834 (N_35834,N_32330,N_30298);
or U35835 (N_35835,N_31289,N_30945);
nor U35836 (N_35836,N_32368,N_33890);
xor U35837 (N_35837,N_32159,N_33650);
or U35838 (N_35838,N_33451,N_33843);
nand U35839 (N_35839,N_32142,N_30811);
or U35840 (N_35840,N_32575,N_33472);
nor U35841 (N_35841,N_33931,N_30466);
and U35842 (N_35842,N_34391,N_30386);
and U35843 (N_35843,N_34873,N_32921);
or U35844 (N_35844,N_33156,N_33137);
nor U35845 (N_35845,N_31168,N_33071);
or U35846 (N_35846,N_33963,N_32907);
and U35847 (N_35847,N_32748,N_33771);
nand U35848 (N_35848,N_34846,N_34790);
nand U35849 (N_35849,N_30033,N_33934);
and U35850 (N_35850,N_34164,N_31695);
xor U35851 (N_35851,N_31018,N_30210);
and U35852 (N_35852,N_32668,N_34546);
xor U35853 (N_35853,N_30037,N_32759);
and U35854 (N_35854,N_32133,N_31887);
nand U35855 (N_35855,N_31023,N_33051);
and U35856 (N_35856,N_30060,N_31354);
nand U35857 (N_35857,N_33545,N_31069);
and U35858 (N_35858,N_34276,N_30861);
nor U35859 (N_35859,N_33097,N_30479);
and U35860 (N_35860,N_31799,N_33112);
nand U35861 (N_35861,N_31556,N_33591);
xor U35862 (N_35862,N_31606,N_30143);
nor U35863 (N_35863,N_33679,N_33442);
or U35864 (N_35864,N_30944,N_30156);
nand U35865 (N_35865,N_33341,N_34226);
or U35866 (N_35866,N_34486,N_32627);
nor U35867 (N_35867,N_32681,N_33166);
or U35868 (N_35868,N_30606,N_30332);
xor U35869 (N_35869,N_33874,N_32470);
and U35870 (N_35870,N_31475,N_34718);
nor U35871 (N_35871,N_31671,N_32055);
and U35872 (N_35872,N_32022,N_30915);
xor U35873 (N_35873,N_30180,N_31536);
nor U35874 (N_35874,N_31046,N_34577);
nand U35875 (N_35875,N_31612,N_33671);
nor U35876 (N_35876,N_31323,N_34055);
or U35877 (N_35877,N_31937,N_32357);
or U35878 (N_35878,N_34163,N_33531);
and U35879 (N_35879,N_33619,N_32115);
nor U35880 (N_35880,N_34039,N_30354);
or U35881 (N_35881,N_34885,N_32480);
and U35882 (N_35882,N_34559,N_34328);
nor U35883 (N_35883,N_33537,N_32951);
nand U35884 (N_35884,N_34495,N_33190);
and U35885 (N_35885,N_33710,N_34337);
xor U35886 (N_35886,N_30077,N_30026);
or U35887 (N_35887,N_31058,N_31094);
or U35888 (N_35888,N_31681,N_30488);
nand U35889 (N_35889,N_34909,N_31975);
nand U35890 (N_35890,N_30342,N_30100);
or U35891 (N_35891,N_32822,N_32538);
or U35892 (N_35892,N_34297,N_32979);
nand U35893 (N_35893,N_32156,N_32170);
nand U35894 (N_35894,N_31962,N_31662);
nor U35895 (N_35895,N_31047,N_33785);
or U35896 (N_35896,N_33275,N_34714);
nor U35897 (N_35897,N_34041,N_30034);
or U35898 (N_35898,N_30222,N_30736);
xor U35899 (N_35899,N_34373,N_31144);
or U35900 (N_35900,N_33904,N_30258);
nor U35901 (N_35901,N_33654,N_32388);
nand U35902 (N_35902,N_33608,N_30498);
nor U35903 (N_35903,N_32393,N_33042);
nand U35904 (N_35904,N_32165,N_30228);
or U35905 (N_35905,N_30830,N_34122);
or U35906 (N_35906,N_33274,N_31700);
nor U35907 (N_35907,N_33188,N_34605);
and U35908 (N_35908,N_30934,N_32825);
and U35909 (N_35909,N_31078,N_31432);
and U35910 (N_35910,N_31816,N_34502);
or U35911 (N_35911,N_32266,N_32518);
and U35912 (N_35912,N_30735,N_31329);
nor U35913 (N_35913,N_32816,N_34413);
xor U35914 (N_35914,N_31068,N_34575);
nand U35915 (N_35915,N_34951,N_31248);
xnor U35916 (N_35916,N_33388,N_34919);
or U35917 (N_35917,N_33902,N_31919);
nand U35918 (N_35918,N_32533,N_33369);
and U35919 (N_35919,N_30192,N_33770);
nor U35920 (N_35920,N_31706,N_31900);
nand U35921 (N_35921,N_33047,N_30547);
nand U35922 (N_35922,N_30075,N_34093);
xnor U35923 (N_35923,N_32002,N_31867);
nand U35924 (N_35924,N_30776,N_32998);
xor U35925 (N_35925,N_31609,N_33350);
nand U35926 (N_35926,N_33181,N_30892);
or U35927 (N_35927,N_34892,N_34825);
nand U35928 (N_35928,N_30716,N_31705);
and U35929 (N_35929,N_31589,N_31668);
nand U35930 (N_35930,N_32450,N_33072);
xor U35931 (N_35931,N_33289,N_31687);
nor U35932 (N_35932,N_32919,N_33459);
xnor U35933 (N_35933,N_33329,N_30224);
xor U35934 (N_35934,N_34631,N_30503);
xor U35935 (N_35935,N_32644,N_34275);
nor U35936 (N_35936,N_31339,N_33456);
nand U35937 (N_35937,N_33302,N_31718);
and U35938 (N_35938,N_31573,N_30340);
and U35939 (N_35939,N_32398,N_30117);
nor U35940 (N_35940,N_34535,N_32332);
nand U35941 (N_35941,N_33217,N_31514);
nand U35942 (N_35942,N_32122,N_34832);
or U35943 (N_35943,N_30686,N_31796);
nand U35944 (N_35944,N_31406,N_34214);
xnor U35945 (N_35945,N_32983,N_33120);
or U35946 (N_35946,N_33103,N_30778);
nand U35947 (N_35947,N_30773,N_30334);
nor U35948 (N_35948,N_32796,N_30625);
xor U35949 (N_35949,N_31441,N_31559);
and U35950 (N_35950,N_31575,N_33087);
nand U35951 (N_35951,N_31948,N_32043);
or U35952 (N_35952,N_33612,N_30573);
and U35953 (N_35953,N_33276,N_33185);
nor U35954 (N_35954,N_30389,N_32449);
nor U35955 (N_35955,N_30303,N_34618);
xnor U35956 (N_35956,N_34622,N_33741);
nor U35957 (N_35957,N_32909,N_31250);
nor U35958 (N_35958,N_34765,N_34756);
xor U35959 (N_35959,N_33130,N_30803);
and U35960 (N_35960,N_33402,N_34578);
xor U35961 (N_35961,N_30370,N_31942);
and U35962 (N_35962,N_34889,N_33530);
xor U35963 (N_35963,N_32631,N_33317);
nand U35964 (N_35964,N_32240,N_33469);
xor U35965 (N_35965,N_33094,N_34497);
nand U35966 (N_35966,N_31059,N_34799);
xnor U35967 (N_35967,N_34545,N_31511);
nand U35968 (N_35968,N_32380,N_30362);
xnor U35969 (N_35969,N_31928,N_31829);
nand U35970 (N_35970,N_30300,N_30620);
and U35971 (N_35971,N_32824,N_32261);
nor U35972 (N_35972,N_34455,N_31410);
xnor U35973 (N_35973,N_30351,N_31126);
xnor U35974 (N_35974,N_34078,N_33368);
and U35975 (N_35975,N_30137,N_34198);
nand U35976 (N_35976,N_33209,N_34418);
and U35977 (N_35977,N_32532,N_33899);
xor U35978 (N_35978,N_34983,N_33630);
nand U35979 (N_35979,N_33961,N_31582);
nand U35980 (N_35980,N_32526,N_31754);
nor U35981 (N_35981,N_33391,N_33582);
or U35982 (N_35982,N_32116,N_33657);
nand U35983 (N_35983,N_30670,N_34724);
nand U35984 (N_35984,N_33122,N_32544);
nand U35985 (N_35985,N_30690,N_32609);
or U35986 (N_35986,N_33606,N_31282);
or U35987 (N_35987,N_33680,N_32551);
and U35988 (N_35988,N_32089,N_31061);
nand U35989 (N_35989,N_33622,N_30405);
nor U35990 (N_35990,N_33316,N_33607);
or U35991 (N_35991,N_33403,N_32701);
and U35992 (N_35992,N_34207,N_33497);
or U35993 (N_35993,N_33922,N_30981);
nand U35994 (N_35994,N_32203,N_32995);
nand U35995 (N_35995,N_34178,N_30814);
and U35996 (N_35996,N_31328,N_33875);
nor U35997 (N_35997,N_34308,N_30722);
xnor U35998 (N_35998,N_33568,N_32734);
xnor U35999 (N_35999,N_33343,N_31510);
and U36000 (N_36000,N_30629,N_30783);
nor U36001 (N_36001,N_33123,N_34301);
and U36002 (N_36002,N_33183,N_34530);
xnor U36003 (N_36003,N_30657,N_31933);
nor U36004 (N_36004,N_34044,N_32443);
or U36005 (N_36005,N_34607,N_31781);
or U36006 (N_36006,N_34063,N_32457);
xor U36007 (N_36007,N_33438,N_33645);
and U36008 (N_36008,N_32185,N_34382);
xor U36009 (N_36009,N_31833,N_31335);
nand U36010 (N_36010,N_33334,N_32517);
and U36011 (N_36011,N_31823,N_34362);
nor U36012 (N_36012,N_30563,N_33851);
or U36013 (N_36013,N_34684,N_33159);
nand U36014 (N_36014,N_33483,N_30297);
nor U36015 (N_36015,N_30040,N_33314);
xnor U36016 (N_36016,N_32107,N_33754);
xor U36017 (N_36017,N_32581,N_33610);
and U36018 (N_36018,N_34356,N_33040);
and U36019 (N_36019,N_32445,N_33806);
nor U36020 (N_36020,N_30096,N_31219);
nand U36021 (N_36021,N_34543,N_34188);
nor U36022 (N_36022,N_33292,N_33794);
nor U36023 (N_36023,N_31093,N_33743);
nor U36024 (N_36024,N_31553,N_31587);
or U36025 (N_36025,N_31505,N_33749);
nor U36026 (N_36026,N_32500,N_34309);
and U36027 (N_36027,N_33237,N_31786);
and U36028 (N_36028,N_31028,N_33985);
nand U36029 (N_36029,N_32573,N_32506);
nand U36030 (N_36030,N_34399,N_30099);
or U36031 (N_36031,N_33572,N_31997);
nand U36032 (N_36032,N_33937,N_32195);
nand U36033 (N_36033,N_33385,N_30682);
nor U36034 (N_36034,N_31119,N_32085);
or U36035 (N_36035,N_33300,N_31517);
nand U36036 (N_36036,N_33141,N_34961);
nand U36037 (N_36037,N_34237,N_30139);
and U36038 (N_36038,N_30444,N_33297);
xnor U36039 (N_36039,N_34872,N_30747);
nand U36040 (N_36040,N_33101,N_31121);
nand U36041 (N_36041,N_32395,N_34708);
nor U36042 (N_36042,N_34752,N_32404);
and U36043 (N_36043,N_33029,N_31272);
nand U36044 (N_36044,N_34124,N_33876);
nand U36045 (N_36045,N_33789,N_30310);
nor U36046 (N_36046,N_30941,N_31355);
xor U36047 (N_36047,N_31542,N_32933);
nor U36048 (N_36048,N_30913,N_33760);
nor U36049 (N_36049,N_31411,N_33017);
and U36050 (N_36050,N_32638,N_30975);
and U36051 (N_36051,N_34210,N_32547);
or U36052 (N_36052,N_30650,N_33485);
nor U36053 (N_36053,N_30448,N_30622);
nand U36054 (N_36054,N_30153,N_34493);
or U36055 (N_36055,N_33418,N_32858);
or U36056 (N_36056,N_32224,N_31957);
nor U36057 (N_36057,N_33414,N_33091);
xnor U36058 (N_36058,N_32886,N_34340);
nand U36059 (N_36059,N_33523,N_33358);
and U36060 (N_36060,N_30838,N_34583);
xor U36061 (N_36061,N_33090,N_34514);
nand U36062 (N_36062,N_34536,N_31082);
xor U36063 (N_36063,N_30423,N_34045);
nand U36064 (N_36064,N_31270,N_32343);
xor U36065 (N_36065,N_34256,N_31180);
or U36066 (N_36066,N_30806,N_31383);
or U36067 (N_36067,N_30195,N_31041);
xor U36068 (N_36068,N_31805,N_31696);
nor U36069 (N_36069,N_32642,N_31890);
xnor U36070 (N_36070,N_33192,N_30083);
nor U36071 (N_36071,N_34563,N_34993);
and U36072 (N_36072,N_34651,N_34867);
nor U36073 (N_36073,N_32950,N_32515);
nand U36074 (N_36074,N_30757,N_34255);
or U36075 (N_36075,N_31261,N_34921);
nand U36076 (N_36076,N_33263,N_32232);
nand U36077 (N_36077,N_32770,N_34195);
and U36078 (N_36078,N_32783,N_33001);
and U36079 (N_36079,N_30056,N_32484);
xor U36080 (N_36080,N_34950,N_32678);
xnor U36081 (N_36081,N_32377,N_30589);
or U36082 (N_36082,N_34453,N_31438);
nand U36083 (N_36083,N_33526,N_32015);
nand U36084 (N_36084,N_31768,N_30590);
xnor U36085 (N_36085,N_33844,N_34411);
nand U36086 (N_36086,N_32079,N_30612);
and U36087 (N_36087,N_34624,N_32582);
xnor U36088 (N_36088,N_34982,N_33473);
xnor U36089 (N_36089,N_32894,N_33430);
or U36090 (N_36090,N_31003,N_30599);
nand U36091 (N_36091,N_32465,N_33449);
nor U36092 (N_36092,N_34019,N_34527);
and U36093 (N_36093,N_30749,N_34459);
or U36094 (N_36094,N_34048,N_30630);
xnor U36095 (N_36095,N_31989,N_34800);
nor U36096 (N_36096,N_33638,N_34184);
or U36097 (N_36097,N_33979,N_30457);
xor U36098 (N_36098,N_34112,N_32006);
nor U36099 (N_36099,N_31977,N_34876);
xnor U36100 (N_36100,N_34760,N_34152);
nand U36101 (N_36101,N_32961,N_31898);
xor U36102 (N_36102,N_30091,N_34762);
nor U36103 (N_36103,N_34691,N_31854);
xnor U36104 (N_36104,N_34022,N_34608);
or U36105 (N_36105,N_31027,N_31968);
xnor U36106 (N_36106,N_33554,N_31961);
nand U36107 (N_36107,N_33578,N_31985);
xnor U36108 (N_36108,N_34952,N_32306);
and U36109 (N_36109,N_32810,N_33663);
or U36110 (N_36110,N_33725,N_33140);
and U36111 (N_36111,N_33852,N_30194);
nand U36112 (N_36112,N_34142,N_31037);
nand U36113 (N_36113,N_31367,N_32364);
nor U36114 (N_36114,N_31307,N_32360);
or U36115 (N_36115,N_32037,N_34116);
nor U36116 (N_36116,N_33924,N_32238);
nor U36117 (N_36117,N_33066,N_33832);
nand U36118 (N_36118,N_31435,N_34334);
nand U36119 (N_36119,N_33059,N_31288);
and U36120 (N_36120,N_30809,N_32131);
xor U36121 (N_36121,N_32899,N_34228);
or U36122 (N_36122,N_34512,N_33833);
nor U36123 (N_36123,N_30914,N_31234);
xor U36124 (N_36124,N_34730,N_32458);
nand U36125 (N_36125,N_31895,N_33692);
nor U36126 (N_36126,N_33936,N_31717);
or U36127 (N_36127,N_32113,N_33191);
xnor U36128 (N_36128,N_31466,N_34871);
xor U36129 (N_36129,N_32331,N_33658);
or U36130 (N_36130,N_32172,N_34257);
or U36131 (N_36131,N_30787,N_30958);
xor U36132 (N_36132,N_34511,N_31667);
nand U36133 (N_36133,N_31979,N_30183);
nand U36134 (N_36134,N_30078,N_33900);
and U36135 (N_36135,N_30234,N_34676);
nor U36136 (N_36136,N_34485,N_32982);
xor U36137 (N_36137,N_33344,N_33535);
xor U36138 (N_36138,N_30043,N_34011);
or U36139 (N_36139,N_30608,N_31443);
and U36140 (N_36140,N_34389,N_32413);
nand U36141 (N_36141,N_31545,N_30714);
nor U36142 (N_36142,N_32965,N_33733);
nand U36143 (N_36143,N_32510,N_30217);
nor U36144 (N_36144,N_33910,N_31610);
nor U36145 (N_36145,N_34038,N_34061);
or U36146 (N_36146,N_30681,N_30446);
and U36147 (N_36147,N_30252,N_32528);
and U36148 (N_36148,N_32248,N_32095);
nor U36149 (N_36149,N_31740,N_31347);
and U36150 (N_36150,N_31361,N_32389);
and U36151 (N_36151,N_34886,N_30728);
nand U36152 (N_36152,N_31216,N_30952);
or U36153 (N_36153,N_33433,N_33394);
and U36154 (N_36154,N_32656,N_33458);
xor U36155 (N_36155,N_32868,N_31871);
xor U36156 (N_36156,N_34864,N_32173);
or U36157 (N_36157,N_32543,N_34269);
or U36158 (N_36158,N_32725,N_32996);
nand U36159 (N_36159,N_32530,N_33515);
nand U36160 (N_36160,N_30377,N_31035);
xnor U36161 (N_36161,N_34960,N_33257);
nor U36162 (N_36162,N_31346,N_33411);
or U36163 (N_36163,N_30484,N_33764);
nand U36164 (N_36164,N_33160,N_32596);
xor U36165 (N_36165,N_32439,N_33840);
nor U36166 (N_36166,N_33816,N_32572);
nand U36167 (N_36167,N_34926,N_33309);
xnor U36168 (N_36168,N_31490,N_30159);
xor U36169 (N_36169,N_32578,N_31735);
nor U36170 (N_36170,N_34147,N_34140);
and U36171 (N_36171,N_31852,N_33652);
nand U36172 (N_36172,N_30187,N_31684);
nor U36173 (N_36173,N_33873,N_33579);
or U36174 (N_36174,N_31324,N_30415);
xor U36175 (N_36175,N_33492,N_31488);
nor U36176 (N_36176,N_31218,N_30461);
and U36177 (N_36177,N_34481,N_32436);
or U36178 (N_36178,N_32496,N_31073);
nand U36179 (N_36179,N_32070,N_30805);
xor U36180 (N_36180,N_33686,N_33540);
or U36181 (N_36181,N_34058,N_32036);
nor U36182 (N_36182,N_30049,N_33386);
xor U36183 (N_36183,N_30702,N_30154);
nor U36184 (N_36184,N_34114,N_34695);
nand U36185 (N_36185,N_31841,N_33631);
nor U36186 (N_36186,N_34404,N_30596);
or U36187 (N_36187,N_34458,N_33839);
and U36188 (N_36188,N_34773,N_34261);
and U36189 (N_36189,N_32774,N_30637);
nand U36190 (N_36190,N_30521,N_34743);
nor U36191 (N_36191,N_32106,N_31133);
xor U36192 (N_36192,N_33909,N_30059);
nor U36193 (N_36193,N_33218,N_34558);
or U36194 (N_36194,N_33577,N_31746);
nor U36195 (N_36195,N_31421,N_31143);
nor U36196 (N_36196,N_30022,N_33031);
nor U36197 (N_36197,N_32589,N_31205);
or U36198 (N_36198,N_33677,N_32920);
nand U36199 (N_36199,N_30221,N_34003);
and U36200 (N_36200,N_33941,N_33792);
or U36201 (N_36201,N_32760,N_32914);
or U36202 (N_36202,N_30042,N_34036);
xor U36203 (N_36203,N_31223,N_30689);
nand U36204 (N_36204,N_30203,N_32255);
xor U36205 (N_36205,N_30052,N_30950);
and U36206 (N_36206,N_34492,N_31187);
and U36207 (N_36207,N_33146,N_30442);
or U36208 (N_36208,N_30496,N_31031);
xnor U36209 (N_36209,N_33980,N_31563);
nor U36210 (N_36210,N_33614,N_30816);
and U36211 (N_36211,N_32665,N_34330);
nor U36212 (N_36212,N_31552,N_31000);
and U36213 (N_36213,N_30942,N_33104);
xor U36214 (N_36214,N_33662,N_31557);
and U36215 (N_36215,N_30492,N_32958);
or U36216 (N_36216,N_31921,N_32687);
xor U36217 (N_36217,N_31162,N_30999);
nor U36218 (N_36218,N_30598,N_30701);
nand U36219 (N_36219,N_33331,N_31150);
nor U36220 (N_36220,N_31413,N_33161);
and U36221 (N_36221,N_33699,N_32212);
xor U36222 (N_36222,N_34723,N_32041);
and U36223 (N_36223,N_30989,N_33375);
nor U36224 (N_36224,N_34704,N_33048);
xor U36225 (N_36225,N_32495,N_33594);
and U36226 (N_36226,N_32804,N_31847);
nand U36227 (N_36227,N_32194,N_32598);
nor U36228 (N_36228,N_31029,N_34917);
xor U36229 (N_36229,N_33681,N_32966);
or U36230 (N_36230,N_30545,N_34347);
nor U36231 (N_36231,N_30500,N_30638);
nand U36232 (N_36232,N_34997,N_34021);
nand U36233 (N_36233,N_33511,N_32580);
or U36234 (N_36234,N_33100,N_32268);
nor U36235 (N_36235,N_32689,N_34774);
and U36236 (N_36236,N_30276,N_31951);
xnor U36237 (N_36237,N_32703,N_34144);
nand U36238 (N_36238,N_34408,N_33082);
nand U36239 (N_36239,N_31214,N_33182);
and U36240 (N_36240,N_31981,N_33786);
and U36241 (N_36241,N_34865,N_32430);
xnor U36242 (N_36242,N_34996,N_33807);
and U36243 (N_36243,N_32535,N_32350);
and U36244 (N_36244,N_32391,N_32872);
xor U36245 (N_36245,N_33842,N_30212);
xnor U36246 (N_36246,N_30707,N_31857);
nor U36247 (N_36247,N_34468,N_33949);
and U36248 (N_36248,N_31263,N_31480);
or U36249 (N_36249,N_30754,N_33731);
xnor U36250 (N_36250,N_30575,N_33142);
nand U36251 (N_36251,N_31603,N_32150);
nand U36252 (N_36252,N_34972,N_33262);
xnor U36253 (N_36253,N_32381,N_31913);
nand U36254 (N_36254,N_33023,N_33324);
nand U36255 (N_36255,N_31015,N_32019);
nor U36256 (N_36256,N_31672,N_33005);
or U36257 (N_36257,N_31512,N_30504);
nand U36258 (N_36258,N_32509,N_32366);
xor U36259 (N_36259,N_31244,N_30911);
nor U36260 (N_36260,N_34985,N_31332);
or U36261 (N_36261,N_34363,N_33165);
nand U36262 (N_36262,N_32747,N_31727);
nor U36263 (N_36263,N_30883,N_32520);
or U36264 (N_36264,N_30028,N_32583);
nor U36265 (N_36265,N_31761,N_31708);
or U36266 (N_36266,N_30661,N_33021);
or U36267 (N_36267,N_30471,N_34197);
nand U36268 (N_36268,N_32103,N_32568);
nand U36269 (N_36269,N_30188,N_30635);
nor U36270 (N_36270,N_31627,N_30849);
or U36271 (N_36271,N_31381,N_34643);
or U36272 (N_36272,N_33559,N_31153);
and U36273 (N_36273,N_32797,N_30454);
and U36274 (N_36274,N_31762,N_32717);
or U36275 (N_36275,N_31699,N_31291);
nand U36276 (N_36276,N_30866,N_30935);
nand U36277 (N_36277,N_30344,N_34060);
or U36278 (N_36278,N_34318,N_30328);
and U36279 (N_36279,N_33012,N_34801);
or U36280 (N_36280,N_33057,N_34623);
nand U36281 (N_36281,N_31922,N_32422);
nor U36282 (N_36282,N_33069,N_32806);
and U36283 (N_36283,N_34134,N_30880);
nand U36284 (N_36284,N_31744,N_33153);
nand U36285 (N_36285,N_33895,N_34532);
nor U36286 (N_36286,N_33872,N_30404);
xnor U36287 (N_36287,N_32925,N_30057);
nor U36288 (N_36288,N_31001,N_33707);
nand U36289 (N_36289,N_33678,N_31009);
and U36290 (N_36290,N_32152,N_32379);
and U36291 (N_36291,N_34670,N_30925);
xnor U36292 (N_36292,N_30086,N_31865);
nand U36293 (N_36293,N_34742,N_32231);
or U36294 (N_36294,N_30881,N_31966);
and U36295 (N_36295,N_34681,N_34384);
nor U36296 (N_36296,N_31751,N_33064);
or U36297 (N_36297,N_30712,N_31131);
xor U36298 (N_36298,N_34108,N_33312);
or U36299 (N_36299,N_31592,N_32731);
nand U36300 (N_36300,N_34499,N_32786);
or U36301 (N_36301,N_34191,N_34883);
nand U36302 (N_36302,N_32262,N_30453);
and U36303 (N_36303,N_34034,N_32944);
nor U36304 (N_36304,N_30241,N_34271);
nor U36305 (N_36305,N_33034,N_31193);
xnor U36306 (N_36306,N_31644,N_31207);
or U36307 (N_36307,N_31499,N_30333);
nand U36308 (N_36308,N_34780,N_32190);
or U36309 (N_36309,N_30063,N_34813);
xor U36310 (N_36310,N_34345,N_32501);
xnor U36311 (N_36311,N_31300,N_31108);
nor U36312 (N_36312,N_34338,N_30011);
xor U36313 (N_36313,N_31020,N_32513);
nand U36314 (N_36314,N_31101,N_34898);
and U36315 (N_36315,N_34973,N_31775);
nand U36316 (N_36316,N_30398,N_32700);
nand U36317 (N_36317,N_30474,N_32910);
nor U36318 (N_36318,N_33491,N_33139);
and U36319 (N_36319,N_31793,N_30870);
and U36320 (N_36320,N_30771,N_31390);
and U36321 (N_36321,N_33721,N_32127);
nor U36322 (N_36322,N_32281,N_33669);
xor U36323 (N_36323,N_30984,N_32479);
or U36324 (N_36324,N_31032,N_32428);
nor U36325 (N_36325,N_33616,N_33866);
and U36326 (N_36326,N_32074,N_34854);
and U36327 (N_36327,N_32709,N_32083);
and U36328 (N_36328,N_33007,N_31802);
xnor U36329 (N_36329,N_32387,N_33413);
or U36330 (N_36330,N_33079,N_33261);
nand U36331 (N_36331,N_32730,N_34259);
nor U36332 (N_36332,N_34971,N_31888);
nand U36333 (N_36333,N_32298,N_34562);
and U36334 (N_36334,N_32383,N_30312);
or U36335 (N_36335,N_33011,N_32512);
xnor U36336 (N_36336,N_33668,N_34815);
or U36337 (N_36337,N_33694,N_33549);
and U36338 (N_36338,N_30832,N_31851);
nand U36339 (N_36339,N_34835,N_32911);
nand U36340 (N_36340,N_34837,N_30094);
xnor U36341 (N_36341,N_30114,N_32168);
xor U36342 (N_36342,N_31436,N_32522);
or U36343 (N_36343,N_32323,N_33756);
and U36344 (N_36344,N_30392,N_32239);
xor U36345 (N_36345,N_30381,N_34990);
nand U36346 (N_36346,N_31189,N_32763);
or U36347 (N_36347,N_30745,N_31591);
nand U36348 (N_36348,N_33206,N_34810);
xnor U36349 (N_36349,N_33958,N_33964);
xnor U36350 (N_36350,N_34007,N_30567);
xnor U36351 (N_36351,N_33955,N_34561);
nor U36352 (N_36352,N_34857,N_33584);
or U36353 (N_36353,N_33211,N_31679);
or U36354 (N_36354,N_34246,N_32219);
or U36355 (N_36355,N_30741,N_32857);
xor U36356 (N_36356,N_34581,N_30960);
or U36357 (N_36357,N_32038,N_34833);
nor U36358 (N_36358,N_34117,N_32333);
and U36359 (N_36359,N_31258,N_31400);
nand U36360 (N_36360,N_33815,N_30104);
and U36361 (N_36361,N_33179,N_33151);
nand U36362 (N_36362,N_32953,N_31166);
xor U36363 (N_36363,N_33996,N_31042);
or U36364 (N_36364,N_33959,N_32632);
nand U36365 (N_36365,N_30536,N_32593);
or U36366 (N_36366,N_34710,N_31491);
and U36367 (N_36367,N_30788,N_34094);
nor U36368 (N_36368,N_33306,N_30317);
xor U36369 (N_36369,N_32851,N_31154);
xnor U36370 (N_36370,N_31021,N_30269);
xnor U36371 (N_36371,N_34930,N_30937);
and U36372 (N_36372,N_33682,N_32247);
or U36373 (N_36373,N_30485,N_34657);
xor U36374 (N_36374,N_31186,N_30768);
nor U36375 (N_36375,N_31451,N_31881);
and U36376 (N_36376,N_30654,N_33552);
nand U36377 (N_36377,N_34100,N_32848);
nand U36378 (N_36378,N_34484,N_31468);
and U36379 (N_36379,N_32494,N_34722);
nor U36380 (N_36380,N_32679,N_32421);
nand U36381 (N_36381,N_30358,N_33213);
or U36382 (N_36382,N_31936,N_30093);
nand U36383 (N_36383,N_31593,N_33248);
xor U36384 (N_36384,N_33111,N_31554);
nand U36385 (N_36385,N_32014,N_30615);
or U36386 (N_36386,N_33599,N_30103);
or U36387 (N_36387,N_32304,N_33997);
and U36388 (N_36388,N_31215,N_34445);
nand U36389 (N_36389,N_30169,N_33431);
nor U36390 (N_36390,N_34171,N_32067);
or U36391 (N_36391,N_30106,N_34595);
and U36392 (N_36392,N_30717,N_33089);
nand U36393 (N_36393,N_34557,N_30263);
xnor U36394 (N_36394,N_32905,N_30624);
and U36395 (N_36395,N_34980,N_33009);
nand U36396 (N_36396,N_34054,N_33661);
and U36397 (N_36397,N_32625,N_34394);
nand U36398 (N_36398,N_31113,N_34665);
nor U36399 (N_36399,N_32464,N_30477);
nor U36400 (N_36400,N_30706,N_30523);
and U36401 (N_36401,N_33709,N_30835);
nand U36402 (N_36402,N_32791,N_30281);
nor U36403 (N_36403,N_31824,N_31298);
and U36404 (N_36404,N_32481,N_33543);
nand U36405 (N_36405,N_34987,N_34288);
nand U36406 (N_36406,N_34477,N_33296);
or U36407 (N_36407,N_31128,N_34274);
nand U36408 (N_36408,N_32189,N_33162);
and U36409 (N_36409,N_33499,N_34388);
nand U36410 (N_36410,N_34490,N_32039);
and U36411 (N_36411,N_33081,N_33327);
nand U36412 (N_36412,N_32502,N_32447);
and U36413 (N_36413,N_32635,N_33814);
xnor U36414 (N_36414,N_30073,N_33326);
and U36415 (N_36415,N_31127,N_32802);
nand U36416 (N_36416,N_32916,N_32082);
nor U36417 (N_36417,N_33639,N_33242);
and U36418 (N_36418,N_30828,N_33423);
or U36419 (N_36419,N_32795,N_32758);
and U36420 (N_36420,N_32836,N_31147);
nor U36421 (N_36421,N_32764,N_33542);
nor U36422 (N_36422,N_32072,N_33539);
nor U36423 (N_36423,N_32926,N_30839);
xnor U36424 (N_36424,N_34855,N_33769);
or U36425 (N_36425,N_33948,N_30202);
and U36426 (N_36426,N_31129,N_32348);
and U36427 (N_36427,N_34849,N_34976);
nand U36428 (N_36428,N_30408,N_30459);
nand U36429 (N_36429,N_34427,N_31693);
xor U36430 (N_36430,N_31581,N_33044);
nor U36431 (N_36431,N_33664,N_34594);
nor U36432 (N_36432,N_34296,N_30238);
and U36433 (N_36433,N_34083,N_34305);
xnor U36434 (N_36434,N_32686,N_33947);
nand U36435 (N_36435,N_34076,N_30798);
nand U36436 (N_36436,N_31175,N_31273);
or U36437 (N_36437,N_33831,N_32302);
and U36438 (N_36438,N_32288,N_30204);
nand U36439 (N_36439,N_32244,N_34590);
nor U36440 (N_36440,N_30628,N_32378);
or U36441 (N_36441,N_30138,N_31620);
nor U36442 (N_36442,N_30223,N_30120);
nor U36443 (N_36443,N_32620,N_32418);
and U36444 (N_36444,N_32912,N_31584);
nor U36445 (N_36445,N_32716,N_34630);
or U36446 (N_36446,N_33566,N_33513);
xnor U36447 (N_36447,N_34160,N_32135);
nor U36448 (N_36448,N_32801,N_31220);
or U36449 (N_36449,N_31090,N_33887);
nor U36450 (N_36450,N_30177,N_30774);
nor U36451 (N_36451,N_30065,N_30385);
xor U36452 (N_36452,N_31753,N_33371);
xor U36453 (N_36453,N_32342,N_31461);
and U36454 (N_36454,N_31673,N_32145);
nor U36455 (N_36455,N_30095,N_30700);
nand U36456 (N_36456,N_30245,N_34938);
nand U36457 (N_36457,N_33452,N_34962);
nor U36458 (N_36458,N_32064,N_31585);
nor U36459 (N_36459,N_34130,N_34314);
and U36460 (N_36460,N_30254,N_32779);
nor U36461 (N_36461,N_31808,N_30924);
and U36462 (N_36462,N_32234,N_34636);
xnor U36463 (N_36463,N_34106,N_31097);
nor U36464 (N_36464,N_34491,N_33118);
xor U36465 (N_36465,N_31719,N_30131);
nand U36466 (N_36466,N_34737,N_30782);
or U36467 (N_36467,N_31527,N_31086);
or U36468 (N_36468,N_30412,N_34289);
nor U36469 (N_36469,N_31326,N_34183);
nor U36470 (N_36470,N_32698,N_33116);
nand U36471 (N_36471,N_32301,N_34062);
and U36472 (N_36472,N_32073,N_34955);
and U36473 (N_36473,N_32552,N_30561);
nand U36474 (N_36474,N_32676,N_33915);
nand U36475 (N_36475,N_31980,N_30619);
xor U36476 (N_36476,N_33175,N_32309);
nand U36477 (N_36477,N_31709,N_30864);
nand U36478 (N_36478,N_33157,N_32337);
and U36479 (N_36479,N_30437,N_32312);
nand U36480 (N_36480,N_32870,N_34279);
or U36481 (N_36481,N_33868,N_32291);
nor U36482 (N_36482,N_30480,N_33846);
xor U36483 (N_36483,N_34311,N_31765);
and U36484 (N_36484,N_30595,N_31815);
xor U36485 (N_36485,N_30191,N_33885);
nor U36486 (N_36486,N_34395,N_30983);
or U36487 (N_36487,N_33058,N_32063);
or U36488 (N_36488,N_34943,N_34397);
nor U36489 (N_36489,N_32986,N_32865);
or U36490 (N_36490,N_30515,N_34287);
nor U36491 (N_36491,N_33735,N_34223);
nor U36492 (N_36492,N_34568,N_34588);
or U36493 (N_36493,N_34149,N_31814);
nand U36494 (N_36494,N_34818,N_32892);
or U36495 (N_36495,N_31412,N_31642);
xnor U36496 (N_36496,N_31092,N_30213);
and U36497 (N_36497,N_30394,N_34736);
nor U36498 (N_36498,N_32557,N_30530);
nand U36499 (N_36499,N_32883,N_33855);
or U36500 (N_36500,N_32283,N_34639);
or U36501 (N_36501,N_34187,N_33667);
xnor U36502 (N_36502,N_33360,N_31026);
nand U36503 (N_36503,N_33693,N_30691);
nor U36504 (N_36504,N_33853,N_31148);
nand U36505 (N_36505,N_30283,N_30993);
and U36506 (N_36506,N_34059,N_32478);
nor U36507 (N_36507,N_33503,N_34107);
or U36508 (N_36508,N_30115,N_33338);
and U36509 (N_36509,N_33019,N_30296);
or U36510 (N_36510,N_32431,N_33264);
nor U36511 (N_36511,N_33016,N_34675);
and U36512 (N_36512,N_34121,N_30588);
nand U36513 (N_36513,N_31976,N_30039);
xnor U36514 (N_36514,N_34000,N_34161);
xnor U36515 (N_36515,N_30127,N_30016);
and U36516 (N_36516,N_31632,N_32929);
xor U36517 (N_36517,N_31858,N_34866);
nor U36518 (N_36518,N_32273,N_32536);
nor U36519 (N_36519,N_31457,N_31384);
or U36520 (N_36520,N_30694,N_30506);
or U36521 (N_36521,N_31938,N_30349);
nand U36522 (N_36522,N_33043,N_34658);
xor U36523 (N_36523,N_34321,N_31722);
xnor U36524 (N_36524,N_30014,N_34461);
nand U36525 (N_36525,N_34847,N_34212);
or U36526 (N_36526,N_32279,N_33712);
or U36527 (N_36527,N_33295,N_31647);
and U36528 (N_36528,N_34716,N_31562);
or U36529 (N_36529,N_32237,N_31725);
xnor U36530 (N_36530,N_33500,N_34591);
or U36531 (N_36531,N_33099,N_34463);
xnor U36532 (N_36532,N_30259,N_30123);
nor U36533 (N_36533,N_30366,N_34024);
or U36534 (N_36534,N_34361,N_30978);
xnor U36535 (N_36535,N_30410,N_31915);
nand U36536 (N_36536,N_31605,N_33022);
or U36537 (N_36537,N_30165,N_30373);
or U36538 (N_36538,N_33854,N_34693);
and U36539 (N_36539,N_32504,N_30994);
nor U36540 (N_36540,N_30644,N_30852);
and U36541 (N_36541,N_33407,N_34975);
or U36542 (N_36542,N_32438,N_34757);
xnor U36543 (N_36543,N_30872,N_32169);
nand U36544 (N_36544,N_34186,N_30134);
or U36545 (N_36545,N_33982,N_34989);
xnor U36546 (N_36546,N_31405,N_31637);
xor U36547 (N_36547,N_30855,N_30711);
xnor U36548 (N_36548,N_32741,N_30050);
xnor U36549 (N_36549,N_31130,N_31891);
nand U36550 (N_36550,N_33170,N_30961);
nor U36551 (N_36551,N_34635,N_33625);
or U36552 (N_36552,N_34834,N_30921);
nor U36553 (N_36553,N_33443,N_33441);
or U36554 (N_36554,N_32141,N_33134);
nor U36555 (N_36555,N_32469,N_33943);
nand U36556 (N_36556,N_31362,N_30072);
or U36557 (N_36557,N_30092,N_34672);
nor U36558 (N_36558,N_33234,N_30288);
and U36559 (N_36559,N_33878,N_34934);
nand U36560 (N_36560,N_30051,N_31638);
nand U36561 (N_36561,N_34098,N_30497);
and U36562 (N_36562,N_32102,N_30443);
and U36563 (N_36563,N_33353,N_31826);
or U36564 (N_36564,N_32821,N_32614);
or U36565 (N_36565,N_34179,N_30867);
and U36566 (N_36566,N_32292,N_34754);
and U36567 (N_36567,N_32895,N_31567);
and U36568 (N_36568,N_32862,N_30584);
xor U36569 (N_36569,N_30968,N_34327);
or U36570 (N_36570,N_31903,N_34336);
nor U36571 (N_36571,N_33415,N_31160);
nor U36572 (N_36572,N_33701,N_32319);
or U36573 (N_36573,N_30455,N_30375);
and U36574 (N_36574,N_34138,N_30791);
nand U36575 (N_36575,N_31103,N_34928);
and U36576 (N_36576,N_33776,N_34133);
nor U36577 (N_36577,N_34884,N_32487);
nor U36578 (N_36578,N_31049,N_30850);
or U36579 (N_36579,N_34331,N_30379);
xnor U36580 (N_36580,N_30002,N_32692);
xnor U36581 (N_36581,N_34103,N_32108);
or U36582 (N_36582,N_30639,N_32277);
and U36583 (N_36583,N_30205,N_33278);
nor U36584 (N_36584,N_31064,N_32587);
or U36585 (N_36585,N_31052,N_30035);
xor U36586 (N_36586,N_32118,N_31142);
or U36587 (N_36587,N_32125,N_30001);
nor U36588 (N_36588,N_32403,N_33144);
nand U36589 (N_36589,N_33320,N_32163);
or U36590 (N_36590,N_33282,N_34653);
nor U36591 (N_36591,N_34759,N_31191);
xor U36592 (N_36592,N_34436,N_34221);
or U36593 (N_36593,N_31343,N_30280);
nand U36594 (N_36594,N_31313,N_33564);
nor U36595 (N_36595,N_30822,N_33428);
or U36596 (N_36596,N_34325,N_32652);
nor U36597 (N_36597,N_31558,N_31209);
xnor U36598 (N_36598,N_33184,N_31967);
nand U36599 (N_36599,N_31036,N_31908);
nand U36600 (N_36600,N_33283,N_33346);
and U36601 (N_36601,N_32210,N_33277);
or U36602 (N_36602,N_34200,N_32456);
xnor U36603 (N_36603,N_34906,N_32803);
xor U36604 (N_36604,N_34771,N_31713);
xnor U36605 (N_36605,N_34095,N_32661);
nor U36606 (N_36606,N_30292,N_30304);
xor U36607 (N_36607,N_30239,N_30897);
nor U36608 (N_36608,N_30971,N_33204);
nand U36609 (N_36609,N_34071,N_33052);
or U36610 (N_36610,N_32313,N_30546);
or U36611 (N_36611,N_32094,N_32252);
or U36612 (N_36612,N_34727,N_31702);
nor U36613 (N_36613,N_31515,N_34285);
xnor U36614 (N_36614,N_30289,N_33828);
and U36615 (N_36615,N_30698,N_34119);
and U36616 (N_36616,N_34424,N_30013);
nand U36617 (N_36617,N_30697,N_31038);
nand U36618 (N_36618,N_30469,N_34838);
or U36619 (N_36619,N_31689,N_34662);
nor U36620 (N_36620,N_30196,N_30677);
and U36621 (N_36621,N_31792,N_34263);
and U36622 (N_36622,N_33354,N_34025);
nand U36623 (N_36623,N_33255,N_33684);
nor U36624 (N_36624,N_30341,N_30185);
or U36625 (N_36625,N_34621,N_30287);
nor U36626 (N_36626,N_32164,N_32991);
and U36627 (N_36627,N_34586,N_33219);
and U36628 (N_36628,N_34349,N_34629);
xnor U36629 (N_36629,N_34009,N_32789);
or U36630 (N_36630,N_32845,N_30141);
and U36631 (N_36631,N_32626,N_33826);
and U36632 (N_36632,N_34251,N_34074);
or U36633 (N_36633,N_31963,N_33041);
and U36634 (N_36634,N_30046,N_32011);
and U36635 (N_36635,N_31204,N_32931);
and U36636 (N_36636,N_30465,N_31899);
or U36637 (N_36637,N_34705,N_33726);
or U36638 (N_36638,N_32672,N_32859);
and U36639 (N_36639,N_34352,N_32809);
nor U36640 (N_36640,N_31305,N_34649);
nor U36641 (N_36641,N_34250,N_30668);
and U36642 (N_36642,N_33083,N_32945);
nand U36643 (N_36643,N_31659,N_33780);
nand U36644 (N_36644,N_33690,N_30440);
and U36645 (N_36645,N_32891,N_32664);
xnor U36646 (N_36646,N_31660,N_34026);
xnor U36647 (N_36647,N_34428,N_31885);
xnor U36648 (N_36648,N_31523,N_32386);
or U36649 (N_36649,N_31472,N_34537);
nand U36650 (N_36650,N_34812,N_30335);
or U36651 (N_36651,N_30900,N_33171);
and U36652 (N_36652,N_34082,N_31238);
and U36653 (N_36653,N_30128,N_31676);
and U36654 (N_36654,N_30108,N_32091);
xnor U36655 (N_36655,N_32160,N_32674);
xor U36656 (N_36656,N_34450,N_30441);
xnor U36657 (N_36657,N_31663,N_33293);
nor U36658 (N_36658,N_30767,N_31024);
xnor U36659 (N_36659,N_34266,N_34879);
and U36660 (N_36660,N_31403,N_30662);
and U36661 (N_36661,N_30763,N_33002);
and U36662 (N_36662,N_34913,N_31050);
nor U36663 (N_36663,N_32566,N_34159);
nand U36664 (N_36664,N_33194,N_30430);
nor U36665 (N_36665,N_31463,N_34802);
nor U36666 (N_36666,N_33558,N_34304);
xor U36667 (N_36667,N_30456,N_34821);
and U36668 (N_36668,N_33689,N_31357);
and U36669 (N_36669,N_33106,N_32226);
and U36670 (N_36670,N_32290,N_30330);
nand U36671 (N_36671,N_30261,N_30243);
nand U36672 (N_36672,N_31566,N_34729);
nand U36673 (N_36673,N_32021,N_32276);
and U36674 (N_36674,N_31167,N_33285);
nand U36675 (N_36675,N_31292,N_34135);
xnor U36676 (N_36676,N_34877,N_33779);
and U36677 (N_36677,N_33751,N_32554);
and U36678 (N_36678,N_32849,N_30607);
nand U36679 (N_36679,N_30600,N_32788);
xnor U36680 (N_36680,N_34845,N_32752);
or U36681 (N_36681,N_30495,N_31402);
nor U36682 (N_36682,N_33467,N_34574);
nand U36683 (N_36683,N_32521,N_32270);
and U36684 (N_36684,N_34819,N_31694);
nand U36685 (N_36685,N_31203,N_34023);
nor U36686 (N_36686,N_31947,N_31371);
or U36687 (N_36687,N_34776,N_34415);
nor U36688 (N_36688,N_30399,N_31363);
and U36689 (N_36689,N_32629,N_33304);
nand U36690 (N_36690,N_31941,N_31991);
and U36691 (N_36691,N_34115,N_31039);
xnor U36692 (N_36692,N_30119,N_30965);
and U36693 (N_36693,N_31901,N_32508);
and U36694 (N_36694,N_34850,N_32397);
or U36695 (N_36695,N_34010,N_32497);
nor U36696 (N_36696,N_34264,N_32670);
and U36697 (N_36697,N_33045,N_34359);
nor U36698 (N_36698,N_30996,N_34920);
and U36699 (N_36699,N_30982,N_30517);
and U36700 (N_36700,N_31993,N_30543);
nor U36701 (N_36701,N_32243,N_34749);
nor U36702 (N_36702,N_30322,N_30136);
xnor U36703 (N_36703,N_30282,N_31456);
nand U36704 (N_36704,N_34933,N_30843);
or U36705 (N_36705,N_31276,N_34216);
xnor U36706 (N_36706,N_33601,N_32376);
nand U36707 (N_36707,N_33653,N_34633);
nor U36708 (N_36708,N_34335,N_31010);
nand U36709 (N_36709,N_30727,N_31016);
nand U36710 (N_36710,N_34748,N_32088);
nor U36711 (N_36711,N_32928,N_32046);
xor U36712 (N_36712,N_32812,N_32599);
nand U36713 (N_36713,N_33466,N_30846);
nor U36714 (N_36714,N_32607,N_34439);
nor U36715 (N_36715,N_33880,N_33465);
or U36716 (N_36716,N_34358,N_30820);
xnor U36717 (N_36717,N_33812,N_30427);
xnor U36718 (N_36718,N_31604,N_30082);
nor U36719 (N_36719,N_34556,N_31379);
and U36720 (N_36720,N_34203,N_30551);
and U36721 (N_36721,N_33867,N_30066);
and U36722 (N_36722,N_31551,N_31135);
nor U36723 (N_36723,N_30739,N_31831);
nor U36724 (N_36724,N_32565,N_30731);
and U36725 (N_36725,N_33970,N_31327);
xnor U36726 (N_36726,N_31011,N_30576);
nand U36727 (N_36727,N_30329,N_30685);
or U36728 (N_36728,N_32090,N_34329);
or U36729 (N_36729,N_31071,N_32294);
nand U36730 (N_36730,N_32191,N_33174);
xnor U36731 (N_36731,N_33349,N_33761);
xnor U36732 (N_36732,N_31830,N_34213);
xor U36733 (N_36733,N_34229,N_33927);
or U36734 (N_36734,N_31372,N_32316);
nand U36735 (N_36735,N_31767,N_34685);
xnor U36736 (N_36736,N_30819,N_34579);
nand U36737 (N_36737,N_30434,N_30568);
nor U36738 (N_36738,N_34470,N_34564);
nand U36739 (N_36739,N_31910,N_34841);
and U36740 (N_36740,N_31640,N_30537);
nand U36741 (N_36741,N_32732,N_34430);
and U36742 (N_36742,N_30756,N_34102);
or U36743 (N_36743,N_34230,N_30481);
nand U36744 (N_36744,N_32890,N_30792);
nor U36745 (N_36745,N_32267,N_31239);
or U36746 (N_36746,N_33337,N_34958);
xor U36747 (N_36747,N_31655,N_31040);
nor U36748 (N_36748,N_30360,N_30302);
xor U36749 (N_36749,N_30923,N_31474);
or U36750 (N_36750,N_30554,N_32680);
nor U36751 (N_36751,N_31397,N_30970);
xor U36752 (N_36752,N_32772,N_32177);
nor U36753 (N_36753,N_30726,N_33436);
or U36754 (N_36754,N_31504,N_30733);
and U36755 (N_36755,N_34942,N_30369);
nand U36756 (N_36756,N_31982,N_33796);
nor U36757 (N_36757,N_30294,N_32546);
or U36758 (N_36758,N_32188,N_34406);
xor U36759 (N_36759,N_33917,N_30470);
and U36760 (N_36760,N_31428,N_34483);
or U36761 (N_36761,N_31972,N_33723);
and U36762 (N_36762,N_34111,N_32051);
nand U36763 (N_36763,N_30859,N_33311);
xnor U36764 (N_36764,N_34073,N_33642);
or U36765 (N_36765,N_32808,N_33655);
or U36766 (N_36766,N_30393,N_32799);
or U36767 (N_36767,N_31615,N_34496);
and U36768 (N_36768,N_33462,N_30181);
nand U36769 (N_36769,N_34922,N_30256);
or U36770 (N_36770,N_32942,N_31579);
and U36771 (N_36771,N_33673,N_34150);
or U36772 (N_36772,N_32303,N_33919);
nor U36773 (N_36773,N_32755,N_30943);
nor U36774 (N_36774,N_32355,N_30125);
nor U36775 (N_36775,N_30491,N_30102);
and U36776 (N_36776,N_31336,N_30467);
nand U36777 (N_36777,N_34615,N_31208);
xor U36778 (N_36778,N_32735,N_31423);
or U36779 (N_36779,N_33240,N_33946);
or U36780 (N_36780,N_33027,N_33763);
nor U36781 (N_36781,N_31782,N_31330);
nor U36782 (N_36782,N_30327,N_31548);
or U36783 (N_36783,N_34869,N_30857);
nand U36784 (N_36784,N_30149,N_30887);
and U36785 (N_36785,N_32462,N_32643);
nand U36786 (N_36786,N_33888,N_30917);
nor U36787 (N_36787,N_32749,N_31055);
xnor U36788 (N_36788,N_34262,N_32326);
or U36789 (N_36789,N_33396,N_30321);
or U36790 (N_36790,N_31136,N_34488);
nand U36791 (N_36791,N_34692,N_31106);
or U36792 (N_36792,N_33487,N_31315);
xor U36793 (N_36793,N_30647,N_30525);
or U36794 (N_36794,N_34956,N_33364);
nand U36795 (N_36795,N_32807,N_33729);
or U36796 (N_36796,N_30306,N_32835);
or U36797 (N_36797,N_30854,N_31859);
xor U36798 (N_36798,N_32840,N_33580);
nand U36799 (N_36799,N_30147,N_33953);
or U36800 (N_36800,N_30081,N_30107);
nor U36801 (N_36801,N_33747,N_30278);
xor U36802 (N_36802,N_30361,N_31252);
nand U36803 (N_36803,N_31561,N_31598);
xor U36804 (N_36804,N_30436,N_31025);
and U36805 (N_36805,N_34796,N_34028);
nor U36806 (N_36806,N_31565,N_32829);
nor U36807 (N_36807,N_30946,N_32287);
or U36808 (N_36808,N_34642,N_34862);
or U36809 (N_36809,N_31807,N_30687);
nor U36810 (N_36810,N_33759,N_31230);
and U36811 (N_36811,N_34764,N_30129);
nand U36812 (N_36812,N_34126,N_31497);
and U36813 (N_36813,N_30144,N_34741);
xor U36814 (N_36814,N_31139,N_30313);
and U36815 (N_36815,N_32061,N_31912);
and U36816 (N_36816,N_32433,N_34638);
and U36817 (N_36817,N_32204,N_33898);
or U36818 (N_36818,N_33647,N_30627);
nor U36819 (N_36819,N_32029,N_34826);
nand U36820 (N_36820,N_30710,N_33720);
xnor U36821 (N_36821,N_33976,N_31862);
and U36822 (N_36822,N_32852,N_34233);
or U36823 (N_36823,N_30462,N_32621);
or U36824 (N_36824,N_31217,N_34310);
or U36825 (N_36825,N_31731,N_33381);
xnor U36826 (N_36826,N_33824,N_34302);
xnor U36827 (N_36827,N_32785,N_30074);
xnor U36828 (N_36828,N_33032,N_30740);
nand U36829 (N_36829,N_32149,N_31733);
nand U36830 (N_36830,N_34944,N_30008);
xor U36831 (N_36831,N_33207,N_32956);
xor U36832 (N_36832,N_32519,N_33036);
nand U36833 (N_36833,N_33932,N_32843);
nand U36834 (N_36834,N_31502,N_34284);
nand U36835 (N_36835,N_31501,N_34319);
nand U36836 (N_36836,N_31578,N_32814);
nor U36837 (N_36837,N_33397,N_34031);
and U36838 (N_36838,N_30715,N_32658);
xor U36839 (N_36839,N_32442,N_33068);
and U36840 (N_36840,N_33688,N_32675);
or U36841 (N_36841,N_34370,N_34793);
nor U36842 (N_36842,N_32260,N_30886);
and U36843 (N_36843,N_30179,N_31631);
and U36844 (N_36844,N_32753,N_32123);
or U36845 (N_36845,N_33208,N_32904);
and U36846 (N_36846,N_34949,N_30660);
or U36847 (N_36847,N_34510,N_32861);
or U36848 (N_36848,N_34703,N_32751);
nand U36849 (N_36849,N_34713,N_31134);
xor U36850 (N_36850,N_31574,N_34205);
or U36851 (N_36851,N_31157,N_34386);
and U36852 (N_36852,N_32713,N_33811);
nor U36853 (N_36853,N_33962,N_30549);
xnor U36854 (N_36854,N_33220,N_32139);
nor U36855 (N_36855,N_31800,N_30824);
nor U36856 (N_36856,N_31616,N_34868);
xor U36857 (N_36857,N_34918,N_31571);
nor U36858 (N_36858,N_32415,N_33762);
nand U36859 (N_36859,N_30719,N_33845);
or U36860 (N_36860,N_30836,N_32459);
nor U36861 (N_36861,N_31923,N_33352);
and U36862 (N_36862,N_33942,N_32841);
xor U36863 (N_36863,N_33829,N_31284);
and U36864 (N_36864,N_30684,N_33752);
and U36865 (N_36865,N_31465,N_34322);
nor U36866 (N_36866,N_31378,N_30235);
nand U36867 (N_36867,N_30197,N_34043);
or U36868 (N_36868,N_31682,N_31110);
xor U36869 (N_36869,N_31087,N_31360);
nor U36870 (N_36870,N_31537,N_33766);
nor U36871 (N_36871,N_33379,N_33901);
nand U36872 (N_36872,N_33378,N_33231);
nor U36873 (N_36873,N_33687,N_34567);
or U36874 (N_36874,N_33903,N_31070);
and U36875 (N_36875,N_31492,N_34199);
nor U36876 (N_36876,N_33921,N_31433);
nand U36877 (N_36877,N_31177,N_34524);
nand U36878 (N_36878,N_30645,N_30250);
xnor U36879 (N_36879,N_31407,N_32293);
xnor U36880 (N_36880,N_30738,N_31452);
xnor U36881 (N_36881,N_33944,N_33716);
xor U36882 (N_36882,N_31791,N_30216);
xor U36883 (N_36883,N_30636,N_33421);
xnor U36884 (N_36884,N_32699,N_32705);
and U36885 (N_36885,N_31935,N_33124);
or U36886 (N_36886,N_32032,N_31146);
and U36887 (N_36887,N_30227,N_30064);
xor U36888 (N_36888,N_30919,N_32407);
nand U36889 (N_36889,N_30438,N_32178);
nand U36890 (N_36890,N_31759,N_32256);
xor U36891 (N_36891,N_32733,N_34067);
nand U36892 (N_36892,N_32217,N_33538);
nor U36893 (N_36893,N_32767,N_30041);
nor U36894 (N_36894,N_33525,N_31726);
nor U36895 (N_36895,N_32592,N_34632);
or U36896 (N_36896,N_30190,N_30266);
nand U36897 (N_36897,N_33366,N_31984);
nor U36898 (N_36898,N_33809,N_32782);
nor U36899 (N_36899,N_34912,N_32351);
and U36900 (N_36900,N_34540,N_32111);
nand U36901 (N_36901,N_32392,N_32228);
xor U36902 (N_36902,N_32490,N_32683);
and U36903 (N_36903,N_34523,N_34368);
or U36904 (N_36904,N_32346,N_33879);
xor U36905 (N_36905,N_32050,N_33470);
xnor U36906 (N_36906,N_30582,N_31955);
and U36907 (N_36907,N_33950,N_34209);
nor U36908 (N_36908,N_33222,N_33164);
and U36909 (N_36909,N_34239,N_31648);
xnor U36910 (N_36910,N_31721,N_34786);
nand U36911 (N_36911,N_33429,N_34687);
and U36912 (N_36912,N_32887,N_30464);
nand U36913 (N_36913,N_34084,N_34249);
nand U36914 (N_36914,N_33383,N_31965);
nor U36915 (N_36915,N_31995,N_34429);
xor U36916 (N_36916,N_32585,N_30566);
or U36917 (N_36917,N_31458,N_33562);
xnor U36918 (N_36918,N_34606,N_34984);
xnor U36919 (N_36919,N_31626,N_32742);
nor U36920 (N_36920,N_30902,N_31243);
nand U36921 (N_36921,N_32013,N_31188);
nor U36922 (N_36922,N_33076,N_34035);
xor U36923 (N_36923,N_33589,N_32778);
nand U36924 (N_36924,N_33863,N_33488);
or U36925 (N_36925,N_34431,N_31077);
or U36926 (N_36926,N_34277,N_32493);
and U36927 (N_36927,N_31279,N_34654);
xor U36928 (N_36928,N_31225,N_33269);
nand U36929 (N_36929,N_30374,N_31084);
xor U36930 (N_36930,N_30080,N_33372);
nor U36931 (N_36931,N_30053,N_30672);
nor U36932 (N_36932,N_31692,N_34235);
nand U36933 (N_36933,N_32694,N_30005);
xnor U36934 (N_36934,N_30242,N_30155);
or U36935 (N_36935,N_30863,N_33532);
xor U36936 (N_36936,N_30006,N_34887);
nor U36937 (N_36937,N_32086,N_34725);
nand U36938 (N_36938,N_34905,N_31385);
and U36939 (N_36939,N_31882,N_33420);
xor U36940 (N_36940,N_30345,N_33412);
and U36941 (N_36941,N_33676,N_32193);
xnor U36942 (N_36942,N_30161,N_31293);
or U36943 (N_36943,N_33363,N_30906);
or U36944 (N_36944,N_30643,N_30813);
nand U36945 (N_36945,N_32166,N_30318);
or U36946 (N_36946,N_34785,N_31608);
xnor U36947 (N_36947,N_30355,N_32867);
xnor U36948 (N_36948,N_34479,N_31960);
nor U36949 (N_36949,N_30198,N_34585);
and U36950 (N_36950,N_30910,N_34141);
xor U36951 (N_36951,N_30247,N_33636);
nand U36952 (N_36952,N_32065,N_34201);
nor U36953 (N_36953,N_34839,N_32372);
nor U36954 (N_36954,N_30024,N_31460);
nor U36955 (N_36955,N_32034,N_31268);
nand U36956 (N_36956,N_30413,N_31267);
nor U36957 (N_36957,N_34503,N_31404);
nand U36958 (N_36958,N_32001,N_33119);
xnor U36959 (N_36959,N_34600,N_32952);
or U36960 (N_36960,N_34422,N_33251);
nor U36961 (N_36961,N_33370,N_31729);
or U36962 (N_36962,N_32215,N_32026);
and U36963 (N_36963,N_32615,N_30133);
nor U36964 (N_36964,N_32662,N_34610);
nand U36965 (N_36965,N_34326,N_30980);
nor U36966 (N_36966,N_31237,N_34500);
nand U36967 (N_36967,N_31247,N_34292);
or U36968 (N_36968,N_34593,N_31053);
or U36969 (N_36969,N_33986,N_34788);
and U36970 (N_36970,N_34344,N_34604);
nand U36971 (N_36971,N_33640,N_31803);
and U36972 (N_36972,N_33520,N_34824);
nand U36973 (N_36973,N_30967,N_34941);
nand U36974 (N_36974,N_33755,N_32202);
xor U36975 (N_36975,N_30829,N_33998);
and U36976 (N_36976,N_31549,N_30478);
or U36977 (N_36977,N_31012,N_32727);
and U36978 (N_36978,N_32542,N_31117);
or U36979 (N_36979,N_30765,N_34673);
nor U36980 (N_36980,N_31251,N_31464);
nand U36981 (N_36981,N_31817,N_34434);
nand U36982 (N_36982,N_34805,N_31621);
nor U36983 (N_36983,N_32976,N_30976);
xnor U36984 (N_36984,N_31091,N_33877);
xnor U36985 (N_36985,N_30642,N_34804);
xor U36986 (N_36986,N_32373,N_31543);
xnor U36987 (N_36987,N_32427,N_30240);
nand U36988 (N_36988,N_30760,N_34355);
and U36989 (N_36989,N_33117,N_33553);
xnor U36990 (N_36990,N_30882,N_34433);
nor U36991 (N_36991,N_30818,N_32176);
or U36992 (N_36992,N_33319,N_31630);
xnor U36993 (N_36993,N_32800,N_30142);
or U36994 (N_36994,N_32856,N_31758);
or U36995 (N_36995,N_30157,N_34129);
xor U36996 (N_36996,N_31853,N_33871);
nand U36997 (N_36997,N_34977,N_31645);
xnor U36998 (N_36998,N_33138,N_31469);
nand U36999 (N_36999,N_34072,N_30587);
nor U37000 (N_37000,N_31206,N_34937);
and U37001 (N_37001,N_34620,N_31309);
or U37002 (N_37002,N_32722,N_30679);
nand U37003 (N_37003,N_34169,N_33434);
nand U37004 (N_37004,N_34584,N_31422);
nor U37005 (N_37005,N_32031,N_32009);
or U37006 (N_37006,N_34534,N_31877);
nor U37007 (N_37007,N_30359,N_31886);
nor U37008 (N_37008,N_32690,N_30284);
and U37009 (N_37009,N_31839,N_33365);
nor U37010 (N_37010,N_34452,N_31994);
or U37011 (N_37011,N_33567,N_32154);
nand U37012 (N_37012,N_33102,N_32162);
and U37013 (N_37013,N_34211,N_34202);
nor U37014 (N_37014,N_33548,N_34248);
nand U37015 (N_37015,N_33708,N_30618);
or U37016 (N_37016,N_34701,N_34769);
xnor U37017 (N_37017,N_31199,N_33198);
or U37018 (N_37018,N_32967,N_32040);
or U37019 (N_37019,N_33427,N_33897);
and U37020 (N_37020,N_34923,N_30699);
nand U37021 (N_37021,N_32475,N_34423);
and U37022 (N_37022,N_33214,N_33390);
nor U37023 (N_37023,N_32486,N_32468);
nor U37024 (N_37024,N_31540,N_33935);
nor U37025 (N_37025,N_31739,N_33325);
and U37026 (N_37026,N_32973,N_32241);
or U37027 (N_37027,N_30669,N_30061);
nor U37028 (N_37028,N_33460,N_31389);
or U37029 (N_37029,N_32426,N_33357);
or U37030 (N_37030,N_30409,N_33163);
or U37031 (N_37031,N_30786,N_32884);
xor U37032 (N_37032,N_33797,N_31988);
nand U37033 (N_37033,N_33857,N_30858);
or U37034 (N_37034,N_31356,N_34146);
xor U37035 (N_37035,N_34032,N_30494);
and U37036 (N_37036,N_34004,N_31266);
or U37037 (N_37037,N_32608,N_30411);
nor U37038 (N_37038,N_31532,N_30089);
nor U37039 (N_37039,N_31819,N_34381);
and U37040 (N_37040,N_34472,N_32746);
and U37041 (N_37041,N_34056,N_34957);
and U37042 (N_37042,N_32058,N_31622);
and U37043 (N_37043,N_33055,N_31145);
or U37044 (N_37044,N_32315,N_32707);
or U37045 (N_37045,N_34979,N_34601);
and U37046 (N_37046,N_31311,N_33516);
and U37047 (N_37047,N_31747,N_34751);
xor U37048 (N_37048,N_33557,N_32684);
and U37049 (N_37049,N_32066,N_31619);
nor U37050 (N_37050,N_31806,N_31674);
and U37051 (N_37051,N_34988,N_34224);
and U37052 (N_37052,N_32363,N_34597);
and U37053 (N_37053,N_31930,N_30407);
and U37054 (N_37054,N_31929,N_34348);
nand U37055 (N_37055,N_31185,N_34617);
and U37056 (N_37056,N_33613,N_31798);
nand U37057 (N_37057,N_34986,N_33728);
or U37058 (N_37058,N_31100,N_31476);
xor U37059 (N_37059,N_34012,N_32842);
nor U37060 (N_37060,N_34416,N_32655);
nor U37061 (N_37061,N_31299,N_33279);
and U37062 (N_37062,N_32308,N_33808);
xor U37063 (N_37063,N_32008,N_33075);
nor U37064 (N_37064,N_32711,N_30810);
and U37065 (N_37065,N_34655,N_32151);
nor U37066 (N_37066,N_31449,N_30825);
and U37067 (N_37067,N_30246,N_31998);
nand U37068 (N_37068,N_30988,N_34772);
nand U37069 (N_37069,N_33496,N_33778);
xnor U37070 (N_37070,N_34747,N_30452);
and U37071 (N_37071,N_33896,N_32474);
nand U37072 (N_37072,N_32186,N_30931);
xnor U37073 (N_37073,N_30295,N_34970);
nand U37074 (N_37074,N_34405,N_30531);
xor U37075 (N_37075,N_34717,N_32370);
nor U37076 (N_37076,N_31618,N_34295);
nor U37077 (N_37077,N_30482,N_30621);
or U37078 (N_37078,N_32514,N_31259);
nor U37079 (N_37079,N_32272,N_30616);
xor U37080 (N_37080,N_32406,N_32347);
nor U37081 (N_37081,N_33107,N_31939);
xnor U37082 (N_37082,N_31586,N_33440);
xnor U37083 (N_37083,N_32400,N_31485);
nor U37084 (N_37084,N_32394,N_32087);
nor U37085 (N_37085,N_33860,N_31017);
nand U37086 (N_37086,N_32743,N_30199);
and U37087 (N_37087,N_33603,N_32871);
or U37088 (N_37088,N_31652,N_33409);
nor U37089 (N_37089,N_30140,N_32128);
nand U37090 (N_37090,N_33573,N_31594);
xor U37091 (N_37091,N_31447,N_33108);
nor U37092 (N_37092,N_33802,N_31096);
and U37093 (N_37093,N_33384,N_31884);
or U37094 (N_37094,N_30372,N_33294);
nor U37095 (N_37095,N_33221,N_31771);
nor U37096 (N_37096,N_32737,N_32455);
xnor U37097 (N_37097,N_30893,N_30207);
xor U37098 (N_37098,N_33147,N_32790);
and U37099 (N_37099,N_31294,N_32358);
nor U37100 (N_37100,N_33504,N_32959);
nand U37101 (N_37101,N_33335,N_32984);
or U37102 (N_37102,N_34831,N_33884);
nor U37103 (N_37103,N_32828,N_34426);
nand U37104 (N_37104,N_31748,N_34137);
or U37105 (N_37105,N_34783,N_32888);
xor U37106 (N_37106,N_34267,N_32651);
xor U37107 (N_37107,N_30273,N_30617);
nor U37108 (N_37108,N_33046,N_32200);
and U37109 (N_37109,N_34131,N_30426);
xor U37110 (N_37110,N_30930,N_34939);
or U37111 (N_37111,N_34874,N_33570);
nand U37112 (N_37112,N_32576,N_33703);
xnor U37113 (N_37113,N_33836,N_31255);
xnor U37114 (N_37114,N_30800,N_30918);
nand U37115 (N_37115,N_30439,N_32444);
nor U37116 (N_37116,N_30744,N_31701);
and U37117 (N_37117,N_34069,N_30891);
or U37118 (N_37118,N_30580,N_32560);
xnor U37119 (N_37119,N_33280,N_33602);
xor U37120 (N_37120,N_32329,N_32461);
xor U37121 (N_37121,N_30279,N_31691);
nand U37122 (N_37122,N_32027,N_34401);
or U37123 (N_37123,N_33224,N_30018);
nor U37124 (N_37124,N_34441,N_32761);
nand U37125 (N_37125,N_33939,N_33724);
xnor U37126 (N_37126,N_34365,N_32466);
nor U37127 (N_37127,N_32798,N_32463);
nand U37128 (N_37128,N_30640,N_30912);
nor U37129 (N_37129,N_32726,N_32084);
and U37130 (N_37130,N_32126,N_31607);
xnor U37131 (N_37131,N_32773,N_32591);
xnor U37132 (N_37132,N_32604,N_33015);
nor U37133 (N_37133,N_30264,N_34566);
and U37134 (N_37134,N_34120,N_31904);
or U37135 (N_37135,N_31697,N_32569);
nand U37136 (N_37136,N_32666,N_32739);
nor U37137 (N_37137,N_31849,N_32913);
nor U37138 (N_37138,N_34070,N_31455);
and U37139 (N_37139,N_31661,N_34893);
and U37140 (N_37140,N_33695,N_30384);
nand U37141 (N_37141,N_34745,N_30244);
nor U37142 (N_37142,N_34339,N_32775);
or U37143 (N_37143,N_31287,N_33215);
nand U37144 (N_37144,N_31810,N_33298);
and U37145 (N_37145,N_31641,N_34698);
xor U37146 (N_37146,N_30879,N_34666);
or U37147 (N_37147,N_32453,N_33813);
xor U37148 (N_37148,N_32511,N_30794);
or U37149 (N_37149,N_30483,N_32414);
or U37150 (N_37150,N_33096,N_30758);
or U37151 (N_37151,N_34101,N_33820);
and U37152 (N_37152,N_34089,N_33177);
or U37153 (N_37153,N_31200,N_30166);
xor U37154 (N_37154,N_34053,N_32985);
nor U37155 (N_37155,N_33605,N_30673);
and U37156 (N_37156,N_30397,N_32697);
xnor U37157 (N_37157,N_31192,N_33882);
nand U37158 (N_37158,N_34156,N_30631);
nor U37159 (N_37159,N_31067,N_32053);
xnor U37160 (N_37160,N_30267,N_31959);
xnor U37161 (N_37161,N_33632,N_32549);
and U37162 (N_37162,N_34697,N_30927);
or U37163 (N_37163,N_31004,N_32740);
nor U37164 (N_37164,N_30513,N_33841);
nor U37165 (N_37165,N_31445,N_34417);
nand U37166 (N_37166,N_34312,N_34744);
xnor U37167 (N_37167,N_31194,N_33983);
nand U37168 (N_37168,N_34706,N_34696);
and U37169 (N_37169,N_33517,N_34435);
nand U37170 (N_37170,N_33453,N_34830);
nor U37171 (N_37171,N_34086,N_32440);
nor U37172 (N_37172,N_34170,N_33479);
or U37173 (N_37173,N_32338,N_34377);
nor U37174 (N_37174,N_32981,N_34809);
xnor U37175 (N_37175,N_34393,N_32550);
or U37176 (N_37176,N_30395,N_34827);
and U37177 (N_37177,N_34241,N_32936);
and U37178 (N_37178,N_33908,N_33547);
or U37179 (N_37179,N_33641,N_34127);
nor U37180 (N_37180,N_31926,N_34602);
or U37181 (N_37181,N_30579,N_32671);
xor U37182 (N_37182,N_31285,N_31448);
and U37183 (N_37183,N_31666,N_30031);
nand U37184 (N_37184,N_30253,N_31163);
nand U37185 (N_37185,N_32434,N_32080);
nor U37186 (N_37186,N_34364,N_31074);
or U37187 (N_37187,N_32744,N_31141);
xor U37188 (N_37188,N_32636,N_31917);
nand U37189 (N_37189,N_34753,N_34609);
nand U37190 (N_37190,N_31508,N_30432);
nand U37191 (N_37191,N_31489,N_32284);
and U37192 (N_37192,N_33777,N_31944);
or U37193 (N_37193,N_32715,N_33990);
nor U37194 (N_37194,N_30869,N_32940);
nor U37195 (N_37195,N_31943,N_31429);
nor U37196 (N_37196,N_31295,N_33232);
or U37197 (N_37197,N_32371,N_31664);
and U37198 (N_37198,N_31467,N_34758);
and U37199 (N_37199,N_33957,N_32567);
and U37200 (N_37200,N_33121,N_31716);
xor U37201 (N_37201,N_34139,N_34910);
nand U37202 (N_37202,N_32941,N_32327);
xor U37203 (N_37203,N_31415,N_32586);
xnor U37204 (N_37204,N_30431,N_30848);
or U37205 (N_37205,N_33823,N_34299);
xnor U37206 (N_37206,N_34959,N_33200);
nand U37207 (N_37207,N_34020,N_34294);
or U37208 (N_37208,N_33038,N_32179);
nor U37209 (N_37209,N_33717,N_30762);
and U37210 (N_37210,N_33149,N_32299);
nand U37211 (N_37211,N_33243,N_34808);
and U37212 (N_37212,N_30808,N_31934);
xnor U37213 (N_37213,N_30633,N_32714);
or U37214 (N_37214,N_31066,N_33714);
or U37215 (N_37215,N_33310,N_32491);
nor U37216 (N_37216,N_31408,N_32993);
nand U37217 (N_37217,N_34341,N_31414);
xnor U37218 (N_37218,N_31297,N_33444);
nand U37219 (N_37219,N_33734,N_31198);
nand U37220 (N_37220,N_32278,N_32004);
or U37221 (N_37221,N_34218,N_33115);
xor U37222 (N_37222,N_33495,N_32605);
and U37223 (N_37223,N_33330,N_31776);
nand U37224 (N_37224,N_32352,N_34390);
xnor U37225 (N_37225,N_31848,N_34555);
or U37226 (N_37226,N_30753,N_30940);
nor U37227 (N_37227,N_30790,N_31677);
nand U37228 (N_37228,N_34775,N_30146);
or U37229 (N_37229,N_33798,N_34603);
nor U37230 (N_37230,N_34088,N_33437);
nor U37231 (N_37231,N_33835,N_31161);
nand U37232 (N_37232,N_34173,N_30175);
xnor U37233 (N_37233,N_31528,N_32750);
and U37234 (N_37234,N_34324,N_31138);
nor U37235 (N_37235,N_34407,N_32429);
nor U37236 (N_37236,N_33634,N_31085);
nor U37237 (N_37237,N_32927,N_34851);
xor U37238 (N_37238,N_31118,N_32650);
and U37239 (N_37239,N_30601,N_31114);
and U37240 (N_37240,N_31617,N_32877);
nand U37241 (N_37241,N_30290,N_32045);
nor U37242 (N_37242,N_31986,N_33698);
and U37243 (N_37243,N_32473,N_31596);
nor U37244 (N_37244,N_30364,N_32745);
nor U37245 (N_37245,N_31636,N_30732);
xor U37246 (N_37246,N_31821,N_34712);
nor U37247 (N_37247,N_33180,N_30683);
and U37248 (N_37248,N_31124,N_33583);
nand U37249 (N_37249,N_34634,N_31062);
nand U37250 (N_37250,N_33972,N_33730);
nor U37251 (N_37251,N_30688,N_30540);
or U37252 (N_37252,N_34505,N_32863);
and U37253 (N_37253,N_33417,N_31137);
nor U37254 (N_37254,N_32477,N_32136);
or U37255 (N_37255,N_31577,N_31007);
or U37256 (N_37256,N_32263,N_32850);
nand U37257 (N_37257,N_33290,N_33229);
nand U37258 (N_37258,N_33918,N_31183);
nand U37259 (N_37259,N_30734,N_31173);
nand U37260 (N_37260,N_32507,N_32975);
or U37261 (N_37261,N_33864,N_30268);
or U37262 (N_37262,N_34118,N_34508);
xnor U37263 (N_37263,N_30785,N_32353);
or U37264 (N_37264,N_31398,N_34946);
and U37265 (N_37265,N_33508,N_34414);
nand U37266 (N_37266,N_34080,N_32057);
and U37267 (N_37267,N_32555,N_34968);
nor U37268 (N_37268,N_34599,N_33404);
xor U37269 (N_37269,N_32972,N_34660);
xnor U37270 (N_37270,N_30067,N_32574);
xnor U37271 (N_37271,N_33303,N_34735);
nand U37272 (N_37272,N_31952,N_31088);
or U37273 (N_37273,N_32610,N_31048);
or U37274 (N_37274,N_31369,N_30277);
nor U37275 (N_37275,N_33706,N_32199);
xor U37276 (N_37276,N_30111,N_32060);
nand U37277 (N_37277,N_32837,N_31918);
nand U37278 (N_37278,N_31572,N_30909);
or U37279 (N_37279,N_31495,N_33291);
xnor U37280 (N_37280,N_33527,N_31779);
or U37281 (N_37281,N_34231,N_33018);
or U37282 (N_37282,N_30260,N_34554);
and U37283 (N_37283,N_34208,N_32425);
nor U37284 (N_37284,N_30178,N_32813);
xor U37285 (N_37285,N_31470,N_32396);
nand U37286 (N_37286,N_31425,N_31320);
nand U37287 (N_37287,N_32864,N_30871);
nor U37288 (N_37288,N_30020,N_30421);
and U37289 (N_37289,N_32649,N_31590);
nor U37290 (N_37290,N_32577,N_31804);
and U37291 (N_37291,N_32875,N_32885);
nand U37292 (N_37292,N_30538,N_31301);
nor U37293 (N_37293,N_34375,N_34244);
xnor U37294 (N_37294,N_33336,N_31112);
and U37295 (N_37295,N_31280,N_32784);
xnor U37296 (N_37296,N_34087,N_31122);
nor U37297 (N_37297,N_30265,N_34077);
nand U37298 (N_37298,N_32977,N_33889);
xor U37299 (N_37299,N_33425,N_32600);
xor U37300 (N_37300,N_33765,N_34746);
and U37301 (N_37301,N_31228,N_30860);
nor U37302 (N_37302,N_32335,N_30812);
nand U37303 (N_37303,N_34828,N_33595);
and U37304 (N_37304,N_34456,N_33913);
and U37305 (N_37305,N_31132,N_33254);
nor U37306 (N_37306,N_33493,N_33266);
nor U37307 (N_37307,N_33086,N_32183);
nor U37308 (N_37308,N_34668,N_31724);
xor U37309 (N_37309,N_33920,N_31525);
and U37310 (N_37310,N_30649,N_32634);
nor U37311 (N_37311,N_32167,N_33006);
nor U37312 (N_37312,N_31105,N_33178);
or U37313 (N_37313,N_33244,N_34895);
nand U37314 (N_37314,N_31265,N_30851);
xnor U37315 (N_37315,N_32896,N_31366);
nand U37316 (N_37316,N_32880,N_30324);
nor U37317 (N_37317,N_34571,N_32898);
or U37318 (N_37318,N_33464,N_31496);
or U37319 (N_37319,N_32640,N_32613);
nand U37320 (N_37320,N_32483,N_34667);
and U37321 (N_37321,N_30962,N_32832);
and U37322 (N_37322,N_31797,N_33856);
or U37323 (N_37323,N_32595,N_34014);
xnor U37324 (N_37324,N_34539,N_30036);
and U37325 (N_37325,N_33989,N_30023);
nand U37326 (N_37326,N_34409,N_33154);
or U37327 (N_37327,N_32101,N_32866);
or U37328 (N_37328,N_34177,N_34533);
nand U37329 (N_37329,N_31658,N_30514);
xor U37330 (N_37330,N_31440,N_30449);
nand U37331 (N_37331,N_30326,N_30486);
xnor U37332 (N_37332,N_30705,N_32988);
or U37333 (N_37333,N_30703,N_30475);
or U37334 (N_37334,N_34351,N_30121);
and U37335 (N_37335,N_31690,N_33971);
and U37336 (N_37336,N_32385,N_33529);
xnor U37337 (N_37337,N_32559,N_34064);
and U37338 (N_37338,N_30225,N_34637);
nor U37339 (N_37339,N_33793,N_30907);
and U37340 (N_37340,N_31909,N_30780);
or U37341 (N_37341,N_33258,N_31033);
nor U37342 (N_37342,N_34945,N_30150);
xor U37343 (N_37343,N_32285,N_32096);
and U37344 (N_37344,N_34440,N_34037);
nand U37345 (N_37345,N_33392,N_33810);
xnor U37346 (N_37346,N_30781,N_30583);
and U37347 (N_37347,N_31564,N_32180);
xor U37348 (N_37348,N_34529,N_31089);
and U37349 (N_37349,N_32954,N_34030);
and U37350 (N_37350,N_30088,N_34927);
nand U37351 (N_37351,N_32673,N_30315);
xnor U37352 (N_37352,N_31115,N_34779);
or U37353 (N_37353,N_34015,N_33026);
or U37354 (N_37354,N_32534,N_31902);
nor U37355 (N_37355,N_34258,N_34091);
and U37356 (N_37356,N_32922,N_31043);
or U37357 (N_37357,N_32934,N_30145);
nand U37358 (N_37358,N_30904,N_31056);
nor U37359 (N_37359,N_30928,N_31749);
nand U37360 (N_37360,N_32104,N_34143);
nand U37361 (N_37361,N_30652,N_32382);
nor U37362 (N_37362,N_34396,N_32405);
nand U37363 (N_37363,N_33401,N_34616);
and U37364 (N_37364,N_30721,N_30070);
or U37365 (N_37365,N_32435,N_30737);
nand U37366 (N_37366,N_33347,N_32482);
nand U37367 (N_37367,N_30122,N_34542);
and U37368 (N_37368,N_31907,N_32402);
xnor U37369 (N_37369,N_34192,N_32257);
nor U37370 (N_37370,N_32097,N_30837);
nor U37371 (N_37371,N_34222,N_30611);
nor U37372 (N_37372,N_31547,N_34820);
nor U37373 (N_37373,N_31602,N_33239);
nand U37374 (N_37374,N_31095,N_31521);
xnor U37375 (N_37375,N_33973,N_32280);
or U37376 (N_37376,N_32157,N_33592);
or U37377 (N_37377,N_30403,N_33978);
nor U37378 (N_37378,N_31334,N_30709);
and U37379 (N_37379,N_34125,N_31969);
or U37380 (N_37380,N_31172,N_32757);
or U37381 (N_37381,N_32017,N_32622);
or U37382 (N_37382,N_31245,N_31945);
and U37383 (N_37383,N_34268,N_33965);
nor U37384 (N_37384,N_34914,N_34360);
nand U37385 (N_37385,N_33212,N_34449);
or U37386 (N_37386,N_34469,N_34715);
and U37387 (N_37387,N_31670,N_30084);
xnor U37388 (N_37388,N_32489,N_34017);
and U37389 (N_37389,N_34528,N_33799);
nand U37390 (N_37390,N_32446,N_30535);
nor U37391 (N_37391,N_31459,N_33426);
nor U37392 (N_37392,N_31992,N_32704);
nand U37393 (N_37393,N_34999,N_32712);
or U37394 (N_37394,N_30571,N_34371);
nand U37395 (N_37395,N_34690,N_34565);
or U37396 (N_37396,N_34513,N_33643);
or U37397 (N_37397,N_30834,N_33585);
xor U37398 (N_37398,N_34878,N_32221);
nand U37399 (N_37399,N_32078,N_32042);
and U37400 (N_37400,N_31766,N_31827);
or U37401 (N_37401,N_32968,N_30713);
or U37402 (N_37402,N_32964,N_34260);
xor U37403 (N_37403,N_31820,N_30875);
or U37404 (N_37404,N_31837,N_32823);
xnor U37405 (N_37405,N_30770,N_32838);
xnor U37406 (N_37406,N_34085,N_31973);
and U37407 (N_37407,N_31624,N_32099);
and U37408 (N_37408,N_32854,N_34220);
or U37409 (N_37409,N_33615,N_32010);
or U37410 (N_37410,N_33176,N_30963);
and U37411 (N_37411,N_31864,N_33000);
or U37412 (N_37412,N_34817,N_34569);
or U37413 (N_37413,N_32645,N_33788);
or U37414 (N_37414,N_34641,N_32531);
nand U37415 (N_37415,N_34016,N_31635);
or U37416 (N_37416,N_30743,N_33307);
and U37417 (N_37417,N_32932,N_33967);
and U37418 (N_37418,N_32618,N_31964);
nand U37419 (N_37419,N_34619,N_31569);
nand U37420 (N_37420,N_30815,N_34180);
or U37421 (N_37421,N_32120,N_33596);
nor U37422 (N_37422,N_31109,N_34047);
nand U37423 (N_37423,N_32437,N_31075);
nand U37424 (N_37424,N_31783,N_31812);
xnor U37425 (N_37425,N_30569,N_34155);
and U37426 (N_37426,N_34739,N_33574);
and U37427 (N_37427,N_31894,N_33738);
xor U37428 (N_37428,N_33233,N_31174);
nor U37429 (N_37429,N_33800,N_31861);
xor U37430 (N_37430,N_30275,N_31625);
and U37431 (N_37431,N_33010,N_30249);
or U37432 (N_37432,N_31358,N_34614);
or U37433 (N_37433,N_34580,N_30045);
and U37434 (N_37434,N_31855,N_32328);
xnor U37435 (N_37435,N_31151,N_34516);
xnor U37436 (N_37436,N_33382,N_31477);
xor U37437 (N_37437,N_34194,N_31319);
or U37438 (N_37438,N_30796,N_32948);
nor U37439 (N_37439,N_32349,N_33235);
nand U37440 (N_37440,N_33646,N_33084);
and U37441 (N_37441,N_31940,N_31516);
nand U37442 (N_37442,N_31044,N_31030);
nand U37443 (N_37443,N_30338,N_31813);
xnor U37444 (N_37444,N_32485,N_32100);
and U37445 (N_37445,N_34013,N_32503);
and U37446 (N_37446,N_30998,N_30058);
and U37447 (N_37447,N_32558,N_32148);
nand U37448 (N_37448,N_30172,N_34027);
nand U37449 (N_37449,N_31714,N_30118);
xnor U37450 (N_37450,N_33457,N_34316);
and U37451 (N_37451,N_31931,N_33938);
nand U37452 (N_37452,N_33481,N_30802);
xnor U37453 (N_37453,N_30055,N_31999);
xnor U37454 (N_37454,N_31387,N_31318);
nor U37455 (N_37455,N_33074,N_32242);
nand U37456 (N_37456,N_32230,N_31836);
nor U37457 (N_37457,N_30090,N_30676);
or U37458 (N_37458,N_30047,N_33551);
xor U37459 (N_37459,N_30025,N_30529);
or U37460 (N_37460,N_34123,N_31675);
or U37461 (N_37461,N_31568,N_33722);
xnor U37462 (N_37462,N_32222,N_34176);
or U37463 (N_37463,N_32310,N_34478);
xor U37464 (N_37464,N_30391,N_32054);
nand U37465 (N_37465,N_34193,N_34844);
xnor U37466 (N_37466,N_33004,N_30987);
or U37467 (N_37467,N_30562,N_31498);
nor U37468 (N_37468,N_33911,N_34489);
xnor U37469 (N_37469,N_34518,N_33230);
nand U37470 (N_37470,N_34454,N_32641);
nand U37471 (N_37471,N_33063,N_33339);
xor U37472 (N_37472,N_33886,N_30951);
nand U37473 (N_37473,N_31409,N_34132);
and U37474 (N_37474,N_30992,N_34995);
or U37475 (N_37475,N_33644,N_31375);
and U37476 (N_37476,N_33132,N_30038);
or U37477 (N_37477,N_32720,N_33598);
nand U37478 (N_37478,N_32197,N_32860);
and U37479 (N_37479,N_30648,N_33476);
nand U37480 (N_37480,N_34272,N_34967);
nor U37481 (N_37481,N_32957,N_32906);
or U37482 (N_37482,N_30186,N_31856);
and U37483 (N_37483,N_30000,N_32472);
nand U37484 (N_37484,N_31102,N_30939);
or U37485 (N_37485,N_30959,N_34227);
or U37486 (N_37486,N_32071,N_33805);
or U37487 (N_37487,N_31054,N_30532);
xor U37488 (N_37488,N_31868,N_30548);
or U37489 (N_37489,N_34688,N_30251);
and U37490 (N_37490,N_31202,N_30003);
xor U37491 (N_37491,N_30908,N_30352);
nor U37492 (N_37492,N_31743,N_33746);
and U37493 (N_37493,N_32677,N_30076);
nor U37494 (N_37494,N_31417,N_32603);
nor U37495 (N_37495,N_30613,N_32047);
xnor U37496 (N_37496,N_33847,N_30799);
or U37497 (N_37497,N_32855,N_34217);
or U37498 (N_37498,N_30433,N_30926);
and U37499 (N_37499,N_32834,N_31493);
xor U37500 (N_37500,N_30236,N_32968);
nand U37501 (N_37501,N_32943,N_34864);
nand U37502 (N_37502,N_32067,N_34263);
or U37503 (N_37503,N_32624,N_30388);
or U37504 (N_37504,N_34851,N_31955);
or U37505 (N_37505,N_32347,N_34647);
or U37506 (N_37506,N_33103,N_30088);
nor U37507 (N_37507,N_31212,N_32265);
xor U37508 (N_37508,N_34413,N_33738);
and U37509 (N_37509,N_31100,N_30283);
xnor U37510 (N_37510,N_30872,N_32293);
nor U37511 (N_37511,N_33497,N_34986);
xnor U37512 (N_37512,N_31459,N_30085);
and U37513 (N_37513,N_31166,N_30977);
and U37514 (N_37514,N_31085,N_34404);
nor U37515 (N_37515,N_33186,N_33263);
xnor U37516 (N_37516,N_31762,N_33032);
or U37517 (N_37517,N_31068,N_34043);
and U37518 (N_37518,N_34838,N_31706);
and U37519 (N_37519,N_32683,N_31750);
xor U37520 (N_37520,N_34879,N_32985);
and U37521 (N_37521,N_34617,N_34373);
xnor U37522 (N_37522,N_33249,N_33419);
xor U37523 (N_37523,N_31422,N_32949);
and U37524 (N_37524,N_33248,N_30404);
nor U37525 (N_37525,N_32395,N_31932);
and U37526 (N_37526,N_31058,N_33430);
and U37527 (N_37527,N_32384,N_30779);
nand U37528 (N_37528,N_32908,N_33768);
nand U37529 (N_37529,N_32957,N_34085);
xnor U37530 (N_37530,N_32558,N_33967);
nor U37531 (N_37531,N_31522,N_34988);
xor U37532 (N_37532,N_32508,N_33335);
and U37533 (N_37533,N_34460,N_33898);
or U37534 (N_37534,N_31156,N_34559);
xor U37535 (N_37535,N_32710,N_31107);
nor U37536 (N_37536,N_33260,N_33429);
or U37537 (N_37537,N_32905,N_30580);
or U37538 (N_37538,N_30367,N_33604);
and U37539 (N_37539,N_32758,N_32216);
and U37540 (N_37540,N_33533,N_31272);
xnor U37541 (N_37541,N_34685,N_33540);
nor U37542 (N_37542,N_32327,N_33345);
nand U37543 (N_37543,N_31878,N_34503);
or U37544 (N_37544,N_33953,N_31098);
xnor U37545 (N_37545,N_32486,N_32202);
or U37546 (N_37546,N_34721,N_32213);
xnor U37547 (N_37547,N_34512,N_30494);
and U37548 (N_37548,N_33086,N_33001);
and U37549 (N_37549,N_33264,N_31361);
xnor U37550 (N_37550,N_34985,N_30396);
and U37551 (N_37551,N_30490,N_30337);
or U37552 (N_37552,N_32089,N_34350);
and U37553 (N_37553,N_34534,N_33347);
or U37554 (N_37554,N_34267,N_33413);
and U37555 (N_37555,N_31814,N_31636);
and U37556 (N_37556,N_34947,N_32148);
nand U37557 (N_37557,N_32954,N_30176);
and U37558 (N_37558,N_31288,N_34555);
nor U37559 (N_37559,N_34772,N_32671);
nand U37560 (N_37560,N_32560,N_34916);
or U37561 (N_37561,N_32872,N_30249);
and U37562 (N_37562,N_33062,N_33207);
nor U37563 (N_37563,N_33587,N_34950);
and U37564 (N_37564,N_30367,N_32603);
and U37565 (N_37565,N_30979,N_31739);
nor U37566 (N_37566,N_31922,N_34510);
or U37567 (N_37567,N_32440,N_34281);
xor U37568 (N_37568,N_33189,N_31098);
nand U37569 (N_37569,N_33435,N_34468);
or U37570 (N_37570,N_30915,N_33382);
xnor U37571 (N_37571,N_34356,N_32694);
and U37572 (N_37572,N_34219,N_34732);
nand U37573 (N_37573,N_31409,N_33498);
xor U37574 (N_37574,N_32885,N_34290);
and U37575 (N_37575,N_34471,N_32991);
nor U37576 (N_37576,N_31764,N_31327);
nor U37577 (N_37577,N_32298,N_30003);
or U37578 (N_37578,N_34084,N_32102);
and U37579 (N_37579,N_34756,N_34269);
nor U37580 (N_37580,N_34929,N_32201);
xor U37581 (N_37581,N_34812,N_30115);
or U37582 (N_37582,N_33845,N_32824);
nand U37583 (N_37583,N_31968,N_31264);
xor U37584 (N_37584,N_34538,N_30029);
and U37585 (N_37585,N_31956,N_34303);
and U37586 (N_37586,N_32689,N_31434);
or U37587 (N_37587,N_34304,N_34940);
and U37588 (N_37588,N_31470,N_33481);
and U37589 (N_37589,N_30720,N_34788);
nand U37590 (N_37590,N_31754,N_34075);
or U37591 (N_37591,N_31811,N_33515);
or U37592 (N_37592,N_33256,N_33103);
xnor U37593 (N_37593,N_32485,N_34252);
or U37594 (N_37594,N_33120,N_32237);
or U37595 (N_37595,N_32237,N_31075);
xor U37596 (N_37596,N_33625,N_32383);
xnor U37597 (N_37597,N_30207,N_30067);
and U37598 (N_37598,N_32456,N_33449);
or U37599 (N_37599,N_32959,N_34854);
and U37600 (N_37600,N_32233,N_34927);
and U37601 (N_37601,N_30773,N_34125);
xor U37602 (N_37602,N_30005,N_32182);
and U37603 (N_37603,N_32256,N_33072);
nor U37604 (N_37604,N_34021,N_34459);
nor U37605 (N_37605,N_34230,N_32016);
or U37606 (N_37606,N_32843,N_30618);
xor U37607 (N_37607,N_31035,N_34757);
or U37608 (N_37608,N_31800,N_31965);
nor U37609 (N_37609,N_30217,N_34186);
nor U37610 (N_37610,N_34724,N_30119);
nand U37611 (N_37611,N_31594,N_31515);
nor U37612 (N_37612,N_33456,N_33763);
nand U37613 (N_37613,N_33577,N_34259);
and U37614 (N_37614,N_32856,N_34531);
nor U37615 (N_37615,N_34908,N_30464);
nand U37616 (N_37616,N_33014,N_33716);
nor U37617 (N_37617,N_31572,N_32031);
xor U37618 (N_37618,N_31963,N_32947);
and U37619 (N_37619,N_30121,N_30073);
nor U37620 (N_37620,N_32693,N_32607);
xnor U37621 (N_37621,N_33875,N_34951);
xnor U37622 (N_37622,N_33820,N_34344);
nor U37623 (N_37623,N_33583,N_32508);
and U37624 (N_37624,N_30553,N_33483);
nor U37625 (N_37625,N_33276,N_30633);
and U37626 (N_37626,N_30340,N_31075);
and U37627 (N_37627,N_32683,N_33326);
nor U37628 (N_37628,N_31899,N_34093);
nand U37629 (N_37629,N_34410,N_33889);
and U37630 (N_37630,N_33778,N_31231);
nand U37631 (N_37631,N_30074,N_33252);
and U37632 (N_37632,N_32831,N_34136);
nand U37633 (N_37633,N_33216,N_33635);
or U37634 (N_37634,N_30243,N_34388);
or U37635 (N_37635,N_32024,N_30558);
nor U37636 (N_37636,N_33665,N_30656);
nor U37637 (N_37637,N_33202,N_33091);
and U37638 (N_37638,N_33124,N_34958);
xnor U37639 (N_37639,N_30003,N_31894);
nor U37640 (N_37640,N_34943,N_34597);
xor U37641 (N_37641,N_30303,N_31935);
xor U37642 (N_37642,N_30512,N_30715);
and U37643 (N_37643,N_33847,N_30722);
or U37644 (N_37644,N_30113,N_31790);
xnor U37645 (N_37645,N_30243,N_34501);
nand U37646 (N_37646,N_34504,N_33460);
nor U37647 (N_37647,N_33265,N_33233);
nand U37648 (N_37648,N_30492,N_30418);
xor U37649 (N_37649,N_34155,N_32170);
nor U37650 (N_37650,N_33353,N_32760);
and U37651 (N_37651,N_33047,N_32425);
or U37652 (N_37652,N_32197,N_30059);
xnor U37653 (N_37653,N_34052,N_34534);
or U37654 (N_37654,N_30635,N_30864);
nand U37655 (N_37655,N_31635,N_34261);
xor U37656 (N_37656,N_34313,N_30146);
nand U37657 (N_37657,N_31960,N_33885);
and U37658 (N_37658,N_30404,N_33901);
or U37659 (N_37659,N_34374,N_30204);
nor U37660 (N_37660,N_32869,N_34557);
nor U37661 (N_37661,N_33025,N_34876);
nand U37662 (N_37662,N_33440,N_32034);
or U37663 (N_37663,N_30777,N_32645);
or U37664 (N_37664,N_32390,N_33214);
nand U37665 (N_37665,N_30725,N_33525);
and U37666 (N_37666,N_34673,N_34109);
and U37667 (N_37667,N_34014,N_32994);
xnor U37668 (N_37668,N_31262,N_31597);
and U37669 (N_37669,N_33972,N_30838);
or U37670 (N_37670,N_34250,N_33857);
nand U37671 (N_37671,N_30037,N_33192);
nand U37672 (N_37672,N_33690,N_33578);
and U37673 (N_37673,N_31584,N_31049);
and U37674 (N_37674,N_32900,N_30648);
xor U37675 (N_37675,N_33209,N_30247);
xnor U37676 (N_37676,N_31559,N_33772);
nor U37677 (N_37677,N_33773,N_32880);
or U37678 (N_37678,N_31450,N_33696);
and U37679 (N_37679,N_33667,N_30800);
nor U37680 (N_37680,N_31322,N_33426);
and U37681 (N_37681,N_30802,N_34324);
nor U37682 (N_37682,N_30484,N_34667);
and U37683 (N_37683,N_30125,N_33363);
nand U37684 (N_37684,N_34959,N_34789);
nand U37685 (N_37685,N_34191,N_31026);
or U37686 (N_37686,N_30601,N_30633);
xor U37687 (N_37687,N_30732,N_31032);
nand U37688 (N_37688,N_31192,N_34989);
nand U37689 (N_37689,N_30644,N_31514);
nor U37690 (N_37690,N_34506,N_30319);
nor U37691 (N_37691,N_34661,N_34475);
xnor U37692 (N_37692,N_30708,N_32173);
xnor U37693 (N_37693,N_31493,N_32775);
xnor U37694 (N_37694,N_34364,N_31993);
nand U37695 (N_37695,N_30202,N_31422);
or U37696 (N_37696,N_31708,N_32155);
and U37697 (N_37697,N_32223,N_32252);
nand U37698 (N_37698,N_33982,N_30780);
and U37699 (N_37699,N_34279,N_34385);
or U37700 (N_37700,N_34553,N_31869);
and U37701 (N_37701,N_31852,N_34251);
nand U37702 (N_37702,N_33721,N_34828);
or U37703 (N_37703,N_30032,N_30101);
xnor U37704 (N_37704,N_33069,N_30537);
nor U37705 (N_37705,N_30032,N_30535);
nor U37706 (N_37706,N_34366,N_31278);
or U37707 (N_37707,N_33789,N_31493);
and U37708 (N_37708,N_33439,N_34305);
nand U37709 (N_37709,N_33195,N_32705);
or U37710 (N_37710,N_33028,N_33940);
nand U37711 (N_37711,N_30868,N_30228);
nand U37712 (N_37712,N_31043,N_34745);
and U37713 (N_37713,N_31689,N_32586);
and U37714 (N_37714,N_30579,N_34840);
xnor U37715 (N_37715,N_34908,N_30843);
nand U37716 (N_37716,N_33295,N_34453);
and U37717 (N_37717,N_32851,N_32036);
xor U37718 (N_37718,N_32877,N_33345);
nor U37719 (N_37719,N_30000,N_31573);
nand U37720 (N_37720,N_30030,N_32949);
xnor U37721 (N_37721,N_33883,N_32640);
or U37722 (N_37722,N_34689,N_30116);
xnor U37723 (N_37723,N_34678,N_34858);
and U37724 (N_37724,N_30099,N_34116);
xor U37725 (N_37725,N_31649,N_31834);
nor U37726 (N_37726,N_31683,N_34521);
or U37727 (N_37727,N_33283,N_30558);
or U37728 (N_37728,N_30047,N_34270);
or U37729 (N_37729,N_34031,N_31072);
or U37730 (N_37730,N_30859,N_30918);
xnor U37731 (N_37731,N_30543,N_34009);
xnor U37732 (N_37732,N_34492,N_34943);
and U37733 (N_37733,N_34539,N_31577);
nand U37734 (N_37734,N_32549,N_33690);
nand U37735 (N_37735,N_30070,N_30103);
or U37736 (N_37736,N_32961,N_32718);
and U37737 (N_37737,N_34311,N_30024);
or U37738 (N_37738,N_33756,N_33716);
nand U37739 (N_37739,N_34256,N_32769);
nor U37740 (N_37740,N_30471,N_33859);
nand U37741 (N_37741,N_34829,N_30583);
nor U37742 (N_37742,N_30037,N_31070);
or U37743 (N_37743,N_32885,N_33944);
or U37744 (N_37744,N_34608,N_31089);
xnor U37745 (N_37745,N_31107,N_30933);
nand U37746 (N_37746,N_32756,N_30544);
nor U37747 (N_37747,N_30240,N_33924);
and U37748 (N_37748,N_30089,N_31079);
or U37749 (N_37749,N_32491,N_34186);
xnor U37750 (N_37750,N_33432,N_33965);
xor U37751 (N_37751,N_30563,N_33700);
nor U37752 (N_37752,N_34789,N_33747);
and U37753 (N_37753,N_32708,N_30022);
nor U37754 (N_37754,N_31111,N_33694);
nand U37755 (N_37755,N_32106,N_34561);
nor U37756 (N_37756,N_34638,N_34697);
nor U37757 (N_37757,N_32541,N_33113);
or U37758 (N_37758,N_30563,N_30835);
and U37759 (N_37759,N_30139,N_34397);
or U37760 (N_37760,N_32103,N_34398);
and U37761 (N_37761,N_31813,N_32356);
and U37762 (N_37762,N_31427,N_32383);
xor U37763 (N_37763,N_34684,N_30264);
xor U37764 (N_37764,N_31235,N_30924);
and U37765 (N_37765,N_30159,N_33334);
or U37766 (N_37766,N_34486,N_31680);
or U37767 (N_37767,N_32429,N_32870);
nor U37768 (N_37768,N_33245,N_30020);
or U37769 (N_37769,N_32330,N_30757);
or U37770 (N_37770,N_30367,N_31319);
nand U37771 (N_37771,N_33958,N_34623);
xnor U37772 (N_37772,N_32560,N_33549);
or U37773 (N_37773,N_30375,N_30573);
nor U37774 (N_37774,N_31263,N_34524);
xor U37775 (N_37775,N_34403,N_34528);
nor U37776 (N_37776,N_30435,N_33227);
or U37777 (N_37777,N_32010,N_34430);
or U37778 (N_37778,N_31664,N_34396);
nand U37779 (N_37779,N_32892,N_34954);
and U37780 (N_37780,N_34354,N_33858);
xnor U37781 (N_37781,N_31708,N_32544);
xor U37782 (N_37782,N_31191,N_32618);
nand U37783 (N_37783,N_34929,N_32015);
or U37784 (N_37784,N_34810,N_30395);
and U37785 (N_37785,N_32247,N_34588);
nand U37786 (N_37786,N_34489,N_30477);
nand U37787 (N_37787,N_30863,N_33591);
xnor U37788 (N_37788,N_30520,N_34560);
nand U37789 (N_37789,N_32654,N_32726);
nand U37790 (N_37790,N_31678,N_34032);
nand U37791 (N_37791,N_33002,N_31261);
or U37792 (N_37792,N_30404,N_33366);
xnor U37793 (N_37793,N_33279,N_32784);
and U37794 (N_37794,N_30041,N_31256);
xor U37795 (N_37795,N_31475,N_30581);
and U37796 (N_37796,N_34398,N_33065);
and U37797 (N_37797,N_31855,N_32130);
nand U37798 (N_37798,N_34212,N_30914);
nor U37799 (N_37799,N_32159,N_30889);
and U37800 (N_37800,N_30337,N_31763);
nor U37801 (N_37801,N_31076,N_30404);
or U37802 (N_37802,N_30307,N_30176);
xnor U37803 (N_37803,N_32178,N_33148);
xor U37804 (N_37804,N_33211,N_34028);
nor U37805 (N_37805,N_33008,N_34517);
nor U37806 (N_37806,N_34337,N_34688);
xnor U37807 (N_37807,N_32412,N_33485);
and U37808 (N_37808,N_30838,N_33621);
nand U37809 (N_37809,N_31081,N_34214);
or U37810 (N_37810,N_31156,N_34098);
and U37811 (N_37811,N_33657,N_34993);
and U37812 (N_37812,N_32751,N_30231);
nor U37813 (N_37813,N_34350,N_33142);
nand U37814 (N_37814,N_34758,N_30430);
or U37815 (N_37815,N_30838,N_34027);
nor U37816 (N_37816,N_32251,N_30942);
and U37817 (N_37817,N_30430,N_31303);
and U37818 (N_37818,N_30717,N_34228);
xor U37819 (N_37819,N_32470,N_33776);
or U37820 (N_37820,N_34831,N_32902);
xnor U37821 (N_37821,N_32128,N_33307);
xor U37822 (N_37822,N_33347,N_31742);
nand U37823 (N_37823,N_34686,N_33776);
nor U37824 (N_37824,N_31664,N_30134);
or U37825 (N_37825,N_31419,N_32994);
or U37826 (N_37826,N_31069,N_32259);
or U37827 (N_37827,N_34628,N_30441);
xor U37828 (N_37828,N_33468,N_31449);
or U37829 (N_37829,N_31877,N_30382);
nor U37830 (N_37830,N_31389,N_34195);
or U37831 (N_37831,N_34343,N_31355);
and U37832 (N_37832,N_32267,N_31342);
xor U37833 (N_37833,N_33911,N_31757);
and U37834 (N_37834,N_31964,N_33764);
or U37835 (N_37835,N_31221,N_32674);
nor U37836 (N_37836,N_32046,N_30329);
and U37837 (N_37837,N_34841,N_32947);
and U37838 (N_37838,N_30589,N_30936);
nor U37839 (N_37839,N_31430,N_32294);
nand U37840 (N_37840,N_31611,N_33542);
or U37841 (N_37841,N_33075,N_30766);
xnor U37842 (N_37842,N_30756,N_31622);
nor U37843 (N_37843,N_30431,N_30658);
nand U37844 (N_37844,N_34276,N_31999);
xor U37845 (N_37845,N_34423,N_31089);
and U37846 (N_37846,N_33195,N_32649);
xnor U37847 (N_37847,N_31850,N_31136);
or U37848 (N_37848,N_32102,N_34656);
nor U37849 (N_37849,N_31699,N_31950);
or U37850 (N_37850,N_34805,N_31583);
nand U37851 (N_37851,N_32178,N_30856);
xnor U37852 (N_37852,N_31152,N_34464);
nor U37853 (N_37853,N_34781,N_31622);
or U37854 (N_37854,N_33930,N_31327);
nand U37855 (N_37855,N_32129,N_34049);
and U37856 (N_37856,N_34929,N_33955);
and U37857 (N_37857,N_34981,N_31516);
and U37858 (N_37858,N_32509,N_33606);
nand U37859 (N_37859,N_30336,N_32544);
or U37860 (N_37860,N_34359,N_34158);
and U37861 (N_37861,N_31860,N_31446);
xor U37862 (N_37862,N_30749,N_30158);
nand U37863 (N_37863,N_30628,N_31007);
and U37864 (N_37864,N_30595,N_32490);
nor U37865 (N_37865,N_32556,N_32618);
and U37866 (N_37866,N_31827,N_30566);
nor U37867 (N_37867,N_31973,N_33233);
xnor U37868 (N_37868,N_30444,N_34049);
and U37869 (N_37869,N_32295,N_34185);
nor U37870 (N_37870,N_32698,N_34831);
or U37871 (N_37871,N_34309,N_33971);
or U37872 (N_37872,N_32447,N_33914);
nor U37873 (N_37873,N_31584,N_33874);
nor U37874 (N_37874,N_30578,N_32630);
nand U37875 (N_37875,N_33782,N_33555);
or U37876 (N_37876,N_32979,N_34709);
nand U37877 (N_37877,N_34188,N_32424);
or U37878 (N_37878,N_33055,N_33424);
or U37879 (N_37879,N_34557,N_34708);
nor U37880 (N_37880,N_32078,N_33574);
nor U37881 (N_37881,N_32977,N_30947);
nor U37882 (N_37882,N_30313,N_33845);
nand U37883 (N_37883,N_33179,N_31208);
nand U37884 (N_37884,N_31669,N_33468);
or U37885 (N_37885,N_32713,N_33038);
nand U37886 (N_37886,N_34006,N_31176);
or U37887 (N_37887,N_31102,N_30087);
nand U37888 (N_37888,N_33358,N_33105);
nand U37889 (N_37889,N_31933,N_34975);
and U37890 (N_37890,N_32854,N_31686);
nand U37891 (N_37891,N_32570,N_31362);
nand U37892 (N_37892,N_31028,N_34095);
xnor U37893 (N_37893,N_34115,N_34924);
nor U37894 (N_37894,N_32835,N_31592);
xnor U37895 (N_37895,N_34349,N_32369);
or U37896 (N_37896,N_30463,N_33415);
or U37897 (N_37897,N_30828,N_32382);
nand U37898 (N_37898,N_31151,N_33580);
nor U37899 (N_37899,N_32573,N_34181);
nor U37900 (N_37900,N_32326,N_33977);
nor U37901 (N_37901,N_31491,N_31322);
nor U37902 (N_37902,N_33327,N_30140);
and U37903 (N_37903,N_34532,N_30560);
and U37904 (N_37904,N_34357,N_33209);
nand U37905 (N_37905,N_34971,N_31947);
or U37906 (N_37906,N_34148,N_30655);
and U37907 (N_37907,N_32747,N_30796);
and U37908 (N_37908,N_31616,N_32097);
nand U37909 (N_37909,N_32961,N_32054);
and U37910 (N_37910,N_33991,N_34543);
nor U37911 (N_37911,N_31155,N_34716);
nand U37912 (N_37912,N_32161,N_34125);
or U37913 (N_37913,N_33311,N_32617);
xnor U37914 (N_37914,N_31227,N_30197);
xor U37915 (N_37915,N_32405,N_31760);
and U37916 (N_37916,N_30389,N_32674);
nand U37917 (N_37917,N_34364,N_30060);
and U37918 (N_37918,N_34990,N_33739);
nor U37919 (N_37919,N_34471,N_33015);
nor U37920 (N_37920,N_30574,N_32353);
and U37921 (N_37921,N_31977,N_32297);
and U37922 (N_37922,N_33143,N_31641);
and U37923 (N_37923,N_31999,N_31186);
nor U37924 (N_37924,N_32408,N_30446);
nand U37925 (N_37925,N_33900,N_33091);
xnor U37926 (N_37926,N_34022,N_32825);
or U37927 (N_37927,N_34255,N_33276);
or U37928 (N_37928,N_30065,N_31209);
nand U37929 (N_37929,N_33423,N_31633);
nand U37930 (N_37930,N_30993,N_32827);
nor U37931 (N_37931,N_32752,N_30881);
or U37932 (N_37932,N_30155,N_34476);
xnor U37933 (N_37933,N_30357,N_32504);
or U37934 (N_37934,N_31776,N_34811);
nand U37935 (N_37935,N_34802,N_33206);
and U37936 (N_37936,N_30891,N_30300);
and U37937 (N_37937,N_34763,N_30663);
nor U37938 (N_37938,N_33235,N_34107);
and U37939 (N_37939,N_31205,N_30985);
nor U37940 (N_37940,N_33621,N_32768);
or U37941 (N_37941,N_33852,N_31271);
or U37942 (N_37942,N_34370,N_34381);
nor U37943 (N_37943,N_30270,N_30662);
nand U37944 (N_37944,N_30458,N_32086);
xor U37945 (N_37945,N_33590,N_32582);
nor U37946 (N_37946,N_34492,N_30900);
nor U37947 (N_37947,N_31108,N_31961);
and U37948 (N_37948,N_33215,N_32556);
nor U37949 (N_37949,N_32804,N_30302);
nor U37950 (N_37950,N_31123,N_30743);
nand U37951 (N_37951,N_31957,N_30521);
nand U37952 (N_37952,N_34940,N_34058);
and U37953 (N_37953,N_31584,N_30296);
nand U37954 (N_37954,N_32349,N_33149);
or U37955 (N_37955,N_32540,N_30195);
and U37956 (N_37956,N_30601,N_33870);
xnor U37957 (N_37957,N_33910,N_30486);
nor U37958 (N_37958,N_30496,N_31900);
nor U37959 (N_37959,N_32438,N_30789);
nor U37960 (N_37960,N_33046,N_30361);
xor U37961 (N_37961,N_31425,N_34858);
or U37962 (N_37962,N_31339,N_30952);
nand U37963 (N_37963,N_31550,N_30128);
or U37964 (N_37964,N_34334,N_32945);
xor U37965 (N_37965,N_32381,N_34468);
nand U37966 (N_37966,N_34069,N_33432);
nand U37967 (N_37967,N_33087,N_31412);
and U37968 (N_37968,N_32272,N_30952);
or U37969 (N_37969,N_30637,N_31080);
and U37970 (N_37970,N_32717,N_33133);
nand U37971 (N_37971,N_30988,N_34823);
nor U37972 (N_37972,N_31091,N_32839);
nor U37973 (N_37973,N_34648,N_30198);
and U37974 (N_37974,N_31608,N_32867);
xnor U37975 (N_37975,N_30614,N_30444);
nor U37976 (N_37976,N_30737,N_33070);
xor U37977 (N_37977,N_32157,N_32487);
xnor U37978 (N_37978,N_32181,N_34951);
or U37979 (N_37979,N_33619,N_32896);
nor U37980 (N_37980,N_32723,N_34432);
nor U37981 (N_37981,N_34924,N_30042);
and U37982 (N_37982,N_34894,N_33860);
and U37983 (N_37983,N_34983,N_30320);
nand U37984 (N_37984,N_30767,N_33397);
nand U37985 (N_37985,N_31407,N_31725);
and U37986 (N_37986,N_34353,N_33284);
or U37987 (N_37987,N_31044,N_32985);
nor U37988 (N_37988,N_32043,N_33687);
or U37989 (N_37989,N_30661,N_34532);
and U37990 (N_37990,N_31559,N_31447);
xor U37991 (N_37991,N_33932,N_33857);
nand U37992 (N_37992,N_32316,N_30695);
and U37993 (N_37993,N_34588,N_30377);
xnor U37994 (N_37994,N_31135,N_31621);
and U37995 (N_37995,N_32153,N_34110);
xnor U37996 (N_37996,N_33338,N_33445);
nand U37997 (N_37997,N_30146,N_33762);
and U37998 (N_37998,N_33683,N_30514);
nor U37999 (N_37999,N_33686,N_31229);
nand U38000 (N_38000,N_31922,N_31548);
and U38001 (N_38001,N_31875,N_33126);
or U38002 (N_38002,N_32505,N_32037);
or U38003 (N_38003,N_31354,N_32498);
nand U38004 (N_38004,N_33894,N_32468);
xnor U38005 (N_38005,N_33671,N_31207);
nor U38006 (N_38006,N_34259,N_32094);
and U38007 (N_38007,N_32174,N_30898);
xor U38008 (N_38008,N_30601,N_32133);
xnor U38009 (N_38009,N_34979,N_34341);
nand U38010 (N_38010,N_30891,N_32397);
xnor U38011 (N_38011,N_34149,N_30291);
xnor U38012 (N_38012,N_31363,N_32932);
nand U38013 (N_38013,N_34045,N_30786);
xor U38014 (N_38014,N_33509,N_34367);
xor U38015 (N_38015,N_33057,N_30906);
nand U38016 (N_38016,N_31609,N_32810);
and U38017 (N_38017,N_32421,N_34596);
or U38018 (N_38018,N_33441,N_30491);
nor U38019 (N_38019,N_31814,N_32575);
nor U38020 (N_38020,N_32916,N_30417);
or U38021 (N_38021,N_30668,N_31205);
nand U38022 (N_38022,N_34428,N_30890);
nor U38023 (N_38023,N_32763,N_33164);
and U38024 (N_38024,N_30693,N_31932);
and U38025 (N_38025,N_32714,N_31755);
and U38026 (N_38026,N_30139,N_30132);
and U38027 (N_38027,N_31809,N_34073);
nor U38028 (N_38028,N_33015,N_34523);
nand U38029 (N_38029,N_30559,N_34027);
or U38030 (N_38030,N_34776,N_32651);
nand U38031 (N_38031,N_33062,N_32356);
nor U38032 (N_38032,N_32942,N_32659);
nand U38033 (N_38033,N_34041,N_34611);
or U38034 (N_38034,N_32685,N_31286);
xnor U38035 (N_38035,N_30219,N_34284);
xor U38036 (N_38036,N_30635,N_34736);
nor U38037 (N_38037,N_32848,N_34415);
nor U38038 (N_38038,N_31574,N_30556);
and U38039 (N_38039,N_30980,N_32376);
nand U38040 (N_38040,N_30972,N_31944);
or U38041 (N_38041,N_34439,N_32997);
nand U38042 (N_38042,N_32125,N_31218);
and U38043 (N_38043,N_32805,N_33847);
and U38044 (N_38044,N_32351,N_32925);
nor U38045 (N_38045,N_33168,N_31134);
and U38046 (N_38046,N_31623,N_33349);
nand U38047 (N_38047,N_32795,N_34323);
xor U38048 (N_38048,N_32526,N_31127);
or U38049 (N_38049,N_33330,N_31616);
nor U38050 (N_38050,N_32184,N_32185);
or U38051 (N_38051,N_30153,N_31862);
and U38052 (N_38052,N_32663,N_33131);
nand U38053 (N_38053,N_32877,N_34620);
and U38054 (N_38054,N_31339,N_32621);
xnor U38055 (N_38055,N_30941,N_30124);
and U38056 (N_38056,N_34608,N_34658);
nor U38057 (N_38057,N_30310,N_30687);
nand U38058 (N_38058,N_31117,N_34912);
nand U38059 (N_38059,N_34993,N_30413);
and U38060 (N_38060,N_30537,N_32553);
xnor U38061 (N_38061,N_34124,N_32343);
nor U38062 (N_38062,N_32934,N_33402);
xor U38063 (N_38063,N_32130,N_34785);
and U38064 (N_38064,N_31484,N_31460);
nor U38065 (N_38065,N_33309,N_34664);
nor U38066 (N_38066,N_34255,N_33781);
or U38067 (N_38067,N_31588,N_33858);
nand U38068 (N_38068,N_33449,N_32742);
and U38069 (N_38069,N_30729,N_32570);
nor U38070 (N_38070,N_31368,N_32928);
or U38071 (N_38071,N_33678,N_31470);
and U38072 (N_38072,N_33613,N_33517);
and U38073 (N_38073,N_32445,N_32603);
or U38074 (N_38074,N_33147,N_33643);
nor U38075 (N_38075,N_30384,N_32835);
nor U38076 (N_38076,N_30915,N_32711);
and U38077 (N_38077,N_32597,N_30163);
nor U38078 (N_38078,N_34966,N_31432);
or U38079 (N_38079,N_30122,N_32093);
nand U38080 (N_38080,N_30267,N_34055);
or U38081 (N_38081,N_32486,N_33919);
xor U38082 (N_38082,N_31740,N_32970);
nand U38083 (N_38083,N_33467,N_33549);
or U38084 (N_38084,N_34487,N_33682);
nand U38085 (N_38085,N_31726,N_34473);
or U38086 (N_38086,N_30314,N_30500);
or U38087 (N_38087,N_32975,N_31833);
or U38088 (N_38088,N_33396,N_30075);
or U38089 (N_38089,N_33677,N_31174);
and U38090 (N_38090,N_33321,N_30637);
or U38091 (N_38091,N_31274,N_33893);
and U38092 (N_38092,N_32643,N_33064);
or U38093 (N_38093,N_33789,N_33227);
or U38094 (N_38094,N_32820,N_33904);
nor U38095 (N_38095,N_33977,N_30392);
nor U38096 (N_38096,N_34257,N_32728);
and U38097 (N_38097,N_34406,N_31799);
nor U38098 (N_38098,N_32032,N_32015);
nor U38099 (N_38099,N_32681,N_34171);
xnor U38100 (N_38100,N_34982,N_31430);
xnor U38101 (N_38101,N_34471,N_34057);
or U38102 (N_38102,N_31422,N_32487);
or U38103 (N_38103,N_30561,N_31210);
and U38104 (N_38104,N_32960,N_32483);
xnor U38105 (N_38105,N_31541,N_31434);
and U38106 (N_38106,N_31455,N_30435);
nand U38107 (N_38107,N_32226,N_32164);
xor U38108 (N_38108,N_33703,N_33964);
nor U38109 (N_38109,N_30303,N_31123);
nor U38110 (N_38110,N_31699,N_34457);
xor U38111 (N_38111,N_33288,N_31887);
or U38112 (N_38112,N_30649,N_30439);
xor U38113 (N_38113,N_33410,N_30113);
nand U38114 (N_38114,N_32639,N_31915);
and U38115 (N_38115,N_34441,N_31521);
nand U38116 (N_38116,N_31433,N_30800);
and U38117 (N_38117,N_30531,N_34589);
and U38118 (N_38118,N_34707,N_32921);
and U38119 (N_38119,N_31349,N_32702);
nand U38120 (N_38120,N_32597,N_30843);
and U38121 (N_38121,N_31964,N_30527);
xnor U38122 (N_38122,N_32778,N_34744);
xnor U38123 (N_38123,N_34649,N_34730);
nand U38124 (N_38124,N_34811,N_31496);
and U38125 (N_38125,N_32997,N_34850);
xnor U38126 (N_38126,N_34470,N_34372);
and U38127 (N_38127,N_33861,N_30080);
or U38128 (N_38128,N_34317,N_34398);
xor U38129 (N_38129,N_31564,N_32708);
nor U38130 (N_38130,N_32991,N_34334);
or U38131 (N_38131,N_33923,N_32050);
nor U38132 (N_38132,N_30162,N_30223);
or U38133 (N_38133,N_30878,N_31484);
or U38134 (N_38134,N_32370,N_31921);
and U38135 (N_38135,N_30667,N_32235);
xnor U38136 (N_38136,N_30922,N_30375);
and U38137 (N_38137,N_33082,N_30486);
xnor U38138 (N_38138,N_34380,N_30530);
and U38139 (N_38139,N_33613,N_32793);
nor U38140 (N_38140,N_30832,N_34453);
nor U38141 (N_38141,N_30136,N_33296);
and U38142 (N_38142,N_34968,N_30016);
and U38143 (N_38143,N_30181,N_32153);
nand U38144 (N_38144,N_33235,N_30249);
or U38145 (N_38145,N_31978,N_31221);
xor U38146 (N_38146,N_33459,N_33504);
or U38147 (N_38147,N_30287,N_31771);
or U38148 (N_38148,N_30152,N_32089);
nor U38149 (N_38149,N_34361,N_33693);
and U38150 (N_38150,N_30298,N_33921);
nor U38151 (N_38151,N_30799,N_32297);
and U38152 (N_38152,N_32011,N_33982);
or U38153 (N_38153,N_31505,N_34071);
and U38154 (N_38154,N_33760,N_30542);
xnor U38155 (N_38155,N_34652,N_33177);
nand U38156 (N_38156,N_33387,N_31670);
nor U38157 (N_38157,N_31137,N_34042);
or U38158 (N_38158,N_33889,N_31094);
xor U38159 (N_38159,N_30656,N_34980);
or U38160 (N_38160,N_34425,N_33295);
nor U38161 (N_38161,N_33791,N_33038);
nor U38162 (N_38162,N_30847,N_33482);
or U38163 (N_38163,N_31173,N_30006);
nand U38164 (N_38164,N_30718,N_30354);
nor U38165 (N_38165,N_34454,N_31406);
or U38166 (N_38166,N_32325,N_34688);
nand U38167 (N_38167,N_32870,N_30771);
and U38168 (N_38168,N_30367,N_30056);
and U38169 (N_38169,N_32583,N_33631);
xor U38170 (N_38170,N_31452,N_30778);
nor U38171 (N_38171,N_33601,N_33257);
xnor U38172 (N_38172,N_30840,N_33153);
nor U38173 (N_38173,N_31570,N_31202);
nand U38174 (N_38174,N_31499,N_33413);
or U38175 (N_38175,N_32952,N_33995);
nor U38176 (N_38176,N_30296,N_33533);
and U38177 (N_38177,N_31619,N_34096);
nor U38178 (N_38178,N_34030,N_30218);
nand U38179 (N_38179,N_31137,N_32957);
or U38180 (N_38180,N_30923,N_34410);
nand U38181 (N_38181,N_32665,N_33554);
or U38182 (N_38182,N_30263,N_31419);
nor U38183 (N_38183,N_32255,N_32744);
or U38184 (N_38184,N_30205,N_31151);
xnor U38185 (N_38185,N_33807,N_32661);
xor U38186 (N_38186,N_32907,N_31030);
or U38187 (N_38187,N_30434,N_30942);
or U38188 (N_38188,N_31623,N_30406);
nor U38189 (N_38189,N_33943,N_34546);
nor U38190 (N_38190,N_30324,N_32169);
nand U38191 (N_38191,N_30324,N_34795);
xnor U38192 (N_38192,N_30286,N_34495);
or U38193 (N_38193,N_32408,N_32065);
and U38194 (N_38194,N_33681,N_34233);
or U38195 (N_38195,N_30689,N_32152);
nor U38196 (N_38196,N_33006,N_32225);
xor U38197 (N_38197,N_33005,N_33508);
or U38198 (N_38198,N_32583,N_30095);
nand U38199 (N_38199,N_31537,N_30429);
nor U38200 (N_38200,N_31396,N_33677);
xnor U38201 (N_38201,N_34928,N_34927);
and U38202 (N_38202,N_33737,N_33106);
nand U38203 (N_38203,N_31101,N_34737);
xor U38204 (N_38204,N_30201,N_30736);
xor U38205 (N_38205,N_32254,N_34873);
and U38206 (N_38206,N_33798,N_32448);
or U38207 (N_38207,N_32951,N_30671);
xor U38208 (N_38208,N_30193,N_31255);
and U38209 (N_38209,N_30854,N_31199);
and U38210 (N_38210,N_30763,N_32821);
or U38211 (N_38211,N_32790,N_34519);
nand U38212 (N_38212,N_30822,N_34491);
and U38213 (N_38213,N_30613,N_34733);
nand U38214 (N_38214,N_34735,N_31277);
nor U38215 (N_38215,N_32997,N_31928);
and U38216 (N_38216,N_32604,N_31280);
nor U38217 (N_38217,N_30927,N_33482);
xnor U38218 (N_38218,N_31351,N_34012);
and U38219 (N_38219,N_34758,N_32279);
nand U38220 (N_38220,N_30256,N_31145);
xor U38221 (N_38221,N_33426,N_34484);
and U38222 (N_38222,N_33015,N_34289);
xnor U38223 (N_38223,N_31568,N_33705);
xnor U38224 (N_38224,N_30874,N_32203);
xnor U38225 (N_38225,N_32908,N_32117);
xnor U38226 (N_38226,N_30468,N_34748);
and U38227 (N_38227,N_33583,N_33994);
nand U38228 (N_38228,N_34348,N_31826);
xor U38229 (N_38229,N_30029,N_30072);
xor U38230 (N_38230,N_34278,N_33352);
and U38231 (N_38231,N_32307,N_30374);
nand U38232 (N_38232,N_31605,N_34372);
nand U38233 (N_38233,N_30830,N_33381);
nand U38234 (N_38234,N_34096,N_33244);
xor U38235 (N_38235,N_31795,N_32334);
or U38236 (N_38236,N_34335,N_34156);
nor U38237 (N_38237,N_33379,N_30087);
nor U38238 (N_38238,N_32659,N_32138);
xor U38239 (N_38239,N_31012,N_33934);
and U38240 (N_38240,N_33258,N_33245);
nor U38241 (N_38241,N_30102,N_32951);
nor U38242 (N_38242,N_33490,N_33076);
or U38243 (N_38243,N_32079,N_30734);
nor U38244 (N_38244,N_33567,N_32494);
xor U38245 (N_38245,N_33937,N_33535);
xnor U38246 (N_38246,N_30576,N_33510);
and U38247 (N_38247,N_32230,N_33323);
nand U38248 (N_38248,N_32972,N_30823);
or U38249 (N_38249,N_32186,N_33502);
nand U38250 (N_38250,N_30537,N_30678);
and U38251 (N_38251,N_30519,N_32326);
or U38252 (N_38252,N_30806,N_30813);
or U38253 (N_38253,N_30857,N_30460);
nor U38254 (N_38254,N_33413,N_30001);
or U38255 (N_38255,N_32404,N_34361);
or U38256 (N_38256,N_30144,N_31790);
nand U38257 (N_38257,N_30794,N_32594);
nand U38258 (N_38258,N_32935,N_30683);
nor U38259 (N_38259,N_30742,N_31284);
and U38260 (N_38260,N_32669,N_30924);
and U38261 (N_38261,N_34128,N_33670);
or U38262 (N_38262,N_33526,N_33479);
or U38263 (N_38263,N_32927,N_30197);
xnor U38264 (N_38264,N_32247,N_34948);
xor U38265 (N_38265,N_33993,N_34150);
xor U38266 (N_38266,N_34399,N_33222);
nor U38267 (N_38267,N_31962,N_31427);
and U38268 (N_38268,N_31739,N_34622);
nand U38269 (N_38269,N_32707,N_34446);
nor U38270 (N_38270,N_31429,N_30818);
and U38271 (N_38271,N_33216,N_34579);
or U38272 (N_38272,N_32737,N_34807);
nand U38273 (N_38273,N_30409,N_32479);
and U38274 (N_38274,N_34394,N_34938);
or U38275 (N_38275,N_33974,N_30621);
and U38276 (N_38276,N_34005,N_31373);
or U38277 (N_38277,N_32169,N_30182);
nand U38278 (N_38278,N_33472,N_33575);
nor U38279 (N_38279,N_33398,N_34180);
nor U38280 (N_38280,N_34626,N_34215);
nand U38281 (N_38281,N_33221,N_33473);
and U38282 (N_38282,N_34202,N_34270);
and U38283 (N_38283,N_34275,N_30119);
and U38284 (N_38284,N_33837,N_31522);
or U38285 (N_38285,N_31079,N_33571);
nand U38286 (N_38286,N_34494,N_32040);
and U38287 (N_38287,N_33867,N_31255);
xor U38288 (N_38288,N_32601,N_30043);
xnor U38289 (N_38289,N_31836,N_32290);
nor U38290 (N_38290,N_30266,N_30511);
and U38291 (N_38291,N_32303,N_34137);
xor U38292 (N_38292,N_33734,N_33569);
xnor U38293 (N_38293,N_30832,N_30849);
or U38294 (N_38294,N_30349,N_30849);
nor U38295 (N_38295,N_31841,N_34428);
or U38296 (N_38296,N_31937,N_30150);
nand U38297 (N_38297,N_34888,N_30512);
or U38298 (N_38298,N_30729,N_32106);
or U38299 (N_38299,N_33928,N_30824);
nand U38300 (N_38300,N_31937,N_34369);
nand U38301 (N_38301,N_30341,N_31882);
nand U38302 (N_38302,N_31613,N_30427);
nand U38303 (N_38303,N_33594,N_32352);
nand U38304 (N_38304,N_34325,N_33993);
xnor U38305 (N_38305,N_33060,N_33058);
nand U38306 (N_38306,N_31759,N_32698);
and U38307 (N_38307,N_30356,N_33865);
nor U38308 (N_38308,N_30731,N_32733);
and U38309 (N_38309,N_33321,N_30974);
and U38310 (N_38310,N_33505,N_33831);
or U38311 (N_38311,N_33633,N_31022);
xor U38312 (N_38312,N_31631,N_31750);
nor U38313 (N_38313,N_31265,N_33978);
xnor U38314 (N_38314,N_32070,N_30964);
and U38315 (N_38315,N_32667,N_31121);
or U38316 (N_38316,N_31657,N_33961);
nor U38317 (N_38317,N_33849,N_32423);
or U38318 (N_38318,N_31607,N_31293);
and U38319 (N_38319,N_30750,N_32636);
or U38320 (N_38320,N_34696,N_31737);
and U38321 (N_38321,N_33600,N_31374);
nor U38322 (N_38322,N_33783,N_33157);
nor U38323 (N_38323,N_32661,N_31061);
nor U38324 (N_38324,N_31453,N_34506);
and U38325 (N_38325,N_34176,N_33834);
nor U38326 (N_38326,N_32043,N_30729);
xor U38327 (N_38327,N_30501,N_32633);
nand U38328 (N_38328,N_33575,N_34608);
nand U38329 (N_38329,N_32870,N_34659);
nor U38330 (N_38330,N_31389,N_32095);
nor U38331 (N_38331,N_30555,N_30989);
nand U38332 (N_38332,N_33773,N_31957);
and U38333 (N_38333,N_34283,N_33196);
nand U38334 (N_38334,N_31929,N_30944);
xnor U38335 (N_38335,N_30099,N_32556);
or U38336 (N_38336,N_31679,N_32229);
nor U38337 (N_38337,N_34632,N_34053);
nand U38338 (N_38338,N_30043,N_33913);
nor U38339 (N_38339,N_32289,N_31085);
or U38340 (N_38340,N_32660,N_31780);
xor U38341 (N_38341,N_31075,N_32033);
xor U38342 (N_38342,N_31958,N_33558);
and U38343 (N_38343,N_30824,N_31565);
xor U38344 (N_38344,N_34838,N_33835);
xnor U38345 (N_38345,N_31163,N_33671);
xnor U38346 (N_38346,N_32411,N_32491);
or U38347 (N_38347,N_31894,N_33634);
nand U38348 (N_38348,N_34370,N_34353);
xnor U38349 (N_38349,N_32524,N_30531);
or U38350 (N_38350,N_34446,N_32603);
xnor U38351 (N_38351,N_32811,N_32391);
and U38352 (N_38352,N_34866,N_34970);
xor U38353 (N_38353,N_30709,N_32903);
and U38354 (N_38354,N_30411,N_34196);
xnor U38355 (N_38355,N_32704,N_33959);
or U38356 (N_38356,N_31925,N_34813);
or U38357 (N_38357,N_34131,N_30665);
nor U38358 (N_38358,N_30261,N_32142);
nor U38359 (N_38359,N_34319,N_32562);
nand U38360 (N_38360,N_34129,N_34135);
nand U38361 (N_38361,N_34821,N_31691);
xnor U38362 (N_38362,N_33991,N_30964);
or U38363 (N_38363,N_30653,N_32407);
or U38364 (N_38364,N_32119,N_34206);
nor U38365 (N_38365,N_33262,N_30828);
and U38366 (N_38366,N_34176,N_34637);
nor U38367 (N_38367,N_33825,N_30056);
nand U38368 (N_38368,N_31870,N_33326);
or U38369 (N_38369,N_34134,N_32215);
nor U38370 (N_38370,N_32578,N_34449);
or U38371 (N_38371,N_33724,N_34138);
xor U38372 (N_38372,N_34847,N_30359);
nand U38373 (N_38373,N_30901,N_32220);
and U38374 (N_38374,N_30344,N_31167);
nand U38375 (N_38375,N_31045,N_32890);
or U38376 (N_38376,N_32367,N_32434);
xor U38377 (N_38377,N_34060,N_30276);
and U38378 (N_38378,N_33602,N_32096);
nand U38379 (N_38379,N_32745,N_34368);
xor U38380 (N_38380,N_30071,N_33991);
or U38381 (N_38381,N_33100,N_33180);
nor U38382 (N_38382,N_33476,N_32910);
or U38383 (N_38383,N_30123,N_31059);
nand U38384 (N_38384,N_34955,N_34943);
or U38385 (N_38385,N_30924,N_31086);
nor U38386 (N_38386,N_34844,N_30620);
or U38387 (N_38387,N_34100,N_33765);
and U38388 (N_38388,N_31694,N_32973);
nand U38389 (N_38389,N_30263,N_32471);
nor U38390 (N_38390,N_30913,N_31367);
nand U38391 (N_38391,N_31039,N_33832);
and U38392 (N_38392,N_34960,N_32353);
nand U38393 (N_38393,N_30609,N_32811);
or U38394 (N_38394,N_31440,N_31821);
xor U38395 (N_38395,N_34104,N_33951);
nand U38396 (N_38396,N_31742,N_33668);
or U38397 (N_38397,N_33393,N_34833);
nand U38398 (N_38398,N_31997,N_32342);
or U38399 (N_38399,N_32316,N_31951);
nor U38400 (N_38400,N_33230,N_31097);
and U38401 (N_38401,N_33050,N_33836);
or U38402 (N_38402,N_34514,N_34227);
nand U38403 (N_38403,N_32060,N_31645);
nand U38404 (N_38404,N_34287,N_33681);
and U38405 (N_38405,N_33696,N_31520);
xnor U38406 (N_38406,N_34380,N_34126);
xor U38407 (N_38407,N_33070,N_30764);
and U38408 (N_38408,N_31509,N_31542);
or U38409 (N_38409,N_34319,N_31952);
nor U38410 (N_38410,N_33891,N_34980);
nor U38411 (N_38411,N_33092,N_34106);
or U38412 (N_38412,N_33753,N_34826);
xor U38413 (N_38413,N_34485,N_33236);
nor U38414 (N_38414,N_32707,N_32518);
and U38415 (N_38415,N_31081,N_32017);
and U38416 (N_38416,N_33853,N_30116);
nand U38417 (N_38417,N_34853,N_30241);
xnor U38418 (N_38418,N_32719,N_33982);
nor U38419 (N_38419,N_32671,N_30013);
nor U38420 (N_38420,N_32451,N_33102);
nand U38421 (N_38421,N_32719,N_31775);
nand U38422 (N_38422,N_32579,N_32070);
xor U38423 (N_38423,N_33916,N_32230);
xor U38424 (N_38424,N_30170,N_31629);
and U38425 (N_38425,N_33345,N_31823);
or U38426 (N_38426,N_34857,N_31465);
and U38427 (N_38427,N_32428,N_34798);
nor U38428 (N_38428,N_34733,N_30444);
nand U38429 (N_38429,N_30912,N_31182);
or U38430 (N_38430,N_34068,N_34728);
nand U38431 (N_38431,N_33671,N_30994);
nor U38432 (N_38432,N_31215,N_32750);
xor U38433 (N_38433,N_33570,N_33611);
and U38434 (N_38434,N_32555,N_31303);
xor U38435 (N_38435,N_30586,N_32508);
nand U38436 (N_38436,N_30075,N_30990);
nand U38437 (N_38437,N_31374,N_31953);
nand U38438 (N_38438,N_32833,N_32835);
or U38439 (N_38439,N_34909,N_32928);
nand U38440 (N_38440,N_34010,N_33516);
nand U38441 (N_38441,N_32824,N_33166);
xor U38442 (N_38442,N_30136,N_31310);
nand U38443 (N_38443,N_33984,N_33432);
nand U38444 (N_38444,N_33194,N_32994);
xnor U38445 (N_38445,N_31737,N_34217);
xor U38446 (N_38446,N_34393,N_34505);
nand U38447 (N_38447,N_30202,N_33308);
or U38448 (N_38448,N_32240,N_32523);
nand U38449 (N_38449,N_33685,N_34699);
nand U38450 (N_38450,N_34037,N_32488);
or U38451 (N_38451,N_30128,N_33489);
or U38452 (N_38452,N_32151,N_34496);
nand U38453 (N_38453,N_30907,N_30365);
and U38454 (N_38454,N_30375,N_31458);
or U38455 (N_38455,N_33094,N_34900);
nand U38456 (N_38456,N_33256,N_32633);
or U38457 (N_38457,N_30397,N_32445);
nand U38458 (N_38458,N_34956,N_31027);
xor U38459 (N_38459,N_33797,N_33913);
nor U38460 (N_38460,N_31474,N_30677);
and U38461 (N_38461,N_32008,N_32916);
nor U38462 (N_38462,N_32523,N_33595);
or U38463 (N_38463,N_33693,N_34344);
nand U38464 (N_38464,N_31193,N_34579);
and U38465 (N_38465,N_33768,N_31184);
nor U38466 (N_38466,N_33276,N_31689);
nor U38467 (N_38467,N_32780,N_31525);
nor U38468 (N_38468,N_31337,N_32095);
or U38469 (N_38469,N_32673,N_34287);
nor U38470 (N_38470,N_32362,N_32008);
nor U38471 (N_38471,N_33190,N_34732);
and U38472 (N_38472,N_31881,N_34241);
and U38473 (N_38473,N_34450,N_32163);
nand U38474 (N_38474,N_32715,N_32004);
and U38475 (N_38475,N_31698,N_34723);
or U38476 (N_38476,N_30480,N_33226);
and U38477 (N_38477,N_30394,N_31238);
xnor U38478 (N_38478,N_31179,N_33489);
nand U38479 (N_38479,N_32377,N_30782);
nor U38480 (N_38480,N_33125,N_30902);
or U38481 (N_38481,N_34858,N_33343);
or U38482 (N_38482,N_30239,N_34261);
xor U38483 (N_38483,N_33039,N_30990);
nor U38484 (N_38484,N_34968,N_30438);
nor U38485 (N_38485,N_34245,N_31336);
or U38486 (N_38486,N_31766,N_30985);
or U38487 (N_38487,N_34810,N_30072);
nor U38488 (N_38488,N_31614,N_31401);
and U38489 (N_38489,N_31455,N_31199);
nand U38490 (N_38490,N_31143,N_30177);
xor U38491 (N_38491,N_30469,N_32429);
and U38492 (N_38492,N_33153,N_31827);
or U38493 (N_38493,N_30201,N_30696);
nand U38494 (N_38494,N_32035,N_33263);
xor U38495 (N_38495,N_31962,N_31536);
xnor U38496 (N_38496,N_34967,N_32187);
nand U38497 (N_38497,N_31109,N_34650);
nor U38498 (N_38498,N_30176,N_32940);
xor U38499 (N_38499,N_31293,N_30254);
nor U38500 (N_38500,N_30201,N_32550);
xor U38501 (N_38501,N_33365,N_32787);
nand U38502 (N_38502,N_31967,N_31672);
nor U38503 (N_38503,N_31834,N_33301);
or U38504 (N_38504,N_32762,N_31402);
xor U38505 (N_38505,N_31309,N_32712);
nor U38506 (N_38506,N_30957,N_32996);
xor U38507 (N_38507,N_34820,N_31333);
xnor U38508 (N_38508,N_32327,N_32040);
xor U38509 (N_38509,N_32902,N_34172);
and U38510 (N_38510,N_34096,N_33267);
or U38511 (N_38511,N_32375,N_32453);
and U38512 (N_38512,N_30554,N_33910);
or U38513 (N_38513,N_31372,N_30394);
and U38514 (N_38514,N_32577,N_30129);
xnor U38515 (N_38515,N_32669,N_34562);
or U38516 (N_38516,N_31027,N_34760);
xor U38517 (N_38517,N_34380,N_34895);
nand U38518 (N_38518,N_33271,N_32467);
nor U38519 (N_38519,N_34285,N_30885);
or U38520 (N_38520,N_30632,N_34835);
nand U38521 (N_38521,N_34605,N_32579);
or U38522 (N_38522,N_34416,N_32948);
or U38523 (N_38523,N_32980,N_33608);
or U38524 (N_38524,N_30873,N_33326);
nor U38525 (N_38525,N_33544,N_34917);
and U38526 (N_38526,N_34111,N_31978);
nor U38527 (N_38527,N_33732,N_30220);
xor U38528 (N_38528,N_31494,N_32539);
nor U38529 (N_38529,N_34422,N_30066);
and U38530 (N_38530,N_33514,N_30848);
or U38531 (N_38531,N_33936,N_34538);
xor U38532 (N_38532,N_34360,N_30597);
xor U38533 (N_38533,N_34067,N_34740);
xnor U38534 (N_38534,N_31219,N_30269);
or U38535 (N_38535,N_31968,N_31910);
nand U38536 (N_38536,N_34027,N_30618);
nor U38537 (N_38537,N_32365,N_34847);
xor U38538 (N_38538,N_33796,N_32891);
and U38539 (N_38539,N_32056,N_31510);
nand U38540 (N_38540,N_30173,N_31960);
nor U38541 (N_38541,N_33971,N_33454);
nor U38542 (N_38542,N_30213,N_30894);
nand U38543 (N_38543,N_34019,N_30231);
xnor U38544 (N_38544,N_33227,N_31288);
or U38545 (N_38545,N_33873,N_31965);
and U38546 (N_38546,N_32680,N_32223);
and U38547 (N_38547,N_32048,N_32199);
nor U38548 (N_38548,N_34682,N_34354);
and U38549 (N_38549,N_32888,N_33252);
nor U38550 (N_38550,N_34042,N_33962);
xnor U38551 (N_38551,N_33554,N_32271);
or U38552 (N_38552,N_32486,N_33965);
and U38553 (N_38553,N_34673,N_31598);
or U38554 (N_38554,N_33210,N_34739);
nor U38555 (N_38555,N_33406,N_30762);
nor U38556 (N_38556,N_34456,N_31947);
xnor U38557 (N_38557,N_34791,N_32892);
and U38558 (N_38558,N_30108,N_30995);
and U38559 (N_38559,N_30278,N_30479);
or U38560 (N_38560,N_33344,N_34278);
and U38561 (N_38561,N_34294,N_34590);
and U38562 (N_38562,N_34569,N_31157);
and U38563 (N_38563,N_34201,N_30176);
and U38564 (N_38564,N_31761,N_32637);
and U38565 (N_38565,N_30883,N_30583);
nand U38566 (N_38566,N_32643,N_33308);
nand U38567 (N_38567,N_34939,N_30732);
xor U38568 (N_38568,N_32361,N_34317);
xor U38569 (N_38569,N_33288,N_31598);
nor U38570 (N_38570,N_31075,N_31448);
nand U38571 (N_38571,N_31956,N_30390);
and U38572 (N_38572,N_34533,N_30170);
and U38573 (N_38573,N_31044,N_34492);
nand U38574 (N_38574,N_33087,N_30198);
and U38575 (N_38575,N_32720,N_33331);
nand U38576 (N_38576,N_32589,N_34438);
xnor U38577 (N_38577,N_32039,N_33315);
nor U38578 (N_38578,N_31281,N_32892);
nor U38579 (N_38579,N_33471,N_34790);
and U38580 (N_38580,N_33039,N_30168);
nor U38581 (N_38581,N_31212,N_34145);
xnor U38582 (N_38582,N_34397,N_33900);
nand U38583 (N_38583,N_34146,N_34131);
or U38584 (N_38584,N_34780,N_32720);
nor U38585 (N_38585,N_34563,N_34281);
or U38586 (N_38586,N_32912,N_31337);
xor U38587 (N_38587,N_33296,N_33028);
xnor U38588 (N_38588,N_31597,N_33464);
and U38589 (N_38589,N_32237,N_34573);
nor U38590 (N_38590,N_33327,N_32078);
and U38591 (N_38591,N_31428,N_34470);
or U38592 (N_38592,N_34225,N_30411);
xnor U38593 (N_38593,N_33705,N_32552);
and U38594 (N_38594,N_32067,N_33232);
nor U38595 (N_38595,N_30963,N_31988);
and U38596 (N_38596,N_32963,N_32926);
nand U38597 (N_38597,N_33432,N_34769);
or U38598 (N_38598,N_31289,N_31804);
and U38599 (N_38599,N_32539,N_33624);
or U38600 (N_38600,N_30207,N_32094);
nor U38601 (N_38601,N_33806,N_33012);
nor U38602 (N_38602,N_30754,N_32997);
or U38603 (N_38603,N_34567,N_34524);
or U38604 (N_38604,N_32306,N_34697);
xnor U38605 (N_38605,N_32074,N_32356);
xor U38606 (N_38606,N_32626,N_31427);
and U38607 (N_38607,N_31871,N_32647);
xnor U38608 (N_38608,N_34544,N_34947);
or U38609 (N_38609,N_31887,N_32349);
nor U38610 (N_38610,N_30709,N_32767);
xor U38611 (N_38611,N_32424,N_32196);
and U38612 (N_38612,N_31699,N_33856);
nand U38613 (N_38613,N_30459,N_34673);
nor U38614 (N_38614,N_32808,N_32974);
xor U38615 (N_38615,N_33522,N_33238);
or U38616 (N_38616,N_31643,N_30302);
and U38617 (N_38617,N_33079,N_32870);
and U38618 (N_38618,N_32266,N_31702);
or U38619 (N_38619,N_34525,N_34368);
nor U38620 (N_38620,N_34554,N_31143);
nor U38621 (N_38621,N_32095,N_31528);
or U38622 (N_38622,N_34738,N_33376);
or U38623 (N_38623,N_33456,N_33701);
xor U38624 (N_38624,N_34717,N_31288);
nor U38625 (N_38625,N_34287,N_32271);
nand U38626 (N_38626,N_34355,N_33178);
and U38627 (N_38627,N_33749,N_32808);
nand U38628 (N_38628,N_31921,N_33408);
nor U38629 (N_38629,N_34993,N_32252);
or U38630 (N_38630,N_34550,N_33793);
nor U38631 (N_38631,N_30859,N_34779);
nor U38632 (N_38632,N_33525,N_34094);
nor U38633 (N_38633,N_33516,N_30895);
nor U38634 (N_38634,N_31348,N_30298);
nor U38635 (N_38635,N_32873,N_30617);
xnor U38636 (N_38636,N_34775,N_33551);
or U38637 (N_38637,N_34639,N_31162);
nor U38638 (N_38638,N_33602,N_30465);
xnor U38639 (N_38639,N_32618,N_32720);
nand U38640 (N_38640,N_31191,N_30684);
or U38641 (N_38641,N_31597,N_30370);
nor U38642 (N_38642,N_30690,N_30264);
or U38643 (N_38643,N_31451,N_31077);
and U38644 (N_38644,N_31612,N_31364);
nand U38645 (N_38645,N_32059,N_31710);
and U38646 (N_38646,N_33599,N_30543);
and U38647 (N_38647,N_33631,N_33869);
and U38648 (N_38648,N_32199,N_32703);
xnor U38649 (N_38649,N_30475,N_33937);
nor U38650 (N_38650,N_32480,N_30526);
and U38651 (N_38651,N_31271,N_31581);
xnor U38652 (N_38652,N_31282,N_34391);
xor U38653 (N_38653,N_32917,N_34793);
or U38654 (N_38654,N_34433,N_31571);
nand U38655 (N_38655,N_34127,N_34315);
xnor U38656 (N_38656,N_30021,N_34084);
and U38657 (N_38657,N_32628,N_32352);
and U38658 (N_38658,N_32964,N_31134);
nand U38659 (N_38659,N_32289,N_31265);
xnor U38660 (N_38660,N_30232,N_30260);
or U38661 (N_38661,N_34568,N_33292);
nor U38662 (N_38662,N_32744,N_34642);
nor U38663 (N_38663,N_33660,N_34915);
or U38664 (N_38664,N_33782,N_32943);
or U38665 (N_38665,N_33194,N_34633);
xnor U38666 (N_38666,N_31037,N_30138);
nand U38667 (N_38667,N_30016,N_31266);
and U38668 (N_38668,N_33733,N_33832);
xor U38669 (N_38669,N_30011,N_33819);
nor U38670 (N_38670,N_30560,N_33226);
nand U38671 (N_38671,N_31090,N_30218);
or U38672 (N_38672,N_31866,N_34072);
or U38673 (N_38673,N_31785,N_30922);
nand U38674 (N_38674,N_33281,N_30205);
and U38675 (N_38675,N_33531,N_33485);
xor U38676 (N_38676,N_30604,N_31443);
and U38677 (N_38677,N_30819,N_31663);
and U38678 (N_38678,N_31843,N_34488);
nor U38679 (N_38679,N_34891,N_31339);
or U38680 (N_38680,N_30544,N_32036);
and U38681 (N_38681,N_31635,N_32475);
xor U38682 (N_38682,N_31146,N_34768);
xnor U38683 (N_38683,N_34917,N_30715);
and U38684 (N_38684,N_31981,N_33514);
nand U38685 (N_38685,N_34374,N_33125);
xnor U38686 (N_38686,N_30198,N_32101);
nor U38687 (N_38687,N_34828,N_33291);
nor U38688 (N_38688,N_33769,N_30695);
or U38689 (N_38689,N_33277,N_30487);
xnor U38690 (N_38690,N_31444,N_32435);
nand U38691 (N_38691,N_33849,N_30672);
nor U38692 (N_38692,N_33662,N_32243);
nand U38693 (N_38693,N_31804,N_30707);
and U38694 (N_38694,N_31944,N_32213);
nand U38695 (N_38695,N_33789,N_33408);
or U38696 (N_38696,N_34815,N_34427);
or U38697 (N_38697,N_32688,N_34983);
xnor U38698 (N_38698,N_33901,N_33249);
nor U38699 (N_38699,N_32460,N_33595);
nand U38700 (N_38700,N_31843,N_34898);
xor U38701 (N_38701,N_34340,N_30921);
or U38702 (N_38702,N_31840,N_33932);
and U38703 (N_38703,N_31640,N_30022);
nand U38704 (N_38704,N_30525,N_31295);
xnor U38705 (N_38705,N_31607,N_31471);
nand U38706 (N_38706,N_32991,N_30713);
or U38707 (N_38707,N_30753,N_33021);
xor U38708 (N_38708,N_30149,N_31218);
or U38709 (N_38709,N_32239,N_34822);
and U38710 (N_38710,N_30315,N_33495);
xor U38711 (N_38711,N_32725,N_30468);
and U38712 (N_38712,N_30637,N_31459);
and U38713 (N_38713,N_31145,N_34180);
and U38714 (N_38714,N_31587,N_33857);
xnor U38715 (N_38715,N_32657,N_34524);
or U38716 (N_38716,N_33260,N_32948);
nand U38717 (N_38717,N_30940,N_34887);
or U38718 (N_38718,N_31052,N_34374);
or U38719 (N_38719,N_33191,N_30166);
nor U38720 (N_38720,N_31387,N_32846);
nor U38721 (N_38721,N_34795,N_31918);
nand U38722 (N_38722,N_34624,N_34716);
nor U38723 (N_38723,N_30124,N_34328);
nor U38724 (N_38724,N_30566,N_33431);
and U38725 (N_38725,N_33923,N_34557);
or U38726 (N_38726,N_30409,N_30756);
xnor U38727 (N_38727,N_32765,N_34699);
or U38728 (N_38728,N_30008,N_33981);
and U38729 (N_38729,N_32939,N_33174);
or U38730 (N_38730,N_34010,N_32735);
nand U38731 (N_38731,N_30333,N_31293);
or U38732 (N_38732,N_32777,N_31317);
and U38733 (N_38733,N_32902,N_31686);
or U38734 (N_38734,N_31817,N_32382);
and U38735 (N_38735,N_33575,N_32815);
nand U38736 (N_38736,N_30642,N_34848);
nand U38737 (N_38737,N_30770,N_30971);
xnor U38738 (N_38738,N_32745,N_30023);
nand U38739 (N_38739,N_31349,N_30706);
xor U38740 (N_38740,N_30874,N_34120);
nor U38741 (N_38741,N_30260,N_33157);
and U38742 (N_38742,N_33039,N_32497);
and U38743 (N_38743,N_31962,N_30018);
or U38744 (N_38744,N_31927,N_31321);
xnor U38745 (N_38745,N_33028,N_32452);
or U38746 (N_38746,N_31011,N_33106);
nor U38747 (N_38747,N_33617,N_30462);
xnor U38748 (N_38748,N_30580,N_33716);
and U38749 (N_38749,N_30215,N_33857);
nand U38750 (N_38750,N_32408,N_30083);
xnor U38751 (N_38751,N_33025,N_30559);
nand U38752 (N_38752,N_30475,N_32917);
or U38753 (N_38753,N_33407,N_34570);
nor U38754 (N_38754,N_34402,N_31079);
nand U38755 (N_38755,N_34795,N_30427);
nand U38756 (N_38756,N_34051,N_32313);
nor U38757 (N_38757,N_30935,N_30687);
nand U38758 (N_38758,N_30649,N_30601);
nand U38759 (N_38759,N_32512,N_31225);
nor U38760 (N_38760,N_32952,N_32215);
or U38761 (N_38761,N_34494,N_30113);
or U38762 (N_38762,N_30454,N_34836);
xnor U38763 (N_38763,N_30341,N_30019);
xor U38764 (N_38764,N_30689,N_32453);
nor U38765 (N_38765,N_31345,N_34746);
nand U38766 (N_38766,N_32998,N_34499);
nor U38767 (N_38767,N_33713,N_33386);
and U38768 (N_38768,N_32323,N_31751);
and U38769 (N_38769,N_34285,N_31934);
xnor U38770 (N_38770,N_34663,N_34801);
nand U38771 (N_38771,N_30007,N_33732);
nor U38772 (N_38772,N_30763,N_31774);
nor U38773 (N_38773,N_31033,N_34368);
nor U38774 (N_38774,N_31621,N_30895);
xnor U38775 (N_38775,N_33476,N_32457);
or U38776 (N_38776,N_34073,N_30225);
nor U38777 (N_38777,N_33528,N_30952);
or U38778 (N_38778,N_32471,N_30400);
nand U38779 (N_38779,N_31759,N_32950);
or U38780 (N_38780,N_31691,N_30591);
and U38781 (N_38781,N_32122,N_33865);
and U38782 (N_38782,N_30214,N_31338);
and U38783 (N_38783,N_30927,N_32304);
and U38784 (N_38784,N_32233,N_32426);
and U38785 (N_38785,N_32854,N_34638);
and U38786 (N_38786,N_34920,N_30079);
nor U38787 (N_38787,N_32333,N_33647);
or U38788 (N_38788,N_31279,N_32886);
nor U38789 (N_38789,N_32167,N_31167);
xnor U38790 (N_38790,N_31648,N_33531);
nor U38791 (N_38791,N_32439,N_33476);
nand U38792 (N_38792,N_33793,N_33047);
xnor U38793 (N_38793,N_31760,N_31737);
nand U38794 (N_38794,N_32643,N_34116);
nor U38795 (N_38795,N_30911,N_33119);
or U38796 (N_38796,N_31403,N_30072);
or U38797 (N_38797,N_30513,N_30475);
nor U38798 (N_38798,N_34097,N_33326);
or U38799 (N_38799,N_32680,N_31150);
xnor U38800 (N_38800,N_34059,N_34241);
and U38801 (N_38801,N_34141,N_32177);
or U38802 (N_38802,N_31750,N_30062);
nand U38803 (N_38803,N_34295,N_30491);
xor U38804 (N_38804,N_34976,N_30596);
and U38805 (N_38805,N_33996,N_34581);
nor U38806 (N_38806,N_32188,N_31461);
xor U38807 (N_38807,N_34573,N_31556);
xnor U38808 (N_38808,N_34640,N_30982);
nor U38809 (N_38809,N_31857,N_33063);
nand U38810 (N_38810,N_31712,N_32001);
and U38811 (N_38811,N_33123,N_32398);
or U38812 (N_38812,N_33808,N_33689);
nand U38813 (N_38813,N_33351,N_30974);
nand U38814 (N_38814,N_33488,N_32231);
or U38815 (N_38815,N_34913,N_32692);
or U38816 (N_38816,N_34510,N_33291);
nor U38817 (N_38817,N_33356,N_31554);
nor U38818 (N_38818,N_33987,N_30557);
or U38819 (N_38819,N_33714,N_30708);
nor U38820 (N_38820,N_32838,N_32140);
or U38821 (N_38821,N_30682,N_32193);
xnor U38822 (N_38822,N_30184,N_34383);
xor U38823 (N_38823,N_33810,N_34350);
nand U38824 (N_38824,N_30487,N_31233);
nand U38825 (N_38825,N_33631,N_33029);
nand U38826 (N_38826,N_33951,N_31322);
and U38827 (N_38827,N_31131,N_32763);
or U38828 (N_38828,N_30127,N_32206);
or U38829 (N_38829,N_34224,N_32619);
nor U38830 (N_38830,N_33765,N_33050);
nand U38831 (N_38831,N_30472,N_30095);
and U38832 (N_38832,N_31806,N_31726);
or U38833 (N_38833,N_31834,N_34501);
nand U38834 (N_38834,N_33857,N_32758);
nand U38835 (N_38835,N_32960,N_31095);
nand U38836 (N_38836,N_33424,N_34556);
or U38837 (N_38837,N_30624,N_30951);
or U38838 (N_38838,N_33842,N_33099);
or U38839 (N_38839,N_32445,N_34272);
nand U38840 (N_38840,N_34646,N_32034);
or U38841 (N_38841,N_33003,N_34350);
or U38842 (N_38842,N_31295,N_31681);
or U38843 (N_38843,N_31611,N_32847);
or U38844 (N_38844,N_33294,N_30481);
and U38845 (N_38845,N_32561,N_33551);
or U38846 (N_38846,N_30392,N_33182);
or U38847 (N_38847,N_32719,N_32403);
nor U38848 (N_38848,N_34238,N_34959);
xnor U38849 (N_38849,N_33524,N_33600);
and U38850 (N_38850,N_30723,N_34616);
xor U38851 (N_38851,N_33016,N_30301);
nand U38852 (N_38852,N_32026,N_33369);
xor U38853 (N_38853,N_32446,N_32478);
xor U38854 (N_38854,N_32772,N_32864);
or U38855 (N_38855,N_34318,N_31281);
xor U38856 (N_38856,N_30894,N_32148);
xor U38857 (N_38857,N_30876,N_31228);
or U38858 (N_38858,N_30169,N_34820);
xor U38859 (N_38859,N_30242,N_31839);
nand U38860 (N_38860,N_31822,N_34291);
nand U38861 (N_38861,N_34317,N_30756);
nand U38862 (N_38862,N_31044,N_33734);
xor U38863 (N_38863,N_32548,N_34437);
and U38864 (N_38864,N_30895,N_34589);
nor U38865 (N_38865,N_31058,N_34668);
xor U38866 (N_38866,N_31582,N_32378);
xor U38867 (N_38867,N_30655,N_31053);
or U38868 (N_38868,N_31918,N_30524);
nand U38869 (N_38869,N_32021,N_33118);
nor U38870 (N_38870,N_32086,N_34757);
nand U38871 (N_38871,N_30203,N_32178);
or U38872 (N_38872,N_31174,N_31296);
xnor U38873 (N_38873,N_30668,N_33338);
nand U38874 (N_38874,N_33854,N_33823);
nor U38875 (N_38875,N_30454,N_32179);
and U38876 (N_38876,N_32452,N_31173);
and U38877 (N_38877,N_33757,N_31301);
nand U38878 (N_38878,N_33461,N_34193);
nand U38879 (N_38879,N_34936,N_34574);
or U38880 (N_38880,N_34708,N_34300);
nor U38881 (N_38881,N_30008,N_33097);
or U38882 (N_38882,N_31895,N_31139);
nand U38883 (N_38883,N_31549,N_32487);
xor U38884 (N_38884,N_32151,N_34908);
and U38885 (N_38885,N_33662,N_33224);
or U38886 (N_38886,N_31040,N_34773);
nor U38887 (N_38887,N_30499,N_30103);
or U38888 (N_38888,N_30923,N_32528);
and U38889 (N_38889,N_30020,N_32805);
and U38890 (N_38890,N_31560,N_31637);
and U38891 (N_38891,N_34315,N_32018);
or U38892 (N_38892,N_34764,N_33333);
xnor U38893 (N_38893,N_30906,N_31451);
and U38894 (N_38894,N_30928,N_33035);
xor U38895 (N_38895,N_31540,N_33620);
xor U38896 (N_38896,N_34997,N_31079);
and U38897 (N_38897,N_31834,N_30194);
nand U38898 (N_38898,N_31570,N_31696);
and U38899 (N_38899,N_31162,N_32826);
nor U38900 (N_38900,N_31746,N_32293);
xor U38901 (N_38901,N_33705,N_31564);
nor U38902 (N_38902,N_30543,N_32472);
or U38903 (N_38903,N_33460,N_33412);
nand U38904 (N_38904,N_32238,N_31917);
or U38905 (N_38905,N_32610,N_32503);
and U38906 (N_38906,N_30877,N_31416);
nand U38907 (N_38907,N_33166,N_30011);
and U38908 (N_38908,N_32554,N_30918);
nand U38909 (N_38909,N_31168,N_30686);
or U38910 (N_38910,N_30271,N_31940);
or U38911 (N_38911,N_33227,N_33845);
or U38912 (N_38912,N_30940,N_33567);
or U38913 (N_38913,N_32536,N_30707);
and U38914 (N_38914,N_33895,N_31361);
and U38915 (N_38915,N_32219,N_32913);
and U38916 (N_38916,N_31453,N_33901);
nor U38917 (N_38917,N_34357,N_34009);
and U38918 (N_38918,N_30179,N_34119);
xnor U38919 (N_38919,N_34237,N_31555);
xnor U38920 (N_38920,N_34762,N_33276);
or U38921 (N_38921,N_34048,N_31538);
and U38922 (N_38922,N_30041,N_31548);
nand U38923 (N_38923,N_30586,N_31598);
or U38924 (N_38924,N_30472,N_32090);
and U38925 (N_38925,N_31641,N_32545);
nand U38926 (N_38926,N_30620,N_31137);
nand U38927 (N_38927,N_33713,N_31381);
and U38928 (N_38928,N_33248,N_33988);
nor U38929 (N_38929,N_34926,N_33415);
nand U38930 (N_38930,N_30096,N_33362);
nand U38931 (N_38931,N_34468,N_31833);
nor U38932 (N_38932,N_32026,N_32081);
or U38933 (N_38933,N_30994,N_30157);
or U38934 (N_38934,N_30099,N_30328);
nand U38935 (N_38935,N_32375,N_33222);
nand U38936 (N_38936,N_33891,N_32904);
xnor U38937 (N_38937,N_33105,N_30458);
and U38938 (N_38938,N_34543,N_32997);
nor U38939 (N_38939,N_34057,N_32740);
xor U38940 (N_38940,N_31997,N_32273);
and U38941 (N_38941,N_33865,N_30156);
nor U38942 (N_38942,N_31792,N_34367);
and U38943 (N_38943,N_33178,N_30987);
and U38944 (N_38944,N_34466,N_34989);
nor U38945 (N_38945,N_34815,N_30881);
nor U38946 (N_38946,N_30995,N_32722);
nand U38947 (N_38947,N_34351,N_33680);
nand U38948 (N_38948,N_32933,N_34243);
and U38949 (N_38949,N_30136,N_31945);
and U38950 (N_38950,N_34869,N_34577);
xnor U38951 (N_38951,N_33161,N_30169);
xnor U38952 (N_38952,N_34118,N_34645);
nor U38953 (N_38953,N_34113,N_34620);
or U38954 (N_38954,N_30677,N_30782);
and U38955 (N_38955,N_31324,N_33103);
and U38956 (N_38956,N_33911,N_34925);
or U38957 (N_38957,N_34458,N_34589);
nor U38958 (N_38958,N_34188,N_31701);
and U38959 (N_38959,N_33803,N_33474);
and U38960 (N_38960,N_32341,N_32529);
nor U38961 (N_38961,N_31700,N_34385);
and U38962 (N_38962,N_32194,N_32277);
or U38963 (N_38963,N_31798,N_33855);
nand U38964 (N_38964,N_30651,N_31913);
nand U38965 (N_38965,N_31520,N_30798);
nor U38966 (N_38966,N_31555,N_30448);
and U38967 (N_38967,N_30915,N_31489);
nor U38968 (N_38968,N_32091,N_34202);
nand U38969 (N_38969,N_30236,N_34468);
xnor U38970 (N_38970,N_32709,N_30334);
nor U38971 (N_38971,N_34198,N_34292);
nand U38972 (N_38972,N_32124,N_31303);
xor U38973 (N_38973,N_31535,N_34623);
nor U38974 (N_38974,N_30006,N_31466);
or U38975 (N_38975,N_31479,N_34708);
or U38976 (N_38976,N_32753,N_33398);
nor U38977 (N_38977,N_33860,N_34732);
nand U38978 (N_38978,N_31801,N_33846);
and U38979 (N_38979,N_31136,N_32003);
and U38980 (N_38980,N_34791,N_33533);
xnor U38981 (N_38981,N_33873,N_34076);
and U38982 (N_38982,N_31234,N_33790);
xor U38983 (N_38983,N_33127,N_30466);
xor U38984 (N_38984,N_33362,N_30446);
nor U38985 (N_38985,N_32758,N_34170);
xor U38986 (N_38986,N_32459,N_33777);
and U38987 (N_38987,N_31757,N_31789);
xnor U38988 (N_38988,N_34358,N_30375);
nor U38989 (N_38989,N_34699,N_34872);
nor U38990 (N_38990,N_30240,N_32655);
nor U38991 (N_38991,N_31958,N_31910);
nor U38992 (N_38992,N_31241,N_33115);
nand U38993 (N_38993,N_31635,N_31287);
nor U38994 (N_38994,N_33421,N_30828);
and U38995 (N_38995,N_30791,N_31473);
and U38996 (N_38996,N_34393,N_32559);
and U38997 (N_38997,N_33232,N_31718);
and U38998 (N_38998,N_33201,N_32413);
nand U38999 (N_38999,N_32452,N_33874);
xor U39000 (N_39000,N_34460,N_32613);
nand U39001 (N_39001,N_33374,N_34210);
and U39002 (N_39002,N_33806,N_34166);
and U39003 (N_39003,N_34286,N_34465);
xor U39004 (N_39004,N_32397,N_34456);
xor U39005 (N_39005,N_34637,N_32015);
nand U39006 (N_39006,N_33489,N_33859);
xnor U39007 (N_39007,N_33467,N_33324);
nand U39008 (N_39008,N_30667,N_33223);
nand U39009 (N_39009,N_32583,N_34124);
xor U39010 (N_39010,N_34418,N_33697);
nand U39011 (N_39011,N_34805,N_32019);
and U39012 (N_39012,N_34387,N_34172);
and U39013 (N_39013,N_30952,N_33650);
xnor U39014 (N_39014,N_34133,N_31561);
or U39015 (N_39015,N_34838,N_30527);
or U39016 (N_39016,N_32430,N_34414);
and U39017 (N_39017,N_30821,N_31165);
and U39018 (N_39018,N_34546,N_30001);
nand U39019 (N_39019,N_31222,N_34992);
and U39020 (N_39020,N_32024,N_32101);
xnor U39021 (N_39021,N_32389,N_33102);
or U39022 (N_39022,N_32895,N_30370);
or U39023 (N_39023,N_31862,N_32937);
xor U39024 (N_39024,N_30384,N_31149);
nor U39025 (N_39025,N_34346,N_34875);
nor U39026 (N_39026,N_30691,N_33783);
or U39027 (N_39027,N_33285,N_30429);
nor U39028 (N_39028,N_31391,N_31033);
and U39029 (N_39029,N_34356,N_31508);
nand U39030 (N_39030,N_31483,N_32008);
and U39031 (N_39031,N_31696,N_31106);
and U39032 (N_39032,N_31555,N_33770);
and U39033 (N_39033,N_31040,N_33698);
nand U39034 (N_39034,N_32953,N_30606);
or U39035 (N_39035,N_31630,N_31182);
nor U39036 (N_39036,N_31382,N_34532);
xnor U39037 (N_39037,N_31920,N_30995);
or U39038 (N_39038,N_31867,N_30657);
nor U39039 (N_39039,N_30190,N_34029);
nor U39040 (N_39040,N_34767,N_31778);
nor U39041 (N_39041,N_33114,N_32866);
xnor U39042 (N_39042,N_32583,N_31097);
or U39043 (N_39043,N_33505,N_30152);
or U39044 (N_39044,N_33375,N_32101);
and U39045 (N_39045,N_34896,N_30722);
nor U39046 (N_39046,N_30812,N_32800);
nand U39047 (N_39047,N_33925,N_34714);
nor U39048 (N_39048,N_32779,N_31458);
nand U39049 (N_39049,N_31299,N_30998);
nor U39050 (N_39050,N_34429,N_34353);
xor U39051 (N_39051,N_30017,N_32921);
nand U39052 (N_39052,N_31496,N_32411);
or U39053 (N_39053,N_34997,N_34877);
nand U39054 (N_39054,N_34084,N_31620);
nand U39055 (N_39055,N_30004,N_30654);
xor U39056 (N_39056,N_34754,N_34156);
and U39057 (N_39057,N_30957,N_30058);
xor U39058 (N_39058,N_30440,N_30539);
xnor U39059 (N_39059,N_34249,N_32749);
nand U39060 (N_39060,N_30817,N_32567);
nand U39061 (N_39061,N_30848,N_31725);
nor U39062 (N_39062,N_31002,N_34288);
or U39063 (N_39063,N_31819,N_30399);
nand U39064 (N_39064,N_34839,N_30991);
xor U39065 (N_39065,N_30217,N_30765);
and U39066 (N_39066,N_33650,N_34339);
or U39067 (N_39067,N_33870,N_32582);
nor U39068 (N_39068,N_30571,N_31826);
or U39069 (N_39069,N_30078,N_32733);
or U39070 (N_39070,N_34022,N_32985);
xnor U39071 (N_39071,N_32282,N_30075);
xor U39072 (N_39072,N_33242,N_31207);
nor U39073 (N_39073,N_34227,N_34352);
xnor U39074 (N_39074,N_31143,N_33544);
xnor U39075 (N_39075,N_31341,N_34833);
nand U39076 (N_39076,N_33809,N_31859);
nand U39077 (N_39077,N_34508,N_31664);
or U39078 (N_39078,N_33525,N_34760);
and U39079 (N_39079,N_34850,N_31692);
xnor U39080 (N_39080,N_33965,N_30333);
xor U39081 (N_39081,N_33495,N_31758);
nand U39082 (N_39082,N_32275,N_31895);
and U39083 (N_39083,N_34868,N_33785);
xor U39084 (N_39084,N_32934,N_30942);
or U39085 (N_39085,N_31617,N_32700);
and U39086 (N_39086,N_30865,N_34718);
or U39087 (N_39087,N_31226,N_30445);
nor U39088 (N_39088,N_34884,N_34067);
xor U39089 (N_39089,N_33915,N_32870);
xnor U39090 (N_39090,N_30688,N_32077);
and U39091 (N_39091,N_34833,N_34604);
and U39092 (N_39092,N_30687,N_32992);
nand U39093 (N_39093,N_30496,N_30775);
nand U39094 (N_39094,N_32985,N_30324);
and U39095 (N_39095,N_32812,N_32996);
nor U39096 (N_39096,N_30184,N_30954);
or U39097 (N_39097,N_34631,N_32746);
xnor U39098 (N_39098,N_33594,N_31718);
nand U39099 (N_39099,N_34737,N_34847);
xor U39100 (N_39100,N_31823,N_31955);
nor U39101 (N_39101,N_34223,N_32191);
xnor U39102 (N_39102,N_31871,N_34350);
and U39103 (N_39103,N_31475,N_30731);
or U39104 (N_39104,N_32375,N_34690);
nor U39105 (N_39105,N_30956,N_34157);
xnor U39106 (N_39106,N_32567,N_32171);
or U39107 (N_39107,N_33247,N_31209);
nand U39108 (N_39108,N_31448,N_32001);
or U39109 (N_39109,N_30635,N_34561);
xor U39110 (N_39110,N_30623,N_31296);
or U39111 (N_39111,N_34382,N_32447);
nand U39112 (N_39112,N_32706,N_30427);
or U39113 (N_39113,N_34228,N_32055);
and U39114 (N_39114,N_33751,N_33716);
or U39115 (N_39115,N_34541,N_30070);
nand U39116 (N_39116,N_34374,N_33860);
or U39117 (N_39117,N_32688,N_30338);
nand U39118 (N_39118,N_31630,N_34605);
xor U39119 (N_39119,N_32764,N_31848);
nor U39120 (N_39120,N_32155,N_30356);
xor U39121 (N_39121,N_33213,N_32482);
and U39122 (N_39122,N_31426,N_34266);
nor U39123 (N_39123,N_32501,N_30075);
nor U39124 (N_39124,N_31964,N_30916);
or U39125 (N_39125,N_32314,N_34427);
or U39126 (N_39126,N_34579,N_32918);
nand U39127 (N_39127,N_34571,N_31731);
nor U39128 (N_39128,N_31770,N_33048);
nor U39129 (N_39129,N_30429,N_33386);
or U39130 (N_39130,N_32062,N_34685);
nor U39131 (N_39131,N_31752,N_32698);
nor U39132 (N_39132,N_30544,N_33496);
xor U39133 (N_39133,N_30828,N_34168);
nor U39134 (N_39134,N_31536,N_32927);
xnor U39135 (N_39135,N_30592,N_31195);
and U39136 (N_39136,N_32204,N_32053);
xnor U39137 (N_39137,N_30910,N_33781);
xnor U39138 (N_39138,N_32236,N_34786);
nor U39139 (N_39139,N_34010,N_30561);
nand U39140 (N_39140,N_30105,N_33276);
and U39141 (N_39141,N_30400,N_31603);
or U39142 (N_39142,N_31664,N_34420);
and U39143 (N_39143,N_30760,N_32956);
or U39144 (N_39144,N_34661,N_33708);
xor U39145 (N_39145,N_30279,N_33569);
nand U39146 (N_39146,N_30368,N_30085);
nand U39147 (N_39147,N_34639,N_32804);
nand U39148 (N_39148,N_31921,N_33970);
nand U39149 (N_39149,N_33390,N_34519);
nor U39150 (N_39150,N_34647,N_30714);
nor U39151 (N_39151,N_30033,N_34553);
xnor U39152 (N_39152,N_34494,N_30000);
nand U39153 (N_39153,N_30850,N_34680);
or U39154 (N_39154,N_31698,N_30408);
nand U39155 (N_39155,N_34672,N_34491);
or U39156 (N_39156,N_33574,N_32213);
and U39157 (N_39157,N_34652,N_30547);
and U39158 (N_39158,N_32463,N_33019);
nand U39159 (N_39159,N_34794,N_31147);
nand U39160 (N_39160,N_30752,N_32952);
or U39161 (N_39161,N_33384,N_30842);
xor U39162 (N_39162,N_34794,N_32731);
nand U39163 (N_39163,N_30358,N_33140);
xor U39164 (N_39164,N_32807,N_33642);
and U39165 (N_39165,N_34606,N_34555);
or U39166 (N_39166,N_32401,N_33858);
nor U39167 (N_39167,N_33332,N_33293);
or U39168 (N_39168,N_31767,N_31687);
xnor U39169 (N_39169,N_32875,N_34443);
or U39170 (N_39170,N_32939,N_33757);
nand U39171 (N_39171,N_32705,N_31146);
and U39172 (N_39172,N_31160,N_30444);
and U39173 (N_39173,N_32654,N_31118);
or U39174 (N_39174,N_30163,N_31025);
xnor U39175 (N_39175,N_33456,N_34146);
xor U39176 (N_39176,N_30732,N_32317);
nand U39177 (N_39177,N_33613,N_33193);
nand U39178 (N_39178,N_33435,N_34613);
nor U39179 (N_39179,N_34853,N_31956);
nand U39180 (N_39180,N_34805,N_33616);
nor U39181 (N_39181,N_33071,N_30830);
nor U39182 (N_39182,N_32391,N_32940);
nand U39183 (N_39183,N_32715,N_32764);
and U39184 (N_39184,N_33282,N_33973);
nor U39185 (N_39185,N_32078,N_31319);
and U39186 (N_39186,N_34204,N_30727);
nor U39187 (N_39187,N_32257,N_34928);
and U39188 (N_39188,N_32460,N_34774);
nand U39189 (N_39189,N_34814,N_34658);
or U39190 (N_39190,N_32987,N_31880);
nand U39191 (N_39191,N_30013,N_34147);
and U39192 (N_39192,N_30099,N_31134);
nand U39193 (N_39193,N_34655,N_33474);
nor U39194 (N_39194,N_30757,N_30636);
or U39195 (N_39195,N_32054,N_31445);
nor U39196 (N_39196,N_34716,N_34220);
xnor U39197 (N_39197,N_32131,N_30665);
and U39198 (N_39198,N_33300,N_32400);
and U39199 (N_39199,N_33267,N_30277);
nor U39200 (N_39200,N_30789,N_33662);
and U39201 (N_39201,N_30387,N_31924);
nor U39202 (N_39202,N_34628,N_33459);
or U39203 (N_39203,N_34190,N_31403);
nand U39204 (N_39204,N_33774,N_30795);
nand U39205 (N_39205,N_33767,N_30003);
nor U39206 (N_39206,N_31461,N_32793);
xnor U39207 (N_39207,N_32430,N_33018);
and U39208 (N_39208,N_32962,N_33941);
nand U39209 (N_39209,N_33935,N_34517);
nor U39210 (N_39210,N_34661,N_32312);
and U39211 (N_39211,N_34995,N_34086);
nor U39212 (N_39212,N_33934,N_34207);
or U39213 (N_39213,N_32232,N_30985);
or U39214 (N_39214,N_30063,N_30367);
nand U39215 (N_39215,N_34834,N_34068);
nand U39216 (N_39216,N_30209,N_30021);
nand U39217 (N_39217,N_34571,N_30688);
or U39218 (N_39218,N_32370,N_30614);
nand U39219 (N_39219,N_34666,N_34319);
xor U39220 (N_39220,N_31337,N_32711);
nor U39221 (N_39221,N_32436,N_31349);
and U39222 (N_39222,N_32167,N_32609);
and U39223 (N_39223,N_32193,N_31295);
nor U39224 (N_39224,N_32494,N_31009);
nor U39225 (N_39225,N_34447,N_31764);
nand U39226 (N_39226,N_33459,N_30957);
and U39227 (N_39227,N_30050,N_30113);
or U39228 (N_39228,N_33056,N_34129);
or U39229 (N_39229,N_32786,N_33600);
or U39230 (N_39230,N_30512,N_33103);
nor U39231 (N_39231,N_32114,N_34605);
xor U39232 (N_39232,N_31105,N_33728);
or U39233 (N_39233,N_34556,N_33688);
and U39234 (N_39234,N_34562,N_31253);
and U39235 (N_39235,N_34567,N_31947);
nor U39236 (N_39236,N_34167,N_32808);
nand U39237 (N_39237,N_31841,N_32056);
nand U39238 (N_39238,N_34583,N_33499);
and U39239 (N_39239,N_31400,N_34292);
nand U39240 (N_39240,N_34900,N_32320);
nand U39241 (N_39241,N_31592,N_33674);
or U39242 (N_39242,N_32476,N_32386);
xnor U39243 (N_39243,N_32219,N_32302);
nand U39244 (N_39244,N_32939,N_33239);
and U39245 (N_39245,N_34360,N_32101);
nor U39246 (N_39246,N_34898,N_32755);
nor U39247 (N_39247,N_31159,N_34733);
or U39248 (N_39248,N_33070,N_34490);
xor U39249 (N_39249,N_30892,N_30944);
or U39250 (N_39250,N_34573,N_32426);
nand U39251 (N_39251,N_33563,N_31048);
or U39252 (N_39252,N_32980,N_32271);
nor U39253 (N_39253,N_34492,N_32426);
xnor U39254 (N_39254,N_32740,N_30421);
xnor U39255 (N_39255,N_32878,N_30168);
nand U39256 (N_39256,N_31666,N_32189);
and U39257 (N_39257,N_34726,N_31670);
xnor U39258 (N_39258,N_34029,N_31897);
nor U39259 (N_39259,N_33960,N_30136);
or U39260 (N_39260,N_30396,N_32843);
and U39261 (N_39261,N_33725,N_33158);
or U39262 (N_39262,N_34999,N_32294);
nor U39263 (N_39263,N_32239,N_30402);
and U39264 (N_39264,N_31063,N_33500);
xor U39265 (N_39265,N_33071,N_33887);
or U39266 (N_39266,N_31588,N_33876);
or U39267 (N_39267,N_31406,N_30004);
or U39268 (N_39268,N_32988,N_30012);
nor U39269 (N_39269,N_32917,N_31183);
nor U39270 (N_39270,N_31854,N_31852);
nand U39271 (N_39271,N_30154,N_32515);
or U39272 (N_39272,N_34128,N_34134);
and U39273 (N_39273,N_33433,N_32343);
nand U39274 (N_39274,N_34655,N_33701);
or U39275 (N_39275,N_32628,N_32576);
and U39276 (N_39276,N_31593,N_31327);
nor U39277 (N_39277,N_33289,N_31662);
nor U39278 (N_39278,N_30918,N_34238);
xor U39279 (N_39279,N_34965,N_32794);
nor U39280 (N_39280,N_34007,N_31892);
and U39281 (N_39281,N_33608,N_31668);
or U39282 (N_39282,N_33214,N_33168);
or U39283 (N_39283,N_31508,N_32945);
and U39284 (N_39284,N_32741,N_33459);
nor U39285 (N_39285,N_30145,N_34346);
nand U39286 (N_39286,N_33621,N_30920);
xnor U39287 (N_39287,N_30894,N_30092);
and U39288 (N_39288,N_30011,N_34388);
xnor U39289 (N_39289,N_32700,N_34756);
nand U39290 (N_39290,N_32069,N_33255);
nor U39291 (N_39291,N_33862,N_31584);
and U39292 (N_39292,N_33583,N_30840);
nor U39293 (N_39293,N_31733,N_31340);
nor U39294 (N_39294,N_34154,N_32089);
nand U39295 (N_39295,N_34523,N_33477);
nand U39296 (N_39296,N_30494,N_34076);
xnor U39297 (N_39297,N_33835,N_31119);
nand U39298 (N_39298,N_34847,N_30880);
nand U39299 (N_39299,N_31198,N_32440);
and U39300 (N_39300,N_30437,N_31183);
and U39301 (N_39301,N_34774,N_32535);
or U39302 (N_39302,N_30173,N_30227);
nand U39303 (N_39303,N_30475,N_34173);
nand U39304 (N_39304,N_31291,N_34409);
nand U39305 (N_39305,N_30670,N_32505);
nand U39306 (N_39306,N_33616,N_31475);
or U39307 (N_39307,N_30461,N_32405);
xnor U39308 (N_39308,N_30990,N_33197);
xor U39309 (N_39309,N_33774,N_32475);
nand U39310 (N_39310,N_32095,N_34106);
or U39311 (N_39311,N_32631,N_32170);
nor U39312 (N_39312,N_34958,N_31817);
xor U39313 (N_39313,N_31592,N_30375);
or U39314 (N_39314,N_30775,N_31358);
nand U39315 (N_39315,N_34637,N_31998);
xor U39316 (N_39316,N_30378,N_31569);
xor U39317 (N_39317,N_30196,N_34727);
xor U39318 (N_39318,N_33501,N_30344);
xnor U39319 (N_39319,N_31251,N_34363);
xor U39320 (N_39320,N_32955,N_31452);
nor U39321 (N_39321,N_30501,N_31927);
nor U39322 (N_39322,N_34315,N_33381);
nand U39323 (N_39323,N_34609,N_31626);
xnor U39324 (N_39324,N_33586,N_31932);
xnor U39325 (N_39325,N_34369,N_30779);
xnor U39326 (N_39326,N_33860,N_34577);
and U39327 (N_39327,N_34785,N_33150);
and U39328 (N_39328,N_32915,N_34715);
or U39329 (N_39329,N_31622,N_32914);
xnor U39330 (N_39330,N_34203,N_32977);
or U39331 (N_39331,N_32294,N_34091);
nor U39332 (N_39332,N_34019,N_30132);
and U39333 (N_39333,N_34236,N_30131);
or U39334 (N_39334,N_30719,N_34514);
nand U39335 (N_39335,N_33313,N_33644);
nor U39336 (N_39336,N_34067,N_32281);
nand U39337 (N_39337,N_32466,N_33039);
nand U39338 (N_39338,N_34749,N_32182);
xor U39339 (N_39339,N_31579,N_34473);
nor U39340 (N_39340,N_34726,N_33089);
nor U39341 (N_39341,N_33660,N_30884);
nand U39342 (N_39342,N_30876,N_34988);
or U39343 (N_39343,N_31939,N_31459);
or U39344 (N_39344,N_32604,N_31156);
or U39345 (N_39345,N_34906,N_34320);
xor U39346 (N_39346,N_32080,N_30971);
nor U39347 (N_39347,N_31351,N_33634);
and U39348 (N_39348,N_30995,N_33360);
nand U39349 (N_39349,N_33969,N_31429);
nor U39350 (N_39350,N_33637,N_30411);
xnor U39351 (N_39351,N_30661,N_32196);
nor U39352 (N_39352,N_31417,N_30546);
or U39353 (N_39353,N_33774,N_32148);
nor U39354 (N_39354,N_30084,N_33367);
xor U39355 (N_39355,N_32645,N_30068);
or U39356 (N_39356,N_33289,N_32655);
or U39357 (N_39357,N_31968,N_31608);
nor U39358 (N_39358,N_30338,N_32388);
nor U39359 (N_39359,N_33303,N_30234);
xor U39360 (N_39360,N_30152,N_34029);
xor U39361 (N_39361,N_32288,N_34680);
xor U39362 (N_39362,N_34497,N_33189);
or U39363 (N_39363,N_31103,N_30525);
and U39364 (N_39364,N_33723,N_33172);
nand U39365 (N_39365,N_31592,N_33634);
nor U39366 (N_39366,N_32169,N_30488);
xor U39367 (N_39367,N_34452,N_34116);
nand U39368 (N_39368,N_33591,N_31740);
and U39369 (N_39369,N_33009,N_33649);
xnor U39370 (N_39370,N_30468,N_31395);
nand U39371 (N_39371,N_32118,N_32770);
and U39372 (N_39372,N_30059,N_31249);
xor U39373 (N_39373,N_34060,N_34949);
nor U39374 (N_39374,N_32482,N_30671);
or U39375 (N_39375,N_30781,N_32299);
nor U39376 (N_39376,N_32830,N_34640);
xnor U39377 (N_39377,N_34306,N_31682);
xnor U39378 (N_39378,N_33470,N_30529);
nand U39379 (N_39379,N_34618,N_30636);
or U39380 (N_39380,N_33790,N_30379);
nor U39381 (N_39381,N_31822,N_31044);
nand U39382 (N_39382,N_32043,N_34728);
nand U39383 (N_39383,N_33188,N_31456);
or U39384 (N_39384,N_34226,N_32552);
xnor U39385 (N_39385,N_32775,N_33500);
nand U39386 (N_39386,N_33279,N_32424);
or U39387 (N_39387,N_33555,N_34640);
and U39388 (N_39388,N_33576,N_30078);
and U39389 (N_39389,N_32591,N_30590);
nand U39390 (N_39390,N_30701,N_32241);
and U39391 (N_39391,N_33670,N_31629);
and U39392 (N_39392,N_30535,N_31819);
or U39393 (N_39393,N_31572,N_31031);
nor U39394 (N_39394,N_34646,N_31803);
nor U39395 (N_39395,N_32827,N_34994);
and U39396 (N_39396,N_32059,N_34867);
nand U39397 (N_39397,N_30637,N_34680);
nand U39398 (N_39398,N_30209,N_34146);
or U39399 (N_39399,N_33924,N_30701);
nand U39400 (N_39400,N_31589,N_31242);
and U39401 (N_39401,N_30302,N_34051);
xor U39402 (N_39402,N_34515,N_32551);
or U39403 (N_39403,N_33146,N_31087);
and U39404 (N_39404,N_31694,N_34028);
xor U39405 (N_39405,N_32967,N_31829);
nor U39406 (N_39406,N_33723,N_31633);
nor U39407 (N_39407,N_34460,N_30409);
or U39408 (N_39408,N_34673,N_31175);
nor U39409 (N_39409,N_31775,N_31167);
and U39410 (N_39410,N_33054,N_33723);
and U39411 (N_39411,N_32094,N_32047);
xor U39412 (N_39412,N_31817,N_31782);
nor U39413 (N_39413,N_32897,N_32684);
and U39414 (N_39414,N_34699,N_34776);
and U39415 (N_39415,N_30031,N_32475);
and U39416 (N_39416,N_30680,N_33216);
and U39417 (N_39417,N_31274,N_32694);
nor U39418 (N_39418,N_30911,N_34448);
and U39419 (N_39419,N_30379,N_32785);
nand U39420 (N_39420,N_30561,N_34248);
xor U39421 (N_39421,N_32404,N_33461);
nand U39422 (N_39422,N_33177,N_34597);
nor U39423 (N_39423,N_30392,N_34198);
xor U39424 (N_39424,N_30422,N_34046);
nor U39425 (N_39425,N_33883,N_31465);
or U39426 (N_39426,N_34521,N_33797);
nor U39427 (N_39427,N_30067,N_31851);
or U39428 (N_39428,N_30334,N_32894);
and U39429 (N_39429,N_33018,N_32695);
nor U39430 (N_39430,N_30175,N_34091);
xnor U39431 (N_39431,N_34393,N_30845);
xnor U39432 (N_39432,N_30465,N_32540);
nor U39433 (N_39433,N_33821,N_30068);
and U39434 (N_39434,N_34453,N_34801);
nand U39435 (N_39435,N_30325,N_33102);
or U39436 (N_39436,N_31778,N_33765);
nand U39437 (N_39437,N_34174,N_34477);
nor U39438 (N_39438,N_30455,N_31099);
nor U39439 (N_39439,N_31641,N_33489);
xnor U39440 (N_39440,N_30384,N_30592);
or U39441 (N_39441,N_31954,N_34066);
and U39442 (N_39442,N_30514,N_32389);
xnor U39443 (N_39443,N_32567,N_32761);
nor U39444 (N_39444,N_34915,N_33950);
or U39445 (N_39445,N_34343,N_31401);
nor U39446 (N_39446,N_30739,N_34476);
nor U39447 (N_39447,N_32906,N_30366);
and U39448 (N_39448,N_30925,N_34969);
xor U39449 (N_39449,N_31851,N_31090);
or U39450 (N_39450,N_33670,N_31910);
or U39451 (N_39451,N_30665,N_33740);
nand U39452 (N_39452,N_32425,N_33247);
xor U39453 (N_39453,N_33528,N_31439);
xnor U39454 (N_39454,N_33584,N_31323);
nand U39455 (N_39455,N_31621,N_30097);
and U39456 (N_39456,N_31071,N_33406);
or U39457 (N_39457,N_31962,N_30458);
and U39458 (N_39458,N_30454,N_32946);
or U39459 (N_39459,N_30221,N_34027);
nor U39460 (N_39460,N_32720,N_30624);
nand U39461 (N_39461,N_31008,N_33334);
nand U39462 (N_39462,N_31396,N_34625);
nand U39463 (N_39463,N_31838,N_33139);
nor U39464 (N_39464,N_33893,N_32856);
or U39465 (N_39465,N_34290,N_34950);
nor U39466 (N_39466,N_34328,N_30715);
and U39467 (N_39467,N_32581,N_31592);
and U39468 (N_39468,N_32600,N_32699);
and U39469 (N_39469,N_34155,N_30551);
and U39470 (N_39470,N_31362,N_30920);
nand U39471 (N_39471,N_31006,N_31527);
nand U39472 (N_39472,N_31744,N_31741);
nand U39473 (N_39473,N_34482,N_32587);
and U39474 (N_39474,N_34573,N_30689);
and U39475 (N_39475,N_31434,N_34349);
and U39476 (N_39476,N_34213,N_33951);
nor U39477 (N_39477,N_30277,N_30464);
xnor U39478 (N_39478,N_33553,N_33084);
nand U39479 (N_39479,N_34745,N_32479);
or U39480 (N_39480,N_30829,N_31022);
xnor U39481 (N_39481,N_34497,N_31379);
and U39482 (N_39482,N_34283,N_30836);
nor U39483 (N_39483,N_33495,N_34760);
xor U39484 (N_39484,N_30384,N_32995);
or U39485 (N_39485,N_33522,N_30186);
nand U39486 (N_39486,N_30465,N_32182);
and U39487 (N_39487,N_33478,N_33402);
nand U39488 (N_39488,N_31298,N_30344);
xor U39489 (N_39489,N_31345,N_30796);
nor U39490 (N_39490,N_33583,N_30773);
nand U39491 (N_39491,N_33422,N_30434);
and U39492 (N_39492,N_32403,N_33031);
or U39493 (N_39493,N_32910,N_31008);
nor U39494 (N_39494,N_30119,N_30227);
nand U39495 (N_39495,N_31988,N_32088);
nand U39496 (N_39496,N_30276,N_31952);
nor U39497 (N_39497,N_31963,N_33524);
xnor U39498 (N_39498,N_32664,N_31870);
or U39499 (N_39499,N_31021,N_34196);
and U39500 (N_39500,N_31045,N_30156);
xnor U39501 (N_39501,N_31844,N_34147);
or U39502 (N_39502,N_30367,N_34649);
nor U39503 (N_39503,N_32845,N_32760);
xor U39504 (N_39504,N_34626,N_31622);
nor U39505 (N_39505,N_32583,N_31993);
or U39506 (N_39506,N_32928,N_32731);
nor U39507 (N_39507,N_30567,N_33385);
xor U39508 (N_39508,N_31244,N_33093);
xnor U39509 (N_39509,N_30739,N_32194);
or U39510 (N_39510,N_33573,N_30979);
xor U39511 (N_39511,N_33601,N_31812);
nor U39512 (N_39512,N_33891,N_30198);
and U39513 (N_39513,N_30935,N_32306);
nand U39514 (N_39514,N_34140,N_33434);
xnor U39515 (N_39515,N_34185,N_31013);
and U39516 (N_39516,N_30237,N_30141);
nand U39517 (N_39517,N_34973,N_34158);
or U39518 (N_39518,N_34033,N_31510);
or U39519 (N_39519,N_34193,N_33650);
or U39520 (N_39520,N_33744,N_34971);
xnor U39521 (N_39521,N_31530,N_31363);
or U39522 (N_39522,N_33692,N_30733);
nand U39523 (N_39523,N_32791,N_33098);
xnor U39524 (N_39524,N_30124,N_32245);
nand U39525 (N_39525,N_31751,N_31223);
xor U39526 (N_39526,N_33372,N_33155);
and U39527 (N_39527,N_30408,N_34719);
nor U39528 (N_39528,N_34234,N_33733);
or U39529 (N_39529,N_32779,N_34589);
nand U39530 (N_39530,N_33108,N_31414);
nand U39531 (N_39531,N_32401,N_30436);
nor U39532 (N_39532,N_32442,N_33963);
or U39533 (N_39533,N_32000,N_34060);
nor U39534 (N_39534,N_30627,N_30518);
and U39535 (N_39535,N_34733,N_33901);
nand U39536 (N_39536,N_30403,N_31109);
xor U39537 (N_39537,N_34111,N_30534);
or U39538 (N_39538,N_31563,N_33021);
and U39539 (N_39539,N_34750,N_32481);
nor U39540 (N_39540,N_32022,N_30627);
xor U39541 (N_39541,N_31099,N_31745);
xnor U39542 (N_39542,N_30135,N_33348);
or U39543 (N_39543,N_30393,N_33835);
xor U39544 (N_39544,N_33229,N_31283);
nor U39545 (N_39545,N_30676,N_33412);
xnor U39546 (N_39546,N_33769,N_34465);
nand U39547 (N_39547,N_32185,N_34635);
nand U39548 (N_39548,N_33281,N_32062);
xnor U39549 (N_39549,N_32221,N_32657);
xor U39550 (N_39550,N_33350,N_31790);
nor U39551 (N_39551,N_30424,N_34581);
and U39552 (N_39552,N_31774,N_30795);
or U39553 (N_39553,N_34189,N_32125);
nand U39554 (N_39554,N_34752,N_32762);
nand U39555 (N_39555,N_34499,N_34475);
and U39556 (N_39556,N_34157,N_31531);
and U39557 (N_39557,N_33557,N_33668);
or U39558 (N_39558,N_32460,N_32145);
xnor U39559 (N_39559,N_34387,N_34150);
or U39560 (N_39560,N_31153,N_30079);
xnor U39561 (N_39561,N_32286,N_33537);
or U39562 (N_39562,N_32736,N_30731);
nand U39563 (N_39563,N_32852,N_34964);
nand U39564 (N_39564,N_33240,N_31837);
xnor U39565 (N_39565,N_32402,N_32816);
and U39566 (N_39566,N_32169,N_30251);
nand U39567 (N_39567,N_31182,N_33437);
or U39568 (N_39568,N_33209,N_33106);
nor U39569 (N_39569,N_30707,N_34475);
nor U39570 (N_39570,N_30595,N_33399);
nor U39571 (N_39571,N_31548,N_31181);
or U39572 (N_39572,N_32340,N_32435);
or U39573 (N_39573,N_33405,N_30693);
nand U39574 (N_39574,N_31315,N_32432);
or U39575 (N_39575,N_34581,N_31651);
nand U39576 (N_39576,N_34101,N_32042);
nand U39577 (N_39577,N_34656,N_33425);
or U39578 (N_39578,N_31009,N_33055);
or U39579 (N_39579,N_32352,N_33372);
xor U39580 (N_39580,N_31394,N_32964);
nor U39581 (N_39581,N_34833,N_30376);
xnor U39582 (N_39582,N_30599,N_30160);
nor U39583 (N_39583,N_34424,N_31363);
nor U39584 (N_39584,N_32354,N_31012);
or U39585 (N_39585,N_34964,N_34160);
and U39586 (N_39586,N_34917,N_32052);
nor U39587 (N_39587,N_33844,N_33194);
xor U39588 (N_39588,N_31794,N_34580);
and U39589 (N_39589,N_30570,N_30747);
xor U39590 (N_39590,N_31087,N_32324);
or U39591 (N_39591,N_33213,N_31097);
xor U39592 (N_39592,N_33627,N_33341);
and U39593 (N_39593,N_34289,N_30486);
or U39594 (N_39594,N_30890,N_30128);
and U39595 (N_39595,N_33731,N_31696);
and U39596 (N_39596,N_31666,N_34454);
xor U39597 (N_39597,N_32940,N_31267);
xnor U39598 (N_39598,N_30025,N_30485);
or U39599 (N_39599,N_30800,N_33793);
and U39600 (N_39600,N_34723,N_34639);
nand U39601 (N_39601,N_30191,N_30126);
or U39602 (N_39602,N_34556,N_31973);
nor U39603 (N_39603,N_31541,N_34310);
nand U39604 (N_39604,N_34831,N_30585);
and U39605 (N_39605,N_32002,N_30283);
or U39606 (N_39606,N_30178,N_30697);
nor U39607 (N_39607,N_34111,N_30924);
and U39608 (N_39608,N_34343,N_32304);
and U39609 (N_39609,N_31753,N_30240);
or U39610 (N_39610,N_32862,N_30695);
and U39611 (N_39611,N_31207,N_30702);
nand U39612 (N_39612,N_33150,N_31330);
or U39613 (N_39613,N_34270,N_31471);
nor U39614 (N_39614,N_33832,N_32511);
and U39615 (N_39615,N_32088,N_31884);
nor U39616 (N_39616,N_33007,N_33106);
and U39617 (N_39617,N_33009,N_33038);
or U39618 (N_39618,N_31010,N_32712);
and U39619 (N_39619,N_33118,N_30970);
nand U39620 (N_39620,N_30016,N_31831);
xor U39621 (N_39621,N_31106,N_33333);
and U39622 (N_39622,N_34373,N_30250);
nor U39623 (N_39623,N_33562,N_31116);
and U39624 (N_39624,N_30314,N_30038);
or U39625 (N_39625,N_32395,N_32782);
and U39626 (N_39626,N_32791,N_34402);
nor U39627 (N_39627,N_34412,N_33599);
xnor U39628 (N_39628,N_31570,N_31323);
nor U39629 (N_39629,N_34774,N_33690);
nand U39630 (N_39630,N_33897,N_30959);
nor U39631 (N_39631,N_34335,N_33754);
and U39632 (N_39632,N_30294,N_34826);
and U39633 (N_39633,N_31086,N_34955);
and U39634 (N_39634,N_34934,N_30114);
or U39635 (N_39635,N_33063,N_31982);
xnor U39636 (N_39636,N_34658,N_34494);
nand U39637 (N_39637,N_33353,N_32832);
or U39638 (N_39638,N_34690,N_31360);
nor U39639 (N_39639,N_32842,N_31237);
nand U39640 (N_39640,N_31004,N_32184);
nand U39641 (N_39641,N_31313,N_31325);
xor U39642 (N_39642,N_33647,N_32127);
or U39643 (N_39643,N_34891,N_33628);
nand U39644 (N_39644,N_30315,N_30113);
or U39645 (N_39645,N_34125,N_33974);
nand U39646 (N_39646,N_31593,N_33657);
or U39647 (N_39647,N_33641,N_31644);
and U39648 (N_39648,N_33775,N_30309);
xor U39649 (N_39649,N_34119,N_30751);
nand U39650 (N_39650,N_31479,N_32597);
nor U39651 (N_39651,N_33788,N_30552);
xnor U39652 (N_39652,N_32055,N_32169);
nor U39653 (N_39653,N_33102,N_31245);
and U39654 (N_39654,N_32491,N_31475);
and U39655 (N_39655,N_34044,N_32391);
and U39656 (N_39656,N_31312,N_33222);
or U39657 (N_39657,N_30446,N_31210);
nand U39658 (N_39658,N_31151,N_31941);
or U39659 (N_39659,N_31724,N_33495);
or U39660 (N_39660,N_32605,N_32587);
or U39661 (N_39661,N_31115,N_33361);
nand U39662 (N_39662,N_34027,N_33298);
xnor U39663 (N_39663,N_31209,N_33415);
or U39664 (N_39664,N_31531,N_33996);
xnor U39665 (N_39665,N_32146,N_32157);
nor U39666 (N_39666,N_32958,N_32645);
xor U39667 (N_39667,N_33164,N_31174);
and U39668 (N_39668,N_33593,N_31954);
and U39669 (N_39669,N_33555,N_34154);
nor U39670 (N_39670,N_33763,N_34772);
nand U39671 (N_39671,N_32691,N_30327);
and U39672 (N_39672,N_30020,N_33473);
nor U39673 (N_39673,N_34895,N_33386);
nor U39674 (N_39674,N_30948,N_31587);
or U39675 (N_39675,N_32607,N_34748);
nand U39676 (N_39676,N_33002,N_33848);
nand U39677 (N_39677,N_33834,N_34541);
nand U39678 (N_39678,N_30783,N_31171);
nand U39679 (N_39679,N_30968,N_33038);
xnor U39680 (N_39680,N_31635,N_31276);
nor U39681 (N_39681,N_30946,N_34417);
xor U39682 (N_39682,N_33651,N_32127);
xnor U39683 (N_39683,N_31546,N_33336);
nor U39684 (N_39684,N_33092,N_32122);
or U39685 (N_39685,N_32041,N_33641);
nand U39686 (N_39686,N_33690,N_31077);
and U39687 (N_39687,N_34465,N_33783);
xor U39688 (N_39688,N_32658,N_34817);
or U39689 (N_39689,N_33367,N_30738);
xnor U39690 (N_39690,N_30233,N_31955);
xor U39691 (N_39691,N_31336,N_32174);
nor U39692 (N_39692,N_31939,N_32027);
xnor U39693 (N_39693,N_30073,N_32808);
xnor U39694 (N_39694,N_31952,N_32482);
nor U39695 (N_39695,N_33518,N_33482);
or U39696 (N_39696,N_33564,N_32188);
and U39697 (N_39697,N_32750,N_32588);
nand U39698 (N_39698,N_31108,N_34560);
nand U39699 (N_39699,N_32393,N_32408);
or U39700 (N_39700,N_33949,N_33664);
or U39701 (N_39701,N_33961,N_30739);
nor U39702 (N_39702,N_30185,N_32452);
xnor U39703 (N_39703,N_33482,N_32379);
nand U39704 (N_39704,N_30183,N_30369);
nand U39705 (N_39705,N_30164,N_30436);
nor U39706 (N_39706,N_31590,N_34920);
nor U39707 (N_39707,N_34170,N_31374);
nand U39708 (N_39708,N_31266,N_31473);
nand U39709 (N_39709,N_34829,N_33835);
xor U39710 (N_39710,N_33083,N_33422);
and U39711 (N_39711,N_30232,N_31502);
nor U39712 (N_39712,N_30643,N_32399);
and U39713 (N_39713,N_32255,N_31491);
nand U39714 (N_39714,N_32109,N_31522);
nor U39715 (N_39715,N_30805,N_32476);
or U39716 (N_39716,N_34603,N_31773);
nand U39717 (N_39717,N_32491,N_30845);
nand U39718 (N_39718,N_31631,N_31125);
xor U39719 (N_39719,N_33585,N_30652);
nor U39720 (N_39720,N_32612,N_34447);
xnor U39721 (N_39721,N_33528,N_32614);
nand U39722 (N_39722,N_30624,N_32485);
xor U39723 (N_39723,N_32141,N_31314);
nor U39724 (N_39724,N_34718,N_33915);
or U39725 (N_39725,N_30958,N_33835);
nand U39726 (N_39726,N_30300,N_33190);
and U39727 (N_39727,N_33083,N_34822);
xnor U39728 (N_39728,N_30285,N_30951);
nand U39729 (N_39729,N_32695,N_34436);
xor U39730 (N_39730,N_33690,N_33638);
or U39731 (N_39731,N_32460,N_33121);
and U39732 (N_39732,N_33014,N_30447);
nand U39733 (N_39733,N_33615,N_33110);
nor U39734 (N_39734,N_31699,N_34346);
or U39735 (N_39735,N_33094,N_33778);
xor U39736 (N_39736,N_33315,N_31730);
xnor U39737 (N_39737,N_34717,N_34517);
xnor U39738 (N_39738,N_31303,N_32430);
xnor U39739 (N_39739,N_34055,N_33211);
nor U39740 (N_39740,N_33496,N_33714);
xnor U39741 (N_39741,N_32459,N_34582);
nor U39742 (N_39742,N_34315,N_34815);
nand U39743 (N_39743,N_30431,N_34140);
nand U39744 (N_39744,N_31637,N_30538);
xnor U39745 (N_39745,N_34893,N_32616);
and U39746 (N_39746,N_33046,N_34126);
xnor U39747 (N_39747,N_30405,N_31265);
nor U39748 (N_39748,N_32732,N_33831);
nand U39749 (N_39749,N_34612,N_30491);
nand U39750 (N_39750,N_33259,N_34672);
or U39751 (N_39751,N_30768,N_32198);
and U39752 (N_39752,N_30177,N_32599);
nand U39753 (N_39753,N_32520,N_32126);
xor U39754 (N_39754,N_31167,N_32515);
or U39755 (N_39755,N_30715,N_30224);
and U39756 (N_39756,N_31977,N_31944);
xor U39757 (N_39757,N_34833,N_34532);
xor U39758 (N_39758,N_32059,N_30862);
nand U39759 (N_39759,N_34408,N_30977);
nand U39760 (N_39760,N_31219,N_30320);
nor U39761 (N_39761,N_34374,N_31560);
nand U39762 (N_39762,N_33384,N_30533);
xnor U39763 (N_39763,N_33846,N_33917);
nand U39764 (N_39764,N_33116,N_30202);
nor U39765 (N_39765,N_33494,N_30146);
or U39766 (N_39766,N_33683,N_30521);
and U39767 (N_39767,N_32246,N_31870);
nand U39768 (N_39768,N_32619,N_30048);
nand U39769 (N_39769,N_31078,N_33398);
or U39770 (N_39770,N_32717,N_31147);
xnor U39771 (N_39771,N_33467,N_34303);
and U39772 (N_39772,N_30402,N_34928);
and U39773 (N_39773,N_33855,N_33869);
and U39774 (N_39774,N_33600,N_34930);
or U39775 (N_39775,N_34821,N_30902);
or U39776 (N_39776,N_33266,N_32284);
and U39777 (N_39777,N_31544,N_33003);
and U39778 (N_39778,N_30297,N_33062);
nor U39779 (N_39779,N_34979,N_33098);
xnor U39780 (N_39780,N_30576,N_31045);
or U39781 (N_39781,N_32007,N_33508);
nor U39782 (N_39782,N_34042,N_32232);
nor U39783 (N_39783,N_33367,N_33848);
nand U39784 (N_39784,N_34302,N_30193);
or U39785 (N_39785,N_30562,N_33167);
xnor U39786 (N_39786,N_30214,N_32873);
xor U39787 (N_39787,N_34453,N_32359);
and U39788 (N_39788,N_31215,N_33422);
or U39789 (N_39789,N_32696,N_30007);
nand U39790 (N_39790,N_33402,N_32329);
nor U39791 (N_39791,N_34429,N_31959);
xor U39792 (N_39792,N_33126,N_34502);
nand U39793 (N_39793,N_34590,N_30037);
nor U39794 (N_39794,N_31441,N_31599);
or U39795 (N_39795,N_31082,N_31319);
and U39796 (N_39796,N_33513,N_32201);
nand U39797 (N_39797,N_32084,N_33545);
nand U39798 (N_39798,N_31358,N_32280);
nor U39799 (N_39799,N_31273,N_34126);
xnor U39800 (N_39800,N_34810,N_33408);
and U39801 (N_39801,N_32518,N_31762);
and U39802 (N_39802,N_31932,N_31244);
xnor U39803 (N_39803,N_33363,N_34457);
and U39804 (N_39804,N_30599,N_32477);
nor U39805 (N_39805,N_30552,N_31397);
xnor U39806 (N_39806,N_31062,N_34083);
nor U39807 (N_39807,N_30120,N_30651);
nor U39808 (N_39808,N_31918,N_30409);
and U39809 (N_39809,N_32848,N_34515);
or U39810 (N_39810,N_34051,N_32274);
or U39811 (N_39811,N_30357,N_31002);
and U39812 (N_39812,N_30679,N_33120);
nand U39813 (N_39813,N_33690,N_32662);
nand U39814 (N_39814,N_33887,N_34548);
nand U39815 (N_39815,N_33311,N_31340);
or U39816 (N_39816,N_32296,N_30030);
nor U39817 (N_39817,N_32054,N_34905);
nand U39818 (N_39818,N_34712,N_30275);
or U39819 (N_39819,N_33690,N_31080);
nor U39820 (N_39820,N_30815,N_30965);
nand U39821 (N_39821,N_30093,N_32517);
nor U39822 (N_39822,N_33621,N_31705);
or U39823 (N_39823,N_33611,N_33059);
and U39824 (N_39824,N_34111,N_34495);
nor U39825 (N_39825,N_33036,N_31298);
nor U39826 (N_39826,N_34846,N_31346);
xnor U39827 (N_39827,N_30591,N_34334);
or U39828 (N_39828,N_34929,N_33184);
and U39829 (N_39829,N_32417,N_30306);
or U39830 (N_39830,N_31376,N_34559);
and U39831 (N_39831,N_34601,N_31329);
xor U39832 (N_39832,N_30345,N_31717);
nor U39833 (N_39833,N_30088,N_32095);
and U39834 (N_39834,N_33957,N_32632);
nor U39835 (N_39835,N_31780,N_33414);
and U39836 (N_39836,N_30465,N_30764);
and U39837 (N_39837,N_33072,N_30335);
nor U39838 (N_39838,N_31013,N_30448);
or U39839 (N_39839,N_30401,N_33209);
nand U39840 (N_39840,N_33333,N_33711);
or U39841 (N_39841,N_33912,N_34059);
and U39842 (N_39842,N_30461,N_32360);
xor U39843 (N_39843,N_30855,N_30494);
nor U39844 (N_39844,N_32125,N_31522);
and U39845 (N_39845,N_34103,N_34595);
xnor U39846 (N_39846,N_32093,N_30750);
nand U39847 (N_39847,N_30282,N_33009);
nor U39848 (N_39848,N_32355,N_32226);
or U39849 (N_39849,N_33761,N_32429);
nand U39850 (N_39850,N_32709,N_30247);
nor U39851 (N_39851,N_32076,N_32052);
and U39852 (N_39852,N_31100,N_31013);
nor U39853 (N_39853,N_34180,N_32477);
nor U39854 (N_39854,N_32006,N_33662);
and U39855 (N_39855,N_34426,N_34791);
nand U39856 (N_39856,N_30669,N_30529);
or U39857 (N_39857,N_34829,N_33081);
or U39858 (N_39858,N_30581,N_32293);
xor U39859 (N_39859,N_31297,N_31508);
nor U39860 (N_39860,N_32643,N_33161);
nor U39861 (N_39861,N_32575,N_32975);
xnor U39862 (N_39862,N_30311,N_34113);
nand U39863 (N_39863,N_32615,N_32456);
nand U39864 (N_39864,N_32219,N_31189);
nor U39865 (N_39865,N_32102,N_30586);
or U39866 (N_39866,N_32005,N_34146);
nor U39867 (N_39867,N_32403,N_33748);
nand U39868 (N_39868,N_30505,N_34155);
nor U39869 (N_39869,N_33492,N_32730);
nand U39870 (N_39870,N_30783,N_30774);
nand U39871 (N_39871,N_31933,N_33541);
nor U39872 (N_39872,N_33817,N_30157);
nor U39873 (N_39873,N_32969,N_32562);
nand U39874 (N_39874,N_31516,N_31377);
and U39875 (N_39875,N_32866,N_34783);
nor U39876 (N_39876,N_32538,N_31056);
xnor U39877 (N_39877,N_32047,N_34493);
or U39878 (N_39878,N_34075,N_30337);
nand U39879 (N_39879,N_32446,N_30471);
xor U39880 (N_39880,N_33607,N_30903);
or U39881 (N_39881,N_31522,N_31200);
and U39882 (N_39882,N_34789,N_34265);
nor U39883 (N_39883,N_34804,N_32740);
and U39884 (N_39884,N_32925,N_32030);
nor U39885 (N_39885,N_34798,N_33177);
xnor U39886 (N_39886,N_34905,N_32206);
nand U39887 (N_39887,N_33951,N_30484);
xor U39888 (N_39888,N_31167,N_31616);
nor U39889 (N_39889,N_32478,N_30586);
or U39890 (N_39890,N_34373,N_30499);
xnor U39891 (N_39891,N_34958,N_32630);
nor U39892 (N_39892,N_33433,N_31443);
and U39893 (N_39893,N_33596,N_31470);
nand U39894 (N_39894,N_30907,N_31017);
nor U39895 (N_39895,N_32045,N_31314);
and U39896 (N_39896,N_32376,N_32355);
nor U39897 (N_39897,N_34251,N_33724);
or U39898 (N_39898,N_34361,N_32915);
nand U39899 (N_39899,N_31146,N_32874);
nor U39900 (N_39900,N_34131,N_34683);
and U39901 (N_39901,N_30229,N_33647);
and U39902 (N_39902,N_34871,N_31405);
nor U39903 (N_39903,N_31174,N_30293);
nand U39904 (N_39904,N_33751,N_30723);
and U39905 (N_39905,N_33113,N_30413);
and U39906 (N_39906,N_31754,N_32376);
and U39907 (N_39907,N_31295,N_32755);
xor U39908 (N_39908,N_30273,N_34564);
nand U39909 (N_39909,N_31623,N_30974);
nand U39910 (N_39910,N_34398,N_34646);
and U39911 (N_39911,N_33465,N_33805);
and U39912 (N_39912,N_32274,N_33401);
and U39913 (N_39913,N_33640,N_30680);
and U39914 (N_39914,N_32634,N_34343);
nor U39915 (N_39915,N_33545,N_32861);
nor U39916 (N_39916,N_33845,N_30644);
or U39917 (N_39917,N_34915,N_33356);
nor U39918 (N_39918,N_34139,N_34181);
or U39919 (N_39919,N_30961,N_32088);
and U39920 (N_39920,N_32923,N_31992);
and U39921 (N_39921,N_34986,N_34701);
and U39922 (N_39922,N_30485,N_30652);
or U39923 (N_39923,N_32786,N_30394);
nand U39924 (N_39924,N_30566,N_33868);
xnor U39925 (N_39925,N_32560,N_30110);
nand U39926 (N_39926,N_31133,N_32619);
nand U39927 (N_39927,N_34290,N_33275);
nand U39928 (N_39928,N_31302,N_33546);
nor U39929 (N_39929,N_34844,N_34222);
xnor U39930 (N_39930,N_34008,N_30186);
nor U39931 (N_39931,N_30755,N_33467);
and U39932 (N_39932,N_32386,N_33483);
nor U39933 (N_39933,N_31801,N_34356);
nand U39934 (N_39934,N_30622,N_32998);
and U39935 (N_39935,N_31622,N_33030);
or U39936 (N_39936,N_33323,N_34244);
and U39937 (N_39937,N_30412,N_30396);
or U39938 (N_39938,N_34408,N_34866);
nand U39939 (N_39939,N_32210,N_32691);
and U39940 (N_39940,N_33793,N_32285);
or U39941 (N_39941,N_32549,N_33714);
xor U39942 (N_39942,N_34765,N_30043);
or U39943 (N_39943,N_30666,N_34942);
nand U39944 (N_39944,N_32325,N_33060);
and U39945 (N_39945,N_33333,N_34561);
nor U39946 (N_39946,N_33676,N_34739);
and U39947 (N_39947,N_33492,N_30355);
or U39948 (N_39948,N_33682,N_31867);
and U39949 (N_39949,N_30515,N_30472);
nand U39950 (N_39950,N_33646,N_31730);
and U39951 (N_39951,N_33301,N_31764);
xnor U39952 (N_39952,N_33070,N_32125);
nand U39953 (N_39953,N_34296,N_30087);
or U39954 (N_39954,N_31599,N_34637);
and U39955 (N_39955,N_33766,N_32650);
xor U39956 (N_39956,N_31779,N_30480);
and U39957 (N_39957,N_34555,N_32760);
and U39958 (N_39958,N_33653,N_33727);
xnor U39959 (N_39959,N_32420,N_34065);
xnor U39960 (N_39960,N_30385,N_34631);
nand U39961 (N_39961,N_33405,N_32797);
nand U39962 (N_39962,N_34368,N_30930);
or U39963 (N_39963,N_33377,N_33997);
nor U39964 (N_39964,N_30301,N_32985);
xnor U39965 (N_39965,N_30018,N_32727);
and U39966 (N_39966,N_32754,N_31189);
nand U39967 (N_39967,N_31710,N_31775);
xor U39968 (N_39968,N_32624,N_30856);
nand U39969 (N_39969,N_30075,N_32689);
nand U39970 (N_39970,N_32486,N_34102);
and U39971 (N_39971,N_32379,N_32065);
nand U39972 (N_39972,N_31250,N_31173);
nor U39973 (N_39973,N_33954,N_32664);
nand U39974 (N_39974,N_33910,N_34272);
or U39975 (N_39975,N_32041,N_34494);
or U39976 (N_39976,N_32559,N_33787);
or U39977 (N_39977,N_33452,N_33253);
nand U39978 (N_39978,N_34982,N_31202);
and U39979 (N_39979,N_33147,N_30275);
nor U39980 (N_39980,N_30774,N_30568);
or U39981 (N_39981,N_33795,N_30858);
or U39982 (N_39982,N_33149,N_33543);
xor U39983 (N_39983,N_32000,N_30743);
nand U39984 (N_39984,N_32318,N_34688);
nand U39985 (N_39985,N_30987,N_34522);
or U39986 (N_39986,N_33922,N_32533);
xnor U39987 (N_39987,N_32639,N_30012);
nor U39988 (N_39988,N_33760,N_32977);
xor U39989 (N_39989,N_33153,N_31760);
nor U39990 (N_39990,N_33442,N_33670);
or U39991 (N_39991,N_34796,N_30708);
or U39992 (N_39992,N_34901,N_34923);
xor U39993 (N_39993,N_31518,N_31560);
xnor U39994 (N_39994,N_32327,N_33124);
xnor U39995 (N_39995,N_34774,N_34080);
and U39996 (N_39996,N_34499,N_33624);
or U39997 (N_39997,N_34551,N_31085);
or U39998 (N_39998,N_31365,N_33952);
xor U39999 (N_39999,N_34298,N_34112);
nor U40000 (N_40000,N_35964,N_35383);
nand U40001 (N_40001,N_37307,N_37332);
and U40002 (N_40002,N_38982,N_37877);
and U40003 (N_40003,N_38815,N_36745);
and U40004 (N_40004,N_39690,N_35620);
or U40005 (N_40005,N_35651,N_35727);
xor U40006 (N_40006,N_36403,N_39679);
and U40007 (N_40007,N_39120,N_39812);
xnor U40008 (N_40008,N_38302,N_35874);
nand U40009 (N_40009,N_38887,N_36656);
xor U40010 (N_40010,N_35487,N_39963);
and U40011 (N_40011,N_39699,N_39653);
nor U40012 (N_40012,N_37158,N_36918);
nand U40013 (N_40013,N_35406,N_37760);
and U40014 (N_40014,N_35098,N_37812);
and U40015 (N_40015,N_36687,N_38252);
xnor U40016 (N_40016,N_36516,N_35732);
nor U40017 (N_40017,N_39965,N_37287);
nand U40018 (N_40018,N_35291,N_37295);
nor U40019 (N_40019,N_39429,N_39234);
nand U40020 (N_40020,N_37666,N_37777);
nand U40021 (N_40021,N_35841,N_36291);
nand U40022 (N_40022,N_35925,N_39005);
and U40023 (N_40023,N_38674,N_37847);
nor U40024 (N_40024,N_36222,N_39416);
nor U40025 (N_40025,N_38439,N_38695);
nor U40026 (N_40026,N_38005,N_36762);
xnor U40027 (N_40027,N_38200,N_35354);
nor U40028 (N_40028,N_39177,N_37586);
nand U40029 (N_40029,N_37425,N_36337);
nor U40030 (N_40030,N_36318,N_39146);
and U40031 (N_40031,N_35879,N_36966);
xor U40032 (N_40032,N_37589,N_38763);
and U40033 (N_40033,N_37284,N_38469);
or U40034 (N_40034,N_36430,N_35920);
and U40035 (N_40035,N_36047,N_39706);
nand U40036 (N_40036,N_36755,N_36088);
xnor U40037 (N_40037,N_35373,N_35361);
and U40038 (N_40038,N_35049,N_38744);
nor U40039 (N_40039,N_35972,N_36915);
or U40040 (N_40040,N_37981,N_38682);
nor U40041 (N_40041,N_38407,N_39869);
nand U40042 (N_40042,N_38412,N_37836);
xor U40043 (N_40043,N_35808,N_37257);
nor U40044 (N_40044,N_36532,N_35193);
nor U40045 (N_40045,N_38890,N_35061);
or U40046 (N_40046,N_38280,N_36339);
and U40047 (N_40047,N_37041,N_38352);
nand U40048 (N_40048,N_36346,N_37514);
nor U40049 (N_40049,N_37357,N_36085);
xnor U40050 (N_40050,N_37634,N_37173);
or U40051 (N_40051,N_37242,N_38765);
nor U40052 (N_40052,N_37545,N_38038);
nand U40053 (N_40053,N_36932,N_39619);
and U40054 (N_40054,N_39474,N_37921);
xor U40055 (N_40055,N_35809,N_39825);
and U40056 (N_40056,N_39767,N_35752);
xor U40057 (N_40057,N_38006,N_35054);
nor U40058 (N_40058,N_39654,N_37297);
nor U40059 (N_40059,N_39190,N_39083);
nand U40060 (N_40060,N_39166,N_36174);
nand U40061 (N_40061,N_35516,N_35788);
nor U40062 (N_40062,N_39307,N_37535);
nand U40063 (N_40063,N_35420,N_38715);
and U40064 (N_40064,N_39249,N_38635);
and U40065 (N_40065,N_35960,N_37486);
nand U40066 (N_40066,N_37077,N_39837);
nand U40067 (N_40067,N_36843,N_38400);
nand U40068 (N_40068,N_38366,N_36999);
xnor U40069 (N_40069,N_36816,N_35772);
nor U40070 (N_40070,N_36317,N_37005);
and U40071 (N_40071,N_35648,N_37341);
nor U40072 (N_40072,N_35915,N_37115);
nor U40073 (N_40073,N_39247,N_37048);
or U40074 (N_40074,N_36013,N_38841);
xor U40075 (N_40075,N_37315,N_36863);
nand U40076 (N_40076,N_35942,N_36369);
nor U40077 (N_40077,N_36647,N_35297);
xor U40078 (N_40078,N_39324,N_38546);
nand U40079 (N_40079,N_38466,N_38315);
xor U40080 (N_40080,N_38324,N_38292);
and U40081 (N_40081,N_38095,N_36784);
xor U40082 (N_40082,N_39758,N_35904);
nor U40083 (N_40083,N_38020,N_37478);
xor U40084 (N_40084,N_38909,N_36846);
nor U40085 (N_40085,N_36670,N_37116);
or U40086 (N_40086,N_36009,N_38316);
nor U40087 (N_40087,N_37922,N_35853);
xor U40088 (N_40088,N_36404,N_35932);
or U40089 (N_40089,N_36059,N_37467);
nor U40090 (N_40090,N_39052,N_39788);
or U40091 (N_40091,N_36227,N_37718);
nand U40092 (N_40092,N_38396,N_39674);
nand U40093 (N_40093,N_38073,N_35187);
xor U40094 (N_40094,N_35008,N_38150);
nor U40095 (N_40095,N_36436,N_39523);
xnor U40096 (N_40096,N_35262,N_37905);
nor U40097 (N_40097,N_36795,N_37319);
nor U40098 (N_40098,N_35774,N_35997);
nor U40099 (N_40099,N_36431,N_39150);
xor U40100 (N_40100,N_36472,N_37624);
and U40101 (N_40101,N_38797,N_35047);
xnor U40102 (N_40102,N_37113,N_39872);
or U40103 (N_40103,N_39731,N_38092);
nand U40104 (N_40104,N_38064,N_39535);
nand U40105 (N_40105,N_37529,N_35536);
or U40106 (N_40106,N_38333,N_36434);
xor U40107 (N_40107,N_35407,N_36287);
nor U40108 (N_40108,N_36207,N_39849);
and U40109 (N_40109,N_35566,N_35756);
or U40110 (N_40110,N_36993,N_39387);
xor U40111 (N_40111,N_36695,N_36831);
nor U40112 (N_40112,N_35987,N_37261);
xnor U40113 (N_40113,N_37794,N_37952);
xor U40114 (N_40114,N_39283,N_38217);
nand U40115 (N_40115,N_35303,N_38372);
or U40116 (N_40116,N_37194,N_35348);
nand U40117 (N_40117,N_38055,N_36374);
xnor U40118 (N_40118,N_35132,N_35873);
and U40119 (N_40119,N_39348,N_38694);
xor U40120 (N_40120,N_38941,N_39286);
nand U40121 (N_40121,N_37442,N_35835);
xnor U40122 (N_40122,N_39040,N_37738);
and U40123 (N_40123,N_39204,N_39484);
and U40124 (N_40124,N_39569,N_37903);
nor U40125 (N_40125,N_37958,N_38732);
xor U40126 (N_40126,N_35424,N_36806);
or U40127 (N_40127,N_37675,N_39148);
or U40128 (N_40128,N_36746,N_37415);
nand U40129 (N_40129,N_38883,N_38937);
nor U40130 (N_40130,N_36355,N_36113);
or U40131 (N_40131,N_36652,N_37983);
nor U40132 (N_40132,N_35497,N_37094);
and U40133 (N_40133,N_38996,N_39514);
nor U40134 (N_40134,N_39284,N_36916);
xnor U40135 (N_40135,N_39054,N_35466);
or U40136 (N_40136,N_38168,N_35454);
and U40137 (N_40137,N_38123,N_39675);
nand U40138 (N_40138,N_38461,N_35699);
or U40139 (N_40139,N_35021,N_39353);
nand U40140 (N_40140,N_39330,N_38985);
and U40141 (N_40141,N_36127,N_35577);
nand U40142 (N_40142,N_36944,N_38170);
and U40143 (N_40143,N_37202,N_36739);
or U40144 (N_40144,N_37197,N_36248);
or U40145 (N_40145,N_35686,N_36734);
nand U40146 (N_40146,N_39102,N_38182);
nand U40147 (N_40147,N_38404,N_39055);
nand U40148 (N_40148,N_35689,N_35502);
nor U40149 (N_40149,N_39343,N_37108);
nor U40150 (N_40150,N_37410,N_36552);
or U40151 (N_40151,N_38047,N_37728);
and U40152 (N_40152,N_36775,N_36428);
and U40153 (N_40153,N_38299,N_37265);
xor U40154 (N_40154,N_37079,N_39843);
xnor U40155 (N_40155,N_36074,N_38606);
or U40156 (N_40156,N_36061,N_38048);
nor U40157 (N_40157,N_36189,N_36931);
xnor U40158 (N_40158,N_38801,N_36273);
xnor U40159 (N_40159,N_37886,N_38238);
nand U40160 (N_40160,N_38183,N_38338);
and U40161 (N_40161,N_39496,N_35740);
or U40162 (N_40162,N_38178,N_37676);
nor U40163 (N_40163,N_38339,N_39199);
xnor U40164 (N_40164,N_38519,N_36353);
xor U40165 (N_40165,N_37608,N_36783);
and U40166 (N_40166,N_35555,N_36922);
and U40167 (N_40167,N_37959,N_36073);
xnor U40168 (N_40168,N_39665,N_37405);
nor U40169 (N_40169,N_38179,N_38709);
xor U40170 (N_40170,N_37244,N_37021);
nor U40171 (N_40171,N_37204,N_39473);
or U40172 (N_40172,N_38533,N_39615);
nand U40173 (N_40173,N_37837,N_36890);
nor U40174 (N_40174,N_38022,N_38158);
and U40175 (N_40175,N_37571,N_39573);
nand U40176 (N_40176,N_35445,N_38241);
nor U40177 (N_40177,N_36104,N_37092);
nor U40178 (N_40178,N_36402,N_38872);
nand U40179 (N_40179,N_35831,N_38211);
xor U40180 (N_40180,N_38290,N_38652);
nor U40181 (N_40181,N_35825,N_36630);
or U40182 (N_40182,N_35485,N_38912);
or U40183 (N_40183,N_38470,N_37432);
nand U40184 (N_40184,N_38271,N_35171);
nor U40185 (N_40185,N_38782,N_37653);
xor U40186 (N_40186,N_37632,N_38714);
or U40187 (N_40187,N_39076,N_37692);
nand U40188 (N_40188,N_36939,N_37440);
nor U40189 (N_40189,N_39013,N_36473);
nand U40190 (N_40190,N_35814,N_38403);
nor U40191 (N_40191,N_35733,N_35030);
nor U40192 (N_40192,N_37208,N_35387);
or U40193 (N_40193,N_35690,N_35881);
xor U40194 (N_40194,N_39003,N_36251);
nor U40195 (N_40195,N_35544,N_36348);
xnor U40196 (N_40196,N_38457,N_35267);
or U40197 (N_40197,N_36870,N_37835);
nor U40198 (N_40198,N_37895,N_36505);
or U40199 (N_40199,N_35575,N_38193);
xnor U40200 (N_40200,N_38645,N_38813);
xnor U40201 (N_40201,N_36850,N_39807);
or U40202 (N_40202,N_38460,N_38831);
or U40203 (N_40203,N_36896,N_35705);
xor U40204 (N_40204,N_37593,N_38787);
nand U40205 (N_40205,N_39263,N_35545);
or U40206 (N_40206,N_38676,N_38573);
xnor U40207 (N_40207,N_38382,N_37125);
and U40208 (N_40208,N_35244,N_36439);
nor U40209 (N_40209,N_35617,N_36672);
or U40210 (N_40210,N_35003,N_35020);
and U40211 (N_40211,N_37627,N_37516);
xnor U40212 (N_40212,N_36096,N_37266);
nand U40213 (N_40213,N_37599,N_39881);
or U40214 (N_40214,N_35463,N_39351);
xor U40215 (N_40215,N_39051,N_37303);
or U40216 (N_40216,N_36016,N_35693);
and U40217 (N_40217,N_36959,N_39585);
xnor U40218 (N_40218,N_37147,N_39396);
xnor U40219 (N_40219,N_37160,N_37117);
and U40220 (N_40220,N_35358,N_37397);
and U40221 (N_40221,N_35556,N_38675);
nand U40222 (N_40222,N_35687,N_38504);
or U40223 (N_40223,N_39490,N_37166);
nor U40224 (N_40224,N_37640,N_36954);
or U40225 (N_40225,N_39411,N_37664);
nor U40226 (N_40226,N_39684,N_37822);
nor U40227 (N_40227,N_38938,N_39913);
nand U40228 (N_40228,N_36570,N_37681);
or U40229 (N_40229,N_36155,N_39250);
nor U40230 (N_40230,N_36362,N_37396);
xnor U40231 (N_40231,N_38216,N_36464);
nand U40232 (N_40232,N_37230,N_39647);
and U40233 (N_40233,N_39538,N_35309);
or U40234 (N_40234,N_37550,N_35522);
nand U40235 (N_40235,N_36773,N_35869);
and U40236 (N_40236,N_38899,N_39466);
nand U40237 (N_40237,N_39791,N_36089);
nor U40238 (N_40238,N_35965,N_37657);
nor U40239 (N_40239,N_36536,N_36512);
nor U40240 (N_40240,N_36469,N_35074);
and U40241 (N_40241,N_37036,N_39157);
nor U40242 (N_40242,N_36810,N_37018);
nand U40243 (N_40243,N_36848,N_38525);
or U40244 (N_40244,N_36812,N_37468);
or U40245 (N_40245,N_38214,N_37190);
nand U40246 (N_40246,N_39281,N_39427);
or U40247 (N_40247,N_39225,N_36470);
and U40248 (N_40248,N_36530,N_35966);
or U40249 (N_40249,N_39532,N_39959);
or U40250 (N_40250,N_36090,N_38791);
nand U40251 (N_40251,N_39093,N_39238);
or U40252 (N_40252,N_36706,N_35338);
nor U40253 (N_40253,N_36692,N_35294);
xor U40254 (N_40254,N_35618,N_38219);
or U40255 (N_40255,N_39754,N_35728);
nand U40256 (N_40256,N_37789,N_36608);
xor U40257 (N_40257,N_37485,N_37459);
or U40258 (N_40258,N_38993,N_35156);
or U40259 (N_40259,N_39046,N_36114);
and U40260 (N_40260,N_36343,N_37621);
xnor U40261 (N_40261,N_36020,N_37540);
nand U40262 (N_40262,N_36575,N_39109);
nor U40263 (N_40263,N_38229,N_36804);
nand U40264 (N_40264,N_39705,N_37626);
and U40265 (N_40265,N_39709,N_36751);
or U40266 (N_40266,N_36933,N_36057);
and U40267 (N_40267,N_37652,N_36069);
nor U40268 (N_40268,N_36603,N_38903);
nor U40269 (N_40269,N_35713,N_38431);
nor U40270 (N_40270,N_36830,N_36418);
or U40271 (N_40271,N_39349,N_36507);
nor U40272 (N_40272,N_38383,N_35432);
or U40273 (N_40273,N_39802,N_35683);
or U40274 (N_40274,N_37806,N_37370);
nand U40275 (N_40275,N_39776,N_35855);
or U40276 (N_40276,N_36129,N_38049);
xor U40277 (N_40277,N_37391,N_36278);
or U40278 (N_40278,N_39126,N_38177);
xnor U40279 (N_40279,N_39629,N_36025);
nor U40280 (N_40280,N_37040,N_35051);
nand U40281 (N_40281,N_39049,N_38343);
nor U40282 (N_40282,N_35860,N_36393);
nand U40283 (N_40283,N_39982,N_35847);
nand U40284 (N_40284,N_35902,N_36881);
or U40285 (N_40285,N_39071,N_39724);
and U40286 (N_40286,N_38161,N_35255);
xor U40287 (N_40287,N_38281,N_37200);
or U40288 (N_40288,N_35684,N_35498);
nor U40289 (N_40289,N_37049,N_35937);
nor U40290 (N_40290,N_39394,N_35608);
nor U40291 (N_40291,N_35196,N_39118);
nor U40292 (N_40292,N_36917,N_38794);
nand U40293 (N_40293,N_35658,N_35359);
and U40294 (N_40294,N_35718,N_35946);
or U40295 (N_40295,N_36257,N_36845);
nand U40296 (N_40296,N_39379,N_35489);
or U40297 (N_40297,N_37351,N_35521);
nand U40298 (N_40298,N_36477,N_38629);
nor U40299 (N_40299,N_37504,N_38206);
and U40300 (N_40300,N_37180,N_38873);
or U40301 (N_40301,N_36313,N_35242);
nand U40302 (N_40302,N_37600,N_36640);
and U40303 (N_40303,N_38423,N_35711);
xnor U40304 (N_40304,N_37778,N_36054);
xor U40305 (N_40305,N_39727,N_39056);
nand U40306 (N_40306,N_39252,N_38735);
nand U40307 (N_40307,N_36225,N_36261);
or U40308 (N_40308,N_35706,N_35264);
and U40309 (N_40309,N_37583,N_39518);
and U40310 (N_40310,N_39625,N_38154);
or U40311 (N_40311,N_38011,N_38349);
and U40312 (N_40312,N_39441,N_38253);
and U40313 (N_40313,N_39676,N_37034);
or U40314 (N_40314,N_35958,N_35823);
nand U40315 (N_40315,N_35908,N_36501);
or U40316 (N_40316,N_37068,N_36951);
nand U40317 (N_40317,N_35231,N_38348);
nand U40318 (N_40318,N_39301,N_35273);
nand U40319 (N_40319,N_38432,N_37126);
or U40320 (N_40320,N_37022,N_35628);
nor U40321 (N_40321,N_37654,N_39189);
nor U40322 (N_40322,N_37637,N_36441);
nor U40323 (N_40323,N_37365,N_37349);
nand U40324 (N_40324,N_38931,N_36923);
and U40325 (N_40325,N_37454,N_37517);
nand U40326 (N_40326,N_39472,N_37274);
nand U40327 (N_40327,N_38991,N_38294);
or U40328 (N_40328,N_38897,N_35458);
and U40329 (N_40329,N_39522,N_38900);
xor U40330 (N_40330,N_37706,N_39403);
or U40331 (N_40331,N_39814,N_37098);
or U40332 (N_40332,N_35675,N_38388);
or U40333 (N_40333,N_36829,N_35222);
and U40334 (N_40334,N_36290,N_37787);
nand U40335 (N_40335,N_39710,N_39392);
nor U40336 (N_40336,N_37017,N_36712);
nand U40337 (N_40337,N_37723,N_35765);
or U40338 (N_40338,N_39001,N_37544);
xnor U40339 (N_40339,N_38494,N_39509);
or U40340 (N_40340,N_37704,N_36970);
and U40341 (N_40341,N_36002,N_39021);
xnor U40342 (N_40342,N_36480,N_38820);
or U40343 (N_40343,N_37590,N_36503);
nand U40344 (N_40344,N_38809,N_37838);
nor U40345 (N_40345,N_37603,N_39289);
xor U40346 (N_40346,N_39431,N_37570);
and U40347 (N_40347,N_37286,N_36569);
nand U40348 (N_40348,N_39402,N_35571);
nor U40349 (N_40349,N_36323,N_35583);
nand U40350 (N_40350,N_37920,N_39744);
xor U40351 (N_40351,N_35990,N_39988);
and U40352 (N_40352,N_35165,N_38990);
xor U40353 (N_40353,N_39091,N_35661);
xor U40354 (N_40354,N_35982,N_38152);
nand U40355 (N_40355,N_35306,N_39748);
or U40356 (N_40356,N_38538,N_37890);
nor U40357 (N_40357,N_35475,N_38600);
and U40358 (N_40358,N_39065,N_35708);
and U40359 (N_40359,N_36904,N_39242);
and U40360 (N_40360,N_39012,N_35325);
nor U40361 (N_40361,N_39422,N_38823);
xnor U40362 (N_40362,N_38223,N_37631);
and U40363 (N_40363,N_38313,N_36022);
nor U40364 (N_40364,N_36188,N_35532);
or U40365 (N_40365,N_37975,N_35897);
nor U40366 (N_40366,N_36794,N_39438);
or U40367 (N_40367,N_37299,N_37594);
and U40368 (N_40368,N_36875,N_38942);
and U40369 (N_40369,N_39401,N_36466);
and U40370 (N_40370,N_35327,N_35069);
and U40371 (N_40371,N_37325,N_38826);
or U40372 (N_40372,N_39898,N_35593);
and U40373 (N_40373,N_35143,N_39185);
and U40374 (N_40374,N_36345,N_39634);
nor U40375 (N_40375,N_36754,N_38035);
nor U40376 (N_40376,N_36181,N_37572);
and U40377 (N_40377,N_35252,N_39677);
nand U40378 (N_40378,N_35213,N_39607);
and U40379 (N_40379,N_36112,N_37699);
or U40380 (N_40380,N_36731,N_37393);
or U40381 (N_40381,N_35922,N_36003);
nand U40382 (N_40382,N_36052,N_35096);
nand U40383 (N_40383,N_39099,N_36124);
nor U40384 (N_40384,N_37526,N_39639);
xor U40385 (N_40385,N_38384,N_35806);
xor U40386 (N_40386,N_37219,N_38967);
nand U40387 (N_40387,N_39486,N_35111);
xor U40388 (N_40388,N_36130,N_36252);
and U40389 (N_40389,N_36209,N_37830);
nor U40390 (N_40390,N_38307,N_36793);
xnor U40391 (N_40391,N_38148,N_39041);
or U40392 (N_40392,N_37999,N_38074);
xnor U40393 (N_40393,N_39385,N_36215);
nor U40394 (N_40394,N_37177,N_37974);
xnor U40395 (N_40395,N_39471,N_38522);
and U40396 (N_40396,N_35892,N_38895);
and U40397 (N_40397,N_38818,N_38187);
and U40398 (N_40398,N_39646,N_35924);
and U40399 (N_40399,N_39506,N_39213);
xnor U40400 (N_40400,N_37604,N_38854);
or U40401 (N_40401,N_38567,N_37502);
nor U40402 (N_40402,N_39752,N_36254);
xnor U40403 (N_40403,N_38118,N_36102);
or U40404 (N_40404,N_37655,N_38127);
nand U40405 (N_40405,N_38594,N_38246);
or U40406 (N_40406,N_36468,N_36325);
nand U40407 (N_40407,N_37580,N_39830);
nand U40408 (N_40408,N_35889,N_38590);
xnor U40409 (N_40409,N_39124,N_38534);
and U40410 (N_40410,N_35933,N_37076);
xnor U40411 (N_40411,N_36178,N_35533);
nor U40412 (N_40412,N_36737,N_36067);
or U40413 (N_40413,N_37344,N_38130);
or U40414 (N_40414,N_35245,N_37457);
xor U40415 (N_40415,N_35207,N_35416);
nand U40416 (N_40416,N_36150,N_39333);
or U40417 (N_40417,N_37617,N_36839);
nor U40418 (N_40418,N_35033,N_38162);
or U40419 (N_40419,N_37118,N_36239);
xnor U40420 (N_40420,N_39191,N_39681);
nor U40421 (N_40421,N_38926,N_35603);
nand U40422 (N_40422,N_37088,N_35175);
nand U40423 (N_40423,N_36985,N_37871);
or U40424 (N_40424,N_37917,N_38669);
or U40425 (N_40425,N_37611,N_35610);
nor U40426 (N_40426,N_39412,N_39482);
xor U40427 (N_40427,N_35017,N_36892);
xnor U40428 (N_40428,N_37527,N_35313);
nand U40429 (N_40429,N_35319,N_38019);
and U40430 (N_40430,N_38257,N_36095);
xnor U40431 (N_40431,N_36789,N_35040);
or U40432 (N_40432,N_35585,N_37138);
xor U40433 (N_40433,N_35646,N_37372);
nand U40434 (N_40434,N_37164,N_38122);
xor U40435 (N_40435,N_38848,N_39133);
xnor U40436 (N_40436,N_38446,N_35395);
or U40437 (N_40437,N_37821,N_37354);
nor U40438 (N_40438,N_35431,N_38711);
or U40439 (N_40439,N_39989,N_39846);
or U40440 (N_40440,N_37969,N_37398);
and U40441 (N_40441,N_35048,N_38163);
and U40442 (N_40442,N_38584,N_39785);
nand U40443 (N_40443,N_39105,N_37199);
nor U40444 (N_40444,N_36498,N_37157);
and U40445 (N_40445,N_35146,N_38998);
and U40446 (N_40446,N_39186,N_35016);
xnor U40447 (N_40447,N_36349,N_35094);
xnor U40448 (N_40448,N_35762,N_35018);
or U40449 (N_40449,N_38227,N_38133);
or U40450 (N_40450,N_39664,N_38070);
or U40451 (N_40451,N_39810,N_37563);
and U40452 (N_40452,N_35562,N_37046);
nand U40453 (N_40453,N_38719,N_38566);
and U40454 (N_40454,N_35611,N_38088);
nor U40455 (N_40455,N_37027,N_37926);
and U40456 (N_40456,N_39875,N_38952);
nand U40457 (N_40457,N_37311,N_38616);
nor U40458 (N_40458,N_37534,N_37900);
nand U40459 (N_40459,N_38345,N_38658);
nor U40460 (N_40460,N_35388,N_39449);
xor U40461 (N_40461,N_39075,N_37107);
nor U40462 (N_40462,N_36565,N_36037);
nand U40463 (N_40463,N_38795,N_35259);
nand U40464 (N_40464,N_37316,N_37375);
nor U40465 (N_40465,N_38951,N_38838);
nor U40466 (N_40466,N_39043,N_38012);
or U40467 (N_40467,N_38305,N_35916);
nor U40468 (N_40468,N_35977,N_35704);
nor U40469 (N_40469,N_36015,N_39426);
xor U40470 (N_40470,N_37128,N_37156);
xor U40471 (N_40471,N_39920,N_38499);
xnor U40472 (N_40472,N_35737,N_38081);
or U40473 (N_40473,N_38822,N_38078);
xnor U40474 (N_40474,N_39736,N_39891);
nor U40475 (N_40475,N_37834,N_39098);
nor U40476 (N_40476,N_38475,N_39106);
nand U40477 (N_40477,N_36133,N_35336);
nand U40478 (N_40478,N_35081,N_36243);
or U40479 (N_40479,N_37114,N_37024);
and U40480 (N_40480,N_38309,N_36727);
and U40481 (N_40481,N_37512,N_36617);
nor U40482 (N_40482,N_37802,N_38041);
and U40483 (N_40483,N_35408,N_39009);
nand U40484 (N_40484,N_36056,N_38016);
nor U40485 (N_40485,N_39620,N_37995);
xor U40486 (N_40486,N_36832,N_37025);
nand U40487 (N_40487,N_35211,N_36666);
nand U40488 (N_40488,N_39085,N_36032);
xnor U40489 (N_40489,N_35261,N_35055);
nor U40490 (N_40490,N_37301,N_35189);
nand U40491 (N_40491,N_39010,N_39217);
or U40492 (N_40492,N_38727,N_39971);
or U40493 (N_40493,N_38752,N_38103);
and U40494 (N_40494,N_37111,N_37121);
or U40495 (N_40495,N_38537,N_39018);
or U40496 (N_40496,N_36545,N_36533);
nand U40497 (N_40497,N_35632,N_36541);
xnor U40498 (N_40498,N_35052,N_38507);
or U40499 (N_40499,N_37436,N_39079);
nor U40500 (N_40500,N_35280,N_39338);
nand U40501 (N_40501,N_35275,N_39764);
or U40502 (N_40502,N_36483,N_37609);
nand U40503 (N_40503,N_35345,N_35460);
and U40504 (N_40504,N_35479,N_36078);
nand U40505 (N_40505,N_38028,N_36447);
nand U40506 (N_40506,N_38124,N_38135);
nand U40507 (N_40507,N_35993,N_37807);
xor U40508 (N_40508,N_39142,N_37314);
or U40509 (N_40509,N_35221,N_36696);
or U40510 (N_40510,N_38582,N_36091);
or U40511 (N_40511,N_37788,N_36156);
and U40512 (N_40512,N_36455,N_36555);
or U40513 (N_40513,N_38766,N_39511);
nand U40514 (N_40514,N_35923,N_35645);
xnor U40515 (N_40515,N_36108,N_36620);
nand U40516 (N_40516,N_39197,N_39445);
or U40517 (N_40517,N_37790,N_39893);
and U40518 (N_40518,N_36833,N_35596);
xor U40519 (N_40519,N_36818,N_38091);
nand U40520 (N_40520,N_35337,N_39708);
xor U40521 (N_40521,N_37072,N_39002);
nor U40522 (N_40522,N_36711,N_37970);
or U40523 (N_40523,N_35926,N_35863);
and U40524 (N_40524,N_36573,N_37809);
or U40525 (N_40525,N_35164,N_37923);
and U40526 (N_40526,N_37188,N_38802);
nand U40527 (N_40527,N_36504,N_36397);
xnor U40528 (N_40528,N_36785,N_35862);
xnor U40529 (N_40529,N_35630,N_38443);
and U40530 (N_40530,N_35285,N_38474);
or U40531 (N_40531,N_35380,N_39955);
or U40532 (N_40532,N_37612,N_35991);
and U40533 (N_40533,N_36866,N_35674);
xnor U40534 (N_40534,N_39400,N_38667);
or U40535 (N_40535,N_35947,N_35582);
nand U40536 (N_40536,N_38426,N_38391);
nor U40537 (N_40537,N_36551,N_39382);
nand U40538 (N_40538,N_35493,N_37231);
or U40539 (N_40539,N_37236,N_39373);
or U40540 (N_40540,N_39826,N_36906);
and U40541 (N_40541,N_35905,N_38596);
and U40542 (N_40542,N_37187,N_35506);
and U40543 (N_40543,N_37169,N_38101);
nor U40544 (N_40544,N_35071,N_38867);
or U40545 (N_40545,N_36905,N_37428);
xor U40546 (N_40546,N_38551,N_35782);
xor U40547 (N_40547,N_36285,N_37735);
nand U40548 (N_40548,N_37988,N_37985);
xor U40549 (N_40549,N_37963,N_36322);
nor U40550 (N_40550,N_38433,N_35557);
nor U40551 (N_40551,N_36299,N_36886);
nor U40552 (N_40552,N_35790,N_37960);
and U40553 (N_40553,N_39337,N_38999);
or U40554 (N_40554,N_39824,N_36406);
or U40555 (N_40555,N_35075,N_38317);
xnor U40556 (N_40556,N_39087,N_36474);
and U40557 (N_40557,N_38236,N_35311);
and U40558 (N_40558,N_37424,N_37889);
nor U40559 (N_40559,N_39593,N_36366);
or U40560 (N_40560,N_35959,N_39564);
nor U40561 (N_40561,N_37929,N_37263);
or U40562 (N_40562,N_35981,N_36619);
xor U40563 (N_40563,N_37145,N_35482);
and U40564 (N_40564,N_35486,N_35810);
nor U40565 (N_40565,N_35378,N_39510);
and U40566 (N_40566,N_35550,N_37235);
or U40567 (N_40567,N_35097,N_35678);
xnor U40568 (N_40568,N_36820,N_37814);
nand U40569 (N_40569,N_38569,N_37376);
nand U40570 (N_40570,N_38416,N_38293);
nor U40571 (N_40571,N_39545,N_35656);
or U40572 (N_40572,N_37496,N_39323);
nor U40573 (N_40573,N_37279,N_36813);
and U40574 (N_40574,N_39188,N_36855);
xor U40575 (N_40575,N_39769,N_38611);
or U40576 (N_40576,N_38258,N_36861);
or U40577 (N_40577,N_35272,N_37195);
and U40578 (N_40578,N_36284,N_38979);
nand U40579 (N_40579,N_35090,N_36852);
nor U40580 (N_40580,N_35625,N_35574);
and U40581 (N_40581,N_39863,N_37002);
nand U40582 (N_40582,N_36650,N_38583);
nor U40583 (N_40583,N_35917,N_39308);
and U40584 (N_40584,N_36996,N_36338);
or U40585 (N_40585,N_39182,N_37091);
nor U40586 (N_40586,N_36700,N_36158);
nand U40587 (N_40587,N_36459,N_38986);
and U40588 (N_40588,N_35885,N_38067);
xor U40589 (N_40589,N_39424,N_39703);
and U40590 (N_40590,N_38393,N_37585);
and U40591 (N_40591,N_35320,N_36006);
nand U40592 (N_40592,N_39437,N_39369);
or U40593 (N_40593,N_35443,N_38556);
xnor U40594 (N_40594,N_37613,N_37097);
and U40595 (N_40595,N_39784,N_37941);
or U40596 (N_40596,N_35206,N_35316);
nand U40597 (N_40597,N_38344,N_35232);
nand U40598 (N_40598,N_38448,N_37224);
and U40599 (N_40599,N_36001,N_36216);
or U40600 (N_40600,N_38462,N_35882);
nand U40601 (N_40601,N_36030,N_36041);
and U40602 (N_40602,N_38435,N_37135);
xnor U40603 (N_40603,N_35531,N_38984);
or U40604 (N_40604,N_35694,N_38061);
or U40605 (N_40605,N_38828,N_36901);
nor U40606 (N_40606,N_35374,N_38160);
xor U40607 (N_40607,N_36321,N_39936);
and U40608 (N_40608,N_36077,N_37909);
xor U40609 (N_40609,N_39549,N_38318);
and U40610 (N_40610,N_38930,N_37687);
and U40611 (N_40611,N_37957,N_37288);
and U40612 (N_40612,N_35537,N_38717);
xnor U40613 (N_40613,N_37423,N_36626);
nor U40614 (N_40614,N_37096,N_39865);
nor U40615 (N_40615,N_36058,N_37946);
xnor U40616 (N_40616,N_36561,N_38688);
or U40617 (N_40617,N_38275,N_36398);
xnor U40618 (N_40618,N_36241,N_37084);
and U40619 (N_40619,N_38935,N_35271);
or U40620 (N_40620,N_39360,N_37745);
nand U40621 (N_40621,N_39592,N_35426);
nor U40622 (N_40622,N_35935,N_39887);
and U40623 (N_40623,N_35682,N_38425);
nand U40624 (N_40624,N_36513,N_37665);
nor U40625 (N_40625,N_35089,N_35775);
nand U40626 (N_40626,N_36475,N_36422);
nor U40627 (N_40627,N_35103,N_35251);
or U40628 (N_40628,N_36673,N_36546);
and U40629 (N_40629,N_39742,N_38785);
nand U40630 (N_40630,N_38268,N_35240);
and U40631 (N_40631,N_39173,N_36157);
xor U40632 (N_40632,N_39315,N_39332);
xor U40633 (N_40633,N_37764,N_38481);
nand U40634 (N_40634,N_39656,N_39314);
or U40635 (N_40635,N_38276,N_38399);
xnor U40636 (N_40636,N_36212,N_38649);
and U40637 (N_40637,N_35070,N_38562);
and U40638 (N_40638,N_36246,N_37862);
or U40639 (N_40639,N_35843,N_35672);
xnor U40640 (N_40640,N_35208,N_36910);
nand U40641 (N_40641,N_38919,N_37775);
or U40642 (N_40642,N_38906,N_38958);
and U40643 (N_40643,N_36680,N_36840);
and U40644 (N_40644,N_37859,N_38778);
nor U40645 (N_40645,N_38167,N_35913);
xnor U40646 (N_40646,N_37656,N_38613);
or U40647 (N_40647,N_38228,N_39107);
and U40648 (N_40648,N_39697,N_39808);
nand U40649 (N_40649,N_38455,N_37881);
xor U40650 (N_40650,N_36869,N_38776);
nand U40651 (N_40651,N_36601,N_35735);
nand U40652 (N_40652,N_38505,N_36857);
nand U40653 (N_40653,N_37435,N_38780);
or U40654 (N_40654,N_36274,N_36490);
and U40655 (N_40655,N_36256,N_35787);
xnor U40656 (N_40656,N_37074,N_39751);
and U40657 (N_40657,N_37702,N_39329);
nand U40658 (N_40658,N_35148,N_35014);
xor U40659 (N_40659,N_35541,N_36421);
and U40660 (N_40660,N_36332,N_36767);
xnor U40661 (N_40661,N_38622,N_38080);
xnor U40662 (N_40662,N_39080,N_36401);
or U40663 (N_40663,N_37402,N_36106);
nor U40664 (N_40664,N_37694,N_36134);
xnor U40665 (N_40665,N_38547,N_39398);
xnor U40666 (N_40666,N_39925,N_37732);
nor U40667 (N_40667,N_37447,N_39555);
xnor U40668 (N_40668,N_36876,N_39290);
or U40669 (N_40669,N_39687,N_35591);
nand U40670 (N_40670,N_37832,N_37891);
or U40671 (N_40671,N_36704,N_35481);
xor U40672 (N_40672,N_39880,N_38115);
nand U40673 (N_40673,N_37008,N_38301);
nor U40674 (N_40674,N_38697,N_38402);
nand U40675 (N_40675,N_36796,N_36279);
xnor U40676 (N_40676,N_39832,N_39730);
xor U40677 (N_40677,N_36965,N_36525);
nand U40678 (N_40678,N_38262,N_39179);
nor U40679 (N_40679,N_36065,N_36000);
nor U40680 (N_40680,N_38171,N_36247);
nand U40681 (N_40681,N_37464,N_39960);
and U40682 (N_40682,N_35159,N_35087);
and U40683 (N_40683,N_39014,N_35857);
nand U40684 (N_40684,N_37384,N_35376);
xor U40685 (N_40685,N_39858,N_38001);
xor U40686 (N_40686,N_36117,N_39479);
or U40687 (N_40687,N_36948,N_36774);
and U40688 (N_40688,N_35429,N_36370);
xnor U40689 (N_40689,N_35085,N_38968);
and U40690 (N_40690,N_36233,N_35007);
or U40691 (N_40691,N_37825,N_38176);
xnor U40692 (N_40692,N_37573,N_36538);
xnor U40693 (N_40693,N_37796,N_39048);
nor U40694 (N_40694,N_38297,N_37054);
xor U40695 (N_40695,N_36713,N_39906);
xor U40696 (N_40696,N_36733,N_38605);
xor U40697 (N_40697,N_38273,N_37660);
xor U40698 (N_40698,N_37591,N_37466);
or U40699 (N_40699,N_35158,N_37935);
nor U40700 (N_40700,N_37256,N_39240);
or U40701 (N_40701,N_38024,N_36740);
nand U40702 (N_40702,N_37259,N_38029);
and U40703 (N_40703,N_35548,N_39516);
xnor U40704 (N_40704,N_39326,N_35195);
nand U40705 (N_40705,N_36265,N_39128);
and U40706 (N_40706,N_38517,N_36008);
and U40707 (N_40707,N_39198,N_36145);
xor U40708 (N_40708,N_36384,N_39980);
xnor U40709 (N_40709,N_37218,N_36506);
and U40710 (N_40710,N_35235,N_36940);
or U40711 (N_40711,N_38445,N_37548);
nor U40712 (N_40712,N_35887,N_37110);
nor U40713 (N_40713,N_35204,N_36655);
nand U40714 (N_40714,N_37439,N_36979);
or U40715 (N_40715,N_36648,N_38213);
and U40716 (N_40716,N_36023,N_37737);
nand U40717 (N_40717,N_35928,N_36983);
nand U40718 (N_40718,N_36179,N_36729);
nor U40719 (N_40719,N_38050,N_38398);
and U40720 (N_40720,N_39756,N_35392);
nand U40721 (N_40721,N_35169,N_35241);
xnor U40722 (N_40722,N_35401,N_38981);
and U40723 (N_40723,N_39854,N_35010);
nor U40724 (N_40724,N_35581,N_37456);
xor U40725 (N_40725,N_35805,N_39377);
and U40726 (N_40726,N_37086,N_38165);
nor U40727 (N_40727,N_36099,N_39860);
or U40728 (N_40728,N_36588,N_35579);
nand U40729 (N_40729,N_37123,N_39391);
and U40730 (N_40730,N_39707,N_37475);
xnor U40731 (N_40731,N_35939,N_37927);
nor U40732 (N_40732,N_38137,N_38243);
nand U40733 (N_40733,N_38117,N_38577);
nand U40734 (N_40734,N_39318,N_36497);
and U40735 (N_40735,N_37215,N_38554);
xor U40736 (N_40736,N_35622,N_39493);
xor U40737 (N_40737,N_35440,N_35697);
nand U40738 (N_40738,N_38205,N_39203);
xor U40739 (N_40739,N_35745,N_37211);
or U40740 (N_40740,N_35650,N_39926);
or U40741 (N_40741,N_36154,N_38877);
nor U40742 (N_40742,N_39551,N_38185);
nand U40743 (N_40743,N_39174,N_39669);
or U40744 (N_40744,N_35588,N_36709);
nor U40745 (N_40745,N_35621,N_39317);
nand U40746 (N_40746,N_38052,N_37416);
nor U40747 (N_40747,N_37741,N_36103);
nor U40748 (N_40748,N_39541,N_37058);
nor U40749 (N_40749,N_37321,N_36364);
nand U40750 (N_40750,N_36132,N_35614);
nor U40751 (N_40751,N_35141,N_37914);
and U40752 (N_40752,N_36162,N_35710);
xnor U40753 (N_40753,N_36702,N_37925);
xor U40754 (N_40754,N_39594,N_36304);
nor U40755 (N_40755,N_37551,N_35602);
or U40756 (N_40756,N_39877,N_35281);
nand U40757 (N_40757,N_35750,N_36136);
nand U40758 (N_40758,N_38610,N_38510);
nor U40759 (N_40759,N_35587,N_37761);
nand U40760 (N_40760,N_36381,N_35865);
and U40761 (N_40761,N_37977,N_37966);
nand U40762 (N_40762,N_36514,N_36269);
nor U40763 (N_40763,N_35462,N_36543);
nand U40764 (N_40764,N_38978,N_39929);
nand U40765 (N_40765,N_35864,N_37294);
and U40766 (N_40766,N_37524,N_38833);
nor U40767 (N_40767,N_39853,N_39038);
xnor U40768 (N_40768,N_37191,N_35284);
nor U40769 (N_40769,N_38363,N_39178);
or U40770 (N_40770,N_39216,N_35856);
nor U40771 (N_40771,N_37403,N_35779);
nor U40772 (N_40772,N_39902,N_39956);
or U40773 (N_40773,N_38498,N_38209);
xor U40774 (N_40774,N_39570,N_36378);
nor U40775 (N_40775,N_35494,N_36891);
or U40776 (N_40776,N_38442,N_38136);
and U40777 (N_40777,N_38234,N_36125);
nand U40778 (N_40778,N_36347,N_37848);
and U40779 (N_40779,N_35613,N_36043);
and U40780 (N_40780,N_39856,N_38893);
nor U40781 (N_40781,N_36577,N_35641);
xnor U40782 (N_40782,N_39806,N_38032);
or U40783 (N_40783,N_39998,N_35296);
nand U40784 (N_40784,N_38821,N_38757);
xor U40785 (N_40785,N_35594,N_35970);
and U40786 (N_40786,N_38746,N_39302);
nand U40787 (N_40787,N_37677,N_37352);
xnor U40788 (N_40788,N_36834,N_37134);
or U40789 (N_40789,N_39721,N_36511);
nor U40790 (N_40790,N_39968,N_39950);
xnor U40791 (N_40791,N_36749,N_39187);
xor U40792 (N_40792,N_36149,N_39840);
nor U40793 (N_40793,N_37359,N_35438);
nand U40794 (N_40794,N_37201,N_38870);
and U40795 (N_40795,N_35334,N_36087);
or U40796 (N_40796,N_37720,N_39269);
or U40797 (N_40797,N_39239,N_35365);
xor U40798 (N_40798,N_38980,N_37588);
or U40799 (N_40799,N_39964,N_35877);
or U40800 (N_40800,N_35609,N_38015);
nor U40801 (N_40801,N_35505,N_35549);
xnor U40802 (N_40802,N_37394,N_36139);
nand U40803 (N_40803,N_38249,N_38406);
nor U40804 (N_40804,N_38595,N_35936);
and U40805 (N_40805,N_36519,N_37887);
xnor U40806 (N_40806,N_35002,N_38858);
nand U40807 (N_40807,N_38885,N_35796);
nand U40808 (N_40808,N_38698,N_37753);
or U40809 (N_40809,N_37013,N_36674);
and U40810 (N_40810,N_39470,N_39192);
xnor U40811 (N_40811,N_38575,N_38279);
nor U40812 (N_40812,N_38729,N_35104);
nor U40813 (N_40813,N_35638,N_36678);
or U40814 (N_40814,N_35278,N_36580);
nor U40815 (N_40815,N_35260,N_39945);
nand U40816 (N_40816,N_36522,N_37522);
nor U40817 (N_40817,N_39548,N_35471);
nor U40818 (N_40818,N_38287,N_36574);
or U40819 (N_40819,N_36271,N_37329);
nand U40820 (N_40820,N_36772,N_38329);
nand U40821 (N_40821,N_36836,N_36760);
xnor U40822 (N_40822,N_36476,N_36801);
or U40823 (N_40823,N_39375,N_36425);
nand U40824 (N_40824,N_39508,N_37385);
and U40825 (N_40825,N_38767,N_35328);
nor U40826 (N_40826,N_37019,N_36244);
nor U40827 (N_40827,N_38748,N_35845);
or U40828 (N_40828,N_36851,N_35473);
and U40829 (N_40829,N_36732,N_37710);
xor U40830 (N_40830,N_35490,N_38480);
xor U40831 (N_40831,N_35215,N_36405);
and U40832 (N_40832,N_38721,N_36427);
or U40833 (N_40833,N_35053,N_36485);
nand U40834 (N_40834,N_37172,N_37682);
xor U40835 (N_40835,N_38572,N_39047);
and U40836 (N_40836,N_38501,N_35755);
and U40837 (N_40837,N_38149,N_35722);
and U40838 (N_40838,N_35597,N_35988);
or U40839 (N_40839,N_35707,N_37030);
nand U40840 (N_40840,N_39066,N_36646);
nand U40841 (N_40841,N_37912,N_35804);
nand U40842 (N_40842,N_38197,N_37607);
nand U40843 (N_40843,N_38512,N_36377);
or U40844 (N_40844,N_39169,N_38843);
and U40845 (N_40845,N_37680,N_39717);
nand U40846 (N_40846,N_37080,N_36309);
or U40847 (N_40847,N_39357,N_39786);
or U40848 (N_40848,N_39948,N_39032);
xor U40849 (N_40849,N_35852,N_36977);
xor U40850 (N_40850,N_36571,N_35600);
and U40851 (N_40851,N_36168,N_38166);
nor U40852 (N_40852,N_39224,N_39309);
and U40853 (N_40853,N_38479,N_39140);
xor U40854 (N_40854,N_38788,N_39678);
or U40855 (N_40855,N_39255,N_39673);
xor U40856 (N_40856,N_39850,N_35015);
or U40857 (N_40857,N_36941,N_36187);
nand U40858 (N_40858,N_37815,N_38201);
xnor U40859 (N_40859,N_36210,N_39193);
and U40860 (N_40860,N_36639,N_36142);
and U40861 (N_40861,N_38905,N_35212);
and U40862 (N_40862,N_38030,N_38769);
nor U40863 (N_40863,N_35802,N_39864);
or U40864 (N_40864,N_39341,N_35180);
xnor U40865 (N_40865,N_39642,N_37953);
nor U40866 (N_40866,N_35341,N_38689);
nand U40867 (N_40867,N_35784,N_35967);
nand U40868 (N_40868,N_37389,N_37366);
xnor U40869 (N_40869,N_38362,N_39367);
and U40870 (N_40870,N_38368,N_39243);
nor U40871 (N_40871,N_37387,N_35530);
nor U40872 (N_40872,N_38553,N_37222);
xnor U40873 (N_40873,N_36159,N_35023);
xor U40874 (N_40874,N_36824,N_35721);
nor U40875 (N_40875,N_36564,N_38497);
or U40876 (N_40876,N_37818,N_38260);
xnor U40877 (N_40877,N_37707,N_39696);
nand U40878 (N_40878,N_38096,N_35829);
nand U40879 (N_40879,N_38051,N_35700);
nor U40880 (N_40880,N_37196,N_37558);
xor U40881 (N_40881,N_37968,N_35749);
and U40882 (N_40882,N_37523,N_37453);
and U40883 (N_40883,N_36471,N_35934);
nand U40884 (N_40884,N_39139,N_35734);
xor U40885 (N_40885,N_39108,N_37568);
or U40886 (N_40886,N_35116,N_39206);
xnor U40887 (N_40887,N_35999,N_37532);
or U40888 (N_40888,N_38774,N_37876);
xnor U40889 (N_40889,N_35517,N_36350);
and U40890 (N_40890,N_38601,N_35754);
nand U40891 (N_40891,N_38394,N_37364);
xnor U40892 (N_40892,N_38155,N_39246);
nor U40893 (N_40893,N_37998,N_36899);
or U40894 (N_40894,N_36192,N_37465);
nor U40895 (N_40895,N_39407,N_38397);
and U40896 (N_40896,N_38369,N_35405);
xnor U40897 (N_40897,N_38761,N_39170);
or U40898 (N_40898,N_38738,N_36980);
nand U40899 (N_40899,N_37248,N_36211);
xnor U40900 (N_40900,N_39694,N_38751);
and U40901 (N_40901,N_37395,N_38266);
or U40902 (N_40902,N_36718,N_39316);
nand U40903 (N_40903,N_37407,N_38589);
or U40904 (N_40904,N_39328,N_39641);
nor U40905 (N_40905,N_39130,N_36627);
nand U40906 (N_40906,N_39233,N_38247);
nor U40907 (N_40907,N_39024,N_35969);
and U40908 (N_40908,N_37885,N_35302);
xnor U40909 (N_40909,N_36387,N_37717);
and U40910 (N_40910,N_37487,N_38272);
nand U40911 (N_40911,N_38413,N_37993);
nor U40912 (N_40912,N_38705,N_38712);
nor U40913 (N_40913,N_39529,N_36638);
nand U40914 (N_40914,N_37742,N_39430);
and U40915 (N_40915,N_37669,N_38087);
xor U40916 (N_40916,N_37615,N_38742);
nand U40917 (N_40917,N_36467,N_38259);
nor U40918 (N_40918,N_37509,N_39078);
nand U40919 (N_40919,N_36903,N_37997);
nand U40920 (N_40920,N_36955,N_37443);
xor U40921 (N_40921,N_36379,N_36584);
nand U40922 (N_40922,N_36736,N_39253);
and U40923 (N_40923,N_36107,N_36606);
xnor U40924 (N_40924,N_36297,N_35179);
xnor U40925 (N_40925,N_37056,N_39713);
nand U40926 (N_40926,N_36893,N_37671);
and U40927 (N_40927,N_37833,N_38955);
nor U40928 (N_40928,N_39624,N_35228);
xor U40929 (N_40929,N_36808,N_35813);
nand U40930 (N_40930,N_38849,N_35113);
nand U40931 (N_40931,N_36815,N_37763);
xnor U40932 (N_40932,N_36679,N_37819);
or U40933 (N_40933,N_39399,N_35276);
or U40934 (N_40934,N_36437,N_37785);
nand U40935 (N_40935,N_39645,N_37630);
or U40936 (N_40936,N_37538,N_39452);
xor U40937 (N_40937,N_35624,N_37146);
nor U40938 (N_40938,N_35685,N_35789);
xnor U40939 (N_40939,N_37899,N_37644);
and U40940 (N_40940,N_35382,N_36604);
xor U40941 (N_40941,N_38330,N_35751);
nor U40942 (N_40942,N_39409,N_39978);
nor U40943 (N_40943,N_36330,N_36976);
nor U40944 (N_40944,N_37127,N_38741);
xor U40945 (N_40945,N_35270,N_39755);
or U40946 (N_40946,N_39911,N_37063);
nand U40947 (N_40947,N_35063,N_37154);
nor U40948 (N_40948,N_39042,N_39325);
xnor U40949 (N_40949,N_35435,N_38141);
nand U40950 (N_40950,N_38040,N_36383);
xor U40951 (N_40951,N_39237,N_36590);
xor U40952 (N_40952,N_36887,N_39125);
or U40953 (N_40953,N_35914,N_35287);
xor U40954 (N_40954,N_37064,N_36957);
nand U40955 (N_40955,N_39468,N_35781);
nand U40956 (N_40956,N_36994,N_36426);
xor U40957 (N_40957,N_39595,N_38811);
or U40958 (N_40958,N_36971,N_36634);
nor U40959 (N_40959,N_36797,N_36641);
or U40960 (N_40960,N_37769,N_39421);
and U40961 (N_40961,N_39847,N_35996);
nor U40962 (N_40962,N_37964,N_37893);
nor U40963 (N_40963,N_38037,N_36724);
and U40964 (N_40964,N_38371,N_35367);
and U40965 (N_40965,N_39274,N_36487);
or U40966 (N_40966,N_36578,N_39259);
and U40967 (N_40967,N_36080,N_37347);
and U40968 (N_40968,N_36799,N_38323);
and U40969 (N_40969,N_35310,N_36877);
or U40970 (N_40970,N_39280,N_35256);
xor U40971 (N_40971,N_36645,N_39588);
nand U40972 (N_40972,N_38189,N_36266);
xnor U40973 (N_40973,N_39793,N_36324);
or U40974 (N_40974,N_35900,N_36624);
xor U40975 (N_40975,N_37283,N_39138);
and U40976 (N_40976,N_38354,N_36165);
nor U40977 (N_40977,N_36486,N_38286);
nand U40978 (N_40978,N_35076,N_36218);
or U40979 (N_40979,N_39732,N_36722);
xor U40980 (N_40980,N_39181,N_37850);
nor U40981 (N_40981,N_38875,N_38696);
and U40982 (N_40982,N_38660,N_36978);
and U40983 (N_40983,N_39540,N_35188);
or U40984 (N_40984,N_35379,N_39524);
nand U40985 (N_40985,N_35767,N_38678);
xor U40986 (N_40986,N_39630,N_39718);
or U40987 (N_40987,N_38451,N_37181);
xor U40988 (N_40988,N_39070,N_38871);
xor U40989 (N_40989,N_38492,N_35442);
and U40990 (N_40990,N_35346,N_39567);
nor U40991 (N_40991,N_35009,N_39970);
nand U40992 (N_40992,N_35839,N_36390);
nand U40993 (N_40993,N_37978,N_36263);
or U40994 (N_40994,N_35949,N_35944);
nor U40995 (N_40995,N_36440,N_35216);
nor U40996 (N_40996,N_39918,N_38405);
xnor U40997 (N_40997,N_37636,N_39111);
nor U40998 (N_40998,N_38627,N_37043);
nand U40999 (N_40999,N_36391,N_36549);
nand U41000 (N_41000,N_35724,N_36780);
nand U41001 (N_41001,N_38956,N_36205);
or U41002 (N_41002,N_37601,N_39770);
or U41003 (N_41003,N_36874,N_37693);
xor U41004 (N_41004,N_35976,N_38342);
or U41005 (N_41005,N_38954,N_37438);
nand U41006 (N_41006,N_37672,N_38618);
and U41007 (N_41007,N_38829,N_38277);
or U41008 (N_41008,N_39094,N_37781);
xnor U41009 (N_41009,N_38146,N_39158);
and U41010 (N_41010,N_35821,N_39082);
or U41011 (N_41011,N_36166,N_36493);
and U41012 (N_41012,N_39794,N_36123);
nor U41013 (N_41013,N_35129,N_36220);
or U41014 (N_41014,N_36281,N_37996);
nor U41015 (N_41015,N_36457,N_36991);
and U41016 (N_41016,N_36598,N_39626);
nor U41017 (N_41017,N_36697,N_35518);
nor U41018 (N_41018,N_38552,N_35635);
xnor U41019 (N_41019,N_39175,N_36879);
or U41020 (N_41020,N_38997,N_35006);
nor U41021 (N_41021,N_37625,N_38059);
xnor U41022 (N_41022,N_37400,N_35037);
nand U41023 (N_41023,N_38509,N_36214);
nand U41024 (N_41024,N_36028,N_36326);
nor U41025 (N_41025,N_38617,N_38869);
or U41026 (N_41026,N_37417,N_39347);
nor U41027 (N_41027,N_39829,N_38453);
or U41028 (N_41028,N_37026,N_36520);
nand U41029 (N_41029,N_38646,N_37906);
nand U41030 (N_41030,N_39519,N_36311);
nor U41031 (N_41031,N_37304,N_35592);
xnor U41032 (N_41032,N_35715,N_38545);
or U41033 (N_41033,N_39113,N_38500);
xnor U41034 (N_41034,N_38218,N_39924);
xnor U41035 (N_41035,N_36842,N_39580);
xor U41036 (N_41036,N_39882,N_37543);
or U41037 (N_41037,N_37840,N_38068);
nand U41038 (N_41038,N_38341,N_35249);
xor U41039 (N_41039,N_39589,N_39542);
xnor U41040 (N_41040,N_38456,N_37746);
xor U41041 (N_41041,N_39053,N_38539);
or U41042 (N_41042,N_37539,N_37162);
nand U41043 (N_41043,N_38250,N_38520);
or U41044 (N_41044,N_36612,N_38332);
nand U41045 (N_41045,N_36365,N_36495);
or U41046 (N_41046,N_38430,N_36275);
and U41047 (N_41047,N_36100,N_38106);
and U41048 (N_41048,N_38673,N_36382);
or U41049 (N_41049,N_38111,N_39915);
xor U41050 (N_41050,N_36615,N_37765);
xnor U41051 (N_41051,N_35833,N_39571);
or U41052 (N_41052,N_37031,N_38704);
nand U41053 (N_41053,N_37980,N_35332);
nand U41054 (N_41054,N_35024,N_37569);
or U41055 (N_41055,N_37167,N_37994);
nor U41056 (N_41056,N_38288,N_37674);
or U41057 (N_41057,N_37185,N_37842);
and U41058 (N_41058,N_35417,N_36039);
nand U41059 (N_41059,N_39818,N_37050);
nand U41060 (N_41060,N_39057,N_39483);
or U41061 (N_41061,N_38380,N_39026);
nor U41062 (N_41062,N_39453,N_38789);
xor U41063 (N_41063,N_36097,N_37100);
xor U41064 (N_41064,N_37401,N_37328);
and U41065 (N_41065,N_38644,N_36310);
or U41066 (N_41066,N_38503,N_36897);
or U41067 (N_41067,N_36372,N_38578);
xor U41068 (N_41068,N_36657,N_38409);
or U41069 (N_41069,N_35499,N_35068);
nor U41070 (N_41070,N_35119,N_36853);
and U41071 (N_41071,N_38003,N_39168);
and U41072 (N_41072,N_37441,N_38528);
or U41073 (N_41073,N_39037,N_37755);
xor U41074 (N_41074,N_37549,N_39648);
nand U41075 (N_41075,N_37371,N_39352);
nor U41076 (N_41076,N_39934,N_38370);
or U41077 (N_41077,N_35277,N_39659);
xor U41078 (N_41078,N_39581,N_35453);
nor U41079 (N_41079,N_36408,N_39735);
nand U41080 (N_41080,N_35044,N_36312);
xor U41081 (N_41081,N_38772,N_35844);
nand U41082 (N_41082,N_35439,N_35569);
or U41083 (N_41083,N_38929,N_37951);
xnor U41084 (N_41084,N_36867,N_37771);
nand U41085 (N_41085,N_38850,N_35607);
and U41086 (N_41086,N_36635,N_38245);
nand U41087 (N_41087,N_39531,N_39141);
nor U41088 (N_41088,N_35357,N_36395);
xor U41089 (N_41089,N_37446,N_36936);
nor U41090 (N_41090,N_35793,N_37689);
nand U41091 (N_41091,N_38265,N_38608);
or U41092 (N_41092,N_38876,N_37638);
or U41093 (N_41093,N_35637,N_36914);
nand U41094 (N_41094,N_39940,N_38312);
xnor U41095 (N_41095,N_36703,N_39783);
or U41096 (N_41096,N_38056,N_37153);
xnor U41097 (N_41097,N_37602,N_35197);
nand U41098 (N_41098,N_37839,N_36195);
and U41099 (N_41099,N_37703,N_37061);
nand U41100 (N_41100,N_37567,N_35340);
and U41101 (N_41101,N_36787,N_36161);
xnor U41102 (N_41102,N_37553,N_37374);
nand U41103 (N_41103,N_36741,N_36292);
xnor U41104 (N_41104,N_36597,N_39268);
and U41105 (N_41105,N_35527,N_37356);
and U41106 (N_41106,N_39932,N_39698);
nand U41107 (N_41107,N_39914,N_38240);
or U41108 (N_41108,N_38374,N_35160);
xnor U41109 (N_41109,N_35803,N_35151);
and U41110 (N_41110,N_38634,N_37479);
nor U41111 (N_41111,N_35163,N_38089);
nor U41112 (N_41112,N_39723,N_39753);
or U41113 (N_41113,N_38643,N_39097);
and U41114 (N_41114,N_36961,N_39395);
nand U41115 (N_41115,N_36800,N_39905);
nand U41116 (N_41116,N_39901,N_36454);
or U41117 (N_41117,N_37223,N_36517);
nand U41118 (N_41118,N_39127,N_36066);
nor U41119 (N_41119,N_39194,N_38834);
and U41120 (N_41120,N_38321,N_38591);
nor U41121 (N_41121,N_37786,N_39362);
or U41122 (N_41122,N_36660,N_39720);
nand U41123 (N_41123,N_36542,N_37948);
nand U41124 (N_41124,N_35099,N_39797);
or U41125 (N_41125,N_35318,N_38847);
nor U41126 (N_41126,N_39313,N_36822);
nand U41127 (N_41127,N_36081,N_38879);
xnor U41128 (N_41128,N_37333,N_37698);
and U41129 (N_41129,N_36050,N_37075);
nand U41130 (N_41130,N_39161,N_37132);
xnor U41131 (N_41131,N_38560,N_35147);
and U41132 (N_41132,N_36942,N_35133);
nor U41133 (N_41133,N_36316,N_35872);
or U41134 (N_41134,N_39658,N_38222);
nor U41135 (N_41135,N_35107,N_36862);
and U41136 (N_41136,N_36562,N_39886);
or U41137 (N_41137,N_38800,N_36301);
nand U41138 (N_41138,N_38147,N_39384);
or U41139 (N_41139,N_35880,N_35540);
nor U41140 (N_41140,N_36764,N_38361);
xnor U41141 (N_41141,N_35626,N_36462);
nand U41142 (N_41142,N_38856,N_35056);
nand U41143 (N_41143,N_36386,N_39215);
nand U41144 (N_41144,N_37990,N_38328);
xor U41145 (N_41145,N_39927,N_38633);
nand U41146 (N_41146,N_38077,N_37592);
or U41147 (N_41147,N_37619,N_39652);
nand U41148 (N_41148,N_36927,N_37237);
and U41149 (N_41149,N_36083,N_35041);
nor U41150 (N_41150,N_39069,N_36276);
nor U41151 (N_41151,N_38677,N_39404);
xor U41152 (N_41152,N_36409,N_38593);
and U41153 (N_41153,N_35954,N_36585);
and U41154 (N_41154,N_35265,N_39688);
or U41155 (N_41155,N_36082,N_38017);
nand U41156 (N_41156,N_38747,N_38473);
or U41157 (N_41157,N_36116,N_35459);
or U41158 (N_41158,N_38777,N_39878);
and U41159 (N_41159,N_37016,N_38959);
nand U41160 (N_41160,N_35576,N_35299);
xnor U41161 (N_41161,N_35647,N_35124);
nand U41162 (N_41162,N_35911,N_39475);
and U41163 (N_41163,N_35411,N_36838);
nor U41164 (N_41164,N_36669,N_39061);
nand U41165 (N_41165,N_35218,N_38190);
nand U41166 (N_41166,N_39897,N_37823);
nor U41167 (N_41167,N_38387,N_37860);
xnor U41168 (N_41168,N_36024,N_39798);
and U41169 (N_41169,N_35161,N_39543);
xor U41170 (N_41170,N_38226,N_37506);
or U41171 (N_41171,N_38267,N_36170);
or U41172 (N_41172,N_38683,N_35670);
and U41173 (N_41173,N_38599,N_38527);
and U41174 (N_41174,N_37291,N_38702);
xnor U41175 (N_41175,N_39232,N_37353);
and U41176 (N_41176,N_38389,N_37944);
nor U41177 (N_41177,N_38631,N_36515);
or U41178 (N_41178,N_35894,N_35470);
or U41179 (N_41179,N_36111,N_38506);
nor U41180 (N_41180,N_35875,N_39298);
nand U41181 (N_41181,N_35633,N_37318);
nand U41182 (N_41182,N_37820,N_38134);
xnor U41183 (N_41183,N_38518,N_36190);
nor U41184 (N_41184,N_35168,N_38514);
and U41185 (N_41185,N_38726,N_39734);
or U41186 (N_41186,N_39119,N_38563);
nand U41187 (N_41187,N_39561,N_36750);
nor U41188 (N_41188,N_37991,N_39534);
nor U41189 (N_41189,N_39584,N_37972);
xnor U41190 (N_41190,N_35945,N_38783);
nor U41191 (N_41191,N_36200,N_36967);
xor U41192 (N_41192,N_37734,N_37736);
nor U41193 (N_41193,N_37989,N_37310);
nor U41194 (N_41194,N_35664,N_39312);
and U41195 (N_41195,N_39211,N_39355);
nand U41196 (N_41196,N_37175,N_35289);
and U41197 (N_41197,N_39896,N_37992);
xnor U41198 (N_41198,N_39984,N_39749);
and U41199 (N_41199,N_36622,N_36203);
nor U41200 (N_41200,N_37883,N_39006);
or U41201 (N_41201,N_35729,N_38880);
nor U41202 (N_41202,N_37557,N_35326);
xnor U41203 (N_41203,N_37178,N_37062);
xor U41204 (N_41204,N_39062,N_35673);
and U41205 (N_41205,N_39817,N_35776);
and U41206 (N_41206,N_35848,N_39136);
and U41207 (N_41207,N_37429,N_36027);
xor U41208 (N_41208,N_37870,N_36946);
nand U41209 (N_41209,N_36186,N_35250);
or U41210 (N_41210,N_39746,N_39771);
nand U41211 (N_41211,N_37343,N_37009);
xor U41212 (N_41212,N_39979,N_36790);
nand U41213 (N_41213,N_35717,N_37663);
xnor U41214 (N_41214,N_39469,N_35542);
xnor U41215 (N_41215,N_36907,N_35134);
or U41216 (N_41216,N_36628,N_39306);
and U41217 (N_41217,N_36989,N_39933);
nor U41218 (N_41218,N_35768,N_38119);
xor U41219 (N_41219,N_39311,N_38988);
and U41220 (N_41220,N_35983,N_35409);
xor U41221 (N_41221,N_37209,N_39371);
and U41222 (N_41222,N_37262,N_35832);
nor U41223 (N_41223,N_36295,N_37106);
nor U41224 (N_41224,N_36223,N_35372);
or U41225 (N_41225,N_36226,N_37936);
xnor U41226 (N_41226,N_37149,N_39952);
xnor U41227 (N_41227,N_38977,N_36553);
nor U41228 (N_41228,N_35677,N_36119);
nor U41229 (N_41229,N_38069,N_36925);
nor U41230 (N_41230,N_38478,N_38220);
nand U41231 (N_41231,N_35660,N_38125);
and U41232 (N_41232,N_38916,N_38105);
or U41233 (N_41233,N_37622,N_37628);
or U41234 (N_41234,N_38692,N_39167);
and U41235 (N_41235,N_39045,N_38561);
nor U41236 (N_41236,N_36092,N_37618);
nand U41237 (N_41237,N_35112,N_39319);
nor U41238 (N_41238,N_39135,N_39986);
nor U41239 (N_41239,N_36053,N_38289);
or U41240 (N_41240,N_38365,N_38739);
and U41241 (N_41241,N_39739,N_37907);
and U41242 (N_41242,N_35317,N_36194);
and U41243 (N_41243,N_38549,N_38685);
xnor U41244 (N_41244,N_39862,N_35838);
nand U41245 (N_41245,N_37700,N_38202);
or U41246 (N_41246,N_38304,N_38784);
nor U41247 (N_41247,N_38367,N_37495);
xnor U41248 (N_41248,N_37102,N_39485);
nor U41249 (N_41249,N_36705,N_35989);
nand U41250 (N_41250,N_39356,N_36094);
nand U41251 (N_41251,N_37878,N_37239);
and U41252 (N_41252,N_37684,N_37695);
xnor U41253 (N_41253,N_36375,N_36456);
nand U41254 (N_41254,N_37460,N_35364);
nor U41255 (N_41255,N_39517,N_37312);
or U41256 (N_41256,N_39288,N_37874);
or U41257 (N_41257,N_39873,N_37803);
xor U41258 (N_41258,N_37647,N_37606);
xor U41259 (N_41259,N_37937,N_39155);
and U41260 (N_41260,N_38099,N_38571);
nor U41261 (N_41261,N_35503,N_37752);
nand U41262 (N_41262,N_35122,N_35962);
and U41263 (N_41263,N_35363,N_37320);
nand U41264 (N_41264,N_38014,N_37377);
and U41265 (N_41265,N_35723,N_35816);
xor U41266 (N_41266,N_38860,N_35106);
nand U41267 (N_41267,N_38060,N_37494);
or U41268 (N_41268,N_35186,N_38891);
nand U41269 (N_41269,N_37105,N_35452);
and U41270 (N_41270,N_37651,N_35763);
nand U41271 (N_41271,N_37254,N_38114);
xor U41272 (N_41272,N_36872,N_37227);
nor U41273 (N_41273,N_35393,N_35248);
nor U41274 (N_41274,N_35091,N_37962);
or U41275 (N_41275,N_36331,N_35780);
and U41276 (N_41276,N_39804,N_35940);
xnor U41277 (N_41277,N_39408,N_37661);
or U41278 (N_41278,N_36548,N_38917);
nor U41279 (N_41279,N_35269,N_37133);
and U41280 (N_41280,N_37578,N_38428);
or U41281 (N_41281,N_39358,N_37552);
nor U41282 (N_41282,N_38004,N_38144);
nand U41283 (N_41283,N_36415,N_39604);
xor U41284 (N_41284,N_35026,N_35410);
xor U41285 (N_41285,N_39463,N_37841);
and U41286 (N_41286,N_37369,N_37961);
nand U41287 (N_41287,N_36010,N_38225);
nor U41288 (N_41288,N_35963,N_38248);
nand U41289 (N_41289,N_36319,N_36521);
nand U41290 (N_41290,N_36478,N_36668);
xnor U41291 (N_41291,N_37729,N_38844);
or U41292 (N_41292,N_36607,N_35013);
xor U41293 (N_41293,N_38109,N_39039);
xnor U41294 (N_41294,N_35861,N_36250);
or U41295 (N_41295,N_38093,N_35131);
xor U41296 (N_41296,N_37866,N_36990);
nor U41297 (N_41297,N_37350,N_38680);
nor U41298 (N_41298,N_38693,N_39544);
and U41299 (N_41299,N_35595,N_39715);
nor U41300 (N_41300,N_38656,N_39722);
nand U41301 (N_41301,N_38945,N_36354);
or U41302 (N_41302,N_35980,N_37852);
and U41303 (N_41303,N_35000,N_37620);
nand U41304 (N_41304,N_38256,N_37434);
xor U41305 (N_41305,N_36021,N_37722);
or U41306 (N_41306,N_37070,N_36206);
nor U41307 (N_41307,N_39207,N_36637);
nand U41308 (N_41308,N_38944,N_38034);
nand U41309 (N_41309,N_38604,N_35110);
xor U41310 (N_41310,N_37750,N_37791);
xnor U41311 (N_41311,N_39036,N_39144);
xor U41312 (N_41312,N_39442,N_38920);
nand U41313 (N_41313,N_39020,N_39613);
nand U41314 (N_41314,N_36667,N_35551);
nor U41315 (N_41315,N_35909,N_36544);
nand U41316 (N_41316,N_37171,N_37073);
and U41317 (N_41317,N_35644,N_36062);
or U41318 (N_41318,N_36138,N_36960);
xor U41319 (N_41319,N_35227,N_35102);
nor U41320 (N_41320,N_35012,N_37846);
nor U41321 (N_41321,N_35876,N_38508);
xnor U41322 (N_41322,N_35474,N_39741);
and U41323 (N_41323,N_37829,N_35461);
xor U41324 (N_41324,N_37766,N_39916);
nand U41325 (N_41325,N_39912,N_37234);
xnor U41326 (N_41326,N_35344,N_37001);
nand U41327 (N_41327,N_37330,N_36463);
or U41328 (N_41328,N_39526,N_38806);
nand U41329 (N_41329,N_37176,N_35743);
nor U41330 (N_41330,N_38817,N_39321);
nor U41331 (N_41331,N_39340,N_37976);
or U41332 (N_41332,N_36368,N_38386);
nand U41333 (N_41333,N_39405,N_37493);
nor U41334 (N_41334,N_38720,N_36197);
nand U41335 (N_41335,N_38814,N_36411);
nor U41336 (N_41336,N_39937,N_37650);
nor U41337 (N_41337,N_39389,N_37470);
nand U41338 (N_41338,N_38138,N_38204);
and U41339 (N_41339,N_38488,N_37250);
and U41340 (N_41340,N_37744,N_37217);
nand U41341 (N_41341,N_35307,N_36776);
and U41342 (N_41342,N_37053,N_38463);
and U41343 (N_41343,N_37170,N_38340);
nand U41344 (N_41344,N_39574,N_39464);
and U41345 (N_41345,N_39376,N_37085);
nand U41346 (N_41346,N_37144,N_38989);
and U41347 (N_41347,N_36420,N_39366);
nand U41348 (N_41348,N_38932,N_35203);
or U41349 (N_41349,N_36527,N_35801);
nor U41350 (N_41350,N_37501,N_39559);
or U41351 (N_41351,N_36414,N_37035);
nor U41352 (N_41352,N_38335,N_38857);
and U41353 (N_41353,N_37270,N_38564);
nor U41354 (N_41354,N_39205,N_39504);
xnor U41355 (N_41355,N_38928,N_39928);
or U41356 (N_41356,N_39867,N_38703);
and U41357 (N_41357,N_38251,N_37412);
nor U41358 (N_41358,N_37892,N_38750);
and U41359 (N_41359,N_39342,N_37482);
and U41360 (N_41360,N_38156,N_36433);
nand U41361 (N_41361,N_37758,N_35084);
and U41362 (N_41362,N_38359,N_37071);
nor U41363 (N_41363,N_38221,N_39525);
nor U41364 (N_41364,N_35878,N_39994);
xnor U41365 (N_41365,N_39180,N_39226);
or U41366 (N_41366,N_35901,N_37305);
or U41367 (N_41367,N_37816,N_38707);
nand U41368 (N_41368,N_38132,N_39666);
or U41369 (N_41369,N_35298,N_39244);
nand U41370 (N_41370,N_39805,N_37721);
and U41371 (N_41371,N_36761,N_39737);
or U41372 (N_41372,N_37865,N_35377);
and U41373 (N_41373,N_37233,N_39435);
or U41374 (N_41374,N_38230,N_35371);
nor U41375 (N_41375,N_39241,N_39222);
nand U41376 (N_41376,N_35174,N_37087);
or U41377 (N_41377,N_37225,N_35771);
and U41378 (N_41378,N_39941,N_37898);
nor U41379 (N_41379,N_35092,N_35992);
and U41380 (N_41380,N_38621,N_37340);
and U41381 (N_41381,N_39425,N_37285);
nand U41382 (N_41382,N_36193,N_37533);
nor U41383 (N_41383,N_39461,N_39537);
xor U41384 (N_41384,N_38023,N_35210);
nor U41385 (N_41385,N_39477,N_38936);
and U41386 (N_41386,N_39973,N_36924);
nor U41387 (N_41387,N_37272,N_38239);
nor U41388 (N_41388,N_39500,N_36591);
nand U41389 (N_41389,N_35846,N_37861);
or U41390 (N_41390,N_37610,N_37444);
nand U41391 (N_41391,N_36633,N_39861);
nor U41392 (N_41392,N_37383,N_36164);
xnor U41393 (N_41393,N_35554,N_38000);
and U41394 (N_41394,N_39300,N_38452);
xor U41395 (N_41395,N_37730,N_37800);
nand U41396 (N_41396,N_37282,N_37633);
nor U41397 (N_41397,N_39842,N_37576);
or U41398 (N_41398,N_36707,N_35022);
nand U41399 (N_41399,N_38458,N_39691);
nor U41400 (N_41400,N_38966,N_38756);
nand U41401 (N_41401,N_37451,N_39636);
nor U41402 (N_41402,N_35072,N_38790);
xnor U41403 (N_41403,N_38173,N_35135);
nand U41404 (N_41404,N_39743,N_39254);
or U41405 (N_41405,N_37813,N_37759);
nand U41406 (N_41406,N_39650,N_38254);
nand U41407 (N_41407,N_39359,N_37373);
xnor U41408 (N_41408,N_38760,N_35930);
or U41409 (N_41409,N_35243,N_39775);
xnor U41410 (N_41410,N_36758,N_35080);
nor U41411 (N_41411,N_35834,N_39599);
xor U41412 (N_41412,N_37280,N_35330);
xnor U41413 (N_41413,N_38008,N_35350);
xor U41414 (N_41414,N_37530,N_37528);
xnor U41415 (N_41415,N_38524,N_37336);
nand U41416 (N_41416,N_36410,N_37575);
xor U41417 (N_41417,N_36691,N_36534);
xor U41418 (N_41418,N_35564,N_36177);
nand U41419 (N_41419,N_38172,N_38157);
nor U41420 (N_41420,N_38624,N_39121);
nor U41421 (N_41421,N_37598,N_36358);
and U41422 (N_41422,N_39747,N_37103);
and U41423 (N_41423,N_38378,N_35665);
xnor U41424 (N_41424,N_37566,N_37934);
nand U41425 (N_41425,N_37635,N_37258);
nand U41426 (N_41426,N_37246,N_38401);
or U41427 (N_41427,N_38408,N_39910);
xnor U41428 (N_41428,N_36237,N_38364);
nand U41429 (N_41429,N_39923,N_38291);
and U41430 (N_41430,N_37784,N_35884);
nor U41431 (N_41431,N_38987,N_35719);
nor U41432 (N_41432,N_36935,N_35938);
nand U41433 (N_41433,N_39773,N_37965);
nor U41434 (N_41434,N_37731,N_37161);
and U41435 (N_41435,N_39716,N_35100);
xnor U41436 (N_41436,N_36625,N_37503);
or U41437 (N_41437,N_38840,N_37797);
xnor U41438 (N_41438,N_37289,N_38331);
or U41439 (N_41439,N_38687,N_37474);
or U41440 (N_41440,N_38169,N_38904);
xnor U41441 (N_41441,N_35118,N_35230);
xnor U41442 (N_41442,N_38058,N_39335);
nand U41443 (N_41443,N_37564,N_37213);
xnor U41444 (N_41444,N_38716,N_35390);
nand U41445 (N_41445,N_37943,N_38295);
nor U41446 (N_41446,N_39145,N_37678);
nand U41447 (N_41447,N_38586,N_37168);
xnor U41448 (N_41448,N_37854,N_37518);
xnor U41449 (N_41449,N_35067,N_38894);
nand U41450 (N_41450,N_38620,N_39848);
nand U41451 (N_41451,N_35868,N_39201);
nor U41452 (N_41452,N_39132,N_39444);
nor U41453 (N_41453,N_38708,N_37186);
or U41454 (N_41454,N_38065,N_38934);
or U41455 (N_41455,N_37012,N_37955);
or U41456 (N_41456,N_39077,N_39789);
nor U41457 (N_41457,N_36714,N_37708);
or U41458 (N_41458,N_36407,N_38723);
nand U41459 (N_41459,N_39465,N_38588);
xnor U41460 (N_41460,N_39809,N_37659);
and U41461 (N_41461,N_38263,N_39467);
nor U41462 (N_41462,N_36688,N_39279);
nor U41463 (N_41463,N_36567,N_35423);
xor U41464 (N_41464,N_36623,N_37252);
or U41465 (N_41465,N_38530,N_39487);
nand U41466 (N_41466,N_38021,N_38653);
or U41467 (N_41467,N_38436,N_35866);
nand U41468 (N_41468,N_38681,N_39733);
or U41469 (N_41469,N_37954,N_37709);
xnor U41470 (N_41470,N_37490,N_36779);
xor U41471 (N_41471,N_38625,N_35450);
nand U41472 (N_41472,N_38550,N_35057);
nand U41473 (N_41473,N_36771,N_38054);
and U41474 (N_41474,N_39372,N_39248);
nor U41475 (N_41475,N_36055,N_36004);
nand U41476 (N_41476,N_35919,N_35433);
or U41477 (N_41477,N_36947,N_35800);
and U41478 (N_41478,N_39660,N_35343);
and U41479 (N_41479,N_39576,N_36981);
xor U41480 (N_41480,N_35237,N_39156);
or U41481 (N_41481,N_36998,N_38755);
or U41482 (N_41482,N_39889,N_35777);
nor U41483 (N_41483,N_35867,N_36777);
and U41484 (N_41484,N_39494,N_36728);
and U41485 (N_41485,N_39000,N_39892);
and U41486 (N_41486,N_38496,N_35528);
nand U41487 (N_41487,N_39874,N_37826);
nor U41488 (N_41488,N_37309,N_35500);
xnor U41489 (N_41489,N_39883,N_38923);
xnor U41490 (N_41490,N_36438,N_38827);
and U41491 (N_41491,N_37782,N_35668);
xnor U41492 (N_41492,N_37047,N_38961);
or U41493 (N_41493,N_37554,N_38585);
and U41494 (N_41494,N_35830,N_35282);
nor U41495 (N_41495,N_38013,N_35441);
and U41496 (N_41496,N_36953,N_39221);
xor U41497 (N_41497,N_37489,N_37851);
nor U41498 (N_41498,N_37492,N_37725);
xnor U41499 (N_41499,N_36305,N_37913);
and U41500 (N_41500,N_38842,N_38076);
nand U41501 (N_41501,N_38285,N_36849);
nand U41502 (N_41502,N_36809,N_38511);
or U41503 (N_41503,N_39208,N_35726);
and U41504 (N_41504,N_35820,N_39433);
xnor U41505 (N_41505,N_36360,N_35077);
xnor U41506 (N_41506,N_36060,N_38736);
nor U41507 (N_41507,N_39331,N_39084);
xor U41508 (N_41508,N_37251,N_36327);
nor U41509 (N_41509,N_36721,N_36169);
nor U41510 (N_41510,N_38100,N_35329);
and U41511 (N_41511,N_38570,N_35283);
nor U41512 (N_41512,N_35663,N_35293);
and U41513 (N_41513,N_35598,N_35692);
xnor U41514 (N_41514,N_38235,N_38910);
nor U41515 (N_41515,N_38116,N_36394);
and U41516 (N_41516,N_39361,N_35095);
xor U41517 (N_41517,N_36293,N_37882);
or U41518 (N_41518,N_35652,N_37984);
nand U41519 (N_41519,N_35766,N_36300);
nor U41520 (N_41520,N_35339,N_39781);
nor U41521 (N_41521,N_36253,N_38284);
xnor U41522 (N_41522,N_37060,N_38580);
nand U41523 (N_41523,N_38145,N_37203);
nor U41524 (N_41524,N_35170,N_36442);
or U41525 (N_41525,N_38175,N_38922);
nand U41526 (N_41526,N_37165,N_37037);
xor U41527 (N_41527,N_36715,N_38973);
nand U41528 (N_41528,N_37326,N_37480);
or U41529 (N_41529,N_39462,N_39938);
xor U41530 (N_41530,N_37260,N_36201);
xnor U41531 (N_41531,N_38992,N_37595);
or U41532 (N_41532,N_38532,N_35748);
and U41533 (N_41533,N_39931,N_38434);
or U41534 (N_41534,N_35115,N_36529);
nand U41535 (N_41535,N_35912,N_36911);
nand U41536 (N_41536,N_36723,N_35640);
and U41537 (N_41537,N_36217,N_36424);
xnor U41538 (N_41538,N_35353,N_35871);
xor U41539 (N_41539,N_36572,N_37521);
nor U41540 (N_41540,N_38043,N_37511);
or U41541 (N_41541,N_38544,N_39729);
and U41542 (N_41542,N_38889,N_38612);
nand U41543 (N_41543,N_36763,N_38753);
or U41544 (N_41544,N_39507,N_35381);
nand U41545 (N_41545,N_36208,N_39728);
nor U41546 (N_41546,N_36051,N_39879);
nor U41547 (N_41547,N_37346,N_35523);
or U41548 (N_41548,N_35125,N_37302);
nor U41549 (N_41549,N_37205,N_36445);
nor U41550 (N_41550,N_35394,N_37739);
or U41551 (N_41551,N_36072,N_36482);
xnor U41552 (N_41552,N_37334,N_36270);
or U41553 (N_41553,N_36791,N_35952);
or U41554 (N_41554,N_39667,N_36649);
and U41555 (N_41555,N_35233,N_35898);
and U41556 (N_41556,N_39278,N_36973);
nand U41557 (N_41557,N_38471,N_39586);
xor U41558 (N_41558,N_35437,N_35360);
or U41559 (N_41559,N_38298,N_39947);
xor U41560 (N_41560,N_39835,N_36258);
nor U41561 (N_41561,N_39627,N_39611);
or U41562 (N_41562,N_37300,N_39162);
nor U41563 (N_41563,N_38731,N_36143);
and U41564 (N_41564,N_35495,N_38576);
or U41565 (N_41565,N_37715,N_37290);
nor U41566 (N_41566,N_38775,N_37915);
nor U41567 (N_41567,N_37536,N_39219);
nor U41568 (N_41568,N_38855,N_37868);
nand U41569 (N_41569,N_39261,N_38410);
or U41570 (N_41570,N_35355,N_39546);
xnor U41571 (N_41571,N_36518,N_35504);
or U41572 (N_41572,N_36110,N_37629);
nor U41573 (N_41573,N_38237,N_39214);
xor U41574 (N_41574,N_39028,N_39609);
or U41575 (N_41575,N_38754,N_38414);
and U41576 (N_41576,N_37498,N_35984);
xnor U41577 (N_41577,N_36213,N_38207);
nand U41578 (N_41578,N_36778,N_37430);
xnor U41579 (N_41579,N_37519,N_37455);
nor U41580 (N_41580,N_39285,N_38648);
xnor U41581 (N_41581,N_35176,N_38969);
xor U41582 (N_41582,N_39603,N_37561);
nand U41583 (N_41583,N_39655,N_35153);
nand U41584 (N_41584,N_35623,N_39820);
or U41585 (N_41585,N_37461,N_36753);
nand U41586 (N_41586,N_36614,N_35027);
nand U41587 (N_41587,N_36644,N_38194);
or U41588 (N_41588,N_35370,N_36419);
or U41589 (N_41589,N_36725,N_37845);
or U41590 (N_41590,N_36921,N_36823);
nand U41591 (N_41591,N_39374,N_37335);
xor U41592 (N_41592,N_37226,N_37390);
or U41593 (N_41593,N_37006,N_38437);
nor U41594 (N_41594,N_38007,N_38637);
xor U41595 (N_41595,N_39661,N_37804);
nor U41596 (N_41596,N_37793,N_39184);
or U41597 (N_41597,N_37481,N_39088);
and U41598 (N_41598,N_38046,N_39845);
nand U41599 (N_41599,N_37712,N_38837);
and U41600 (N_41600,N_37555,N_35258);
nor U41601 (N_41601,N_37267,N_35586);
nand U41602 (N_41602,N_36992,N_35192);
xor U41603 (N_41603,N_37614,N_36900);
nand U41604 (N_41604,N_35465,N_39089);
nor U41605 (N_41605,N_38444,N_39521);
and U41606 (N_41606,N_36864,N_37331);
xnor U41607 (N_41607,N_39556,N_37269);
nand U41608 (N_41608,N_36296,N_35323);
nand U41609 (N_41609,N_38107,N_37360);
or U41610 (N_41610,N_35226,N_39590);
or U41611 (N_41611,N_38810,N_35224);
xor U41612 (N_41612,N_38946,N_35599);
nor U41613 (N_41613,N_36909,N_35266);
or U41614 (N_41614,N_37904,N_38598);
nand U41615 (N_41615,N_37382,N_39414);
nand U41616 (N_41616,N_38438,N_38730);
nand U41617 (N_41617,N_37616,N_39434);
or U41618 (N_41618,N_38485,N_37367);
and U41619 (N_41619,N_37673,N_35739);
nand U41620 (N_41620,N_37867,N_35384);
xnor U41621 (N_41621,N_37045,N_36333);
or U41622 (N_41622,N_35157,N_37507);
xor U41623 (N_41623,N_38184,N_36677);
and U41624 (N_41624,N_38962,N_36341);
or U41625 (N_41625,N_36643,N_37406);
nand U41626 (N_41626,N_39417,N_38609);
nand U41627 (N_41627,N_39951,N_39074);
or U41628 (N_41628,N_37924,N_38581);
and U41629 (N_41629,N_35088,N_38650);
and U41630 (N_41630,N_36873,N_39644);
nor U41631 (N_41631,N_37932,N_39997);
xnor U41632 (N_41632,N_39063,N_37089);
or U41633 (N_41633,N_36122,N_39795);
xnor U41634 (N_41634,N_38597,N_37433);
or U41635 (N_41635,N_36146,N_36888);
or U41636 (N_41636,N_37919,N_39383);
nor U41637 (N_41637,N_39750,N_39600);
nor U41638 (N_41638,N_36448,N_37241);
nand U41639 (N_41639,N_36526,N_37207);
nor U41640 (N_41640,N_39777,N_39336);
and U41641 (N_41641,N_35155,N_37667);
nand U41642 (N_41642,N_37956,N_39513);
nand U41643 (N_41643,N_35162,N_36589);
xor U41644 (N_41644,N_38640,N_38713);
nor U41645 (N_41645,N_37582,N_37109);
nand U41646 (N_41646,N_39303,N_37770);
nand U41647 (N_41647,N_36488,N_38083);
and U41648 (N_41648,N_39700,N_38523);
or U41649 (N_41649,N_38745,N_35078);
nand U41650 (N_41650,N_39610,N_39129);
xor U41651 (N_41651,N_36595,N_38208);
nor U41652 (N_41652,N_39163,N_37386);
nor U41653 (N_41653,N_35605,N_38487);
nor U41654 (N_41654,N_39030,N_35827);
nand U41655 (N_41655,N_39492,N_38623);
xnor U41656 (N_41656,N_36191,N_39388);
xnor U41657 (N_41657,N_38592,N_39064);
and U41658 (N_41658,N_39868,N_35720);
or U41659 (N_41659,N_38921,N_39962);
nor U41660 (N_41660,N_38427,N_35064);
or U41661 (N_41661,N_38663,N_38320);
xnor U41662 (N_41662,N_37795,N_36759);
nor U41663 (N_41663,N_38830,N_37355);
nand U41664 (N_41664,N_36676,N_35695);
xnor U41665 (N_41665,N_39617,N_39841);
or U41666 (N_41666,N_36172,N_36492);
and U41667 (N_41667,N_38852,N_38261);
nand U41668 (N_41668,N_38108,N_38215);
nand U41669 (N_41669,N_38010,N_36240);
and U41670 (N_41670,N_36196,N_37939);
or U41671 (N_41671,N_38866,N_35173);
xnor U41672 (N_41672,N_37193,N_38447);
nor U41673 (N_41673,N_37500,N_38943);
xor U41674 (N_41674,N_37052,N_39975);
xnor U41675 (N_41675,N_37093,N_35101);
and U41676 (N_41676,N_36500,N_39560);
nor U41677 (N_41677,N_39907,N_35578);
nor U41678 (N_41678,N_37198,N_35229);
nor U41679 (N_41679,N_36566,N_37431);
nand U41680 (N_41680,N_36964,N_35199);
nor U41681 (N_41681,N_37119,N_37505);
or U41682 (N_41682,N_39212,N_38042);
xnor U41683 (N_41683,N_39200,N_36262);
nor U41684 (N_41684,N_35402,N_36042);
or U41685 (N_41685,N_36229,N_36599);
nor U41686 (N_41686,N_37452,N_38390);
xnor U41687 (N_41687,N_35491,N_39380);
nor U41688 (N_41688,N_37916,N_36929);
nand U41689 (N_41689,N_36131,N_39149);
nand U41690 (N_41690,N_37033,N_38053);
or U41691 (N_41691,N_36264,N_35524);
nand U41692 (N_41692,N_39816,N_38326);
nor U41693 (N_41693,N_39799,N_37930);
nor U41694 (N_41694,N_36592,N_38308);
and U41695 (N_41695,N_38543,N_38375);
and U41696 (N_41696,N_37278,N_36231);
and U41697 (N_41697,N_39614,N_39904);
or U41698 (N_41698,N_36689,N_39967);
and U41699 (N_41699,N_36509,N_35507);
or U41700 (N_41700,N_35109,N_37662);
nand U41701 (N_41701,N_38773,N_35736);
and U41702 (N_41702,N_37342,N_38212);
xor U41703 (N_41703,N_36937,N_38282);
xor U41704 (N_41704,N_37011,N_37253);
nor U41705 (N_41705,N_35455,N_36086);
or U41706 (N_41706,N_35712,N_36417);
xnor U41707 (N_41707,N_35130,N_36871);
and U41708 (N_41708,N_39498,N_35986);
and U41709 (N_41709,N_36974,N_36204);
nand U41710 (N_41710,N_35347,N_39231);
and U41711 (N_41711,N_35634,N_36171);
and U41712 (N_41712,N_35004,N_39558);
and U41713 (N_41713,N_39220,N_39528);
nor U41714 (N_41714,N_38079,N_36934);
and U41715 (N_41715,N_39235,N_38679);
nor U41716 (N_41716,N_37856,N_35315);
or U41717 (N_41717,N_35534,N_38062);
nand U41718 (N_41718,N_37422,N_39822);
nor U41719 (N_41719,N_37014,N_39112);
and U41720 (N_41720,N_38429,N_38950);
or U41721 (N_41721,N_39778,N_37065);
xnor U41722 (N_41722,N_36596,N_36631);
and U41723 (N_41723,N_36286,N_38224);
and U41724 (N_41724,N_37751,N_36798);
or U41725 (N_41725,N_36735,N_37817);
xnor U41726 (N_41726,N_36019,N_37559);
or U41727 (N_41727,N_38310,N_38846);
nor U41728 (N_41728,N_38558,N_36450);
or U41729 (N_41729,N_38441,N_35741);
xnor U41730 (N_41730,N_38796,N_35526);
or U41731 (N_41731,N_36508,N_35488);
and U41732 (N_41732,N_35655,N_36581);
and U41733 (N_41733,N_36826,N_36975);
xnor U41734 (N_41734,N_39081,N_39116);
or U41735 (N_41735,N_35301,N_38417);
and U41736 (N_41736,N_36788,N_37136);
nand U41737 (N_41737,N_39344,N_37643);
or U41738 (N_41738,N_35019,N_39294);
nand U41739 (N_41739,N_37277,N_36045);
xnor U41740 (N_41740,N_39670,N_36786);
or U41741 (N_41741,N_35058,N_39365);
or U41742 (N_41742,N_35025,N_38868);
nand U41743 (N_41743,N_36413,N_38574);
nor U41744 (N_41744,N_39839,N_39790);
and U41745 (N_41745,N_39772,N_39443);
nor U41746 (N_41746,N_36412,N_39782);
or U41747 (N_41747,N_36962,N_35818);
or U41748 (N_41748,N_36036,N_39553);
or U41749 (N_41749,N_39616,N_38557);
and U41750 (N_41750,N_39575,N_36683);
nand U41751 (N_41751,N_38636,N_37010);
nor U41752 (N_41752,N_36582,N_37408);
nor U41753 (N_41753,N_35604,N_37293);
nand U41754 (N_41754,N_38805,N_37773);
nand U41755 (N_41755,N_39137,N_36894);
nor U41756 (N_41756,N_38255,N_38940);
and U41757 (N_41757,N_35201,N_39828);
xor U41758 (N_41758,N_37142,N_36260);
and U41759 (N_41759,N_39499,N_39267);
xor U41760 (N_41760,N_39563,N_39682);
xnor U41761 (N_41761,N_36344,N_38839);
nand U41762 (N_41762,N_35456,N_38799);
nor U41763 (N_41763,N_35791,N_38832);
nor U41764 (N_41764,N_39460,N_37853);
xor U41765 (N_41765,N_39072,N_35995);
nand U41766 (N_41766,N_38139,N_35120);
xor U41767 (N_41767,N_36854,N_37159);
xor U41768 (N_41768,N_36163,N_39295);
nand U41769 (N_41769,N_35643,N_35760);
and U41770 (N_41770,N_35035,N_37249);
nand U41771 (N_41771,N_36388,N_37697);
nand U41772 (N_41772,N_37696,N_39811);
nor U41773 (N_41773,N_36101,N_36949);
xnor U41774 (N_41774,N_39151,N_35331);
nor U41775 (N_41775,N_38607,N_38541);
nor U41776 (N_41776,N_37473,N_39339);
xor U41777 (N_41777,N_39110,N_37525);
nor U41778 (N_41778,N_39823,N_39618);
or U41779 (N_41779,N_37897,N_35538);
nand U41780 (N_41780,N_36600,N_36898);
xor U41781 (N_41781,N_35138,N_37945);
and U41782 (N_41782,N_37404,N_39245);
and U41783 (N_41783,N_35421,N_37726);
nand U41784 (N_41784,N_35953,N_35469);
xor U41785 (N_41785,N_35391,N_35191);
and U41786 (N_41786,N_36895,N_39015);
nand U41787 (N_41787,N_38094,N_39643);
and U41788 (N_41788,N_36757,N_38180);
or U41789 (N_41789,N_35890,N_36076);
and U41790 (N_41790,N_39763,N_37727);
or U41791 (N_41791,N_37101,N_39275);
nand U41792 (N_41792,N_36770,N_36230);
xnor U41793 (N_41793,N_37419,N_35477);
and U41794 (N_41794,N_36380,N_35758);
nand U41795 (N_41795,N_36882,N_36720);
and U41796 (N_41796,N_37756,N_35449);
nand U41797 (N_41797,N_35778,N_35066);
nand U41798 (N_41798,N_38662,N_37565);
nor U41799 (N_41799,N_36576,N_38018);
nand U41800 (N_41800,N_35209,N_39439);
xor U41801 (N_41801,N_36653,N_38825);
xnor U41802 (N_41802,N_38090,N_37605);
xor U41803 (N_41803,N_36328,N_36175);
nand U41804 (N_41804,N_35619,N_37979);
nor U41805 (N_41805,N_36912,N_36499);
xor U41806 (N_41806,N_39350,N_37445);
nand U41807 (N_41807,N_39983,N_38192);
nand U41808 (N_41808,N_38965,N_36079);
nand U41809 (N_41809,N_39512,N_36636);
and U41810 (N_41810,N_36563,N_38486);
and U41811 (N_41811,N_37931,N_37066);
nand U41812 (N_41812,N_37679,N_35414);
nor U41813 (N_41813,N_39587,N_37067);
and U41814 (N_41814,N_36335,N_38725);
and U41815 (N_41815,N_36280,N_35223);
nor U41816 (N_41816,N_35039,N_36449);
nand U41817 (N_41817,N_37872,N_36128);
nor U41818 (N_41818,N_36173,N_39264);
nor U41819 (N_41819,N_39502,N_38626);
xnor U41820 (N_41820,N_37541,N_35172);
xnor U41821 (N_41821,N_35413,N_35998);
and U41822 (N_41822,N_39228,N_35139);
xnor U41823 (N_41823,N_36708,N_38911);
or U41824 (N_41824,N_35680,N_36782);
nor U41825 (N_41825,N_36068,N_39649);
nand U41826 (N_41826,N_39974,N_37888);
and U41827 (N_41827,N_38781,N_37042);
and U41828 (N_41828,N_39702,N_37427);
nor U41829 (N_41829,N_35764,N_35511);
or U41830 (N_41830,N_39505,N_38722);
nand U41831 (N_41831,N_39305,N_36302);
or U41832 (N_41832,N_37003,N_37296);
and U41833 (N_41833,N_38812,N_36202);
nor U41834 (N_41834,N_39903,N_35627);
xor U41835 (N_41835,N_39930,N_39565);
xor U41836 (N_41836,N_39909,N_36148);
nor U41837 (N_41837,N_35045,N_38057);
xnor U41838 (N_41838,N_35046,N_39354);
or U41839 (N_41839,N_35725,N_37792);
xnor U41840 (N_41840,N_38770,N_36554);
nor U41841 (N_41841,N_36802,N_39019);
xor U41842 (N_41842,N_39304,N_36035);
xnor U41843 (N_41843,N_39672,N_36084);
xor U41844 (N_41844,N_39230,N_37023);
nor U41845 (N_41845,N_36160,N_37306);
or U41846 (N_41846,N_36465,N_35144);
nand U41847 (N_41847,N_38306,N_37458);
or U41848 (N_41848,N_39262,N_39759);
nand U41849 (N_41849,N_37243,N_38140);
or U41850 (N_41850,N_36167,N_35166);
nor U41851 (N_41851,N_35854,N_37015);
nor U41852 (N_41852,N_37857,N_38186);
and U41853 (N_41853,N_37379,N_39547);
and U41854 (N_41854,N_39870,N_37130);
and U41855 (N_41855,N_38356,N_38957);
xor U41856 (N_41856,N_38718,N_38322);
and U41857 (N_41857,N_37831,N_37597);
nor U41858 (N_41858,N_37749,N_37039);
or U41859 (N_41859,N_39134,N_38244);
nand U41860 (N_41860,N_36738,N_36385);
nand U41861 (N_41861,N_35295,N_36268);
nand U41862 (N_41862,N_38467,N_37762);
or U41863 (N_41863,N_39160,N_36963);
or U41864 (N_41864,N_38668,N_35136);
and U41865 (N_41865,N_36860,N_35849);
or U41866 (N_41866,N_35563,N_38129);
nand U41867 (N_41867,N_36198,N_37143);
xnor U41868 (N_41868,N_36654,N_37967);
nand U41869 (N_41869,N_38924,N_35546);
nand U41870 (N_41870,N_35415,N_37317);
or U41871 (N_41871,N_37508,N_37214);
or U41872 (N_41872,N_38614,N_36752);
xnor U41873 (N_41873,N_38424,N_38376);
and U41874 (N_41874,N_37348,N_38638);
or U41875 (N_41875,N_38983,N_39159);
nand U41876 (N_41876,N_37462,N_35214);
or U41877 (N_41877,N_35747,N_36453);
nand U41878 (N_41878,N_38602,N_38947);
nor U41879 (N_41879,N_36044,N_38232);
xor U41880 (N_41880,N_35590,N_38824);
or U41881 (N_41881,N_38672,N_35126);
nor U41882 (N_41882,N_35666,N_35529);
nor U41883 (N_41883,N_39202,N_37104);
and U41884 (N_41884,N_36817,N_37129);
nor U41885 (N_41885,N_35086,N_36594);
nand U41886 (N_41886,N_38131,N_38142);
nor U41887 (N_41887,N_35746,N_37380);
xor U41888 (N_41888,N_35851,N_39765);
nor U41889 (N_41889,N_39386,N_39229);
nor U41890 (N_41890,N_36952,N_35893);
nor U41891 (N_41891,N_38121,N_38381);
nand U41892 (N_41892,N_37642,N_37808);
or U41893 (N_41893,N_37768,N_36458);
xnor U41894 (N_41894,N_39095,N_36012);
and U41895 (N_41895,N_38657,N_39060);
and U41896 (N_41896,N_36958,N_38651);
nor U41897 (N_41897,N_35430,N_36719);
nand U41898 (N_41898,N_35895,N_39944);
or U41899 (N_41899,N_39297,N_39257);
or U41900 (N_41900,N_38143,N_36115);
and U41901 (N_41901,N_39815,N_35978);
and U41902 (N_41902,N_38164,N_35753);
nor U41903 (N_41903,N_39004,N_37245);
xor U41904 (N_41904,N_37918,N_35167);
or U41905 (N_41905,N_39803,N_38933);
or U41906 (N_41906,N_39101,N_36314);
and U41907 (N_41907,N_39533,N_36747);
nor U41908 (N_41908,N_39050,N_36007);
nand U41909 (N_41909,N_39995,N_37083);
or U41910 (N_41910,N_38159,N_36400);
and U41911 (N_41911,N_39851,N_39935);
and U41912 (N_41912,N_36259,N_39320);
nor U41913 (N_41913,N_37414,N_35451);
nand U41914 (N_41914,N_38960,N_35950);
nor U41915 (N_41915,N_38044,N_38568);
nor U41916 (N_41916,N_36289,N_36093);
or U41917 (N_41917,N_37212,N_36807);
nor U41918 (N_41918,N_38472,N_36856);
or U41919 (N_41919,N_36539,N_36686);
and U41920 (N_41920,N_38803,N_37338);
and U41921 (N_41921,N_36642,N_37124);
and U41922 (N_41922,N_39819,N_38862);
and U41923 (N_41923,N_39578,N_37411);
and U41924 (N_41924,N_39410,N_36972);
xor U41925 (N_41925,N_35427,N_36559);
and U41926 (N_41926,N_37174,N_38639);
nand U41927 (N_41927,N_38907,N_38699);
and U41928 (N_41928,N_38764,N_35447);
nor U41929 (N_41929,N_35510,N_37004);
and U41930 (N_41930,N_37950,N_39866);
and U41931 (N_41931,N_35356,N_35399);
xnor U41932 (N_41932,N_38097,N_37292);
xor U41933 (N_41933,N_36632,N_36232);
or U41934 (N_41934,N_39552,N_35744);
or U41935 (N_41935,N_36841,N_38392);
xnor U41936 (N_41936,N_35580,N_35509);
xor U41937 (N_41937,N_36664,N_35842);
nand U41938 (N_41938,N_37810,N_38642);
xnor U41939 (N_41939,N_35769,N_35761);
or U41940 (N_41940,N_39495,N_38710);
nor U41941 (N_41941,N_36835,N_36120);
and U41942 (N_41942,N_39568,N_39086);
nand U41943 (N_41943,N_37264,N_35921);
or U41944 (N_41944,N_39834,N_36987);
and U41945 (N_41945,N_35539,N_36063);
nand U41946 (N_41946,N_37152,N_36742);
or U41947 (N_41947,N_38351,N_38411);
and U41948 (N_41948,N_37884,N_36583);
and U41949 (N_41949,N_39440,N_35177);
nor U41950 (N_41950,N_39557,N_38513);
xnor U41951 (N_41951,N_37776,N_39152);
nor U41952 (N_41952,N_38994,N_39011);
and U41953 (N_41953,N_39859,N_35567);
nor U41954 (N_41954,N_36884,N_38762);
or U41955 (N_41955,N_36814,N_39760);
xor U41956 (N_41956,N_37421,N_35478);
and U41957 (N_41957,N_39635,N_39515);
xor U41958 (N_41958,N_38734,N_36452);
nor U41959 (N_41959,N_36821,N_39704);
xor U41960 (N_41960,N_39044,N_35043);
and U41961 (N_41961,N_37649,N_37137);
xor U41962 (N_41962,N_35194,N_38379);
or U41963 (N_41963,N_35253,N_37757);
nor U41964 (N_41964,N_38914,N_37141);
nand U41965 (N_41965,N_36185,N_39762);
nand U41966 (N_41966,N_37858,N_37189);
nand U41967 (N_41967,N_37491,N_36825);
xor U41968 (N_41968,N_36255,N_37148);
and U41969 (N_41969,N_39680,N_38031);
nand U41970 (N_41970,N_35028,N_36451);
or U41971 (N_41971,N_39651,N_38976);
nor U41972 (N_41972,N_35654,N_36558);
nand U41973 (N_41973,N_36769,N_39346);
nand U41974 (N_41974,N_36491,N_38686);
and U41975 (N_41975,N_36064,N_37055);
nand U41976 (N_41976,N_39291,N_39176);
xnor U41977 (N_41977,N_39165,N_37368);
xnor U41978 (N_41978,N_37690,N_39059);
or U41979 (N_41979,N_35322,N_38395);
xor U41980 (N_41980,N_38270,N_37743);
xnor U41981 (N_41981,N_37210,N_37844);
xnor U41982 (N_41982,N_36792,N_36234);
nand U41983 (N_41983,N_36373,N_35154);
nand U41984 (N_41984,N_39117,N_35559);
or U41985 (N_41985,N_35492,N_39612);
nand U41986 (N_41986,N_36930,N_39605);
or U41987 (N_41987,N_38026,N_35899);
nor U41988 (N_41988,N_35184,N_38337);
nor U41989 (N_41989,N_37327,N_36547);
xor U41990 (N_41990,N_38422,N_36945);
xnor U41991 (N_41991,N_37323,N_35202);
xor U41992 (N_41992,N_36376,N_35178);
xor U41993 (N_41993,N_36858,N_38737);
xor U41994 (N_41994,N_38861,N_38851);
or U41995 (N_41995,N_39633,N_37824);
nor U41996 (N_41996,N_38743,N_35005);
xnor U41997 (N_41997,N_38949,N_38536);
nand U41998 (N_41998,N_38798,N_36699);
xnor U41999 (N_41999,N_38373,N_39419);
nand U42000 (N_42000,N_35701,N_35572);
and U42001 (N_42001,N_36105,N_38865);
nand U42002 (N_42002,N_38974,N_35123);
nor U42003 (N_42003,N_35036,N_39711);
or U42004 (N_42004,N_36489,N_35807);
xnor U42005 (N_42005,N_39310,N_36847);
or U42006 (N_42006,N_39210,N_35659);
nand U42007 (N_42007,N_36969,N_38882);
nand U42008 (N_42008,N_35759,N_35636);
or U42009 (N_42009,N_39539,N_35464);
or U42010 (N_42010,N_39821,N_39976);
nand U42011 (N_42011,N_35616,N_36033);
nor U42012 (N_42012,N_37399,N_37869);
xnor U42013 (N_42013,N_37345,N_37247);
nor U42014 (N_42014,N_37497,N_35979);
nor U42015 (N_42015,N_38559,N_35837);
nor U42016 (N_42016,N_36140,N_38526);
and U42017 (N_42017,N_36658,N_35425);
xor U42018 (N_42018,N_36242,N_35943);
or U42019 (N_42019,N_38415,N_36618);
and U42020 (N_42020,N_35629,N_38684);
or U42021 (N_42021,N_39447,N_38082);
nor U42022 (N_42022,N_35903,N_36460);
or U42023 (N_42023,N_35446,N_39946);
or U42024 (N_42024,N_38807,N_39693);
xnor U42025 (N_42025,N_39566,N_35688);
and U42026 (N_42026,N_37155,N_37713);
or U42027 (N_42027,N_38892,N_35038);
nor U42028 (N_42028,N_36070,N_36446);
xor U42029 (N_42029,N_36531,N_38353);
and U42030 (N_42030,N_39689,N_35105);
and U42031 (N_42031,N_39363,N_39236);
xor U42032 (N_42032,N_36363,N_36662);
nand U42033 (N_42033,N_37229,N_38908);
or U42034 (N_42034,N_35730,N_36029);
nand U42035 (N_42035,N_39265,N_39623);
nand U42036 (N_42036,N_35691,N_39668);
nor U42037 (N_42037,N_35397,N_37783);
and U42038 (N_42038,N_36046,N_37477);
nor U42039 (N_42039,N_36982,N_38491);
nor U42040 (N_42040,N_37476,N_39436);
nand U42041 (N_42041,N_39276,N_36663);
and U42042 (N_42042,N_39153,N_39985);
and U42043 (N_42043,N_38346,N_36135);
xnor U42044 (N_42044,N_36416,N_35263);
and U42045 (N_42045,N_36540,N_37183);
and U42046 (N_42046,N_38025,N_38884);
nand U42047 (N_42047,N_39757,N_38808);
nand U42048 (N_42048,N_37082,N_35183);
or U42049 (N_42049,N_35448,N_35888);
or U42050 (N_42050,N_38233,N_37531);
nor U42051 (N_42051,N_39637,N_35975);
xor U42052 (N_42052,N_35257,N_35886);
nor U42053 (N_42053,N_39270,N_39100);
nand U42054 (N_42054,N_37361,N_38336);
xnor U42055 (N_42055,N_39969,N_35034);
and U42056 (N_42056,N_38274,N_37437);
and U42057 (N_42057,N_37513,N_36928);
xor U42058 (N_42058,N_35667,N_36283);
or U42059 (N_42059,N_37911,N_39943);
and U42060 (N_42060,N_38665,N_36277);
nand U42061 (N_42061,N_36744,N_39582);
nor U42062 (N_42062,N_38579,N_39602);
or U42063 (N_42063,N_37450,N_35570);
nand U42064 (N_42064,N_35140,N_35121);
nand U42065 (N_42065,N_36837,N_36665);
nand U42066 (N_42066,N_35400,N_36238);
xnor U42067 (N_42067,N_38925,N_39497);
nor U42068 (N_42068,N_35149,N_35601);
xor U42069 (N_42069,N_38542,N_37982);
nand U42070 (N_42070,N_36885,N_35543);
or U42071 (N_42071,N_39957,N_35457);
nor U42072 (N_42072,N_36392,N_39122);
xor U42073 (N_42073,N_39844,N_37510);
or U42074 (N_42074,N_35792,N_35525);
or U42075 (N_42075,N_38269,N_36611);
nand U42076 (N_42076,N_37879,N_35386);
xnor U42077 (N_42077,N_38199,N_36651);
xor U42078 (N_42078,N_35312,N_37163);
xor U42079 (N_42079,N_36913,N_38174);
xnor U42080 (N_42080,N_37828,N_35702);
nand U42081 (N_42081,N_35182,N_37562);
xnor U42082 (N_42082,N_39370,N_37560);
and U42083 (N_42083,N_35957,N_38898);
nor U42084 (N_42084,N_39451,N_37902);
nor U42085 (N_42085,N_37308,N_35300);
and U42086 (N_42086,N_35029,N_35181);
and U42087 (N_42087,N_35404,N_35247);
xor U42088 (N_42088,N_37670,N_36031);
xor U42089 (N_42089,N_39292,N_39766);
nand U42090 (N_42090,N_35274,N_37668);
nor U42091 (N_42091,N_36768,N_35639);
nand U42092 (N_42092,N_39857,N_36479);
xor U42093 (N_42093,N_37767,N_35389);
or U42094 (N_42094,N_39415,N_39917);
or U42095 (N_42095,N_36557,N_38278);
and U42096 (N_42096,N_39638,N_36698);
or U42097 (N_42097,N_38948,N_36018);
xnor U42098 (N_42098,N_35050,N_38666);
nand U42099 (N_42099,N_38311,N_35929);
nor U42100 (N_42100,N_37901,N_38502);
xnor U42101 (N_42101,N_35128,N_37472);
nor U42102 (N_42102,N_38793,N_39092);
nor U42103 (N_42103,N_35512,N_38853);
nor U42104 (N_42104,N_35501,N_36389);
and U42105 (N_42105,N_37150,N_38881);
and U42106 (N_42106,N_36593,N_35941);
nand U42107 (N_42107,N_39632,N_36510);
xnor U42108 (N_42108,N_39900,N_36926);
or U42109 (N_42109,N_39800,N_37711);
nand U42110 (N_42110,N_36743,N_38104);
or U42111 (N_42111,N_35467,N_38084);
nor U42112 (N_42112,N_39608,N_38419);
and U42113 (N_42113,N_36889,N_39899);
and U42114 (N_42114,N_39685,N_39143);
xor U42115 (N_42115,N_36144,N_35150);
nand U42116 (N_42116,N_35657,N_39418);
nor U42117 (N_42117,N_37038,N_38072);
nand U42118 (N_42118,N_39745,N_36484);
nand U42119 (N_42119,N_36075,N_35117);
xnor U42120 (N_42120,N_38360,N_38670);
and U42121 (N_42121,N_38098,N_37471);
nor U42122 (N_42122,N_39450,N_37238);
and U42123 (N_42123,N_39657,N_39273);
or U42124 (N_42124,N_37232,N_39598);
xor U42125 (N_42125,N_39432,N_35519);
nand U42126 (N_42126,N_39457,N_39406);
xnor U42127 (N_42127,N_36461,N_37880);
nand U42128 (N_42128,N_36399,N_35065);
or U42129 (N_42129,N_35059,N_39031);
xor U42130 (N_42130,N_35794,N_38792);
nand U42131 (N_42131,N_35676,N_39787);
nand U42132 (N_42132,N_37221,N_38296);
nor U42133 (N_42133,N_39961,N_38027);
nand U42134 (N_42134,N_39256,N_36616);
nor U42135 (N_42135,N_36356,N_36342);
nor U42136 (N_42136,N_38066,N_39972);
xnor U42137 (N_42137,N_36152,N_39390);
nor U42138 (N_42138,N_35483,N_37933);
nor U42139 (N_42139,N_38045,N_37683);
and U42140 (N_42140,N_38548,N_38700);
or U42141 (N_42141,N_36040,N_39577);
nand U42142 (N_42142,N_39621,N_36329);
nand U42143 (N_42143,N_37469,N_37324);
nand U42144 (N_42144,N_39218,N_39977);
nand U42145 (N_42145,N_38647,N_35254);
xor U42146 (N_42146,N_39530,N_39103);
nand U42147 (N_42147,N_35631,N_35716);
or U42148 (N_42148,N_36556,N_37268);
nand U42149 (N_42149,N_39686,N_36359);
nor U42150 (N_42150,N_36717,N_39322);
nand U42151 (N_42151,N_37099,N_35797);
nand U42152 (N_42152,N_37896,N_36272);
nand U42153 (N_42153,N_37855,N_36995);
xor U42154 (N_42154,N_37714,N_39768);
nand U42155 (N_42155,N_35419,N_35333);
nor U42156 (N_42156,N_36224,N_35480);
xnor U42157 (N_42157,N_38483,N_36109);
and U42158 (N_42158,N_36049,N_35292);
nor U42159 (N_42159,N_37987,N_38664);
nand U42160 (N_42160,N_36038,N_37971);
nand U42161 (N_42161,N_39692,N_38420);
nor U42162 (N_42162,N_38655,N_35366);
xnor U42163 (N_42163,N_36997,N_39293);
nor U42164 (N_42164,N_35951,N_35246);
or U42165 (N_42165,N_35927,N_36228);
nand U42166 (N_42166,N_37032,N_35836);
nor U42167 (N_42167,N_37029,N_37658);
and U42168 (N_42168,N_36444,N_38749);
nand U42169 (N_42169,N_39033,N_39628);
and U42170 (N_42170,N_39364,N_36684);
xnor U42171 (N_42171,N_39966,N_39455);
nor U42172 (N_42172,N_38126,N_38771);
and U42173 (N_42173,N_39345,N_36827);
xnor U42174 (N_42174,N_37639,N_39895);
xor U42175 (N_42175,N_38535,N_37772);
or U42176 (N_42176,N_39227,N_38540);
or U42177 (N_42177,N_38733,N_37240);
and U42178 (N_42178,N_38355,N_39029);
or U42179 (N_42179,N_39035,N_37051);
or U42180 (N_42180,N_36282,N_39981);
nand U42181 (N_42181,N_36306,N_38995);
or U42182 (N_42182,N_35795,N_36014);
nand U42183 (N_42183,N_37059,N_39195);
nor U42184 (N_42184,N_36984,N_35349);
nor U42185 (N_42185,N_35369,N_37547);
nand U42186 (N_42186,N_39579,N_36502);
nor U42187 (N_42187,N_35679,N_37641);
nand U42188 (N_42188,N_39894,N_39999);
xnor U42189 (N_42189,N_35403,N_37112);
xnor U42190 (N_42190,N_35535,N_36748);
xnor U42191 (N_42191,N_37747,N_39488);
or U42192 (N_42192,N_36586,N_38804);
xnor U42193 (N_42193,N_35219,N_37409);
and U42194 (N_42194,N_38464,N_38970);
and U42195 (N_42195,N_38009,N_39287);
or U42196 (N_42196,N_36956,N_39740);
nor U42197 (N_42197,N_38659,N_37648);
xnor U42198 (N_42198,N_39172,N_38482);
nand U42199 (N_42199,N_35362,N_36147);
and U42200 (N_42200,N_38521,N_36351);
nand U42201 (N_42201,N_39428,N_38603);
and U42202 (N_42202,N_35615,N_35891);
or U42203 (N_42203,N_38334,N_36048);
nand U42204 (N_42204,N_36685,N_36235);
and U42205 (N_42205,N_36361,N_35565);
nand U42206 (N_42206,N_38864,N_37418);
nand U42207 (N_42207,N_36320,N_37192);
and U42208 (N_42208,N_36236,N_35508);
or U42209 (N_42209,N_36690,N_36494);
nor U42210 (N_42210,N_35434,N_35142);
or U42211 (N_42211,N_35108,N_35468);
nor U42212 (N_42212,N_38819,N_36844);
nor U42213 (N_42213,N_35785,N_36153);
xnor U42214 (N_42214,N_36726,N_36267);
and U42215 (N_42215,N_35198,N_39801);
xor U42216 (N_42216,N_36435,N_39695);
nand U42217 (N_42217,N_38927,N_36868);
or U42218 (N_42218,N_36182,N_35696);
nand U42219 (N_42219,N_37894,N_36950);
nor U42220 (N_42220,N_35589,N_36245);
nor U42221 (N_42221,N_35385,N_37520);
nand U42222 (N_42222,N_38859,N_35513);
nor U42223 (N_42223,N_39550,N_39096);
or U42224 (N_42224,N_37426,N_38314);
xor U42225 (N_42225,N_36137,N_36587);
or U42226 (N_42226,N_37849,N_38493);
nand U42227 (N_42227,N_35918,N_38816);
xnor U42228 (N_42228,N_35681,N_35896);
xor U42229 (N_42229,N_35956,N_35428);
or U42230 (N_42230,N_39454,N_35290);
and U42231 (N_42231,N_35514,N_36681);
and U42232 (N_42232,N_39327,N_39939);
nand U42233 (N_42233,N_35082,N_38421);
and U42234 (N_42234,N_37028,N_38495);
nand U42235 (N_42235,N_35288,N_39831);
xor U42236 (N_42236,N_38036,N_37179);
nor U42237 (N_42237,N_38939,N_35662);
or U42238 (N_42238,N_36610,N_36883);
nand U42239 (N_42239,N_38203,N_39536);
nand U42240 (N_42240,N_38440,N_39296);
nor U42241 (N_42241,N_37748,N_39953);
or U42242 (N_42242,N_38113,N_37182);
nor U42243 (N_42243,N_38971,N_37131);
nor U42244 (N_42244,N_39780,N_38628);
xor U42245 (N_42245,N_35137,N_36011);
and U42246 (N_42246,N_39725,N_37057);
or U42247 (N_42247,N_39104,N_38728);
or U42248 (N_42248,N_37281,N_39719);
nand U42249 (N_42249,N_37298,N_37448);
or U42250 (N_42250,N_38264,N_38515);
or U42251 (N_42251,N_39622,N_38071);
nand U42252 (N_42252,N_39520,N_35342);
xnor U42253 (N_42253,N_36730,N_36605);
and U42254 (N_42254,N_37151,N_38632);
nor U42255 (N_42255,N_39640,N_39662);
nand U42256 (N_42256,N_39996,N_37363);
nor U42257 (N_42257,N_38489,N_39919);
or U42258 (N_42258,N_37780,N_35742);
and U42259 (N_42259,N_37220,N_39987);
nand U42260 (N_42260,N_35850,N_38325);
nand U42261 (N_42261,N_39271,N_39299);
xnor U42262 (N_42262,N_35859,N_38377);
nand U42263 (N_42263,N_38691,N_36034);
and U42264 (N_42264,N_39458,N_36819);
nand U42265 (N_42265,N_37805,N_36432);
nand U42266 (N_42266,N_35910,N_38319);
or U42267 (N_42267,N_35073,N_39631);
nand U42268 (N_42268,N_38615,N_38918);
nor U42269 (N_42269,N_38347,N_35324);
nor U42270 (N_42270,N_37537,N_37646);
nand U42271 (N_42271,N_37095,N_35114);
or U42272 (N_42272,N_39852,N_35828);
and U42273 (N_42273,N_36118,N_36803);
nand U42274 (N_42274,N_36661,N_38724);
nor U42275 (N_42275,N_35145,N_39260);
nor U42276 (N_42276,N_36756,N_39562);
or U42277 (N_42277,N_36352,N_35304);
nor U42278 (N_42278,N_39503,N_35994);
xnor U42279 (N_42279,N_38874,N_35220);
xor U42280 (N_42280,N_37686,N_37020);
xor U42281 (N_42281,N_35239,N_37938);
or U42282 (N_42282,N_35496,N_36176);
or U42283 (N_42283,N_38358,N_39381);
and U42284 (N_42284,N_36579,N_38110);
and U42285 (N_42285,N_35217,N_36693);
nor U42286 (N_42286,N_37584,N_38654);
nand U42287 (N_42287,N_36396,N_36180);
nor U42288 (N_42288,N_36481,N_38181);
or U42289 (N_42289,N_36308,N_39459);
nand U42290 (N_42290,N_37081,N_38191);
nor U42291 (N_42291,N_39591,N_39068);
xnor U42292 (N_42292,N_39774,N_39922);
nand U42293 (N_42293,N_38231,N_39884);
nor U42294 (N_42294,N_35955,N_39813);
and U42295 (N_42295,N_35709,N_37420);
nand U42296 (N_42296,N_37691,N_36716);
nor U42297 (N_42297,N_35484,N_39885);
xnor U42298 (N_42298,N_35560,N_35314);
nand U42299 (N_42299,N_38350,N_37740);
nand U42300 (N_42300,N_35238,N_36357);
or U42301 (N_42301,N_38835,N_35824);
nor U42302 (N_42302,N_37484,N_38075);
nand U42303 (N_42303,N_35127,N_38845);
xor U42304 (N_42304,N_37206,N_37337);
or U42305 (N_42305,N_39456,N_37754);
xor U42306 (N_42306,N_35268,N_37623);
and U42307 (N_42307,N_39016,N_37488);
nor U42308 (N_42308,N_39480,N_39601);
and U42309 (N_42309,N_39017,N_35883);
and U42310 (N_42310,N_39827,N_37322);
nand U42311 (N_42311,N_38188,N_38671);
or U42312 (N_42312,N_37577,N_36986);
nor U42313 (N_42313,N_35799,N_39921);
nand U42314 (N_42314,N_39836,N_35973);
or U42315 (N_42315,N_36535,N_35396);
or U42316 (N_42316,N_37413,N_37184);
xnor U42317 (N_42317,N_36303,N_35308);
and U42318 (N_42318,N_38195,N_39991);
and U42319 (N_42319,N_39258,N_39393);
or U42320 (N_42320,N_38888,N_35811);
and U42321 (N_42321,N_37044,N_35961);
xor U42322 (N_42322,N_35870,N_35305);
nor U42323 (N_42323,N_36629,N_39023);
nand U42324 (N_42324,N_39481,N_37774);
nand U42325 (N_42325,N_35757,N_37705);
nor U42326 (N_42326,N_37701,N_39792);
and U42327 (N_42327,N_36859,N_37942);
and U42328 (N_42328,N_36524,N_39423);
or U42329 (N_42329,N_36908,N_37483);
nor U42330 (N_42330,N_38484,N_35858);
and U42331 (N_42331,N_38476,N_37216);
xor U42332 (N_42332,N_39871,N_35783);
nor U42333 (N_42333,N_36005,N_39726);
nor U42334 (N_42334,N_36071,N_38283);
nand U42335 (N_42335,N_39073,N_37873);
xor U42336 (N_42336,N_39478,N_39183);
nor U42337 (N_42337,N_36865,N_36919);
nand U42338 (N_42338,N_39712,N_35671);
nand U42339 (N_42339,N_35931,N_36902);
and U42340 (N_42340,N_35826,N_38972);
and U42341 (N_42341,N_36336,N_36765);
or U42342 (N_42342,N_35573,N_38630);
xor U42343 (N_42343,N_39448,N_36659);
xor U42344 (N_42344,N_38085,N_39115);
or U42345 (N_42345,N_39027,N_36609);
and U42346 (N_42346,N_35561,N_37139);
or U42347 (N_42347,N_36294,N_39663);
nand U42348 (N_42348,N_38902,N_35568);
and U42349 (N_42349,N_36528,N_39992);
and U42350 (N_42350,N_39164,N_35907);
nor U42351 (N_42351,N_35351,N_37276);
nand U42352 (N_42352,N_38300,N_35042);
or U42353 (N_42353,N_39888,N_39058);
or U42354 (N_42354,N_38151,N_37645);
or U42355 (N_42355,N_35352,N_36121);
or U42356 (N_42356,N_36568,N_37973);
and U42357 (N_42357,N_37581,N_36199);
and U42358 (N_42358,N_35786,N_35079);
and U42359 (N_42359,N_37596,N_35436);
and U42360 (N_42360,N_37574,N_35093);
xnor U42361 (N_42361,N_37120,N_35205);
nor U42362 (N_42362,N_38587,N_38661);
nand U42363 (N_42363,N_39761,N_38468);
nor U42364 (N_42364,N_35444,N_36613);
xor U42365 (N_42365,N_35398,N_37449);
and U42366 (N_42366,N_37724,N_36675);
or U42367 (N_42367,N_35612,N_36811);
xor U42368 (N_42368,N_37273,N_35321);
or U42369 (N_42369,N_36315,N_39958);
xnor U42370 (N_42370,N_37864,N_37271);
or U42371 (N_42371,N_35515,N_39701);
xor U42372 (N_42372,N_39501,N_39855);
and U42373 (N_42373,N_39114,N_35714);
nand U42374 (N_42374,N_35422,N_37733);
nor U42375 (N_42375,N_35812,N_38112);
or U42376 (N_42376,N_35552,N_37799);
nand U42377 (N_42377,N_38975,N_39251);
or U42378 (N_42378,N_35225,N_39413);
or U42379 (N_42379,N_38964,N_38128);
or U42380 (N_42380,N_35236,N_35815);
and U42381 (N_42381,N_38303,N_36288);
xor U42382 (N_42382,N_36968,N_37362);
nand U42383 (N_42383,N_35418,N_36367);
nand U42384 (N_42384,N_39572,N_38327);
and U42385 (N_42385,N_39277,N_37801);
nor U42386 (N_42386,N_39008,N_36151);
or U42387 (N_42387,N_39196,N_36298);
or U42388 (N_42388,N_35584,N_38863);
nor U42389 (N_42389,N_35060,N_39838);
or U42390 (N_42390,N_38477,N_36026);
nand U42391 (N_42391,N_35279,N_37875);
and U42392 (N_42392,N_38896,N_38901);
nand U42393 (N_42393,N_37688,N_35558);
and U42394 (N_42394,N_39209,N_35234);
nand U42395 (N_42395,N_39147,N_39491);
nor U42396 (N_42396,N_37000,N_36496);
nor U42397 (N_42397,N_38153,N_36219);
xnor U42398 (N_42398,N_39007,N_36550);
nand U42399 (N_42399,N_37499,N_37928);
or U42400 (N_42400,N_35185,N_39554);
nand U42401 (N_42401,N_39606,N_35669);
or U42402 (N_42402,N_36920,N_38102);
or U42403 (N_42403,N_39954,N_37090);
and U42404 (N_42404,N_35738,N_38465);
xnor U42405 (N_42405,N_38836,N_37515);
nor U42406 (N_42406,N_37339,N_35974);
nand U42407 (N_42407,N_39123,N_39596);
and U42408 (N_42408,N_37228,N_37910);
and U42409 (N_42409,N_38706,N_38768);
nor U42410 (N_42410,N_39942,N_37392);
and U42411 (N_42411,N_38357,N_37811);
nor U42412 (N_42412,N_35642,N_38490);
or U42413 (N_42413,N_35906,N_39272);
nor U42414 (N_42414,N_37069,N_39990);
or U42415 (N_42415,N_38516,N_35190);
and U42416 (N_42416,N_37078,N_39420);
nand U42417 (N_42417,N_35031,N_36334);
nand U42418 (N_42418,N_39022,N_37843);
or U42419 (N_42419,N_39476,N_37587);
nand U42420 (N_42420,N_36828,N_35649);
or U42421 (N_42421,N_35698,N_39067);
or U42422 (N_42422,N_36429,N_36340);
xor U42423 (N_42423,N_39397,N_35606);
or U42424 (N_42424,N_38210,N_36221);
nor U42425 (N_42425,N_38454,N_38740);
xor U42426 (N_42426,N_35968,N_39034);
xor U42427 (N_42427,N_39334,N_39223);
or U42428 (N_42428,N_39683,N_35375);
xor U42429 (N_42429,N_37719,N_35200);
or U42430 (N_42430,N_39025,N_37716);
or U42431 (N_42431,N_35819,N_35703);
and U42432 (N_42432,N_36988,N_35731);
xnor U42433 (N_42433,N_36602,N_37863);
nand U42434 (N_42434,N_36781,N_36943);
or U42435 (N_42435,N_37275,N_37779);
nor U42436 (N_42436,N_36443,N_35840);
and U42437 (N_42437,N_39833,N_35152);
nand U42438 (N_42438,N_39796,N_39171);
nor U42439 (N_42439,N_38459,N_36249);
nand U42440 (N_42440,N_39738,N_36307);
nand U42441 (N_42441,N_37542,N_39266);
nor U42442 (N_42442,N_36682,N_38529);
nor U42443 (N_42443,N_39446,N_37947);
nand U42444 (N_42444,N_38786,N_36621);
nand U42445 (N_42445,N_38033,N_35798);
nor U42446 (N_42446,N_38886,N_38555);
nor U42447 (N_42447,N_36878,N_38913);
nor U42448 (N_42448,N_35062,N_35412);
nand U42449 (N_42449,N_36126,N_35335);
nor U42450 (N_42450,N_37007,N_38449);
nor U42451 (N_42451,N_35286,N_38701);
and U42452 (N_42452,N_36701,N_37949);
xnor U42453 (N_42453,N_39779,N_36184);
and U42454 (N_42454,N_38385,N_38758);
nor U42455 (N_42455,N_38198,N_37827);
and U42456 (N_42456,N_35770,N_39949);
nand U42457 (N_42457,N_35971,N_38531);
and U42458 (N_42458,N_38641,N_37122);
and U42459 (N_42459,N_35822,N_38963);
nand U42460 (N_42460,N_39527,N_37798);
nand U42461 (N_42461,N_35553,N_37378);
nor U42462 (N_42462,N_37358,N_35653);
nand U42463 (N_42463,N_39993,N_39282);
or U42464 (N_42464,N_39908,N_38002);
and U42465 (N_42465,N_37986,N_38779);
nor U42466 (N_42466,N_35948,N_36423);
or U42467 (N_42467,N_39876,N_37463);
or U42468 (N_42468,N_36710,N_35472);
nand U42469 (N_42469,N_36805,N_39154);
and U42470 (N_42470,N_36141,N_39890);
or U42471 (N_42471,N_36880,N_37388);
and U42472 (N_42472,N_39090,N_36671);
nand U42473 (N_42473,N_38878,N_35520);
or U42474 (N_42474,N_35001,N_38196);
nor U42475 (N_42475,N_37908,N_36183);
xor U42476 (N_42476,N_35368,N_37313);
and U42477 (N_42477,N_38039,N_36098);
or U42478 (N_42478,N_38120,N_38759);
xnor U42479 (N_42479,N_36371,N_38063);
and U42480 (N_42480,N_38953,N_37685);
and U42481 (N_42481,N_37940,N_39489);
or U42482 (N_42482,N_38086,N_35011);
nor U42483 (N_42483,N_35773,N_35817);
nand U42484 (N_42484,N_36766,N_38450);
and U42485 (N_42485,N_39714,N_39583);
nand U42486 (N_42486,N_36017,N_39597);
and U42487 (N_42487,N_38418,N_37255);
nor U42488 (N_42488,N_36537,N_35476);
xor U42489 (N_42489,N_39671,N_36938);
nand U42490 (N_42490,N_35032,N_39131);
and U42491 (N_42491,N_37140,N_39368);
nand U42492 (N_42492,N_38915,N_38690);
or U42493 (N_42493,N_37381,N_37579);
nor U42494 (N_42494,N_36560,N_38242);
and U42495 (N_42495,N_38565,N_35547);
and U42496 (N_42496,N_35985,N_36523);
nand U42497 (N_42497,N_38619,N_35083);
xor U42498 (N_42498,N_39378,N_37556);
nand U42499 (N_42499,N_36694,N_37546);
and U42500 (N_42500,N_39971,N_38718);
nand U42501 (N_42501,N_35906,N_39694);
xor U42502 (N_42502,N_39461,N_36325);
nor U42503 (N_42503,N_38737,N_39256);
and U42504 (N_42504,N_37930,N_35297);
or U42505 (N_42505,N_36855,N_37653);
xnor U42506 (N_42506,N_35921,N_36774);
xnor U42507 (N_42507,N_38139,N_39468);
nor U42508 (N_42508,N_39745,N_37573);
or U42509 (N_42509,N_36021,N_39699);
xnor U42510 (N_42510,N_35115,N_36057);
and U42511 (N_42511,N_39268,N_36903);
or U42512 (N_42512,N_38284,N_37396);
xnor U42513 (N_42513,N_37009,N_39843);
and U42514 (N_42514,N_38860,N_37388);
nand U42515 (N_42515,N_35466,N_38214);
and U42516 (N_42516,N_39573,N_39486);
and U42517 (N_42517,N_37887,N_35189);
or U42518 (N_42518,N_37802,N_36235);
or U42519 (N_42519,N_38208,N_38699);
nor U42520 (N_42520,N_37527,N_35142);
nor U42521 (N_42521,N_35043,N_36894);
xor U42522 (N_42522,N_38212,N_37245);
xor U42523 (N_42523,N_39398,N_38451);
and U42524 (N_42524,N_39983,N_39615);
nor U42525 (N_42525,N_39304,N_35109);
nand U42526 (N_42526,N_39678,N_39092);
nand U42527 (N_42527,N_38036,N_36212);
xor U42528 (N_42528,N_39826,N_38211);
or U42529 (N_42529,N_37653,N_35956);
or U42530 (N_42530,N_36305,N_38798);
and U42531 (N_42531,N_36770,N_37358);
nor U42532 (N_42532,N_37325,N_38495);
nor U42533 (N_42533,N_35176,N_37182);
or U42534 (N_42534,N_35634,N_35852);
nor U42535 (N_42535,N_38287,N_38268);
or U42536 (N_42536,N_37117,N_39653);
or U42537 (N_42537,N_39123,N_37002);
and U42538 (N_42538,N_37262,N_35888);
and U42539 (N_42539,N_37643,N_37195);
nor U42540 (N_42540,N_38794,N_38827);
nor U42541 (N_42541,N_36765,N_38793);
or U42542 (N_42542,N_36661,N_35650);
or U42543 (N_42543,N_36832,N_35657);
xnor U42544 (N_42544,N_38098,N_36947);
and U42545 (N_42545,N_38087,N_39854);
xnor U42546 (N_42546,N_36216,N_35636);
nor U42547 (N_42547,N_37040,N_35008);
and U42548 (N_42548,N_35207,N_38497);
or U42549 (N_42549,N_39914,N_35729);
xor U42550 (N_42550,N_36545,N_35692);
xor U42551 (N_42551,N_36957,N_35852);
nor U42552 (N_42552,N_38831,N_37602);
and U42553 (N_42553,N_36482,N_35030);
nor U42554 (N_42554,N_38952,N_38306);
xnor U42555 (N_42555,N_35500,N_36572);
and U42556 (N_42556,N_39594,N_39606);
or U42557 (N_42557,N_36713,N_37823);
and U42558 (N_42558,N_38363,N_35015);
nand U42559 (N_42559,N_36718,N_39579);
nand U42560 (N_42560,N_38172,N_37629);
or U42561 (N_42561,N_38818,N_35103);
xor U42562 (N_42562,N_39022,N_39807);
or U42563 (N_42563,N_36299,N_39546);
or U42564 (N_42564,N_38032,N_36235);
nor U42565 (N_42565,N_35015,N_37405);
or U42566 (N_42566,N_39961,N_36954);
nor U42567 (N_42567,N_35490,N_39116);
nor U42568 (N_42568,N_39501,N_39866);
and U42569 (N_42569,N_39062,N_35759);
nand U42570 (N_42570,N_37693,N_37762);
nor U42571 (N_42571,N_39486,N_39653);
nand U42572 (N_42572,N_39107,N_38052);
or U42573 (N_42573,N_36854,N_36298);
or U42574 (N_42574,N_36248,N_37556);
xor U42575 (N_42575,N_38682,N_38409);
and U42576 (N_42576,N_37136,N_35591);
and U42577 (N_42577,N_39459,N_39637);
or U42578 (N_42578,N_39451,N_36310);
or U42579 (N_42579,N_38098,N_37640);
nand U42580 (N_42580,N_39463,N_37894);
nor U42581 (N_42581,N_39581,N_39364);
nor U42582 (N_42582,N_39987,N_37862);
and U42583 (N_42583,N_39274,N_39191);
xor U42584 (N_42584,N_38676,N_36012);
and U42585 (N_42585,N_38957,N_35099);
nor U42586 (N_42586,N_38607,N_35857);
xnor U42587 (N_42587,N_38269,N_37916);
xnor U42588 (N_42588,N_39823,N_38574);
xnor U42589 (N_42589,N_37963,N_37324);
and U42590 (N_42590,N_39096,N_39728);
and U42591 (N_42591,N_36310,N_35893);
nor U42592 (N_42592,N_35421,N_35607);
or U42593 (N_42593,N_35264,N_39047);
or U42594 (N_42594,N_36906,N_36022);
xor U42595 (N_42595,N_39068,N_38588);
xnor U42596 (N_42596,N_37015,N_36160);
and U42597 (N_42597,N_39880,N_35415);
nand U42598 (N_42598,N_35560,N_38410);
and U42599 (N_42599,N_35619,N_39591);
xnor U42600 (N_42600,N_38309,N_37401);
or U42601 (N_42601,N_37244,N_38465);
or U42602 (N_42602,N_35118,N_35773);
nand U42603 (N_42603,N_39411,N_37777);
or U42604 (N_42604,N_38728,N_36373);
or U42605 (N_42605,N_37197,N_35755);
or U42606 (N_42606,N_39695,N_37032);
and U42607 (N_42607,N_38262,N_35329);
nand U42608 (N_42608,N_38334,N_35092);
or U42609 (N_42609,N_37349,N_38000);
nand U42610 (N_42610,N_39267,N_38320);
or U42611 (N_42611,N_37131,N_37747);
or U42612 (N_42612,N_36058,N_39670);
and U42613 (N_42613,N_37383,N_37995);
and U42614 (N_42614,N_38428,N_37198);
nor U42615 (N_42615,N_37468,N_38857);
and U42616 (N_42616,N_35174,N_37256);
nand U42617 (N_42617,N_39891,N_39038);
nand U42618 (N_42618,N_36216,N_39207);
xor U42619 (N_42619,N_38212,N_36622);
nand U42620 (N_42620,N_38267,N_35155);
xor U42621 (N_42621,N_38301,N_39029);
nand U42622 (N_42622,N_38169,N_39453);
and U42623 (N_42623,N_36915,N_37363);
and U42624 (N_42624,N_35043,N_39695);
nor U42625 (N_42625,N_37211,N_35242);
nand U42626 (N_42626,N_35950,N_35254);
nor U42627 (N_42627,N_37154,N_38841);
nand U42628 (N_42628,N_35151,N_38945);
nand U42629 (N_42629,N_38313,N_37655);
nand U42630 (N_42630,N_38799,N_37085);
or U42631 (N_42631,N_35000,N_38296);
and U42632 (N_42632,N_36117,N_38606);
xnor U42633 (N_42633,N_35650,N_39303);
nor U42634 (N_42634,N_39392,N_36479);
nor U42635 (N_42635,N_39843,N_35919);
and U42636 (N_42636,N_37382,N_38558);
or U42637 (N_42637,N_36992,N_35048);
nor U42638 (N_42638,N_38909,N_37619);
nand U42639 (N_42639,N_37553,N_38467);
nand U42640 (N_42640,N_37296,N_36621);
nor U42641 (N_42641,N_35945,N_37755);
and U42642 (N_42642,N_37996,N_36645);
and U42643 (N_42643,N_36567,N_38882);
or U42644 (N_42644,N_36477,N_36327);
nand U42645 (N_42645,N_36185,N_38455);
and U42646 (N_42646,N_36001,N_37977);
and U42647 (N_42647,N_36968,N_35215);
and U42648 (N_42648,N_37938,N_36904);
xor U42649 (N_42649,N_35089,N_36154);
xor U42650 (N_42650,N_36141,N_35910);
or U42651 (N_42651,N_39741,N_37224);
nor U42652 (N_42652,N_35956,N_36173);
nand U42653 (N_42653,N_36337,N_38058);
nand U42654 (N_42654,N_38141,N_37221);
and U42655 (N_42655,N_35967,N_35987);
xnor U42656 (N_42656,N_37347,N_37152);
and U42657 (N_42657,N_39002,N_38110);
nor U42658 (N_42658,N_35762,N_35341);
nor U42659 (N_42659,N_39655,N_36927);
or U42660 (N_42660,N_36555,N_38884);
xor U42661 (N_42661,N_39258,N_37552);
nand U42662 (N_42662,N_39272,N_36650);
nand U42663 (N_42663,N_38691,N_39066);
or U42664 (N_42664,N_37184,N_38070);
or U42665 (N_42665,N_38823,N_39977);
nor U42666 (N_42666,N_36931,N_37555);
and U42667 (N_42667,N_36837,N_36040);
and U42668 (N_42668,N_36719,N_37788);
or U42669 (N_42669,N_35127,N_37361);
nand U42670 (N_42670,N_37923,N_37542);
xor U42671 (N_42671,N_37869,N_37225);
xnor U42672 (N_42672,N_38079,N_38721);
nand U42673 (N_42673,N_38241,N_39321);
xor U42674 (N_42674,N_36754,N_37706);
xnor U42675 (N_42675,N_36741,N_38223);
nor U42676 (N_42676,N_38451,N_36549);
xnor U42677 (N_42677,N_39108,N_38974);
nand U42678 (N_42678,N_36446,N_38105);
or U42679 (N_42679,N_35491,N_37973);
nor U42680 (N_42680,N_39691,N_39709);
or U42681 (N_42681,N_36124,N_38427);
and U42682 (N_42682,N_37743,N_36709);
xor U42683 (N_42683,N_37638,N_36229);
xor U42684 (N_42684,N_36852,N_35110);
or U42685 (N_42685,N_39670,N_38943);
or U42686 (N_42686,N_37893,N_38429);
xnor U42687 (N_42687,N_37468,N_36725);
nand U42688 (N_42688,N_38992,N_35300);
and U42689 (N_42689,N_37930,N_36598);
nor U42690 (N_42690,N_38217,N_39343);
xnor U42691 (N_42691,N_36172,N_38772);
nor U42692 (N_42692,N_36712,N_36072);
nand U42693 (N_42693,N_35934,N_35093);
nand U42694 (N_42694,N_39056,N_37497);
or U42695 (N_42695,N_38231,N_39998);
nor U42696 (N_42696,N_35577,N_35978);
or U42697 (N_42697,N_35868,N_36586);
nand U42698 (N_42698,N_37922,N_36998);
or U42699 (N_42699,N_36156,N_38373);
or U42700 (N_42700,N_36635,N_38976);
and U42701 (N_42701,N_38120,N_39417);
nand U42702 (N_42702,N_39791,N_36398);
nand U42703 (N_42703,N_38307,N_39511);
and U42704 (N_42704,N_37184,N_38744);
or U42705 (N_42705,N_38716,N_36925);
nor U42706 (N_42706,N_38558,N_35552);
nand U42707 (N_42707,N_39599,N_39586);
nand U42708 (N_42708,N_36198,N_36249);
nor U42709 (N_42709,N_35559,N_38769);
nand U42710 (N_42710,N_38604,N_36016);
or U42711 (N_42711,N_37408,N_36352);
or U42712 (N_42712,N_38723,N_35779);
nand U42713 (N_42713,N_38026,N_38551);
nor U42714 (N_42714,N_38375,N_39106);
xor U42715 (N_42715,N_39904,N_36696);
nand U42716 (N_42716,N_35476,N_37454);
nand U42717 (N_42717,N_38968,N_36029);
nand U42718 (N_42718,N_39675,N_37804);
nand U42719 (N_42719,N_35972,N_36706);
xnor U42720 (N_42720,N_39559,N_35424);
or U42721 (N_42721,N_38184,N_39815);
xnor U42722 (N_42722,N_38310,N_37259);
nand U42723 (N_42723,N_37186,N_35300);
or U42724 (N_42724,N_36911,N_37625);
or U42725 (N_42725,N_39506,N_36743);
xor U42726 (N_42726,N_35817,N_37130);
and U42727 (N_42727,N_36952,N_35618);
nor U42728 (N_42728,N_35266,N_36126);
nand U42729 (N_42729,N_37032,N_36047);
or U42730 (N_42730,N_36127,N_39039);
and U42731 (N_42731,N_36715,N_35989);
or U42732 (N_42732,N_38936,N_38035);
nor U42733 (N_42733,N_36177,N_36690);
nand U42734 (N_42734,N_38697,N_37086);
nand U42735 (N_42735,N_35414,N_39952);
and U42736 (N_42736,N_37147,N_38561);
and U42737 (N_42737,N_35466,N_35702);
and U42738 (N_42738,N_37869,N_36216);
nor U42739 (N_42739,N_38555,N_35364);
nor U42740 (N_42740,N_37780,N_36194);
or U42741 (N_42741,N_39228,N_35827);
or U42742 (N_42742,N_39878,N_38811);
and U42743 (N_42743,N_39684,N_37057);
and U42744 (N_42744,N_36942,N_35238);
xor U42745 (N_42745,N_37987,N_35582);
xnor U42746 (N_42746,N_36211,N_37370);
nand U42747 (N_42747,N_37957,N_36829);
nor U42748 (N_42748,N_36053,N_35424);
or U42749 (N_42749,N_36215,N_38777);
xor U42750 (N_42750,N_36254,N_37499);
nor U42751 (N_42751,N_35918,N_39257);
nor U42752 (N_42752,N_35799,N_38975);
xor U42753 (N_42753,N_38608,N_36597);
xor U42754 (N_42754,N_38743,N_36468);
and U42755 (N_42755,N_35003,N_36755);
nor U42756 (N_42756,N_38813,N_38073);
xnor U42757 (N_42757,N_35551,N_37835);
nor U42758 (N_42758,N_38381,N_38610);
nor U42759 (N_42759,N_36475,N_36540);
xor U42760 (N_42760,N_37484,N_38630);
nor U42761 (N_42761,N_39807,N_36466);
or U42762 (N_42762,N_36921,N_38030);
and U42763 (N_42763,N_38297,N_39126);
and U42764 (N_42764,N_39575,N_36629);
nand U42765 (N_42765,N_36025,N_35046);
and U42766 (N_42766,N_36679,N_35166);
or U42767 (N_42767,N_36402,N_36671);
xor U42768 (N_42768,N_38733,N_39906);
nand U42769 (N_42769,N_39556,N_35891);
xor U42770 (N_42770,N_37438,N_36347);
or U42771 (N_42771,N_37767,N_36204);
nor U42772 (N_42772,N_38986,N_39228);
nand U42773 (N_42773,N_35670,N_39372);
and U42774 (N_42774,N_39899,N_37537);
or U42775 (N_42775,N_37532,N_36063);
nand U42776 (N_42776,N_37516,N_37948);
or U42777 (N_42777,N_36993,N_35438);
nor U42778 (N_42778,N_35863,N_38559);
xnor U42779 (N_42779,N_36051,N_37015);
xnor U42780 (N_42780,N_39289,N_39228);
nor U42781 (N_42781,N_39585,N_39702);
nor U42782 (N_42782,N_36430,N_36580);
and U42783 (N_42783,N_39648,N_38938);
and U42784 (N_42784,N_36689,N_38000);
nand U42785 (N_42785,N_38826,N_37719);
or U42786 (N_42786,N_36362,N_38748);
and U42787 (N_42787,N_38530,N_35101);
nand U42788 (N_42788,N_36063,N_37871);
and U42789 (N_42789,N_36894,N_35318);
xnor U42790 (N_42790,N_38303,N_35392);
and U42791 (N_42791,N_37424,N_38552);
xor U42792 (N_42792,N_39199,N_36452);
xor U42793 (N_42793,N_36789,N_36614);
or U42794 (N_42794,N_38428,N_37797);
and U42795 (N_42795,N_38611,N_35944);
and U42796 (N_42796,N_36122,N_39348);
or U42797 (N_42797,N_38227,N_38370);
or U42798 (N_42798,N_37333,N_37464);
nor U42799 (N_42799,N_35595,N_39580);
nor U42800 (N_42800,N_39165,N_36598);
or U42801 (N_42801,N_38490,N_35598);
nand U42802 (N_42802,N_35207,N_37051);
nand U42803 (N_42803,N_35491,N_39222);
xor U42804 (N_42804,N_37860,N_39069);
nor U42805 (N_42805,N_38900,N_35194);
and U42806 (N_42806,N_36292,N_37758);
nor U42807 (N_42807,N_37150,N_39697);
or U42808 (N_42808,N_37039,N_37872);
nor U42809 (N_42809,N_37245,N_37919);
xnor U42810 (N_42810,N_37539,N_38226);
nand U42811 (N_42811,N_37390,N_36639);
or U42812 (N_42812,N_35132,N_39171);
nand U42813 (N_42813,N_36671,N_35914);
and U42814 (N_42814,N_39063,N_38572);
nand U42815 (N_42815,N_38475,N_37293);
xnor U42816 (N_42816,N_39600,N_39278);
nand U42817 (N_42817,N_35263,N_38325);
nand U42818 (N_42818,N_35275,N_39473);
xnor U42819 (N_42819,N_36027,N_35942);
nor U42820 (N_42820,N_38539,N_37837);
nand U42821 (N_42821,N_36241,N_39585);
xnor U42822 (N_42822,N_39210,N_36651);
nor U42823 (N_42823,N_35655,N_35467);
and U42824 (N_42824,N_37382,N_39172);
or U42825 (N_42825,N_36213,N_37021);
and U42826 (N_42826,N_39381,N_36997);
or U42827 (N_42827,N_36781,N_37303);
and U42828 (N_42828,N_38617,N_38805);
nand U42829 (N_42829,N_39426,N_35709);
xnor U42830 (N_42830,N_38792,N_35057);
nor U42831 (N_42831,N_37107,N_35078);
nor U42832 (N_42832,N_36933,N_36546);
or U42833 (N_42833,N_37243,N_37028);
nand U42834 (N_42834,N_38709,N_36954);
or U42835 (N_42835,N_35918,N_39226);
nand U42836 (N_42836,N_38504,N_39935);
nor U42837 (N_42837,N_36065,N_36048);
or U42838 (N_42838,N_38092,N_36032);
nand U42839 (N_42839,N_36045,N_37630);
xor U42840 (N_42840,N_36477,N_37776);
and U42841 (N_42841,N_38675,N_36169);
or U42842 (N_42842,N_35736,N_38284);
and U42843 (N_42843,N_38899,N_38037);
nor U42844 (N_42844,N_37761,N_36090);
and U42845 (N_42845,N_39667,N_39323);
nor U42846 (N_42846,N_37948,N_36328);
xor U42847 (N_42847,N_36097,N_35304);
or U42848 (N_42848,N_37927,N_39050);
and U42849 (N_42849,N_36994,N_37821);
nor U42850 (N_42850,N_39134,N_35393);
nor U42851 (N_42851,N_39378,N_36445);
nand U42852 (N_42852,N_35091,N_38661);
and U42853 (N_42853,N_39554,N_35005);
xnor U42854 (N_42854,N_39516,N_36533);
nor U42855 (N_42855,N_39687,N_38473);
and U42856 (N_42856,N_36130,N_37116);
nand U42857 (N_42857,N_38360,N_38431);
nor U42858 (N_42858,N_37879,N_37833);
nor U42859 (N_42859,N_38779,N_37398);
nand U42860 (N_42860,N_37874,N_35719);
and U42861 (N_42861,N_37394,N_37656);
nand U42862 (N_42862,N_37487,N_36987);
and U42863 (N_42863,N_37121,N_37852);
nor U42864 (N_42864,N_35347,N_39290);
nor U42865 (N_42865,N_36987,N_39263);
and U42866 (N_42866,N_38210,N_35995);
and U42867 (N_42867,N_35172,N_37642);
xor U42868 (N_42868,N_37399,N_35446);
and U42869 (N_42869,N_37278,N_36444);
nor U42870 (N_42870,N_35325,N_39621);
and U42871 (N_42871,N_35997,N_38788);
and U42872 (N_42872,N_35371,N_38061);
or U42873 (N_42873,N_37407,N_35098);
nand U42874 (N_42874,N_36250,N_35134);
and U42875 (N_42875,N_39953,N_39755);
nand U42876 (N_42876,N_35733,N_35919);
or U42877 (N_42877,N_36930,N_37554);
xnor U42878 (N_42878,N_36814,N_36335);
nor U42879 (N_42879,N_39840,N_36129);
nor U42880 (N_42880,N_37353,N_39469);
nand U42881 (N_42881,N_36481,N_36165);
nand U42882 (N_42882,N_36608,N_37645);
nand U42883 (N_42883,N_36319,N_38415);
or U42884 (N_42884,N_37900,N_36666);
nand U42885 (N_42885,N_38694,N_39420);
xor U42886 (N_42886,N_39369,N_35095);
or U42887 (N_42887,N_36650,N_35451);
nor U42888 (N_42888,N_35777,N_35247);
and U42889 (N_42889,N_38898,N_37248);
nand U42890 (N_42890,N_37410,N_39539);
xor U42891 (N_42891,N_37122,N_35515);
xnor U42892 (N_42892,N_37582,N_35190);
or U42893 (N_42893,N_37900,N_38687);
xor U42894 (N_42894,N_38949,N_39413);
and U42895 (N_42895,N_37502,N_38240);
nor U42896 (N_42896,N_39988,N_35928);
or U42897 (N_42897,N_39319,N_38272);
xor U42898 (N_42898,N_35654,N_39373);
and U42899 (N_42899,N_35854,N_38469);
nor U42900 (N_42900,N_35804,N_35090);
or U42901 (N_42901,N_36633,N_36229);
nand U42902 (N_42902,N_35098,N_36700);
xor U42903 (N_42903,N_35394,N_39239);
nor U42904 (N_42904,N_37813,N_37294);
xnor U42905 (N_42905,N_35527,N_35138);
xnor U42906 (N_42906,N_37008,N_36244);
xnor U42907 (N_42907,N_39559,N_37458);
nand U42908 (N_42908,N_36780,N_35480);
nand U42909 (N_42909,N_37842,N_37558);
and U42910 (N_42910,N_35078,N_38395);
and U42911 (N_42911,N_38715,N_37649);
xnor U42912 (N_42912,N_38910,N_37942);
and U42913 (N_42913,N_36028,N_36777);
nand U42914 (N_42914,N_39104,N_38802);
nand U42915 (N_42915,N_35973,N_35500);
or U42916 (N_42916,N_38553,N_35664);
nor U42917 (N_42917,N_39374,N_35467);
nand U42918 (N_42918,N_37169,N_35388);
xnor U42919 (N_42919,N_37118,N_36920);
or U42920 (N_42920,N_35568,N_38618);
nor U42921 (N_42921,N_37630,N_36969);
nor U42922 (N_42922,N_39375,N_35553);
nor U42923 (N_42923,N_37383,N_36201);
xnor U42924 (N_42924,N_39196,N_35915);
xnor U42925 (N_42925,N_36979,N_35031);
nor U42926 (N_42926,N_36265,N_39933);
and U42927 (N_42927,N_39141,N_35412);
and U42928 (N_42928,N_37991,N_39111);
or U42929 (N_42929,N_38484,N_38824);
or U42930 (N_42930,N_38753,N_37213);
or U42931 (N_42931,N_39568,N_38059);
nand U42932 (N_42932,N_37239,N_35682);
and U42933 (N_42933,N_35519,N_38485);
nor U42934 (N_42934,N_35030,N_36973);
or U42935 (N_42935,N_36702,N_39824);
nand U42936 (N_42936,N_37171,N_36860);
xor U42937 (N_42937,N_35337,N_39248);
and U42938 (N_42938,N_37016,N_39979);
nor U42939 (N_42939,N_38639,N_39368);
nand U42940 (N_42940,N_36948,N_35016);
nand U42941 (N_42941,N_35788,N_37809);
and U42942 (N_42942,N_38199,N_39985);
nor U42943 (N_42943,N_36171,N_38138);
and U42944 (N_42944,N_37040,N_36680);
nor U42945 (N_42945,N_36933,N_38177);
and U42946 (N_42946,N_36013,N_39926);
nor U42947 (N_42947,N_38747,N_38864);
nand U42948 (N_42948,N_39333,N_38618);
nor U42949 (N_42949,N_38163,N_35047);
nor U42950 (N_42950,N_39852,N_38550);
nand U42951 (N_42951,N_38548,N_37986);
or U42952 (N_42952,N_35295,N_35075);
and U42953 (N_42953,N_37341,N_38635);
and U42954 (N_42954,N_36926,N_38654);
or U42955 (N_42955,N_36693,N_35973);
nor U42956 (N_42956,N_39617,N_37166);
nand U42957 (N_42957,N_35061,N_39466);
nand U42958 (N_42958,N_36046,N_35059);
or U42959 (N_42959,N_39519,N_35786);
or U42960 (N_42960,N_37088,N_38882);
and U42961 (N_42961,N_36121,N_35869);
or U42962 (N_42962,N_36159,N_38627);
and U42963 (N_42963,N_35438,N_38131);
nor U42964 (N_42964,N_37000,N_35223);
or U42965 (N_42965,N_36082,N_35771);
and U42966 (N_42966,N_37328,N_39064);
and U42967 (N_42967,N_36851,N_37776);
or U42968 (N_42968,N_38688,N_36156);
nor U42969 (N_42969,N_38609,N_37356);
and U42970 (N_42970,N_35401,N_35890);
xnor U42971 (N_42971,N_35959,N_36784);
nor U42972 (N_42972,N_35649,N_36942);
or U42973 (N_42973,N_35357,N_35431);
xnor U42974 (N_42974,N_36807,N_37623);
nor U42975 (N_42975,N_38202,N_37310);
nand U42976 (N_42976,N_38709,N_35810);
nor U42977 (N_42977,N_39315,N_39004);
xnor U42978 (N_42978,N_36659,N_39554);
and U42979 (N_42979,N_37937,N_39974);
and U42980 (N_42980,N_35038,N_35742);
or U42981 (N_42981,N_38311,N_35001);
nand U42982 (N_42982,N_39704,N_39241);
nand U42983 (N_42983,N_36251,N_38804);
nor U42984 (N_42984,N_37459,N_35362);
nor U42985 (N_42985,N_37006,N_38353);
and U42986 (N_42986,N_37709,N_37350);
or U42987 (N_42987,N_36305,N_35958);
and U42988 (N_42988,N_38625,N_37265);
nor U42989 (N_42989,N_38451,N_39729);
nor U42990 (N_42990,N_36123,N_35820);
xnor U42991 (N_42991,N_39742,N_38497);
or U42992 (N_42992,N_39315,N_38591);
nor U42993 (N_42993,N_38148,N_39308);
nand U42994 (N_42994,N_37435,N_39623);
or U42995 (N_42995,N_38892,N_35235);
nand U42996 (N_42996,N_38143,N_37740);
nor U42997 (N_42997,N_39167,N_37367);
xnor U42998 (N_42998,N_39023,N_37450);
xor U42999 (N_42999,N_36650,N_36452);
and U43000 (N_43000,N_39439,N_39232);
or U43001 (N_43001,N_35990,N_36635);
or U43002 (N_43002,N_37775,N_37079);
nand U43003 (N_43003,N_38276,N_37165);
nand U43004 (N_43004,N_39424,N_36265);
nand U43005 (N_43005,N_35525,N_36664);
and U43006 (N_43006,N_39501,N_37583);
or U43007 (N_43007,N_39994,N_38574);
and U43008 (N_43008,N_37830,N_39823);
or U43009 (N_43009,N_37268,N_37778);
or U43010 (N_43010,N_39729,N_39252);
and U43011 (N_43011,N_35788,N_36962);
nor U43012 (N_43012,N_37892,N_38821);
and U43013 (N_43013,N_37728,N_36369);
and U43014 (N_43014,N_38528,N_35446);
or U43015 (N_43015,N_39144,N_37375);
and U43016 (N_43016,N_39394,N_36754);
or U43017 (N_43017,N_37879,N_35475);
or U43018 (N_43018,N_38103,N_37880);
or U43019 (N_43019,N_36195,N_35953);
nand U43020 (N_43020,N_38793,N_36135);
nor U43021 (N_43021,N_35583,N_35886);
or U43022 (N_43022,N_38067,N_35155);
nor U43023 (N_43023,N_37133,N_36165);
and U43024 (N_43024,N_36613,N_36714);
xnor U43025 (N_43025,N_37648,N_35308);
or U43026 (N_43026,N_39312,N_35998);
and U43027 (N_43027,N_36574,N_39182);
and U43028 (N_43028,N_37845,N_39846);
xor U43029 (N_43029,N_36200,N_37751);
nor U43030 (N_43030,N_37232,N_35712);
or U43031 (N_43031,N_39657,N_36132);
and U43032 (N_43032,N_35991,N_35467);
xnor U43033 (N_43033,N_39935,N_36330);
xor U43034 (N_43034,N_38304,N_38689);
nor U43035 (N_43035,N_35876,N_39408);
xnor U43036 (N_43036,N_36488,N_36680);
nand U43037 (N_43037,N_38023,N_37859);
nor U43038 (N_43038,N_38942,N_39473);
nor U43039 (N_43039,N_35166,N_37125);
nor U43040 (N_43040,N_35886,N_36718);
xnor U43041 (N_43041,N_37823,N_35519);
nor U43042 (N_43042,N_38000,N_37242);
nand U43043 (N_43043,N_36615,N_37586);
nand U43044 (N_43044,N_35606,N_36018);
xor U43045 (N_43045,N_36746,N_38694);
and U43046 (N_43046,N_37851,N_38021);
and U43047 (N_43047,N_38421,N_39690);
xor U43048 (N_43048,N_37653,N_36466);
nor U43049 (N_43049,N_36309,N_39257);
nor U43050 (N_43050,N_36042,N_36037);
xnor U43051 (N_43051,N_39947,N_38333);
nand U43052 (N_43052,N_39691,N_35882);
nor U43053 (N_43053,N_35068,N_35242);
or U43054 (N_43054,N_35585,N_38388);
nor U43055 (N_43055,N_36841,N_38890);
nand U43056 (N_43056,N_37863,N_38856);
nor U43057 (N_43057,N_36715,N_35495);
and U43058 (N_43058,N_36693,N_38506);
nor U43059 (N_43059,N_38655,N_35520);
xnor U43060 (N_43060,N_37326,N_35603);
xor U43061 (N_43061,N_39516,N_35336);
nor U43062 (N_43062,N_39866,N_37045);
nor U43063 (N_43063,N_39545,N_36746);
xnor U43064 (N_43064,N_37482,N_37390);
or U43065 (N_43065,N_38079,N_39277);
xor U43066 (N_43066,N_36017,N_37988);
nor U43067 (N_43067,N_36812,N_38126);
nor U43068 (N_43068,N_37347,N_35958);
xor U43069 (N_43069,N_39953,N_36395);
nand U43070 (N_43070,N_39953,N_37193);
xor U43071 (N_43071,N_39075,N_38877);
xor U43072 (N_43072,N_36381,N_38145);
or U43073 (N_43073,N_35380,N_37007);
and U43074 (N_43074,N_37883,N_39247);
nor U43075 (N_43075,N_39486,N_35242);
nand U43076 (N_43076,N_38484,N_38926);
or U43077 (N_43077,N_38126,N_35773);
xnor U43078 (N_43078,N_36190,N_37680);
nor U43079 (N_43079,N_39124,N_37903);
nor U43080 (N_43080,N_36503,N_35449);
nand U43081 (N_43081,N_38336,N_39951);
and U43082 (N_43082,N_38724,N_39200);
or U43083 (N_43083,N_38889,N_38046);
nor U43084 (N_43084,N_38174,N_36847);
nand U43085 (N_43085,N_37652,N_38237);
or U43086 (N_43086,N_35885,N_36165);
or U43087 (N_43087,N_38710,N_36667);
nand U43088 (N_43088,N_36568,N_37617);
nand U43089 (N_43089,N_36546,N_38758);
xnor U43090 (N_43090,N_39298,N_36994);
nor U43091 (N_43091,N_35517,N_39631);
nand U43092 (N_43092,N_37497,N_39793);
and U43093 (N_43093,N_35123,N_36671);
nor U43094 (N_43094,N_37586,N_38178);
nor U43095 (N_43095,N_37872,N_35089);
and U43096 (N_43096,N_37144,N_39438);
nor U43097 (N_43097,N_36086,N_39674);
or U43098 (N_43098,N_37156,N_39412);
nor U43099 (N_43099,N_36554,N_38510);
xnor U43100 (N_43100,N_39315,N_35655);
xnor U43101 (N_43101,N_36873,N_39467);
and U43102 (N_43102,N_38900,N_36112);
xnor U43103 (N_43103,N_35629,N_35797);
xnor U43104 (N_43104,N_36313,N_38432);
nor U43105 (N_43105,N_37810,N_36499);
xnor U43106 (N_43106,N_35485,N_39529);
nand U43107 (N_43107,N_37528,N_37447);
nand U43108 (N_43108,N_38739,N_35298);
or U43109 (N_43109,N_39754,N_38245);
xnor U43110 (N_43110,N_37443,N_39908);
xnor U43111 (N_43111,N_37763,N_38824);
xor U43112 (N_43112,N_37230,N_35494);
or U43113 (N_43113,N_35993,N_39163);
nor U43114 (N_43114,N_35011,N_36881);
nor U43115 (N_43115,N_37397,N_35889);
nand U43116 (N_43116,N_39201,N_38727);
nand U43117 (N_43117,N_36192,N_39402);
nand U43118 (N_43118,N_35674,N_39388);
nand U43119 (N_43119,N_35945,N_37988);
and U43120 (N_43120,N_35359,N_38720);
nand U43121 (N_43121,N_37084,N_38100);
and U43122 (N_43122,N_39229,N_36668);
or U43123 (N_43123,N_35825,N_39824);
or U43124 (N_43124,N_36582,N_39684);
nand U43125 (N_43125,N_35260,N_37288);
and U43126 (N_43126,N_35046,N_39715);
nor U43127 (N_43127,N_38746,N_35397);
xor U43128 (N_43128,N_35928,N_36355);
or U43129 (N_43129,N_37627,N_37906);
nor U43130 (N_43130,N_38226,N_37139);
nor U43131 (N_43131,N_39370,N_36740);
or U43132 (N_43132,N_39730,N_37090);
and U43133 (N_43133,N_39362,N_38973);
xor U43134 (N_43134,N_39218,N_36027);
nand U43135 (N_43135,N_37509,N_37401);
nand U43136 (N_43136,N_37806,N_39643);
or U43137 (N_43137,N_39010,N_38565);
or U43138 (N_43138,N_35276,N_38110);
and U43139 (N_43139,N_39591,N_37114);
or U43140 (N_43140,N_39769,N_39122);
or U43141 (N_43141,N_36450,N_35993);
and U43142 (N_43142,N_38345,N_39882);
or U43143 (N_43143,N_35570,N_37932);
or U43144 (N_43144,N_39538,N_39464);
and U43145 (N_43145,N_38657,N_37333);
nand U43146 (N_43146,N_35642,N_37931);
nor U43147 (N_43147,N_36103,N_38862);
or U43148 (N_43148,N_38307,N_35517);
nor U43149 (N_43149,N_37785,N_36619);
or U43150 (N_43150,N_35145,N_37000);
and U43151 (N_43151,N_35830,N_37188);
and U43152 (N_43152,N_37040,N_37448);
nand U43153 (N_43153,N_37720,N_37557);
and U43154 (N_43154,N_35002,N_39410);
xor U43155 (N_43155,N_38264,N_38612);
xnor U43156 (N_43156,N_39406,N_36144);
and U43157 (N_43157,N_39168,N_38919);
and U43158 (N_43158,N_36928,N_36825);
nor U43159 (N_43159,N_37398,N_35744);
xor U43160 (N_43160,N_39296,N_37142);
or U43161 (N_43161,N_38481,N_36753);
and U43162 (N_43162,N_39492,N_35004);
nand U43163 (N_43163,N_38557,N_37698);
nor U43164 (N_43164,N_39192,N_39943);
or U43165 (N_43165,N_39839,N_37446);
or U43166 (N_43166,N_36432,N_37981);
nor U43167 (N_43167,N_35962,N_39451);
xor U43168 (N_43168,N_38394,N_38725);
or U43169 (N_43169,N_35128,N_37010);
nand U43170 (N_43170,N_38652,N_37991);
nand U43171 (N_43171,N_39040,N_36041);
nand U43172 (N_43172,N_35033,N_36418);
xnor U43173 (N_43173,N_36409,N_37413);
nor U43174 (N_43174,N_35236,N_39982);
and U43175 (N_43175,N_35025,N_38842);
xor U43176 (N_43176,N_39635,N_37863);
xnor U43177 (N_43177,N_39678,N_37176);
or U43178 (N_43178,N_35750,N_37351);
nor U43179 (N_43179,N_35095,N_37985);
nand U43180 (N_43180,N_39287,N_38195);
xnor U43181 (N_43181,N_39743,N_35800);
nor U43182 (N_43182,N_36782,N_36377);
or U43183 (N_43183,N_35120,N_37106);
nor U43184 (N_43184,N_35762,N_36309);
nor U43185 (N_43185,N_35216,N_35268);
nor U43186 (N_43186,N_36414,N_36381);
xor U43187 (N_43187,N_37119,N_35751);
nand U43188 (N_43188,N_36008,N_39092);
nor U43189 (N_43189,N_36128,N_36961);
nand U43190 (N_43190,N_35310,N_36508);
and U43191 (N_43191,N_39421,N_37941);
nand U43192 (N_43192,N_37351,N_37040);
nor U43193 (N_43193,N_39334,N_35987);
nor U43194 (N_43194,N_39529,N_39850);
xnor U43195 (N_43195,N_38991,N_37787);
nand U43196 (N_43196,N_39334,N_35042);
nor U43197 (N_43197,N_39570,N_36466);
or U43198 (N_43198,N_38257,N_38148);
nor U43199 (N_43199,N_38785,N_35474);
nand U43200 (N_43200,N_38229,N_35502);
nand U43201 (N_43201,N_39180,N_38661);
or U43202 (N_43202,N_39079,N_39686);
nand U43203 (N_43203,N_35764,N_35356);
and U43204 (N_43204,N_38003,N_38152);
nand U43205 (N_43205,N_38147,N_37503);
or U43206 (N_43206,N_39722,N_37634);
or U43207 (N_43207,N_35809,N_36986);
nand U43208 (N_43208,N_36721,N_35234);
and U43209 (N_43209,N_36200,N_37715);
xnor U43210 (N_43210,N_35653,N_36141);
nor U43211 (N_43211,N_35898,N_35909);
and U43212 (N_43212,N_37421,N_38635);
or U43213 (N_43213,N_38017,N_39819);
xor U43214 (N_43214,N_38290,N_39823);
and U43215 (N_43215,N_37173,N_38219);
nand U43216 (N_43216,N_36381,N_38120);
or U43217 (N_43217,N_38041,N_36297);
xor U43218 (N_43218,N_38272,N_39488);
nand U43219 (N_43219,N_35263,N_35856);
and U43220 (N_43220,N_38186,N_38066);
nor U43221 (N_43221,N_38816,N_36626);
nor U43222 (N_43222,N_37515,N_39182);
or U43223 (N_43223,N_39785,N_35710);
nand U43224 (N_43224,N_39565,N_36030);
and U43225 (N_43225,N_37183,N_36440);
xor U43226 (N_43226,N_39050,N_37579);
and U43227 (N_43227,N_37329,N_37893);
and U43228 (N_43228,N_38535,N_38010);
and U43229 (N_43229,N_35598,N_36993);
and U43230 (N_43230,N_36600,N_35728);
nor U43231 (N_43231,N_35336,N_39566);
or U43232 (N_43232,N_37963,N_39100);
and U43233 (N_43233,N_39132,N_37206);
nand U43234 (N_43234,N_37277,N_36103);
xor U43235 (N_43235,N_37085,N_37679);
nor U43236 (N_43236,N_39141,N_37336);
nand U43237 (N_43237,N_35602,N_38265);
and U43238 (N_43238,N_35443,N_35461);
nand U43239 (N_43239,N_35542,N_39474);
and U43240 (N_43240,N_36498,N_39086);
nand U43241 (N_43241,N_38858,N_36118);
and U43242 (N_43242,N_37358,N_36647);
nand U43243 (N_43243,N_39949,N_38953);
nand U43244 (N_43244,N_36556,N_36598);
nand U43245 (N_43245,N_36253,N_35562);
nor U43246 (N_43246,N_39337,N_37801);
and U43247 (N_43247,N_39441,N_38162);
or U43248 (N_43248,N_37237,N_35619);
and U43249 (N_43249,N_35339,N_38720);
nor U43250 (N_43250,N_39778,N_39649);
nor U43251 (N_43251,N_36690,N_39596);
nor U43252 (N_43252,N_35493,N_37267);
nor U43253 (N_43253,N_36543,N_35984);
xor U43254 (N_43254,N_38432,N_35986);
or U43255 (N_43255,N_38303,N_38552);
xor U43256 (N_43256,N_37948,N_35368);
nand U43257 (N_43257,N_35103,N_36508);
xor U43258 (N_43258,N_39264,N_35863);
and U43259 (N_43259,N_37181,N_37355);
xor U43260 (N_43260,N_39759,N_38148);
and U43261 (N_43261,N_36713,N_38684);
xnor U43262 (N_43262,N_39060,N_39597);
xor U43263 (N_43263,N_39904,N_35242);
nor U43264 (N_43264,N_37811,N_39123);
nor U43265 (N_43265,N_39414,N_38323);
or U43266 (N_43266,N_39442,N_35798);
xnor U43267 (N_43267,N_35965,N_35246);
nor U43268 (N_43268,N_35677,N_39300);
xor U43269 (N_43269,N_35859,N_38307);
and U43270 (N_43270,N_36311,N_39137);
xor U43271 (N_43271,N_39647,N_39840);
or U43272 (N_43272,N_35081,N_35206);
xor U43273 (N_43273,N_39162,N_38635);
nand U43274 (N_43274,N_39634,N_37813);
nand U43275 (N_43275,N_36907,N_36417);
xor U43276 (N_43276,N_37001,N_35663);
nor U43277 (N_43277,N_37015,N_36136);
xor U43278 (N_43278,N_38279,N_39613);
nand U43279 (N_43279,N_38125,N_36044);
nor U43280 (N_43280,N_36948,N_39801);
and U43281 (N_43281,N_39453,N_35688);
nor U43282 (N_43282,N_35604,N_35613);
or U43283 (N_43283,N_35784,N_38963);
nor U43284 (N_43284,N_36897,N_36050);
nand U43285 (N_43285,N_38188,N_39864);
and U43286 (N_43286,N_37760,N_37564);
nand U43287 (N_43287,N_37111,N_39868);
xnor U43288 (N_43288,N_35308,N_35561);
nor U43289 (N_43289,N_36258,N_35420);
and U43290 (N_43290,N_38101,N_37917);
or U43291 (N_43291,N_37367,N_37237);
nor U43292 (N_43292,N_35005,N_39953);
nor U43293 (N_43293,N_35656,N_37320);
nand U43294 (N_43294,N_36299,N_36354);
xnor U43295 (N_43295,N_39311,N_39084);
nor U43296 (N_43296,N_37880,N_36765);
nand U43297 (N_43297,N_36320,N_38828);
and U43298 (N_43298,N_36928,N_36828);
xnor U43299 (N_43299,N_36813,N_36173);
xor U43300 (N_43300,N_36261,N_39483);
xor U43301 (N_43301,N_35260,N_36673);
xor U43302 (N_43302,N_37319,N_38753);
nor U43303 (N_43303,N_38371,N_38881);
or U43304 (N_43304,N_37594,N_39563);
xnor U43305 (N_43305,N_36988,N_36392);
and U43306 (N_43306,N_35058,N_38943);
and U43307 (N_43307,N_37658,N_38853);
xnor U43308 (N_43308,N_38193,N_35659);
or U43309 (N_43309,N_37221,N_39391);
or U43310 (N_43310,N_37992,N_39147);
or U43311 (N_43311,N_35776,N_39169);
xnor U43312 (N_43312,N_36322,N_37332);
nor U43313 (N_43313,N_37921,N_36038);
nor U43314 (N_43314,N_35159,N_39215);
nand U43315 (N_43315,N_36778,N_38072);
nor U43316 (N_43316,N_35144,N_36572);
and U43317 (N_43317,N_37489,N_36551);
and U43318 (N_43318,N_37052,N_38331);
nand U43319 (N_43319,N_35455,N_35776);
or U43320 (N_43320,N_36262,N_39970);
or U43321 (N_43321,N_35616,N_36730);
and U43322 (N_43322,N_37328,N_37872);
xor U43323 (N_43323,N_37775,N_38773);
xor U43324 (N_43324,N_38791,N_39827);
and U43325 (N_43325,N_37559,N_39673);
xor U43326 (N_43326,N_37354,N_38518);
nor U43327 (N_43327,N_39920,N_39673);
nand U43328 (N_43328,N_36251,N_39998);
and U43329 (N_43329,N_39210,N_36607);
and U43330 (N_43330,N_35278,N_36911);
nor U43331 (N_43331,N_37388,N_35587);
or U43332 (N_43332,N_38004,N_35984);
xnor U43333 (N_43333,N_38955,N_39434);
nor U43334 (N_43334,N_36276,N_38332);
nand U43335 (N_43335,N_36826,N_39461);
nor U43336 (N_43336,N_36455,N_37954);
nor U43337 (N_43337,N_38959,N_37316);
xnor U43338 (N_43338,N_38197,N_37223);
xnor U43339 (N_43339,N_35880,N_36450);
or U43340 (N_43340,N_38841,N_37860);
xnor U43341 (N_43341,N_36500,N_37756);
nand U43342 (N_43342,N_38552,N_35066);
nand U43343 (N_43343,N_38632,N_39944);
nand U43344 (N_43344,N_37167,N_37302);
or U43345 (N_43345,N_35618,N_39388);
nand U43346 (N_43346,N_37437,N_36648);
nand U43347 (N_43347,N_39764,N_37845);
nor U43348 (N_43348,N_37778,N_35159);
nand U43349 (N_43349,N_35312,N_38105);
or U43350 (N_43350,N_36251,N_39601);
nor U43351 (N_43351,N_37594,N_36578);
and U43352 (N_43352,N_37192,N_35445);
nor U43353 (N_43353,N_35549,N_39611);
xor U43354 (N_43354,N_39392,N_39913);
nor U43355 (N_43355,N_36305,N_35181);
nor U43356 (N_43356,N_37236,N_36533);
nand U43357 (N_43357,N_38144,N_37000);
nand U43358 (N_43358,N_36615,N_35000);
or U43359 (N_43359,N_39072,N_38217);
or U43360 (N_43360,N_38264,N_37029);
or U43361 (N_43361,N_36205,N_39264);
nand U43362 (N_43362,N_35588,N_38817);
and U43363 (N_43363,N_37463,N_38630);
and U43364 (N_43364,N_37748,N_39510);
nor U43365 (N_43365,N_39583,N_35584);
xor U43366 (N_43366,N_36432,N_39216);
nor U43367 (N_43367,N_37113,N_38365);
nor U43368 (N_43368,N_35306,N_36173);
or U43369 (N_43369,N_36796,N_38726);
and U43370 (N_43370,N_36968,N_37783);
and U43371 (N_43371,N_35369,N_38335);
nand U43372 (N_43372,N_39375,N_39352);
or U43373 (N_43373,N_37236,N_35329);
nand U43374 (N_43374,N_37318,N_36316);
or U43375 (N_43375,N_38487,N_36483);
nand U43376 (N_43376,N_36730,N_39281);
nand U43377 (N_43377,N_38078,N_37165);
xor U43378 (N_43378,N_35058,N_36631);
or U43379 (N_43379,N_36040,N_35574);
and U43380 (N_43380,N_38295,N_38656);
xor U43381 (N_43381,N_39289,N_35980);
nand U43382 (N_43382,N_37077,N_37786);
xor U43383 (N_43383,N_39402,N_39581);
nor U43384 (N_43384,N_38041,N_37037);
and U43385 (N_43385,N_36255,N_36783);
or U43386 (N_43386,N_37460,N_38722);
nor U43387 (N_43387,N_36696,N_38824);
nor U43388 (N_43388,N_36628,N_38394);
or U43389 (N_43389,N_38032,N_39325);
nor U43390 (N_43390,N_37093,N_39495);
or U43391 (N_43391,N_37953,N_35785);
nand U43392 (N_43392,N_36102,N_35530);
nor U43393 (N_43393,N_37832,N_36104);
and U43394 (N_43394,N_38713,N_36274);
or U43395 (N_43395,N_39568,N_39150);
and U43396 (N_43396,N_36094,N_35572);
nand U43397 (N_43397,N_38080,N_35084);
nand U43398 (N_43398,N_35445,N_36267);
nor U43399 (N_43399,N_36952,N_37419);
or U43400 (N_43400,N_38945,N_39870);
nand U43401 (N_43401,N_38480,N_37304);
or U43402 (N_43402,N_39377,N_35889);
nor U43403 (N_43403,N_36972,N_38227);
or U43404 (N_43404,N_35770,N_35567);
and U43405 (N_43405,N_35212,N_36139);
nand U43406 (N_43406,N_36730,N_36611);
nor U43407 (N_43407,N_37166,N_39978);
nand U43408 (N_43408,N_38509,N_39616);
and U43409 (N_43409,N_35426,N_39420);
nand U43410 (N_43410,N_35925,N_36877);
xnor U43411 (N_43411,N_39525,N_39219);
or U43412 (N_43412,N_36734,N_38314);
nor U43413 (N_43413,N_37192,N_35941);
and U43414 (N_43414,N_38433,N_38127);
and U43415 (N_43415,N_39767,N_38871);
nand U43416 (N_43416,N_39661,N_38163);
xnor U43417 (N_43417,N_39026,N_36795);
or U43418 (N_43418,N_36725,N_39641);
nand U43419 (N_43419,N_35302,N_35824);
nor U43420 (N_43420,N_35451,N_35220);
xor U43421 (N_43421,N_35485,N_38166);
nor U43422 (N_43422,N_37028,N_39432);
xnor U43423 (N_43423,N_35538,N_39891);
and U43424 (N_43424,N_38994,N_39786);
nand U43425 (N_43425,N_36638,N_35029);
nor U43426 (N_43426,N_35905,N_38621);
and U43427 (N_43427,N_37925,N_37168);
and U43428 (N_43428,N_37123,N_37331);
nor U43429 (N_43429,N_35949,N_39021);
nor U43430 (N_43430,N_37385,N_36578);
or U43431 (N_43431,N_37207,N_37298);
nand U43432 (N_43432,N_37935,N_37610);
nor U43433 (N_43433,N_38957,N_37475);
nand U43434 (N_43434,N_37805,N_37927);
xor U43435 (N_43435,N_35051,N_39501);
or U43436 (N_43436,N_38501,N_38380);
nor U43437 (N_43437,N_37123,N_37223);
or U43438 (N_43438,N_37745,N_39708);
or U43439 (N_43439,N_36841,N_35573);
nor U43440 (N_43440,N_39356,N_36605);
xnor U43441 (N_43441,N_39738,N_35362);
nor U43442 (N_43442,N_39441,N_35510);
or U43443 (N_43443,N_37435,N_36544);
nor U43444 (N_43444,N_35883,N_39820);
nor U43445 (N_43445,N_39994,N_35777);
nand U43446 (N_43446,N_35266,N_35875);
xor U43447 (N_43447,N_39833,N_36696);
nor U43448 (N_43448,N_35112,N_36461);
or U43449 (N_43449,N_39829,N_35658);
nor U43450 (N_43450,N_37355,N_35821);
nor U43451 (N_43451,N_36635,N_37408);
nor U43452 (N_43452,N_36608,N_39211);
nor U43453 (N_43453,N_39343,N_37520);
xnor U43454 (N_43454,N_38918,N_39571);
nand U43455 (N_43455,N_39081,N_39878);
nor U43456 (N_43456,N_36775,N_39815);
nand U43457 (N_43457,N_39129,N_37951);
and U43458 (N_43458,N_35064,N_37253);
and U43459 (N_43459,N_38737,N_38552);
nor U43460 (N_43460,N_38232,N_36689);
nand U43461 (N_43461,N_36819,N_35179);
or U43462 (N_43462,N_36219,N_38003);
nand U43463 (N_43463,N_37221,N_37157);
or U43464 (N_43464,N_38521,N_37378);
and U43465 (N_43465,N_36307,N_38619);
or U43466 (N_43466,N_38887,N_36847);
xor U43467 (N_43467,N_37688,N_36322);
nor U43468 (N_43468,N_36590,N_39827);
and U43469 (N_43469,N_37267,N_36662);
nor U43470 (N_43470,N_37529,N_36346);
xnor U43471 (N_43471,N_36305,N_36546);
and U43472 (N_43472,N_36448,N_36724);
xor U43473 (N_43473,N_35284,N_37825);
or U43474 (N_43474,N_36995,N_35259);
or U43475 (N_43475,N_39955,N_37934);
xnor U43476 (N_43476,N_39782,N_37237);
xor U43477 (N_43477,N_35881,N_35519);
and U43478 (N_43478,N_36689,N_35311);
nand U43479 (N_43479,N_37679,N_35200);
nand U43480 (N_43480,N_38727,N_36827);
and U43481 (N_43481,N_39028,N_39206);
xor U43482 (N_43482,N_38567,N_35807);
or U43483 (N_43483,N_37864,N_38445);
nand U43484 (N_43484,N_36337,N_37639);
xnor U43485 (N_43485,N_38826,N_36404);
nand U43486 (N_43486,N_35363,N_35015);
and U43487 (N_43487,N_37435,N_36432);
or U43488 (N_43488,N_35236,N_39245);
or U43489 (N_43489,N_36615,N_39593);
nor U43490 (N_43490,N_35928,N_35926);
nand U43491 (N_43491,N_39742,N_35653);
and U43492 (N_43492,N_38783,N_38401);
nor U43493 (N_43493,N_38699,N_39660);
and U43494 (N_43494,N_39913,N_37512);
and U43495 (N_43495,N_36655,N_35800);
nand U43496 (N_43496,N_37483,N_39377);
xnor U43497 (N_43497,N_35393,N_39584);
xnor U43498 (N_43498,N_39902,N_35468);
or U43499 (N_43499,N_36693,N_36945);
and U43500 (N_43500,N_35804,N_35015);
nand U43501 (N_43501,N_36094,N_35154);
nor U43502 (N_43502,N_35688,N_39678);
and U43503 (N_43503,N_37258,N_37416);
or U43504 (N_43504,N_39511,N_35131);
nor U43505 (N_43505,N_39234,N_38245);
nand U43506 (N_43506,N_38902,N_39180);
nand U43507 (N_43507,N_37962,N_36386);
nand U43508 (N_43508,N_36780,N_36944);
xor U43509 (N_43509,N_39756,N_39040);
nand U43510 (N_43510,N_39077,N_38392);
nand U43511 (N_43511,N_39112,N_39674);
xnor U43512 (N_43512,N_37111,N_36712);
xnor U43513 (N_43513,N_38379,N_39685);
or U43514 (N_43514,N_36639,N_35779);
and U43515 (N_43515,N_39988,N_39094);
nor U43516 (N_43516,N_35085,N_38095);
xnor U43517 (N_43517,N_39353,N_35928);
nand U43518 (N_43518,N_39921,N_35629);
and U43519 (N_43519,N_36846,N_35560);
and U43520 (N_43520,N_37492,N_37846);
nand U43521 (N_43521,N_37594,N_37640);
and U43522 (N_43522,N_39726,N_38103);
or U43523 (N_43523,N_39100,N_37606);
nand U43524 (N_43524,N_39337,N_37779);
xor U43525 (N_43525,N_35512,N_38713);
nand U43526 (N_43526,N_38665,N_39705);
or U43527 (N_43527,N_36805,N_39993);
nor U43528 (N_43528,N_38436,N_39415);
nand U43529 (N_43529,N_38626,N_39749);
nor U43530 (N_43530,N_39475,N_36346);
nand U43531 (N_43531,N_35991,N_38972);
or U43532 (N_43532,N_39079,N_35094);
nand U43533 (N_43533,N_38230,N_36199);
or U43534 (N_43534,N_38367,N_37257);
nor U43535 (N_43535,N_36694,N_35875);
and U43536 (N_43536,N_37768,N_37229);
and U43537 (N_43537,N_39843,N_39064);
or U43538 (N_43538,N_35184,N_38145);
nor U43539 (N_43539,N_36097,N_38906);
or U43540 (N_43540,N_35457,N_36126);
or U43541 (N_43541,N_37209,N_35263);
nand U43542 (N_43542,N_37652,N_38012);
nor U43543 (N_43543,N_35061,N_37043);
and U43544 (N_43544,N_35389,N_37908);
nor U43545 (N_43545,N_36915,N_39703);
and U43546 (N_43546,N_37177,N_35806);
nand U43547 (N_43547,N_35407,N_37018);
xor U43548 (N_43548,N_35319,N_39536);
nand U43549 (N_43549,N_39775,N_35533);
xnor U43550 (N_43550,N_39793,N_39154);
nor U43551 (N_43551,N_35120,N_37875);
nor U43552 (N_43552,N_39078,N_37907);
nand U43553 (N_43553,N_37410,N_36509);
nor U43554 (N_43554,N_35358,N_38742);
xor U43555 (N_43555,N_39269,N_36291);
or U43556 (N_43556,N_37142,N_36689);
nand U43557 (N_43557,N_35612,N_39610);
or U43558 (N_43558,N_39723,N_39939);
and U43559 (N_43559,N_39258,N_39672);
nor U43560 (N_43560,N_37619,N_39563);
and U43561 (N_43561,N_39505,N_35791);
nor U43562 (N_43562,N_38799,N_36812);
nor U43563 (N_43563,N_38071,N_39056);
and U43564 (N_43564,N_36036,N_36145);
or U43565 (N_43565,N_36580,N_38627);
and U43566 (N_43566,N_37444,N_37583);
xnor U43567 (N_43567,N_37660,N_38147);
xnor U43568 (N_43568,N_39022,N_35518);
nand U43569 (N_43569,N_39683,N_36263);
or U43570 (N_43570,N_35540,N_37043);
and U43571 (N_43571,N_38873,N_35146);
xor U43572 (N_43572,N_36225,N_38127);
nor U43573 (N_43573,N_37778,N_37347);
xor U43574 (N_43574,N_36647,N_38668);
nor U43575 (N_43575,N_37207,N_35585);
xnor U43576 (N_43576,N_37643,N_37211);
xor U43577 (N_43577,N_37681,N_39892);
and U43578 (N_43578,N_38521,N_38968);
or U43579 (N_43579,N_37404,N_38071);
nor U43580 (N_43580,N_37672,N_36774);
or U43581 (N_43581,N_37088,N_35900);
or U43582 (N_43582,N_35156,N_38437);
and U43583 (N_43583,N_35824,N_35712);
nand U43584 (N_43584,N_37062,N_39844);
nand U43585 (N_43585,N_37812,N_35238);
or U43586 (N_43586,N_38771,N_37233);
nor U43587 (N_43587,N_35546,N_37895);
xor U43588 (N_43588,N_39201,N_38425);
xnor U43589 (N_43589,N_39514,N_35114);
or U43590 (N_43590,N_37509,N_39392);
and U43591 (N_43591,N_36307,N_39830);
and U43592 (N_43592,N_35543,N_38379);
nor U43593 (N_43593,N_39742,N_39168);
nor U43594 (N_43594,N_39449,N_35652);
xor U43595 (N_43595,N_36356,N_36206);
nor U43596 (N_43596,N_35249,N_36788);
nor U43597 (N_43597,N_39602,N_38716);
or U43598 (N_43598,N_38139,N_39034);
nand U43599 (N_43599,N_35053,N_39496);
or U43600 (N_43600,N_37285,N_36352);
nor U43601 (N_43601,N_35650,N_39216);
nand U43602 (N_43602,N_38277,N_35800);
xor U43603 (N_43603,N_35437,N_37324);
or U43604 (N_43604,N_38430,N_35221);
xnor U43605 (N_43605,N_39795,N_35511);
nand U43606 (N_43606,N_35161,N_38797);
nand U43607 (N_43607,N_39594,N_38424);
and U43608 (N_43608,N_35468,N_36759);
nor U43609 (N_43609,N_36067,N_37374);
nor U43610 (N_43610,N_37322,N_35275);
and U43611 (N_43611,N_37171,N_38227);
nor U43612 (N_43612,N_39124,N_38161);
xnor U43613 (N_43613,N_37540,N_38623);
xnor U43614 (N_43614,N_37419,N_37431);
and U43615 (N_43615,N_37424,N_35084);
xnor U43616 (N_43616,N_38629,N_35156);
xnor U43617 (N_43617,N_36298,N_36624);
nor U43618 (N_43618,N_39050,N_35980);
nand U43619 (N_43619,N_35016,N_37912);
and U43620 (N_43620,N_39098,N_36644);
or U43621 (N_43621,N_39320,N_38815);
nand U43622 (N_43622,N_35546,N_36124);
xnor U43623 (N_43623,N_37854,N_39859);
nand U43624 (N_43624,N_39360,N_38428);
and U43625 (N_43625,N_38015,N_38869);
xor U43626 (N_43626,N_39616,N_38403);
nor U43627 (N_43627,N_37475,N_35014);
and U43628 (N_43628,N_39325,N_38739);
or U43629 (N_43629,N_35041,N_38947);
nor U43630 (N_43630,N_35704,N_35290);
nand U43631 (N_43631,N_37029,N_37549);
or U43632 (N_43632,N_36358,N_36184);
and U43633 (N_43633,N_35727,N_37013);
xnor U43634 (N_43634,N_36305,N_39946);
xor U43635 (N_43635,N_39122,N_39367);
and U43636 (N_43636,N_37149,N_35688);
and U43637 (N_43637,N_38041,N_38842);
or U43638 (N_43638,N_35160,N_35021);
or U43639 (N_43639,N_36063,N_35161);
and U43640 (N_43640,N_36015,N_39075);
nor U43641 (N_43641,N_37816,N_38923);
or U43642 (N_43642,N_39042,N_38513);
nand U43643 (N_43643,N_38705,N_39456);
xnor U43644 (N_43644,N_38976,N_38014);
nor U43645 (N_43645,N_35805,N_38379);
nor U43646 (N_43646,N_35093,N_38366);
and U43647 (N_43647,N_39194,N_36644);
xnor U43648 (N_43648,N_39772,N_35295);
nor U43649 (N_43649,N_39356,N_39157);
nor U43650 (N_43650,N_36564,N_38656);
and U43651 (N_43651,N_39073,N_39868);
or U43652 (N_43652,N_38381,N_38153);
nand U43653 (N_43653,N_37700,N_35273);
nor U43654 (N_43654,N_38385,N_36379);
or U43655 (N_43655,N_37483,N_36600);
and U43656 (N_43656,N_38826,N_39889);
and U43657 (N_43657,N_37571,N_39749);
nor U43658 (N_43658,N_37377,N_39751);
nor U43659 (N_43659,N_37739,N_38766);
or U43660 (N_43660,N_39491,N_38174);
nand U43661 (N_43661,N_36708,N_36174);
or U43662 (N_43662,N_38887,N_38753);
or U43663 (N_43663,N_38297,N_38018);
nand U43664 (N_43664,N_36217,N_38445);
xnor U43665 (N_43665,N_35183,N_39950);
xnor U43666 (N_43666,N_36181,N_39928);
xor U43667 (N_43667,N_39905,N_35432);
nor U43668 (N_43668,N_37863,N_35951);
xnor U43669 (N_43669,N_35724,N_37228);
or U43670 (N_43670,N_37321,N_37714);
nand U43671 (N_43671,N_38070,N_37933);
or U43672 (N_43672,N_35091,N_39078);
nand U43673 (N_43673,N_35394,N_36440);
or U43674 (N_43674,N_39366,N_35195);
nor U43675 (N_43675,N_37886,N_38623);
xnor U43676 (N_43676,N_36941,N_37189);
xor U43677 (N_43677,N_39951,N_37035);
nand U43678 (N_43678,N_35156,N_36144);
nand U43679 (N_43679,N_36698,N_35506);
and U43680 (N_43680,N_37136,N_36340);
and U43681 (N_43681,N_35828,N_38127);
and U43682 (N_43682,N_38841,N_36027);
xnor U43683 (N_43683,N_38336,N_35826);
and U43684 (N_43684,N_36354,N_35055);
and U43685 (N_43685,N_36407,N_38316);
or U43686 (N_43686,N_37494,N_37295);
or U43687 (N_43687,N_37032,N_38711);
xnor U43688 (N_43688,N_36053,N_37388);
xnor U43689 (N_43689,N_39189,N_36370);
and U43690 (N_43690,N_38511,N_37098);
xnor U43691 (N_43691,N_38770,N_36765);
nand U43692 (N_43692,N_37183,N_39466);
xnor U43693 (N_43693,N_39453,N_39384);
xnor U43694 (N_43694,N_36171,N_35181);
and U43695 (N_43695,N_38200,N_38960);
and U43696 (N_43696,N_39936,N_37872);
and U43697 (N_43697,N_35156,N_39594);
xnor U43698 (N_43698,N_36134,N_39049);
nor U43699 (N_43699,N_36685,N_35952);
nor U43700 (N_43700,N_38250,N_37576);
xor U43701 (N_43701,N_35990,N_39002);
nor U43702 (N_43702,N_37123,N_35538);
and U43703 (N_43703,N_37399,N_37889);
or U43704 (N_43704,N_35074,N_38929);
and U43705 (N_43705,N_39223,N_38229);
or U43706 (N_43706,N_35810,N_36512);
nand U43707 (N_43707,N_39618,N_39195);
nor U43708 (N_43708,N_36387,N_38619);
xor U43709 (N_43709,N_39669,N_36640);
and U43710 (N_43710,N_35377,N_36395);
and U43711 (N_43711,N_38053,N_36619);
xnor U43712 (N_43712,N_35732,N_37457);
or U43713 (N_43713,N_37854,N_36393);
nor U43714 (N_43714,N_35977,N_35145);
xnor U43715 (N_43715,N_36514,N_38197);
or U43716 (N_43716,N_36535,N_39112);
nor U43717 (N_43717,N_35330,N_37825);
or U43718 (N_43718,N_36917,N_39683);
and U43719 (N_43719,N_36711,N_37828);
or U43720 (N_43720,N_36464,N_37401);
nor U43721 (N_43721,N_37262,N_35841);
nand U43722 (N_43722,N_38347,N_38190);
nand U43723 (N_43723,N_35015,N_35146);
xor U43724 (N_43724,N_38381,N_35280);
nor U43725 (N_43725,N_38558,N_38736);
and U43726 (N_43726,N_35101,N_38154);
nand U43727 (N_43727,N_36539,N_39912);
nand U43728 (N_43728,N_39737,N_37930);
xor U43729 (N_43729,N_39893,N_36769);
and U43730 (N_43730,N_36844,N_36585);
nor U43731 (N_43731,N_38428,N_36219);
nor U43732 (N_43732,N_37621,N_38355);
nand U43733 (N_43733,N_37975,N_35630);
nand U43734 (N_43734,N_39152,N_38570);
and U43735 (N_43735,N_35817,N_38991);
and U43736 (N_43736,N_35883,N_38894);
xor U43737 (N_43737,N_35041,N_39954);
or U43738 (N_43738,N_38287,N_38863);
nor U43739 (N_43739,N_38498,N_37513);
nand U43740 (N_43740,N_35069,N_35690);
and U43741 (N_43741,N_36419,N_36989);
nand U43742 (N_43742,N_37694,N_36710);
nand U43743 (N_43743,N_37140,N_37710);
and U43744 (N_43744,N_37102,N_36638);
xnor U43745 (N_43745,N_36632,N_36176);
and U43746 (N_43746,N_35505,N_35725);
nand U43747 (N_43747,N_38658,N_35418);
nand U43748 (N_43748,N_37401,N_38383);
nand U43749 (N_43749,N_39394,N_35137);
xor U43750 (N_43750,N_37756,N_39889);
xnor U43751 (N_43751,N_35375,N_36336);
nor U43752 (N_43752,N_37963,N_36912);
or U43753 (N_43753,N_38389,N_38489);
xor U43754 (N_43754,N_38314,N_37103);
nand U43755 (N_43755,N_37282,N_37587);
and U43756 (N_43756,N_35069,N_37971);
or U43757 (N_43757,N_37468,N_35388);
xnor U43758 (N_43758,N_37602,N_35852);
nor U43759 (N_43759,N_39120,N_39545);
or U43760 (N_43760,N_39282,N_36147);
and U43761 (N_43761,N_36919,N_37800);
nand U43762 (N_43762,N_37429,N_39747);
and U43763 (N_43763,N_36279,N_38010);
or U43764 (N_43764,N_39741,N_36746);
or U43765 (N_43765,N_36383,N_38179);
nor U43766 (N_43766,N_35875,N_36233);
or U43767 (N_43767,N_37583,N_38033);
nor U43768 (N_43768,N_37029,N_35431);
and U43769 (N_43769,N_35674,N_36067);
or U43770 (N_43770,N_35274,N_39895);
and U43771 (N_43771,N_36868,N_35145);
and U43772 (N_43772,N_35115,N_38602);
nand U43773 (N_43773,N_37458,N_38894);
xnor U43774 (N_43774,N_38115,N_35386);
nor U43775 (N_43775,N_35313,N_39673);
nor U43776 (N_43776,N_37025,N_37300);
and U43777 (N_43777,N_39759,N_36176);
nor U43778 (N_43778,N_36643,N_37312);
and U43779 (N_43779,N_39957,N_35132);
and U43780 (N_43780,N_36964,N_35260);
nand U43781 (N_43781,N_35605,N_38178);
or U43782 (N_43782,N_37025,N_38461);
or U43783 (N_43783,N_35605,N_36600);
xor U43784 (N_43784,N_38112,N_37430);
xor U43785 (N_43785,N_39560,N_37991);
nand U43786 (N_43786,N_38302,N_39704);
xor U43787 (N_43787,N_36903,N_36120);
and U43788 (N_43788,N_39679,N_35951);
nor U43789 (N_43789,N_35046,N_39527);
and U43790 (N_43790,N_35840,N_35296);
nand U43791 (N_43791,N_35506,N_39841);
or U43792 (N_43792,N_35522,N_35835);
nand U43793 (N_43793,N_36224,N_39903);
and U43794 (N_43794,N_39248,N_35874);
xnor U43795 (N_43795,N_35309,N_37398);
nand U43796 (N_43796,N_36610,N_39615);
nand U43797 (N_43797,N_35709,N_37986);
and U43798 (N_43798,N_35944,N_37657);
and U43799 (N_43799,N_36101,N_36396);
xor U43800 (N_43800,N_39902,N_37494);
and U43801 (N_43801,N_39627,N_36019);
nand U43802 (N_43802,N_35827,N_36602);
or U43803 (N_43803,N_36020,N_38298);
xnor U43804 (N_43804,N_37764,N_35640);
or U43805 (N_43805,N_35726,N_39843);
or U43806 (N_43806,N_38017,N_39421);
or U43807 (N_43807,N_35437,N_36310);
and U43808 (N_43808,N_36166,N_37139);
and U43809 (N_43809,N_38494,N_39906);
or U43810 (N_43810,N_37665,N_36910);
or U43811 (N_43811,N_39731,N_39009);
nand U43812 (N_43812,N_38525,N_36406);
xnor U43813 (N_43813,N_38522,N_39387);
nor U43814 (N_43814,N_38265,N_39166);
and U43815 (N_43815,N_35538,N_36964);
nor U43816 (N_43816,N_36584,N_37002);
and U43817 (N_43817,N_37981,N_35918);
and U43818 (N_43818,N_36243,N_38684);
or U43819 (N_43819,N_37267,N_39401);
or U43820 (N_43820,N_39320,N_36145);
nor U43821 (N_43821,N_36186,N_39424);
nor U43822 (N_43822,N_35907,N_38270);
nand U43823 (N_43823,N_35706,N_37874);
and U43824 (N_43824,N_36485,N_39523);
nor U43825 (N_43825,N_36567,N_39686);
xor U43826 (N_43826,N_38000,N_36966);
nand U43827 (N_43827,N_39152,N_39431);
or U43828 (N_43828,N_38763,N_35252);
xnor U43829 (N_43829,N_38693,N_36379);
and U43830 (N_43830,N_36731,N_36602);
and U43831 (N_43831,N_37873,N_35195);
nand U43832 (N_43832,N_37624,N_38471);
nand U43833 (N_43833,N_39074,N_37196);
or U43834 (N_43834,N_37056,N_37247);
and U43835 (N_43835,N_37839,N_38499);
or U43836 (N_43836,N_39883,N_38731);
nor U43837 (N_43837,N_35326,N_39131);
xnor U43838 (N_43838,N_38057,N_38754);
and U43839 (N_43839,N_37500,N_38985);
xor U43840 (N_43840,N_38455,N_39162);
or U43841 (N_43841,N_39139,N_37296);
and U43842 (N_43842,N_35623,N_39790);
xnor U43843 (N_43843,N_35079,N_39439);
xor U43844 (N_43844,N_37706,N_37946);
xnor U43845 (N_43845,N_35230,N_36180);
nand U43846 (N_43846,N_37113,N_35854);
and U43847 (N_43847,N_35850,N_35544);
and U43848 (N_43848,N_39779,N_38847);
xor U43849 (N_43849,N_35311,N_39768);
xnor U43850 (N_43850,N_35329,N_35146);
nor U43851 (N_43851,N_39414,N_39987);
and U43852 (N_43852,N_35459,N_37352);
xor U43853 (N_43853,N_38387,N_37987);
nor U43854 (N_43854,N_39741,N_39787);
or U43855 (N_43855,N_35511,N_36547);
and U43856 (N_43856,N_36692,N_35077);
or U43857 (N_43857,N_35085,N_37818);
nor U43858 (N_43858,N_35395,N_35138);
nor U43859 (N_43859,N_35094,N_39576);
nand U43860 (N_43860,N_38468,N_35389);
nor U43861 (N_43861,N_38744,N_37320);
nor U43862 (N_43862,N_39225,N_37364);
or U43863 (N_43863,N_37772,N_37369);
nor U43864 (N_43864,N_39524,N_37674);
and U43865 (N_43865,N_38927,N_39452);
nand U43866 (N_43866,N_39737,N_37363);
and U43867 (N_43867,N_37758,N_36421);
nor U43868 (N_43868,N_35991,N_36290);
nor U43869 (N_43869,N_35425,N_39969);
xnor U43870 (N_43870,N_35386,N_37875);
nor U43871 (N_43871,N_35576,N_36403);
nor U43872 (N_43872,N_35942,N_36134);
nand U43873 (N_43873,N_36836,N_35182);
xnor U43874 (N_43874,N_36291,N_36527);
and U43875 (N_43875,N_39434,N_36759);
xor U43876 (N_43876,N_38879,N_35885);
or U43877 (N_43877,N_38850,N_38321);
nand U43878 (N_43878,N_37427,N_35234);
or U43879 (N_43879,N_35283,N_36222);
nor U43880 (N_43880,N_35157,N_39859);
or U43881 (N_43881,N_39005,N_38956);
nor U43882 (N_43882,N_36840,N_38267);
nand U43883 (N_43883,N_39892,N_37503);
nand U43884 (N_43884,N_35025,N_35960);
xor U43885 (N_43885,N_35565,N_35720);
and U43886 (N_43886,N_36503,N_39999);
xor U43887 (N_43887,N_37450,N_35101);
xor U43888 (N_43888,N_36010,N_35483);
xor U43889 (N_43889,N_38004,N_37667);
xor U43890 (N_43890,N_38961,N_36177);
and U43891 (N_43891,N_39968,N_37280);
or U43892 (N_43892,N_36437,N_36659);
or U43893 (N_43893,N_37819,N_37488);
nor U43894 (N_43894,N_37917,N_39474);
nand U43895 (N_43895,N_38527,N_37591);
nor U43896 (N_43896,N_35461,N_35416);
or U43897 (N_43897,N_38404,N_35129);
and U43898 (N_43898,N_35130,N_37067);
or U43899 (N_43899,N_35947,N_36265);
or U43900 (N_43900,N_39054,N_35570);
or U43901 (N_43901,N_37590,N_36764);
nand U43902 (N_43902,N_36857,N_35015);
or U43903 (N_43903,N_39231,N_39159);
nand U43904 (N_43904,N_37464,N_36802);
nor U43905 (N_43905,N_38287,N_35355);
nor U43906 (N_43906,N_38215,N_39336);
or U43907 (N_43907,N_39088,N_36048);
nor U43908 (N_43908,N_35921,N_38847);
and U43909 (N_43909,N_37675,N_39388);
and U43910 (N_43910,N_35284,N_35840);
nand U43911 (N_43911,N_36490,N_38491);
xor U43912 (N_43912,N_37122,N_36205);
and U43913 (N_43913,N_38557,N_38510);
nor U43914 (N_43914,N_35973,N_39266);
or U43915 (N_43915,N_37527,N_37227);
or U43916 (N_43916,N_39773,N_36433);
and U43917 (N_43917,N_36488,N_37471);
xor U43918 (N_43918,N_38273,N_39305);
nor U43919 (N_43919,N_36973,N_38850);
or U43920 (N_43920,N_38063,N_39915);
nand U43921 (N_43921,N_35718,N_35387);
xnor U43922 (N_43922,N_37055,N_37401);
and U43923 (N_43923,N_37405,N_39712);
xnor U43924 (N_43924,N_36424,N_39443);
or U43925 (N_43925,N_36842,N_36679);
xor U43926 (N_43926,N_37514,N_37794);
and U43927 (N_43927,N_36219,N_37019);
nor U43928 (N_43928,N_38341,N_38479);
or U43929 (N_43929,N_39437,N_38338);
nand U43930 (N_43930,N_36719,N_38790);
nor U43931 (N_43931,N_35485,N_37577);
xor U43932 (N_43932,N_39252,N_39811);
and U43933 (N_43933,N_37313,N_38057);
nor U43934 (N_43934,N_35334,N_38977);
and U43935 (N_43935,N_35136,N_38295);
and U43936 (N_43936,N_37937,N_38557);
nor U43937 (N_43937,N_37142,N_37776);
nand U43938 (N_43938,N_37412,N_38828);
xor U43939 (N_43939,N_35000,N_36986);
nand U43940 (N_43940,N_38237,N_38958);
nand U43941 (N_43941,N_35280,N_39633);
or U43942 (N_43942,N_35578,N_36939);
xor U43943 (N_43943,N_35784,N_39469);
or U43944 (N_43944,N_39228,N_36409);
nand U43945 (N_43945,N_37066,N_35956);
nor U43946 (N_43946,N_38761,N_38198);
nand U43947 (N_43947,N_36022,N_36121);
and U43948 (N_43948,N_39000,N_37907);
nand U43949 (N_43949,N_36152,N_39941);
or U43950 (N_43950,N_39175,N_36902);
and U43951 (N_43951,N_39062,N_37019);
or U43952 (N_43952,N_38645,N_36630);
nor U43953 (N_43953,N_36672,N_37028);
nor U43954 (N_43954,N_35567,N_36390);
nand U43955 (N_43955,N_39549,N_35605);
nor U43956 (N_43956,N_35570,N_35617);
and U43957 (N_43957,N_37781,N_39938);
or U43958 (N_43958,N_38954,N_36556);
nor U43959 (N_43959,N_35373,N_37917);
nand U43960 (N_43960,N_37200,N_39711);
and U43961 (N_43961,N_35407,N_35621);
nand U43962 (N_43962,N_37952,N_35466);
and U43963 (N_43963,N_36113,N_38450);
or U43964 (N_43964,N_39674,N_35145);
nor U43965 (N_43965,N_39712,N_36888);
or U43966 (N_43966,N_37822,N_36713);
or U43967 (N_43967,N_36095,N_35285);
nand U43968 (N_43968,N_35444,N_37445);
or U43969 (N_43969,N_36310,N_37221);
xnor U43970 (N_43970,N_37460,N_37246);
xor U43971 (N_43971,N_37116,N_36847);
nor U43972 (N_43972,N_38198,N_39848);
and U43973 (N_43973,N_36878,N_35288);
or U43974 (N_43974,N_35014,N_37838);
xor U43975 (N_43975,N_36000,N_35760);
nor U43976 (N_43976,N_37251,N_37438);
nor U43977 (N_43977,N_38976,N_35875);
xnor U43978 (N_43978,N_37427,N_35155);
and U43979 (N_43979,N_36261,N_36860);
nand U43980 (N_43980,N_35977,N_37951);
xor U43981 (N_43981,N_36730,N_37562);
or U43982 (N_43982,N_37646,N_37812);
xnor U43983 (N_43983,N_38719,N_38090);
and U43984 (N_43984,N_36676,N_36754);
nor U43985 (N_43985,N_36726,N_39557);
nor U43986 (N_43986,N_39800,N_37158);
or U43987 (N_43987,N_38259,N_37792);
or U43988 (N_43988,N_38311,N_39566);
nand U43989 (N_43989,N_38180,N_37605);
or U43990 (N_43990,N_38517,N_35793);
or U43991 (N_43991,N_35714,N_39652);
and U43992 (N_43992,N_39117,N_39965);
or U43993 (N_43993,N_37643,N_35724);
and U43994 (N_43994,N_35633,N_37271);
nand U43995 (N_43995,N_38969,N_38068);
xnor U43996 (N_43996,N_36644,N_36827);
nand U43997 (N_43997,N_36566,N_39551);
nand U43998 (N_43998,N_35812,N_36843);
nand U43999 (N_43999,N_36978,N_39411);
nor U44000 (N_44000,N_36834,N_39578);
or U44001 (N_44001,N_39872,N_39260);
xor U44002 (N_44002,N_38207,N_35516);
or U44003 (N_44003,N_38993,N_36625);
nand U44004 (N_44004,N_39884,N_38350);
and U44005 (N_44005,N_37661,N_39764);
xnor U44006 (N_44006,N_39508,N_35633);
or U44007 (N_44007,N_35222,N_35536);
and U44008 (N_44008,N_39319,N_38921);
and U44009 (N_44009,N_35550,N_37121);
xnor U44010 (N_44010,N_39505,N_35673);
xor U44011 (N_44011,N_39154,N_35025);
xnor U44012 (N_44012,N_36240,N_36062);
nor U44013 (N_44013,N_38157,N_37897);
and U44014 (N_44014,N_36902,N_36996);
nand U44015 (N_44015,N_37257,N_39835);
and U44016 (N_44016,N_39238,N_36569);
nand U44017 (N_44017,N_36973,N_35506);
or U44018 (N_44018,N_39248,N_35161);
or U44019 (N_44019,N_37648,N_39574);
or U44020 (N_44020,N_35100,N_35299);
and U44021 (N_44021,N_39411,N_35884);
nor U44022 (N_44022,N_38308,N_39349);
or U44023 (N_44023,N_38422,N_38765);
nor U44024 (N_44024,N_38167,N_36992);
nand U44025 (N_44025,N_38705,N_38184);
xor U44026 (N_44026,N_37967,N_38024);
nor U44027 (N_44027,N_35851,N_37655);
nor U44028 (N_44028,N_36532,N_36299);
nand U44029 (N_44029,N_37369,N_35515);
and U44030 (N_44030,N_36845,N_36665);
or U44031 (N_44031,N_39605,N_36871);
or U44032 (N_44032,N_39015,N_39226);
nand U44033 (N_44033,N_36659,N_38113);
and U44034 (N_44034,N_39979,N_39977);
xor U44035 (N_44035,N_35806,N_35032);
or U44036 (N_44036,N_39505,N_35066);
nor U44037 (N_44037,N_39941,N_36692);
or U44038 (N_44038,N_36263,N_36291);
nor U44039 (N_44039,N_38341,N_36801);
and U44040 (N_44040,N_36220,N_38085);
nand U44041 (N_44041,N_39436,N_36551);
nand U44042 (N_44042,N_35284,N_38848);
and U44043 (N_44043,N_38743,N_35899);
and U44044 (N_44044,N_35972,N_39974);
xnor U44045 (N_44045,N_36041,N_35555);
xnor U44046 (N_44046,N_36146,N_38914);
xor U44047 (N_44047,N_35590,N_35030);
and U44048 (N_44048,N_39408,N_39361);
nor U44049 (N_44049,N_35284,N_36863);
or U44050 (N_44050,N_37309,N_39665);
xor U44051 (N_44051,N_37643,N_39397);
or U44052 (N_44052,N_38793,N_35807);
or U44053 (N_44053,N_37446,N_35875);
and U44054 (N_44054,N_36836,N_39624);
or U44055 (N_44055,N_39548,N_37219);
nand U44056 (N_44056,N_35067,N_39534);
nand U44057 (N_44057,N_38562,N_36999);
xor U44058 (N_44058,N_38472,N_37403);
nor U44059 (N_44059,N_36598,N_37818);
xnor U44060 (N_44060,N_35111,N_35531);
and U44061 (N_44061,N_37257,N_37922);
xnor U44062 (N_44062,N_38561,N_35734);
and U44063 (N_44063,N_36298,N_36493);
or U44064 (N_44064,N_35505,N_39589);
xor U44065 (N_44065,N_38301,N_38887);
nor U44066 (N_44066,N_35038,N_36852);
or U44067 (N_44067,N_38161,N_37818);
or U44068 (N_44068,N_39585,N_38145);
nand U44069 (N_44069,N_36156,N_37590);
or U44070 (N_44070,N_35272,N_39632);
and U44071 (N_44071,N_38544,N_38399);
xor U44072 (N_44072,N_38480,N_37173);
and U44073 (N_44073,N_37826,N_37774);
nor U44074 (N_44074,N_39242,N_35888);
nand U44075 (N_44075,N_35395,N_37326);
and U44076 (N_44076,N_35914,N_39394);
xor U44077 (N_44077,N_36581,N_35503);
nor U44078 (N_44078,N_35254,N_36205);
and U44079 (N_44079,N_39568,N_35150);
nand U44080 (N_44080,N_35489,N_37186);
nand U44081 (N_44081,N_36244,N_36134);
and U44082 (N_44082,N_35739,N_38476);
or U44083 (N_44083,N_36868,N_38941);
and U44084 (N_44084,N_37845,N_35922);
xor U44085 (N_44085,N_36980,N_37190);
xor U44086 (N_44086,N_37373,N_36008);
xor U44087 (N_44087,N_36010,N_39107);
or U44088 (N_44088,N_35732,N_36382);
nand U44089 (N_44089,N_37970,N_35049);
or U44090 (N_44090,N_35616,N_35690);
xor U44091 (N_44091,N_38926,N_39244);
xnor U44092 (N_44092,N_38280,N_37934);
xnor U44093 (N_44093,N_38874,N_39415);
xor U44094 (N_44094,N_36115,N_39288);
nand U44095 (N_44095,N_39986,N_35131);
and U44096 (N_44096,N_38453,N_36416);
or U44097 (N_44097,N_39845,N_37357);
nand U44098 (N_44098,N_36510,N_35091);
nand U44099 (N_44099,N_35520,N_37220);
and U44100 (N_44100,N_39199,N_39898);
or U44101 (N_44101,N_36162,N_38853);
xnor U44102 (N_44102,N_37258,N_38522);
xnor U44103 (N_44103,N_38311,N_39763);
nor U44104 (N_44104,N_36155,N_36897);
or U44105 (N_44105,N_36486,N_36647);
and U44106 (N_44106,N_36691,N_38529);
nor U44107 (N_44107,N_36777,N_39896);
or U44108 (N_44108,N_37502,N_35895);
nor U44109 (N_44109,N_38080,N_35146);
nand U44110 (N_44110,N_37927,N_39385);
and U44111 (N_44111,N_39149,N_38161);
nand U44112 (N_44112,N_37190,N_39821);
xnor U44113 (N_44113,N_37096,N_39879);
nor U44114 (N_44114,N_37517,N_37109);
or U44115 (N_44115,N_36443,N_37409);
nor U44116 (N_44116,N_39201,N_36201);
and U44117 (N_44117,N_38090,N_38259);
nand U44118 (N_44118,N_39684,N_38733);
xor U44119 (N_44119,N_39731,N_38336);
xor U44120 (N_44120,N_35810,N_38486);
nor U44121 (N_44121,N_35360,N_37110);
and U44122 (N_44122,N_35549,N_37078);
nor U44123 (N_44123,N_37661,N_35049);
nor U44124 (N_44124,N_38173,N_39167);
nand U44125 (N_44125,N_39957,N_38492);
and U44126 (N_44126,N_39831,N_35080);
nand U44127 (N_44127,N_37087,N_37202);
or U44128 (N_44128,N_37401,N_38140);
or U44129 (N_44129,N_39809,N_39408);
and U44130 (N_44130,N_38860,N_38835);
nand U44131 (N_44131,N_38805,N_37164);
nand U44132 (N_44132,N_35279,N_39407);
nor U44133 (N_44133,N_35195,N_39536);
or U44134 (N_44134,N_36499,N_35029);
nor U44135 (N_44135,N_39061,N_36856);
nand U44136 (N_44136,N_37036,N_36806);
or U44137 (N_44137,N_37000,N_39622);
nand U44138 (N_44138,N_35943,N_39881);
and U44139 (N_44139,N_36733,N_37994);
and U44140 (N_44140,N_39504,N_37189);
nand U44141 (N_44141,N_39056,N_38462);
and U44142 (N_44142,N_35160,N_37666);
xor U44143 (N_44143,N_37961,N_35216);
and U44144 (N_44144,N_39194,N_38001);
and U44145 (N_44145,N_35097,N_36096);
and U44146 (N_44146,N_36076,N_39246);
xnor U44147 (N_44147,N_39837,N_38566);
nand U44148 (N_44148,N_37272,N_36683);
xnor U44149 (N_44149,N_37707,N_39806);
nand U44150 (N_44150,N_35532,N_38866);
nand U44151 (N_44151,N_35837,N_35146);
and U44152 (N_44152,N_38749,N_36212);
or U44153 (N_44153,N_38152,N_39986);
or U44154 (N_44154,N_38291,N_38956);
xnor U44155 (N_44155,N_35249,N_35757);
and U44156 (N_44156,N_37499,N_39221);
and U44157 (N_44157,N_37622,N_37690);
xnor U44158 (N_44158,N_38085,N_39501);
or U44159 (N_44159,N_39790,N_37759);
or U44160 (N_44160,N_38515,N_35217);
and U44161 (N_44161,N_36997,N_37508);
nand U44162 (N_44162,N_36657,N_36023);
nor U44163 (N_44163,N_36580,N_37181);
nor U44164 (N_44164,N_37716,N_36434);
xor U44165 (N_44165,N_37428,N_37308);
nor U44166 (N_44166,N_35956,N_38102);
or U44167 (N_44167,N_36806,N_39398);
and U44168 (N_44168,N_38177,N_39877);
or U44169 (N_44169,N_37084,N_35743);
nand U44170 (N_44170,N_39792,N_38765);
nand U44171 (N_44171,N_37281,N_38866);
nand U44172 (N_44172,N_38669,N_35179);
xor U44173 (N_44173,N_38330,N_36954);
or U44174 (N_44174,N_36225,N_39368);
or U44175 (N_44175,N_38761,N_36648);
or U44176 (N_44176,N_36673,N_35918);
and U44177 (N_44177,N_35872,N_35338);
nor U44178 (N_44178,N_39490,N_37446);
and U44179 (N_44179,N_39279,N_36888);
or U44180 (N_44180,N_37885,N_36991);
nand U44181 (N_44181,N_37352,N_38866);
xnor U44182 (N_44182,N_38690,N_35669);
nor U44183 (N_44183,N_38102,N_39491);
nand U44184 (N_44184,N_39490,N_37488);
nand U44185 (N_44185,N_39596,N_38980);
and U44186 (N_44186,N_35150,N_39102);
and U44187 (N_44187,N_39871,N_36461);
or U44188 (N_44188,N_38204,N_36639);
nor U44189 (N_44189,N_38908,N_39272);
nor U44190 (N_44190,N_39331,N_35534);
nor U44191 (N_44191,N_35388,N_36251);
or U44192 (N_44192,N_38444,N_36339);
and U44193 (N_44193,N_38255,N_39521);
nand U44194 (N_44194,N_36662,N_39451);
and U44195 (N_44195,N_36173,N_38158);
nor U44196 (N_44196,N_39054,N_38963);
and U44197 (N_44197,N_35554,N_38209);
and U44198 (N_44198,N_38867,N_35404);
xnor U44199 (N_44199,N_39197,N_35105);
nand U44200 (N_44200,N_38669,N_35401);
or U44201 (N_44201,N_39097,N_39705);
and U44202 (N_44202,N_35016,N_36792);
nor U44203 (N_44203,N_35704,N_39802);
or U44204 (N_44204,N_35837,N_38766);
xor U44205 (N_44205,N_35024,N_35491);
or U44206 (N_44206,N_37135,N_36302);
xnor U44207 (N_44207,N_36734,N_35231);
and U44208 (N_44208,N_36058,N_39524);
or U44209 (N_44209,N_36595,N_36989);
nand U44210 (N_44210,N_38244,N_35685);
or U44211 (N_44211,N_39470,N_39854);
nand U44212 (N_44212,N_37024,N_37371);
xnor U44213 (N_44213,N_35496,N_38233);
or U44214 (N_44214,N_36845,N_35871);
nor U44215 (N_44215,N_39542,N_36436);
nand U44216 (N_44216,N_35706,N_36539);
or U44217 (N_44217,N_37173,N_37507);
and U44218 (N_44218,N_37900,N_37172);
or U44219 (N_44219,N_36803,N_39860);
xnor U44220 (N_44220,N_35471,N_36884);
nor U44221 (N_44221,N_35830,N_36849);
xnor U44222 (N_44222,N_39461,N_35919);
or U44223 (N_44223,N_39419,N_35931);
xor U44224 (N_44224,N_38322,N_38041);
or U44225 (N_44225,N_35605,N_38558);
xor U44226 (N_44226,N_37236,N_35401);
and U44227 (N_44227,N_38428,N_35161);
xor U44228 (N_44228,N_39132,N_35739);
and U44229 (N_44229,N_36003,N_37460);
and U44230 (N_44230,N_37560,N_36480);
nand U44231 (N_44231,N_36251,N_38445);
or U44232 (N_44232,N_36013,N_38145);
nor U44233 (N_44233,N_39232,N_36552);
or U44234 (N_44234,N_38526,N_37868);
nor U44235 (N_44235,N_36919,N_35516);
xnor U44236 (N_44236,N_35682,N_37342);
nand U44237 (N_44237,N_35154,N_38444);
xor U44238 (N_44238,N_39979,N_37294);
nand U44239 (N_44239,N_35560,N_35444);
and U44240 (N_44240,N_38391,N_36650);
and U44241 (N_44241,N_36578,N_38668);
and U44242 (N_44242,N_38794,N_37602);
nor U44243 (N_44243,N_37302,N_37987);
xnor U44244 (N_44244,N_39010,N_37271);
nor U44245 (N_44245,N_36376,N_39138);
xnor U44246 (N_44246,N_36677,N_39853);
or U44247 (N_44247,N_38149,N_39287);
nor U44248 (N_44248,N_39851,N_38235);
xnor U44249 (N_44249,N_37018,N_35408);
nor U44250 (N_44250,N_36941,N_38196);
and U44251 (N_44251,N_36472,N_35633);
xnor U44252 (N_44252,N_37913,N_37055);
or U44253 (N_44253,N_36998,N_38695);
nor U44254 (N_44254,N_39395,N_36515);
or U44255 (N_44255,N_39345,N_35478);
xor U44256 (N_44256,N_37558,N_39308);
nor U44257 (N_44257,N_36886,N_38548);
or U44258 (N_44258,N_38477,N_39388);
xnor U44259 (N_44259,N_36284,N_38947);
and U44260 (N_44260,N_38579,N_36598);
or U44261 (N_44261,N_38858,N_38800);
and U44262 (N_44262,N_36234,N_36958);
xor U44263 (N_44263,N_36020,N_39634);
and U44264 (N_44264,N_35931,N_37327);
xnor U44265 (N_44265,N_39585,N_35277);
or U44266 (N_44266,N_37832,N_37661);
or U44267 (N_44267,N_35124,N_37514);
xor U44268 (N_44268,N_36214,N_38207);
nand U44269 (N_44269,N_39147,N_39397);
nand U44270 (N_44270,N_39365,N_37465);
and U44271 (N_44271,N_39492,N_39567);
or U44272 (N_44272,N_38447,N_36697);
nand U44273 (N_44273,N_36293,N_35378);
or U44274 (N_44274,N_37852,N_35768);
and U44275 (N_44275,N_35512,N_39359);
nor U44276 (N_44276,N_37779,N_37774);
and U44277 (N_44277,N_39873,N_36757);
nand U44278 (N_44278,N_37249,N_37496);
or U44279 (N_44279,N_37804,N_35035);
nand U44280 (N_44280,N_36238,N_35386);
and U44281 (N_44281,N_35545,N_38312);
nand U44282 (N_44282,N_39159,N_37880);
nor U44283 (N_44283,N_35364,N_39761);
or U44284 (N_44284,N_39846,N_37311);
nor U44285 (N_44285,N_36291,N_35776);
xor U44286 (N_44286,N_38407,N_36778);
nor U44287 (N_44287,N_37660,N_35837);
or U44288 (N_44288,N_39097,N_36416);
xor U44289 (N_44289,N_38148,N_38354);
xor U44290 (N_44290,N_35043,N_37095);
or U44291 (N_44291,N_37307,N_37340);
nor U44292 (N_44292,N_35739,N_35873);
and U44293 (N_44293,N_38097,N_35996);
nor U44294 (N_44294,N_38689,N_38841);
nor U44295 (N_44295,N_39074,N_37697);
nor U44296 (N_44296,N_36023,N_35236);
or U44297 (N_44297,N_35580,N_39002);
and U44298 (N_44298,N_37812,N_37366);
nor U44299 (N_44299,N_38332,N_35076);
nand U44300 (N_44300,N_38202,N_39246);
nor U44301 (N_44301,N_36049,N_36390);
nand U44302 (N_44302,N_37583,N_37683);
or U44303 (N_44303,N_37159,N_39066);
xor U44304 (N_44304,N_36604,N_36333);
or U44305 (N_44305,N_36112,N_39308);
and U44306 (N_44306,N_37866,N_39627);
nand U44307 (N_44307,N_38013,N_38167);
and U44308 (N_44308,N_36903,N_37554);
or U44309 (N_44309,N_39630,N_35938);
nand U44310 (N_44310,N_39035,N_38068);
xnor U44311 (N_44311,N_39645,N_36900);
or U44312 (N_44312,N_39756,N_36281);
nor U44313 (N_44313,N_39473,N_35247);
xor U44314 (N_44314,N_36762,N_37380);
and U44315 (N_44315,N_39775,N_37861);
nand U44316 (N_44316,N_36963,N_36436);
and U44317 (N_44317,N_36044,N_38703);
nor U44318 (N_44318,N_37279,N_39251);
or U44319 (N_44319,N_38869,N_35989);
nor U44320 (N_44320,N_36632,N_36881);
nand U44321 (N_44321,N_37692,N_36199);
nand U44322 (N_44322,N_38805,N_35104);
nor U44323 (N_44323,N_36933,N_38374);
and U44324 (N_44324,N_39913,N_39804);
nor U44325 (N_44325,N_36912,N_35660);
and U44326 (N_44326,N_35389,N_38990);
nor U44327 (N_44327,N_36659,N_39779);
nor U44328 (N_44328,N_36996,N_35770);
and U44329 (N_44329,N_37526,N_36758);
and U44330 (N_44330,N_39335,N_35847);
or U44331 (N_44331,N_35673,N_37123);
nor U44332 (N_44332,N_35341,N_39021);
nor U44333 (N_44333,N_36920,N_37269);
nor U44334 (N_44334,N_36164,N_37172);
and U44335 (N_44335,N_39841,N_37152);
xnor U44336 (N_44336,N_37419,N_39358);
xnor U44337 (N_44337,N_39269,N_39195);
xnor U44338 (N_44338,N_37069,N_37601);
xnor U44339 (N_44339,N_37732,N_37677);
and U44340 (N_44340,N_37271,N_39000);
or U44341 (N_44341,N_38216,N_36015);
nand U44342 (N_44342,N_35926,N_35055);
nor U44343 (N_44343,N_39249,N_36431);
nor U44344 (N_44344,N_39033,N_35197);
nor U44345 (N_44345,N_36828,N_35731);
nand U44346 (N_44346,N_38529,N_39053);
nand U44347 (N_44347,N_39695,N_35597);
nor U44348 (N_44348,N_39989,N_39157);
and U44349 (N_44349,N_39889,N_37509);
xnor U44350 (N_44350,N_39922,N_36485);
and U44351 (N_44351,N_35629,N_39513);
xor U44352 (N_44352,N_36356,N_39880);
nor U44353 (N_44353,N_36787,N_36418);
nand U44354 (N_44354,N_38280,N_35335);
xor U44355 (N_44355,N_36749,N_36610);
or U44356 (N_44356,N_38014,N_39871);
and U44357 (N_44357,N_37221,N_35456);
nor U44358 (N_44358,N_39574,N_38461);
or U44359 (N_44359,N_36392,N_35794);
nand U44360 (N_44360,N_39981,N_36023);
or U44361 (N_44361,N_37255,N_39361);
or U44362 (N_44362,N_38037,N_37077);
xor U44363 (N_44363,N_35781,N_36262);
nand U44364 (N_44364,N_36150,N_36832);
and U44365 (N_44365,N_35436,N_35827);
or U44366 (N_44366,N_38211,N_39170);
nor U44367 (N_44367,N_36661,N_39667);
xnor U44368 (N_44368,N_37540,N_35269);
or U44369 (N_44369,N_39135,N_36299);
and U44370 (N_44370,N_36513,N_35426);
nand U44371 (N_44371,N_35835,N_37601);
nor U44372 (N_44372,N_39890,N_38340);
nand U44373 (N_44373,N_39632,N_39091);
and U44374 (N_44374,N_35454,N_37920);
and U44375 (N_44375,N_37700,N_36479);
nand U44376 (N_44376,N_38473,N_39526);
nand U44377 (N_44377,N_37434,N_39064);
xnor U44378 (N_44378,N_35162,N_39412);
and U44379 (N_44379,N_38400,N_35023);
and U44380 (N_44380,N_35755,N_39200);
xor U44381 (N_44381,N_38936,N_39500);
or U44382 (N_44382,N_38957,N_37862);
nor U44383 (N_44383,N_38827,N_35664);
or U44384 (N_44384,N_38660,N_35548);
or U44385 (N_44385,N_36176,N_37140);
nor U44386 (N_44386,N_36293,N_39883);
nand U44387 (N_44387,N_35997,N_36206);
nor U44388 (N_44388,N_37487,N_39631);
xor U44389 (N_44389,N_38956,N_36882);
or U44390 (N_44390,N_35398,N_37837);
nor U44391 (N_44391,N_36864,N_38271);
and U44392 (N_44392,N_36742,N_36876);
and U44393 (N_44393,N_35258,N_35277);
and U44394 (N_44394,N_36645,N_38995);
or U44395 (N_44395,N_39277,N_39226);
or U44396 (N_44396,N_36112,N_36762);
or U44397 (N_44397,N_36281,N_37341);
or U44398 (N_44398,N_35755,N_38336);
or U44399 (N_44399,N_39333,N_36015);
or U44400 (N_44400,N_37194,N_35917);
or U44401 (N_44401,N_36554,N_38891);
and U44402 (N_44402,N_35821,N_37894);
or U44403 (N_44403,N_35243,N_35228);
xor U44404 (N_44404,N_35881,N_36115);
nor U44405 (N_44405,N_39068,N_39240);
nor U44406 (N_44406,N_35445,N_36228);
nand U44407 (N_44407,N_37293,N_39366);
xor U44408 (N_44408,N_39055,N_35211);
nor U44409 (N_44409,N_39789,N_36201);
or U44410 (N_44410,N_38208,N_36378);
or U44411 (N_44411,N_36333,N_36279);
or U44412 (N_44412,N_35066,N_39475);
nor U44413 (N_44413,N_37377,N_39694);
or U44414 (N_44414,N_35082,N_37359);
nand U44415 (N_44415,N_37583,N_36405);
or U44416 (N_44416,N_35861,N_36970);
nand U44417 (N_44417,N_37656,N_36276);
and U44418 (N_44418,N_37829,N_37320);
or U44419 (N_44419,N_35680,N_37050);
nand U44420 (N_44420,N_38479,N_37656);
nand U44421 (N_44421,N_36847,N_39031);
and U44422 (N_44422,N_39831,N_35362);
nand U44423 (N_44423,N_37226,N_38458);
nor U44424 (N_44424,N_35288,N_36005);
xor U44425 (N_44425,N_39925,N_39423);
nand U44426 (N_44426,N_39017,N_35560);
xnor U44427 (N_44427,N_39606,N_36117);
nand U44428 (N_44428,N_38477,N_37081);
or U44429 (N_44429,N_38645,N_39433);
and U44430 (N_44430,N_37399,N_36652);
and U44431 (N_44431,N_36671,N_35306);
or U44432 (N_44432,N_36919,N_36888);
or U44433 (N_44433,N_36187,N_39573);
xor U44434 (N_44434,N_35557,N_39998);
or U44435 (N_44435,N_36652,N_39340);
nand U44436 (N_44436,N_39919,N_37130);
or U44437 (N_44437,N_36742,N_35004);
nor U44438 (N_44438,N_35409,N_37267);
nor U44439 (N_44439,N_36877,N_36368);
xor U44440 (N_44440,N_38466,N_37302);
xnor U44441 (N_44441,N_37972,N_38517);
and U44442 (N_44442,N_39000,N_35285);
or U44443 (N_44443,N_38159,N_37588);
nor U44444 (N_44444,N_38133,N_38001);
and U44445 (N_44445,N_36017,N_39457);
or U44446 (N_44446,N_39531,N_35019);
nand U44447 (N_44447,N_36183,N_39903);
nand U44448 (N_44448,N_39250,N_38512);
nand U44449 (N_44449,N_37530,N_35583);
xor U44450 (N_44450,N_37064,N_37086);
and U44451 (N_44451,N_37597,N_36043);
and U44452 (N_44452,N_37835,N_36860);
or U44453 (N_44453,N_37028,N_36866);
nor U44454 (N_44454,N_36442,N_38812);
or U44455 (N_44455,N_35603,N_38571);
or U44456 (N_44456,N_39619,N_39916);
nand U44457 (N_44457,N_36045,N_38366);
nor U44458 (N_44458,N_37047,N_36485);
nor U44459 (N_44459,N_35965,N_39533);
and U44460 (N_44460,N_35498,N_37322);
or U44461 (N_44461,N_36901,N_37399);
nor U44462 (N_44462,N_35554,N_39919);
xnor U44463 (N_44463,N_38165,N_39783);
nand U44464 (N_44464,N_36749,N_38695);
nor U44465 (N_44465,N_36457,N_39569);
xnor U44466 (N_44466,N_35925,N_36863);
nand U44467 (N_44467,N_37334,N_38269);
xor U44468 (N_44468,N_37524,N_38343);
nand U44469 (N_44469,N_37656,N_37517);
and U44470 (N_44470,N_39892,N_38786);
nor U44471 (N_44471,N_37014,N_37038);
or U44472 (N_44472,N_38680,N_35079);
and U44473 (N_44473,N_37690,N_37129);
nand U44474 (N_44474,N_36269,N_38963);
xor U44475 (N_44475,N_38574,N_36908);
or U44476 (N_44476,N_36339,N_38100);
nor U44477 (N_44477,N_35596,N_38520);
nor U44478 (N_44478,N_36379,N_37138);
nand U44479 (N_44479,N_35673,N_37074);
xor U44480 (N_44480,N_39195,N_38131);
nand U44481 (N_44481,N_37351,N_37500);
nand U44482 (N_44482,N_39670,N_37925);
or U44483 (N_44483,N_37212,N_39862);
and U44484 (N_44484,N_39798,N_39929);
or U44485 (N_44485,N_37732,N_36437);
nand U44486 (N_44486,N_36682,N_39537);
and U44487 (N_44487,N_36643,N_39601);
nand U44488 (N_44488,N_37503,N_35506);
nand U44489 (N_44489,N_35482,N_35199);
and U44490 (N_44490,N_36783,N_38631);
nand U44491 (N_44491,N_37019,N_35732);
nand U44492 (N_44492,N_38929,N_38461);
nand U44493 (N_44493,N_39118,N_36727);
xnor U44494 (N_44494,N_35599,N_39709);
or U44495 (N_44495,N_35419,N_39661);
nor U44496 (N_44496,N_39638,N_39572);
xor U44497 (N_44497,N_39676,N_35249);
or U44498 (N_44498,N_38759,N_35434);
and U44499 (N_44499,N_36626,N_39485);
and U44500 (N_44500,N_39523,N_35835);
nor U44501 (N_44501,N_36738,N_35664);
xor U44502 (N_44502,N_38082,N_37314);
nand U44503 (N_44503,N_37470,N_38052);
and U44504 (N_44504,N_35536,N_35637);
nand U44505 (N_44505,N_38136,N_37496);
and U44506 (N_44506,N_35069,N_39641);
nor U44507 (N_44507,N_38310,N_35768);
nand U44508 (N_44508,N_36739,N_39389);
nand U44509 (N_44509,N_35076,N_39214);
and U44510 (N_44510,N_38065,N_37800);
xor U44511 (N_44511,N_38813,N_36231);
xor U44512 (N_44512,N_36430,N_38185);
or U44513 (N_44513,N_36280,N_38166);
xor U44514 (N_44514,N_38624,N_35060);
or U44515 (N_44515,N_36866,N_35422);
nand U44516 (N_44516,N_39186,N_36815);
xnor U44517 (N_44517,N_35457,N_38429);
xor U44518 (N_44518,N_37881,N_35794);
nand U44519 (N_44519,N_36160,N_39112);
nand U44520 (N_44520,N_38046,N_36069);
nor U44521 (N_44521,N_37048,N_36072);
and U44522 (N_44522,N_39561,N_37269);
xor U44523 (N_44523,N_37718,N_36646);
or U44524 (N_44524,N_39210,N_37819);
nor U44525 (N_44525,N_39518,N_36791);
and U44526 (N_44526,N_37956,N_37343);
nor U44527 (N_44527,N_39317,N_35475);
or U44528 (N_44528,N_36138,N_38071);
nand U44529 (N_44529,N_37204,N_35938);
and U44530 (N_44530,N_35770,N_37284);
and U44531 (N_44531,N_36470,N_38020);
nor U44532 (N_44532,N_37633,N_36830);
xor U44533 (N_44533,N_37426,N_36523);
and U44534 (N_44534,N_35049,N_35266);
and U44535 (N_44535,N_39589,N_39018);
or U44536 (N_44536,N_36498,N_39488);
and U44537 (N_44537,N_36248,N_39965);
nor U44538 (N_44538,N_35135,N_36895);
nand U44539 (N_44539,N_37696,N_37052);
nand U44540 (N_44540,N_35588,N_39753);
or U44541 (N_44541,N_37666,N_37231);
nor U44542 (N_44542,N_36788,N_38735);
or U44543 (N_44543,N_39845,N_38569);
or U44544 (N_44544,N_35280,N_37056);
nand U44545 (N_44545,N_38347,N_38928);
xor U44546 (N_44546,N_36312,N_35160);
nand U44547 (N_44547,N_35932,N_38665);
nand U44548 (N_44548,N_37760,N_37490);
nand U44549 (N_44549,N_39356,N_36552);
xor U44550 (N_44550,N_36181,N_35616);
or U44551 (N_44551,N_36967,N_39785);
or U44552 (N_44552,N_37267,N_38157);
and U44553 (N_44553,N_38109,N_35098);
and U44554 (N_44554,N_39209,N_37769);
or U44555 (N_44555,N_39706,N_37199);
and U44556 (N_44556,N_37941,N_38830);
or U44557 (N_44557,N_38436,N_37012);
and U44558 (N_44558,N_36297,N_36727);
and U44559 (N_44559,N_35283,N_35329);
nand U44560 (N_44560,N_35270,N_38485);
or U44561 (N_44561,N_35087,N_36363);
or U44562 (N_44562,N_35776,N_39689);
nor U44563 (N_44563,N_39261,N_36119);
xnor U44564 (N_44564,N_38079,N_38579);
xor U44565 (N_44565,N_38179,N_35053);
and U44566 (N_44566,N_36785,N_37757);
nand U44567 (N_44567,N_36732,N_36764);
nand U44568 (N_44568,N_37746,N_38242);
nand U44569 (N_44569,N_35328,N_39320);
nor U44570 (N_44570,N_39763,N_36193);
xnor U44571 (N_44571,N_36060,N_37064);
nor U44572 (N_44572,N_39140,N_36668);
and U44573 (N_44573,N_35014,N_35693);
or U44574 (N_44574,N_39747,N_38015);
xor U44575 (N_44575,N_36787,N_37351);
xnor U44576 (N_44576,N_36833,N_36055);
xnor U44577 (N_44577,N_37758,N_37295);
nor U44578 (N_44578,N_37086,N_38487);
xor U44579 (N_44579,N_38821,N_37042);
xor U44580 (N_44580,N_39570,N_39385);
nand U44581 (N_44581,N_35754,N_37275);
and U44582 (N_44582,N_36473,N_38380);
nand U44583 (N_44583,N_38754,N_36369);
nand U44584 (N_44584,N_37641,N_38810);
nor U44585 (N_44585,N_35919,N_37203);
nor U44586 (N_44586,N_36239,N_35781);
xor U44587 (N_44587,N_36086,N_39304);
xor U44588 (N_44588,N_36020,N_38095);
nor U44589 (N_44589,N_37623,N_38293);
nand U44590 (N_44590,N_35636,N_36654);
nor U44591 (N_44591,N_39072,N_39682);
xnor U44592 (N_44592,N_39868,N_36325);
or U44593 (N_44593,N_36354,N_38952);
and U44594 (N_44594,N_38316,N_39314);
or U44595 (N_44595,N_38724,N_36571);
xor U44596 (N_44596,N_39934,N_35422);
nand U44597 (N_44597,N_39438,N_35053);
nor U44598 (N_44598,N_38123,N_39983);
nand U44599 (N_44599,N_36042,N_37028);
xnor U44600 (N_44600,N_35779,N_36792);
or U44601 (N_44601,N_36811,N_35092);
xor U44602 (N_44602,N_38282,N_37255);
nand U44603 (N_44603,N_38588,N_35190);
and U44604 (N_44604,N_39023,N_36215);
xnor U44605 (N_44605,N_36177,N_37822);
or U44606 (N_44606,N_37034,N_37471);
xnor U44607 (N_44607,N_38670,N_35836);
and U44608 (N_44608,N_37221,N_39113);
nor U44609 (N_44609,N_36083,N_37093);
nor U44610 (N_44610,N_35059,N_35949);
nor U44611 (N_44611,N_39206,N_36970);
nand U44612 (N_44612,N_37723,N_37957);
xnor U44613 (N_44613,N_38290,N_37203);
nor U44614 (N_44614,N_36093,N_37923);
nor U44615 (N_44615,N_39921,N_37505);
xor U44616 (N_44616,N_39240,N_35478);
and U44617 (N_44617,N_37764,N_39119);
and U44618 (N_44618,N_39722,N_36208);
or U44619 (N_44619,N_35881,N_35479);
nand U44620 (N_44620,N_39147,N_35830);
nand U44621 (N_44621,N_36272,N_35172);
nand U44622 (N_44622,N_35352,N_35208);
or U44623 (N_44623,N_38325,N_37223);
xor U44624 (N_44624,N_37476,N_36891);
nor U44625 (N_44625,N_35217,N_36207);
nor U44626 (N_44626,N_37556,N_35678);
xor U44627 (N_44627,N_38438,N_37846);
xor U44628 (N_44628,N_39737,N_36229);
xnor U44629 (N_44629,N_39850,N_37224);
nor U44630 (N_44630,N_36485,N_36924);
and U44631 (N_44631,N_35928,N_35622);
or U44632 (N_44632,N_38692,N_39202);
nor U44633 (N_44633,N_36875,N_39225);
nor U44634 (N_44634,N_36217,N_36512);
nor U44635 (N_44635,N_39495,N_36808);
nor U44636 (N_44636,N_35485,N_39814);
xor U44637 (N_44637,N_37332,N_39831);
and U44638 (N_44638,N_35900,N_36689);
or U44639 (N_44639,N_39791,N_39749);
nand U44640 (N_44640,N_39237,N_38351);
nand U44641 (N_44641,N_37587,N_36891);
nand U44642 (N_44642,N_39255,N_38894);
nor U44643 (N_44643,N_37658,N_37013);
nand U44644 (N_44644,N_35736,N_37212);
and U44645 (N_44645,N_36232,N_39683);
xnor U44646 (N_44646,N_39910,N_35990);
nor U44647 (N_44647,N_37489,N_39280);
nand U44648 (N_44648,N_35123,N_35587);
nor U44649 (N_44649,N_37416,N_39905);
nand U44650 (N_44650,N_35937,N_39354);
nand U44651 (N_44651,N_35349,N_36660);
nor U44652 (N_44652,N_37029,N_35763);
and U44653 (N_44653,N_39267,N_38154);
nor U44654 (N_44654,N_39091,N_38769);
and U44655 (N_44655,N_35235,N_35757);
or U44656 (N_44656,N_38980,N_37650);
and U44657 (N_44657,N_38983,N_36327);
or U44658 (N_44658,N_36955,N_36102);
nor U44659 (N_44659,N_38298,N_36365);
nor U44660 (N_44660,N_35003,N_36292);
nor U44661 (N_44661,N_39646,N_38086);
xor U44662 (N_44662,N_35941,N_39148);
nand U44663 (N_44663,N_36863,N_39777);
xnor U44664 (N_44664,N_39880,N_37523);
xnor U44665 (N_44665,N_36230,N_35366);
nand U44666 (N_44666,N_39980,N_35202);
nor U44667 (N_44667,N_35574,N_35381);
xnor U44668 (N_44668,N_38164,N_39300);
and U44669 (N_44669,N_36823,N_38734);
nand U44670 (N_44670,N_36224,N_36712);
nor U44671 (N_44671,N_35515,N_38419);
nor U44672 (N_44672,N_38304,N_36506);
nand U44673 (N_44673,N_36980,N_38366);
and U44674 (N_44674,N_36013,N_39493);
or U44675 (N_44675,N_38564,N_38837);
xnor U44676 (N_44676,N_36564,N_38985);
or U44677 (N_44677,N_37793,N_36694);
nor U44678 (N_44678,N_38885,N_37777);
nor U44679 (N_44679,N_38290,N_38585);
nor U44680 (N_44680,N_37708,N_36929);
nor U44681 (N_44681,N_35837,N_35111);
or U44682 (N_44682,N_39160,N_38207);
and U44683 (N_44683,N_35202,N_38555);
and U44684 (N_44684,N_37321,N_39309);
xor U44685 (N_44685,N_39440,N_39801);
nand U44686 (N_44686,N_39332,N_37234);
and U44687 (N_44687,N_35423,N_35892);
and U44688 (N_44688,N_38138,N_36050);
nand U44689 (N_44689,N_35299,N_38717);
and U44690 (N_44690,N_35104,N_39794);
or U44691 (N_44691,N_36805,N_38962);
nand U44692 (N_44692,N_37239,N_38929);
nand U44693 (N_44693,N_35982,N_36878);
or U44694 (N_44694,N_38360,N_37643);
nor U44695 (N_44695,N_36435,N_37119);
and U44696 (N_44696,N_38152,N_38944);
nand U44697 (N_44697,N_36238,N_35789);
or U44698 (N_44698,N_36837,N_37187);
xor U44699 (N_44699,N_37950,N_35169);
nor U44700 (N_44700,N_39165,N_37427);
nand U44701 (N_44701,N_38944,N_35780);
xor U44702 (N_44702,N_38688,N_35096);
or U44703 (N_44703,N_38148,N_39033);
xnor U44704 (N_44704,N_37300,N_39286);
or U44705 (N_44705,N_39554,N_37243);
nor U44706 (N_44706,N_37771,N_35407);
xor U44707 (N_44707,N_38439,N_39358);
and U44708 (N_44708,N_38653,N_39189);
or U44709 (N_44709,N_37287,N_38957);
and U44710 (N_44710,N_39304,N_35191);
nand U44711 (N_44711,N_35205,N_38398);
and U44712 (N_44712,N_38342,N_37606);
nor U44713 (N_44713,N_37714,N_36024);
nand U44714 (N_44714,N_38652,N_38730);
or U44715 (N_44715,N_35888,N_39067);
xor U44716 (N_44716,N_35376,N_36165);
and U44717 (N_44717,N_39696,N_38570);
and U44718 (N_44718,N_38047,N_38195);
nand U44719 (N_44719,N_39255,N_38820);
xor U44720 (N_44720,N_36398,N_38658);
and U44721 (N_44721,N_35110,N_36815);
nand U44722 (N_44722,N_35777,N_38551);
xnor U44723 (N_44723,N_35264,N_36595);
or U44724 (N_44724,N_39049,N_35825);
nor U44725 (N_44725,N_38400,N_35929);
xor U44726 (N_44726,N_39213,N_37362);
or U44727 (N_44727,N_38960,N_36432);
xor U44728 (N_44728,N_35901,N_37264);
and U44729 (N_44729,N_38864,N_38476);
nor U44730 (N_44730,N_37738,N_37187);
and U44731 (N_44731,N_39498,N_39945);
xor U44732 (N_44732,N_39588,N_35699);
nand U44733 (N_44733,N_35857,N_35676);
nand U44734 (N_44734,N_38998,N_35063);
nand U44735 (N_44735,N_35171,N_35576);
and U44736 (N_44736,N_36321,N_35408);
xor U44737 (N_44737,N_37704,N_35129);
nand U44738 (N_44738,N_36778,N_37985);
xnor U44739 (N_44739,N_35702,N_37356);
or U44740 (N_44740,N_39999,N_37269);
nand U44741 (N_44741,N_35139,N_39849);
nor U44742 (N_44742,N_37682,N_36682);
xor U44743 (N_44743,N_37086,N_38864);
and U44744 (N_44744,N_37204,N_37176);
nor U44745 (N_44745,N_37940,N_35340);
nand U44746 (N_44746,N_39815,N_38838);
or U44747 (N_44747,N_35105,N_35388);
and U44748 (N_44748,N_36920,N_39410);
nand U44749 (N_44749,N_37802,N_39688);
xor U44750 (N_44750,N_36881,N_39621);
nor U44751 (N_44751,N_39297,N_39181);
nand U44752 (N_44752,N_36702,N_38248);
nor U44753 (N_44753,N_37082,N_37982);
xnor U44754 (N_44754,N_39193,N_38326);
or U44755 (N_44755,N_35109,N_37208);
nand U44756 (N_44756,N_38582,N_38973);
xor U44757 (N_44757,N_37210,N_38572);
nor U44758 (N_44758,N_37042,N_37362);
nand U44759 (N_44759,N_38604,N_38241);
nand U44760 (N_44760,N_35223,N_39406);
nor U44761 (N_44761,N_37774,N_39463);
or U44762 (N_44762,N_38194,N_38508);
nand U44763 (N_44763,N_39030,N_37893);
nor U44764 (N_44764,N_36315,N_39132);
nand U44765 (N_44765,N_37827,N_36092);
and U44766 (N_44766,N_37518,N_38199);
nor U44767 (N_44767,N_36635,N_37944);
xor U44768 (N_44768,N_38671,N_39067);
nand U44769 (N_44769,N_36886,N_39720);
xnor U44770 (N_44770,N_39570,N_36918);
xor U44771 (N_44771,N_39829,N_35407);
and U44772 (N_44772,N_39582,N_38609);
or U44773 (N_44773,N_37356,N_39760);
or U44774 (N_44774,N_37330,N_39763);
and U44775 (N_44775,N_37404,N_36672);
or U44776 (N_44776,N_37664,N_37233);
xnor U44777 (N_44777,N_39200,N_39005);
or U44778 (N_44778,N_35860,N_39164);
nand U44779 (N_44779,N_36940,N_35114);
and U44780 (N_44780,N_36543,N_37039);
nor U44781 (N_44781,N_35722,N_35987);
and U44782 (N_44782,N_39187,N_36198);
and U44783 (N_44783,N_36839,N_37087);
nor U44784 (N_44784,N_36195,N_35869);
and U44785 (N_44785,N_36274,N_38449);
and U44786 (N_44786,N_38051,N_39531);
or U44787 (N_44787,N_38139,N_35622);
nand U44788 (N_44788,N_36379,N_37984);
and U44789 (N_44789,N_39761,N_36557);
nand U44790 (N_44790,N_37943,N_37957);
nand U44791 (N_44791,N_39573,N_36549);
nor U44792 (N_44792,N_35109,N_35908);
xnor U44793 (N_44793,N_35850,N_38653);
xnor U44794 (N_44794,N_39245,N_37894);
or U44795 (N_44795,N_35737,N_38485);
nor U44796 (N_44796,N_38395,N_35817);
nand U44797 (N_44797,N_35841,N_36967);
nand U44798 (N_44798,N_35418,N_39162);
xor U44799 (N_44799,N_37224,N_38637);
or U44800 (N_44800,N_36977,N_36768);
xnor U44801 (N_44801,N_38714,N_38931);
or U44802 (N_44802,N_38555,N_38216);
or U44803 (N_44803,N_38161,N_39760);
and U44804 (N_44804,N_38420,N_38482);
nor U44805 (N_44805,N_35200,N_37500);
nand U44806 (N_44806,N_35620,N_35633);
nand U44807 (N_44807,N_37506,N_36782);
nor U44808 (N_44808,N_38293,N_38007);
xnor U44809 (N_44809,N_37897,N_35379);
xor U44810 (N_44810,N_38598,N_38441);
nand U44811 (N_44811,N_37045,N_35954);
xnor U44812 (N_44812,N_36901,N_37847);
nor U44813 (N_44813,N_35475,N_38383);
xnor U44814 (N_44814,N_36508,N_39927);
and U44815 (N_44815,N_37798,N_39504);
and U44816 (N_44816,N_39042,N_35228);
xnor U44817 (N_44817,N_37605,N_37126);
nor U44818 (N_44818,N_35365,N_36936);
or U44819 (N_44819,N_38535,N_36701);
xor U44820 (N_44820,N_36252,N_38900);
xor U44821 (N_44821,N_36155,N_36357);
or U44822 (N_44822,N_36713,N_35368);
nand U44823 (N_44823,N_35035,N_39797);
and U44824 (N_44824,N_36862,N_36519);
xor U44825 (N_44825,N_36856,N_39288);
or U44826 (N_44826,N_39248,N_37511);
and U44827 (N_44827,N_37580,N_36645);
nand U44828 (N_44828,N_35508,N_36745);
or U44829 (N_44829,N_36223,N_36919);
or U44830 (N_44830,N_38752,N_36648);
nand U44831 (N_44831,N_38928,N_37065);
or U44832 (N_44832,N_36037,N_36644);
xnor U44833 (N_44833,N_37575,N_39100);
xor U44834 (N_44834,N_35709,N_35790);
and U44835 (N_44835,N_39598,N_39895);
and U44836 (N_44836,N_36846,N_39712);
nand U44837 (N_44837,N_35545,N_38680);
or U44838 (N_44838,N_39897,N_38529);
xnor U44839 (N_44839,N_36687,N_37616);
and U44840 (N_44840,N_37282,N_36120);
and U44841 (N_44841,N_36317,N_35834);
nand U44842 (N_44842,N_39295,N_38952);
and U44843 (N_44843,N_37009,N_39877);
nand U44844 (N_44844,N_37804,N_35287);
and U44845 (N_44845,N_39224,N_36652);
xor U44846 (N_44846,N_36371,N_36556);
and U44847 (N_44847,N_39090,N_37214);
or U44848 (N_44848,N_39965,N_38053);
or U44849 (N_44849,N_36701,N_36798);
and U44850 (N_44850,N_39363,N_36373);
xnor U44851 (N_44851,N_36687,N_38338);
or U44852 (N_44852,N_38856,N_38132);
and U44853 (N_44853,N_39771,N_37148);
or U44854 (N_44854,N_36360,N_37950);
xor U44855 (N_44855,N_39971,N_37915);
xor U44856 (N_44856,N_36525,N_37173);
xnor U44857 (N_44857,N_35827,N_37233);
nor U44858 (N_44858,N_36289,N_39672);
and U44859 (N_44859,N_36832,N_37926);
or U44860 (N_44860,N_39096,N_37277);
nor U44861 (N_44861,N_35223,N_37505);
and U44862 (N_44862,N_36310,N_39731);
nand U44863 (N_44863,N_36389,N_39690);
nor U44864 (N_44864,N_37317,N_39549);
and U44865 (N_44865,N_37186,N_39638);
nor U44866 (N_44866,N_38362,N_35725);
nor U44867 (N_44867,N_36736,N_39494);
and U44868 (N_44868,N_38818,N_35168);
nand U44869 (N_44869,N_35345,N_39809);
or U44870 (N_44870,N_37406,N_39519);
nand U44871 (N_44871,N_36262,N_36878);
nor U44872 (N_44872,N_36813,N_37606);
and U44873 (N_44873,N_39592,N_39093);
nand U44874 (N_44874,N_37283,N_35988);
or U44875 (N_44875,N_36056,N_39607);
nor U44876 (N_44876,N_37046,N_37798);
or U44877 (N_44877,N_35097,N_39506);
or U44878 (N_44878,N_39927,N_36045);
nor U44879 (N_44879,N_35693,N_37562);
xor U44880 (N_44880,N_36427,N_38593);
xor U44881 (N_44881,N_37359,N_38776);
or U44882 (N_44882,N_35124,N_37837);
and U44883 (N_44883,N_35537,N_35463);
nor U44884 (N_44884,N_35583,N_38722);
xor U44885 (N_44885,N_39306,N_37978);
xor U44886 (N_44886,N_37179,N_36640);
nor U44887 (N_44887,N_37661,N_39944);
and U44888 (N_44888,N_37185,N_36151);
and U44889 (N_44889,N_35422,N_37339);
nand U44890 (N_44890,N_39984,N_38592);
or U44891 (N_44891,N_38946,N_36397);
xor U44892 (N_44892,N_35848,N_36767);
or U44893 (N_44893,N_35507,N_37528);
or U44894 (N_44894,N_39467,N_39369);
or U44895 (N_44895,N_35742,N_36660);
nand U44896 (N_44896,N_36730,N_37726);
nor U44897 (N_44897,N_38975,N_35538);
nor U44898 (N_44898,N_36399,N_39736);
and U44899 (N_44899,N_36826,N_35978);
nand U44900 (N_44900,N_37771,N_35913);
nand U44901 (N_44901,N_39494,N_35257);
nand U44902 (N_44902,N_35409,N_37886);
nor U44903 (N_44903,N_35174,N_36855);
xor U44904 (N_44904,N_37280,N_39282);
and U44905 (N_44905,N_35867,N_39977);
and U44906 (N_44906,N_37330,N_39724);
nand U44907 (N_44907,N_35942,N_37673);
and U44908 (N_44908,N_36334,N_37835);
nand U44909 (N_44909,N_37325,N_36618);
xnor U44910 (N_44910,N_39991,N_35608);
and U44911 (N_44911,N_39038,N_38670);
or U44912 (N_44912,N_37176,N_35144);
nand U44913 (N_44913,N_35372,N_36583);
nand U44914 (N_44914,N_35786,N_39556);
xnor U44915 (N_44915,N_39038,N_38060);
nor U44916 (N_44916,N_38765,N_39613);
nand U44917 (N_44917,N_39341,N_38406);
nand U44918 (N_44918,N_38108,N_39906);
nor U44919 (N_44919,N_38594,N_39902);
nand U44920 (N_44920,N_39273,N_35570);
nand U44921 (N_44921,N_35735,N_36910);
and U44922 (N_44922,N_38785,N_36406);
or U44923 (N_44923,N_36455,N_38155);
xnor U44924 (N_44924,N_35547,N_36633);
and U44925 (N_44925,N_39998,N_38550);
xnor U44926 (N_44926,N_39938,N_38965);
nand U44927 (N_44927,N_37780,N_37731);
nand U44928 (N_44928,N_38594,N_35896);
and U44929 (N_44929,N_35710,N_36840);
or U44930 (N_44930,N_35719,N_36256);
and U44931 (N_44931,N_36355,N_39181);
xnor U44932 (N_44932,N_35615,N_35863);
or U44933 (N_44933,N_37844,N_36459);
xor U44934 (N_44934,N_38473,N_37934);
nor U44935 (N_44935,N_38823,N_37256);
nand U44936 (N_44936,N_36295,N_36042);
or U44937 (N_44937,N_38172,N_35413);
or U44938 (N_44938,N_37091,N_35099);
nor U44939 (N_44939,N_38812,N_38154);
nor U44940 (N_44940,N_35575,N_35268);
xnor U44941 (N_44941,N_36973,N_39052);
nor U44942 (N_44942,N_37118,N_36997);
nor U44943 (N_44943,N_39211,N_39587);
xnor U44944 (N_44944,N_36517,N_36782);
or U44945 (N_44945,N_36881,N_37718);
and U44946 (N_44946,N_35456,N_38657);
nor U44947 (N_44947,N_39011,N_39888);
nand U44948 (N_44948,N_37335,N_35080);
or U44949 (N_44949,N_39439,N_35722);
nand U44950 (N_44950,N_39798,N_37153);
nor U44951 (N_44951,N_39887,N_35016);
nand U44952 (N_44952,N_37190,N_37369);
nor U44953 (N_44953,N_36597,N_39007);
and U44954 (N_44954,N_38489,N_39508);
nor U44955 (N_44955,N_38362,N_37806);
nor U44956 (N_44956,N_36797,N_38784);
xnor U44957 (N_44957,N_38601,N_35687);
or U44958 (N_44958,N_38671,N_36678);
nand U44959 (N_44959,N_35980,N_39251);
xor U44960 (N_44960,N_37453,N_38670);
nor U44961 (N_44961,N_35784,N_38051);
xor U44962 (N_44962,N_36829,N_38226);
nand U44963 (N_44963,N_39945,N_37465);
xor U44964 (N_44964,N_36160,N_36207);
xor U44965 (N_44965,N_35071,N_38246);
nor U44966 (N_44966,N_37712,N_37487);
and U44967 (N_44967,N_35611,N_36963);
or U44968 (N_44968,N_35336,N_36308);
nor U44969 (N_44969,N_37174,N_35691);
and U44970 (N_44970,N_38422,N_37561);
or U44971 (N_44971,N_37756,N_37300);
and U44972 (N_44972,N_36087,N_36313);
xor U44973 (N_44973,N_36322,N_36781);
xnor U44974 (N_44974,N_37288,N_35370);
or U44975 (N_44975,N_37803,N_35347);
xnor U44976 (N_44976,N_35746,N_38471);
and U44977 (N_44977,N_38024,N_36731);
and U44978 (N_44978,N_38604,N_37403);
and U44979 (N_44979,N_36916,N_37362);
or U44980 (N_44980,N_38316,N_35210);
nand U44981 (N_44981,N_37252,N_35785);
nand U44982 (N_44982,N_39427,N_38361);
xor U44983 (N_44983,N_36627,N_37075);
nand U44984 (N_44984,N_37571,N_36164);
nor U44985 (N_44985,N_37998,N_35048);
and U44986 (N_44986,N_39684,N_37508);
and U44987 (N_44987,N_37817,N_36184);
and U44988 (N_44988,N_36458,N_35636);
and U44989 (N_44989,N_36113,N_35898);
and U44990 (N_44990,N_39125,N_36479);
and U44991 (N_44991,N_36997,N_35307);
and U44992 (N_44992,N_35641,N_37013);
xnor U44993 (N_44993,N_36930,N_35212);
xnor U44994 (N_44994,N_38062,N_39315);
nand U44995 (N_44995,N_39058,N_37350);
or U44996 (N_44996,N_37649,N_37895);
xnor U44997 (N_44997,N_36766,N_37471);
nand U44998 (N_44998,N_36318,N_38504);
and U44999 (N_44999,N_35321,N_37018);
and U45000 (N_45000,N_40070,N_41095);
xor U45001 (N_45001,N_41139,N_42860);
xnor U45002 (N_45002,N_44073,N_40560);
nor U45003 (N_45003,N_42162,N_41797);
and U45004 (N_45004,N_40399,N_41169);
and U45005 (N_45005,N_40916,N_41524);
xnor U45006 (N_45006,N_44954,N_42509);
nand U45007 (N_45007,N_42103,N_44172);
xnor U45008 (N_45008,N_42858,N_42245);
or U45009 (N_45009,N_40310,N_43910);
and U45010 (N_45010,N_42733,N_44080);
nor U45011 (N_45011,N_40313,N_43589);
nor U45012 (N_45012,N_43332,N_42738);
xnor U45013 (N_45013,N_42898,N_43281);
nor U45014 (N_45014,N_42277,N_44499);
nor U45015 (N_45015,N_44150,N_40872);
xor U45016 (N_45016,N_44759,N_40015);
or U45017 (N_45017,N_44998,N_41000);
or U45018 (N_45018,N_42346,N_43338);
nand U45019 (N_45019,N_43487,N_40573);
and U45020 (N_45020,N_41057,N_40711);
or U45021 (N_45021,N_42338,N_43585);
nor U45022 (N_45022,N_40473,N_44001);
nor U45023 (N_45023,N_43812,N_44734);
nor U45024 (N_45024,N_42035,N_42658);
nand U45025 (N_45025,N_41570,N_41036);
nand U45026 (N_45026,N_40813,N_41677);
or U45027 (N_45027,N_43969,N_40315);
nand U45028 (N_45028,N_44394,N_41703);
xnor U45029 (N_45029,N_41603,N_44859);
and U45030 (N_45030,N_44406,N_41492);
xnor U45031 (N_45031,N_43798,N_41455);
nand U45032 (N_45032,N_42529,N_41035);
xor U45033 (N_45033,N_44855,N_43086);
nor U45034 (N_45034,N_41412,N_44061);
nand U45035 (N_45035,N_42314,N_41737);
and U45036 (N_45036,N_41209,N_41094);
xnor U45037 (N_45037,N_41715,N_40631);
nand U45038 (N_45038,N_40254,N_40505);
nand U45039 (N_45039,N_40027,N_41919);
nand U45040 (N_45040,N_41761,N_44478);
nand U45041 (N_45041,N_44757,N_41587);
nand U45042 (N_45042,N_42391,N_41378);
and U45043 (N_45043,N_42696,N_42850);
and U45044 (N_45044,N_44371,N_44673);
and U45045 (N_45045,N_42533,N_40527);
or U45046 (N_45046,N_40763,N_42697);
and U45047 (N_45047,N_42319,N_44528);
xnor U45048 (N_45048,N_44659,N_41565);
xnor U45049 (N_45049,N_42645,N_42115);
nor U45050 (N_45050,N_42229,N_40046);
or U45051 (N_45051,N_43699,N_41701);
and U45052 (N_45052,N_40892,N_43441);
nor U45053 (N_45053,N_40346,N_42952);
xor U45054 (N_45054,N_42836,N_43764);
nand U45055 (N_45055,N_44186,N_43405);
xor U45056 (N_45056,N_44986,N_44536);
xnor U45057 (N_45057,N_41323,N_40695);
and U45058 (N_45058,N_42655,N_41177);
nor U45059 (N_45059,N_41241,N_44652);
or U45060 (N_45060,N_40798,N_41503);
nand U45061 (N_45061,N_42688,N_44723);
or U45062 (N_45062,N_42454,N_43496);
nand U45063 (N_45063,N_42653,N_41040);
nand U45064 (N_45064,N_42067,N_41397);
and U45065 (N_45065,N_40260,N_44194);
nor U45066 (N_45066,N_41243,N_41066);
nor U45067 (N_45067,N_41778,N_42192);
xor U45068 (N_45068,N_43689,N_44380);
or U45069 (N_45069,N_42197,N_44549);
nor U45070 (N_45070,N_41775,N_41527);
and U45071 (N_45071,N_43390,N_44917);
nor U45072 (N_45072,N_42181,N_41058);
xor U45073 (N_45073,N_41684,N_42424);
and U45074 (N_45074,N_40969,N_44485);
and U45075 (N_45075,N_44355,N_42522);
and U45076 (N_45076,N_40326,N_42867);
xnor U45077 (N_45077,N_41907,N_42154);
xnor U45078 (N_45078,N_40924,N_43903);
xor U45079 (N_45079,N_43518,N_40583);
xnor U45080 (N_45080,N_40441,N_42851);
and U45081 (N_45081,N_40903,N_42014);
xnor U45082 (N_45082,N_43670,N_40443);
xnor U45083 (N_45083,N_41428,N_40189);
xnor U45084 (N_45084,N_44166,N_42341);
nand U45085 (N_45085,N_42300,N_42134);
and U45086 (N_45086,N_42152,N_42825);
or U45087 (N_45087,N_44650,N_42877);
or U45088 (N_45088,N_42007,N_41357);
nor U45089 (N_45089,N_42040,N_43613);
nand U45090 (N_45090,N_41666,N_41215);
and U45091 (N_45091,N_43606,N_40710);
or U45092 (N_45092,N_44192,N_43173);
xor U45093 (N_45093,N_44788,N_41188);
nand U45094 (N_45094,N_40931,N_40165);
nor U45095 (N_45095,N_42973,N_44346);
or U45096 (N_45096,N_42905,N_43758);
nor U45097 (N_45097,N_41765,N_40153);
xor U45098 (N_45098,N_44087,N_44252);
or U45099 (N_45099,N_40411,N_41659);
and U45100 (N_45100,N_42046,N_42216);
nand U45101 (N_45101,N_44382,N_44390);
nand U45102 (N_45102,N_43945,N_41187);
or U45103 (N_45103,N_44690,N_43276);
nand U45104 (N_45104,N_44191,N_41848);
nand U45105 (N_45105,N_41405,N_44991);
and U45106 (N_45106,N_41173,N_42213);
and U45107 (N_45107,N_41005,N_43342);
nand U45108 (N_45108,N_40414,N_43459);
and U45109 (N_45109,N_41767,N_40747);
xor U45110 (N_45110,N_43269,N_43070);
or U45111 (N_45111,N_41998,N_42751);
and U45112 (N_45112,N_41128,N_41225);
nand U45113 (N_45113,N_41687,N_42966);
xor U45114 (N_45114,N_43251,N_42617);
and U45115 (N_45115,N_44432,N_40580);
or U45116 (N_45116,N_44676,N_44487);
nand U45117 (N_45117,N_40345,N_44678);
xnor U45118 (N_45118,N_43561,N_40790);
nand U45119 (N_45119,N_44140,N_40507);
xnor U45120 (N_45120,N_40698,N_42122);
nor U45121 (N_45121,N_40836,N_44318);
nor U45122 (N_45122,N_42743,N_44333);
nand U45123 (N_45123,N_44383,N_41490);
or U45124 (N_45124,N_43452,N_40146);
nand U45125 (N_45125,N_41846,N_43241);
or U45126 (N_45126,N_42353,N_43597);
xnor U45127 (N_45127,N_41594,N_40614);
xor U45128 (N_45128,N_43743,N_43638);
and U45129 (N_45129,N_43448,N_41012);
and U45130 (N_45130,N_43470,N_42578);
xnor U45131 (N_45131,N_44553,N_42818);
and U45132 (N_45132,N_42336,N_43063);
xor U45133 (N_45133,N_42083,N_43372);
or U45134 (N_45134,N_41271,N_40244);
xnor U45135 (N_45135,N_43476,N_42254);
nor U45136 (N_45136,N_40392,N_41063);
xnor U45137 (N_45137,N_41955,N_41985);
and U45138 (N_45138,N_43895,N_43734);
nand U45139 (N_45139,N_44115,N_40524);
or U45140 (N_45140,N_44148,N_44983);
nor U45141 (N_45141,N_41449,N_41023);
nand U45142 (N_45142,N_41895,N_40882);
or U45143 (N_45143,N_41543,N_40003);
nor U45144 (N_45144,N_44065,N_42884);
or U45145 (N_45145,N_42010,N_40318);
nor U45146 (N_45146,N_40004,N_43971);
nor U45147 (N_45147,N_43984,N_42158);
nor U45148 (N_45148,N_41514,N_40201);
nor U45149 (N_45149,N_42703,N_44654);
nor U45150 (N_45150,N_41520,N_43694);
and U45151 (N_45151,N_44544,N_41431);
and U45152 (N_45152,N_41123,N_41402);
and U45153 (N_45153,N_43471,N_41026);
xnor U45154 (N_45154,N_40336,N_44017);
nor U45155 (N_45155,N_43472,N_41902);
xor U45156 (N_45156,N_43396,N_42561);
nand U45157 (N_45157,N_40139,N_43748);
nor U45158 (N_45158,N_44743,N_40736);
nand U45159 (N_45159,N_41471,N_44294);
nand U45160 (N_45160,N_42176,N_44488);
or U45161 (N_45161,N_42273,N_41843);
nand U45162 (N_45162,N_40429,N_41185);
xor U45163 (N_45163,N_44736,N_44058);
and U45164 (N_45164,N_41320,N_41360);
nor U45165 (N_45165,N_44096,N_43465);
nand U45166 (N_45166,N_43235,N_40277);
or U45167 (N_45167,N_44292,N_42599);
or U45168 (N_45168,N_43300,N_43335);
and U45169 (N_45169,N_42762,N_44279);
nor U45170 (N_45170,N_40298,N_41560);
nand U45171 (N_45171,N_41588,N_41769);
nand U45172 (N_45172,N_40486,N_42185);
nand U45173 (N_45173,N_41105,N_40495);
or U45174 (N_45174,N_42530,N_40198);
nand U45175 (N_45175,N_42777,N_41084);
and U45176 (N_45176,N_44989,N_42059);
nand U45177 (N_45177,N_42430,N_44854);
xnor U45178 (N_45178,N_43376,N_41838);
xnor U45179 (N_45179,N_43663,N_42663);
and U45180 (N_45180,N_41523,N_44126);
and U45181 (N_45181,N_41297,N_42641);
and U45182 (N_45182,N_43581,N_40839);
nor U45183 (N_45183,N_44183,N_42908);
nand U45184 (N_45184,N_43307,N_43968);
or U45185 (N_45185,N_42794,N_44624);
and U45186 (N_45186,N_41125,N_41091);
xor U45187 (N_45187,N_43815,N_43103);
nand U45188 (N_45188,N_44814,N_43757);
or U45189 (N_45189,N_40131,N_40817);
nand U45190 (N_45190,N_44152,N_42342);
or U45191 (N_45191,N_40772,N_40841);
nand U45192 (N_45192,N_42586,N_43728);
xnor U45193 (N_45193,N_41699,N_42717);
and U45194 (N_45194,N_43192,N_44532);
and U45195 (N_45195,N_44283,N_44914);
or U45196 (N_45196,N_43776,N_44204);
nor U45197 (N_45197,N_41615,N_40152);
or U45198 (N_45198,N_41711,N_41067);
or U45199 (N_45199,N_41255,N_42823);
xnor U45200 (N_45200,N_40179,N_42475);
nor U45201 (N_45201,N_43744,N_40502);
or U45202 (N_45202,N_43479,N_42331);
nor U45203 (N_45203,N_42995,N_40941);
or U45204 (N_45204,N_43989,N_41736);
and U45205 (N_45205,N_43535,N_43891);
xnor U45206 (N_45206,N_40001,N_41980);
nand U45207 (N_45207,N_40630,N_43838);
and U45208 (N_45208,N_41132,N_44786);
nand U45209 (N_45209,N_41211,N_40619);
or U45210 (N_45210,N_43933,N_43117);
and U45211 (N_45211,N_42837,N_41695);
and U45212 (N_45212,N_44530,N_43206);
nand U45213 (N_45213,N_44173,N_43398);
nor U45214 (N_45214,N_42360,N_44149);
xor U45215 (N_45215,N_44187,N_44376);
nand U45216 (N_45216,N_41375,N_41430);
xnor U45217 (N_45217,N_41507,N_44589);
nor U45218 (N_45218,N_40229,N_44889);
nor U45219 (N_45219,N_44339,N_42135);
and U45220 (N_45220,N_43793,N_40245);
nand U45221 (N_45221,N_41438,N_41511);
nor U45222 (N_45222,N_44362,N_40012);
nor U45223 (N_45223,N_42439,N_42283);
nand U45224 (N_45224,N_43783,N_41180);
and U45225 (N_45225,N_40632,N_41710);
nor U45226 (N_45226,N_41167,N_42280);
and U45227 (N_45227,N_44324,N_43138);
nor U45228 (N_45228,N_42309,N_40601);
nand U45229 (N_45229,N_41601,N_44254);
nand U45230 (N_45230,N_40460,N_44260);
or U45231 (N_45231,N_43028,N_41676);
nand U45232 (N_45232,N_42726,N_42897);
nand U45233 (N_45233,N_40060,N_41254);
xor U45234 (N_45234,N_44908,N_43221);
nand U45235 (N_45235,N_40019,N_43571);
or U45236 (N_45236,N_42782,N_41855);
nand U45237 (N_45237,N_41693,N_43854);
nor U45238 (N_45238,N_44347,N_40320);
xnor U45239 (N_45239,N_41253,N_44540);
nand U45240 (N_45240,N_43920,N_40167);
nor U45241 (N_45241,N_42787,N_40217);
xor U45242 (N_45242,N_40528,N_43572);
xnor U45243 (N_45243,N_42951,N_40879);
nand U45244 (N_45244,N_41033,N_41111);
and U45245 (N_45245,N_43443,N_42290);
or U45246 (N_45246,N_41181,N_41022);
nor U45247 (N_45247,N_41409,N_42597);
or U45248 (N_45248,N_42619,N_44871);
or U45249 (N_45249,N_41999,N_44291);
nand U45250 (N_45250,N_43078,N_43990);
xnor U45251 (N_45251,N_40683,N_43799);
or U45252 (N_45252,N_42676,N_40812);
nand U45253 (N_45253,N_41714,N_42074);
and U45254 (N_45254,N_43876,N_42426);
nor U45255 (N_45255,N_43233,N_40390);
nor U45256 (N_45256,N_44562,N_42175);
nor U45257 (N_45257,N_44276,N_44030);
nor U45258 (N_45258,N_42584,N_44699);
nand U45259 (N_45259,N_41549,N_42043);
or U45260 (N_45260,N_43368,N_40541);
xor U45261 (N_45261,N_42301,N_40735);
nand U45262 (N_45262,N_41551,N_40562);
or U45263 (N_45263,N_42079,N_44209);
or U45264 (N_45264,N_41075,N_41162);
nor U45265 (N_45265,N_41704,N_43770);
and U45266 (N_45266,N_40365,N_40403);
xnor U45267 (N_45267,N_44715,N_43213);
nor U45268 (N_45268,N_44812,N_40026);
and U45269 (N_45269,N_40934,N_43807);
nand U45270 (N_45270,N_40523,N_41011);
xnor U45271 (N_45271,N_42345,N_43143);
and U45272 (N_45272,N_41528,N_43291);
nor U45273 (N_45273,N_44887,N_40926);
and U45274 (N_45274,N_41893,N_42725);
xnor U45275 (N_45275,N_42332,N_42206);
or U45276 (N_45276,N_42894,N_41505);
and U45277 (N_45277,N_43015,N_41239);
or U45278 (N_45278,N_44595,N_43871);
xor U45279 (N_45279,N_40163,N_44960);
nor U45280 (N_45280,N_41109,N_40119);
xor U45281 (N_45281,N_40897,N_44329);
and U45282 (N_45282,N_40362,N_42455);
or U45283 (N_45283,N_44733,N_44978);
nor U45284 (N_45284,N_41906,N_44825);
nor U45285 (N_45285,N_43239,N_42555);
nand U45286 (N_45286,N_40883,N_40258);
nand U45287 (N_45287,N_41080,N_43832);
nand U45288 (N_45288,N_42996,N_43668);
nor U45289 (N_45289,N_42467,N_40187);
and U45290 (N_45290,N_40049,N_44884);
xnor U45291 (N_45291,N_44344,N_43666);
nand U45292 (N_45292,N_43827,N_41130);
nand U45293 (N_45293,N_43530,N_43558);
nand U45294 (N_45294,N_43381,N_42684);
nor U45295 (N_45295,N_42070,N_42226);
nand U45296 (N_45296,N_42880,N_40234);
nor U45297 (N_45297,N_40123,N_40481);
xor U45298 (N_45298,N_40180,N_40255);
nor U45299 (N_45299,N_42065,N_42321);
nand U45300 (N_45300,N_41439,N_43682);
or U45301 (N_45301,N_40886,N_41085);
nor U45302 (N_45302,N_43655,N_40397);
xnor U45303 (N_45303,N_44490,N_40376);
nor U45304 (N_45304,N_40008,N_41990);
nor U45305 (N_45305,N_41763,N_41073);
xor U45306 (N_45306,N_41450,N_41531);
and U45307 (N_45307,N_44489,N_43419);
nor U45308 (N_45308,N_42285,N_43611);
or U45309 (N_45309,N_40014,N_40085);
and U45310 (N_45310,N_43965,N_43413);
and U45311 (N_45311,N_44133,N_43992);
and U45312 (N_45312,N_42604,N_41606);
or U45313 (N_45313,N_40555,N_41788);
or U45314 (N_45314,N_43565,N_43841);
xor U45315 (N_45315,N_43049,N_42559);
and U45316 (N_45316,N_42133,N_41388);
nor U45317 (N_45317,N_44874,N_42883);
or U45318 (N_45318,N_44106,N_44464);
and U45319 (N_45319,N_44193,N_44742);
xor U45320 (N_45320,N_43163,N_42769);
nor U45321 (N_45321,N_42396,N_43707);
nand U45322 (N_45322,N_41262,N_42616);
and U45323 (N_45323,N_42998,N_42150);
nand U45324 (N_45324,N_41122,N_42340);
or U45325 (N_45325,N_40294,N_41460);
nor U45326 (N_45326,N_40618,N_40337);
and U45327 (N_45327,N_40321,N_42297);
or U45328 (N_45328,N_44145,N_42514);
nor U45329 (N_45329,N_41809,N_42381);
xnor U45330 (N_45330,N_44995,N_40760);
nand U45331 (N_45331,N_40993,N_40251);
nand U45332 (N_45332,N_41422,N_42802);
nor U45333 (N_45333,N_40928,N_43296);
or U45334 (N_45334,N_40448,N_41231);
xnor U45335 (N_45335,N_41787,N_40453);
or U45336 (N_45336,N_40635,N_42208);
nor U45337 (N_45337,N_42575,N_42253);
nor U45338 (N_45338,N_44226,N_44076);
or U45339 (N_45339,N_41213,N_43014);
and U45340 (N_45340,N_41831,N_41489);
nand U45341 (N_45341,N_44768,N_42852);
or U45342 (N_45342,N_43787,N_42261);
and U45343 (N_45343,N_41708,N_42881);
xor U45344 (N_45344,N_44642,N_44900);
and U45345 (N_45345,N_42459,N_40723);
and U45346 (N_45346,N_44920,N_42512);
xor U45347 (N_45347,N_43897,N_41009);
or U45348 (N_45348,N_40218,N_41477);
or U45349 (N_45349,N_43096,N_42975);
or U45350 (N_45350,N_42879,N_43142);
or U45351 (N_45351,N_41914,N_43639);
nand U45352 (N_45352,N_44229,N_44778);
or U45353 (N_45353,N_41706,N_40821);
xor U45354 (N_45354,N_40518,N_41930);
nor U45355 (N_45355,N_43801,N_42936);
and U45356 (N_45356,N_44100,N_44300);
nor U45357 (N_45357,N_43603,N_42824);
nand U45358 (N_45358,N_43979,N_44691);
and U45359 (N_45359,N_43362,N_43231);
and U45360 (N_45360,N_43642,N_41716);
xnor U45361 (N_45361,N_42146,N_42325);
and U45362 (N_45362,N_42276,N_44906);
nand U45363 (N_45363,N_43119,N_40018);
nand U45364 (N_45364,N_43115,N_44615);
xnor U45365 (N_45365,N_40780,N_43914);
or U45366 (N_45366,N_42462,N_44793);
and U45367 (N_45367,N_43195,N_42031);
nor U45368 (N_45368,N_44568,N_40076);
or U45369 (N_45369,N_41106,N_42814);
nor U45370 (N_45370,N_42193,N_43742);
nor U45371 (N_45371,N_44205,N_42507);
xnor U45372 (N_45372,N_44309,N_43872);
nand U45373 (N_45373,N_40782,N_42800);
nand U45374 (N_45374,N_44741,N_40352);
and U45375 (N_45375,N_42131,N_41440);
and U45376 (N_45376,N_40730,N_40725);
nand U45377 (N_45377,N_42144,N_43228);
nor U45378 (N_45378,N_43194,N_44181);
nor U45379 (N_45379,N_42844,N_40987);
and U45380 (N_45380,N_43991,N_41366);
nor U45381 (N_45381,N_43918,N_42406);
xnor U45382 (N_45382,N_44513,N_42552);
and U45383 (N_45383,N_42127,N_42964);
nand U45384 (N_45384,N_43763,N_41121);
xnor U45385 (N_45385,N_41633,N_40285);
xnor U45386 (N_45386,N_41296,N_43833);
nor U45387 (N_45387,N_42491,N_44119);
or U45388 (N_45388,N_42310,N_42323);
and U45389 (N_45389,N_43881,N_44466);
or U45390 (N_45390,N_40353,N_43686);
or U45391 (N_45391,N_41926,N_42773);
nand U45392 (N_45392,N_43462,N_44199);
xnor U45393 (N_45393,N_43485,N_42215);
or U45394 (N_45394,N_41242,N_41237);
or U45395 (N_45395,N_42739,N_42210);
and U45396 (N_45396,N_44160,N_44894);
nand U45397 (N_45397,N_40145,N_43280);
and U45398 (N_45398,N_44103,N_44046);
xnor U45399 (N_45399,N_44483,N_40126);
xor U45400 (N_45400,N_42393,N_40671);
xor U45401 (N_45401,N_44599,N_43406);
and U45402 (N_45402,N_43200,N_41068);
nor U45403 (N_45403,N_40870,N_42212);
nand U45404 (N_45404,N_43484,N_44677);
nand U45405 (N_45405,N_41729,N_40830);
and U45406 (N_45406,N_43710,N_41671);
and U45407 (N_45407,N_43355,N_40980);
xor U45408 (N_45408,N_41314,N_40446);
nand U45409 (N_45409,N_44433,N_40522);
nand U45410 (N_45410,N_40264,N_44542);
and U45411 (N_45411,N_40843,N_43848);
nor U45412 (N_45412,N_43256,N_42030);
or U45413 (N_45413,N_42091,N_40617);
nand U45414 (N_45414,N_43574,N_42049);
or U45415 (N_45415,N_43576,N_40044);
nor U45416 (N_45416,N_40262,N_43041);
or U45417 (N_45417,N_40547,N_41119);
nand U45418 (N_45418,N_43125,N_41277);
xnor U45419 (N_45419,N_42807,N_42577);
or U45420 (N_45420,N_43442,N_44591);
or U45421 (N_45421,N_44569,N_40111);
xor U45422 (N_45422,N_43002,N_40973);
nor U45423 (N_45423,N_41987,N_41101);
nand U45424 (N_45424,N_42644,N_43247);
or U45425 (N_45425,N_44154,N_44321);
xor U45426 (N_45426,N_40374,N_42677);
nor U45427 (N_45427,N_44262,N_43698);
nor U45428 (N_45428,N_41750,N_44751);
and U45429 (N_45429,N_44110,N_40013);
or U45430 (N_45430,N_43943,N_43430);
nand U45431 (N_45431,N_40641,N_43508);
nand U45432 (N_45432,N_44468,N_41029);
xor U45433 (N_45433,N_42005,N_43087);
nor U45434 (N_45434,N_43510,N_44086);
and U45435 (N_45435,N_44566,N_43948);
nand U45436 (N_45436,N_42592,N_41686);
or U45437 (N_45437,N_42923,N_43075);
nor U45438 (N_45438,N_44518,N_42812);
and U45439 (N_45439,N_40133,N_43491);
and U45440 (N_45440,N_43534,N_44946);
or U45441 (N_45441,N_43382,N_44665);
nand U45442 (N_45442,N_44040,N_44416);
nand U45443 (N_45443,N_40366,N_43236);
xor U45444 (N_45444,N_40552,N_40597);
nand U45445 (N_45445,N_44559,N_42937);
nor U45446 (N_45446,N_44307,N_41042);
and U45447 (N_45447,N_44575,N_41915);
xor U45448 (N_45448,N_44656,N_43538);
xnor U45449 (N_45449,N_43211,N_43171);
nand U45450 (N_45450,N_43284,N_44310);
xnor U45451 (N_45451,N_44312,N_44074);
nor U45452 (N_45452,N_44824,N_42129);
nand U45453 (N_45453,N_42246,N_41961);
xor U45454 (N_45454,N_42929,N_41293);
or U45455 (N_45455,N_43165,N_44964);
nand U45456 (N_45456,N_42352,N_42191);
xor U45457 (N_45457,N_42941,N_43309);
nand U45458 (N_45458,N_40373,N_44661);
xnor U45459 (N_45459,N_41723,N_43853);
nor U45460 (N_45460,N_42147,N_44128);
or U45461 (N_45461,N_40770,N_42412);
nand U45462 (N_45462,N_43295,N_44403);
nand U45463 (N_45463,N_40144,N_44737);
or U45464 (N_45464,N_40256,N_43108);
or U45465 (N_45465,N_42084,N_44840);
and U45466 (N_45466,N_40933,N_43395);
or U45467 (N_45467,N_44669,N_41103);
nor U45468 (N_45468,N_42902,N_40203);
xnor U45469 (N_45469,N_44857,N_43752);
xor U45470 (N_45470,N_40214,N_41593);
and U45471 (N_45471,N_44724,N_43759);
nand U45472 (N_45472,N_43489,N_41513);
and U45473 (N_45473,N_43847,N_40192);
xor U45474 (N_45474,N_41444,N_44012);
and U45475 (N_45475,N_41604,N_40579);
nor U45476 (N_45476,N_40602,N_43375);
xor U45477 (N_45477,N_44535,N_41090);
nand U45478 (N_45478,N_44379,N_40894);
xnor U45479 (N_45479,N_44412,N_42354);
nor U45480 (N_45480,N_43665,N_40427);
and U45481 (N_45481,N_42476,N_41027);
or U45482 (N_45482,N_43416,N_44411);
nand U45483 (N_45483,N_44929,N_44430);
nand U45484 (N_45484,N_43708,N_41696);
or U45485 (N_45485,N_41636,N_41651);
or U45486 (N_45486,N_44558,N_42913);
or U45487 (N_45487,N_43012,N_43136);
nand U45488 (N_45488,N_40236,N_43450);
nor U45489 (N_45489,N_41847,N_42453);
nand U45490 (N_45490,N_42055,N_44278);
xnor U45491 (N_45491,N_43466,N_44853);
or U45492 (N_45492,N_40286,N_43123);
xnor U45493 (N_45493,N_43046,N_43440);
xor U45494 (N_45494,N_42389,N_43966);
xnor U45495 (N_45495,N_43870,N_40960);
or U45496 (N_45496,N_42275,N_42237);
or U45497 (N_45497,N_43902,N_42052);
or U45498 (N_45498,N_40824,N_44955);
or U45499 (N_45499,N_44604,N_41335);
nor U45500 (N_45500,N_40077,N_44034);
nand U45501 (N_45501,N_44332,N_41051);
or U45502 (N_45502,N_42008,N_42833);
and U45503 (N_45503,N_42942,N_41287);
or U45504 (N_45504,N_42108,N_43901);
nand U45505 (N_45505,N_40109,N_43511);
nor U45506 (N_45506,N_42926,N_42589);
and U45507 (N_45507,N_44408,N_44985);
nor U45508 (N_45508,N_40450,N_40797);
and U45509 (N_45509,N_42813,N_44109);
nor U45510 (N_45510,N_40738,N_44233);
and U45511 (N_45511,N_44740,N_42225);
or U45512 (N_45512,N_44578,N_41433);
nand U45513 (N_45513,N_44389,N_41039);
nor U45514 (N_45514,N_40775,N_40868);
and U45515 (N_45515,N_43556,N_41235);
or U45516 (N_45516,N_41638,N_42292);
or U45517 (N_45517,N_40516,N_44512);
or U45518 (N_45518,N_42859,N_44289);
or U45519 (N_45519,N_44941,N_41888);
and U45520 (N_45520,N_43240,N_43204);
xor U45521 (N_45521,N_43741,N_43345);
nand U45522 (N_45522,N_43721,N_40006);
nand U45523 (N_45523,N_43314,N_42402);
xnor U45524 (N_45524,N_40116,N_40990);
nor U45525 (N_45525,N_40515,N_40195);
nand U45526 (N_45526,N_44653,N_44870);
nor U45527 (N_45527,N_40715,N_40807);
nor U45528 (N_45528,N_40832,N_44798);
and U45529 (N_45529,N_43409,N_43190);
nor U45530 (N_45530,N_43946,N_40947);
nor U45531 (N_45531,N_44822,N_42609);
nor U45532 (N_45532,N_43003,N_42050);
or U45533 (N_45533,N_44153,N_42039);
xor U45534 (N_45534,N_44703,N_40270);
xnor U45535 (N_45535,N_40067,N_41541);
xnor U45536 (N_45536,N_42900,N_44280);
nand U45537 (N_45537,N_40504,N_42333);
and U45538 (N_45538,N_42251,N_43540);
xnor U45539 (N_45539,N_43122,N_42407);
and U45540 (N_45540,N_42685,N_43973);
xnor U45541 (N_45541,N_40651,N_42885);
and U45542 (N_45542,N_42270,N_40407);
nor U45543 (N_45543,N_42448,N_43702);
xor U45544 (N_45544,N_40606,N_43196);
or U45545 (N_45545,N_40835,N_42786);
nor U45546 (N_45546,N_40061,N_42404);
or U45547 (N_45547,N_43267,N_41841);
nor U45548 (N_45548,N_41652,N_40064);
or U45549 (N_45549,N_41304,N_42487);
nor U45550 (N_45550,N_44495,N_44902);
or U45551 (N_45551,N_40425,N_42960);
xnor U45552 (N_45552,N_41118,N_40744);
xor U45553 (N_45553,N_42694,N_44177);
or U45554 (N_45554,N_41577,N_44471);
xnor U45555 (N_45555,N_41952,N_44049);
nor U45556 (N_45556,N_41960,N_42494);
nand U45557 (N_45557,N_43922,N_43069);
xor U45558 (N_45558,N_40844,N_44237);
or U45559 (N_45559,N_41929,N_44479);
nor U45560 (N_45560,N_40041,N_41041);
xor U45561 (N_45561,N_40732,N_44269);
and U45562 (N_45562,N_43318,N_43816);
and U45563 (N_45563,N_42495,N_44270);
xor U45564 (N_45564,N_44587,N_44572);
or U45565 (N_45565,N_40224,N_41389);
and U45566 (N_45566,N_42822,N_42518);
or U45567 (N_45567,N_42612,N_43057);
and U45568 (N_45568,N_40074,N_44910);
nand U45569 (N_45569,N_40161,N_43421);
or U45570 (N_45570,N_43155,N_42750);
and U45571 (N_45571,N_41858,N_44850);
xnor U45572 (N_45572,N_40854,N_41030);
nor U45573 (N_45573,N_44440,N_41472);
and U45574 (N_45574,N_41545,N_41456);
nor U45575 (N_45575,N_42170,N_41981);
xor U45576 (N_45576,N_42637,N_42286);
nor U45577 (N_45577,N_43915,N_43023);
or U45578 (N_45578,N_42980,N_40509);
nand U45579 (N_45579,N_43788,N_43166);
xnor U45580 (N_45580,N_44522,N_42783);
xor U45581 (N_45581,N_44810,N_42511);
xnor U45582 (N_45582,N_43444,N_44317);
xnor U45583 (N_45583,N_41236,N_42296);
nor U45584 (N_45584,N_44138,N_42411);
and U45585 (N_45585,N_41697,N_44271);
nand U45586 (N_45586,N_40796,N_41059);
nor U45587 (N_45587,N_40052,N_40778);
or U45588 (N_45588,N_40257,N_40645);
xnor U45589 (N_45589,N_40621,N_40086);
and U45590 (N_45590,N_43229,N_40838);
nand U45591 (N_45591,N_40644,N_44377);
nor U45592 (N_45592,N_40789,N_42516);
xnor U45593 (N_45593,N_44721,N_40045);
nand U45594 (N_45594,N_43730,N_40456);
nand U45595 (N_45595,N_43065,N_42136);
or U45596 (N_45596,N_40539,N_44343);
or U45597 (N_45597,N_41772,N_40219);
xor U45598 (N_45598,N_44706,N_40445);
or U45599 (N_45599,N_44286,N_40033);
nor U45600 (N_45600,N_40704,N_42624);
nand U45601 (N_45601,N_43114,N_44225);
nor U45602 (N_45602,N_40433,N_43016);
or U45603 (N_45603,N_44649,N_40084);
and U45604 (N_45604,N_42479,N_40590);
nand U45605 (N_45605,N_41386,N_42198);
and U45606 (N_45606,N_42572,N_42339);
and U45607 (N_45607,N_43527,N_41396);
and U45608 (N_45608,N_40925,N_43216);
xor U45609 (N_45609,N_43560,N_43127);
nor U45610 (N_45610,N_40291,N_42126);
nand U45611 (N_45611,N_40795,N_40490);
xnor U45612 (N_45612,N_43077,N_44732);
nand U45613 (N_45613,N_43843,N_43302);
nor U45614 (N_45614,N_43133,N_43888);
nor U45615 (N_45615,N_41149,N_43674);
nor U45616 (N_45616,N_41074,N_41476);
or U45617 (N_45617,N_43113,N_43305);
and U45618 (N_45618,N_44776,N_44981);
and U45619 (N_45619,N_44157,N_42349);
nand U45620 (N_45620,N_42772,N_43401);
nand U45621 (N_45621,N_44116,N_44378);
and U45622 (N_45622,N_44081,N_43219);
nand U45623 (N_45623,N_42568,N_44580);
or U45624 (N_45624,N_43771,N_43439);
xor U45625 (N_45625,N_42383,N_43588);
and U45626 (N_45626,N_40568,N_44816);
nor U45627 (N_45627,N_44462,N_41365);
nor U45628 (N_45628,N_44972,N_41424);
and U45629 (N_45629,N_43646,N_41001);
nand U45630 (N_45630,N_42853,N_44244);
xor U45631 (N_45631,N_44621,N_41088);
nand U45632 (N_45632,N_43930,N_40211);
xnor U45633 (N_45633,N_43047,N_44125);
nand U45634 (N_45634,N_43469,N_42374);
or U45635 (N_45635,N_43697,N_43579);
nor U45636 (N_45636,N_40766,N_42009);
and U45637 (N_45637,N_44797,N_42643);
nand U45638 (N_45638,N_44965,N_44526);
nor U45639 (N_45639,N_40627,N_40669);
nor U45640 (N_45640,N_42890,N_40565);
or U45641 (N_45641,N_44679,N_41488);
nand U45642 (N_45642,N_40338,N_44645);
nor U45643 (N_45643,N_44790,N_43828);
nor U45644 (N_45644,N_41547,N_41598);
nor U45645 (N_45645,N_43537,N_41530);
nand U45646 (N_45646,N_41584,N_44577);
or U45647 (N_45647,N_43197,N_44878);
nor U45648 (N_45648,N_43813,N_42011);
xnor U45649 (N_45649,N_44176,N_42218);
nor U45650 (N_45650,N_40707,N_41491);
and U45651 (N_45651,N_40132,N_41607);
nand U45652 (N_45652,N_43688,N_44760);
nand U45653 (N_45653,N_44596,N_44327);
xor U45654 (N_45654,N_44235,N_40350);
nor U45655 (N_45655,N_44939,N_42660);
or U45656 (N_45656,N_44057,N_42795);
xnor U45657 (N_45657,N_43913,N_43325);
nand U45658 (N_45658,N_41724,N_41995);
xnor U45659 (N_45659,N_41359,N_42959);
and U45660 (N_45660,N_40332,N_40166);
xnor U45661 (N_45661,N_42699,N_40375);
xnor U45662 (N_45662,N_42528,N_44890);
nand U45663 (N_45663,N_44467,N_40065);
nor U45664 (N_45664,N_43347,N_44556);
nand U45665 (N_45665,N_41554,N_44407);
nor U45666 (N_45666,N_42779,N_41938);
and U45667 (N_45667,N_43536,N_41368);
nor U45668 (N_45668,N_43339,N_40995);
or U45669 (N_45669,N_43883,N_43927);
and U45670 (N_45670,N_44094,N_43999);
nor U45671 (N_45671,N_40949,N_43208);
nand U45672 (N_45672,N_43941,N_43690);
xnor U45673 (N_45673,N_41499,N_40979);
and U45674 (N_45674,N_44473,N_40578);
xnor U45675 (N_45675,N_44427,N_43384);
and U45676 (N_45676,N_42327,N_44633);
nand U45677 (N_45677,N_40512,N_40953);
nand U45678 (N_45678,N_42416,N_40637);
and U45679 (N_45679,N_41166,N_41229);
nor U45680 (N_45680,N_44827,N_41936);
xnor U45681 (N_45681,N_42054,N_44429);
nor U45682 (N_45682,N_42348,N_43380);
xor U45683 (N_45683,N_40623,N_40753);
nor U45684 (N_45684,N_43011,N_42710);
and U45685 (N_45685,N_40740,N_41782);
nor U45686 (N_45686,N_42505,N_40422);
nor U45687 (N_45687,N_42468,N_42569);
xnor U45688 (N_45688,N_44163,N_44883);
xor U45689 (N_45689,N_41274,N_41202);
nand U45690 (N_45690,N_42622,N_43453);
or U45691 (N_45691,N_41310,N_40777);
xor U45692 (N_45692,N_42832,N_40135);
and U45693 (N_45693,N_42087,N_43718);
nor U45694 (N_45694,N_43935,N_40025);
nand U45695 (N_45695,N_43500,N_42291);
nand U45696 (N_45696,N_40867,N_42588);
xor U45697 (N_45697,N_42137,N_42888);
xnor U45698 (N_45698,N_44420,N_44428);
nand U45699 (N_45699,N_43617,N_42256);
nor U45700 (N_45700,N_41657,N_44627);
xor U45701 (N_45701,N_43022,N_41197);
or U45702 (N_45702,N_40743,N_41744);
and U45703 (N_45703,N_43671,N_42234);
nor U45704 (N_45704,N_43423,N_40662);
nor U45705 (N_45705,N_41208,N_43056);
nor U45706 (N_45706,N_43032,N_43623);
nand U45707 (N_45707,N_44421,N_40325);
xor U45708 (N_45708,N_42874,N_41864);
and U45709 (N_45709,N_43066,N_41836);
nand U45710 (N_45710,N_40479,N_42477);
xor U45711 (N_45711,N_40185,N_43408);
xor U45712 (N_45712,N_44682,N_41537);
nor U45713 (N_45713,N_44451,N_43525);
and U45714 (N_45714,N_41678,N_43947);
and U45715 (N_45715,N_44838,N_44533);
and U45716 (N_45716,N_42259,N_41781);
nor U45717 (N_45717,N_43083,N_41908);
nor U45718 (N_45718,N_44719,N_40556);
or U45719 (N_45719,N_41969,N_44631);
nand U45720 (N_45720,N_44928,N_43615);
nor U45721 (N_45721,N_42012,N_42264);
nand U45722 (N_45722,N_41308,N_44534);
and U45723 (N_45723,N_42351,N_40964);
xor U45724 (N_45724,N_41270,N_41493);
nor U45725 (N_45725,N_43907,N_43293);
and U45726 (N_45726,N_42875,N_42729);
and U45727 (N_45727,N_40998,N_42978);
nor U45728 (N_45728,N_42481,N_41196);
or U45729 (N_45729,N_40073,N_43322);
nor U45730 (N_45730,N_40387,N_42017);
or U45731 (N_45731,N_40174,N_42148);
and U45732 (N_45732,N_42673,N_41532);
nor U45733 (N_45733,N_40948,N_44581);
xor U45734 (N_45734,N_42258,N_40997);
and U45735 (N_45735,N_43082,N_42990);
nand U45736 (N_45736,N_40534,N_44146);
and U45737 (N_45737,N_41179,N_42308);
xor U45738 (N_45738,N_42864,N_40545);
and U45739 (N_45739,N_42536,N_42496);
or U45740 (N_45740,N_44780,N_42281);
or U45741 (N_45741,N_43551,N_42249);
and U45742 (N_45742,N_42781,N_41749);
and U45743 (N_45743,N_43543,N_42958);
xor U45744 (N_45744,N_44608,N_42419);
nand U45745 (N_45745,N_43567,N_41660);
xor U45746 (N_45746,N_44885,N_43612);
nand U45747 (N_45747,N_41924,N_40691);
nor U45748 (N_45748,N_40875,N_41951);
nand U45749 (N_45749,N_41644,N_40355);
and U45750 (N_45750,N_43512,N_40902);
or U45751 (N_45751,N_44236,N_40050);
nor U45752 (N_45752,N_43573,N_42910);
nor U45753 (N_45753,N_44249,N_42397);
xnor U45754 (N_45754,N_42432,N_43277);
nor U45755 (N_45755,N_40554,N_41533);
nor U45756 (N_45756,N_41474,N_44019);
or U45757 (N_45757,N_43593,N_44944);
nand U45758 (N_45758,N_40977,N_41909);
and U45759 (N_45759,N_44936,N_42233);
or U45760 (N_45760,N_43675,N_42545);
and U45761 (N_45761,N_41568,N_40398);
or U45762 (N_45762,N_40663,N_40688);
nor U45763 (N_45763,N_44342,N_44612);
or U45764 (N_45764,N_44987,N_42600);
or U45765 (N_45765,N_41759,N_43997);
nor U45766 (N_45766,N_40382,N_40066);
or U45767 (N_45767,N_44053,N_43445);
and U45768 (N_45768,N_44932,N_42842);
nand U45769 (N_45769,N_41193,N_42207);
or U45770 (N_45770,N_42174,N_42525);
xnor U45771 (N_45771,N_44005,N_44622);
or U45772 (N_45772,N_44635,N_42590);
and U45773 (N_45773,N_40232,N_44769);
and U45774 (N_45774,N_41912,N_44228);
and U45775 (N_45775,N_40209,N_42809);
xor U45776 (N_45776,N_42473,N_43102);
nor U45777 (N_45777,N_43139,N_44766);
or U45778 (N_45778,N_44121,N_44895);
xor U45779 (N_45779,N_43242,N_40082);
xnor U45780 (N_45780,N_43227,N_42704);
and U45781 (N_45781,N_40169,N_43311);
or U45782 (N_45782,N_43986,N_44898);
and U45783 (N_45783,N_41819,N_44820);
nor U45784 (N_45784,N_40094,N_43035);
or U45785 (N_45785,N_41931,N_43923);
nand U45786 (N_45786,N_41918,N_40811);
nand U45787 (N_45787,N_44431,N_41794);
or U45788 (N_45788,N_42399,N_42909);
nor U45789 (N_45789,N_42415,N_40113);
xnor U45790 (N_45790,N_43374,N_40042);
nand U45791 (N_45791,N_40147,N_44866);
nand U45792 (N_45792,N_40992,N_41883);
or U45793 (N_45793,N_42806,N_41353);
nand U45794 (N_45794,N_41176,N_41610);
nand U45795 (N_45795,N_41614,N_41061);
nor U45796 (N_45796,N_41717,N_44945);
xor U45797 (N_45797,N_41425,N_42247);
xnor U45798 (N_45798,N_44414,N_44015);
nor U45799 (N_45799,N_42240,N_40815);
nor U45800 (N_45800,N_42168,N_41261);
xnor U45801 (N_45801,N_40510,N_40196);
xor U45802 (N_45802,N_41741,N_42387);
nor U45803 (N_45803,N_40117,N_40679);
nor U45804 (N_45804,N_42120,N_40303);
nor U45805 (N_45805,N_41071,N_41451);
xor U45806 (N_45806,N_42991,N_40913);
nand U45807 (N_45807,N_41845,N_43679);
or U45808 (N_45808,N_42350,N_41583);
xor U45809 (N_45809,N_42527,N_42042);
nand U45810 (N_45810,N_40661,N_41046);
or U45811 (N_45811,N_42033,N_40305);
xnor U45812 (N_45812,N_40199,N_40413);
xor U45813 (N_45813,N_42141,N_40227);
xnor U45814 (N_45814,N_41768,N_40672);
and U45815 (N_45815,N_41989,N_42605);
xor U45816 (N_45816,N_43890,N_43831);
xnor U45817 (N_45817,N_42914,N_41324);
and U45818 (N_45818,N_43391,N_42889);
and U45819 (N_45819,N_41363,N_42865);
nand U45820 (N_45820,N_41756,N_40681);
and U45821 (N_45821,N_41479,N_40988);
xnor U45822 (N_45822,N_41791,N_40063);
nor U45823 (N_45823,N_44171,N_40304);
xnor U45824 (N_45824,N_41963,N_40874);
and U45825 (N_45825,N_41595,N_42939);
and U45826 (N_45826,N_43105,N_44139);
and U45827 (N_45827,N_42094,N_43640);
nand U45828 (N_45828,N_42375,N_44698);
nor U45829 (N_45829,N_42804,N_40648);
or U45830 (N_45830,N_42230,N_41342);
and U45831 (N_45831,N_42664,N_44950);
and U45832 (N_45832,N_40057,N_41340);
nor U45833 (N_45833,N_42994,N_43424);
nor U45834 (N_45834,N_43461,N_41204);
nor U45835 (N_45835,N_41628,N_42971);
nand U45836 (N_45836,N_41755,N_40608);
nand U45837 (N_45837,N_40955,N_43779);
nand U45838 (N_45838,N_40869,N_43932);
nand U45839 (N_45839,N_40557,N_42395);
or U45840 (N_45840,N_40091,N_43756);
nor U45841 (N_45841,N_43684,N_44168);
nor U45842 (N_45842,N_44493,N_42963);
or U45843 (N_45843,N_43438,N_42887);
nor U45844 (N_45844,N_40864,N_43225);
and U45845 (N_45845,N_41138,N_44655);
or U45846 (N_45846,N_43856,N_43412);
or U45847 (N_45847,N_42759,N_44214);
nor U45848 (N_45848,N_44201,N_43931);
nor U45849 (N_45849,N_40323,N_43939);
or U45850 (N_45850,N_43168,N_40364);
nand U45851 (N_45851,N_41273,N_42510);
nor U45852 (N_45852,N_44303,N_42893);
nand U45853 (N_45853,N_41240,N_41948);
or U45854 (N_45854,N_41575,N_40324);
xor U45855 (N_45855,N_43018,N_40702);
and U45856 (N_45856,N_41535,N_41200);
nor U45857 (N_45857,N_41228,N_41352);
nor U45858 (N_45858,N_40930,N_42917);
and U45859 (N_45859,N_40078,N_44841);
nand U45860 (N_45860,N_41435,N_41643);
and U45861 (N_45861,N_44250,N_43619);
or U45862 (N_45862,N_42076,N_44334);
and U45863 (N_45863,N_40474,N_41302);
nor U45864 (N_45864,N_43457,N_40279);
nand U45865 (N_45865,N_44988,N_41445);
nand U45866 (N_45866,N_40756,N_41165);
nor U45867 (N_45867,N_42662,N_43360);
xnor U45868 (N_45868,N_44977,N_40372);
xor U45869 (N_45869,N_41789,N_40092);
or U45870 (N_45870,N_41413,N_40080);
nor U45871 (N_45871,N_40363,N_40468);
xor U45872 (N_45872,N_42715,N_41691);
nor U45873 (N_45873,N_40265,N_44845);
and U45874 (N_45874,N_44957,N_44158);
or U45875 (N_45875,N_43201,N_40488);
nor U45876 (N_45876,N_44085,N_41815);
nand U45877 (N_45877,N_40148,N_44861);
nand U45878 (N_45878,N_44974,N_44370);
or U45879 (N_45879,N_41713,N_44413);
nand U45880 (N_45880,N_44392,N_40771);
nand U45881 (N_45881,N_44222,N_42303);
nor U45882 (N_45882,N_40946,N_43553);
nor U45883 (N_45883,N_43315,N_41004);
nand U45884 (N_45884,N_42596,N_43531);
nor U45885 (N_45885,N_44646,N_42734);
nor U45886 (N_45886,N_43737,N_43425);
nor U45887 (N_45887,N_44975,N_43458);
or U45888 (N_45888,N_42789,N_44337);
or U45889 (N_45889,N_41325,N_44802);
nor U45890 (N_45890,N_41332,N_44882);
and U45891 (N_45891,N_44593,N_44658);
xnor U45892 (N_45892,N_40705,N_40610);
xnor U45893 (N_45893,N_43908,N_42707);
nand U45894 (N_45894,N_43153,N_43693);
or U45895 (N_45895,N_42793,N_43587);
xnor U45896 (N_45896,N_41275,N_40837);
xnor U45897 (N_45897,N_42143,N_40675);
nand U45898 (N_45898,N_40241,N_41550);
nor U45899 (N_45899,N_40386,N_41631);
or U45900 (N_45900,N_43051,N_42719);
xnor U45901 (N_45901,N_40865,N_42370);
nand U45902 (N_45902,N_44141,N_43369);
xnor U45903 (N_45903,N_42027,N_44364);
xor U45904 (N_45904,N_41108,N_40529);
nor U45905 (N_45905,N_40400,N_44357);
or U45906 (N_45906,N_41849,N_44221);
or U45907 (N_45907,N_44501,N_40709);
or U45908 (N_45908,N_42678,N_42896);
nor U45909 (N_45909,N_42138,N_42675);
nor U45910 (N_45910,N_40207,N_41770);
nor U45911 (N_45911,N_43959,N_40765);
or U45912 (N_45912,N_42177,N_42334);
or U45913 (N_45913,N_41783,N_44876);
or U45914 (N_45914,N_41825,N_42110);
nor U45915 (N_45915,N_43704,N_41334);
and U45916 (N_45916,N_40327,N_42598);
xor U45917 (N_45917,N_41928,N_40793);
xnor U45918 (N_45918,N_42845,N_43729);
nand U45919 (N_45919,N_40299,N_42985);
nor U45920 (N_45920,N_44517,N_41653);
and U45921 (N_45921,N_40609,N_43187);
or U45922 (N_45922,N_43111,N_43088);
or U45923 (N_45923,N_40859,N_43132);
nand U45924 (N_45924,N_41238,N_42358);
xnor U45925 (N_45925,N_43885,N_41569);
nand U45926 (N_45926,N_44165,N_42232);
or U45927 (N_45927,N_44931,N_40083);
nor U45928 (N_45928,N_43811,N_42322);
and U45929 (N_45929,N_43726,N_42149);
nor U45930 (N_45930,N_44804,N_40439);
xnor U45931 (N_45931,N_42746,N_42400);
or U45932 (N_45932,N_44801,N_42947);
xor U45933 (N_45933,N_42925,N_42062);
and U45934 (N_45934,N_42640,N_41194);
nor U45935 (N_45935,N_42968,N_44796);
xor U45936 (N_45936,N_40600,N_41467);
nor U45937 (N_45937,N_44924,N_41223);
or U45938 (N_45938,N_40283,N_42478);
nand U45939 (N_45939,N_43181,N_41048);
nor U45940 (N_45940,N_40788,N_40654);
xnor U45941 (N_45941,N_42444,N_42124);
or U45942 (N_45942,N_44508,N_41567);
nor U45943 (N_45943,N_40746,N_41582);
nand U45944 (N_45944,N_41627,N_42922);
or U45945 (N_45945,N_40703,N_42956);
nor U45946 (N_45946,N_40259,N_43917);
and U45947 (N_45947,N_44189,N_42180);
or U45948 (N_45948,N_42546,N_42001);
nor U45949 (N_45949,N_40322,N_42570);
and U45950 (N_45950,N_43128,N_40191);
nor U45951 (N_45951,N_43502,N_40588);
xor U45952 (N_45952,N_41333,N_42648);
or U45953 (N_45953,N_44385,N_43008);
nand U45954 (N_45954,N_44210,N_44775);
and U45955 (N_45955,N_44925,N_42161);
nor U45956 (N_45956,N_41392,N_44255);
and U45957 (N_45957,N_40233,N_44693);
nor U45958 (N_45958,N_40569,N_41937);
xor U45959 (N_45959,N_41641,N_44539);
nand U45960 (N_45960,N_40208,N_43773);
and U45961 (N_45961,N_41134,N_40596);
nand U45962 (N_45962,N_40757,N_40739);
nand U45963 (N_45963,N_43820,N_44600);
or U45964 (N_45964,N_40104,N_41892);
xnor U45965 (N_45965,N_43962,N_44259);
nor U45966 (N_45966,N_43602,N_42970);
and U45967 (N_45967,N_40994,N_40576);
or U45968 (N_45968,N_44395,N_40714);
nor U45969 (N_45969,N_42668,N_40656);
and U45970 (N_45970,N_41184,N_42681);
or U45971 (N_45971,N_42139,N_42497);
nor U45972 (N_45972,N_44829,N_43000);
xor U45973 (N_45973,N_44401,N_44461);
nand U45974 (N_45974,N_42295,N_44088);
nor U45975 (N_45975,N_40857,N_40974);
nand U45976 (N_45976,N_43010,N_44184);
nand U45977 (N_45977,N_44537,N_44311);
nand U45978 (N_45978,N_44043,N_43263);
xnor U45979 (N_45979,N_41997,N_44055);
nand U45980 (N_45980,N_40963,N_43842);
and U45981 (N_45981,N_40791,N_43072);
nor U45982 (N_45982,N_41414,N_40911);
nor U45983 (N_45983,N_43483,N_44613);
and U45984 (N_45984,N_41837,N_43036);
nand U45985 (N_45985,N_43781,N_41318);
nor U45986 (N_45986,N_43214,N_44079);
nand U45987 (N_45987,N_44817,N_41205);
and U45988 (N_45988,N_42392,N_43791);
and U45989 (N_45989,N_44007,N_40983);
nand U45990 (N_45990,N_44601,N_40676);
or U45991 (N_45991,N_40906,N_40408);
xor U45992 (N_45992,N_43892,N_41076);
nor U45993 (N_45993,N_43621,N_42263);
or U45994 (N_45994,N_41591,N_42287);
or U45995 (N_45995,N_43545,N_43937);
xor U45996 (N_45996,N_40177,N_43170);
nor U45997 (N_45997,N_43632,N_44937);
and U45998 (N_45998,N_43858,N_40143);
xor U45999 (N_45999,N_44273,N_44560);
or U46000 (N_46000,N_42000,N_43618);
nand U46001 (N_46001,N_44815,N_42744);
or U46002 (N_46002,N_43323,N_40749);
nor U46003 (N_46003,N_40650,N_42184);
nand U46004 (N_46004,N_42169,N_44159);
nor U46005 (N_46005,N_44366,N_40646);
nor U46006 (N_46006,N_43563,N_43366);
nand U46007 (N_46007,N_44893,N_43020);
or U46008 (N_46008,N_40261,N_44410);
nand U46009 (N_46009,N_43821,N_44386);
nor U46010 (N_46010,N_43344,N_40622);
nor U46011 (N_46011,N_44135,N_43762);
nand U46012 (N_46012,N_43786,N_41087);
or U46013 (N_46013,N_42935,N_41292);
and U46014 (N_46014,N_43243,N_43100);
nor U46015 (N_46015,N_42157,N_43720);
and U46016 (N_46016,N_40921,N_43687);
or U46017 (N_46017,N_44904,N_41640);
and U46018 (N_46018,N_41147,N_42403);
xnor U46019 (N_46019,N_44023,N_44025);
and U46020 (N_46020,N_40235,N_40432);
nand U46021 (N_46021,N_43905,N_41877);
and U46022 (N_46022,N_41630,N_44118);
and U46023 (N_46023,N_43950,N_42866);
or U46024 (N_46024,N_40616,N_40984);
xor U46025 (N_46025,N_41656,N_43659);
or U46026 (N_46026,N_42521,N_40288);
xor U46027 (N_46027,N_40805,N_42854);
nand U46028 (N_46028,N_43157,N_41994);
or U46029 (N_46029,N_44735,N_43435);
nor U46030 (N_46030,N_44640,N_42414);
and U46031 (N_46031,N_44014,N_40665);
xor U46032 (N_46032,N_41682,N_41116);
or U46033 (N_46033,N_42427,N_44922);
xor U46034 (N_46034,N_44992,N_41629);
nand U46035 (N_46035,N_42020,N_43348);
and U46036 (N_46036,N_41283,N_43027);
nor U46037 (N_46037,N_44680,N_43982);
nand U46038 (N_46038,N_44670,N_40781);
nand U46039 (N_46039,N_40985,N_42236);
or U46040 (N_46040,N_43780,N_43972);
xor U46041 (N_46041,N_43808,N_42335);
and U46042 (N_46042,N_43454,N_40833);
nand U46043 (N_46043,N_40381,N_42502);
nand U46044 (N_46044,N_41616,N_43911);
and U46045 (N_46045,N_42451,N_40742);
xor U46046 (N_46046,N_44761,N_44907);
nand U46047 (N_46047,N_42366,N_40564);
and U46048 (N_46048,N_43175,N_41484);
xnor U46049 (N_46049,N_40611,N_41010);
and U46050 (N_46050,N_41083,N_43198);
nand U46051 (N_46051,N_40939,N_40503);
and U46052 (N_46052,N_44520,N_42901);
and U46053 (N_46053,N_41120,N_44452);
and U46054 (N_46054,N_40706,N_41126);
xor U46055 (N_46055,N_42102,N_41672);
and U46056 (N_46056,N_42255,N_41498);
or U46057 (N_46057,N_40487,N_41290);
nand U46058 (N_46058,N_41993,N_40348);
xnor U46059 (N_46059,N_41038,N_44514);
nor U46060 (N_46060,N_44423,N_42841);
and U46061 (N_46061,N_40022,N_43159);
nand U46062 (N_46062,N_44644,N_43747);
or U46063 (N_46063,N_40404,N_42266);
or U46064 (N_46064,N_42630,N_43795);
nor U46065 (N_46065,N_41910,N_44227);
nand U46066 (N_46066,N_40826,N_40745);
or U46067 (N_46067,N_43524,N_43532);
xor U46068 (N_46068,N_44563,N_43288);
nor U46069 (N_46069,N_44836,N_43777);
and U46070 (N_46070,N_43397,N_43658);
xnor U46071 (N_46071,N_41739,N_42436);
nor U46072 (N_46072,N_42943,N_40485);
nor U46073 (N_46073,N_41186,N_41032);
or U46074 (N_46074,N_42499,N_42544);
or U46075 (N_46075,N_42483,N_40599);
nand U46076 (N_46076,N_40039,N_43287);
xor U46077 (N_46077,N_42986,N_41552);
nor U46078 (N_46078,N_42757,N_42593);
and U46079 (N_46079,N_40088,N_43357);
and U46080 (N_46080,N_43503,N_43713);
nor U46081 (N_46081,N_44472,N_42461);
nor U46082 (N_46082,N_40537,N_41115);
nor U46083 (N_46083,N_43614,N_40500);
nor U46084 (N_46084,N_42047,N_43184);
and U46085 (N_46085,N_43365,N_41024);
xor U46086 (N_46086,N_42969,N_41370);
nor U46087 (N_46087,N_42613,N_42019);
xnor U46088 (N_46088,N_40726,N_43549);
or U46089 (N_46089,N_42118,N_41141);
nand U46090 (N_46090,N_41256,N_43899);
xnor U46091 (N_46091,N_43706,N_43131);
or U46092 (N_46092,N_44041,N_42173);
nand U46093 (N_46093,N_40940,N_44756);
nor U46094 (N_46094,N_41733,N_42705);
or U46095 (N_46095,N_44606,N_43909);
xnor U46096 (N_46096,N_44374,N_42420);
nand U46097 (N_46097,N_40513,N_40909);
or U46098 (N_46098,N_43071,N_41055);
nor U46099 (N_46099,N_42904,N_43074);
nand U46100 (N_46100,N_43468,N_42440);
and U46101 (N_46101,N_41681,N_40105);
xnor U46102 (N_46102,N_42727,N_43738);
nor U46103 (N_46103,N_41764,N_42380);
and U46104 (N_46104,N_40278,N_41979);
or U46105 (N_46105,N_41081,N_42930);
nand U46106 (N_46106,N_41487,N_40477);
nand U46107 (N_46107,N_40975,N_40263);
or U46108 (N_46108,N_43608,N_43389);
xnor U46109 (N_46109,N_44930,N_44714);
nand U46110 (N_46110,N_41712,N_44662);
nor U46111 (N_46111,N_40825,N_41796);
and U46112 (N_46112,N_44426,N_44617);
nor U46113 (N_46113,N_41956,N_43431);
nor U46114 (N_46114,N_41619,N_41153);
nor U46115 (N_46115,N_41639,N_44224);
xor U46116 (N_46116,N_41625,N_42449);
nand U46117 (N_46117,N_42768,N_40890);
or U46118 (N_46118,N_41331,N_41178);
or U46119 (N_46119,N_43499,N_41468);
and U46120 (N_46120,N_44215,N_44681);
or U46121 (N_46121,N_43146,N_40751);
xnor U46122 (N_46122,N_42445,N_40563);
nand U46123 (N_46123,N_41862,N_44167);
nor U46124 (N_46124,N_40809,N_41383);
nand U46125 (N_46125,N_41372,N_43952);
or U46126 (N_46126,N_41933,N_41465);
or U46127 (N_46127,N_43924,N_41199);
or U46128 (N_46128,N_41349,N_42687);
nand U46129 (N_46129,N_43110,N_44516);
nand U46130 (N_46130,N_43526,N_44763);
xor U46131 (N_46131,N_41078,N_40908);
nor U46132 (N_46132,N_41872,N_44356);
xor U46133 (N_46133,N_43031,N_42931);
xnor U46134 (N_46134,N_41053,N_40700);
nand U46135 (N_46135,N_40359,N_42611);
nor U46136 (N_46136,N_44045,N_42535);
and U46137 (N_46137,N_43248,N_43790);
nor U46138 (N_46138,N_41802,N_41158);
nand U46139 (N_46139,N_40570,N_43934);
nand U46140 (N_46140,N_41462,N_42911);
nand U46141 (N_46141,N_43299,N_43203);
and U46142 (N_46142,N_42737,N_44561);
or U46143 (N_46143,N_41203,N_42220);
nor U46144 (N_46144,N_42472,N_42077);
nor U46145 (N_46145,N_40029,N_43147);
or U46146 (N_46146,N_43007,N_43054);
or U46147 (N_46147,N_42649,N_44657);
and U46148 (N_46148,N_41808,N_44554);
or U46149 (N_46149,N_40761,N_43834);
nor U46150 (N_46150,N_41486,N_44326);
nor U46151 (N_46151,N_44067,N_41731);
and U46152 (N_46152,N_40384,N_40981);
and U46153 (N_46153,N_44588,N_41129);
xor U46154 (N_46154,N_41504,N_40351);
or U46155 (N_46155,N_42830,N_42799);
xor U46156 (N_46156,N_43900,N_41941);
and U46157 (N_46157,N_44935,N_42878);
and U46158 (N_46158,N_42013,N_41940);
xor U46159 (N_46159,N_40484,N_41307);
or U46160 (N_46160,N_44251,N_44806);
or U46161 (N_46161,N_44257,N_41972);
and U46162 (N_46162,N_43303,N_41669);
or U46163 (N_46163,N_43716,N_44498);
and U46164 (N_46164,N_44439,N_41089);
and U46165 (N_46165,N_41298,N_43152);
and U46166 (N_46166,N_42508,N_40284);
nand U46167 (N_46167,N_44705,N_44777);
nand U46168 (N_46168,N_44830,N_41341);
nor U46169 (N_46169,N_41611,N_43154);
xnor U46170 (N_46170,N_43289,N_42104);
xnor U46171 (N_46171,N_43392,N_41230);
nor U46172 (N_46172,N_42107,N_42827);
nand U46173 (N_46173,N_41381,N_43598);
nand U46174 (N_46174,N_43321,N_42179);
xnor U46175 (N_46175,N_41581,N_41191);
and U46176 (N_46176,N_42709,N_41850);
nand U46177 (N_46177,N_44666,N_43040);
and U46178 (N_46178,N_44122,N_40615);
or U46179 (N_46179,N_43498,N_40942);
and U46180 (N_46180,N_44265,N_42015);
and U46181 (N_46181,N_43383,N_44651);
nand U46182 (N_46182,N_42686,N_41700);
or U46183 (N_46183,N_44918,N_40731);
or U46184 (N_46184,N_42740,N_40402);
xnor U46185 (N_46185,N_44867,N_40643);
nand U46186 (N_46186,N_43260,N_43093);
xnor U46187 (N_46187,N_41182,N_40773);
nand U46188 (N_46188,N_40428,N_41740);
nand U46189 (N_46189,N_40005,N_40112);
nand U46190 (N_46190,N_43064,N_40096);
nand U46191 (N_46191,N_44212,N_41618);
and U46192 (N_46192,N_41028,N_43994);
nand U46193 (N_46193,N_42365,N_40017);
nor U46194 (N_46194,N_41437,N_40491);
and U46195 (N_46195,N_43417,N_40822);
and U46196 (N_46196,N_44455,N_42916);
nand U46197 (N_46197,N_41857,N_40193);
and U46198 (N_46198,N_43601,N_43557);
nor U46199 (N_46199,N_43359,N_43974);
nor U46200 (N_46200,N_40575,N_42659);
or U46201 (N_46201,N_43630,N_42846);
nand U46202 (N_46202,N_40124,N_44630);
xor U46203 (N_46203,N_42028,N_40237);
nand U46204 (N_46204,N_41894,N_42202);
and U46205 (N_46205,N_42187,N_43835);
nand U46206 (N_46206,N_40168,N_43683);
xor U46207 (N_46207,N_40212,N_42183);
xnor U46208 (N_46208,N_44185,N_44868);
nand U46209 (N_46209,N_40031,N_41882);
nand U46210 (N_46210,N_42820,N_43919);
nor U46211 (N_46211,N_42114,N_44083);
xnor U46212 (N_46212,N_42541,N_40810);
nand U46213 (N_46213,N_41854,N_44008);
and U46214 (N_46214,N_43433,N_42700);
nor U46215 (N_46215,N_44131,N_43428);
or U46216 (N_46216,N_43645,N_40915);
or U46217 (N_46217,N_40853,N_44755);
xor U46218 (N_46218,N_42023,N_41824);
or U46219 (N_46219,N_41816,N_42690);
or U46220 (N_46220,N_44393,N_42831);
nand U46221 (N_46221,N_41634,N_40047);
and U46222 (N_46222,N_41408,N_43164);
or U46223 (N_46223,N_44684,N_41748);
or U46224 (N_46224,N_41328,N_40499);
and U46225 (N_46225,N_41875,N_42262);
xnor U46226 (N_46226,N_44582,N_43378);
nor U46227 (N_46227,N_44373,N_42567);
nor U46228 (N_46228,N_40677,N_43861);
nand U46229 (N_46229,N_44102,N_42606);
nand U46230 (N_46230,N_42378,N_41897);
nor U46231 (N_46231,N_42784,N_41168);
and U46232 (N_46232,N_44865,N_43329);
or U46233 (N_46233,N_44482,N_44198);
nor U46234 (N_46234,N_44031,N_43942);
and U46235 (N_46235,N_43592,N_41927);
xor U46236 (N_46236,N_42098,N_40347);
nand U46237 (N_46237,N_42377,N_40923);
nor U46238 (N_46238,N_41945,N_41526);
or U46239 (N_46239,N_42089,N_44834);
and U46240 (N_46240,N_40834,N_43477);
xnor U46241 (N_46241,N_42379,N_44142);
nor U46242 (N_46242,N_44545,N_41754);
and U46243 (N_46243,N_42993,N_42635);
xnor U46244 (N_46244,N_41890,N_42078);
or U46245 (N_46245,N_42045,N_40639);
xnor U46246 (N_46246,N_41538,N_43186);
or U46247 (N_46247,N_44547,N_40438);
nand U46248 (N_46248,N_43746,N_41117);
xor U46249 (N_46249,N_40971,N_43317);
xor U46250 (N_46250,N_41418,N_44282);
nor U46251 (N_46251,N_41805,N_41784);
xor U46252 (N_46252,N_43987,N_41420);
xor U46253 (N_46253,N_43024,N_42081);
or U46254 (N_46254,N_40156,N_40584);
and U46255 (N_46255,N_42945,N_42022);
nand U46256 (N_46256,N_41469,N_40551);
xnor U46257 (N_46257,N_40951,N_44243);
and U46258 (N_46258,N_40098,N_44541);
nand U46259 (N_46259,N_42337,N_40081);
and U46260 (N_46260,N_40068,N_44940);
or U46261 (N_46261,N_41589,N_41221);
nor U46262 (N_46262,N_40991,N_42405);
xor U46263 (N_46263,N_44375,N_44351);
nor U46264 (N_46264,N_43803,N_43951);
xnor U46265 (N_46265,N_44979,N_43719);
nor U46266 (N_46266,N_40242,N_40804);
and U46267 (N_46267,N_42620,N_41351);
and U46268 (N_46268,N_41470,N_40699);
nor U46269 (N_46269,N_44722,N_40134);
nand U46270 (N_46270,N_41086,N_40962);
or U46271 (N_46271,N_40888,N_41548);
xor U46272 (N_46272,N_42519,N_41935);
xnor U46273 (N_46273,N_40204,N_40733);
or U46274 (N_46274,N_42538,N_44576);
nor U46275 (N_46275,N_44971,N_41104);
xor U46276 (N_46276,N_43257,N_42320);
nor U46277 (N_46277,N_40062,N_44839);
or U46278 (N_46278,N_44013,N_43749);
or U46279 (N_46279,N_40230,N_44826);
nand U46280 (N_46280,N_44888,N_42317);
and U46281 (N_46281,N_40462,N_41195);
nor U46282 (N_46282,N_41572,N_44538);
and U46283 (N_46283,N_41019,N_40290);
nor U46284 (N_46284,N_42018,N_42683);
xor U46285 (N_46285,N_40741,N_42539);
and U46286 (N_46286,N_44316,N_40582);
and U46287 (N_46287,N_44266,N_40720);
xnor U46288 (N_46288,N_44525,N_40685);
xor U46289 (N_46289,N_43331,N_40966);
nor U46290 (N_46290,N_42695,N_40638);
or U46291 (N_46291,N_42504,N_44475);
xnor U46292 (N_46292,N_40848,N_43568);
xor U46293 (N_46293,N_41725,N_42840);
or U46294 (N_46294,N_41346,N_42435);
and U46295 (N_46295,N_40787,N_40907);
nand U46296 (N_46296,N_42272,N_43794);
nor U46297 (N_46297,N_44821,N_40712);
and U46298 (N_46298,N_43272,N_40972);
nor U46299 (N_46299,N_43224,N_41150);
and U46300 (N_46300,N_43264,N_40444);
xnor U46301 (N_46301,N_43800,N_44689);
or U46302 (N_46302,N_43988,N_41730);
nor U46303 (N_46303,N_42165,N_42097);
xnor U46304 (N_46304,N_41269,N_42125);
nand U46305 (N_46305,N_43494,N_42106);
and U46306 (N_46306,N_43025,N_42021);
nor U46307 (N_46307,N_41045,N_44927);
xnor U46308 (N_46308,N_42776,N_43691);
nand U46309 (N_46309,N_40818,N_41705);
and U46310 (N_46310,N_44695,N_40176);
nor U46311 (N_46311,N_42227,N_44773);
nand U46312 (N_46312,N_40783,N_41358);
xor U46313 (N_46313,N_41319,N_40889);
and U46314 (N_46314,N_44976,N_41343);
or U46315 (N_46315,N_43161,N_43090);
nor U46316 (N_46316,N_43182,N_42816);
and U46317 (N_46317,N_41390,N_42188);
xor U46318 (N_46318,N_43735,N_42576);
nor U46319 (N_46319,N_43824,N_44239);
and U46320 (N_46320,N_44993,N_42920);
and U46321 (N_46321,N_41303,N_41626);
or U46322 (N_46322,N_42293,N_43852);
nor U46323 (N_46323,N_43377,N_44683);
nand U46324 (N_46324,N_42503,N_41913);
xor U46325 (N_46325,N_42068,N_41732);
and U46326 (N_46326,N_42298,N_41939);
nor U46327 (N_46327,N_43497,N_40937);
nand U46328 (N_46328,N_40271,N_40130);
and U46329 (N_46329,N_44402,N_43495);
or U46330 (N_46330,N_42279,N_43060);
nor U46331 (N_46331,N_43740,N_41881);
nor U46332 (N_46332,N_41959,N_42364);
xor U46333 (N_46333,N_40724,N_43352);
xnor U46334 (N_46334,N_44858,N_44062);
nor U46335 (N_46335,N_42698,N_42101);
xor U46336 (N_46336,N_41171,N_43067);
nor U46337 (N_46337,N_41842,N_44308);
nand U46338 (N_46338,N_44264,N_43769);
nand U46339 (N_46339,N_40861,N_43059);
and U46340 (N_46340,N_40358,N_44949);
nand U46341 (N_46341,N_44460,N_42460);
nor U46342 (N_46342,N_43043,N_44880);
or U46343 (N_46343,N_44823,N_44029);
nand U46344 (N_46344,N_44837,N_44783);
and U46345 (N_46345,N_40457,N_43475);
nand U46346 (N_46346,N_41407,N_43176);
xnor U46347 (N_46347,N_42869,N_40542);
nand U46348 (N_46348,N_44136,N_40957);
nand U46349 (N_46349,N_44903,N_44054);
nor U46350 (N_46350,N_40581,N_42650);
nor U46351 (N_46351,N_43627,N_42140);
nand U46352 (N_46352,N_42221,N_43249);
xnor U46353 (N_46353,N_42486,N_42585);
or U46354 (N_46354,N_41338,N_41403);
and U46355 (N_46355,N_41399,N_41988);
or U46356 (N_46356,N_43244,N_44047);
nor U46357 (N_46357,N_43809,N_42838);
xnor U46358 (N_46358,N_41376,N_43628);
nor U46359 (N_46359,N_42433,N_42357);
nor U46360 (N_46360,N_43696,N_44256);
nand U46361 (N_46361,N_42761,N_40158);
or U46362 (N_46362,N_40494,N_44180);
xor U46363 (N_46363,N_43859,N_41771);
xor U46364 (N_46364,N_41183,N_42758);
or U46365 (N_46365,N_44219,N_41529);
nand U46366 (N_46366,N_43724,N_41459);
xor U46367 (N_46367,N_40649,N_44474);
and U46368 (N_46368,N_40466,N_43106);
xnor U46369 (N_46369,N_43254,N_40125);
nor U46370 (N_46370,N_40566,N_42712);
or U46371 (N_46371,N_40181,N_41885);
xor U46372 (N_46372,N_40965,N_40452);
and U46373 (N_46373,N_42513,N_43490);
nor U46374 (N_46374,N_40340,N_41219);
or U46375 (N_46375,N_40816,N_42373);
nand U46376 (N_46376,N_44851,N_42398);
and U46377 (N_46377,N_41674,N_44042);
or U46378 (N_46378,N_42201,N_44132);
nor U46379 (N_46379,N_44849,N_41852);
or U46380 (N_46380,N_42876,N_40238);
nor U46381 (N_46381,N_44129,N_43714);
nand U46382 (N_46382,N_40175,N_44305);
and U46383 (N_46383,N_41294,N_40470);
nand U46384 (N_46384,N_44598,N_44112);
and U46385 (N_46385,N_43250,N_42657);
and U46386 (N_46386,N_42093,N_41464);
or U46387 (N_46387,N_40341,N_44813);
or U46388 (N_46388,N_41226,N_40970);
nand U46389 (N_46389,N_43849,N_42248);
nor U46390 (N_46390,N_44913,N_40274);
xor U46391 (N_46391,N_43258,N_42796);
nor U46392 (N_46392,N_41192,N_41339);
nor U46393 (N_46393,N_41721,N_40976);
or U46394 (N_46394,N_43162,N_40682);
xnor U46395 (N_46395,N_44447,N_42153);
or U46396 (N_46396,N_43869,N_42250);
nor U46397 (N_46397,N_44828,N_41501);
nor U46398 (N_46398,N_44616,N_44564);
xor U46399 (N_46399,N_43364,N_42862);
and U46400 (N_46400,N_41925,N_43647);
and U46401 (N_46401,N_40385,N_43350);
xor U46402 (N_46402,N_42950,N_41943);
nor U46403 (N_46403,N_41510,N_40996);
or U46404 (N_46404,N_41609,N_41140);
xor U46405 (N_46405,N_42048,N_41650);
nor U46406 (N_46406,N_41316,N_44009);
and U46407 (N_46407,N_44442,N_44050);
nand U46408 (N_46408,N_42284,N_40501);
nor U46409 (N_46409,N_44217,N_43868);
nor U46410 (N_46410,N_41962,N_42299);
xor U46411 (N_46411,N_40567,N_41131);
or U46412 (N_46412,N_42817,N_41508);
nand U46413 (N_46413,N_42810,N_40184);
xor U46414 (N_46414,N_40752,N_43985);
nand U46415 (N_46415,N_42123,N_41367);
nor U46416 (N_46416,N_42421,N_41034);
or U46417 (N_46417,N_42981,N_44842);
xnor U46418 (N_46418,N_44477,N_41807);
nand U46419 (N_46419,N_41013,N_44090);
or U46420 (N_46420,N_41540,N_44519);
and U46421 (N_46421,N_41996,N_43282);
nor U46422 (N_46422,N_41596,N_41234);
xor U46423 (N_46423,N_40482,N_44603);
and U46424 (N_46424,N_43009,N_42615);
xor U46425 (N_46425,N_42517,N_41779);
xnor U46426 (N_46426,N_43625,N_40593);
nand U46427 (N_46427,N_41007,N_43279);
and U46428 (N_46428,N_44068,N_44762);
and U46429 (N_46429,N_44629,N_41947);
or U46430 (N_46430,N_41154,N_41886);
or U46431 (N_46431,N_42735,N_42506);
and U46432 (N_46432,N_42984,N_44409);
and U46433 (N_46433,N_40300,N_42006);
nor U46434 (N_46434,N_44709,N_41330);
nand U46435 (N_46435,N_44805,N_41047);
and U46436 (N_46436,N_42456,N_41859);
nor U46437 (N_46437,N_42834,N_40307);
or U46438 (N_46438,N_40160,N_43371);
and U46439 (N_46439,N_42554,N_44618);
and U46440 (N_46440,N_40896,N_44241);
xnor U46441 (N_46441,N_44003,N_41654);
nor U46442 (N_46442,N_40871,N_44010);
and U46443 (N_46443,N_42565,N_42871);
or U46444 (N_46444,N_43722,N_44454);
xnor U46445 (N_46445,N_44962,N_43297);
or U46446 (N_46446,N_42765,N_44846);
xnor U46447 (N_46447,N_41432,N_44200);
nand U46448 (N_46448,N_42515,N_42982);
nor U46449 (N_46449,N_43044,N_44446);
xor U46450 (N_46450,N_40164,N_41746);
and U46451 (N_46451,N_44648,N_41124);
or U46452 (N_46452,N_42614,N_41110);
nand U46453 (N_46453,N_43607,N_42099);
and U46454 (N_46454,N_41655,N_42671);
xor U46455 (N_46455,N_42086,N_42632);
nand U46456 (N_46456,N_40328,N_44404);
and U46457 (N_46457,N_41573,N_42706);
or U46458 (N_46458,N_44070,N_43765);
and U46459 (N_46459,N_40549,N_43449);
and U46460 (N_46460,N_42989,N_44063);
and U46461 (N_46461,N_42474,N_42056);
and U46462 (N_46462,N_44579,N_40417);
and U46463 (N_46463,N_44077,N_40216);
and U46464 (N_46464,N_40673,N_42749);
or U46465 (N_46465,N_42928,N_43664);
nand U46466 (N_46466,N_42753,N_44258);
or U46467 (N_46467,N_44864,N_44619);
nand U46468 (N_46468,N_41382,N_44869);
xnor U46469 (N_46469,N_43207,N_42463);
and U46470 (N_46470,N_42470,N_44713);
and U46471 (N_46471,N_42243,N_41043);
xnor U46472 (N_46472,N_43662,N_42204);
or U46473 (N_46473,N_41977,N_44984);
or U46474 (N_46474,N_41473,N_42465);
or U46475 (N_46475,N_43547,N_43804);
xnor U46476 (N_46476,N_40692,N_43079);
and U46477 (N_46477,N_43575,N_40058);
xor U46478 (N_46478,N_41679,N_41590);
and U46479 (N_46479,N_43429,N_43261);
nand U46480 (N_46480,N_43887,N_43591);
nand U46481 (N_46481,N_44325,N_41622);
and U46482 (N_46482,N_42848,N_44852);
or U46483 (N_46483,N_40231,N_44387);
xnor U46484 (N_46484,N_43778,N_44004);
xnor U46485 (N_46485,N_44179,N_41745);
or U46486 (N_46486,N_42730,N_43505);
nand U46487 (N_46487,N_41766,N_42024);
and U46488 (N_46488,N_43033,N_43097);
xnor U46489 (N_46489,N_44758,N_43586);
nor U46490 (N_46490,N_42409,N_42537);
or U46491 (N_46491,N_43451,N_40986);
xor U46492 (N_46492,N_40101,N_43880);
nand U46493 (N_46493,N_42058,N_42244);
nand U46494 (N_46494,N_41077,N_40508);
or U46495 (N_46495,N_40295,N_43521);
nor U46496 (N_46496,N_41967,N_44361);
or U46497 (N_46497,N_43836,N_42755);
or U46498 (N_46498,N_43327,N_42304);
nand U46499 (N_46499,N_44819,N_44277);
nand U46500 (N_46500,N_40943,N_44863);
nand U46501 (N_46501,N_42371,N_40269);
and U46502 (N_46502,N_43346,N_44747);
nor U46503 (N_46503,N_44056,N_40287);
nor U46504 (N_46504,N_40653,N_41164);
nand U46505 (N_46505,N_44363,N_40497);
and U46506 (N_46506,N_42797,N_40048);
or U46507 (N_46507,N_44584,N_40708);
and U46508 (N_46508,N_44248,N_42222);
nor U46509 (N_46509,N_43964,N_40110);
nand U46510 (N_46510,N_41663,N_42723);
or U46511 (N_46511,N_42063,N_41878);
nor U46512 (N_46512,N_44779,N_41478);
nand U46513 (N_46513,N_42203,N_42954);
xor U46514 (N_46514,N_43005,N_41602);
nand U46515 (N_46515,N_40806,N_40950);
or U46516 (N_46516,N_42413,N_41097);
or U46517 (N_46517,N_41578,N_42626);
or U46518 (N_46518,N_44418,N_42766);
xor U46519 (N_46519,N_43774,N_41384);
and U46520 (N_46520,N_43446,N_40419);
xnor U46521 (N_46521,N_41916,N_44782);
nand U46522 (N_46522,N_41159,N_40901);
nor U46523 (N_46523,N_42912,N_42891);
nand U46524 (N_46524,N_44704,N_42828);
xnor U46525 (N_46525,N_41827,N_41133);
and U46526 (N_46526,N_40412,N_43677);
or U46527 (N_46527,N_40489,N_42441);
xnor U46528 (N_46528,N_41278,N_40225);
and U46529 (N_46529,N_41758,N_44391);
nand U46530 (N_46530,N_41266,N_44674);
or U46531 (N_46531,N_44417,N_40759);
and U46532 (N_46532,N_42313,N_44245);
and U46533 (N_46533,N_41252,N_40586);
or U46534 (N_46534,N_43509,N_44637);
nand U46535 (N_46535,N_40226,N_44752);
or U46536 (N_46536,N_41612,N_41441);
nor U46537 (N_46537,N_44174,N_44934);
or U46538 (N_46538,N_41728,N_40660);
or U46539 (N_46539,N_40142,N_41911);
xor U46540 (N_46540,N_43940,N_40463);
or U46541 (N_46541,N_41145,N_43676);
xor U46542 (N_46542,N_41891,N_43634);
nand U46543 (N_46543,N_43993,N_42999);
or U46544 (N_46544,N_40640,N_40877);
nand U46545 (N_46545,N_44486,N_42105);
nor U46546 (N_46546,N_40900,N_41649);
or U46547 (N_46547,N_42774,N_44860);
nor U46548 (N_46548,N_42855,N_44527);
xnor U46549 (N_46549,N_42868,N_40538);
nand U46550 (N_46550,N_41306,N_44844);
nor U46551 (N_46551,N_42130,N_43205);
nor U46552 (N_46552,N_40543,N_40171);
nor U46553 (N_46553,N_43648,N_42940);
or U46554 (N_46554,N_42636,N_44565);
nand U46555 (N_46555,N_42623,N_43226);
nand U46556 (N_46556,N_41722,N_41250);
xor U46557 (N_46557,N_42756,N_44956);
and U46558 (N_46558,N_40858,N_42388);
nand U46559 (N_46559,N_42003,N_44075);
xor U46560 (N_46560,N_40764,N_41818);
nand U46561 (N_46561,N_44022,N_41828);
xor U46562 (N_46562,N_42092,N_40401);
nor U46563 (N_46563,N_43144,N_43761);
or U46564 (N_46564,N_44663,N_42564);
nor U46565 (N_46565,N_40628,N_41417);
xnor U46566 (N_46566,N_42359,N_43751);
or U46567 (N_46567,N_44458,N_43936);
nor U46568 (N_46568,N_40335,N_43963);
or U46569 (N_46569,N_40016,N_44770);
xor U46570 (N_46570,N_40594,N_43313);
or U46571 (N_46571,N_44405,N_42882);
and U46572 (N_46572,N_43301,N_41137);
nand U46573 (N_46573,N_41144,N_43493);
nor U46574 (N_46574,N_43422,N_44891);
nor U46575 (N_46575,N_44948,N_43337);
nor U46576 (N_46576,N_43961,N_44748);
nand U46577 (N_46577,N_43817,N_43463);
or U46578 (N_46578,N_44231,N_42547);
or U46579 (N_46579,N_44641,N_43736);
or U46580 (N_46580,N_43089,N_41522);
nor U46581 (N_46581,N_44745,N_41832);
and U46582 (N_46582,N_44459,N_42691);
nor U46583 (N_46583,N_41434,N_41646);
and U46584 (N_46584,N_41021,N_43520);
or U46585 (N_46585,N_40206,N_43818);
nand U46586 (N_46586,N_41539,N_41974);
xor U46587 (N_46587,N_41689,N_41900);
and U46588 (N_46588,N_40718,N_44727);
xor U46589 (N_46589,N_43361,N_44573);
or U46590 (N_46590,N_42355,N_40437);
or U46591 (N_46591,N_41163,N_41964);
nand U46592 (N_46592,N_44164,N_40684);
xor U46593 (N_46593,N_40849,N_43467);
nand U46594 (N_46594,N_41446,N_42344);
and U46595 (N_46595,N_43426,N_43649);
xnor U46596 (N_46596,N_44701,N_41064);
nor U46597 (N_46597,N_41896,N_41233);
nand U46598 (N_46598,N_41443,N_40678);
and U46599 (N_46599,N_43725,N_42770);
or U46600 (N_46600,N_44048,N_44044);
and U46601 (N_46601,N_40794,N_44970);
nor U46602 (N_46602,N_44728,N_42500);
or U46603 (N_46603,N_43351,N_42638);
and U46604 (N_46604,N_41401,N_41785);
and U46605 (N_46605,N_41917,N_44753);
and U46606 (N_46606,N_42713,N_44774);
nand U46607 (N_46607,N_41257,N_44315);
nand U46608 (N_46608,N_43129,N_43156);
nor U46609 (N_46609,N_42785,N_40138);
nor U46610 (N_46610,N_40188,N_42747);
and U46611 (N_46611,N_43529,N_41313);
and U46612 (N_46612,N_43234,N_41835);
and U46613 (N_46613,N_44848,N_44340);
nand U46614 (N_46614,N_42955,N_43456);
nand U46615 (N_46615,N_44424,N_41429);
nand U46616 (N_46616,N_41496,N_44543);
xor U46617 (N_46617,N_43709,N_42760);
and U46618 (N_46618,N_44463,N_43312);
or U46619 (N_46619,N_41874,N_41992);
xnor U46620 (N_46620,N_40478,N_42988);
nand U46621 (N_46621,N_44791,N_44113);
or U46622 (N_46622,N_41136,N_42610);
and U46623 (N_46623,N_42680,N_42457);
nor U46624 (N_46624,N_41050,N_42480);
or U46625 (N_46625,N_42899,N_40536);
nor U46626 (N_46626,N_44436,N_40342);
xnor U46627 (N_46627,N_41965,N_42034);
or U46628 (N_46628,N_40301,N_43460);
or U46629 (N_46629,N_43095,N_41574);
nand U46630 (N_46630,N_41870,N_41562);
or U46631 (N_46631,N_43037,N_44938);
nor U46632 (N_46632,N_44338,N_43006);
or U46633 (N_46633,N_44006,N_44585);
and U46634 (N_46634,N_42401,N_42523);
and U46635 (N_46635,N_43174,N_43855);
nand U46636 (N_46636,N_43544,N_41175);
and U46637 (N_46637,N_44272,N_40642);
xnor U46638 (N_46638,N_42628,N_42602);
nor U46639 (N_46639,N_40037,N_42274);
or U46640 (N_46640,N_44469,N_41774);
and U46641 (N_46641,N_44456,N_41820);
xor U46642 (N_46642,N_43896,N_44348);
and U46643 (N_46643,N_40956,N_41760);
and U46644 (N_46644,N_43879,N_43183);
or U46645 (N_46645,N_40762,N_42803);
nand U46646 (N_46646,N_41982,N_41272);
nor U46647 (N_46647,N_42356,N_43021);
xnor U46648 (N_46648,N_41904,N_42674);
xnor U46649 (N_46649,N_44018,N_41868);
and U46650 (N_46650,N_43191,N_42450);
nor U46651 (N_46651,N_40360,N_40155);
nand U46652 (N_46652,N_40558,N_43081);
nor U46653 (N_46653,N_44246,N_43473);
nor U46654 (N_46654,N_41321,N_42316);
xor U46655 (N_46655,N_41249,N_40658);
nand U46656 (N_46656,N_43889,N_40496);
and U46657 (N_46657,N_42583,N_42843);
nand U46658 (N_46658,N_43784,N_44555);
nor U46659 (N_46659,N_44647,N_41400);
or U46660 (N_46660,N_44832,N_40910);
nand U46661 (N_46661,N_42289,N_43760);
and U46662 (N_46662,N_41398,N_43513);
xor U46663 (N_46663,N_44943,N_40696);
and U46664 (N_46664,N_40121,N_40107);
xor U46665 (N_46665,N_43622,N_41322);
nand U46666 (N_46666,N_40891,N_42408);
nor U46667 (N_46667,N_41839,N_44320);
nand U46668 (N_46668,N_43875,N_44726);
or U46669 (N_46669,N_41621,N_41635);
nand U46670 (N_46670,N_40424,N_43137);
nand U46671 (N_46671,N_42242,N_40389);
xor U46672 (N_46672,N_40511,N_40814);
nor U46673 (N_46673,N_40292,N_42041);
nand U46674 (N_46674,N_43996,N_40932);
and U46675 (N_46675,N_41442,N_40434);
nor U46676 (N_46676,N_44069,N_40842);
xnor U46677 (N_46677,N_40103,N_41792);
and U46678 (N_46678,N_43978,N_42549);
nor U46679 (N_46679,N_44095,N_40122);
xnor U46680 (N_46680,N_44470,N_44952);
nand U46681 (N_46681,N_44319,N_40182);
xnor U46682 (N_46682,N_42268,N_40895);
xnor U46683 (N_46683,N_42423,N_44494);
nor U46684 (N_46684,N_44350,N_42601);
or U46685 (N_46685,N_40792,N_42164);
xnor U46686 (N_46686,N_43237,N_41362);
nand U46687 (N_46687,N_42692,N_40517);
or U46688 (N_46688,N_40471,N_43857);
or U46689 (N_46689,N_40129,N_44397);
nand U46690 (N_46690,N_42607,N_44345);
nor U46691 (N_46691,N_41983,N_43884);
nand U46692 (N_46692,N_41189,N_44365);
xnor U46693 (N_46693,N_44304,N_43667);
xor U46694 (N_46694,N_40210,N_42946);
nand U46695 (N_46695,N_41647,N_44632);
xor U46696 (N_46696,N_44594,N_44388);
and U46697 (N_46697,N_44425,N_43657);
nand U46698 (N_46698,N_42591,N_41190);
and U46699 (N_46699,N_44437,N_40416);
and U46700 (N_46700,N_42429,N_44480);
and U46701 (N_46701,N_42145,N_41380);
nand U46702 (N_46702,N_40458,N_40917);
and U46703 (N_46703,N_44134,N_42808);
or U46704 (N_46704,N_43851,N_41817);
and U46705 (N_46705,N_40927,N_41719);
and U46706 (N_46706,N_42580,N_44800);
nor U46707 (N_46707,N_43517,N_40595);
xnor U46708 (N_46708,N_44738,N_42669);
nor U46709 (N_46709,N_40415,N_44586);
xor U46710 (N_46710,N_40140,N_43085);
nand U46711 (N_46711,N_40410,N_43637);
xor U46712 (N_46712,N_43320,N_41410);
nand U46713 (N_46713,N_42532,N_42742);
or U46714 (N_46714,N_41887,N_41558);
and U46715 (N_46715,N_44602,N_40383);
and U46716 (N_46716,N_43308,N_43864);
nand U46717 (N_46717,N_41426,N_44072);
nand U46718 (N_46718,N_40250,N_42329);
and U46719 (N_46719,N_40734,N_44169);
or U46720 (N_46720,N_44359,N_42736);
nor U46721 (N_46721,N_43732,N_44772);
and U46722 (N_46722,N_40369,N_41222);
nand U46723 (N_46723,N_41821,N_44130);
nand U46724 (N_46724,N_40297,N_41553);
nor U46725 (N_46725,N_44968,N_40072);
xnor U46726 (N_46726,N_42171,N_40141);
nand U46727 (N_46727,N_43559,N_43061);
xor U46728 (N_46728,N_44500,N_44694);
or U46729 (N_46729,N_42417,N_40840);
nand U46730 (N_46730,N_42488,N_43533);
xor U46731 (N_46731,N_40922,N_42863);
or U46732 (N_46732,N_44919,N_44933);
xor U46733 (N_46733,N_40585,N_41201);
nor U46734 (N_46734,N_40371,N_42214);
nor U46735 (N_46735,N_42835,N_43265);
or U46736 (N_46736,N_41423,N_44336);
nand U46737 (N_46737,N_40431,N_43850);
xnor U46738 (N_46738,N_41427,N_43583);
and U46739 (N_46739,N_44803,N_41248);
nand U46740 (N_46740,N_44511,N_41922);
nor U46741 (N_46741,N_40276,N_42974);
nor U46742 (N_46742,N_43705,N_43998);
or U46743 (N_46743,N_42109,N_41556);
nand U46744 (N_46744,N_43504,N_41949);
nand U46745 (N_46745,N_40435,N_41762);
xor U46746 (N_46746,N_44367,N_41448);
nand U46747 (N_46747,N_41889,N_41830);
nand U46748 (N_46748,N_41826,N_40550);
and U46749 (N_46749,N_42987,N_41419);
nor U46750 (N_46750,N_40533,N_44552);
xnor U46751 (N_46751,N_43386,N_43772);
nand U46752 (N_46752,N_40846,N_43711);
xnor U46753 (N_46753,N_43641,N_44368);
nand U46754 (N_46754,N_44127,N_40801);
nor U46755 (N_46755,N_41299,N_44877);
and U46756 (N_46756,N_43539,N_42767);
and U46757 (N_46757,N_40247,N_40535);
nor U46758 (N_46758,N_40899,N_43552);
and U46759 (N_46759,N_43782,N_44510);
xnor U46760 (N_46760,N_42798,N_40945);
nand U46761 (N_46761,N_40272,N_41742);
xnor U46762 (N_46762,N_40159,N_40316);
and U46763 (N_46763,N_41905,N_41662);
or U46764 (N_46764,N_40197,N_44335);
nor U46765 (N_46765,N_43052,N_43652);
xnor U46766 (N_46766,N_41561,N_40069);
nor U46767 (N_46767,N_41743,N_43407);
or U46768 (N_46768,N_41698,N_42603);
xor U46769 (N_46769,N_41070,N_44290);
or U46770 (N_46770,N_41497,N_40774);
nor U46771 (N_46771,N_40737,N_42849);
or U46772 (N_46772,N_40099,N_43278);
and U46773 (N_46773,N_40607,N_44611);
nand U46774 (N_46774,N_44503,N_43845);
xnor U46775 (N_46775,N_40729,N_44197);
nor U46776 (N_46776,N_42661,N_42907);
nor U46777 (N_46777,N_42235,N_43514);
nor U46778 (N_46778,N_40118,N_43434);
xnor U46779 (N_46779,N_44688,N_41752);
or U46780 (N_46780,N_43983,N_41092);
xnor U46781 (N_46781,N_42166,N_43501);
or U46782 (N_46782,N_40178,N_43594);
xor U46783 (N_46783,N_42997,N_44639);
nand U46784 (N_46784,N_42447,N_42082);
nor U46785 (N_46785,N_41515,N_43410);
nand U46786 (N_46786,N_44746,N_44281);
or U46787 (N_46787,N_41113,N_40561);
or U46788 (N_46788,N_41579,N_43681);
xor U46789 (N_46789,N_41600,N_43326);
nand U46790 (N_46790,N_40876,N_43306);
nor U46791 (N_46791,N_41823,N_40087);
and U46792 (N_46792,N_42654,N_40887);
xor U46793 (N_46793,N_41282,N_41350);
or U46794 (N_46794,N_44605,N_44720);
and U46795 (N_46795,N_43255,N_42267);
xor U46796 (N_46796,N_44238,N_44111);
nand U46797 (N_46797,N_42113,N_41880);
xor U46798 (N_46798,N_43898,N_44916);
xor U46799 (N_46799,N_43731,N_41264);
xor U46800 (N_46800,N_44625,N_40449);
xor U46801 (N_46801,N_41637,N_42983);
or U46802 (N_46802,N_43121,N_42095);
or U46803 (N_46803,N_44818,N_42791);
and U46804 (N_46804,N_41096,N_42363);
xor U46805 (N_46805,N_40032,N_44492);
or U46806 (N_46806,N_42805,N_40090);
nor U46807 (N_46807,N_44574,N_43437);
nand U46808 (N_46808,N_44896,N_41518);
and U46809 (N_46809,N_43334,N_43188);
and U46810 (N_46810,N_41798,N_42182);
xor U46811 (N_46811,N_40249,N_41062);
xor U46812 (N_46812,N_40465,N_41174);
or U46813 (N_46813,N_44060,N_42618);
and U46814 (N_46814,N_43328,N_41851);
and U46815 (N_46815,N_42763,N_41394);
or U46816 (N_46816,N_40282,N_44263);
or U46817 (N_46817,N_42667,N_43402);
nand U46818 (N_46818,N_40314,N_44016);
nor U46819 (N_46819,N_41099,N_43775);
nand U46820 (N_46820,N_44967,N_44261);
and U46821 (N_46821,N_40223,N_43893);
nand U46822 (N_46822,N_40319,N_44531);
or U46823 (N_46823,N_43620,N_41605);
or U46824 (N_46824,N_42257,N_43755);
nor U46825 (N_46825,N_40440,N_40357);
nand U46826 (N_46826,N_44024,N_43480);
and U46827 (N_46827,N_43822,N_44626);
xnor U46828 (N_46828,N_43210,N_44381);
xor U46829 (N_46829,N_42384,N_44515);
and U46830 (N_46830,N_42200,N_40587);
or U46831 (N_46831,N_43399,N_41502);
and U46832 (N_46832,N_40162,N_41780);
or U46833 (N_46833,N_44274,N_40755);
or U46834 (N_46834,N_43220,N_41207);
xnor U46835 (N_46835,N_42493,N_41822);
and U46836 (N_46836,N_41385,N_44546);
and U46837 (N_46837,N_41735,N_42369);
xor U46838 (N_46838,N_40451,N_40748);
nor U46839 (N_46839,N_43562,N_43750);
or U46840 (N_46840,N_43995,N_42390);
xor U46841 (N_46841,N_43712,N_41946);
nand U46842 (N_46842,N_40553,N_42972);
and U46843 (N_46843,N_41025,N_42927);
nor U46844 (N_46844,N_41463,N_43212);
nor U46845 (N_46845,N_41738,N_41227);
xor U46846 (N_46846,N_41265,N_40034);
nor U46847 (N_46847,N_43654,N_41876);
nand U46848 (N_46848,N_42873,N_42238);
nor U46849 (N_46849,N_42117,N_44897);
nor U46850 (N_46850,N_41020,N_40136);
nand U46851 (N_46851,N_43379,N_40625);
nand U46852 (N_46852,N_43692,N_40727);
nor U46853 (N_46853,N_44697,N_42711);
and U46854 (N_46854,N_44744,N_43802);
or U46855 (N_46855,N_40598,N_41268);
nand U46856 (N_46856,N_41642,N_43042);
nand U46857 (N_46857,N_44064,N_41049);
and U46858 (N_46858,N_40548,N_43878);
nor U46859 (N_46859,N_42069,N_41901);
or U46860 (N_46860,N_41421,N_42886);
nor U46861 (N_46861,N_40881,N_41957);
and U46862 (N_46862,N_40935,N_40150);
nand U46863 (N_46863,N_41018,N_44496);
nand U46864 (N_46864,N_44872,N_42343);
nor U46865 (N_46865,N_40095,N_43541);
or U46866 (N_46866,N_41281,N_41688);
and U46867 (N_46867,N_44059,N_42720);
xnor U46868 (N_46868,N_43134,N_41871);
nor U46869 (N_46869,N_43001,N_41098);
or U46870 (N_46870,N_44457,N_43810);
and U46871 (N_46871,N_42410,N_44082);
nor U46872 (N_46872,N_43053,N_43492);
or U46873 (N_46873,N_41436,N_41016);
and U46874 (N_46874,N_43929,N_42631);
and U46875 (N_46875,N_43353,N_43977);
and U46876 (N_46876,N_41673,N_41861);
nor U46877 (N_46877,N_44444,N_41347);
or U46878 (N_46878,N_42196,N_40356);
xnor U46879 (N_46879,N_42948,N_41834);
and U46880 (N_46880,N_44301,N_41597);
nor U46881 (N_46881,N_43626,N_43482);
or U46882 (N_46882,N_40394,N_44807);
xor U46883 (N_46883,N_43058,N_44182);
or U46884 (N_46884,N_40694,N_42962);
nand U46885 (N_46885,N_44643,N_44785);
nand U46886 (N_46886,N_44435,N_44000);
or U46887 (N_46887,N_42485,N_41156);
or U46888 (N_46888,N_40055,N_43723);
nand U46889 (N_46889,N_41944,N_43954);
xnor U46890 (N_46890,N_41923,N_43700);
nand U46891 (N_46891,N_44614,N_43616);
and U46892 (N_46892,N_41536,N_43363);
and U46893 (N_46893,N_44947,N_41142);
and U46894 (N_46894,N_41665,N_41288);
nand U46895 (N_46895,N_44211,N_42647);
or U46896 (N_46896,N_41799,N_40253);
nor U46897 (N_46897,N_44242,N_43944);
nor U46898 (N_46898,N_44021,N_42209);
or U46899 (N_46899,N_40312,N_43865);
and U46900 (N_46900,N_44765,N_44306);
nor U46901 (N_46901,N_42368,N_43605);
and U46902 (N_46902,N_44767,N_41151);
or U46903 (N_46903,N_40418,N_41247);
nand U46904 (N_46904,N_40885,N_40330);
and U46905 (N_46905,N_40851,N_42701);
nand U46906 (N_46906,N_41285,N_43179);
nand U46907 (N_46907,N_43172,N_43604);
nand U46908 (N_46908,N_42452,N_40423);
and U46909 (N_46909,N_42434,N_42895);
nor U46910 (N_46910,N_44400,N_43866);
nor U46911 (N_46911,N_40978,N_42542);
or U46912 (N_46912,N_43019,N_43629);
xnor U46913 (N_46913,N_41973,N_41406);
xor U46914 (N_46914,N_44026,N_40020);
nor U46915 (N_46915,N_44216,N_42194);
nor U46916 (N_46916,N_43844,N_40281);
nand U46917 (N_46917,N_44443,N_41356);
and U46918 (N_46918,N_44502,N_44223);
and U46919 (N_46919,N_41082,N_43819);
nor U46920 (N_46920,N_40430,N_42933);
xnor U46921 (N_46921,N_41369,N_43792);
xor U46922 (N_46922,N_41127,N_40102);
nand U46923 (N_46923,N_40633,N_41773);
nand U46924 (N_46924,N_41566,N_44032);
and U46925 (N_46925,N_40912,N_42682);
and U46926 (N_46926,N_44911,N_41800);
xor U46927 (N_46927,N_43921,N_43199);
or U46928 (N_46928,N_43099,N_41276);
and U46929 (N_46929,N_43252,N_42326);
nand U46930 (N_46930,N_43266,N_41143);
or U46931 (N_46931,N_40831,N_44781);
or U46932 (N_46932,N_41903,N_41753);
nor U46933 (N_46933,N_42693,N_41457);
nor U46934 (N_46934,N_42372,N_41037);
and U46935 (N_46935,N_42425,N_43701);
nand U46936 (N_46936,N_43785,N_40863);
xor U46937 (N_46937,N_42501,N_42437);
or U46938 (N_46938,N_44923,N_41244);
or U46939 (N_46939,N_41393,N_42639);
xor U46940 (N_46940,N_42728,N_40866);
and U46941 (N_46941,N_41286,N_41683);
xor U46942 (N_46942,N_41291,N_44287);
nor U46943 (N_46943,N_44352,N_43796);
or U46944 (N_46944,N_41305,N_43167);
nor U46945 (N_46945,N_41102,N_44399);
and U46946 (N_46946,N_44202,N_41135);
or U46947 (N_46947,N_42128,N_40343);
or U46948 (N_46948,N_43805,N_40221);
and U46949 (N_46949,N_40280,N_41899);
nor U46950 (N_46950,N_43050,N_43189);
xnor U46951 (N_46951,N_40289,N_42651);
or U46952 (N_46952,N_42870,N_44234);
nor U46953 (N_46953,N_42431,N_42438);
nor U46954 (N_46954,N_41546,N_41494);
or U46955 (N_46955,N_40719,N_43837);
nand U46956 (N_46956,N_41840,N_42224);
nand U46957 (N_46957,N_43149,N_40115);
or U46958 (N_46958,N_41879,N_40311);
or U46959 (N_46959,N_43949,N_42665);
and U46960 (N_46960,N_41072,N_44144);
and U46961 (N_46961,N_44275,N_44634);
xor U46962 (N_46962,N_44921,N_41623);
nor U46963 (N_46963,N_43141,N_43636);
or U46964 (N_46964,N_40442,N_41709);
xor U46965 (N_46965,N_43522,N_44926);
and U46966 (N_46966,N_44636,N_43273);
xor U46967 (N_46967,N_42915,N_42385);
xnor U46968 (N_46968,N_40455,N_40604);
or U46969 (N_46969,N_44098,N_42112);
nand U46970 (N_46970,N_40634,N_40717);
nand U46971 (N_46971,N_40845,N_41586);
nand U46972 (N_46972,N_43358,N_41069);
nand U46973 (N_46973,N_40768,N_40464);
nor U46974 (N_46974,N_40655,N_41942);
xor U46975 (N_46975,N_40309,N_40624);
nand U46976 (N_46976,N_44037,N_41309);
or U46977 (N_46977,N_42004,N_40689);
and U46978 (N_46978,N_40056,N_40850);
nor U46979 (N_46979,N_41453,N_40591);
nand U46980 (N_46980,N_43938,N_43004);
nand U46981 (N_46981,N_44330,N_40220);
xor U46982 (N_46982,N_44717,N_40784);
and U46983 (N_46983,N_44718,N_44052);
and U46984 (N_46984,N_40961,N_42228);
and U46985 (N_46985,N_40157,N_40572);
nand U46986 (N_46986,N_42826,N_42394);
and U46987 (N_46987,N_43523,N_42656);
xor U46988 (N_46988,N_43098,N_42679);
xor U46989 (N_46989,N_43957,N_41747);
xor U46990 (N_46990,N_42367,N_41670);
and U46991 (N_46991,N_42498,N_42026);
nand U46992 (N_46992,N_41065,N_40914);
nor U46993 (N_46993,N_44299,N_43860);
xnor U46994 (N_46994,N_43270,N_40349);
nor U46995 (N_46995,N_42121,N_40329);
xnor U46996 (N_46996,N_40652,N_44104);
nor U46997 (N_46997,N_42721,N_44354);
xnor U46998 (N_46998,N_43112,N_43222);
nor U46999 (N_46999,N_41608,N_40172);
or U47000 (N_47000,N_44509,N_41585);
nor U47001 (N_47001,N_42938,N_42324);
nand U47002 (N_47002,N_43486,N_42306);
and U47003 (N_47003,N_43766,N_41374);
xor U47004 (N_47004,N_43324,N_40758);
nand U47005 (N_47005,N_42608,N_43073);
or U47006 (N_47006,N_44729,N_44099);
xor U47007 (N_47007,N_40769,N_43294);
or U47008 (N_47008,N_44195,N_40559);
nor U47009 (N_47009,N_44147,N_42771);
or U47010 (N_47010,N_40228,N_43092);
nand U47011 (N_47011,N_44521,N_43789);
nand U47012 (N_47012,N_40750,N_40170);
and U47013 (N_47013,N_43319,N_40480);
or U47014 (N_47014,N_40388,N_44331);
and U47015 (N_47015,N_43754,N_40246);
or U47016 (N_47016,N_42977,N_42231);
xor U47017 (N_47017,N_40799,N_41867);
nor U47018 (N_47018,N_42919,N_40267);
nor U47019 (N_47019,N_43120,N_42965);
xor U47020 (N_47020,N_44033,N_42288);
xor U47021 (N_47021,N_42934,N_41986);
or U47022 (N_47022,N_42557,N_44909);
and U47023 (N_47023,N_41006,N_40613);
nor U47024 (N_47024,N_41580,N_44664);
nor U47025 (N_47025,N_44973,N_42484);
xnor U47026 (N_47026,N_41865,N_40786);
and U47027 (N_47027,N_44298,N_43084);
nor U47028 (N_47028,N_43029,N_42269);
or U47029 (N_47029,N_40361,N_40222);
and U47030 (N_47030,N_44961,N_43341);
or U47031 (N_47031,N_42520,N_41447);
and U47032 (N_47032,N_40880,N_40436);
or U47033 (N_47033,N_43542,N_42953);
nand U47034 (N_47034,N_42708,N_40690);
xor U47035 (N_47035,N_43447,N_42205);
and U47036 (N_47036,N_44997,N_40659);
and U47037 (N_47037,N_43223,N_42548);
nor U47038 (N_47038,N_43080,N_40674);
and U47039 (N_47039,N_42167,N_40852);
nor U47040 (N_47040,N_44101,N_40183);
and U47041 (N_47041,N_40767,N_44749);
and U47042 (N_47042,N_44028,N_43367);
nor U47043 (N_47043,N_43202,N_40526);
and U47044 (N_47044,N_43356,N_42111);
and U47045 (N_47045,N_41970,N_40194);
and U47046 (N_47046,N_42582,N_41968);
xor U47047 (N_47047,N_40043,N_42714);
or U47048 (N_47048,N_44799,N_41326);
and U47049 (N_47049,N_44206,N_41336);
nand U47050 (N_47050,N_42271,N_43478);
and U47051 (N_47051,N_41844,N_41976);
or U47052 (N_47052,N_40856,N_42016);
nand U47053 (N_47053,N_40954,N_43656);
and U47054 (N_47054,N_44230,N_43669);
nor U47055 (N_47055,N_41198,N_41017);
or U47056 (N_47056,N_41485,N_41829);
nor U47057 (N_47057,N_44912,N_40862);
nor U47058 (N_47058,N_41898,N_42775);
nand U47059 (N_47059,N_43135,N_40728);
nor U47060 (N_47060,N_40520,N_43436);
nor U47061 (N_47061,N_41517,N_43333);
or U47062 (N_47062,N_44267,N_42311);
xnor U47063 (N_47063,N_44162,N_41157);
nor U47064 (N_47064,N_41599,N_42857);
xor U47065 (N_47065,N_42829,N_43427);
or U47066 (N_47066,N_42466,N_42563);
nand U47067 (N_47067,N_40186,N_42318);
or U47068 (N_47068,N_40936,N_42778);
and U47069 (N_47069,N_44384,N_42629);
nor U47070 (N_47070,N_40154,N_42571);
nor U47071 (N_47071,N_42211,N_41707);
or U47072 (N_47072,N_43739,N_42847);
or U47073 (N_47073,N_44084,N_43584);
nand U47074 (N_47074,N_41519,N_44667);
nor U47075 (N_47075,N_41853,N_44730);
or U47076 (N_47076,N_40959,N_44886);
nand U47077 (N_47077,N_43516,N_42553);
nor U47078 (N_47078,N_43336,N_40059);
and U47079 (N_47079,N_44881,N_42075);
xor U47080 (N_47080,N_42223,N_44739);
nor U47081 (N_47081,N_42090,N_43151);
nor U47082 (N_47082,N_42792,N_42724);
or U47083 (N_47083,N_40071,N_40302);
xnor U47084 (N_47084,N_41466,N_41361);
and U47085 (N_47085,N_41776,N_41480);
or U47086 (N_47086,N_43548,N_43055);
nor U47087 (N_47087,N_40506,N_40275);
or U47088 (N_47088,N_40128,N_43414);
or U47089 (N_47089,N_40589,N_44108);
or U47090 (N_47090,N_43246,N_43839);
or U47091 (N_47091,N_43862,N_42044);
nor U47092 (N_47092,N_43975,N_41648);
or U47093 (N_47093,N_43515,N_40023);
nor U47094 (N_47094,N_43635,N_43271);
or U47095 (N_47095,N_42976,N_43275);
nand U47096 (N_47096,N_41495,N_41002);
nor U47097 (N_47097,N_43068,N_44314);
or U47098 (N_47098,N_40213,N_44151);
nor U47099 (N_47099,N_44692,N_40379);
and U47100 (N_47100,N_42305,N_44484);
nor U47101 (N_47101,N_44951,N_41311);
and U47102 (N_47102,N_44091,N_43253);
and U47103 (N_47103,N_43958,N_44901);
nand U47104 (N_47104,N_44295,N_41152);
and U47105 (N_47105,N_42918,N_40035);
and U47106 (N_47106,N_40308,N_40475);
or U47107 (N_47107,N_43506,N_44481);
nand U47108 (N_47108,N_44232,N_42646);
and U47109 (N_47109,N_42155,N_40240);
and U47110 (N_47110,N_42064,N_41003);
or U47111 (N_47111,N_43695,N_43218);
xnor U47112 (N_47112,N_43753,N_43767);
or U47113 (N_47113,N_43262,N_42672);
or U47114 (N_47114,N_44638,N_43956);
nor U47115 (N_47115,N_40120,N_41668);
nand U47116 (N_47116,N_40024,N_44873);
and U47117 (N_47117,N_42312,N_43970);
nand U47118 (N_47118,N_40100,N_43177);
nor U47119 (N_47119,N_43633,N_42096);
and U47120 (N_47120,N_41217,N_44203);
xnor U47121 (N_47121,N_42422,N_41506);
nand U47122 (N_47122,N_43873,N_40721);
xnor U47123 (N_47123,N_42801,N_42992);
nand U47124 (N_47124,N_40687,N_43385);
nand U47125 (N_47125,N_41617,N_41563);
or U47126 (N_47126,N_43703,N_40521);
and U47127 (N_47127,N_40667,N_41377);
xor U47128 (N_47128,N_40079,N_44445);
and U47129 (N_47129,N_44313,N_43180);
nor U47130 (N_47130,N_44268,N_42142);
or U47131 (N_47131,N_42702,N_40331);
or U47132 (N_47132,N_43550,N_40127);
xor U47133 (N_47133,N_42085,N_44105);
xor U47134 (N_47134,N_41516,N_43715);
or U47135 (N_47135,N_40823,N_43481);
and U47136 (N_47136,N_40395,N_41031);
or U47137 (N_47137,N_40420,N_40626);
or U47138 (N_47138,N_44687,N_41114);
nor U47139 (N_47139,N_41975,N_42418);
nand U47140 (N_47140,N_42821,N_40920);
xnor U47141 (N_47141,N_42061,N_42872);
nand U47142 (N_47142,N_43595,N_44843);
or U47143 (N_47143,N_44958,N_42634);
or U47144 (N_47144,N_42160,N_43045);
or U47145 (N_47145,N_43316,N_41112);
and U47146 (N_47146,N_40380,N_42315);
or U47147 (N_47147,N_43116,N_41984);
or U47148 (N_47148,N_43030,N_41373);
nand U47149 (N_47149,N_44285,N_40093);
nand U47150 (N_47150,N_42574,N_40967);
nand U47151 (N_47151,N_41869,N_40200);
nor U47152 (N_47152,N_40339,N_44686);
or U47153 (N_47153,N_42745,N_40368);
and U47154 (N_47154,N_42151,N_41284);
or U47155 (N_47155,N_43685,N_42132);
and U47156 (N_47156,N_43886,N_42811);
nand U47157 (N_47157,N_40697,N_44415);
and U47158 (N_47158,N_40873,N_40317);
xnor U47159 (N_47159,N_44143,N_44020);
xnor U47160 (N_47160,N_41482,N_44328);
nand U47161 (N_47161,N_42036,N_40803);
nor U47162 (N_47162,N_41954,N_40393);
nor U47163 (N_47163,N_41806,N_41245);
xnor U47164 (N_47164,N_44240,N_43274);
nand U47165 (N_47165,N_42163,N_43464);
xnor U47166 (N_47166,N_44296,N_42442);
and U47167 (N_47167,N_44341,N_42627);
nand U47168 (N_47168,N_44253,N_41632);
nor U47169 (N_47169,N_42754,N_43432);
nor U47170 (N_47170,N_44349,N_41348);
nand U47171 (N_47171,N_41620,N_42722);
nor U47172 (N_47172,N_43038,N_42156);
and U47173 (N_47173,N_44220,N_40149);
and U47174 (N_47174,N_41355,N_43826);
or U47175 (N_47175,N_41395,N_40009);
and U47176 (N_47176,N_41161,N_42100);
or U47177 (N_47177,N_42903,N_40666);
and U47178 (N_47178,N_43955,N_43104);
nor U47179 (N_47179,N_42731,N_44953);
or U47180 (N_47180,N_43400,N_44685);
nor U47181 (N_47181,N_40421,N_42428);
or U47182 (N_47182,N_41624,N_41576);
xor U47183 (N_47183,N_41812,N_41452);
xor U47184 (N_47184,N_42471,N_40636);
or U47185 (N_47185,N_44623,N_44465);
xor U47186 (N_47186,N_42861,N_42239);
nand U47187 (N_47187,N_40820,N_40467);
nand U47188 (N_47188,N_43094,N_41052);
and U47189 (N_47189,N_43388,N_43415);
xor U47190 (N_47190,N_40893,N_43894);
nor U47191 (N_47191,N_42172,N_42482);
nand U47192 (N_47192,N_43404,N_44196);
or U47193 (N_47193,N_40620,N_41295);
nand U47194 (N_47194,N_40860,N_42241);
and U47195 (N_47195,N_44038,N_43091);
nor U47196 (N_47196,N_44504,N_43238);
nor U47197 (N_47197,N_43150,N_43926);
nand U47198 (N_47198,N_44571,N_40989);
nor U47199 (N_47199,N_41146,N_44794);
and U47200 (N_47200,N_41795,N_43148);
or U47201 (N_47201,N_44856,N_44808);
and U47202 (N_47202,N_41873,N_42376);
or U47203 (N_47203,N_44107,N_44592);
nand U47204 (N_47204,N_44124,N_43644);
or U47205 (N_47205,N_41690,N_41727);
and U47206 (N_47206,N_42037,N_40577);
xnor U47207 (N_47207,N_44708,N_42071);
or U47208 (N_47208,N_44696,N_43418);
and U47209 (N_47209,N_44915,N_43840);
nor U47210 (N_47210,N_43797,N_41932);
nand U47211 (N_47211,N_40668,N_44506);
and U47212 (N_47212,N_43846,N_41258);
and U47213 (N_47213,N_43578,N_44583);
and U47214 (N_47214,N_41260,N_40114);
or U47215 (N_47215,N_43130,N_41364);
xor U47216 (N_47216,N_44398,N_44175);
xor U47217 (N_47217,N_44419,N_43882);
xor U47218 (N_47218,N_43283,N_44980);
or U47219 (N_47219,N_43193,N_44607);
nand U47220 (N_47220,N_44833,N_41014);
or U47221 (N_47221,N_44497,N_41934);
nor U47222 (N_47222,N_42032,N_44905);
or U47223 (N_47223,N_40469,N_41786);
nor U47224 (N_47224,N_43349,N_40333);
xor U47225 (N_47225,N_41793,N_43245);
or U47226 (N_47226,N_43420,N_42540);
or U47227 (N_47227,N_42464,N_41415);
or U47228 (N_47228,N_42764,N_44710);
and U47229 (N_47229,N_43126,N_42788);
nor U47230 (N_47230,N_44570,N_44792);
and U47231 (N_47231,N_43580,N_42961);
xnor U47232 (N_47232,N_44620,N_41757);
nor U47233 (N_47233,N_44784,N_42666);
and U47234 (N_47234,N_41404,N_40952);
xnor U47235 (N_47235,N_43178,N_40248);
or U47236 (N_47236,N_42362,N_42642);
or U47237 (N_47237,N_44700,N_44036);
nor U47238 (N_47238,N_43650,N_43519);
and U47239 (N_47239,N_41345,N_44831);
xnor U47240 (N_47240,N_43916,N_43286);
and U47241 (N_47241,N_41391,N_41833);
xor U47242 (N_47242,N_40670,N_42595);
nand U47243 (N_47243,N_40531,N_40053);
xor U47244 (N_47244,N_44892,N_44218);
xor U47245 (N_47245,N_43394,N_40884);
xor U47246 (N_47246,N_43863,N_44942);
nor U47247 (N_47247,N_42633,N_41525);
xor U47248 (N_47248,N_44711,N_43928);
xnor U47249 (N_47249,N_41416,N_43823);
nand U47250 (N_47250,N_42446,N_44609);
or U47251 (N_47251,N_40038,N_43298);
nor U47252 (N_47252,N_42752,N_44835);
xor U47253 (N_47253,N_41008,N_42490);
xor U47254 (N_47254,N_43733,N_44491);
nor U47255 (N_47255,N_40243,N_40021);
xnor U47256 (N_47256,N_42189,N_42856);
xor U47257 (N_47257,N_41521,N_41790);
nor U47258 (N_47258,N_41411,N_40054);
and U47259 (N_47259,N_40785,N_44207);
nor U47260 (N_47260,N_40519,N_41317);
or U47261 (N_47261,N_40603,N_44093);
xor U47262 (N_47262,N_40958,N_42282);
nand U47263 (N_47263,N_44170,N_44862);
nand U47264 (N_47264,N_42265,N_42562);
xor U47265 (N_47265,N_40036,N_40252);
nand U47266 (N_47266,N_40905,N_42199);
nor U47267 (N_47267,N_41054,N_42748);
nand U47268 (N_47268,N_44999,N_40454);
or U47269 (N_47269,N_42186,N_41726);
nand U47270 (N_47270,N_40492,N_41056);
nor U47271 (N_47271,N_44529,N_40904);
nand U47272 (N_47272,N_44750,N_43118);
or U47273 (N_47273,N_43017,N_42689);
nor U47274 (N_47274,N_40530,N_41210);
or U47275 (N_47275,N_42732,N_44899);
nand U47276 (N_47276,N_44448,N_44323);
nor U47277 (N_47277,N_44671,N_40483);
or U47278 (N_47278,N_42219,N_40693);
nor U47279 (N_47279,N_40493,N_44161);
nor U47280 (N_47280,N_40929,N_42551);
nor U47281 (N_47281,N_44089,N_41148);
or U47282 (N_47282,N_44847,N_43488);
xor U47283 (N_47283,N_41044,N_41863);
or U47284 (N_47284,N_42057,N_43660);
or U47285 (N_47285,N_41804,N_44725);
nand U47286 (N_47286,N_42080,N_40215);
and U47287 (N_47287,N_42921,N_41694);
or U47288 (N_47288,N_42159,N_40202);
or U47289 (N_47289,N_42051,N_41172);
nor U47290 (N_47290,N_42252,N_40007);
and U47291 (N_47291,N_40878,N_44610);
or U47292 (N_47292,N_40190,N_40898);
nor U47293 (N_47293,N_42566,N_44369);
nor U47294 (N_47294,N_43387,N_43340);
or U47295 (N_47295,N_41592,N_43124);
or U47296 (N_47296,N_40680,N_42278);
and U47297 (N_47297,N_42560,N_44039);
nand U47298 (N_47298,N_40461,N_43976);
or U47299 (N_47299,N_44789,N_40525);
and U47300 (N_47300,N_41289,N_43590);
or U47301 (N_47301,N_40754,N_41093);
and U47302 (N_47302,N_43610,N_40266);
nor U47303 (N_47303,N_41312,N_43373);
nand U47304 (N_47304,N_43076,N_44449);
or U47305 (N_47305,N_42066,N_44963);
and U47306 (N_47306,N_42294,N_40647);
nor U47307 (N_47307,N_41379,N_40426);
nand U47308 (N_47308,N_44372,N_41170);
xor U47309 (N_47309,N_42579,N_44764);
xnor U47310 (N_47310,N_42957,N_44668);
nand U47311 (N_47311,N_40982,N_41613);
xor U47312 (N_47312,N_40776,N_41667);
nor U47313 (N_47313,N_42330,N_43370);
nand U47314 (N_47314,N_40605,N_43643);
and U47315 (N_47315,N_40629,N_40089);
nor U47316 (N_47316,N_41664,N_40396);
nor U47317 (N_47317,N_40664,N_43330);
or U47318 (N_47318,N_42526,N_44707);
and U47319 (N_47319,N_42217,N_42741);
nand U47320 (N_47320,N_42979,N_42924);
and U47321 (N_47321,N_43232,N_44002);
xor U47322 (N_47322,N_44066,N_43310);
nor U47323 (N_47323,N_43158,N_44567);
and U47324 (N_47324,N_41571,N_43215);
nor U47325 (N_47325,N_41216,N_43680);
and U47326 (N_47326,N_40040,N_44672);
nor U47327 (N_47327,N_43048,N_44297);
nand U47328 (N_47328,N_41658,N_42119);
nand U47329 (N_47329,N_44996,N_43209);
nand U47330 (N_47330,N_43403,N_44011);
and U47331 (N_47331,N_44120,N_43259);
and U47332 (N_47332,N_40498,N_41481);
nand U47333 (N_47333,N_43745,N_41557);
and U47334 (N_47334,N_43953,N_42531);
xor U47335 (N_47335,N_44208,N_41327);
xor U47336 (N_47336,N_40378,N_44982);
and U47337 (N_47337,N_42260,N_40051);
nand U47338 (N_47338,N_44811,N_41966);
xnor U47339 (N_47339,N_41329,N_41280);
nand U47340 (N_47340,N_41251,N_43570);
or U47341 (N_47341,N_41387,N_40574);
or U47342 (N_47342,N_43727,N_40938);
nor U47343 (N_47343,N_41856,N_40028);
nor U47344 (N_47344,N_42116,N_44628);
nand U47345 (N_47345,N_42190,N_44156);
xor U47346 (N_47346,N_42178,N_41685);
and U47347 (N_47347,N_40409,N_41534);
xor U47348 (N_47348,N_44557,N_40000);
nor U47349 (N_47349,N_43672,N_43673);
or U47350 (N_47350,N_44994,N_43101);
or U47351 (N_47351,N_41803,N_40268);
xor U47352 (N_47352,N_40097,N_44523);
and U47353 (N_47353,N_43768,N_40293);
nor U47354 (N_47354,N_41267,N_42625);
nand U47355 (N_47355,N_40296,N_40544);
nand U47356 (N_47356,N_43582,N_43026);
nor U47357 (N_47357,N_40999,N_43577);
nor U47358 (N_47358,N_41015,N_41971);
or U47359 (N_47359,N_40722,N_40075);
nor U47360 (N_47360,N_43609,N_43829);
xor U47361 (N_47361,N_41107,N_41978);
xnor U47362 (N_47362,N_43555,N_43285);
or U47363 (N_47363,N_40716,N_43474);
nand U47364 (N_47364,N_41259,N_42025);
nand U47365 (N_47365,N_42718,N_44114);
or U47366 (N_47366,N_44422,N_42819);
xnor U47367 (N_47367,N_41661,N_40002);
nor U47368 (N_47368,N_40151,N_42029);
nand U47369 (N_47369,N_44434,N_40944);
nor U47370 (N_47370,N_43912,N_43109);
xor U47371 (N_47371,N_40847,N_41810);
nand U47372 (N_47372,N_41100,N_44188);
or U47373 (N_47373,N_44396,N_42328);
or U47374 (N_47374,N_43230,N_43814);
and U47375 (N_47375,N_43107,N_41680);
nand U47376 (N_47376,N_42361,N_42302);
and U47377 (N_47377,N_42556,N_42443);
nor U47378 (N_47378,N_43960,N_41814);
and U47379 (N_47379,N_43906,N_40334);
xor U47380 (N_47380,N_42489,N_41734);
nand U47381 (N_47381,N_43599,N_43039);
nand U47382 (N_47382,N_43140,N_44123);
and U47383 (N_47383,N_41214,N_43806);
nand U47384 (N_47384,N_42524,N_42652);
or U47385 (N_47385,N_44731,N_43564);
xnor U47386 (N_47386,N_41559,N_44071);
xor U47387 (N_47387,N_41354,N_43292);
xnor U47388 (N_47388,N_43651,N_44550);
xor U47389 (N_47389,N_41212,N_40205);
nand U47390 (N_47390,N_41555,N_40173);
nand U47391 (N_47391,N_41155,N_43393);
or U47392 (N_47392,N_44322,N_41337);
nand U47393 (N_47393,N_40239,N_41801);
nand U47394 (N_47394,N_42550,N_44353);
nor U47395 (N_47395,N_40472,N_40919);
nand U47396 (N_47396,N_44507,N_41675);
nor U47397 (N_47397,N_40137,N_40546);
nor U47398 (N_47398,N_43904,N_42458);
and U47399 (N_47399,N_43013,N_44137);
nor U47400 (N_47400,N_43569,N_42906);
and U47401 (N_47401,N_44969,N_40819);
nand U47402 (N_47402,N_43981,N_41454);
and U47403 (N_47403,N_43160,N_44590);
or U47404 (N_47404,N_42949,N_41751);
nand U47405 (N_47405,N_42621,N_42053);
and U47406 (N_47406,N_40540,N_43507);
xnor U47407 (N_47407,N_42780,N_41279);
or U47408 (N_47408,N_40306,N_43596);
nor U47409 (N_47409,N_44771,N_40828);
and U47410 (N_47410,N_40370,N_44712);
xnor U47411 (N_47411,N_41060,N_41884);
nand U47412 (N_47412,N_41509,N_41160);
and U47413 (N_47413,N_41921,N_42382);
xnor U47414 (N_47414,N_44675,N_41866);
nor U47415 (N_47415,N_41720,N_44875);
and U47416 (N_47416,N_42195,N_40447);
nand U47417 (N_47417,N_44051,N_43268);
or U47418 (N_47418,N_44097,N_42534);
and U47419 (N_47419,N_41953,N_43554);
or U47420 (N_47420,N_40273,N_42944);
and U47421 (N_47421,N_44360,N_43967);
xor U47422 (N_47422,N_43925,N_42716);
nand U47423 (N_47423,N_40968,N_42670);
xnor U47424 (N_47424,N_44293,N_40011);
xor U47425 (N_47425,N_44660,N_43661);
and U47426 (N_47426,N_42892,N_42839);
xnor U47427 (N_47427,N_42587,N_42002);
xor U47428 (N_47428,N_43185,N_42581);
nand U47429 (N_47429,N_42932,N_44302);
nor U47430 (N_47430,N_42073,N_40391);
nand U47431 (N_47431,N_44548,N_40829);
or U47432 (N_47432,N_43528,N_42347);
xor U47433 (N_47433,N_42543,N_42967);
and U47434 (N_47434,N_41475,N_44453);
nor U47435 (N_47435,N_43830,N_40612);
nand U47436 (N_47436,N_43631,N_44035);
nor U47437 (N_47437,N_41344,N_44754);
nor U47438 (N_47438,N_40855,N_44524);
nor U47439 (N_47439,N_42594,N_40713);
nor U47440 (N_47440,N_41263,N_40686);
nand U47441 (N_47441,N_41218,N_43678);
and U47442 (N_47442,N_41371,N_41079);
nor U47443 (N_47443,N_40592,N_41692);
and U47444 (N_47444,N_44438,N_40800);
nor U47445 (N_47445,N_44809,N_43411);
and U47446 (N_47446,N_44990,N_40532);
or U47447 (N_47447,N_44027,N_40344);
xor U47448 (N_47448,N_40657,N_44178);
nand U47449 (N_47449,N_44879,N_42492);
and U47450 (N_47450,N_40827,N_44358);
nand U47451 (N_47451,N_40459,N_43874);
nor U47452 (N_47452,N_40808,N_41950);
nor U47453 (N_47453,N_44450,N_44505);
nor U47454 (N_47454,N_44966,N_43169);
xnor U47455 (N_47455,N_43717,N_44190);
nand U47456 (N_47456,N_41461,N_43145);
xor U47457 (N_47457,N_40377,N_44078);
and U47458 (N_47458,N_43877,N_42815);
or U47459 (N_47459,N_44117,N_44092);
and U47460 (N_47460,N_42307,N_40030);
and U47461 (N_47461,N_41811,N_43867);
nor U47462 (N_47462,N_40779,N_43455);
and U47463 (N_47463,N_42072,N_43034);
nand U47464 (N_47464,N_42573,N_41718);
or U47465 (N_47465,N_42790,N_41813);
or U47466 (N_47466,N_41958,N_44284);
or U47467 (N_47467,N_41224,N_42558);
or U47468 (N_47468,N_40405,N_40476);
nor U47469 (N_47469,N_44795,N_44213);
or U47470 (N_47470,N_44702,N_44551);
nand U47471 (N_47471,N_40918,N_44716);
nor U47472 (N_47472,N_44441,N_40010);
xnor U47473 (N_47473,N_41483,N_43624);
nor U47474 (N_47474,N_41920,N_43290);
xor U47475 (N_47475,N_43217,N_43062);
nand U47476 (N_47476,N_40406,N_41220);
xnor U47477 (N_47477,N_41301,N_43980);
nand U47478 (N_47478,N_40367,N_41544);
nor U47479 (N_47479,N_42469,N_40701);
xnor U47480 (N_47480,N_41246,N_44787);
or U47481 (N_47481,N_43653,N_42088);
and U47482 (N_47482,N_42386,N_41232);
or U47483 (N_47483,N_43546,N_41500);
nand U47484 (N_47484,N_43825,N_43600);
and U47485 (N_47485,N_41860,N_41300);
nand U47486 (N_47486,N_41542,N_44476);
nand U47487 (N_47487,N_40354,N_43566);
or U47488 (N_47488,N_41702,N_41512);
and U47489 (N_47489,N_40802,N_40571);
or U47490 (N_47490,N_41564,N_41645);
nor U47491 (N_47491,N_42060,N_44155);
or U47492 (N_47492,N_44288,N_40108);
xor U47493 (N_47493,N_42038,N_41991);
nor U47494 (N_47494,N_44597,N_44959);
xor U47495 (N_47495,N_40514,N_44247);
nand U47496 (N_47496,N_43343,N_41458);
and U47497 (N_47497,N_41206,N_40106);
nand U47498 (N_47498,N_41315,N_43304);
or U47499 (N_47499,N_41777,N_43354);
or U47500 (N_47500,N_41400,N_40475);
nor U47501 (N_47501,N_41330,N_42491);
nor U47502 (N_47502,N_42182,N_40831);
xor U47503 (N_47503,N_40236,N_43342);
or U47504 (N_47504,N_43579,N_43589);
nand U47505 (N_47505,N_43865,N_41621);
xnor U47506 (N_47506,N_44315,N_44755);
and U47507 (N_47507,N_43028,N_43252);
xor U47508 (N_47508,N_43400,N_44279);
nor U47509 (N_47509,N_40621,N_41433);
nand U47510 (N_47510,N_41280,N_41882);
xnor U47511 (N_47511,N_41284,N_43755);
nor U47512 (N_47512,N_43004,N_41270);
xor U47513 (N_47513,N_40545,N_44217);
and U47514 (N_47514,N_40594,N_40368);
nor U47515 (N_47515,N_43515,N_42478);
nand U47516 (N_47516,N_40391,N_42540);
nor U47517 (N_47517,N_40104,N_42188);
and U47518 (N_47518,N_40766,N_43778);
or U47519 (N_47519,N_43384,N_44649);
or U47520 (N_47520,N_40883,N_41359);
xor U47521 (N_47521,N_43663,N_43556);
nand U47522 (N_47522,N_40511,N_40285);
xor U47523 (N_47523,N_41674,N_44665);
and U47524 (N_47524,N_43252,N_41077);
xnor U47525 (N_47525,N_44948,N_41715);
nor U47526 (N_47526,N_43926,N_42457);
xnor U47527 (N_47527,N_40465,N_43447);
nor U47528 (N_47528,N_40275,N_40550);
nor U47529 (N_47529,N_43863,N_41882);
xnor U47530 (N_47530,N_40040,N_41962);
xor U47531 (N_47531,N_42868,N_42913);
nor U47532 (N_47532,N_41573,N_44505);
xnor U47533 (N_47533,N_40627,N_42487);
xor U47534 (N_47534,N_41357,N_40144);
or U47535 (N_47535,N_42626,N_41580);
nor U47536 (N_47536,N_42923,N_44074);
xnor U47537 (N_47537,N_42319,N_42566);
nand U47538 (N_47538,N_41893,N_40924);
nand U47539 (N_47539,N_43176,N_41427);
nor U47540 (N_47540,N_42917,N_40681);
xnor U47541 (N_47541,N_44632,N_40027);
nor U47542 (N_47542,N_41699,N_43785);
nand U47543 (N_47543,N_44206,N_42137);
nor U47544 (N_47544,N_42057,N_43207);
nand U47545 (N_47545,N_43407,N_44619);
or U47546 (N_47546,N_44059,N_41140);
or U47547 (N_47547,N_43673,N_41586);
nand U47548 (N_47548,N_40295,N_43871);
or U47549 (N_47549,N_44916,N_42683);
nor U47550 (N_47550,N_40886,N_43025);
xor U47551 (N_47551,N_41505,N_42152);
xnor U47552 (N_47552,N_43573,N_43141);
or U47553 (N_47553,N_42132,N_41609);
or U47554 (N_47554,N_41317,N_43098);
or U47555 (N_47555,N_43925,N_40064);
xor U47556 (N_47556,N_43641,N_44489);
xnor U47557 (N_47557,N_41437,N_42924);
xor U47558 (N_47558,N_44579,N_40149);
or U47559 (N_47559,N_41456,N_42346);
nand U47560 (N_47560,N_43367,N_43201);
or U47561 (N_47561,N_42459,N_42623);
and U47562 (N_47562,N_43829,N_40793);
xnor U47563 (N_47563,N_42332,N_43636);
or U47564 (N_47564,N_42626,N_44860);
and U47565 (N_47565,N_44175,N_43629);
and U47566 (N_47566,N_44153,N_43810);
and U47567 (N_47567,N_44595,N_42329);
nand U47568 (N_47568,N_41773,N_41462);
and U47569 (N_47569,N_40451,N_42387);
or U47570 (N_47570,N_42121,N_40094);
and U47571 (N_47571,N_41218,N_40822);
xor U47572 (N_47572,N_44905,N_43433);
nand U47573 (N_47573,N_42460,N_42772);
nor U47574 (N_47574,N_42510,N_43238);
nand U47575 (N_47575,N_43063,N_43428);
nor U47576 (N_47576,N_44322,N_41399);
and U47577 (N_47577,N_44862,N_43585);
nor U47578 (N_47578,N_41628,N_43830);
or U47579 (N_47579,N_43466,N_44294);
nor U47580 (N_47580,N_44392,N_43956);
nand U47581 (N_47581,N_44808,N_40104);
xor U47582 (N_47582,N_44350,N_44570);
nand U47583 (N_47583,N_41572,N_44045);
nand U47584 (N_47584,N_43033,N_40188);
nor U47585 (N_47585,N_40641,N_41132);
or U47586 (N_47586,N_40775,N_40725);
and U47587 (N_47587,N_42755,N_43877);
nor U47588 (N_47588,N_44520,N_43451);
or U47589 (N_47589,N_42166,N_44955);
nand U47590 (N_47590,N_41304,N_44452);
and U47591 (N_47591,N_43045,N_44284);
and U47592 (N_47592,N_44512,N_43168);
xnor U47593 (N_47593,N_41367,N_44143);
and U47594 (N_47594,N_43045,N_40866);
and U47595 (N_47595,N_41596,N_41455);
and U47596 (N_47596,N_44972,N_42890);
and U47597 (N_47597,N_41225,N_44472);
nand U47598 (N_47598,N_43456,N_44036);
or U47599 (N_47599,N_41116,N_43336);
and U47600 (N_47600,N_40134,N_42502);
nand U47601 (N_47601,N_44596,N_42669);
or U47602 (N_47602,N_41315,N_44861);
or U47603 (N_47603,N_44807,N_41876);
xnor U47604 (N_47604,N_42548,N_42250);
or U47605 (N_47605,N_44303,N_40799);
or U47606 (N_47606,N_44090,N_43117);
xnor U47607 (N_47607,N_42983,N_40612);
nor U47608 (N_47608,N_41587,N_42382);
nand U47609 (N_47609,N_40396,N_41731);
nand U47610 (N_47610,N_41665,N_41550);
or U47611 (N_47611,N_42058,N_41242);
and U47612 (N_47612,N_42190,N_44545);
nor U47613 (N_47613,N_43602,N_40082);
and U47614 (N_47614,N_44010,N_40235);
nor U47615 (N_47615,N_41001,N_41404);
nand U47616 (N_47616,N_41657,N_40358);
xor U47617 (N_47617,N_41079,N_44357);
nand U47618 (N_47618,N_44054,N_41595);
nand U47619 (N_47619,N_40917,N_40561);
xnor U47620 (N_47620,N_43000,N_41903);
or U47621 (N_47621,N_43298,N_44301);
nor U47622 (N_47622,N_43748,N_44722);
and U47623 (N_47623,N_41853,N_43343);
xor U47624 (N_47624,N_42566,N_44779);
nand U47625 (N_47625,N_43337,N_40077);
nor U47626 (N_47626,N_40461,N_40849);
xor U47627 (N_47627,N_42606,N_43552);
and U47628 (N_47628,N_40730,N_42639);
and U47629 (N_47629,N_44360,N_41959);
or U47630 (N_47630,N_40894,N_42927);
and U47631 (N_47631,N_43726,N_44371);
xnor U47632 (N_47632,N_40453,N_42860);
nor U47633 (N_47633,N_41922,N_42421);
or U47634 (N_47634,N_40910,N_43075);
nor U47635 (N_47635,N_41610,N_43002);
nor U47636 (N_47636,N_42146,N_41455);
xnor U47637 (N_47637,N_42997,N_41628);
and U47638 (N_47638,N_40434,N_44201);
or U47639 (N_47639,N_41445,N_44384);
nand U47640 (N_47640,N_44363,N_41680);
nor U47641 (N_47641,N_41947,N_41240);
nor U47642 (N_47642,N_40375,N_43150);
and U47643 (N_47643,N_42404,N_42945);
nor U47644 (N_47644,N_41827,N_42642);
xor U47645 (N_47645,N_42252,N_42546);
and U47646 (N_47646,N_44665,N_41519);
nor U47647 (N_47647,N_44121,N_40455);
nor U47648 (N_47648,N_42909,N_40572);
nor U47649 (N_47649,N_41697,N_42547);
nor U47650 (N_47650,N_41997,N_41586);
nor U47651 (N_47651,N_43933,N_41639);
and U47652 (N_47652,N_40562,N_44442);
nand U47653 (N_47653,N_41193,N_42806);
and U47654 (N_47654,N_43450,N_44587);
nor U47655 (N_47655,N_44773,N_40939);
or U47656 (N_47656,N_43600,N_40378);
or U47657 (N_47657,N_43576,N_41268);
or U47658 (N_47658,N_41787,N_42527);
or U47659 (N_47659,N_44332,N_40718);
nor U47660 (N_47660,N_42040,N_44397);
nand U47661 (N_47661,N_40459,N_41176);
nand U47662 (N_47662,N_43497,N_44172);
and U47663 (N_47663,N_42109,N_42616);
or U47664 (N_47664,N_43103,N_40183);
nor U47665 (N_47665,N_40155,N_43922);
nand U47666 (N_47666,N_43114,N_42491);
nand U47667 (N_47667,N_42421,N_40667);
xnor U47668 (N_47668,N_42585,N_43630);
xnor U47669 (N_47669,N_42686,N_41636);
xnor U47670 (N_47670,N_43828,N_42109);
and U47671 (N_47671,N_40060,N_44086);
nand U47672 (N_47672,N_44999,N_41592);
or U47673 (N_47673,N_43206,N_43104);
nor U47674 (N_47674,N_43840,N_43444);
xor U47675 (N_47675,N_44624,N_41061);
or U47676 (N_47676,N_41354,N_40786);
nand U47677 (N_47677,N_44692,N_41527);
xor U47678 (N_47678,N_42448,N_43539);
or U47679 (N_47679,N_41189,N_40564);
nor U47680 (N_47680,N_43028,N_41493);
or U47681 (N_47681,N_44528,N_43333);
nor U47682 (N_47682,N_44275,N_41370);
or U47683 (N_47683,N_44504,N_41863);
or U47684 (N_47684,N_43434,N_43587);
and U47685 (N_47685,N_41535,N_41164);
or U47686 (N_47686,N_41372,N_40527);
and U47687 (N_47687,N_43110,N_40226);
and U47688 (N_47688,N_41675,N_44331);
and U47689 (N_47689,N_43030,N_40119);
xor U47690 (N_47690,N_40753,N_41092);
nand U47691 (N_47691,N_43129,N_44118);
and U47692 (N_47692,N_44284,N_41091);
nor U47693 (N_47693,N_43984,N_43908);
nor U47694 (N_47694,N_44238,N_42151);
nor U47695 (N_47695,N_40107,N_40699);
xor U47696 (N_47696,N_42361,N_42553);
nand U47697 (N_47697,N_43776,N_43982);
nor U47698 (N_47698,N_42011,N_42578);
xnor U47699 (N_47699,N_41699,N_41458);
xor U47700 (N_47700,N_43210,N_40173);
and U47701 (N_47701,N_40960,N_43653);
nand U47702 (N_47702,N_42751,N_43460);
xor U47703 (N_47703,N_40962,N_43845);
nor U47704 (N_47704,N_44909,N_41872);
and U47705 (N_47705,N_41845,N_43228);
nand U47706 (N_47706,N_43718,N_41372);
and U47707 (N_47707,N_41223,N_41063);
and U47708 (N_47708,N_42925,N_42980);
xnor U47709 (N_47709,N_43036,N_40918);
nor U47710 (N_47710,N_41106,N_43620);
and U47711 (N_47711,N_44497,N_42887);
or U47712 (N_47712,N_41002,N_43166);
and U47713 (N_47713,N_44336,N_43322);
and U47714 (N_47714,N_44861,N_42289);
and U47715 (N_47715,N_42103,N_41292);
and U47716 (N_47716,N_42883,N_41395);
nor U47717 (N_47717,N_40023,N_43121);
nor U47718 (N_47718,N_43586,N_40670);
and U47719 (N_47719,N_41301,N_44064);
nor U47720 (N_47720,N_42768,N_43851);
nand U47721 (N_47721,N_43081,N_41861);
nand U47722 (N_47722,N_42667,N_41749);
and U47723 (N_47723,N_43292,N_43297);
and U47724 (N_47724,N_44813,N_42509);
and U47725 (N_47725,N_42024,N_40144);
and U47726 (N_47726,N_40898,N_42305);
nand U47727 (N_47727,N_41541,N_44854);
nor U47728 (N_47728,N_41610,N_43645);
xor U47729 (N_47729,N_40767,N_44275);
and U47730 (N_47730,N_41212,N_42260);
nor U47731 (N_47731,N_40476,N_44064);
xor U47732 (N_47732,N_43837,N_41776);
xor U47733 (N_47733,N_40827,N_40239);
nor U47734 (N_47734,N_40356,N_43857);
or U47735 (N_47735,N_42539,N_43535);
xor U47736 (N_47736,N_41781,N_40736);
nor U47737 (N_47737,N_42859,N_42644);
or U47738 (N_47738,N_40317,N_44249);
nor U47739 (N_47739,N_44216,N_43781);
xnor U47740 (N_47740,N_44083,N_41937);
xor U47741 (N_47741,N_43171,N_41709);
nor U47742 (N_47742,N_44820,N_43238);
nand U47743 (N_47743,N_40873,N_43636);
and U47744 (N_47744,N_44313,N_42256);
xnor U47745 (N_47745,N_40250,N_40813);
or U47746 (N_47746,N_42394,N_42684);
and U47747 (N_47747,N_42542,N_44646);
or U47748 (N_47748,N_43249,N_40332);
or U47749 (N_47749,N_41963,N_40812);
nor U47750 (N_47750,N_40536,N_42022);
nand U47751 (N_47751,N_41451,N_41794);
nand U47752 (N_47752,N_40869,N_40746);
nor U47753 (N_47753,N_40746,N_41138);
xor U47754 (N_47754,N_42908,N_44322);
nand U47755 (N_47755,N_40162,N_40389);
nand U47756 (N_47756,N_40284,N_41613);
nor U47757 (N_47757,N_42091,N_41526);
and U47758 (N_47758,N_43974,N_43402);
nand U47759 (N_47759,N_44966,N_40875);
nand U47760 (N_47760,N_40177,N_42667);
or U47761 (N_47761,N_43797,N_43560);
xnor U47762 (N_47762,N_40282,N_44956);
nand U47763 (N_47763,N_40407,N_40642);
and U47764 (N_47764,N_40586,N_40124);
and U47765 (N_47765,N_43719,N_44049);
nand U47766 (N_47766,N_44691,N_44320);
nand U47767 (N_47767,N_44675,N_43627);
nand U47768 (N_47768,N_43198,N_41461);
or U47769 (N_47769,N_42339,N_44951);
or U47770 (N_47770,N_44594,N_44067);
nand U47771 (N_47771,N_40204,N_40560);
or U47772 (N_47772,N_42372,N_42272);
nor U47773 (N_47773,N_40862,N_42050);
and U47774 (N_47774,N_40721,N_41118);
and U47775 (N_47775,N_42174,N_44944);
xor U47776 (N_47776,N_40032,N_42581);
nand U47777 (N_47777,N_42020,N_43916);
nor U47778 (N_47778,N_44728,N_44145);
and U47779 (N_47779,N_43926,N_43749);
or U47780 (N_47780,N_40960,N_43026);
and U47781 (N_47781,N_42068,N_40578);
xnor U47782 (N_47782,N_41452,N_43003);
or U47783 (N_47783,N_44163,N_41781);
or U47784 (N_47784,N_42194,N_43444);
nand U47785 (N_47785,N_42770,N_40655);
and U47786 (N_47786,N_40111,N_41183);
and U47787 (N_47787,N_44226,N_42539);
xnor U47788 (N_47788,N_41814,N_40429);
nor U47789 (N_47789,N_40836,N_41211);
nand U47790 (N_47790,N_44790,N_41464);
nand U47791 (N_47791,N_40093,N_42465);
and U47792 (N_47792,N_43180,N_43661);
nor U47793 (N_47793,N_43705,N_43168);
nor U47794 (N_47794,N_43690,N_40470);
or U47795 (N_47795,N_40376,N_41416);
and U47796 (N_47796,N_44258,N_43367);
or U47797 (N_47797,N_40291,N_40276);
nand U47798 (N_47798,N_44813,N_41245);
nor U47799 (N_47799,N_42937,N_42535);
and U47800 (N_47800,N_40595,N_44714);
nor U47801 (N_47801,N_40731,N_42588);
nor U47802 (N_47802,N_41929,N_43289);
xnor U47803 (N_47803,N_40042,N_43274);
xnor U47804 (N_47804,N_44895,N_42914);
nand U47805 (N_47805,N_42198,N_41167);
or U47806 (N_47806,N_40868,N_42602);
xnor U47807 (N_47807,N_42659,N_41774);
nand U47808 (N_47808,N_41219,N_43631);
xor U47809 (N_47809,N_41174,N_40904);
and U47810 (N_47810,N_44237,N_43982);
nand U47811 (N_47811,N_44154,N_40476);
xnor U47812 (N_47812,N_42872,N_41599);
and U47813 (N_47813,N_43092,N_44217);
xor U47814 (N_47814,N_44871,N_40589);
and U47815 (N_47815,N_40432,N_43262);
nor U47816 (N_47816,N_44800,N_40175);
nand U47817 (N_47817,N_40457,N_40657);
or U47818 (N_47818,N_44717,N_43462);
nor U47819 (N_47819,N_43839,N_43247);
xor U47820 (N_47820,N_41500,N_40956);
and U47821 (N_47821,N_43862,N_40483);
or U47822 (N_47822,N_43418,N_41166);
or U47823 (N_47823,N_44265,N_44589);
and U47824 (N_47824,N_41071,N_42564);
nand U47825 (N_47825,N_43834,N_40709);
and U47826 (N_47826,N_42168,N_43579);
nand U47827 (N_47827,N_43580,N_42243);
and U47828 (N_47828,N_43079,N_40535);
xnor U47829 (N_47829,N_43648,N_42696);
nor U47830 (N_47830,N_42533,N_43866);
nor U47831 (N_47831,N_42397,N_40623);
xor U47832 (N_47832,N_40448,N_43890);
nor U47833 (N_47833,N_40154,N_40269);
and U47834 (N_47834,N_43551,N_40758);
xnor U47835 (N_47835,N_42634,N_41409);
and U47836 (N_47836,N_44859,N_42631);
or U47837 (N_47837,N_43450,N_42814);
or U47838 (N_47838,N_40405,N_44010);
xor U47839 (N_47839,N_43779,N_44618);
or U47840 (N_47840,N_41163,N_40301);
or U47841 (N_47841,N_43906,N_41770);
nor U47842 (N_47842,N_41333,N_41916);
xnor U47843 (N_47843,N_43957,N_40216);
nand U47844 (N_47844,N_42500,N_41220);
nand U47845 (N_47845,N_43949,N_41276);
nand U47846 (N_47846,N_43237,N_42886);
or U47847 (N_47847,N_42705,N_40453);
nand U47848 (N_47848,N_40285,N_43326);
and U47849 (N_47849,N_43952,N_42512);
nor U47850 (N_47850,N_43099,N_42371);
nand U47851 (N_47851,N_41481,N_40801);
nand U47852 (N_47852,N_40014,N_43395);
xor U47853 (N_47853,N_44490,N_42189);
nor U47854 (N_47854,N_40501,N_43742);
and U47855 (N_47855,N_41266,N_43493);
xnor U47856 (N_47856,N_41881,N_42560);
and U47857 (N_47857,N_42696,N_40477);
nand U47858 (N_47858,N_42093,N_40548);
and U47859 (N_47859,N_40748,N_44204);
nand U47860 (N_47860,N_43015,N_43581);
nand U47861 (N_47861,N_42752,N_42378);
or U47862 (N_47862,N_43622,N_42002);
nor U47863 (N_47863,N_41634,N_40749);
or U47864 (N_47864,N_42311,N_43700);
nand U47865 (N_47865,N_42044,N_41878);
and U47866 (N_47866,N_44069,N_44435);
xor U47867 (N_47867,N_44476,N_43970);
and U47868 (N_47868,N_40614,N_40551);
and U47869 (N_47869,N_42678,N_42423);
xnor U47870 (N_47870,N_42444,N_41149);
nand U47871 (N_47871,N_40821,N_43940);
or U47872 (N_47872,N_42902,N_41115);
nor U47873 (N_47873,N_42820,N_41205);
or U47874 (N_47874,N_44495,N_43666);
or U47875 (N_47875,N_40472,N_44707);
or U47876 (N_47876,N_42903,N_41728);
or U47877 (N_47877,N_42262,N_41617);
xnor U47878 (N_47878,N_40412,N_44371);
xnor U47879 (N_47879,N_41227,N_43993);
and U47880 (N_47880,N_41633,N_43367);
or U47881 (N_47881,N_40875,N_40605);
nand U47882 (N_47882,N_40845,N_43299);
xnor U47883 (N_47883,N_40827,N_41564);
and U47884 (N_47884,N_42733,N_42405);
nor U47885 (N_47885,N_40836,N_42143);
and U47886 (N_47886,N_41217,N_42149);
or U47887 (N_47887,N_44436,N_41133);
xor U47888 (N_47888,N_44201,N_44098);
and U47889 (N_47889,N_44686,N_44225);
and U47890 (N_47890,N_40381,N_44633);
nand U47891 (N_47891,N_42178,N_41929);
xor U47892 (N_47892,N_40710,N_43538);
and U47893 (N_47893,N_42652,N_43577);
or U47894 (N_47894,N_42952,N_41741);
and U47895 (N_47895,N_43549,N_42966);
or U47896 (N_47896,N_42454,N_44777);
and U47897 (N_47897,N_44478,N_42164);
or U47898 (N_47898,N_44540,N_41064);
nor U47899 (N_47899,N_42564,N_44839);
and U47900 (N_47900,N_43045,N_43412);
xnor U47901 (N_47901,N_44027,N_43965);
nand U47902 (N_47902,N_44998,N_43011);
or U47903 (N_47903,N_40510,N_42976);
and U47904 (N_47904,N_42513,N_41653);
and U47905 (N_47905,N_40229,N_41605);
and U47906 (N_47906,N_43451,N_44240);
or U47907 (N_47907,N_44091,N_40773);
and U47908 (N_47908,N_44178,N_42904);
or U47909 (N_47909,N_41730,N_40650);
nor U47910 (N_47910,N_41716,N_44934);
and U47911 (N_47911,N_44453,N_42991);
or U47912 (N_47912,N_44531,N_44774);
nor U47913 (N_47913,N_42118,N_43004);
nor U47914 (N_47914,N_44481,N_42181);
or U47915 (N_47915,N_44825,N_42711);
and U47916 (N_47916,N_40171,N_44269);
xor U47917 (N_47917,N_40443,N_40816);
or U47918 (N_47918,N_44178,N_44709);
or U47919 (N_47919,N_40150,N_42995);
or U47920 (N_47920,N_43619,N_42540);
nand U47921 (N_47921,N_42443,N_41359);
nand U47922 (N_47922,N_42605,N_42639);
or U47923 (N_47923,N_42995,N_40925);
nor U47924 (N_47924,N_41209,N_42709);
or U47925 (N_47925,N_43469,N_40221);
nor U47926 (N_47926,N_44756,N_40550);
and U47927 (N_47927,N_42634,N_42271);
xor U47928 (N_47928,N_40505,N_44893);
and U47929 (N_47929,N_44497,N_40759);
nor U47930 (N_47930,N_40373,N_41022);
or U47931 (N_47931,N_42815,N_43337);
nand U47932 (N_47932,N_43193,N_43269);
nand U47933 (N_47933,N_41810,N_42289);
and U47934 (N_47934,N_40074,N_43363);
and U47935 (N_47935,N_43299,N_40707);
xor U47936 (N_47936,N_43109,N_41631);
nand U47937 (N_47937,N_43241,N_44936);
nor U47938 (N_47938,N_42210,N_44748);
or U47939 (N_47939,N_40027,N_44283);
nand U47940 (N_47940,N_44087,N_44076);
xnor U47941 (N_47941,N_43368,N_42568);
or U47942 (N_47942,N_43092,N_40689);
nand U47943 (N_47943,N_41733,N_40963);
nand U47944 (N_47944,N_43706,N_40480);
nor U47945 (N_47945,N_41359,N_43033);
or U47946 (N_47946,N_41233,N_43838);
or U47947 (N_47947,N_42223,N_40393);
xor U47948 (N_47948,N_40259,N_40316);
xor U47949 (N_47949,N_41843,N_44316);
xnor U47950 (N_47950,N_40968,N_43388);
and U47951 (N_47951,N_42042,N_40641);
nor U47952 (N_47952,N_43983,N_41395);
and U47953 (N_47953,N_40941,N_41828);
nand U47954 (N_47954,N_44760,N_44768);
and U47955 (N_47955,N_42996,N_40527);
and U47956 (N_47956,N_44684,N_40853);
and U47957 (N_47957,N_42186,N_42042);
or U47958 (N_47958,N_40277,N_44230);
nand U47959 (N_47959,N_42068,N_43894);
nor U47960 (N_47960,N_43954,N_41123);
nor U47961 (N_47961,N_42336,N_43047);
or U47962 (N_47962,N_40885,N_41163);
nand U47963 (N_47963,N_44348,N_42288);
and U47964 (N_47964,N_42987,N_43561);
or U47965 (N_47965,N_40268,N_44399);
or U47966 (N_47966,N_41094,N_42325);
xnor U47967 (N_47967,N_43196,N_42170);
or U47968 (N_47968,N_44600,N_44328);
nor U47969 (N_47969,N_41533,N_41149);
nand U47970 (N_47970,N_43850,N_41266);
nor U47971 (N_47971,N_41888,N_43358);
xnor U47972 (N_47972,N_43798,N_40930);
nor U47973 (N_47973,N_44571,N_43617);
xor U47974 (N_47974,N_41630,N_42261);
xor U47975 (N_47975,N_44196,N_43285);
and U47976 (N_47976,N_44385,N_41049);
or U47977 (N_47977,N_40814,N_42216);
and U47978 (N_47978,N_41283,N_44284);
nand U47979 (N_47979,N_43729,N_40409);
xnor U47980 (N_47980,N_42111,N_40980);
nor U47981 (N_47981,N_42986,N_43860);
or U47982 (N_47982,N_43158,N_42264);
xor U47983 (N_47983,N_41007,N_44451);
or U47984 (N_47984,N_42849,N_41429);
or U47985 (N_47985,N_40470,N_40148);
nor U47986 (N_47986,N_42361,N_40210);
and U47987 (N_47987,N_43502,N_42013);
nand U47988 (N_47988,N_43207,N_41437);
xor U47989 (N_47989,N_43981,N_40882);
nor U47990 (N_47990,N_41274,N_43373);
and U47991 (N_47991,N_40798,N_41239);
nor U47992 (N_47992,N_43990,N_44694);
nor U47993 (N_47993,N_42313,N_41774);
nand U47994 (N_47994,N_41374,N_41885);
xor U47995 (N_47995,N_42272,N_40233);
nand U47996 (N_47996,N_40878,N_44785);
nand U47997 (N_47997,N_43089,N_40177);
nand U47998 (N_47998,N_40588,N_40285);
xnor U47999 (N_47999,N_43239,N_42337);
xor U48000 (N_48000,N_44871,N_42976);
xor U48001 (N_48001,N_43719,N_44540);
nand U48002 (N_48002,N_40280,N_40613);
and U48003 (N_48003,N_44497,N_42748);
and U48004 (N_48004,N_42626,N_44144);
nor U48005 (N_48005,N_40027,N_43995);
and U48006 (N_48006,N_42095,N_42603);
nand U48007 (N_48007,N_42445,N_44004);
nor U48008 (N_48008,N_41630,N_42011);
or U48009 (N_48009,N_44165,N_41869);
or U48010 (N_48010,N_40491,N_40755);
and U48011 (N_48011,N_42237,N_41566);
and U48012 (N_48012,N_42558,N_41736);
nor U48013 (N_48013,N_44435,N_40378);
or U48014 (N_48014,N_42095,N_40742);
nand U48015 (N_48015,N_42971,N_42277);
xnor U48016 (N_48016,N_41294,N_43281);
nor U48017 (N_48017,N_42437,N_42777);
or U48018 (N_48018,N_44662,N_42139);
xor U48019 (N_48019,N_44519,N_42608);
and U48020 (N_48020,N_42101,N_44205);
nand U48021 (N_48021,N_40716,N_44466);
nand U48022 (N_48022,N_41892,N_44231);
xor U48023 (N_48023,N_42859,N_40673);
nor U48024 (N_48024,N_44720,N_41267);
or U48025 (N_48025,N_43463,N_42113);
and U48026 (N_48026,N_43080,N_41713);
nor U48027 (N_48027,N_41341,N_43516);
nand U48028 (N_48028,N_40924,N_44910);
or U48029 (N_48029,N_40674,N_41284);
and U48030 (N_48030,N_44125,N_44496);
and U48031 (N_48031,N_43751,N_40409);
nand U48032 (N_48032,N_41901,N_44539);
xor U48033 (N_48033,N_42406,N_44952);
and U48034 (N_48034,N_44914,N_42938);
or U48035 (N_48035,N_44021,N_44193);
and U48036 (N_48036,N_42892,N_44014);
xnor U48037 (N_48037,N_40013,N_41928);
and U48038 (N_48038,N_43384,N_44573);
and U48039 (N_48039,N_44651,N_42455);
xnor U48040 (N_48040,N_40214,N_44789);
or U48041 (N_48041,N_42690,N_44499);
xor U48042 (N_48042,N_40079,N_43882);
and U48043 (N_48043,N_40265,N_41838);
and U48044 (N_48044,N_43069,N_44471);
nor U48045 (N_48045,N_44687,N_40569);
nor U48046 (N_48046,N_44768,N_41876);
and U48047 (N_48047,N_42549,N_40666);
and U48048 (N_48048,N_44520,N_44813);
xnor U48049 (N_48049,N_43038,N_40121);
nand U48050 (N_48050,N_41976,N_44091);
nor U48051 (N_48051,N_42229,N_44892);
nor U48052 (N_48052,N_40137,N_41416);
nor U48053 (N_48053,N_41849,N_42560);
nor U48054 (N_48054,N_40607,N_40853);
nand U48055 (N_48055,N_41722,N_40583);
nor U48056 (N_48056,N_41736,N_43391);
nand U48057 (N_48057,N_42292,N_44969);
nand U48058 (N_48058,N_41964,N_43902);
nand U48059 (N_48059,N_44622,N_40274);
nand U48060 (N_48060,N_42448,N_42038);
xnor U48061 (N_48061,N_42892,N_40677);
or U48062 (N_48062,N_44010,N_41753);
and U48063 (N_48063,N_41199,N_44562);
or U48064 (N_48064,N_43919,N_44531);
or U48065 (N_48065,N_43615,N_41272);
and U48066 (N_48066,N_44517,N_41698);
or U48067 (N_48067,N_42768,N_40322);
and U48068 (N_48068,N_44964,N_44519);
nor U48069 (N_48069,N_41702,N_40932);
nor U48070 (N_48070,N_42776,N_44738);
and U48071 (N_48071,N_40842,N_40936);
nor U48072 (N_48072,N_42743,N_41090);
nand U48073 (N_48073,N_41037,N_40565);
nor U48074 (N_48074,N_43225,N_44838);
or U48075 (N_48075,N_43017,N_43119);
nand U48076 (N_48076,N_43253,N_42335);
and U48077 (N_48077,N_42660,N_44331);
xnor U48078 (N_48078,N_41940,N_43403);
xnor U48079 (N_48079,N_43025,N_44059);
nand U48080 (N_48080,N_44366,N_42958);
xnor U48081 (N_48081,N_40525,N_43616);
nand U48082 (N_48082,N_41818,N_42526);
and U48083 (N_48083,N_44422,N_40132);
xnor U48084 (N_48084,N_44320,N_40834);
nor U48085 (N_48085,N_42805,N_40934);
nor U48086 (N_48086,N_41391,N_41146);
nand U48087 (N_48087,N_43105,N_41538);
nand U48088 (N_48088,N_44860,N_44564);
nor U48089 (N_48089,N_44605,N_40421);
nand U48090 (N_48090,N_44246,N_44816);
nand U48091 (N_48091,N_40434,N_41992);
xnor U48092 (N_48092,N_43467,N_42749);
and U48093 (N_48093,N_41085,N_43420);
xnor U48094 (N_48094,N_42713,N_40099);
nand U48095 (N_48095,N_42140,N_40595);
or U48096 (N_48096,N_42801,N_41844);
nor U48097 (N_48097,N_41088,N_40150);
nor U48098 (N_48098,N_42089,N_41813);
nor U48099 (N_48099,N_43647,N_42116);
and U48100 (N_48100,N_40594,N_42549);
nand U48101 (N_48101,N_42823,N_42184);
or U48102 (N_48102,N_42167,N_42939);
and U48103 (N_48103,N_42200,N_42405);
and U48104 (N_48104,N_44316,N_42820);
xor U48105 (N_48105,N_41056,N_40337);
xor U48106 (N_48106,N_40033,N_44563);
nand U48107 (N_48107,N_40934,N_41748);
nand U48108 (N_48108,N_40474,N_44820);
and U48109 (N_48109,N_44756,N_42813);
nor U48110 (N_48110,N_40707,N_40376);
nor U48111 (N_48111,N_40103,N_40242);
and U48112 (N_48112,N_40843,N_40701);
nor U48113 (N_48113,N_40371,N_43486);
nor U48114 (N_48114,N_41606,N_41169);
nand U48115 (N_48115,N_44348,N_40560);
nand U48116 (N_48116,N_40590,N_40511);
nand U48117 (N_48117,N_42523,N_43078);
xor U48118 (N_48118,N_40344,N_44812);
nor U48119 (N_48119,N_40723,N_40578);
nand U48120 (N_48120,N_42929,N_43243);
or U48121 (N_48121,N_42222,N_43079);
xnor U48122 (N_48122,N_41507,N_43239);
and U48123 (N_48123,N_41333,N_44164);
nor U48124 (N_48124,N_44089,N_42835);
and U48125 (N_48125,N_44514,N_42316);
or U48126 (N_48126,N_44098,N_42291);
nor U48127 (N_48127,N_42111,N_43479);
and U48128 (N_48128,N_42748,N_43153);
and U48129 (N_48129,N_42160,N_43953);
nand U48130 (N_48130,N_44211,N_43279);
nand U48131 (N_48131,N_42130,N_40005);
nor U48132 (N_48132,N_40533,N_44704);
or U48133 (N_48133,N_43005,N_44958);
and U48134 (N_48134,N_42379,N_44178);
nand U48135 (N_48135,N_43699,N_43975);
nand U48136 (N_48136,N_40417,N_40986);
xnor U48137 (N_48137,N_42348,N_44658);
or U48138 (N_48138,N_43035,N_43120);
and U48139 (N_48139,N_44329,N_43729);
or U48140 (N_48140,N_41523,N_41635);
or U48141 (N_48141,N_42024,N_43993);
nor U48142 (N_48142,N_42973,N_42723);
xnor U48143 (N_48143,N_41547,N_41591);
or U48144 (N_48144,N_44083,N_40269);
or U48145 (N_48145,N_41416,N_43385);
nand U48146 (N_48146,N_40312,N_43692);
or U48147 (N_48147,N_40250,N_43292);
or U48148 (N_48148,N_40732,N_42229);
xor U48149 (N_48149,N_40489,N_42816);
xor U48150 (N_48150,N_44275,N_40399);
xor U48151 (N_48151,N_41566,N_41108);
nand U48152 (N_48152,N_41171,N_40796);
nand U48153 (N_48153,N_40433,N_44791);
nand U48154 (N_48154,N_42847,N_42079);
nor U48155 (N_48155,N_40928,N_44783);
xor U48156 (N_48156,N_44614,N_41859);
nor U48157 (N_48157,N_41963,N_44209);
nor U48158 (N_48158,N_40529,N_43176);
and U48159 (N_48159,N_40215,N_44941);
nor U48160 (N_48160,N_41841,N_44731);
nor U48161 (N_48161,N_44369,N_41507);
or U48162 (N_48162,N_42872,N_44401);
or U48163 (N_48163,N_43232,N_44179);
or U48164 (N_48164,N_43385,N_44558);
nand U48165 (N_48165,N_41269,N_44485);
xor U48166 (N_48166,N_42077,N_44222);
nor U48167 (N_48167,N_44535,N_42988);
xnor U48168 (N_48168,N_41548,N_43730);
and U48169 (N_48169,N_43488,N_40575);
nand U48170 (N_48170,N_43451,N_40002);
or U48171 (N_48171,N_42502,N_40192);
nor U48172 (N_48172,N_43704,N_41807);
xnor U48173 (N_48173,N_42240,N_44058);
or U48174 (N_48174,N_42359,N_43001);
and U48175 (N_48175,N_44974,N_42986);
or U48176 (N_48176,N_43580,N_42801);
and U48177 (N_48177,N_42346,N_42405);
xnor U48178 (N_48178,N_44969,N_43481);
nand U48179 (N_48179,N_41990,N_41796);
nand U48180 (N_48180,N_42808,N_40735);
nand U48181 (N_48181,N_42894,N_42497);
nand U48182 (N_48182,N_44518,N_41815);
nor U48183 (N_48183,N_44315,N_44198);
nor U48184 (N_48184,N_41634,N_43696);
nand U48185 (N_48185,N_44142,N_42023);
nand U48186 (N_48186,N_41815,N_41760);
or U48187 (N_48187,N_44172,N_41897);
nor U48188 (N_48188,N_44046,N_42175);
and U48189 (N_48189,N_41660,N_41563);
xor U48190 (N_48190,N_42273,N_41368);
nor U48191 (N_48191,N_41354,N_44319);
xor U48192 (N_48192,N_44300,N_40970);
nor U48193 (N_48193,N_41304,N_41505);
xnor U48194 (N_48194,N_40388,N_44739);
nor U48195 (N_48195,N_44653,N_44022);
xnor U48196 (N_48196,N_41876,N_43911);
or U48197 (N_48197,N_41416,N_44074);
or U48198 (N_48198,N_43886,N_40527);
or U48199 (N_48199,N_42108,N_40236);
nor U48200 (N_48200,N_42878,N_43695);
or U48201 (N_48201,N_40505,N_41100);
or U48202 (N_48202,N_42262,N_43922);
xnor U48203 (N_48203,N_41759,N_44174);
and U48204 (N_48204,N_41938,N_44793);
nand U48205 (N_48205,N_42681,N_41246);
xnor U48206 (N_48206,N_41612,N_44879);
nand U48207 (N_48207,N_44426,N_44981);
nand U48208 (N_48208,N_42933,N_41441);
and U48209 (N_48209,N_40473,N_43446);
nand U48210 (N_48210,N_40951,N_43088);
nand U48211 (N_48211,N_44353,N_41990);
nor U48212 (N_48212,N_44403,N_40266);
nand U48213 (N_48213,N_41836,N_44502);
xor U48214 (N_48214,N_40454,N_44347);
or U48215 (N_48215,N_41382,N_43654);
xor U48216 (N_48216,N_44734,N_42815);
nand U48217 (N_48217,N_44563,N_41473);
and U48218 (N_48218,N_43930,N_43929);
xor U48219 (N_48219,N_42863,N_42228);
xor U48220 (N_48220,N_44361,N_43302);
and U48221 (N_48221,N_40696,N_42826);
xor U48222 (N_48222,N_44235,N_44408);
nand U48223 (N_48223,N_42159,N_43770);
and U48224 (N_48224,N_41851,N_44064);
nor U48225 (N_48225,N_41713,N_41016);
xnor U48226 (N_48226,N_40226,N_40942);
xor U48227 (N_48227,N_43331,N_43547);
and U48228 (N_48228,N_43190,N_40107);
xor U48229 (N_48229,N_44178,N_40314);
and U48230 (N_48230,N_41154,N_40896);
and U48231 (N_48231,N_43882,N_40197);
or U48232 (N_48232,N_40372,N_41411);
nand U48233 (N_48233,N_40899,N_41886);
nand U48234 (N_48234,N_43184,N_41489);
and U48235 (N_48235,N_42221,N_42791);
nand U48236 (N_48236,N_43339,N_42641);
nand U48237 (N_48237,N_43864,N_44429);
or U48238 (N_48238,N_41757,N_42133);
nor U48239 (N_48239,N_42610,N_40113);
and U48240 (N_48240,N_42111,N_42114);
nand U48241 (N_48241,N_44520,N_40507);
and U48242 (N_48242,N_42222,N_44882);
nor U48243 (N_48243,N_40897,N_42875);
xor U48244 (N_48244,N_43190,N_44219);
nor U48245 (N_48245,N_43326,N_40110);
xor U48246 (N_48246,N_41061,N_42758);
nor U48247 (N_48247,N_41077,N_41030);
and U48248 (N_48248,N_43835,N_43423);
nor U48249 (N_48249,N_40462,N_42377);
xnor U48250 (N_48250,N_40796,N_43369);
or U48251 (N_48251,N_42381,N_40148);
or U48252 (N_48252,N_40215,N_41152);
nor U48253 (N_48253,N_42217,N_43193);
xor U48254 (N_48254,N_42549,N_40551);
or U48255 (N_48255,N_42579,N_42905);
and U48256 (N_48256,N_40016,N_44505);
nor U48257 (N_48257,N_44592,N_44052);
xor U48258 (N_48258,N_40319,N_43937);
nand U48259 (N_48259,N_41958,N_43575);
nor U48260 (N_48260,N_44416,N_42370);
and U48261 (N_48261,N_41149,N_41008);
or U48262 (N_48262,N_44966,N_41036);
nor U48263 (N_48263,N_40393,N_41635);
nand U48264 (N_48264,N_44359,N_41649);
nand U48265 (N_48265,N_44063,N_44954);
xor U48266 (N_48266,N_43619,N_42561);
and U48267 (N_48267,N_41818,N_42063);
nand U48268 (N_48268,N_43905,N_43257);
or U48269 (N_48269,N_40206,N_40977);
or U48270 (N_48270,N_43140,N_40479);
or U48271 (N_48271,N_41532,N_43173);
xor U48272 (N_48272,N_44413,N_44419);
nor U48273 (N_48273,N_44704,N_42345);
nor U48274 (N_48274,N_41824,N_40538);
nand U48275 (N_48275,N_41559,N_44375);
xnor U48276 (N_48276,N_41486,N_44237);
nor U48277 (N_48277,N_40879,N_44388);
and U48278 (N_48278,N_40083,N_41272);
nand U48279 (N_48279,N_43415,N_41155);
and U48280 (N_48280,N_43833,N_42029);
or U48281 (N_48281,N_44192,N_42393);
nand U48282 (N_48282,N_41662,N_43559);
and U48283 (N_48283,N_44401,N_43888);
and U48284 (N_48284,N_43346,N_41717);
and U48285 (N_48285,N_40121,N_42178);
or U48286 (N_48286,N_41360,N_44585);
and U48287 (N_48287,N_42121,N_41479);
nand U48288 (N_48288,N_41038,N_41158);
xor U48289 (N_48289,N_42121,N_41219);
and U48290 (N_48290,N_43740,N_40265);
or U48291 (N_48291,N_40601,N_40804);
nor U48292 (N_48292,N_42799,N_40158);
xnor U48293 (N_48293,N_41122,N_40846);
or U48294 (N_48294,N_44142,N_44424);
nor U48295 (N_48295,N_42054,N_43955);
nand U48296 (N_48296,N_41012,N_43416);
nor U48297 (N_48297,N_41064,N_43249);
or U48298 (N_48298,N_43140,N_41924);
nor U48299 (N_48299,N_41226,N_40702);
nor U48300 (N_48300,N_44525,N_44688);
xnor U48301 (N_48301,N_43525,N_40387);
nand U48302 (N_48302,N_40965,N_40293);
nand U48303 (N_48303,N_43640,N_44702);
xnor U48304 (N_48304,N_42760,N_44281);
and U48305 (N_48305,N_44085,N_41185);
nor U48306 (N_48306,N_40416,N_42912);
nand U48307 (N_48307,N_40915,N_42464);
nand U48308 (N_48308,N_43128,N_43724);
or U48309 (N_48309,N_44369,N_42578);
nand U48310 (N_48310,N_42521,N_41097);
or U48311 (N_48311,N_42396,N_41480);
and U48312 (N_48312,N_44938,N_41941);
and U48313 (N_48313,N_40414,N_42329);
and U48314 (N_48314,N_40265,N_42140);
xor U48315 (N_48315,N_42939,N_41994);
nand U48316 (N_48316,N_42039,N_44409);
and U48317 (N_48317,N_40868,N_44160);
or U48318 (N_48318,N_40567,N_41772);
nor U48319 (N_48319,N_43404,N_44290);
nor U48320 (N_48320,N_44851,N_44850);
and U48321 (N_48321,N_42679,N_44810);
or U48322 (N_48322,N_41553,N_41628);
nor U48323 (N_48323,N_40317,N_41099);
and U48324 (N_48324,N_44696,N_40996);
and U48325 (N_48325,N_40386,N_41471);
or U48326 (N_48326,N_40149,N_41751);
xnor U48327 (N_48327,N_41533,N_41785);
or U48328 (N_48328,N_41732,N_42066);
nand U48329 (N_48329,N_43445,N_42537);
nor U48330 (N_48330,N_43955,N_43511);
xnor U48331 (N_48331,N_42610,N_41667);
or U48332 (N_48332,N_44626,N_44684);
or U48333 (N_48333,N_44216,N_44882);
or U48334 (N_48334,N_42733,N_41959);
nor U48335 (N_48335,N_40800,N_41039);
and U48336 (N_48336,N_42241,N_44965);
or U48337 (N_48337,N_40481,N_40125);
or U48338 (N_48338,N_41805,N_44383);
and U48339 (N_48339,N_41384,N_42545);
or U48340 (N_48340,N_42697,N_40443);
xnor U48341 (N_48341,N_43769,N_41651);
nand U48342 (N_48342,N_44814,N_42529);
or U48343 (N_48343,N_44231,N_44406);
and U48344 (N_48344,N_43092,N_43388);
xor U48345 (N_48345,N_44587,N_41593);
or U48346 (N_48346,N_42344,N_44388);
xnor U48347 (N_48347,N_40293,N_41614);
or U48348 (N_48348,N_44109,N_43567);
nand U48349 (N_48349,N_43229,N_43929);
nor U48350 (N_48350,N_44930,N_42153);
nor U48351 (N_48351,N_42211,N_42888);
xor U48352 (N_48352,N_43526,N_43639);
xor U48353 (N_48353,N_42630,N_44438);
or U48354 (N_48354,N_43844,N_44580);
xnor U48355 (N_48355,N_42544,N_42140);
and U48356 (N_48356,N_43885,N_42940);
xnor U48357 (N_48357,N_42633,N_42043);
or U48358 (N_48358,N_43629,N_43522);
nor U48359 (N_48359,N_44725,N_43012);
nor U48360 (N_48360,N_42661,N_40597);
and U48361 (N_48361,N_42264,N_43209);
and U48362 (N_48362,N_42208,N_41020);
or U48363 (N_48363,N_42793,N_43916);
nor U48364 (N_48364,N_43121,N_40444);
and U48365 (N_48365,N_43340,N_42355);
or U48366 (N_48366,N_44784,N_44938);
and U48367 (N_48367,N_43122,N_40633);
or U48368 (N_48368,N_40290,N_41191);
nor U48369 (N_48369,N_43260,N_42182);
and U48370 (N_48370,N_43127,N_44037);
and U48371 (N_48371,N_42084,N_44429);
nor U48372 (N_48372,N_43796,N_41980);
or U48373 (N_48373,N_41390,N_41304);
nor U48374 (N_48374,N_44162,N_40663);
nor U48375 (N_48375,N_43524,N_44336);
nor U48376 (N_48376,N_42816,N_43064);
xor U48377 (N_48377,N_43793,N_42049);
or U48378 (N_48378,N_42870,N_44507);
xor U48379 (N_48379,N_42295,N_42563);
and U48380 (N_48380,N_40860,N_43902);
xnor U48381 (N_48381,N_40125,N_43645);
nor U48382 (N_48382,N_40145,N_43821);
xnor U48383 (N_48383,N_40154,N_41321);
and U48384 (N_48384,N_43147,N_40598);
or U48385 (N_48385,N_41816,N_41520);
and U48386 (N_48386,N_41555,N_44028);
and U48387 (N_48387,N_43944,N_41434);
nand U48388 (N_48388,N_40896,N_43949);
or U48389 (N_48389,N_41048,N_42023);
nor U48390 (N_48390,N_41450,N_44878);
nand U48391 (N_48391,N_44668,N_43518);
nor U48392 (N_48392,N_42264,N_42746);
nand U48393 (N_48393,N_41318,N_41296);
or U48394 (N_48394,N_43515,N_42671);
nand U48395 (N_48395,N_42490,N_43532);
and U48396 (N_48396,N_40075,N_41558);
and U48397 (N_48397,N_41752,N_41530);
nand U48398 (N_48398,N_43077,N_44178);
nor U48399 (N_48399,N_42806,N_43900);
xor U48400 (N_48400,N_44387,N_40649);
nand U48401 (N_48401,N_42492,N_41752);
xnor U48402 (N_48402,N_41107,N_43332);
nand U48403 (N_48403,N_44595,N_41254);
and U48404 (N_48404,N_43248,N_43727);
nand U48405 (N_48405,N_40792,N_44429);
nand U48406 (N_48406,N_43919,N_43042);
and U48407 (N_48407,N_42350,N_44625);
and U48408 (N_48408,N_42692,N_40584);
and U48409 (N_48409,N_40225,N_42541);
xnor U48410 (N_48410,N_40301,N_44635);
nor U48411 (N_48411,N_41727,N_44230);
or U48412 (N_48412,N_40863,N_41709);
or U48413 (N_48413,N_44013,N_42515);
xnor U48414 (N_48414,N_44566,N_44437);
nand U48415 (N_48415,N_44168,N_43215);
xor U48416 (N_48416,N_44843,N_40480);
nor U48417 (N_48417,N_44499,N_41837);
xor U48418 (N_48418,N_41945,N_44335);
and U48419 (N_48419,N_40203,N_40043);
nor U48420 (N_48420,N_44972,N_43923);
and U48421 (N_48421,N_40850,N_42571);
xor U48422 (N_48422,N_42075,N_42375);
or U48423 (N_48423,N_43661,N_43230);
and U48424 (N_48424,N_41922,N_43337);
xor U48425 (N_48425,N_44275,N_40597);
nor U48426 (N_48426,N_43620,N_43919);
nand U48427 (N_48427,N_43450,N_40760);
xnor U48428 (N_48428,N_43018,N_40410);
or U48429 (N_48429,N_44983,N_40217);
xor U48430 (N_48430,N_42049,N_42710);
and U48431 (N_48431,N_42051,N_44967);
xnor U48432 (N_48432,N_44248,N_41231);
nor U48433 (N_48433,N_43296,N_43553);
nand U48434 (N_48434,N_44428,N_43137);
and U48435 (N_48435,N_42045,N_40947);
and U48436 (N_48436,N_41302,N_40670);
nor U48437 (N_48437,N_43491,N_41756);
or U48438 (N_48438,N_41490,N_40533);
nand U48439 (N_48439,N_42026,N_43768);
or U48440 (N_48440,N_41507,N_42670);
and U48441 (N_48441,N_42458,N_41036);
nor U48442 (N_48442,N_42376,N_44685);
nor U48443 (N_48443,N_44398,N_43934);
nor U48444 (N_48444,N_41826,N_43691);
xor U48445 (N_48445,N_43184,N_41425);
and U48446 (N_48446,N_41092,N_43427);
nand U48447 (N_48447,N_41532,N_43812);
xnor U48448 (N_48448,N_43426,N_41765);
and U48449 (N_48449,N_44606,N_43878);
nand U48450 (N_48450,N_42423,N_43569);
nand U48451 (N_48451,N_41604,N_40128);
xor U48452 (N_48452,N_42395,N_44259);
nor U48453 (N_48453,N_44437,N_44225);
nor U48454 (N_48454,N_43802,N_41894);
and U48455 (N_48455,N_44178,N_41897);
xnor U48456 (N_48456,N_40550,N_40722);
nor U48457 (N_48457,N_41685,N_40579);
nor U48458 (N_48458,N_43210,N_43471);
and U48459 (N_48459,N_42060,N_44880);
nor U48460 (N_48460,N_40684,N_41366);
or U48461 (N_48461,N_41193,N_44601);
or U48462 (N_48462,N_44591,N_40358);
nand U48463 (N_48463,N_40669,N_41226);
xor U48464 (N_48464,N_41153,N_41805);
nor U48465 (N_48465,N_41972,N_43513);
xnor U48466 (N_48466,N_44595,N_41548);
xnor U48467 (N_48467,N_42036,N_42923);
nor U48468 (N_48468,N_44874,N_44166);
nand U48469 (N_48469,N_41616,N_41150);
nand U48470 (N_48470,N_42302,N_40634);
nand U48471 (N_48471,N_41920,N_40575);
or U48472 (N_48472,N_41963,N_41475);
xnor U48473 (N_48473,N_43598,N_40850);
and U48474 (N_48474,N_42393,N_43236);
xor U48475 (N_48475,N_44592,N_42462);
and U48476 (N_48476,N_43558,N_40965);
or U48477 (N_48477,N_44795,N_40348);
or U48478 (N_48478,N_42459,N_42128);
or U48479 (N_48479,N_40237,N_43396);
or U48480 (N_48480,N_42958,N_40834);
nand U48481 (N_48481,N_43644,N_43252);
nand U48482 (N_48482,N_41098,N_42808);
or U48483 (N_48483,N_44429,N_42063);
or U48484 (N_48484,N_43627,N_40859);
and U48485 (N_48485,N_40396,N_43237);
nand U48486 (N_48486,N_41992,N_41432);
and U48487 (N_48487,N_42315,N_42545);
nor U48488 (N_48488,N_44553,N_40440);
nand U48489 (N_48489,N_43935,N_41461);
or U48490 (N_48490,N_41129,N_41404);
or U48491 (N_48491,N_44056,N_41184);
nand U48492 (N_48492,N_44658,N_40475);
or U48493 (N_48493,N_42044,N_44731);
xor U48494 (N_48494,N_44913,N_42622);
nand U48495 (N_48495,N_42993,N_41645);
xnor U48496 (N_48496,N_44457,N_40347);
xnor U48497 (N_48497,N_42828,N_43164);
xnor U48498 (N_48498,N_43473,N_40579);
nor U48499 (N_48499,N_41482,N_42405);
or U48500 (N_48500,N_41014,N_41837);
xnor U48501 (N_48501,N_44550,N_43710);
and U48502 (N_48502,N_41122,N_42925);
xnor U48503 (N_48503,N_42514,N_40660);
or U48504 (N_48504,N_44342,N_42965);
and U48505 (N_48505,N_44601,N_40728);
xor U48506 (N_48506,N_40672,N_43202);
nand U48507 (N_48507,N_42271,N_41787);
nand U48508 (N_48508,N_42994,N_41104);
xor U48509 (N_48509,N_43249,N_44609);
nor U48510 (N_48510,N_43611,N_44957);
and U48511 (N_48511,N_42568,N_42457);
nor U48512 (N_48512,N_40203,N_40416);
nand U48513 (N_48513,N_42040,N_40038);
and U48514 (N_48514,N_43625,N_42029);
or U48515 (N_48515,N_42384,N_42037);
xnor U48516 (N_48516,N_44196,N_41336);
or U48517 (N_48517,N_42249,N_44131);
or U48518 (N_48518,N_41400,N_40586);
nor U48519 (N_48519,N_42279,N_44987);
xnor U48520 (N_48520,N_42083,N_41747);
and U48521 (N_48521,N_41840,N_43217);
nand U48522 (N_48522,N_40601,N_43940);
and U48523 (N_48523,N_42640,N_41903);
or U48524 (N_48524,N_44323,N_41645);
or U48525 (N_48525,N_42969,N_44239);
and U48526 (N_48526,N_40472,N_43840);
nand U48527 (N_48527,N_41007,N_42481);
nor U48528 (N_48528,N_40715,N_44321);
and U48529 (N_48529,N_41911,N_40818);
nand U48530 (N_48530,N_42915,N_41345);
nand U48531 (N_48531,N_44060,N_42720);
nand U48532 (N_48532,N_43527,N_43038);
nand U48533 (N_48533,N_40286,N_42177);
nor U48534 (N_48534,N_40589,N_40619);
or U48535 (N_48535,N_41057,N_40905);
and U48536 (N_48536,N_43402,N_44538);
xnor U48537 (N_48537,N_42623,N_41560);
xor U48538 (N_48538,N_43426,N_41948);
or U48539 (N_48539,N_40811,N_40391);
nand U48540 (N_48540,N_43948,N_41723);
xor U48541 (N_48541,N_41601,N_41002);
and U48542 (N_48542,N_42206,N_44051);
xnor U48543 (N_48543,N_40618,N_42513);
nor U48544 (N_48544,N_42681,N_42004);
or U48545 (N_48545,N_42742,N_42416);
nand U48546 (N_48546,N_42120,N_42275);
or U48547 (N_48547,N_41548,N_42222);
and U48548 (N_48548,N_43006,N_44492);
and U48549 (N_48549,N_41889,N_42170);
nor U48550 (N_48550,N_41748,N_42462);
and U48551 (N_48551,N_44993,N_41049);
nor U48552 (N_48552,N_41018,N_40602);
nand U48553 (N_48553,N_44400,N_41649);
nand U48554 (N_48554,N_43419,N_40933);
nor U48555 (N_48555,N_41024,N_41221);
nand U48556 (N_48556,N_44198,N_42165);
nor U48557 (N_48557,N_44250,N_42815);
and U48558 (N_48558,N_40907,N_41689);
and U48559 (N_48559,N_40195,N_44855);
nand U48560 (N_48560,N_41247,N_43882);
nor U48561 (N_48561,N_43054,N_40756);
and U48562 (N_48562,N_44225,N_40806);
nor U48563 (N_48563,N_43319,N_42057);
xor U48564 (N_48564,N_41272,N_40303);
or U48565 (N_48565,N_41011,N_43729);
and U48566 (N_48566,N_41262,N_41598);
or U48567 (N_48567,N_41892,N_44048);
or U48568 (N_48568,N_41844,N_42164);
nor U48569 (N_48569,N_44987,N_44935);
and U48570 (N_48570,N_42090,N_41893);
nand U48571 (N_48571,N_44066,N_41889);
and U48572 (N_48572,N_44158,N_44442);
nand U48573 (N_48573,N_44470,N_42519);
nor U48574 (N_48574,N_43580,N_40943);
nand U48575 (N_48575,N_42702,N_40669);
or U48576 (N_48576,N_42387,N_42473);
and U48577 (N_48577,N_44975,N_41808);
xnor U48578 (N_48578,N_42793,N_40333);
and U48579 (N_48579,N_44602,N_43190);
and U48580 (N_48580,N_43937,N_44231);
nand U48581 (N_48581,N_44902,N_40711);
and U48582 (N_48582,N_44206,N_42337);
nand U48583 (N_48583,N_44780,N_40569);
or U48584 (N_48584,N_41825,N_41195);
nor U48585 (N_48585,N_41817,N_43841);
xor U48586 (N_48586,N_40128,N_42254);
nor U48587 (N_48587,N_41602,N_43609);
nor U48588 (N_48588,N_43616,N_40943);
nor U48589 (N_48589,N_44797,N_43073);
nor U48590 (N_48590,N_41625,N_42470);
or U48591 (N_48591,N_43162,N_44494);
nor U48592 (N_48592,N_43810,N_42882);
and U48593 (N_48593,N_41177,N_42464);
nor U48594 (N_48594,N_42020,N_43293);
or U48595 (N_48595,N_43732,N_44355);
or U48596 (N_48596,N_42090,N_44812);
nand U48597 (N_48597,N_41070,N_43460);
xor U48598 (N_48598,N_44400,N_40219);
or U48599 (N_48599,N_42123,N_42668);
nand U48600 (N_48600,N_41354,N_42926);
nor U48601 (N_48601,N_42256,N_44117);
xnor U48602 (N_48602,N_41530,N_42286);
or U48603 (N_48603,N_41751,N_42473);
nand U48604 (N_48604,N_44182,N_42793);
or U48605 (N_48605,N_42420,N_43738);
nor U48606 (N_48606,N_44418,N_40879);
or U48607 (N_48607,N_42697,N_43444);
nor U48608 (N_48608,N_41572,N_42568);
nor U48609 (N_48609,N_42246,N_41700);
nand U48610 (N_48610,N_44363,N_42170);
or U48611 (N_48611,N_40438,N_44077);
nor U48612 (N_48612,N_40539,N_40361);
nand U48613 (N_48613,N_43128,N_41253);
nor U48614 (N_48614,N_40585,N_41841);
nand U48615 (N_48615,N_41125,N_43718);
or U48616 (N_48616,N_40760,N_43907);
nand U48617 (N_48617,N_40536,N_44540);
nand U48618 (N_48618,N_43554,N_43456);
nor U48619 (N_48619,N_42156,N_43483);
nor U48620 (N_48620,N_43765,N_42308);
nand U48621 (N_48621,N_40741,N_44100);
nor U48622 (N_48622,N_43292,N_41333);
nor U48623 (N_48623,N_42715,N_43368);
or U48624 (N_48624,N_42253,N_41809);
or U48625 (N_48625,N_44386,N_43149);
and U48626 (N_48626,N_44458,N_41527);
nor U48627 (N_48627,N_42690,N_40443);
xnor U48628 (N_48628,N_42189,N_41061);
nor U48629 (N_48629,N_43911,N_42375);
nor U48630 (N_48630,N_43975,N_41398);
and U48631 (N_48631,N_41214,N_44744);
and U48632 (N_48632,N_43592,N_41905);
nor U48633 (N_48633,N_40675,N_40603);
or U48634 (N_48634,N_41638,N_42074);
or U48635 (N_48635,N_44015,N_43124);
nand U48636 (N_48636,N_43191,N_42819);
nor U48637 (N_48637,N_44551,N_40146);
nor U48638 (N_48638,N_41786,N_43168);
and U48639 (N_48639,N_41359,N_42377);
nor U48640 (N_48640,N_40190,N_43717);
xor U48641 (N_48641,N_42452,N_40883);
nor U48642 (N_48642,N_43942,N_43553);
nor U48643 (N_48643,N_40496,N_44575);
nand U48644 (N_48644,N_40481,N_40665);
or U48645 (N_48645,N_43267,N_44890);
and U48646 (N_48646,N_44314,N_43552);
xor U48647 (N_48647,N_44604,N_43251);
or U48648 (N_48648,N_44467,N_44657);
nor U48649 (N_48649,N_43718,N_42973);
nor U48650 (N_48650,N_41918,N_41593);
or U48651 (N_48651,N_40680,N_41986);
and U48652 (N_48652,N_40612,N_41802);
nor U48653 (N_48653,N_41021,N_40994);
and U48654 (N_48654,N_43690,N_40684);
nor U48655 (N_48655,N_44359,N_40004);
xnor U48656 (N_48656,N_41139,N_41030);
and U48657 (N_48657,N_43352,N_41435);
nand U48658 (N_48658,N_40235,N_43000);
nor U48659 (N_48659,N_44471,N_40749);
or U48660 (N_48660,N_44243,N_43417);
and U48661 (N_48661,N_43501,N_42142);
and U48662 (N_48662,N_41068,N_41449);
and U48663 (N_48663,N_44695,N_44065);
nor U48664 (N_48664,N_44621,N_44701);
nor U48665 (N_48665,N_41823,N_41766);
xnor U48666 (N_48666,N_40365,N_41387);
xnor U48667 (N_48667,N_42733,N_42926);
nor U48668 (N_48668,N_40616,N_43096);
xor U48669 (N_48669,N_43011,N_40907);
nand U48670 (N_48670,N_40126,N_43889);
or U48671 (N_48671,N_43383,N_43082);
or U48672 (N_48672,N_43256,N_41798);
nor U48673 (N_48673,N_40134,N_41756);
and U48674 (N_48674,N_40771,N_43864);
xnor U48675 (N_48675,N_41577,N_44803);
nand U48676 (N_48676,N_42476,N_40536);
or U48677 (N_48677,N_40366,N_41583);
xor U48678 (N_48678,N_42103,N_40186);
xor U48679 (N_48679,N_44470,N_42172);
nand U48680 (N_48680,N_44950,N_44467);
or U48681 (N_48681,N_41634,N_40083);
xor U48682 (N_48682,N_42881,N_43934);
nand U48683 (N_48683,N_41279,N_42132);
xor U48684 (N_48684,N_44739,N_42754);
or U48685 (N_48685,N_43653,N_43060);
or U48686 (N_48686,N_41875,N_40403);
nand U48687 (N_48687,N_43014,N_41545);
and U48688 (N_48688,N_40943,N_41234);
or U48689 (N_48689,N_44273,N_43095);
nor U48690 (N_48690,N_43958,N_41312);
nand U48691 (N_48691,N_41333,N_44431);
or U48692 (N_48692,N_41364,N_44423);
xor U48693 (N_48693,N_42007,N_40716);
nand U48694 (N_48694,N_42918,N_44858);
or U48695 (N_48695,N_40408,N_40554);
xor U48696 (N_48696,N_44594,N_44117);
nand U48697 (N_48697,N_43020,N_40014);
xor U48698 (N_48698,N_40304,N_40905);
xor U48699 (N_48699,N_44849,N_40028);
or U48700 (N_48700,N_40439,N_42633);
and U48701 (N_48701,N_44441,N_44706);
nand U48702 (N_48702,N_42498,N_42679);
and U48703 (N_48703,N_41623,N_40024);
nor U48704 (N_48704,N_41429,N_43213);
xor U48705 (N_48705,N_43084,N_42617);
xor U48706 (N_48706,N_44299,N_42102);
and U48707 (N_48707,N_44308,N_44312);
or U48708 (N_48708,N_42230,N_40437);
or U48709 (N_48709,N_44048,N_41553);
nor U48710 (N_48710,N_40806,N_41195);
nor U48711 (N_48711,N_41345,N_43391);
xor U48712 (N_48712,N_41995,N_41308);
nor U48713 (N_48713,N_40840,N_43285);
or U48714 (N_48714,N_41678,N_41937);
and U48715 (N_48715,N_40844,N_43463);
nand U48716 (N_48716,N_43740,N_40735);
or U48717 (N_48717,N_43367,N_42868);
nand U48718 (N_48718,N_43013,N_43745);
nand U48719 (N_48719,N_44825,N_44857);
nor U48720 (N_48720,N_41546,N_42390);
nor U48721 (N_48721,N_40850,N_43760);
and U48722 (N_48722,N_44390,N_40250);
and U48723 (N_48723,N_44545,N_44084);
and U48724 (N_48724,N_44986,N_44719);
and U48725 (N_48725,N_40908,N_43056);
nand U48726 (N_48726,N_40458,N_42340);
or U48727 (N_48727,N_42651,N_42467);
xnor U48728 (N_48728,N_40635,N_42049);
xnor U48729 (N_48729,N_44661,N_40831);
nor U48730 (N_48730,N_42002,N_40832);
or U48731 (N_48731,N_43304,N_44817);
or U48732 (N_48732,N_41344,N_44600);
or U48733 (N_48733,N_44942,N_41360);
or U48734 (N_48734,N_44657,N_42414);
nor U48735 (N_48735,N_40218,N_40366);
nand U48736 (N_48736,N_42674,N_43955);
xor U48737 (N_48737,N_41181,N_42847);
nor U48738 (N_48738,N_42446,N_44799);
xor U48739 (N_48739,N_43802,N_42434);
or U48740 (N_48740,N_44380,N_41222);
nand U48741 (N_48741,N_40820,N_44753);
nor U48742 (N_48742,N_43828,N_44401);
xor U48743 (N_48743,N_42110,N_40736);
nand U48744 (N_48744,N_42451,N_43490);
and U48745 (N_48745,N_42214,N_44952);
xnor U48746 (N_48746,N_44884,N_40821);
nand U48747 (N_48747,N_40788,N_42449);
or U48748 (N_48748,N_42619,N_42659);
and U48749 (N_48749,N_40316,N_41384);
nor U48750 (N_48750,N_41067,N_40864);
and U48751 (N_48751,N_44241,N_41550);
or U48752 (N_48752,N_41143,N_40395);
and U48753 (N_48753,N_40246,N_44525);
and U48754 (N_48754,N_40332,N_43574);
or U48755 (N_48755,N_42614,N_44688);
xor U48756 (N_48756,N_43763,N_41401);
nor U48757 (N_48757,N_44160,N_40898);
nor U48758 (N_48758,N_44856,N_44805);
nand U48759 (N_48759,N_42966,N_43019);
xor U48760 (N_48760,N_42243,N_44446);
and U48761 (N_48761,N_42535,N_41553);
nand U48762 (N_48762,N_41168,N_43492);
or U48763 (N_48763,N_40799,N_43695);
xor U48764 (N_48764,N_41976,N_40325);
nand U48765 (N_48765,N_43671,N_42475);
and U48766 (N_48766,N_43623,N_41441);
and U48767 (N_48767,N_40244,N_43870);
xor U48768 (N_48768,N_42058,N_41091);
nand U48769 (N_48769,N_43206,N_42517);
nor U48770 (N_48770,N_44253,N_41035);
and U48771 (N_48771,N_43759,N_43134);
or U48772 (N_48772,N_43722,N_42903);
nand U48773 (N_48773,N_42451,N_41307);
xnor U48774 (N_48774,N_42231,N_43772);
nor U48775 (N_48775,N_44812,N_42335);
nor U48776 (N_48776,N_44636,N_43870);
nor U48777 (N_48777,N_43401,N_42341);
and U48778 (N_48778,N_42219,N_43740);
nor U48779 (N_48779,N_43106,N_42665);
or U48780 (N_48780,N_44628,N_42406);
or U48781 (N_48781,N_43465,N_44733);
nand U48782 (N_48782,N_41894,N_42200);
and U48783 (N_48783,N_44318,N_44534);
nand U48784 (N_48784,N_42730,N_42842);
nand U48785 (N_48785,N_40699,N_43302);
or U48786 (N_48786,N_43813,N_40253);
and U48787 (N_48787,N_44732,N_40692);
or U48788 (N_48788,N_40645,N_42244);
xor U48789 (N_48789,N_42383,N_40013);
nand U48790 (N_48790,N_40352,N_41562);
and U48791 (N_48791,N_40567,N_43538);
and U48792 (N_48792,N_41669,N_42456);
nor U48793 (N_48793,N_43975,N_41170);
and U48794 (N_48794,N_41719,N_43212);
and U48795 (N_48795,N_41805,N_41078);
xnor U48796 (N_48796,N_42044,N_42085);
or U48797 (N_48797,N_42100,N_41645);
and U48798 (N_48798,N_44882,N_41593);
nand U48799 (N_48799,N_40575,N_43821);
nand U48800 (N_48800,N_44187,N_43520);
xnor U48801 (N_48801,N_44023,N_43738);
nand U48802 (N_48802,N_41653,N_40462);
or U48803 (N_48803,N_41807,N_43524);
xor U48804 (N_48804,N_40751,N_40878);
nor U48805 (N_48805,N_44668,N_42646);
and U48806 (N_48806,N_44364,N_43986);
xor U48807 (N_48807,N_42768,N_42665);
nor U48808 (N_48808,N_40148,N_41538);
xor U48809 (N_48809,N_44274,N_42791);
nand U48810 (N_48810,N_44174,N_43076);
nand U48811 (N_48811,N_42262,N_42066);
xnor U48812 (N_48812,N_43466,N_44543);
nand U48813 (N_48813,N_44939,N_41697);
or U48814 (N_48814,N_41407,N_43756);
xnor U48815 (N_48815,N_41879,N_42999);
xnor U48816 (N_48816,N_43985,N_41928);
nor U48817 (N_48817,N_43109,N_42954);
xnor U48818 (N_48818,N_42784,N_41991);
nor U48819 (N_48819,N_42999,N_43768);
nand U48820 (N_48820,N_44436,N_40687);
or U48821 (N_48821,N_41674,N_44563);
and U48822 (N_48822,N_40654,N_42057);
xnor U48823 (N_48823,N_40914,N_42090);
xnor U48824 (N_48824,N_40472,N_40601);
nor U48825 (N_48825,N_41440,N_43171);
and U48826 (N_48826,N_41492,N_42286);
xnor U48827 (N_48827,N_43773,N_40316);
nor U48828 (N_48828,N_42182,N_41741);
or U48829 (N_48829,N_44229,N_42997);
nand U48830 (N_48830,N_42846,N_44652);
nor U48831 (N_48831,N_44316,N_43394);
and U48832 (N_48832,N_43447,N_44895);
nand U48833 (N_48833,N_44882,N_41256);
xor U48834 (N_48834,N_41408,N_40746);
or U48835 (N_48835,N_43338,N_40294);
nand U48836 (N_48836,N_44930,N_40457);
or U48837 (N_48837,N_43273,N_43919);
and U48838 (N_48838,N_42327,N_41025);
and U48839 (N_48839,N_40004,N_42297);
nor U48840 (N_48840,N_41562,N_43177);
nor U48841 (N_48841,N_42254,N_42345);
and U48842 (N_48842,N_44201,N_44889);
nor U48843 (N_48843,N_44780,N_43004);
nor U48844 (N_48844,N_43514,N_40783);
and U48845 (N_48845,N_44848,N_42045);
nor U48846 (N_48846,N_41737,N_40595);
nor U48847 (N_48847,N_41388,N_40376);
and U48848 (N_48848,N_42260,N_42632);
or U48849 (N_48849,N_42823,N_41310);
or U48850 (N_48850,N_40104,N_41855);
and U48851 (N_48851,N_40451,N_43546);
or U48852 (N_48852,N_40679,N_42514);
nand U48853 (N_48853,N_44929,N_40892);
or U48854 (N_48854,N_40665,N_44694);
or U48855 (N_48855,N_40556,N_43250);
nor U48856 (N_48856,N_42767,N_40484);
nor U48857 (N_48857,N_41253,N_41502);
nor U48858 (N_48858,N_44195,N_44409);
nor U48859 (N_48859,N_40517,N_40286);
nand U48860 (N_48860,N_40723,N_43115);
or U48861 (N_48861,N_41730,N_40663);
nor U48862 (N_48862,N_41085,N_43777);
or U48863 (N_48863,N_43484,N_42722);
nor U48864 (N_48864,N_44975,N_42349);
and U48865 (N_48865,N_44597,N_43067);
nand U48866 (N_48866,N_42790,N_40164);
nor U48867 (N_48867,N_42500,N_44839);
and U48868 (N_48868,N_43765,N_42365);
and U48869 (N_48869,N_41897,N_42136);
or U48870 (N_48870,N_42506,N_40445);
or U48871 (N_48871,N_41385,N_43979);
xnor U48872 (N_48872,N_43684,N_43387);
nand U48873 (N_48873,N_42466,N_42190);
xor U48874 (N_48874,N_40227,N_40643);
and U48875 (N_48875,N_41610,N_43401);
nor U48876 (N_48876,N_40842,N_44181);
nand U48877 (N_48877,N_41294,N_40997);
nand U48878 (N_48878,N_41871,N_44333);
or U48879 (N_48879,N_41406,N_44185);
nand U48880 (N_48880,N_44863,N_44382);
or U48881 (N_48881,N_44944,N_40869);
nor U48882 (N_48882,N_44371,N_42779);
nand U48883 (N_48883,N_40261,N_40300);
and U48884 (N_48884,N_40442,N_42556);
xnor U48885 (N_48885,N_44209,N_43719);
nor U48886 (N_48886,N_44573,N_44245);
or U48887 (N_48887,N_44672,N_43805);
nand U48888 (N_48888,N_42581,N_43065);
or U48889 (N_48889,N_42182,N_43077);
or U48890 (N_48890,N_44103,N_42127);
nand U48891 (N_48891,N_44272,N_42381);
or U48892 (N_48892,N_40123,N_41215);
xor U48893 (N_48893,N_44836,N_40731);
xnor U48894 (N_48894,N_41343,N_41382);
or U48895 (N_48895,N_43056,N_40202);
nor U48896 (N_48896,N_40981,N_42360);
nand U48897 (N_48897,N_41156,N_44482);
and U48898 (N_48898,N_44723,N_44440);
xor U48899 (N_48899,N_42814,N_40677);
nand U48900 (N_48900,N_43697,N_44794);
nand U48901 (N_48901,N_40090,N_40874);
xor U48902 (N_48902,N_44978,N_40298);
nand U48903 (N_48903,N_43687,N_43945);
or U48904 (N_48904,N_42333,N_42940);
and U48905 (N_48905,N_41402,N_42918);
or U48906 (N_48906,N_41822,N_43564);
and U48907 (N_48907,N_42502,N_41444);
xor U48908 (N_48908,N_44227,N_41320);
nand U48909 (N_48909,N_41734,N_40590);
nand U48910 (N_48910,N_41145,N_44349);
or U48911 (N_48911,N_43692,N_42105);
or U48912 (N_48912,N_40673,N_41169);
nand U48913 (N_48913,N_41863,N_43540);
and U48914 (N_48914,N_42537,N_42644);
and U48915 (N_48915,N_44213,N_40399);
and U48916 (N_48916,N_42097,N_44197);
nor U48917 (N_48917,N_40480,N_41059);
xor U48918 (N_48918,N_41837,N_41886);
nand U48919 (N_48919,N_41382,N_44410);
nor U48920 (N_48920,N_42077,N_41678);
nand U48921 (N_48921,N_44300,N_43258);
nand U48922 (N_48922,N_43876,N_42512);
xor U48923 (N_48923,N_44129,N_41500);
nor U48924 (N_48924,N_41746,N_42001);
and U48925 (N_48925,N_41718,N_40789);
nor U48926 (N_48926,N_44400,N_41936);
or U48927 (N_48927,N_44749,N_40243);
and U48928 (N_48928,N_43685,N_42834);
or U48929 (N_48929,N_40070,N_41282);
xnor U48930 (N_48930,N_41921,N_42902);
and U48931 (N_48931,N_41342,N_42046);
or U48932 (N_48932,N_41628,N_44703);
nor U48933 (N_48933,N_40898,N_41759);
xnor U48934 (N_48934,N_42613,N_41297);
xnor U48935 (N_48935,N_41918,N_43820);
xnor U48936 (N_48936,N_42528,N_42405);
nand U48937 (N_48937,N_41531,N_40301);
and U48938 (N_48938,N_40508,N_41740);
nand U48939 (N_48939,N_42686,N_42141);
nor U48940 (N_48940,N_44527,N_43453);
nor U48941 (N_48941,N_42555,N_41717);
or U48942 (N_48942,N_40577,N_43696);
nor U48943 (N_48943,N_41364,N_44742);
nand U48944 (N_48944,N_40516,N_42737);
nor U48945 (N_48945,N_42786,N_40725);
and U48946 (N_48946,N_41320,N_43997);
nand U48947 (N_48947,N_41834,N_40932);
xnor U48948 (N_48948,N_40770,N_42964);
and U48949 (N_48949,N_41770,N_43818);
nand U48950 (N_48950,N_42474,N_40963);
xor U48951 (N_48951,N_41493,N_43096);
nand U48952 (N_48952,N_42747,N_42628);
xnor U48953 (N_48953,N_40855,N_43627);
or U48954 (N_48954,N_40154,N_43235);
xnor U48955 (N_48955,N_41460,N_43695);
nand U48956 (N_48956,N_41558,N_42748);
nor U48957 (N_48957,N_43773,N_40752);
and U48958 (N_48958,N_43562,N_41022);
and U48959 (N_48959,N_40613,N_44833);
nand U48960 (N_48960,N_40499,N_43094);
nand U48961 (N_48961,N_41057,N_44919);
nor U48962 (N_48962,N_42538,N_44667);
or U48963 (N_48963,N_40985,N_41358);
or U48964 (N_48964,N_43153,N_43504);
nor U48965 (N_48965,N_44104,N_40956);
xor U48966 (N_48966,N_40734,N_42665);
and U48967 (N_48967,N_40106,N_41315);
nor U48968 (N_48968,N_40816,N_40533);
or U48969 (N_48969,N_44984,N_44959);
and U48970 (N_48970,N_42007,N_43434);
or U48971 (N_48971,N_44886,N_42579);
or U48972 (N_48972,N_43608,N_42947);
nand U48973 (N_48973,N_44622,N_44434);
or U48974 (N_48974,N_43297,N_40289);
and U48975 (N_48975,N_44136,N_44920);
xor U48976 (N_48976,N_40197,N_41250);
and U48977 (N_48977,N_44501,N_41220);
or U48978 (N_48978,N_42685,N_40197);
and U48979 (N_48979,N_43440,N_40069);
or U48980 (N_48980,N_41296,N_44267);
nor U48981 (N_48981,N_42627,N_42576);
nand U48982 (N_48982,N_41255,N_41994);
xor U48983 (N_48983,N_44757,N_41716);
and U48984 (N_48984,N_43151,N_43475);
nand U48985 (N_48985,N_44099,N_40123);
and U48986 (N_48986,N_42476,N_41038);
nor U48987 (N_48987,N_42556,N_43060);
xnor U48988 (N_48988,N_42785,N_43550);
xor U48989 (N_48989,N_41873,N_43831);
xnor U48990 (N_48990,N_42612,N_41738);
xor U48991 (N_48991,N_43333,N_43991);
xnor U48992 (N_48992,N_41956,N_44639);
xnor U48993 (N_48993,N_42869,N_42281);
xnor U48994 (N_48994,N_43564,N_42167);
nand U48995 (N_48995,N_42124,N_43941);
nor U48996 (N_48996,N_42611,N_43772);
and U48997 (N_48997,N_40532,N_44259);
or U48998 (N_48998,N_44525,N_42496);
or U48999 (N_48999,N_41927,N_40389);
nor U49000 (N_49000,N_42211,N_43767);
and U49001 (N_49001,N_42552,N_42374);
nor U49002 (N_49002,N_40210,N_43086);
and U49003 (N_49003,N_40990,N_43397);
nor U49004 (N_49004,N_42158,N_43605);
xnor U49005 (N_49005,N_41653,N_42933);
or U49006 (N_49006,N_44084,N_40423);
nand U49007 (N_49007,N_44031,N_40726);
nor U49008 (N_49008,N_41691,N_42303);
nand U49009 (N_49009,N_42919,N_40734);
nand U49010 (N_49010,N_40964,N_44323);
xnor U49011 (N_49011,N_41499,N_44180);
nor U49012 (N_49012,N_40156,N_44907);
nand U49013 (N_49013,N_43888,N_41616);
and U49014 (N_49014,N_44139,N_41089);
and U49015 (N_49015,N_43703,N_40948);
and U49016 (N_49016,N_40517,N_40663);
xnor U49017 (N_49017,N_44128,N_40146);
or U49018 (N_49018,N_43399,N_41923);
nand U49019 (N_49019,N_41737,N_42531);
xnor U49020 (N_49020,N_40887,N_41719);
and U49021 (N_49021,N_44105,N_40507);
or U49022 (N_49022,N_41434,N_40185);
or U49023 (N_49023,N_40011,N_44557);
or U49024 (N_49024,N_41307,N_41422);
and U49025 (N_49025,N_43552,N_43501);
nor U49026 (N_49026,N_44714,N_40487);
xor U49027 (N_49027,N_41610,N_43805);
or U49028 (N_49028,N_42845,N_43601);
and U49029 (N_49029,N_40780,N_43539);
and U49030 (N_49030,N_40921,N_42326);
nor U49031 (N_49031,N_41847,N_44115);
xor U49032 (N_49032,N_44836,N_40262);
xor U49033 (N_49033,N_44389,N_41523);
xor U49034 (N_49034,N_43040,N_42338);
nand U49035 (N_49035,N_41491,N_41871);
or U49036 (N_49036,N_40246,N_43862);
nand U49037 (N_49037,N_42583,N_44134);
or U49038 (N_49038,N_43370,N_43628);
xor U49039 (N_49039,N_42946,N_44420);
nor U49040 (N_49040,N_43300,N_41620);
and U49041 (N_49041,N_44401,N_41504);
and U49042 (N_49042,N_41820,N_40659);
and U49043 (N_49043,N_40671,N_42028);
and U49044 (N_49044,N_42731,N_41887);
and U49045 (N_49045,N_42917,N_43913);
xnor U49046 (N_49046,N_42726,N_41080);
or U49047 (N_49047,N_44369,N_44670);
xor U49048 (N_49048,N_41624,N_41786);
or U49049 (N_49049,N_42178,N_44867);
nor U49050 (N_49050,N_41597,N_41964);
or U49051 (N_49051,N_41776,N_43840);
or U49052 (N_49052,N_42399,N_43480);
xnor U49053 (N_49053,N_40046,N_43143);
nor U49054 (N_49054,N_42820,N_42640);
nor U49055 (N_49055,N_44260,N_41637);
xor U49056 (N_49056,N_40652,N_44825);
and U49057 (N_49057,N_40102,N_42476);
nor U49058 (N_49058,N_43663,N_41865);
and U49059 (N_49059,N_44041,N_44614);
and U49060 (N_49060,N_44993,N_41458);
or U49061 (N_49061,N_43771,N_40342);
xnor U49062 (N_49062,N_43180,N_40169);
or U49063 (N_49063,N_41289,N_42433);
nor U49064 (N_49064,N_40768,N_44925);
or U49065 (N_49065,N_42351,N_44961);
and U49066 (N_49066,N_41756,N_44742);
xor U49067 (N_49067,N_42075,N_44926);
nor U49068 (N_49068,N_43520,N_44128);
or U49069 (N_49069,N_40951,N_44834);
nand U49070 (N_49070,N_44309,N_43547);
nor U49071 (N_49071,N_40221,N_43593);
xnor U49072 (N_49072,N_43422,N_41563);
and U49073 (N_49073,N_40438,N_44115);
and U49074 (N_49074,N_43903,N_44634);
nand U49075 (N_49075,N_40500,N_43988);
nor U49076 (N_49076,N_42329,N_43160);
or U49077 (N_49077,N_40842,N_41739);
xor U49078 (N_49078,N_43992,N_44170);
xnor U49079 (N_49079,N_44789,N_44643);
nand U49080 (N_49080,N_40273,N_44987);
and U49081 (N_49081,N_43985,N_41366);
nand U49082 (N_49082,N_43252,N_44769);
nand U49083 (N_49083,N_42651,N_40560);
nor U49084 (N_49084,N_43631,N_42614);
xor U49085 (N_49085,N_42409,N_43523);
nor U49086 (N_49086,N_40777,N_40289);
xor U49087 (N_49087,N_43955,N_40616);
nand U49088 (N_49088,N_42648,N_43047);
and U49089 (N_49089,N_41486,N_41823);
xor U49090 (N_49090,N_43221,N_44157);
nand U49091 (N_49091,N_42508,N_40257);
nand U49092 (N_49092,N_43110,N_43822);
or U49093 (N_49093,N_41786,N_44287);
nand U49094 (N_49094,N_40346,N_40017);
xnor U49095 (N_49095,N_40134,N_41381);
nor U49096 (N_49096,N_41823,N_43206);
nor U49097 (N_49097,N_40440,N_42417);
nor U49098 (N_49098,N_42608,N_44608);
xnor U49099 (N_49099,N_42249,N_41636);
and U49100 (N_49100,N_41652,N_41295);
and U49101 (N_49101,N_41878,N_44624);
and U49102 (N_49102,N_43016,N_41066);
or U49103 (N_49103,N_42628,N_41055);
nor U49104 (N_49104,N_40757,N_40995);
or U49105 (N_49105,N_44178,N_40226);
xor U49106 (N_49106,N_43491,N_41905);
nor U49107 (N_49107,N_41840,N_42568);
xnor U49108 (N_49108,N_41026,N_41451);
nor U49109 (N_49109,N_40011,N_41274);
nor U49110 (N_49110,N_42016,N_40900);
nor U49111 (N_49111,N_44938,N_44936);
xnor U49112 (N_49112,N_43191,N_43444);
and U49113 (N_49113,N_40777,N_44632);
xnor U49114 (N_49114,N_44809,N_41010);
nor U49115 (N_49115,N_40656,N_43130);
and U49116 (N_49116,N_44776,N_42773);
xor U49117 (N_49117,N_41679,N_42386);
or U49118 (N_49118,N_41270,N_42411);
xor U49119 (N_49119,N_43955,N_41419);
xnor U49120 (N_49120,N_40903,N_44226);
and U49121 (N_49121,N_43191,N_40048);
and U49122 (N_49122,N_44682,N_40377);
xnor U49123 (N_49123,N_41849,N_41521);
or U49124 (N_49124,N_44560,N_40141);
nand U49125 (N_49125,N_41169,N_43905);
xnor U49126 (N_49126,N_42162,N_40304);
nand U49127 (N_49127,N_42634,N_41568);
xnor U49128 (N_49128,N_44580,N_41306);
and U49129 (N_49129,N_40918,N_43618);
xor U49130 (N_49130,N_40484,N_43531);
or U49131 (N_49131,N_44028,N_41922);
and U49132 (N_49132,N_41432,N_44018);
nand U49133 (N_49133,N_41425,N_42521);
xor U49134 (N_49134,N_40243,N_42348);
xnor U49135 (N_49135,N_41620,N_42959);
nor U49136 (N_49136,N_43370,N_42333);
or U49137 (N_49137,N_43461,N_44504);
xor U49138 (N_49138,N_40501,N_40086);
xnor U49139 (N_49139,N_41055,N_44464);
nor U49140 (N_49140,N_44072,N_43227);
or U49141 (N_49141,N_41627,N_43187);
xnor U49142 (N_49142,N_42342,N_41666);
or U49143 (N_49143,N_40718,N_40393);
nand U49144 (N_49144,N_44035,N_44890);
nor U49145 (N_49145,N_43763,N_42959);
and U49146 (N_49146,N_43188,N_40389);
or U49147 (N_49147,N_44873,N_40578);
and U49148 (N_49148,N_42285,N_43750);
nand U49149 (N_49149,N_44793,N_40147);
nor U49150 (N_49150,N_42205,N_43750);
xor U49151 (N_49151,N_40776,N_40120);
or U49152 (N_49152,N_41995,N_43164);
nor U49153 (N_49153,N_42440,N_41201);
or U49154 (N_49154,N_40442,N_40595);
and U49155 (N_49155,N_42678,N_43347);
nor U49156 (N_49156,N_44254,N_40071);
nand U49157 (N_49157,N_41168,N_42094);
and U49158 (N_49158,N_44916,N_41581);
and U49159 (N_49159,N_41899,N_44976);
and U49160 (N_49160,N_42971,N_40263);
xnor U49161 (N_49161,N_43035,N_44281);
nand U49162 (N_49162,N_42312,N_41505);
nand U49163 (N_49163,N_44644,N_41760);
nor U49164 (N_49164,N_44048,N_40235);
nand U49165 (N_49165,N_44474,N_40230);
xnor U49166 (N_49166,N_41850,N_41060);
nor U49167 (N_49167,N_41117,N_41934);
or U49168 (N_49168,N_44114,N_42899);
or U49169 (N_49169,N_42813,N_41469);
nand U49170 (N_49170,N_40329,N_44821);
and U49171 (N_49171,N_42941,N_42137);
and U49172 (N_49172,N_43434,N_41180);
or U49173 (N_49173,N_40241,N_41978);
or U49174 (N_49174,N_40505,N_40945);
or U49175 (N_49175,N_43867,N_43070);
nor U49176 (N_49176,N_41231,N_40690);
or U49177 (N_49177,N_43236,N_42203);
or U49178 (N_49178,N_44005,N_43973);
nand U49179 (N_49179,N_41723,N_44655);
xor U49180 (N_49180,N_44395,N_42915);
and U49181 (N_49181,N_44186,N_44211);
or U49182 (N_49182,N_42429,N_40848);
nor U49183 (N_49183,N_44908,N_42685);
and U49184 (N_49184,N_42075,N_41524);
xnor U49185 (N_49185,N_42575,N_44160);
nand U49186 (N_49186,N_40606,N_42122);
nor U49187 (N_49187,N_42052,N_41004);
and U49188 (N_49188,N_42382,N_41305);
xor U49189 (N_49189,N_40455,N_44724);
nand U49190 (N_49190,N_43823,N_44598);
nor U49191 (N_49191,N_42966,N_43409);
and U49192 (N_49192,N_41460,N_40065);
and U49193 (N_49193,N_40980,N_44001);
nor U49194 (N_49194,N_44461,N_41185);
nand U49195 (N_49195,N_43629,N_44570);
nor U49196 (N_49196,N_44672,N_41513);
nor U49197 (N_49197,N_41717,N_42905);
nor U49198 (N_49198,N_40598,N_42658);
and U49199 (N_49199,N_43981,N_40337);
nand U49200 (N_49200,N_42364,N_43993);
nor U49201 (N_49201,N_44758,N_41015);
xor U49202 (N_49202,N_42094,N_40625);
nand U49203 (N_49203,N_40528,N_42727);
or U49204 (N_49204,N_40774,N_40057);
xnor U49205 (N_49205,N_40204,N_42719);
xor U49206 (N_49206,N_40745,N_43598);
and U49207 (N_49207,N_43151,N_44674);
xor U49208 (N_49208,N_41710,N_40108);
or U49209 (N_49209,N_43909,N_42133);
xnor U49210 (N_49210,N_40074,N_43589);
xnor U49211 (N_49211,N_42177,N_42678);
and U49212 (N_49212,N_44555,N_40120);
xor U49213 (N_49213,N_40973,N_42389);
nand U49214 (N_49214,N_43310,N_44335);
xnor U49215 (N_49215,N_43293,N_40707);
xor U49216 (N_49216,N_40843,N_42887);
xor U49217 (N_49217,N_42669,N_43307);
xor U49218 (N_49218,N_41845,N_40520);
nor U49219 (N_49219,N_43314,N_44722);
or U49220 (N_49220,N_44591,N_42101);
nand U49221 (N_49221,N_43486,N_43469);
xor U49222 (N_49222,N_44348,N_43026);
nor U49223 (N_49223,N_40658,N_41075);
and U49224 (N_49224,N_40520,N_44777);
or U49225 (N_49225,N_40014,N_43392);
or U49226 (N_49226,N_44391,N_43944);
nor U49227 (N_49227,N_41187,N_40843);
nand U49228 (N_49228,N_42252,N_41152);
and U49229 (N_49229,N_43318,N_42123);
nand U49230 (N_49230,N_41607,N_40878);
nor U49231 (N_49231,N_44400,N_42102);
nor U49232 (N_49232,N_41432,N_40323);
or U49233 (N_49233,N_44534,N_40742);
and U49234 (N_49234,N_40527,N_43489);
or U49235 (N_49235,N_41578,N_44133);
or U49236 (N_49236,N_43282,N_43548);
xnor U49237 (N_49237,N_43767,N_43324);
nor U49238 (N_49238,N_40089,N_42444);
or U49239 (N_49239,N_44263,N_44063);
nor U49240 (N_49240,N_43339,N_43412);
nand U49241 (N_49241,N_41672,N_40125);
or U49242 (N_49242,N_43727,N_43032);
and U49243 (N_49243,N_42556,N_41592);
nor U49244 (N_49244,N_42568,N_41638);
nor U49245 (N_49245,N_41601,N_41697);
nor U49246 (N_49246,N_43474,N_41969);
xnor U49247 (N_49247,N_41477,N_43119);
and U49248 (N_49248,N_40008,N_42764);
and U49249 (N_49249,N_43002,N_44564);
or U49250 (N_49250,N_41106,N_41088);
and U49251 (N_49251,N_41022,N_43526);
nor U49252 (N_49252,N_41479,N_40678);
xor U49253 (N_49253,N_44481,N_40408);
and U49254 (N_49254,N_41360,N_42602);
nand U49255 (N_49255,N_42794,N_44287);
or U49256 (N_49256,N_40011,N_44033);
or U49257 (N_49257,N_44656,N_40897);
and U49258 (N_49258,N_40961,N_43900);
nand U49259 (N_49259,N_41113,N_43372);
and U49260 (N_49260,N_42630,N_43229);
xor U49261 (N_49261,N_44097,N_42805);
nand U49262 (N_49262,N_41184,N_41956);
or U49263 (N_49263,N_42268,N_41187);
and U49264 (N_49264,N_42972,N_43444);
and U49265 (N_49265,N_42070,N_42266);
nor U49266 (N_49266,N_40293,N_42174);
and U49267 (N_49267,N_43465,N_44995);
or U49268 (N_49268,N_41607,N_40906);
or U49269 (N_49269,N_43491,N_42239);
xor U49270 (N_49270,N_40673,N_43646);
nor U49271 (N_49271,N_43236,N_40509);
or U49272 (N_49272,N_43263,N_43871);
nor U49273 (N_49273,N_44853,N_44830);
or U49274 (N_49274,N_42375,N_43083);
nand U49275 (N_49275,N_44845,N_43854);
nor U49276 (N_49276,N_42009,N_44893);
and U49277 (N_49277,N_42605,N_44421);
nor U49278 (N_49278,N_40242,N_44548);
nand U49279 (N_49279,N_41251,N_41503);
xor U49280 (N_49280,N_44100,N_41403);
xor U49281 (N_49281,N_43953,N_42043);
nor U49282 (N_49282,N_43821,N_43572);
nand U49283 (N_49283,N_41828,N_43923);
nand U49284 (N_49284,N_44258,N_44948);
nand U49285 (N_49285,N_42726,N_44678);
or U49286 (N_49286,N_43379,N_40691);
nand U49287 (N_49287,N_40948,N_41108);
and U49288 (N_49288,N_42372,N_44270);
or U49289 (N_49289,N_44002,N_44870);
xor U49290 (N_49290,N_44506,N_41543);
and U49291 (N_49291,N_41908,N_41434);
nand U49292 (N_49292,N_42864,N_43603);
xnor U49293 (N_49293,N_41875,N_43336);
xor U49294 (N_49294,N_41726,N_44303);
or U49295 (N_49295,N_40149,N_40754);
xnor U49296 (N_49296,N_40042,N_40250);
nand U49297 (N_49297,N_40974,N_43957);
nand U49298 (N_49298,N_44241,N_41740);
xnor U49299 (N_49299,N_40683,N_43305);
nand U49300 (N_49300,N_42529,N_40418);
or U49301 (N_49301,N_40189,N_44299);
or U49302 (N_49302,N_44282,N_40312);
xnor U49303 (N_49303,N_43632,N_40634);
xor U49304 (N_49304,N_41970,N_43764);
nand U49305 (N_49305,N_44693,N_42815);
or U49306 (N_49306,N_44915,N_44692);
and U49307 (N_49307,N_44511,N_42062);
or U49308 (N_49308,N_43632,N_41147);
nor U49309 (N_49309,N_42769,N_43513);
or U49310 (N_49310,N_44469,N_40133);
nor U49311 (N_49311,N_44258,N_43794);
xnor U49312 (N_49312,N_43474,N_41934);
and U49313 (N_49313,N_41130,N_42595);
nor U49314 (N_49314,N_41619,N_41349);
nand U49315 (N_49315,N_43002,N_44668);
or U49316 (N_49316,N_40058,N_43658);
nor U49317 (N_49317,N_42385,N_43429);
and U49318 (N_49318,N_43296,N_41527);
and U49319 (N_49319,N_42333,N_42732);
nor U49320 (N_49320,N_40217,N_43376);
and U49321 (N_49321,N_40319,N_40251);
or U49322 (N_49322,N_40545,N_41586);
xor U49323 (N_49323,N_42818,N_44386);
or U49324 (N_49324,N_42788,N_44036);
or U49325 (N_49325,N_40982,N_43112);
xor U49326 (N_49326,N_40109,N_44990);
nor U49327 (N_49327,N_40545,N_44270);
and U49328 (N_49328,N_44924,N_42042);
nor U49329 (N_49329,N_44307,N_40005);
nand U49330 (N_49330,N_42546,N_41568);
and U49331 (N_49331,N_42087,N_42018);
xor U49332 (N_49332,N_43677,N_43407);
and U49333 (N_49333,N_44712,N_42717);
nand U49334 (N_49334,N_41023,N_43140);
and U49335 (N_49335,N_41550,N_40650);
nor U49336 (N_49336,N_40999,N_40393);
or U49337 (N_49337,N_42913,N_43917);
and U49338 (N_49338,N_42934,N_43740);
or U49339 (N_49339,N_42305,N_44346);
or U49340 (N_49340,N_40400,N_40706);
xor U49341 (N_49341,N_42015,N_41954);
xnor U49342 (N_49342,N_44204,N_42574);
or U49343 (N_49343,N_42012,N_40081);
nor U49344 (N_49344,N_43290,N_41148);
and U49345 (N_49345,N_44890,N_43386);
xor U49346 (N_49346,N_43665,N_40329);
xor U49347 (N_49347,N_43193,N_41905);
nor U49348 (N_49348,N_40272,N_42534);
xor U49349 (N_49349,N_42520,N_41849);
and U49350 (N_49350,N_43394,N_44426);
xnor U49351 (N_49351,N_41796,N_40175);
and U49352 (N_49352,N_44792,N_41157);
nand U49353 (N_49353,N_40803,N_41660);
or U49354 (N_49354,N_40482,N_41290);
xnor U49355 (N_49355,N_42657,N_44002);
and U49356 (N_49356,N_40926,N_40344);
nand U49357 (N_49357,N_43983,N_44670);
nor U49358 (N_49358,N_41518,N_43968);
nor U49359 (N_49359,N_41428,N_43925);
and U49360 (N_49360,N_42151,N_42809);
nor U49361 (N_49361,N_40321,N_42191);
nand U49362 (N_49362,N_41166,N_41771);
nand U49363 (N_49363,N_42898,N_41129);
xor U49364 (N_49364,N_40960,N_41405);
xor U49365 (N_49365,N_42983,N_41736);
or U49366 (N_49366,N_41117,N_42333);
or U49367 (N_49367,N_41023,N_40567);
nand U49368 (N_49368,N_43426,N_44772);
or U49369 (N_49369,N_41212,N_44911);
or U49370 (N_49370,N_40221,N_43096);
or U49371 (N_49371,N_44808,N_40633);
nand U49372 (N_49372,N_42199,N_44694);
and U49373 (N_49373,N_41226,N_43101);
nand U49374 (N_49374,N_43660,N_43760);
nand U49375 (N_49375,N_40979,N_44512);
nor U49376 (N_49376,N_42582,N_44661);
nand U49377 (N_49377,N_42164,N_44810);
xnor U49378 (N_49378,N_40047,N_40383);
and U49379 (N_49379,N_44421,N_41648);
nand U49380 (N_49380,N_40324,N_42696);
nand U49381 (N_49381,N_42879,N_41506);
or U49382 (N_49382,N_44367,N_43391);
nor U49383 (N_49383,N_42218,N_41119);
and U49384 (N_49384,N_44167,N_41007);
nand U49385 (N_49385,N_42052,N_43549);
or U49386 (N_49386,N_41547,N_41943);
nor U49387 (N_49387,N_44186,N_43789);
xor U49388 (N_49388,N_43844,N_42063);
nand U49389 (N_49389,N_41923,N_41602);
nand U49390 (N_49390,N_42764,N_42602);
xnor U49391 (N_49391,N_44964,N_44993);
nand U49392 (N_49392,N_40142,N_41564);
xnor U49393 (N_49393,N_41997,N_43061);
or U49394 (N_49394,N_43387,N_40559);
nand U49395 (N_49395,N_44634,N_40426);
and U49396 (N_49396,N_42450,N_41938);
and U49397 (N_49397,N_41197,N_41983);
nor U49398 (N_49398,N_42620,N_40744);
nor U49399 (N_49399,N_40264,N_40138);
nand U49400 (N_49400,N_42319,N_44831);
and U49401 (N_49401,N_41831,N_42573);
nand U49402 (N_49402,N_43529,N_43359);
nor U49403 (N_49403,N_44366,N_41792);
nor U49404 (N_49404,N_42850,N_44856);
or U49405 (N_49405,N_41382,N_41425);
nand U49406 (N_49406,N_44417,N_43988);
nor U49407 (N_49407,N_41575,N_41078);
or U49408 (N_49408,N_43344,N_42896);
and U49409 (N_49409,N_41248,N_42609);
and U49410 (N_49410,N_42346,N_43275);
or U49411 (N_49411,N_44341,N_42832);
nor U49412 (N_49412,N_43304,N_44201);
nor U49413 (N_49413,N_41262,N_40808);
xnor U49414 (N_49414,N_41548,N_41497);
xnor U49415 (N_49415,N_44557,N_43754);
xor U49416 (N_49416,N_42337,N_40127);
nor U49417 (N_49417,N_43156,N_40129);
xor U49418 (N_49418,N_43786,N_42986);
nor U49419 (N_49419,N_41219,N_43447);
and U49420 (N_49420,N_40501,N_44002);
nor U49421 (N_49421,N_42494,N_42246);
xor U49422 (N_49422,N_41750,N_43658);
and U49423 (N_49423,N_42219,N_42684);
xnor U49424 (N_49424,N_43671,N_44434);
nand U49425 (N_49425,N_42928,N_41352);
nand U49426 (N_49426,N_43393,N_40442);
nor U49427 (N_49427,N_44266,N_43637);
nor U49428 (N_49428,N_43596,N_40536);
nor U49429 (N_49429,N_40876,N_41529);
and U49430 (N_49430,N_42693,N_42245);
nor U49431 (N_49431,N_40020,N_40425);
nand U49432 (N_49432,N_42916,N_43015);
and U49433 (N_49433,N_44951,N_40806);
and U49434 (N_49434,N_42856,N_41703);
nor U49435 (N_49435,N_44693,N_44084);
and U49436 (N_49436,N_44563,N_44188);
or U49437 (N_49437,N_41580,N_40829);
or U49438 (N_49438,N_44124,N_40997);
nor U49439 (N_49439,N_40631,N_41502);
nand U49440 (N_49440,N_43327,N_40519);
or U49441 (N_49441,N_44475,N_43153);
nand U49442 (N_49442,N_42027,N_42885);
xnor U49443 (N_49443,N_41536,N_43279);
or U49444 (N_49444,N_40824,N_44994);
and U49445 (N_49445,N_40162,N_41758);
nand U49446 (N_49446,N_44932,N_41132);
or U49447 (N_49447,N_43612,N_40064);
xnor U49448 (N_49448,N_43822,N_42669);
xor U49449 (N_49449,N_43451,N_42724);
nand U49450 (N_49450,N_42315,N_42046);
xnor U49451 (N_49451,N_44937,N_44356);
or U49452 (N_49452,N_40885,N_43438);
nor U49453 (N_49453,N_43605,N_40194);
nand U49454 (N_49454,N_42207,N_44968);
and U49455 (N_49455,N_40238,N_44535);
nor U49456 (N_49456,N_42171,N_40524);
nand U49457 (N_49457,N_44845,N_43856);
nand U49458 (N_49458,N_44335,N_42739);
xor U49459 (N_49459,N_44148,N_44433);
nor U49460 (N_49460,N_43291,N_40520);
or U49461 (N_49461,N_41819,N_42257);
xnor U49462 (N_49462,N_40401,N_44801);
or U49463 (N_49463,N_40588,N_41527);
and U49464 (N_49464,N_42255,N_44332);
nand U49465 (N_49465,N_43151,N_43793);
or U49466 (N_49466,N_44197,N_41819);
and U49467 (N_49467,N_41927,N_43349);
nor U49468 (N_49468,N_43667,N_40341);
nor U49469 (N_49469,N_44275,N_42480);
xnor U49470 (N_49470,N_40332,N_41597);
nor U49471 (N_49471,N_42477,N_42112);
xnor U49472 (N_49472,N_43234,N_41521);
nor U49473 (N_49473,N_44165,N_43378);
xor U49474 (N_49474,N_43818,N_43363);
xor U49475 (N_49475,N_44471,N_41744);
xnor U49476 (N_49476,N_40664,N_41337);
or U49477 (N_49477,N_40243,N_41602);
and U49478 (N_49478,N_42084,N_40226);
xnor U49479 (N_49479,N_44682,N_43564);
xor U49480 (N_49480,N_43118,N_43159);
or U49481 (N_49481,N_42185,N_44901);
or U49482 (N_49482,N_43731,N_40071);
nor U49483 (N_49483,N_42056,N_41020);
nand U49484 (N_49484,N_44441,N_43327);
nand U49485 (N_49485,N_41785,N_41385);
nand U49486 (N_49486,N_40689,N_41518);
xor U49487 (N_49487,N_41913,N_41882);
and U49488 (N_49488,N_42056,N_42008);
nand U49489 (N_49489,N_40128,N_40174);
or U49490 (N_49490,N_44282,N_40999);
and U49491 (N_49491,N_40033,N_44528);
or U49492 (N_49492,N_42649,N_40043);
nand U49493 (N_49493,N_42278,N_41807);
nor U49494 (N_49494,N_43115,N_41728);
nand U49495 (N_49495,N_44945,N_42327);
xor U49496 (N_49496,N_43707,N_40241);
xnor U49497 (N_49497,N_41304,N_41769);
nor U49498 (N_49498,N_40922,N_41366);
and U49499 (N_49499,N_40089,N_43963);
and U49500 (N_49500,N_40228,N_40552);
xor U49501 (N_49501,N_43212,N_42759);
xnor U49502 (N_49502,N_44126,N_40923);
xnor U49503 (N_49503,N_42449,N_44986);
xnor U49504 (N_49504,N_43121,N_43833);
and U49505 (N_49505,N_42097,N_42700);
nand U49506 (N_49506,N_40516,N_42417);
or U49507 (N_49507,N_43703,N_42843);
xnor U49508 (N_49508,N_41528,N_44296);
or U49509 (N_49509,N_41391,N_43193);
xnor U49510 (N_49510,N_44665,N_42323);
and U49511 (N_49511,N_42227,N_41836);
or U49512 (N_49512,N_40003,N_44754);
nand U49513 (N_49513,N_43127,N_41189);
xor U49514 (N_49514,N_43729,N_44201);
nor U49515 (N_49515,N_44476,N_41649);
nor U49516 (N_49516,N_44902,N_41725);
nor U49517 (N_49517,N_42215,N_41279);
nand U49518 (N_49518,N_40583,N_41165);
nor U49519 (N_49519,N_43093,N_43991);
nand U49520 (N_49520,N_43777,N_43540);
nor U49521 (N_49521,N_44560,N_43871);
or U49522 (N_49522,N_43005,N_41346);
nor U49523 (N_49523,N_41284,N_44125);
xnor U49524 (N_49524,N_41608,N_44482);
xor U49525 (N_49525,N_41716,N_44191);
xor U49526 (N_49526,N_41266,N_44347);
or U49527 (N_49527,N_44920,N_42411);
or U49528 (N_49528,N_42654,N_43338);
and U49529 (N_49529,N_41573,N_44150);
nand U49530 (N_49530,N_42901,N_42084);
xnor U49531 (N_49531,N_41807,N_43363);
xor U49532 (N_49532,N_41412,N_40620);
or U49533 (N_49533,N_42883,N_44003);
nor U49534 (N_49534,N_40343,N_40278);
nand U49535 (N_49535,N_44528,N_41087);
nor U49536 (N_49536,N_40386,N_40342);
nor U49537 (N_49537,N_40927,N_43733);
nor U49538 (N_49538,N_42291,N_40061);
nor U49539 (N_49539,N_42364,N_42845);
xor U49540 (N_49540,N_42056,N_44635);
nand U49541 (N_49541,N_44428,N_40295);
nand U49542 (N_49542,N_42746,N_43377);
nor U49543 (N_49543,N_43116,N_44661);
or U49544 (N_49544,N_40618,N_40667);
nand U49545 (N_49545,N_40259,N_44567);
nor U49546 (N_49546,N_40538,N_41504);
or U49547 (N_49547,N_40531,N_44744);
or U49548 (N_49548,N_40743,N_40315);
and U49549 (N_49549,N_44164,N_41438);
xor U49550 (N_49550,N_40100,N_44099);
xor U49551 (N_49551,N_44498,N_44851);
and U49552 (N_49552,N_41639,N_44283);
or U49553 (N_49553,N_42635,N_43992);
or U49554 (N_49554,N_41690,N_43324);
nand U49555 (N_49555,N_44110,N_44703);
nor U49556 (N_49556,N_44391,N_40112);
xnor U49557 (N_49557,N_41404,N_41639);
nor U49558 (N_49558,N_41593,N_40082);
or U49559 (N_49559,N_42602,N_42491);
nand U49560 (N_49560,N_41520,N_40381);
xnor U49561 (N_49561,N_42270,N_44560);
xor U49562 (N_49562,N_43813,N_41756);
or U49563 (N_49563,N_41047,N_43004);
nand U49564 (N_49564,N_41629,N_42857);
or U49565 (N_49565,N_40454,N_42101);
xor U49566 (N_49566,N_42419,N_43727);
and U49567 (N_49567,N_41670,N_43569);
or U49568 (N_49568,N_44206,N_40412);
nor U49569 (N_49569,N_40883,N_40192);
xor U49570 (N_49570,N_44320,N_44348);
and U49571 (N_49571,N_41740,N_44272);
or U49572 (N_49572,N_44879,N_44046);
or U49573 (N_49573,N_41101,N_43107);
and U49574 (N_49574,N_43469,N_40036);
xnor U49575 (N_49575,N_43174,N_41235);
nand U49576 (N_49576,N_42098,N_40222);
nor U49577 (N_49577,N_43232,N_41580);
and U49578 (N_49578,N_43372,N_41949);
or U49579 (N_49579,N_44606,N_41791);
nand U49580 (N_49580,N_41882,N_41727);
or U49581 (N_49581,N_42409,N_40623);
nor U49582 (N_49582,N_43282,N_40007);
or U49583 (N_49583,N_40469,N_40865);
and U49584 (N_49584,N_43441,N_43219);
xor U49585 (N_49585,N_43092,N_42101);
nand U49586 (N_49586,N_41809,N_40621);
or U49587 (N_49587,N_41844,N_41198);
and U49588 (N_49588,N_43625,N_44789);
nor U49589 (N_49589,N_40893,N_40083);
nand U49590 (N_49590,N_42731,N_40433);
nand U49591 (N_49591,N_40686,N_42457);
or U49592 (N_49592,N_40125,N_42743);
xnor U49593 (N_49593,N_44949,N_41066);
nor U49594 (N_49594,N_43377,N_41855);
xor U49595 (N_49595,N_44938,N_43761);
and U49596 (N_49596,N_41984,N_40479);
and U49597 (N_49597,N_41052,N_40436);
and U49598 (N_49598,N_42419,N_41437);
nor U49599 (N_49599,N_41987,N_44050);
or U49600 (N_49600,N_43020,N_42230);
xor U49601 (N_49601,N_43048,N_44096);
and U49602 (N_49602,N_40702,N_43855);
nand U49603 (N_49603,N_41602,N_41988);
xnor U49604 (N_49604,N_40080,N_43370);
or U49605 (N_49605,N_42037,N_40588);
nand U49606 (N_49606,N_41371,N_42947);
xnor U49607 (N_49607,N_42465,N_40275);
or U49608 (N_49608,N_43479,N_44948);
nor U49609 (N_49609,N_44071,N_44089);
nand U49610 (N_49610,N_44029,N_41093);
nor U49611 (N_49611,N_43211,N_41415);
nor U49612 (N_49612,N_41925,N_40125);
and U49613 (N_49613,N_41696,N_42690);
xor U49614 (N_49614,N_43680,N_43654);
and U49615 (N_49615,N_44195,N_43113);
nor U49616 (N_49616,N_43575,N_40288);
nand U49617 (N_49617,N_44343,N_40991);
nor U49618 (N_49618,N_42695,N_42227);
or U49619 (N_49619,N_42086,N_42577);
nor U49620 (N_49620,N_42994,N_40095);
xor U49621 (N_49621,N_42632,N_44077);
and U49622 (N_49622,N_42385,N_42658);
or U49623 (N_49623,N_41089,N_43152);
or U49624 (N_49624,N_40625,N_42354);
nor U49625 (N_49625,N_40119,N_44626);
and U49626 (N_49626,N_40040,N_43808);
nor U49627 (N_49627,N_42527,N_43719);
nor U49628 (N_49628,N_44511,N_43550);
nand U49629 (N_49629,N_43126,N_44316);
xnor U49630 (N_49630,N_42512,N_40032);
or U49631 (N_49631,N_40546,N_40464);
nand U49632 (N_49632,N_43050,N_41623);
xor U49633 (N_49633,N_44558,N_40497);
nor U49634 (N_49634,N_40304,N_40442);
or U49635 (N_49635,N_41541,N_42521);
nand U49636 (N_49636,N_43223,N_42540);
nor U49637 (N_49637,N_43355,N_42343);
nor U49638 (N_49638,N_44438,N_41876);
and U49639 (N_49639,N_42478,N_44453);
xor U49640 (N_49640,N_41164,N_44531);
and U49641 (N_49641,N_40107,N_43188);
or U49642 (N_49642,N_42062,N_41144);
nand U49643 (N_49643,N_40393,N_43318);
nand U49644 (N_49644,N_42110,N_44793);
and U49645 (N_49645,N_43744,N_41160);
xor U49646 (N_49646,N_40382,N_41778);
nor U49647 (N_49647,N_42618,N_41839);
nand U49648 (N_49648,N_40011,N_41891);
xor U49649 (N_49649,N_41314,N_42103);
or U49650 (N_49650,N_44988,N_43615);
and U49651 (N_49651,N_42386,N_40540);
nor U49652 (N_49652,N_43305,N_40969);
or U49653 (N_49653,N_44161,N_40155);
or U49654 (N_49654,N_44560,N_42574);
or U49655 (N_49655,N_42503,N_41995);
and U49656 (N_49656,N_40587,N_44316);
nor U49657 (N_49657,N_41103,N_41796);
xnor U49658 (N_49658,N_43089,N_40495);
nand U49659 (N_49659,N_40695,N_42731);
and U49660 (N_49660,N_42509,N_41427);
nor U49661 (N_49661,N_44729,N_40171);
xnor U49662 (N_49662,N_41957,N_43256);
or U49663 (N_49663,N_42463,N_42681);
nand U49664 (N_49664,N_41062,N_44135);
or U49665 (N_49665,N_40040,N_41601);
or U49666 (N_49666,N_42016,N_44062);
xor U49667 (N_49667,N_41243,N_41291);
nor U49668 (N_49668,N_43850,N_40208);
nand U49669 (N_49669,N_43970,N_40345);
nand U49670 (N_49670,N_41007,N_43155);
and U49671 (N_49671,N_44614,N_40657);
nand U49672 (N_49672,N_42015,N_40719);
and U49673 (N_49673,N_42893,N_42960);
or U49674 (N_49674,N_44426,N_44567);
and U49675 (N_49675,N_42287,N_42728);
nand U49676 (N_49676,N_44699,N_41245);
nor U49677 (N_49677,N_40175,N_44001);
xnor U49678 (N_49678,N_44639,N_42530);
nand U49679 (N_49679,N_44860,N_42740);
and U49680 (N_49680,N_43546,N_41401);
and U49681 (N_49681,N_42901,N_41068);
nand U49682 (N_49682,N_41413,N_40507);
xnor U49683 (N_49683,N_40684,N_43173);
nor U49684 (N_49684,N_43142,N_44675);
xnor U49685 (N_49685,N_44623,N_40010);
and U49686 (N_49686,N_42701,N_40814);
or U49687 (N_49687,N_44110,N_43964);
xor U49688 (N_49688,N_44221,N_40613);
or U49689 (N_49689,N_41860,N_44659);
nor U49690 (N_49690,N_44411,N_43600);
or U49691 (N_49691,N_44769,N_44711);
and U49692 (N_49692,N_41417,N_41086);
nand U49693 (N_49693,N_40334,N_43305);
xor U49694 (N_49694,N_44526,N_42754);
nand U49695 (N_49695,N_42550,N_44764);
nand U49696 (N_49696,N_42508,N_42385);
xnor U49697 (N_49697,N_41897,N_44774);
nor U49698 (N_49698,N_44293,N_43828);
nor U49699 (N_49699,N_42874,N_42971);
nand U49700 (N_49700,N_40691,N_41254);
or U49701 (N_49701,N_40550,N_40564);
xnor U49702 (N_49702,N_42001,N_41867);
and U49703 (N_49703,N_42887,N_42549);
nand U49704 (N_49704,N_44872,N_44474);
xnor U49705 (N_49705,N_42879,N_42306);
xor U49706 (N_49706,N_40821,N_44005);
nor U49707 (N_49707,N_44444,N_44665);
and U49708 (N_49708,N_44020,N_43195);
nor U49709 (N_49709,N_43440,N_44433);
or U49710 (N_49710,N_42164,N_44495);
xnor U49711 (N_49711,N_44383,N_42311);
and U49712 (N_49712,N_41923,N_42502);
nand U49713 (N_49713,N_40655,N_43560);
nor U49714 (N_49714,N_41104,N_42611);
xnor U49715 (N_49715,N_41922,N_41719);
nor U49716 (N_49716,N_41155,N_41103);
nor U49717 (N_49717,N_42471,N_43076);
nand U49718 (N_49718,N_43714,N_41634);
nor U49719 (N_49719,N_43192,N_41897);
or U49720 (N_49720,N_43460,N_43704);
and U49721 (N_49721,N_44661,N_42738);
xor U49722 (N_49722,N_44586,N_41305);
nor U49723 (N_49723,N_41119,N_44574);
or U49724 (N_49724,N_43404,N_43435);
or U49725 (N_49725,N_42303,N_43709);
and U49726 (N_49726,N_44085,N_43957);
or U49727 (N_49727,N_41612,N_42482);
and U49728 (N_49728,N_43429,N_44200);
or U49729 (N_49729,N_41770,N_40520);
xor U49730 (N_49730,N_44192,N_43048);
nor U49731 (N_49731,N_44186,N_43515);
xor U49732 (N_49732,N_40957,N_41408);
and U49733 (N_49733,N_40667,N_41667);
or U49734 (N_49734,N_42323,N_41164);
nor U49735 (N_49735,N_41120,N_43966);
nor U49736 (N_49736,N_40417,N_44537);
nor U49737 (N_49737,N_41983,N_40958);
nand U49738 (N_49738,N_42068,N_43335);
xor U49739 (N_49739,N_44467,N_40958);
or U49740 (N_49740,N_44205,N_42340);
nand U49741 (N_49741,N_41222,N_40218);
xor U49742 (N_49742,N_40804,N_42409);
nand U49743 (N_49743,N_41563,N_41290);
nor U49744 (N_49744,N_42975,N_44258);
or U49745 (N_49745,N_40717,N_41151);
xor U49746 (N_49746,N_41499,N_42631);
nand U49747 (N_49747,N_43277,N_40609);
nor U49748 (N_49748,N_40642,N_44347);
and U49749 (N_49749,N_42411,N_40903);
xnor U49750 (N_49750,N_42355,N_40348);
nand U49751 (N_49751,N_44057,N_43082);
nor U49752 (N_49752,N_42267,N_43602);
nor U49753 (N_49753,N_42756,N_42605);
nand U49754 (N_49754,N_43134,N_44030);
or U49755 (N_49755,N_44255,N_41615);
nand U49756 (N_49756,N_44231,N_42190);
or U49757 (N_49757,N_44186,N_40563);
nand U49758 (N_49758,N_42920,N_42993);
and U49759 (N_49759,N_40289,N_43629);
nand U49760 (N_49760,N_44693,N_44741);
or U49761 (N_49761,N_42933,N_44472);
xor U49762 (N_49762,N_44973,N_40860);
or U49763 (N_49763,N_42869,N_40403);
or U49764 (N_49764,N_40318,N_43612);
xor U49765 (N_49765,N_41759,N_44398);
nor U49766 (N_49766,N_41714,N_41879);
and U49767 (N_49767,N_44360,N_41583);
nand U49768 (N_49768,N_44636,N_40420);
nand U49769 (N_49769,N_40109,N_44161);
nor U49770 (N_49770,N_43527,N_42932);
and U49771 (N_49771,N_41283,N_41921);
and U49772 (N_49772,N_42096,N_40271);
xor U49773 (N_49773,N_42828,N_40377);
xor U49774 (N_49774,N_42530,N_43804);
nor U49775 (N_49775,N_41075,N_41246);
and U49776 (N_49776,N_44376,N_40643);
nor U49777 (N_49777,N_40620,N_41717);
nor U49778 (N_49778,N_41336,N_40386);
xor U49779 (N_49779,N_44860,N_43477);
or U49780 (N_49780,N_40364,N_42483);
or U49781 (N_49781,N_41146,N_44670);
nand U49782 (N_49782,N_42807,N_41651);
nor U49783 (N_49783,N_40122,N_41692);
xor U49784 (N_49784,N_44587,N_40390);
and U49785 (N_49785,N_42995,N_44924);
or U49786 (N_49786,N_40073,N_41942);
xnor U49787 (N_49787,N_43047,N_43134);
nand U49788 (N_49788,N_44963,N_41726);
nand U49789 (N_49789,N_44992,N_42509);
and U49790 (N_49790,N_44021,N_41383);
nand U49791 (N_49791,N_42922,N_41550);
or U49792 (N_49792,N_40546,N_41273);
and U49793 (N_49793,N_44165,N_44987);
nor U49794 (N_49794,N_43746,N_43484);
or U49795 (N_49795,N_44975,N_40502);
or U49796 (N_49796,N_41841,N_41649);
xor U49797 (N_49797,N_40241,N_40941);
nor U49798 (N_49798,N_41998,N_43131);
and U49799 (N_49799,N_42081,N_42921);
nor U49800 (N_49800,N_44665,N_43500);
nand U49801 (N_49801,N_42795,N_41021);
or U49802 (N_49802,N_44390,N_40281);
or U49803 (N_49803,N_44423,N_43098);
or U49804 (N_49804,N_42132,N_41532);
xor U49805 (N_49805,N_44637,N_41200);
nor U49806 (N_49806,N_40573,N_40234);
nand U49807 (N_49807,N_43699,N_42634);
nor U49808 (N_49808,N_44990,N_41188);
nor U49809 (N_49809,N_44526,N_40477);
or U49810 (N_49810,N_42868,N_42999);
or U49811 (N_49811,N_42900,N_42291);
nor U49812 (N_49812,N_41609,N_44464);
nor U49813 (N_49813,N_41024,N_42684);
and U49814 (N_49814,N_43550,N_41464);
nor U49815 (N_49815,N_43276,N_40901);
xnor U49816 (N_49816,N_40112,N_43967);
or U49817 (N_49817,N_44045,N_44852);
or U49818 (N_49818,N_40824,N_42221);
nand U49819 (N_49819,N_41259,N_43774);
or U49820 (N_49820,N_41888,N_42518);
nand U49821 (N_49821,N_43507,N_42892);
nand U49822 (N_49822,N_41187,N_40570);
nor U49823 (N_49823,N_43463,N_41207);
and U49824 (N_49824,N_44929,N_42376);
or U49825 (N_49825,N_42729,N_42959);
and U49826 (N_49826,N_44052,N_44620);
nor U49827 (N_49827,N_40984,N_40564);
xnor U49828 (N_49828,N_43916,N_43594);
or U49829 (N_49829,N_40220,N_40862);
xor U49830 (N_49830,N_40236,N_44268);
nand U49831 (N_49831,N_42569,N_43542);
or U49832 (N_49832,N_43633,N_40092);
or U49833 (N_49833,N_43225,N_43245);
and U49834 (N_49834,N_42058,N_40137);
or U49835 (N_49835,N_40928,N_42982);
or U49836 (N_49836,N_43422,N_40767);
xnor U49837 (N_49837,N_42544,N_40816);
nor U49838 (N_49838,N_44986,N_41112);
xnor U49839 (N_49839,N_42509,N_42149);
nor U49840 (N_49840,N_43599,N_40497);
nor U49841 (N_49841,N_43174,N_41496);
nor U49842 (N_49842,N_44628,N_40522);
and U49843 (N_49843,N_40244,N_44475);
xor U49844 (N_49844,N_42998,N_44341);
nand U49845 (N_49845,N_42536,N_43988);
nand U49846 (N_49846,N_44007,N_42425);
xor U49847 (N_49847,N_43593,N_42075);
xnor U49848 (N_49848,N_42591,N_40951);
nand U49849 (N_49849,N_41015,N_42337);
xnor U49850 (N_49850,N_41875,N_42545);
or U49851 (N_49851,N_42144,N_43000);
and U49852 (N_49852,N_42973,N_44800);
or U49853 (N_49853,N_44694,N_43056);
nand U49854 (N_49854,N_41407,N_44539);
xnor U49855 (N_49855,N_40910,N_44373);
and U49856 (N_49856,N_41176,N_44839);
nand U49857 (N_49857,N_42463,N_44869);
xnor U49858 (N_49858,N_40380,N_43343);
and U49859 (N_49859,N_41627,N_44742);
nor U49860 (N_49860,N_44781,N_40487);
nand U49861 (N_49861,N_44226,N_43599);
and U49862 (N_49862,N_42190,N_41608);
or U49863 (N_49863,N_43206,N_41262);
or U49864 (N_49864,N_44953,N_43991);
xor U49865 (N_49865,N_41774,N_43958);
or U49866 (N_49866,N_43243,N_42563);
nor U49867 (N_49867,N_43224,N_43082);
nand U49868 (N_49868,N_41985,N_42877);
nand U49869 (N_49869,N_42126,N_43975);
and U49870 (N_49870,N_43443,N_43977);
nor U49871 (N_49871,N_41091,N_42268);
or U49872 (N_49872,N_40845,N_41938);
nor U49873 (N_49873,N_44081,N_40291);
xor U49874 (N_49874,N_41459,N_41477);
nand U49875 (N_49875,N_42930,N_40497);
xnor U49876 (N_49876,N_44125,N_44209);
nor U49877 (N_49877,N_40171,N_43077);
nand U49878 (N_49878,N_42363,N_41115);
or U49879 (N_49879,N_42839,N_42006);
nor U49880 (N_49880,N_41308,N_43173);
xnor U49881 (N_49881,N_44115,N_44706);
and U49882 (N_49882,N_43489,N_43775);
and U49883 (N_49883,N_40630,N_42226);
nor U49884 (N_49884,N_43625,N_41742);
and U49885 (N_49885,N_44785,N_43762);
or U49886 (N_49886,N_41041,N_42924);
and U49887 (N_49887,N_40228,N_41596);
xnor U49888 (N_49888,N_40467,N_43058);
nand U49889 (N_49889,N_40301,N_43043);
and U49890 (N_49890,N_44811,N_43242);
and U49891 (N_49891,N_44049,N_40915);
and U49892 (N_49892,N_42549,N_44730);
xnor U49893 (N_49893,N_43983,N_43825);
or U49894 (N_49894,N_44305,N_42529);
nand U49895 (N_49895,N_40770,N_41992);
or U49896 (N_49896,N_40183,N_40957);
xor U49897 (N_49897,N_43980,N_44230);
and U49898 (N_49898,N_42979,N_41247);
nor U49899 (N_49899,N_43626,N_40361);
or U49900 (N_49900,N_42620,N_41082);
xor U49901 (N_49901,N_40781,N_43021);
nand U49902 (N_49902,N_44636,N_42294);
and U49903 (N_49903,N_42287,N_40803);
and U49904 (N_49904,N_41049,N_43588);
xnor U49905 (N_49905,N_41524,N_43815);
or U49906 (N_49906,N_41145,N_41021);
nor U49907 (N_49907,N_43582,N_43792);
nor U49908 (N_49908,N_42699,N_40473);
or U49909 (N_49909,N_44194,N_40620);
xnor U49910 (N_49910,N_43211,N_42820);
nand U49911 (N_49911,N_42602,N_44328);
nor U49912 (N_49912,N_40284,N_41906);
nor U49913 (N_49913,N_40615,N_41510);
nand U49914 (N_49914,N_44851,N_40856);
xnor U49915 (N_49915,N_42452,N_40296);
xor U49916 (N_49916,N_41250,N_44380);
nand U49917 (N_49917,N_43832,N_41670);
or U49918 (N_49918,N_43494,N_40836);
or U49919 (N_49919,N_44827,N_44060);
nor U49920 (N_49920,N_40345,N_42919);
nand U49921 (N_49921,N_42416,N_43761);
nand U49922 (N_49922,N_43654,N_40612);
or U49923 (N_49923,N_43092,N_43708);
nor U49924 (N_49924,N_41805,N_41087);
nor U49925 (N_49925,N_40797,N_40019);
nand U49926 (N_49926,N_42082,N_43522);
nor U49927 (N_49927,N_41267,N_40377);
nand U49928 (N_49928,N_44303,N_41960);
xnor U49929 (N_49929,N_43528,N_42512);
or U49930 (N_49930,N_41746,N_40318);
nand U49931 (N_49931,N_44628,N_44631);
nor U49932 (N_49932,N_42882,N_43902);
nand U49933 (N_49933,N_42709,N_40434);
and U49934 (N_49934,N_43655,N_43388);
or U49935 (N_49935,N_43199,N_41254);
or U49936 (N_49936,N_43610,N_42608);
xnor U49937 (N_49937,N_41347,N_43805);
or U49938 (N_49938,N_43388,N_44545);
nor U49939 (N_49939,N_43926,N_44849);
nor U49940 (N_49940,N_42031,N_41603);
nor U49941 (N_49941,N_40685,N_42841);
nor U49942 (N_49942,N_44775,N_40469);
nor U49943 (N_49943,N_43116,N_41408);
nand U49944 (N_49944,N_41832,N_41426);
nand U49945 (N_49945,N_42499,N_44422);
and U49946 (N_49946,N_40260,N_43380);
xor U49947 (N_49947,N_42512,N_41887);
and U49948 (N_49948,N_43818,N_43847);
and U49949 (N_49949,N_43756,N_43955);
nor U49950 (N_49950,N_42289,N_41705);
xnor U49951 (N_49951,N_42966,N_42898);
xor U49952 (N_49952,N_43648,N_42573);
xnor U49953 (N_49953,N_40082,N_44005);
nand U49954 (N_49954,N_44816,N_40769);
xnor U49955 (N_49955,N_42313,N_42461);
nand U49956 (N_49956,N_42837,N_42136);
and U49957 (N_49957,N_42602,N_42458);
or U49958 (N_49958,N_42766,N_43435);
xnor U49959 (N_49959,N_44858,N_44516);
nor U49960 (N_49960,N_40024,N_41972);
xor U49961 (N_49961,N_44512,N_42062);
or U49962 (N_49962,N_44027,N_41838);
nor U49963 (N_49963,N_43854,N_42547);
nor U49964 (N_49964,N_41803,N_41146);
or U49965 (N_49965,N_41071,N_42589);
and U49966 (N_49966,N_40418,N_42336);
or U49967 (N_49967,N_40499,N_43267);
or U49968 (N_49968,N_43203,N_42620);
or U49969 (N_49969,N_43507,N_42913);
and U49970 (N_49970,N_42947,N_43312);
xor U49971 (N_49971,N_40427,N_40557);
xnor U49972 (N_49972,N_43018,N_40318);
and U49973 (N_49973,N_40137,N_41866);
nand U49974 (N_49974,N_41921,N_41752);
xnor U49975 (N_49975,N_42984,N_42032);
nor U49976 (N_49976,N_41411,N_41524);
or U49977 (N_49977,N_44556,N_42807);
nand U49978 (N_49978,N_40070,N_41405);
nor U49979 (N_49979,N_42127,N_40928);
or U49980 (N_49980,N_40572,N_44663);
and U49981 (N_49981,N_41242,N_40340);
nor U49982 (N_49982,N_43065,N_43460);
or U49983 (N_49983,N_40635,N_43946);
nor U49984 (N_49984,N_40929,N_40528);
nand U49985 (N_49985,N_40747,N_44121);
or U49986 (N_49986,N_42277,N_42136);
nor U49987 (N_49987,N_44479,N_43362);
nor U49988 (N_49988,N_41595,N_43307);
nand U49989 (N_49989,N_43825,N_41473);
nand U49990 (N_49990,N_42618,N_41784);
and U49991 (N_49991,N_43765,N_41197);
and U49992 (N_49992,N_42325,N_42701);
and U49993 (N_49993,N_42344,N_44873);
nor U49994 (N_49994,N_43121,N_41927);
nand U49995 (N_49995,N_43070,N_43578);
nor U49996 (N_49996,N_42885,N_41672);
nand U49997 (N_49997,N_43304,N_42120);
xnor U49998 (N_49998,N_42839,N_41779);
or U49999 (N_49999,N_40598,N_43123);
nand UO_0 (O_0,N_49826,N_48179);
nor UO_1 (O_1,N_45659,N_49457);
and UO_2 (O_2,N_49126,N_48066);
nand UO_3 (O_3,N_45926,N_47733);
or UO_4 (O_4,N_49767,N_48198);
xnor UO_5 (O_5,N_46045,N_49583);
nand UO_6 (O_6,N_48804,N_45903);
xnor UO_7 (O_7,N_46665,N_46845);
and UO_8 (O_8,N_47462,N_47245);
nor UO_9 (O_9,N_47119,N_49269);
nand UO_10 (O_10,N_48313,N_49213);
nor UO_11 (O_11,N_49756,N_49891);
nor UO_12 (O_12,N_49452,N_46316);
nor UO_13 (O_13,N_45218,N_47173);
or UO_14 (O_14,N_47018,N_47107);
xor UO_15 (O_15,N_46213,N_48797);
xor UO_16 (O_16,N_46044,N_45933);
xnor UO_17 (O_17,N_48594,N_45617);
or UO_18 (O_18,N_49752,N_49405);
and UO_19 (O_19,N_47112,N_47265);
nor UO_20 (O_20,N_49784,N_46298);
or UO_21 (O_21,N_49289,N_46438);
and UO_22 (O_22,N_47717,N_48139);
and UO_23 (O_23,N_49194,N_45840);
or UO_24 (O_24,N_47358,N_46839);
xnor UO_25 (O_25,N_49399,N_47642);
nor UO_26 (O_26,N_49462,N_45458);
or UO_27 (O_27,N_45862,N_47384);
nand UO_28 (O_28,N_48523,N_45615);
nor UO_29 (O_29,N_49667,N_46687);
nor UO_30 (O_30,N_49203,N_45054);
and UO_31 (O_31,N_48688,N_48210);
or UO_32 (O_32,N_49656,N_49993);
or UO_33 (O_33,N_48989,N_45268);
xor UO_34 (O_34,N_49035,N_45121);
or UO_35 (O_35,N_49716,N_49815);
nor UO_36 (O_36,N_45632,N_49950);
or UO_37 (O_37,N_46307,N_49897);
and UO_38 (O_38,N_47643,N_47758);
nand UO_39 (O_39,N_45868,N_46804);
nand UO_40 (O_40,N_49751,N_48143);
nand UO_41 (O_41,N_46155,N_45485);
nand UO_42 (O_42,N_48228,N_47007);
nor UO_43 (O_43,N_48647,N_46874);
nand UO_44 (O_44,N_45379,N_49532);
nor UO_45 (O_45,N_46176,N_45106);
and UO_46 (O_46,N_49140,N_46476);
xor UO_47 (O_47,N_46056,N_47985);
or UO_48 (O_48,N_45854,N_48110);
or UO_49 (O_49,N_49416,N_48632);
xnor UO_50 (O_50,N_45859,N_47676);
and UO_51 (O_51,N_47454,N_48518);
and UO_52 (O_52,N_46009,N_46581);
nand UO_53 (O_53,N_47631,N_49317);
or UO_54 (O_54,N_45896,N_45332);
xnor UO_55 (O_55,N_47593,N_46382);
or UO_56 (O_56,N_48664,N_47945);
and UO_57 (O_57,N_47000,N_46290);
nor UO_58 (O_58,N_48042,N_48165);
xnor UO_59 (O_59,N_48814,N_45735);
and UO_60 (O_60,N_49649,N_48779);
or UO_61 (O_61,N_47276,N_46684);
nor UO_62 (O_62,N_49338,N_48187);
nand UO_63 (O_63,N_46512,N_47486);
nand UO_64 (O_64,N_46251,N_46221);
nand UO_65 (O_65,N_47074,N_48729);
and UO_66 (O_66,N_47139,N_49446);
or UO_67 (O_67,N_45114,N_47960);
xor UO_68 (O_68,N_48233,N_47175);
and UO_69 (O_69,N_46423,N_47669);
nor UO_70 (O_70,N_45845,N_48425);
xnor UO_71 (O_71,N_48996,N_46784);
or UO_72 (O_72,N_45119,N_47162);
xor UO_73 (O_73,N_45810,N_47288);
or UO_74 (O_74,N_45522,N_45222);
and UO_75 (O_75,N_45390,N_48158);
or UO_76 (O_76,N_48380,N_48938);
or UO_77 (O_77,N_48090,N_48633);
nand UO_78 (O_78,N_47863,N_47239);
nor UO_79 (O_79,N_48086,N_48089);
nand UO_80 (O_80,N_45653,N_46544);
xor UO_81 (O_81,N_46878,N_45076);
xor UO_82 (O_82,N_48004,N_47929);
xor UO_83 (O_83,N_45642,N_46773);
xnor UO_84 (O_84,N_47168,N_49620);
or UO_85 (O_85,N_49877,N_48604);
and UO_86 (O_86,N_45606,N_47195);
and UO_87 (O_87,N_48893,N_45831);
nand UO_88 (O_88,N_48911,N_46108);
nand UO_89 (O_89,N_48457,N_46707);
or UO_90 (O_90,N_49166,N_46922);
xnor UO_91 (O_91,N_46623,N_48474);
nand UO_92 (O_92,N_45534,N_47321);
or UO_93 (O_93,N_47295,N_46182);
or UO_94 (O_94,N_46337,N_47138);
nor UO_95 (O_95,N_46153,N_46796);
nor UO_96 (O_96,N_47957,N_48643);
and UO_97 (O_97,N_47774,N_46209);
or UO_98 (O_98,N_45329,N_46724);
nand UO_99 (O_99,N_46670,N_48451);
and UO_100 (O_100,N_45988,N_46865);
and UO_101 (O_101,N_45134,N_49287);
and UO_102 (O_102,N_47932,N_46779);
xor UO_103 (O_103,N_46013,N_45791);
nand UO_104 (O_104,N_45957,N_49415);
nand UO_105 (O_105,N_47330,N_47867);
or UO_106 (O_106,N_46694,N_49308);
xnor UO_107 (O_107,N_46095,N_45045);
xor UO_108 (O_108,N_46855,N_48377);
or UO_109 (O_109,N_45296,N_46094);
nor UO_110 (O_110,N_49169,N_46727);
or UO_111 (O_111,N_48258,N_48416);
or UO_112 (O_112,N_49930,N_49316);
and UO_113 (O_113,N_49661,N_49185);
and UO_114 (O_114,N_48917,N_47645);
and UO_115 (O_115,N_45161,N_49643);
xor UO_116 (O_116,N_47061,N_48391);
nor UO_117 (O_117,N_45473,N_48326);
and UO_118 (O_118,N_47102,N_49600);
nor UO_119 (O_119,N_45984,N_49932);
nor UO_120 (O_120,N_45302,N_49569);
nor UO_121 (O_121,N_46989,N_45729);
nor UO_122 (O_122,N_49113,N_49513);
or UO_123 (O_123,N_46149,N_47280);
or UO_124 (O_124,N_45384,N_48556);
and UO_125 (O_125,N_45861,N_48307);
xnor UO_126 (O_126,N_46870,N_47810);
nor UO_127 (O_127,N_47686,N_46543);
nor UO_128 (O_128,N_46477,N_47011);
or UO_129 (O_129,N_45030,N_46730);
and UO_130 (O_130,N_45915,N_48168);
nor UO_131 (O_131,N_45551,N_47681);
nor UO_132 (O_132,N_47445,N_45187);
or UO_133 (O_133,N_46763,N_45238);
or UO_134 (O_134,N_49760,N_45955);
nor UO_135 (O_135,N_48201,N_49451);
nand UO_136 (O_136,N_45630,N_46043);
or UO_137 (O_137,N_48075,N_48622);
xnor UO_138 (O_138,N_47047,N_47213);
and UO_139 (O_139,N_47339,N_48417);
nand UO_140 (O_140,N_49615,N_47996);
nand UO_141 (O_141,N_48148,N_45746);
xor UO_142 (O_142,N_45479,N_45705);
nand UO_143 (O_143,N_45837,N_46921);
xnor UO_144 (O_144,N_47036,N_45597);
nand UO_145 (O_145,N_46516,N_47380);
xnor UO_146 (O_146,N_47037,N_49910);
nand UO_147 (O_147,N_47582,N_47842);
or UO_148 (O_148,N_47221,N_47357);
nand UO_149 (O_149,N_49020,N_46720);
xor UO_150 (O_150,N_49913,N_45503);
and UO_151 (O_151,N_47950,N_48299);
or UO_152 (O_152,N_45511,N_49616);
xnor UO_153 (O_153,N_46433,N_46678);
xor UO_154 (O_154,N_47560,N_45252);
nand UO_155 (O_155,N_46985,N_46708);
and UO_156 (O_156,N_48085,N_47746);
xor UO_157 (O_157,N_46428,N_47506);
nor UO_158 (O_158,N_48027,N_48792);
or UO_159 (O_159,N_49742,N_46160);
xor UO_160 (O_160,N_47255,N_49801);
nor UO_161 (O_161,N_49201,N_46862);
nor UO_162 (O_162,N_47496,N_48968);
xnor UO_163 (O_163,N_48964,N_46047);
and UO_164 (O_164,N_49714,N_46229);
nand UO_165 (O_165,N_47680,N_46584);
nor UO_166 (O_166,N_46527,N_45707);
nor UO_167 (O_167,N_46318,N_48428);
xnor UO_168 (O_168,N_46256,N_47369);
and UO_169 (O_169,N_48221,N_47527);
xnor UO_170 (O_170,N_47250,N_49633);
and UO_171 (O_171,N_46585,N_45088);
nand UO_172 (O_172,N_49484,N_45279);
and UO_173 (O_173,N_48668,N_45805);
and UO_174 (O_174,N_45870,N_46202);
and UO_175 (O_175,N_46242,N_45936);
nand UO_176 (O_176,N_46051,N_48094);
nor UO_177 (O_177,N_46347,N_48656);
nand UO_178 (O_178,N_46192,N_49432);
nand UO_179 (O_179,N_48419,N_46188);
or UO_180 (O_180,N_49110,N_45658);
and UO_181 (O_181,N_47703,N_48961);
or UO_182 (O_182,N_47936,N_45894);
and UO_183 (O_183,N_46911,N_47001);
xor UO_184 (O_184,N_45600,N_46780);
and UO_185 (O_185,N_47855,N_47508);
nor UO_186 (O_186,N_49837,N_47032);
nand UO_187 (O_187,N_48871,N_48510);
or UO_188 (O_188,N_48734,N_46212);
nand UO_189 (O_189,N_47944,N_46731);
and UO_190 (O_190,N_48883,N_47572);
nor UO_191 (O_191,N_49172,N_46937);
nor UO_192 (O_192,N_45257,N_49739);
xor UO_193 (O_193,N_46394,N_49027);
and UO_194 (O_194,N_48981,N_48300);
xor UO_195 (O_195,N_45507,N_48872);
nor UO_196 (O_196,N_46031,N_47870);
nor UO_197 (O_197,N_47305,N_45717);
nor UO_198 (O_198,N_49453,N_48152);
xnor UO_199 (O_199,N_46408,N_46480);
nand UO_200 (O_200,N_48714,N_49629);
or UO_201 (O_201,N_48584,N_46627);
or UO_202 (O_202,N_47115,N_46513);
or UO_203 (O_203,N_47164,N_49847);
and UO_204 (O_204,N_47992,N_49850);
nor UO_205 (O_205,N_49222,N_45715);
or UO_206 (O_206,N_45993,N_45335);
nand UO_207 (O_207,N_46181,N_49054);
xor UO_208 (O_208,N_45569,N_45244);
or UO_209 (O_209,N_49449,N_47955);
nor UO_210 (O_210,N_48050,N_46161);
nor UO_211 (O_211,N_46086,N_45945);
and UO_212 (O_212,N_47298,N_48954);
or UO_213 (O_213,N_45447,N_45607);
xor UO_214 (O_214,N_49480,N_49087);
nor UO_215 (O_215,N_49732,N_46603);
nand UO_216 (O_216,N_49147,N_49744);
xnor UO_217 (O_217,N_47283,N_47264);
xnor UO_218 (O_218,N_46424,N_47878);
nor UO_219 (O_219,N_46853,N_45970);
nor UO_220 (O_220,N_45820,N_46484);
xor UO_221 (O_221,N_48172,N_46661);
or UO_222 (O_222,N_45145,N_48985);
nor UO_223 (O_223,N_46065,N_46866);
or UO_224 (O_224,N_48645,N_49114);
nor UO_225 (O_225,N_48574,N_45764);
xor UO_226 (O_226,N_48421,N_45528);
nand UO_227 (O_227,N_46082,N_49889);
nand UO_228 (O_228,N_47328,N_46285);
nand UO_229 (O_229,N_47601,N_48735);
nor UO_230 (O_230,N_46036,N_46361);
xnor UO_231 (O_231,N_48061,N_45713);
nor UO_232 (O_232,N_45526,N_47236);
xor UO_233 (O_233,N_49556,N_46322);
nand UO_234 (O_234,N_46452,N_46474);
or UO_235 (O_235,N_48799,N_48011);
or UO_236 (O_236,N_49790,N_48612);
and UO_237 (O_237,N_45835,N_49506);
or UO_238 (O_238,N_49275,N_45014);
and UO_239 (O_239,N_49696,N_48998);
and UO_240 (O_240,N_48199,N_49663);
xor UO_241 (O_241,N_47148,N_46446);
nand UO_242 (O_242,N_46370,N_48738);
or UO_243 (O_243,N_48940,N_47772);
nand UO_244 (O_244,N_46122,N_49386);
nand UO_245 (O_245,N_47602,N_47982);
nor UO_246 (O_246,N_45804,N_49785);
nand UO_247 (O_247,N_48277,N_47006);
and UO_248 (O_248,N_46799,N_49797);
nor UO_249 (O_249,N_46397,N_48443);
or UO_250 (O_250,N_47394,N_48679);
nor UO_251 (O_251,N_46028,N_45246);
or UO_252 (O_252,N_49501,N_45881);
nor UO_253 (O_253,N_49012,N_45683);
xnor UO_254 (O_254,N_49987,N_48121);
and UO_255 (O_255,N_46055,N_46239);
nand UO_256 (O_256,N_48392,N_45101);
and UO_257 (O_257,N_46765,N_49563);
nand UO_258 (O_258,N_45934,N_49566);
or UO_259 (O_259,N_48430,N_49922);
and UO_260 (O_260,N_48945,N_45732);
and UO_261 (O_261,N_47463,N_46310);
nor UO_262 (O_262,N_45093,N_46909);
or UO_263 (O_263,N_48810,N_46733);
nand UO_264 (O_264,N_49156,N_47637);
and UO_265 (O_265,N_45586,N_49969);
xnor UO_266 (O_266,N_45053,N_48155);
xnor UO_267 (O_267,N_48213,N_48133);
xnor UO_268 (O_268,N_49880,N_46455);
xor UO_269 (O_269,N_47923,N_46295);
nor UO_270 (O_270,N_46263,N_49435);
nor UO_271 (O_271,N_49261,N_46217);
or UO_272 (O_272,N_47478,N_49832);
or UO_273 (O_273,N_48189,N_47990);
and UO_274 (O_274,N_47086,N_46454);
or UO_275 (O_275,N_49456,N_45353);
xnor UO_276 (O_276,N_49691,N_48296);
nand UO_277 (O_277,N_45583,N_48209);
nor UO_278 (O_278,N_47302,N_48589);
nand UO_279 (O_279,N_46861,N_46660);
and UO_280 (O_280,N_47015,N_46432);
and UO_281 (O_281,N_47169,N_49438);
or UO_282 (O_282,N_45577,N_46333);
xnor UO_283 (O_283,N_48867,N_47779);
or UO_284 (O_284,N_49843,N_49772);
xnor UO_285 (O_285,N_49690,N_49344);
and UO_286 (O_286,N_48608,N_46672);
xnor UO_287 (O_287,N_48730,N_46133);
nor UO_288 (O_288,N_46726,N_48422);
nor UO_289 (O_289,N_47233,N_49614);
xnor UO_290 (O_290,N_45463,N_47579);
xnor UO_291 (O_291,N_47180,N_49659);
and UO_292 (O_292,N_49581,N_48640);
xor UO_293 (O_293,N_47004,N_45902);
nor UO_294 (O_294,N_49589,N_46167);
nand UO_295 (O_295,N_49018,N_46848);
xor UO_296 (O_296,N_48924,N_47296);
or UO_297 (O_297,N_49793,N_48111);
xnor UO_298 (O_298,N_45057,N_45456);
and UO_299 (O_299,N_45790,N_46963);
and UO_300 (O_300,N_47675,N_49250);
nand UO_301 (O_301,N_49009,N_49887);
nand UO_302 (O_302,N_49398,N_46426);
or UO_303 (O_303,N_45263,N_48698);
nor UO_304 (O_304,N_46425,N_48910);
and UO_305 (O_305,N_49498,N_49901);
nor UO_306 (O_306,N_46901,N_46150);
nor UO_307 (O_307,N_46884,N_45611);
and UO_308 (O_308,N_45289,N_48769);
nand UO_309 (O_309,N_48102,N_49726);
nand UO_310 (O_310,N_48146,N_49144);
xor UO_311 (O_311,N_48483,N_49091);
and UO_312 (O_312,N_47728,N_48896);
xor UO_313 (O_313,N_48588,N_46350);
nand UO_314 (O_314,N_48358,N_49665);
nand UO_315 (O_315,N_46891,N_47204);
nor UO_316 (O_316,N_45514,N_46483);
and UO_317 (O_317,N_49619,N_48934);
and UO_318 (O_318,N_46001,N_47128);
xor UO_319 (O_319,N_49345,N_46388);
nor UO_320 (O_320,N_48344,N_48752);
xnor UO_321 (O_321,N_49911,N_47625);
nor UO_322 (O_322,N_45159,N_49187);
xor UO_323 (O_323,N_49285,N_45216);
and UO_324 (O_324,N_47644,N_48054);
xor UO_325 (O_325,N_49764,N_45085);
nand UO_326 (O_326,N_45667,N_48237);
or UO_327 (O_327,N_49208,N_48508);
or UO_328 (O_328,N_46187,N_45095);
or UO_329 (O_329,N_48543,N_45852);
nand UO_330 (O_330,N_46523,N_49291);
xnor UO_331 (O_331,N_48409,N_47567);
nor UO_332 (O_332,N_47576,N_47721);
nand UO_333 (O_333,N_46649,N_45294);
nand UO_334 (O_334,N_46243,N_45982);
nand UO_335 (O_335,N_48778,N_49970);
xnor UO_336 (O_336,N_47095,N_48573);
or UO_337 (O_337,N_49391,N_46556);
and UO_338 (O_338,N_49924,N_47971);
nand UO_339 (O_339,N_49318,N_45373);
xnor UO_340 (O_340,N_45130,N_49990);
xor UO_341 (O_341,N_47135,N_49768);
xor UO_342 (O_342,N_45442,N_48274);
or UO_343 (O_343,N_49682,N_49870);
nor UO_344 (O_344,N_46999,N_47909);
nor UO_345 (O_345,N_47624,N_45318);
nand UO_346 (O_346,N_46920,N_49786);
and UO_347 (O_347,N_47161,N_47140);
and UO_348 (O_348,N_49999,N_45519);
or UO_349 (O_349,N_47869,N_49834);
xnor UO_350 (O_350,N_46936,N_47038);
nand UO_351 (O_351,N_48545,N_47317);
xnor UO_352 (O_352,N_48957,N_47411);
or UO_353 (O_353,N_48292,N_49628);
xnor UO_354 (O_354,N_46608,N_47356);
and UO_355 (O_355,N_48290,N_48047);
nand UO_356 (O_356,N_45531,N_49996);
or UO_357 (O_357,N_45338,N_45916);
and UO_358 (O_358,N_45151,N_49976);
or UO_359 (O_359,N_46000,N_48639);
or UO_360 (O_360,N_49789,N_48332);
or UO_361 (O_361,N_45662,N_48712);
or UO_362 (O_362,N_47552,N_49518);
xor UO_363 (O_363,N_47663,N_49251);
xnor UO_364 (O_364,N_45111,N_49550);
or UO_365 (O_365,N_48157,N_49298);
or UO_366 (O_366,N_49542,N_46787);
or UO_367 (O_367,N_46732,N_45616);
or UO_368 (O_368,N_47816,N_49640);
nand UO_369 (O_369,N_48696,N_46038);
nand UO_370 (O_370,N_46084,N_45722);
xor UO_371 (O_371,N_48915,N_49270);
nor UO_372 (O_372,N_45529,N_48306);
nor UO_373 (O_373,N_45675,N_49598);
or UO_374 (O_374,N_45265,N_45459);
nor UO_375 (O_375,N_49050,N_47226);
xnor UO_376 (O_376,N_45360,N_49743);
nor UO_377 (O_377,N_45419,N_47791);
nor UO_378 (O_378,N_47654,N_48958);
and UO_379 (O_379,N_46782,N_49070);
and UO_380 (O_380,N_45719,N_46379);
or UO_381 (O_381,N_45486,N_47474);
nor UO_382 (O_382,N_46117,N_47777);
nand UO_383 (O_383,N_49197,N_48141);
nand UO_384 (O_384,N_46274,N_47685);
or UO_385 (O_385,N_47535,N_46300);
nand UO_386 (O_386,N_47993,N_48808);
nor UO_387 (O_387,N_49502,N_47071);
xor UO_388 (O_388,N_48197,N_49671);
xnor UO_389 (O_389,N_47212,N_46561);
and UO_390 (O_390,N_46566,N_49938);
nor UO_391 (O_391,N_46498,N_45762);
or UO_392 (O_392,N_48845,N_45846);
nor UO_393 (O_393,N_45636,N_47215);
nor UO_394 (O_394,N_46233,N_48777);
nand UO_395 (O_395,N_47913,N_48445);
nand UO_396 (O_396,N_46783,N_46745);
nand UO_397 (O_397,N_48458,N_46048);
or UO_398 (O_398,N_48950,N_47067);
xnor UO_399 (O_399,N_47900,N_45770);
nor UO_400 (O_400,N_45598,N_46974);
xnor UO_401 (O_401,N_48101,N_48580);
and UO_402 (O_402,N_46385,N_45201);
or UO_403 (O_403,N_48657,N_47958);
xnor UO_404 (O_404,N_48269,N_48394);
or UO_405 (O_405,N_46450,N_47041);
xnor UO_406 (O_406,N_46528,N_48120);
nand UO_407 (O_407,N_48174,N_45367);
and UO_408 (O_408,N_45680,N_48407);
or UO_409 (O_409,N_46296,N_48878);
nor UO_410 (O_410,N_47801,N_46882);
and UO_411 (O_411,N_45242,N_47235);
nand UO_412 (O_412,N_48951,N_49262);
and UO_413 (O_413,N_49748,N_46435);
or UO_414 (O_414,N_49408,N_49676);
nand UO_415 (O_415,N_45580,N_45376);
or UO_416 (O_416,N_49830,N_49707);
xnor UO_417 (O_417,N_45566,N_45863);
xnor UO_418 (O_418,N_45104,N_49572);
xnor UO_419 (O_419,N_47359,N_48454);
xnor UO_420 (O_420,N_46099,N_48974);
xor UO_421 (O_421,N_49783,N_45195);
xnor UO_422 (O_422,N_46738,N_47124);
xnor UO_423 (O_423,N_45608,N_49662);
xor UO_424 (O_424,N_45260,N_49603);
nor UO_425 (O_425,N_46511,N_47223);
nor UO_426 (O_426,N_46786,N_48150);
xor UO_427 (O_427,N_47492,N_48927);
xor UO_428 (O_428,N_46616,N_48809);
xor UO_429 (O_429,N_47066,N_47117);
and UO_430 (O_430,N_49584,N_47729);
nand UO_431 (O_431,N_45967,N_46264);
nand UO_432 (O_432,N_45372,N_45807);
and UO_433 (O_433,N_49529,N_48859);
and UO_434 (O_434,N_46923,N_45559);
nor UO_435 (O_435,N_45467,N_45427);
nor UO_436 (O_436,N_49454,N_49097);
nand UO_437 (O_437,N_45004,N_49141);
xor UO_438 (O_438,N_47129,N_47403);
xnor UO_439 (O_439,N_46464,N_46342);
and UO_440 (O_440,N_48721,N_45020);
nor UO_441 (O_441,N_49302,N_46916);
nor UO_442 (O_442,N_45696,N_45167);
nand UO_443 (O_443,N_46359,N_47546);
nor UO_444 (O_444,N_46828,N_49129);
or UO_445 (O_445,N_48904,N_49425);
nor UO_446 (O_446,N_48798,N_48281);
or UO_447 (O_447,N_48827,N_47838);
and UO_448 (O_448,N_46026,N_45987);
and UO_449 (O_449,N_47077,N_46163);
xor UO_450 (O_450,N_46795,N_45385);
xor UO_451 (O_451,N_49625,N_48742);
and UO_452 (O_452,N_49003,N_48325);
nor UO_453 (O_453,N_48373,N_46472);
nor UO_454 (O_454,N_46743,N_46170);
xnor UO_455 (O_455,N_49822,N_47400);
or UO_456 (O_456,N_46218,N_45251);
nand UO_457 (O_457,N_47823,N_47827);
nand UO_458 (O_458,N_45833,N_46068);
nand UO_459 (O_459,N_49862,N_46418);
nand UO_460 (O_460,N_48252,N_47182);
nand UO_461 (O_461,N_48317,N_45368);
nor UO_462 (O_462,N_49746,N_46789);
nand UO_463 (O_463,N_49409,N_45788);
nand UO_464 (O_464,N_48737,N_49694);
nand UO_465 (O_465,N_49986,N_46353);
xnor UO_466 (O_466,N_47687,N_46412);
nor UO_467 (O_467,N_49701,N_48944);
nand UO_468 (O_468,N_45978,N_48504);
or UO_469 (O_469,N_47988,N_45708);
xor UO_470 (O_470,N_45858,N_46441);
nand UO_471 (O_471,N_49072,N_47487);
nand UO_472 (O_472,N_45766,N_45871);
nor UO_473 (O_473,N_47354,N_45392);
xnor UO_474 (O_474,N_49787,N_49387);
nand UO_475 (O_475,N_47632,N_48920);
nor UO_476 (O_476,N_48115,N_47500);
xor UO_477 (O_477,N_49375,N_47690);
and UO_478 (O_478,N_49535,N_46635);
xnor UO_479 (O_479,N_45402,N_47565);
or UO_480 (O_480,N_48449,N_48936);
nand UO_481 (O_481,N_49153,N_46716);
nand UO_482 (O_482,N_49668,N_48057);
nand UO_483 (O_483,N_46626,N_47421);
nand UO_484 (O_484,N_49892,N_48558);
and UO_485 (O_485,N_46179,N_47234);
or UO_486 (O_486,N_47639,N_46816);
nand UO_487 (O_487,N_46377,N_46685);
and UO_488 (O_488,N_46625,N_45352);
nand UO_489 (O_489,N_46840,N_46565);
nand UO_490 (O_490,N_46396,N_47415);
nand UO_491 (O_491,N_45750,N_46368);
and UO_492 (O_492,N_49921,N_49234);
xnor UO_493 (O_493,N_45783,N_48024);
nor UO_494 (O_494,N_45823,N_48966);
nor UO_495 (O_495,N_48821,N_48720);
and UO_496 (O_496,N_45530,N_49216);
xnor UO_497 (O_497,N_49492,N_46293);
or UO_498 (O_498,N_45999,N_49695);
nand UO_499 (O_499,N_47844,N_48396);
xnor UO_500 (O_500,N_47748,N_49490);
and UO_501 (O_501,N_49228,N_49046);
xnor UO_502 (O_502,N_46138,N_46468);
nor UO_503 (O_503,N_48685,N_49105);
xor UO_504 (O_504,N_47641,N_48666);
xor UO_505 (O_505,N_47216,N_45585);
nand UO_506 (O_506,N_48820,N_49115);
and UO_507 (O_507,N_49045,N_49039);
nor UO_508 (O_508,N_47068,N_48464);
nand UO_509 (O_509,N_45545,N_45744);
or UO_510 (O_510,N_47407,N_48592);
or UO_511 (O_511,N_47338,N_49749);
nand UO_512 (O_512,N_49127,N_48818);
or UO_513 (O_513,N_47436,N_45283);
xor UO_514 (O_514,N_49758,N_48901);
nand UO_515 (O_515,N_46029,N_48716);
or UO_516 (O_516,N_49680,N_45181);
and UO_517 (O_517,N_47617,N_48505);
and UO_518 (O_518,N_49444,N_46096);
and UO_519 (O_519,N_47587,N_47160);
or UO_520 (O_520,N_47274,N_47891);
and UO_521 (O_521,N_49624,N_45880);
and UO_522 (O_522,N_49099,N_47513);
nor UO_523 (O_523,N_48908,N_45886);
and UO_524 (O_524,N_46115,N_46815);
xnor UO_525 (O_525,N_47270,N_46387);
and UO_526 (O_526,N_47299,N_47123);
and UO_527 (O_527,N_49562,N_48889);
or UO_528 (O_528,N_49521,N_45295);
nor UO_529 (O_529,N_45200,N_47051);
xor UO_530 (O_530,N_47151,N_45068);
or UO_531 (O_531,N_46510,N_47318);
and UO_532 (O_532,N_48613,N_46534);
xnor UO_533 (O_533,N_46760,N_49303);
or UO_534 (O_534,N_48866,N_45375);
nor UO_535 (O_535,N_48286,N_45927);
xnor UO_536 (O_536,N_47155,N_48191);
or UO_537 (O_537,N_46837,N_49981);
and UO_538 (O_538,N_47453,N_47271);
and UO_539 (O_539,N_47704,N_48978);
xnor UO_540 (O_540,N_49833,N_45188);
or UO_541 (O_541,N_48395,N_47708);
or UO_542 (O_542,N_46302,N_48276);
or UO_543 (O_543,N_48975,N_45782);
xnor UO_544 (O_544,N_48776,N_49090);
nor UO_545 (O_545,N_45194,N_45391);
nand UO_546 (O_546,N_47145,N_47266);
or UO_547 (O_547,N_45543,N_47635);
xor UO_548 (O_548,N_49098,N_45796);
nor UO_549 (O_549,N_45098,N_46663);
xor UO_550 (O_550,N_47883,N_48060);
nand UO_551 (O_551,N_48811,N_45909);
or UO_552 (O_552,N_49814,N_48405);
and UO_553 (O_553,N_48329,N_45677);
nand UO_554 (O_554,N_49259,N_46391);
nor UO_555 (O_555,N_49652,N_46895);
xnor UO_556 (O_556,N_46539,N_48648);
nor UO_557 (O_557,N_47987,N_46535);
or UO_558 (O_558,N_47840,N_46466);
nand UO_559 (O_559,N_45142,N_49230);
nand UO_560 (O_560,N_48650,N_47315);
or UO_561 (O_561,N_46244,N_47497);
and UO_562 (O_562,N_47304,N_49552);
and UO_563 (O_563,N_48841,N_48379);
and UO_564 (O_564,N_47079,N_46682);
and UO_565 (O_565,N_46019,N_49106);
nand UO_566 (O_566,N_45760,N_46818);
or UO_567 (O_567,N_47947,N_46317);
xnor UO_568 (O_568,N_45092,N_49470);
nor UO_569 (O_569,N_47633,N_46766);
or UO_570 (O_570,N_49806,N_45966);
or UO_571 (O_571,N_48916,N_46972);
or UO_572 (O_572,N_49182,N_48244);
and UO_573 (O_573,N_46113,N_45147);
nand UO_574 (O_574,N_46223,N_45414);
xnor UO_575 (O_575,N_49985,N_48794);
or UO_576 (O_576,N_46607,N_48138);
or UO_577 (O_577,N_45899,N_45929);
nand UO_578 (O_578,N_47043,N_45964);
nor UO_579 (O_579,N_47677,N_46487);
or UO_580 (O_580,N_46058,N_48970);
nor UO_581 (O_581,N_46140,N_48440);
nand UO_582 (O_582,N_48823,N_48994);
nand UO_583 (O_583,N_48796,N_49528);
nor UO_584 (O_584,N_46851,N_48456);
or UO_585 (O_585,N_45941,N_46386);
and UO_586 (O_586,N_49100,N_45077);
or UO_587 (O_587,N_49074,N_45842);
nor UO_588 (O_588,N_48212,N_46406);
or UO_589 (O_589,N_47342,N_45219);
and UO_590 (O_590,N_49334,N_46505);
nor UO_591 (O_591,N_46380,N_49347);
xor UO_592 (O_592,N_48345,N_45786);
xor UO_593 (O_593,N_48119,N_45231);
and UO_594 (O_594,N_47743,N_48819);
nand UO_595 (O_595,N_46545,N_47845);
nand UO_596 (O_596,N_48616,N_49138);
nor UO_597 (O_597,N_46352,N_46366);
and UO_598 (O_598,N_49853,N_45990);
and UO_599 (O_599,N_45180,N_46802);
and UO_600 (O_600,N_47718,N_45110);
nand UO_601 (O_601,N_49301,N_45347);
nand UO_602 (O_602,N_46105,N_49893);
or UO_603 (O_603,N_45747,N_49235);
nand UO_604 (O_604,N_49031,N_49431);
or UO_605 (O_605,N_47609,N_49549);
or UO_606 (O_606,N_48463,N_45884);
nand UO_607 (O_607,N_49176,N_49149);
nand UO_608 (O_608,N_45772,N_47181);
nand UO_609 (O_609,N_45829,N_48330);
and UO_610 (O_610,N_46281,N_45191);
nor UO_611 (O_611,N_45860,N_45849);
xor UO_612 (O_612,N_49730,N_47809);
and UO_613 (O_613,N_47933,N_46227);
and UO_614 (O_614,N_49621,N_45230);
nand UO_615 (O_615,N_47792,N_47391);
xor UO_616 (O_616,N_45794,N_49381);
and UO_617 (O_617,N_49442,N_47865);
xnor UO_618 (O_618,N_49545,N_49068);
nand UO_619 (O_619,N_47586,N_47904);
nor UO_620 (O_620,N_46645,N_47201);
nand UO_621 (O_621,N_46980,N_45977);
and UO_622 (O_622,N_47662,N_48444);
and UO_623 (O_623,N_45239,N_49421);
or UO_624 (O_624,N_48873,N_47447);
or UO_625 (O_625,N_45876,N_47163);
or UO_626 (O_626,N_47830,N_46902);
nor UO_627 (O_627,N_47970,N_45548);
nand UO_628 (O_628,N_49778,N_48497);
nor UO_629 (O_629,N_49565,N_47554);
nand UO_630 (O_630,N_47227,N_46502);
nand UO_631 (O_631,N_47467,N_45059);
xnor UO_632 (O_632,N_48812,N_49947);
and UO_633 (O_633,N_46116,N_47431);
nor UO_634 (O_634,N_45537,N_48948);
and UO_635 (O_635,N_49173,N_46788);
nor UO_636 (O_636,N_46088,N_47709);
or UO_637 (O_637,N_47382,N_49685);
nor UO_638 (O_638,N_47767,N_47550);
nor UO_639 (O_639,N_45578,N_49145);
nand UO_640 (O_640,N_48470,N_47476);
or UO_641 (O_641,N_45494,N_49904);
nor UO_642 (O_642,N_49361,N_47153);
nand UO_643 (O_643,N_46102,N_47647);
nand UO_644 (O_644,N_45432,N_45451);
and UO_645 (O_645,N_46979,N_45186);
or UO_646 (O_646,N_48862,N_48476);
nand UO_647 (O_647,N_45527,N_46269);
nor UO_648 (O_648,N_49810,N_46049);
xnor UO_649 (O_649,N_47875,N_45574);
or UO_650 (O_650,N_45182,N_47599);
and UO_651 (O_651,N_48971,N_48747);
or UO_652 (O_652,N_47099,N_48621);
nand UO_653 (O_653,N_45673,N_46159);
nor UO_654 (O_654,N_47720,N_46079);
nand UO_655 (O_655,N_49779,N_47837);
xor UO_656 (O_656,N_45890,N_49543);
nor UO_657 (O_657,N_47480,N_45901);
nand UO_658 (O_658,N_45315,N_49807);
or UO_659 (O_659,N_46395,N_46599);
xor UO_660 (O_660,N_45071,N_48528);
and UO_661 (O_661,N_46641,N_45723);
or UO_662 (O_662,N_46723,N_45552);
nor UO_663 (O_663,N_46279,N_47502);
nor UO_664 (O_664,N_48145,N_49326);
and UO_665 (O_665,N_48606,N_49246);
nand UO_666 (O_666,N_48037,N_45016);
and UO_667 (O_667,N_48833,N_49903);
nand UO_668 (O_668,N_47557,N_45072);
or UO_669 (O_669,N_47974,N_47886);
or UO_670 (O_670,N_46691,N_46590);
or UO_671 (O_671,N_45841,N_49311);
xnor UO_672 (O_672,N_45887,N_49085);
and UO_673 (O_673,N_45264,N_47154);
xor UO_674 (O_674,N_49376,N_49049);
or UO_675 (O_675,N_48335,N_45491);
xor UO_676 (O_676,N_46898,N_47914);
nand UO_677 (O_677,N_46106,N_45699);
nand UO_678 (O_678,N_49838,N_47995);
and UO_679 (O_679,N_47997,N_45626);
nand UO_680 (O_680,N_49092,N_47279);
or UO_681 (O_681,N_49660,N_45691);
nor UO_682 (O_682,N_49956,N_45623);
nor UO_683 (O_683,N_45780,N_49044);
xnor UO_684 (O_684,N_45874,N_49471);
or UO_685 (O_685,N_46021,N_45911);
xor UO_686 (O_686,N_47398,N_45350);
nand UO_687 (O_687,N_48577,N_45324);
nor UO_688 (O_688,N_48482,N_49644);
nand UO_689 (O_689,N_49638,N_49839);
nand UO_690 (O_690,N_48642,N_47090);
and UO_691 (O_691,N_45685,N_47232);
and UO_692 (O_692,N_48192,N_49254);
nand UO_693 (O_693,N_48291,N_47664);
nor UO_694 (O_694,N_45650,N_49002);
and UO_695 (O_695,N_49592,N_46569);
xnor UO_696 (O_696,N_46485,N_45325);
xor UO_697 (O_697,N_46249,N_49180);
or UO_698 (O_698,N_48603,N_47636);
and UO_699 (O_699,N_49576,N_48627);
nand UO_700 (O_700,N_47544,N_45867);
xor UO_701 (O_701,N_49519,N_48791);
nor UO_702 (O_702,N_45081,N_46719);
or UO_703 (O_703,N_49781,N_49184);
and UO_704 (O_704,N_48132,N_47033);
and UO_705 (O_705,N_49854,N_46015);
or UO_706 (O_706,N_48973,N_45753);
nor UO_707 (O_707,N_45008,N_46654);
nand UO_708 (O_708,N_49335,N_48617);
and UO_709 (O_709,N_48489,N_48182);
and UO_710 (O_710,N_45209,N_46458);
nand UO_711 (O_711,N_46219,N_49570);
nand UO_712 (O_712,N_45687,N_49623);
nor UO_713 (O_713,N_49440,N_47653);
and UO_714 (O_714,N_45558,N_47930);
and UO_715 (O_715,N_47778,N_46718);
nor UO_716 (O_716,N_49512,N_49007);
nor UO_717 (O_717,N_46284,N_46676);
nand UO_718 (O_718,N_47063,N_45245);
or UO_719 (O_719,N_49151,N_47424);
and UO_720 (O_720,N_45468,N_47699);
nand UO_721 (O_721,N_49217,N_49923);
xnor UO_722 (O_722,N_48382,N_48068);
xnor UO_723 (O_723,N_49079,N_45061);
nor UO_724 (O_724,N_47871,N_47529);
xnor UO_725 (O_725,N_46615,N_47976);
and UO_726 (O_726,N_48595,N_46204);
xnor UO_727 (O_727,N_47665,N_49841);
or UO_728 (O_728,N_48726,N_48376);
xor UO_729 (O_729,N_48903,N_46196);
and UO_730 (O_730,N_45693,N_46538);
or UO_731 (O_731,N_45256,N_45799);
nor UO_732 (O_732,N_46320,N_46681);
nand UO_733 (O_733,N_46039,N_48021);
and UO_734 (O_734,N_46042,N_48270);
xnor UO_735 (O_735,N_45269,N_47695);
or UO_736 (O_736,N_45310,N_49305);
nor UO_737 (O_737,N_45572,N_47114);
and UO_738 (O_738,N_45668,N_48217);
nand UO_739 (O_739,N_47520,N_45154);
and UO_740 (O_740,N_46808,N_45768);
nor UO_741 (O_741,N_48398,N_47956);
xnor UO_742 (O_742,N_46375,N_48517);
xor UO_743 (O_743,N_46710,N_46679);
xor UO_744 (O_744,N_45403,N_49210);
or UO_745 (O_745,N_49631,N_49196);
nor UO_746 (O_746,N_48858,N_48540);
nand UO_747 (O_747,N_49008,N_49170);
nand UO_748 (O_748,N_47705,N_49082);
nor UO_749 (O_749,N_48757,N_47738);
and UO_750 (O_750,N_48039,N_47925);
nand UO_751 (O_751,N_46696,N_49940);
or UO_752 (O_752,N_48695,N_47907);
nand UO_753 (O_753,N_45627,N_45702);
and UO_754 (O_754,N_49445,N_45404);
and UO_755 (O_755,N_46957,N_47242);
or UO_756 (O_756,N_46411,N_46883);
and UO_757 (O_757,N_46276,N_47736);
and UO_758 (O_758,N_45724,N_46653);
or UO_759 (O_759,N_48247,N_46164);
nand UO_760 (O_760,N_46572,N_48890);
nor UO_761 (O_761,N_46114,N_49664);
xor UO_762 (O_762,N_45822,N_47523);
xor UO_763 (O_763,N_47994,N_47563);
or UO_764 (O_764,N_48783,N_45533);
nand UO_765 (O_765,N_48694,N_47773);
nand UO_766 (O_766,N_46111,N_47671);
nor UO_767 (O_767,N_46834,N_45905);
xnor UO_768 (O_768,N_45048,N_45359);
nand UO_769 (O_769,N_47171,N_48646);
nor UO_770 (O_770,N_47952,N_49995);
and UO_771 (O_771,N_45664,N_46514);
and UO_772 (O_772,N_45441,N_45742);
nor UO_773 (O_773,N_47873,N_48654);
and UO_774 (O_774,N_48222,N_46465);
nor UO_775 (O_775,N_48930,N_49882);
nand UO_776 (O_776,N_46203,N_48773);
nor UO_777 (O_777,N_45864,N_48135);
nor UO_778 (O_778,N_45383,N_45663);
xnor UO_779 (O_779,N_47493,N_49757);
nand UO_780 (O_780,N_46076,N_45025);
nor UO_781 (O_781,N_47730,N_49093);
nor UO_782 (O_782,N_49538,N_49315);
or UO_783 (O_783,N_48549,N_48636);
nor UO_784 (O_784,N_49899,N_45313);
xor UO_785 (O_785,N_46364,N_47012);
nand UO_786 (O_786,N_46305,N_48412);
and UO_787 (O_787,N_48156,N_45399);
nor UO_788 (O_788,N_48785,N_48188);
nand UO_789 (O_789,N_45395,N_45633);
nand UO_790 (O_790,N_46807,N_46618);
nor UO_791 (O_791,N_46224,N_47749);
and UO_792 (O_792,N_48723,N_46908);
or UO_793 (O_793,N_49984,N_46984);
xor UO_794 (O_794,N_45670,N_48625);
or UO_795 (O_795,N_45307,N_45602);
and UO_796 (O_796,N_45436,N_49130);
and UO_797 (O_797,N_45339,N_45550);
or UO_798 (O_798,N_47916,N_46063);
nor UO_799 (O_799,N_47692,N_48711);
xnor UO_800 (O_800,N_47859,N_48571);
nor UO_801 (O_801,N_47251,N_49104);
nor UO_802 (O_802,N_45299,N_47045);
or UO_803 (O_803,N_49266,N_47405);
and UO_804 (O_804,N_47207,N_45079);
xnor UO_805 (O_805,N_48851,N_46524);
xnor UO_806 (O_806,N_49064,N_45287);
or UO_807 (O_807,N_48384,N_49975);
or UO_808 (O_808,N_45539,N_46877);
nand UO_809 (O_809,N_47951,N_46756);
nand UO_810 (O_810,N_48739,N_46503);
nor UO_811 (O_811,N_49641,N_45609);
nand UO_812 (O_812,N_49458,N_47511);
and UO_813 (O_813,N_48282,N_47412);
or UO_814 (O_814,N_48137,N_46356);
or UO_815 (O_815,N_48355,N_49799);
nor UO_816 (O_816,N_49609,N_46925);
nor UO_817 (O_817,N_46747,N_45489);
xnor UO_818 (O_818,N_49846,N_46090);
and UO_819 (O_819,N_45297,N_47568);
nor UO_820 (O_820,N_47906,N_48324);
or UO_821 (O_821,N_46286,N_45027);
nand UO_822 (O_822,N_48895,N_47942);
xor UO_823 (O_823,N_46680,N_47282);
or UO_824 (O_824,N_46729,N_45958);
or UO_825 (O_825,N_45455,N_46867);
and UO_826 (O_826,N_48718,N_45243);
nand UO_827 (O_827,N_47765,N_45734);
or UO_828 (O_828,N_48481,N_47395);
nor UO_829 (O_829,N_48551,N_47656);
nor UO_830 (O_830,N_48795,N_48552);
xnor UO_831 (O_831,N_45891,N_45006);
or UO_832 (O_832,N_46894,N_45199);
xnor UO_833 (O_833,N_46819,N_48824);
nor UO_834 (O_834,N_47786,N_47218);
nand UO_835 (O_835,N_48448,N_49865);
nand UO_836 (O_836,N_46500,N_48025);
xnor UO_837 (O_837,N_47524,N_45541);
nor UO_838 (O_838,N_47861,N_45904);
nand UO_839 (O_839,N_46144,N_48733);
or UO_840 (O_840,N_48689,N_45149);
and UO_841 (O_841,N_46314,N_45773);
nand UO_842 (O_842,N_48272,N_45196);
and UO_843 (O_843,N_48837,N_47459);
nand UO_844 (O_844,N_47484,N_46794);
xor UO_845 (O_845,N_45408,N_45888);
or UO_846 (O_846,N_46226,N_48477);
xor UO_847 (O_847,N_46619,N_49514);
and UO_848 (O_848,N_47623,N_47375);
xnor UO_849 (O_849,N_48242,N_46230);
xor UO_850 (O_850,N_48452,N_46962);
xnor UO_851 (O_851,N_47211,N_47127);
or UO_852 (O_852,N_48852,N_46711);
xnor UO_853 (O_853,N_47363,N_46592);
and UO_854 (O_854,N_48842,N_47611);
nand UO_855 (O_855,N_47055,N_48072);
xnor UO_856 (O_856,N_49389,N_49450);
nand UO_857 (O_857,N_46416,N_46968);
nor UO_858 (O_858,N_48186,N_49221);
nand UO_859 (O_859,N_45808,N_48304);
xor UO_860 (O_860,N_45082,N_45652);
nor UO_861 (O_861,N_45116,N_48807);
and UO_862 (O_862,N_45311,N_47648);
and UO_863 (O_863,N_46156,N_45164);
nand UO_864 (O_864,N_47064,N_45176);
and UO_865 (O_865,N_47752,N_48676);
nor UO_866 (O_866,N_49831,N_46648);
nor UO_867 (O_867,N_47847,N_49225);
xor UO_868 (O_868,N_47285,N_49186);
nand UO_869 (O_869,N_49403,N_46205);
or UO_870 (O_870,N_49795,N_49310);
nor UO_871 (O_871,N_47785,N_47828);
and UO_872 (O_872,N_48163,N_46907);
nor UO_873 (O_873,N_48565,N_49544);
nand UO_874 (O_874,N_46549,N_47220);
nand UO_875 (O_875,N_45254,N_49974);
and UO_876 (O_876,N_47423,N_46228);
and UO_877 (O_877,N_45839,N_46200);
and UO_878 (O_878,N_46430,N_48826);
nor UO_879 (O_879,N_47882,N_47607);
and UO_880 (O_880,N_48223,N_45646);
nor UO_881 (O_881,N_49782,N_48240);
nor UO_882 (O_882,N_45298,N_49332);
nor UO_883 (O_883,N_46367,N_47666);
nand UO_884 (O_884,N_48857,N_45107);
xor UO_885 (O_885,N_45220,N_45211);
xor UO_886 (O_886,N_48839,N_46008);
xor UO_887 (O_887,N_46331,N_45144);
and UO_888 (O_888,N_46002,N_48140);
nand UO_889 (O_889,N_48727,N_47512);
xnor UO_890 (O_890,N_45477,N_49349);
xor UO_891 (O_891,N_46308,N_46012);
or UO_892 (O_892,N_47387,N_47367);
xnor UO_893 (O_893,N_46772,N_45232);
and UO_894 (O_894,N_45515,N_46575);
and UO_895 (O_895,N_49674,N_48697);
and UO_896 (O_896,N_45420,N_47488);
or UO_897 (O_897,N_45426,N_48479);
and UO_898 (O_898,N_49527,N_47826);
and UO_899 (O_899,N_47458,N_46240);
or UO_900 (O_900,N_46960,N_47757);
xnor UO_901 (O_901,N_45018,N_46287);
or UO_902 (O_902,N_48122,N_49819);
xor UO_903 (O_903,N_48393,N_46833);
xnor UO_904 (O_904,N_46583,N_45112);
nand UO_905 (O_905,N_46886,N_45688);
or UO_906 (O_906,N_47108,N_47416);
nor UO_907 (O_907,N_46061,N_49926);
nand UO_908 (O_908,N_49812,N_45422);
nor UO_909 (O_909,N_47228,N_47417);
nor UO_910 (O_910,N_47325,N_47857);
nand UO_911 (O_911,N_47998,N_47896);
xnor UO_912 (O_912,N_45951,N_46929);
xnor UO_913 (O_913,N_47351,N_47261);
xnor UO_914 (O_914,N_49296,N_49036);
nand UO_915 (O_915,N_46977,N_45610);
nand UO_916 (O_916,N_49558,N_45163);
nor UO_917 (O_917,N_46606,N_45365);
and UO_918 (O_918,N_48559,N_47573);
and UO_919 (O_919,N_48782,N_47350);
and UO_920 (O_920,N_47471,N_47953);
nor UO_921 (O_921,N_47418,N_46912);
and UO_922 (O_922,N_46074,N_49019);
and UO_923 (O_923,N_47348,N_46559);
xor UO_924 (O_924,N_46686,N_49591);
xor UO_925 (O_925,N_45334,N_47109);
and UO_926 (O_926,N_48283,N_46614);
nor UO_927 (O_927,N_46491,N_49908);
nand UO_928 (O_928,N_46398,N_47009);
and UO_929 (O_929,N_46289,N_48279);
and UO_930 (O_930,N_47770,N_48087);
nor UO_931 (O_931,N_46125,N_48424);
nor UO_932 (O_932,N_46518,N_45170);
nand UO_933 (O_933,N_49057,N_45815);
or UO_934 (O_934,N_45412,N_48728);
xor UO_935 (O_935,N_48999,N_46620);
xor UO_936 (O_936,N_49906,N_49095);
or UO_937 (O_937,N_46103,N_48378);
or UO_938 (O_938,N_48919,N_48933);
xnor UO_939 (O_939,N_48892,N_48251);
or UO_940 (O_940,N_48069,N_48942);
xnor UO_941 (O_941,N_48758,N_47219);
nor UO_942 (O_942,N_48402,N_47888);
xnor UO_943 (O_943,N_46062,N_47443);
xor UO_944 (O_944,N_46238,N_48427);
nor UO_945 (O_945,N_48522,N_46631);
and UO_946 (O_946,N_48943,N_45474);
or UO_947 (O_947,N_48147,N_49602);
xnor UO_948 (O_948,N_45838,N_46246);
or UO_949 (O_949,N_46554,N_48843);
or UO_950 (O_950,N_47693,N_46241);
and UO_951 (O_951,N_49177,N_48012);
xor UO_952 (O_952,N_45599,N_46080);
and UO_953 (O_953,N_45740,N_47031);
and UO_954 (O_954,N_47080,N_46798);
or UO_955 (O_955,N_46360,N_45488);
or UO_956 (O_956,N_48931,N_49112);
or UO_957 (O_957,N_48874,N_49973);
nor UO_958 (O_958,N_49961,N_45060);
and UO_959 (O_959,N_48651,N_45115);
nand UO_960 (O_960,N_46197,N_46101);
nand UO_961 (O_961,N_46393,N_49509);
xnor UO_962 (O_962,N_48830,N_45568);
nor UO_963 (O_963,N_47206,N_49928);
or UO_964 (O_964,N_46896,N_47344);
xnor UO_965 (O_965,N_46410,N_46792);
and UO_966 (O_966,N_46586,N_49547);
and UO_967 (O_967,N_49960,N_46767);
or UO_968 (O_968,N_49835,N_47880);
or UO_969 (O_969,N_47231,N_48962);
xnor UO_970 (O_970,N_47322,N_49120);
nor UO_971 (O_971,N_46750,N_47628);
nand UO_972 (O_972,N_48447,N_49601);
and UO_973 (O_973,N_48610,N_49531);
and UO_974 (O_974,N_49192,N_47795);
nand UO_975 (O_975,N_45410,N_48764);
xnor UO_976 (O_976,N_49152,N_49481);
and UO_977 (O_977,N_46657,N_49655);
and UO_978 (O_978,N_48232,N_48096);
and UO_979 (O_979,N_47818,N_47157);
nor UO_980 (O_980,N_48219,N_47372);
xnor UO_981 (O_981,N_45666,N_45273);
xor UO_982 (O_982,N_48455,N_49382);
and UO_983 (O_983,N_48512,N_48585);
xor UO_984 (O_984,N_46381,N_47903);
xor UO_985 (O_985,N_48123,N_49108);
xnor UO_986 (O_986,N_45737,N_47131);
and UO_987 (O_987,N_48704,N_45443);
xor UO_988 (O_988,N_45411,N_45518);
and UO_989 (O_989,N_48891,N_49336);
xnor UO_990 (O_990,N_46991,N_48560);
or UO_991 (O_991,N_46517,N_48953);
nor UO_992 (O_992,N_48318,N_47537);
and UO_993 (O_993,N_47025,N_47432);
nand UO_994 (O_994,N_49357,N_47187);
and UO_995 (O_995,N_47781,N_47670);
nand UO_996 (O_996,N_49200,N_47452);
nand UO_997 (O_997,N_46222,N_49507);
or UO_998 (O_998,N_46255,N_46073);
xnor UO_999 (O_999,N_45105,N_45676);
and UO_1000 (O_1000,N_47152,N_46859);
nand UO_1001 (O_1001,N_46325,N_48046);
xor UO_1002 (O_1002,N_47149,N_49520);
and UO_1003 (O_1003,N_49232,N_48400);
xnor UO_1004 (O_1004,N_49294,N_48261);
nor UO_1005 (O_1005,N_47058,N_48308);
nor UO_1006 (O_1006,N_45333,N_48888);
or UO_1007 (O_1007,N_48388,N_48401);
or UO_1008 (O_1008,N_47858,N_48838);
and UO_1009 (O_1009,N_48583,N_45525);
or UO_1010 (O_1010,N_48856,N_49883);
or UO_1011 (O_1011,N_47291,N_46928);
nor UO_1012 (O_1012,N_45821,N_48130);
xnor UO_1013 (O_1013,N_47027,N_46934);
xor UO_1014 (O_1014,N_46041,N_48100);
and UO_1015 (O_1015,N_46011,N_48995);
and UO_1016 (O_1016,N_45125,N_45285);
or UO_1017 (O_1017,N_46712,N_48109);
and UO_1018 (O_1018,N_45557,N_48349);
nand UO_1019 (O_1019,N_45262,N_45198);
nand UO_1020 (O_1020,N_47651,N_47620);
nand UO_1021 (O_1021,N_47707,N_46490);
and UO_1022 (O_1022,N_48357,N_46519);
xnor UO_1023 (O_1023,N_47715,N_48390);
nand UO_1024 (O_1024,N_48468,N_49646);
or UO_1025 (O_1025,N_46329,N_46207);
nor UO_1026 (O_1026,N_46402,N_48319);
nor UO_1027 (O_1027,N_45312,N_48498);
xor UO_1028 (O_1028,N_49394,N_48076);
xnor UO_1029 (O_1029,N_45918,N_48992);
xnor UO_1030 (O_1030,N_48224,N_48707);
nor UO_1031 (O_1031,N_49388,N_46593);
nand UO_1032 (O_1032,N_47851,N_48009);
or UO_1033 (O_1033,N_49219,N_49523);
and UO_1034 (O_1034,N_47542,N_49265);
nor UO_1035 (O_1035,N_48118,N_49994);
nor UO_1036 (O_1036,N_47533,N_46950);
nor UO_1037 (O_1037,N_46945,N_48772);
and UO_1038 (O_1038,N_49286,N_49183);
nor UO_1039 (O_1039,N_47336,N_49530);
nand UO_1040 (O_1040,N_48658,N_45681);
nand UO_1041 (O_1041,N_46457,N_49611);
and UO_1042 (O_1042,N_49574,N_45942);
nand UO_1043 (O_1043,N_49935,N_45316);
nor UO_1044 (O_1044,N_46489,N_45022);
nor UO_1045 (O_1045,N_48195,N_47934);
nor UO_1046 (O_1046,N_46178,N_46071);
and UO_1047 (O_1047,N_48914,N_47360);
nand UO_1048 (O_1048,N_49557,N_45797);
nor UO_1049 (O_1049,N_49014,N_45031);
nand UO_1050 (O_1050,N_47788,N_47902);
nor UO_1051 (O_1051,N_49885,N_48670);
nand UO_1052 (O_1052,N_46975,N_47113);
or UO_1053 (O_1053,N_47199,N_48877);
and UO_1054 (O_1054,N_46400,N_45346);
and UO_1055 (O_1055,N_46899,N_46621);
xor UO_1056 (O_1056,N_46378,N_45754);
xnor UO_1057 (O_1057,N_46497,N_49395);
and UO_1058 (O_1058,N_49759,N_49215);
and UO_1059 (O_1059,N_45661,N_45944);
nand UO_1060 (O_1060,N_48848,N_49263);
and UO_1061 (O_1061,N_45710,N_45322);
nand UO_1062 (O_1062,N_47538,N_45971);
nand UO_1063 (O_1063,N_47525,N_45131);
or UO_1064 (O_1064,N_49422,N_47766);
and UO_1065 (O_1065,N_46234,N_47608);
nor UO_1066 (O_1066,N_48693,N_45013);
or UO_1067 (O_1067,N_46904,N_48305);
nand UO_1068 (O_1068,N_49508,N_46384);
and UO_1069 (O_1069,N_48755,N_48828);
and UO_1070 (O_1070,N_45570,N_47088);
and UO_1071 (O_1071,N_46700,N_45781);
or UO_1072 (O_1072,N_47566,N_49016);
xnor UO_1073 (O_1073,N_47734,N_46014);
nor UO_1074 (O_1074,N_46893,N_47605);
xnor UO_1075 (O_1075,N_46130,N_46849);
nor UO_1076 (O_1076,N_47824,N_48703);
xnor UO_1077 (O_1077,N_49418,N_47485);
and UO_1078 (O_1078,N_48691,N_49653);
nor UO_1079 (O_1079,N_46237,N_48997);
or UO_1080 (O_1080,N_45920,N_46939);
nand UO_1081 (O_1081,N_48264,N_45354);
and UO_1082 (O_1082,N_45953,N_48246);
xnor UO_1083 (O_1083,N_46560,N_45153);
xnor UO_1084 (O_1084,N_45039,N_46358);
nand UO_1085 (O_1085,N_45614,N_48488);
nand UO_1086 (O_1086,N_49256,N_47682);
and UO_1087 (O_1087,N_46312,N_49461);
nand UO_1088 (O_1088,N_46601,N_48263);
nand UO_1089 (O_1089,N_45233,N_48771);
nand UO_1090 (O_1090,N_46761,N_45825);
and UO_1091 (O_1091,N_45464,N_47300);
and UO_1092 (O_1092,N_47526,N_48789);
or UO_1093 (O_1093,N_46420,N_49741);
xor UO_1094 (O_1094,N_49417,N_45556);
nand UO_1095 (O_1095,N_48125,N_48091);
nand UO_1096 (O_1096,N_49377,N_48923);
nor UO_1097 (O_1097,N_45290,N_49568);
or UO_1098 (O_1098,N_48245,N_45524);
nor UO_1099 (O_1099,N_49774,N_47072);
or UO_1100 (O_1100,N_45351,N_46171);
nor UO_1101 (O_1101,N_47540,N_45721);
and UO_1102 (O_1102,N_47594,N_49268);
and UO_1103 (O_1103,N_48527,N_48861);
nor UO_1104 (O_1104,N_48905,N_49168);
nor UO_1105 (O_1105,N_45819,N_48206);
xor UO_1106 (O_1106,N_48259,N_47365);
xor UO_1107 (O_1107,N_45417,N_47603);
xnor UO_1108 (O_1108,N_47972,N_47329);
and UO_1109 (O_1109,N_45341,N_49069);
nor UO_1110 (O_1110,N_49273,N_45701);
or UO_1111 (O_1111,N_45793,N_48426);
nor UO_1112 (O_1112,N_48784,N_45097);
nand UO_1113 (O_1113,N_46443,N_47834);
nand UO_1114 (O_1114,N_46650,N_47070);
or UO_1115 (O_1115,N_47962,N_45141);
nor UO_1116 (O_1116,N_48243,N_45189);
xnor UO_1117 (O_1117,N_45853,N_47879);
nand UO_1118 (O_1118,N_47092,N_45813);
and UO_1119 (O_1119,N_49328,N_49933);
nand UO_1120 (O_1120,N_48991,N_49434);
or UO_1121 (O_1121,N_46850,N_45225);
and UO_1122 (O_1122,N_48253,N_46831);
nand UO_1123 (O_1123,N_48983,N_46120);
or UO_1124 (O_1124,N_45877,N_49516);
xor UO_1125 (O_1125,N_46801,N_47105);
or UO_1126 (O_1126,N_46530,N_45986);
nor UO_1127 (O_1127,N_45258,N_49227);
or UO_1128 (O_1128,N_48051,N_45049);
nand UO_1129 (O_1129,N_47710,N_49915);
or UO_1130 (O_1130,N_45579,N_46283);
and UO_1131 (O_1131,N_47370,N_47427);
nor UO_1132 (O_1132,N_45160,N_47660);
and UO_1133 (O_1133,N_48675,N_47915);
and UO_1134 (O_1134,N_49278,N_46214);
and UO_1135 (O_1135,N_49952,N_45343);
nand UO_1136 (O_1136,N_48399,N_46739);
and UO_1137 (O_1137,N_46046,N_48511);
nand UO_1138 (O_1138,N_49704,N_46742);
xor UO_1139 (O_1139,N_47532,N_48673);
or UO_1140 (O_1140,N_48207,N_47340);
and UO_1141 (O_1141,N_45962,N_48485);
xor UO_1142 (O_1142,N_46478,N_45036);
nand UO_1143 (O_1143,N_48467,N_45087);
nand UO_1144 (O_1144,N_48502,N_45669);
xor UO_1145 (O_1145,N_46467,N_45895);
and UO_1146 (O_1146,N_49657,N_45304);
and UO_1147 (O_1147,N_45024,N_46573);
or UO_1148 (O_1148,N_48972,N_47604);
nand UO_1149 (O_1149,N_48367,N_46306);
or UO_1150 (O_1150,N_45362,N_49048);
nand UO_1151 (O_1151,N_49861,N_46033);
and UO_1152 (O_1152,N_48438,N_46677);
xor UO_1153 (O_1153,N_45469,N_46863);
nand UO_1154 (O_1154,N_45438,N_45816);
and UO_1155 (O_1155,N_49033,N_49040);
and UO_1156 (O_1156,N_48297,N_48238);
and UO_1157 (O_1157,N_46577,N_45064);
or UO_1158 (O_1158,N_48986,N_47203);
nor UO_1159 (O_1159,N_48007,N_49279);
nand UO_1160 (O_1160,N_45484,N_47661);
xnor UO_1161 (O_1161,N_46638,N_48315);
and UO_1162 (O_1162,N_46321,N_46169);
xor UO_1163 (O_1163,N_45739,N_47273);
nor UO_1164 (O_1164,N_45425,N_46162);
xnor UO_1165 (O_1165,N_47472,N_46698);
nand UO_1166 (O_1166,N_46995,N_49362);
and UO_1167 (O_1167,N_47172,N_47833);
nand UO_1168 (O_1168,N_49102,N_45593);
nand UO_1169 (O_1169,N_46826,N_49220);
nor UO_1170 (O_1170,N_45989,N_49419);
and UO_1171 (O_1171,N_48103,N_45207);
nor UO_1172 (O_1172,N_49713,N_49276);
nand UO_1173 (O_1173,N_49340,N_46417);
nand UO_1174 (O_1174,N_48002,N_46582);
xor UO_1175 (O_1175,N_49028,N_47668);
and UO_1176 (O_1176,N_49067,N_46721);
or UO_1177 (O_1177,N_45637,N_47696);
xor UO_1178 (O_1178,N_47390,N_48486);
nor UO_1179 (O_1179,N_45434,N_47402);
xnor UO_1180 (O_1180,N_48912,N_46521);
nor UO_1181 (O_1181,N_45466,N_45150);
nand UO_1182 (O_1182,N_47062,N_45733);
nor UO_1183 (O_1183,N_48906,N_45640);
and UO_1184 (O_1184,N_48576,N_47222);
nor UO_1185 (O_1185,N_49406,N_49065);
nor UO_1186 (O_1186,N_46526,N_47927);
nor UO_1187 (O_1187,N_46365,N_48717);
nor UO_1188 (O_1188,N_46822,N_46624);
nand UO_1189 (O_1189,N_46717,N_49738);
and UO_1190 (O_1190,N_47750,N_46966);
nor UO_1191 (O_1191,N_49905,N_47420);
and UO_1192 (O_1192,N_45398,N_46409);
xnor UO_1193 (O_1193,N_46596,N_49745);
xor UO_1194 (O_1194,N_49575,N_49959);
nand UO_1195 (O_1195,N_49577,N_45331);
nor UO_1196 (O_1196,N_46254,N_45875);
nor UO_1197 (O_1197,N_47698,N_47208);
xnor UO_1198 (O_1198,N_46671,N_45995);
or UO_1199 (O_1199,N_49699,N_47073);
nor UO_1200 (O_1200,N_45431,N_47789);
xnor UO_1201 (O_1201,N_49702,N_46349);
nor UO_1202 (O_1202,N_48634,N_48083);
xnor UO_1203 (O_1203,N_45109,N_46964);
and UO_1204 (O_1204,N_47076,N_47286);
and UO_1205 (O_1205,N_49594,N_47754);
nor UO_1206 (O_1206,N_47517,N_45741);
nand UO_1207 (O_1207,N_47755,N_45758);
nor UO_1208 (O_1208,N_46978,N_46827);
and UO_1209 (O_1209,N_49697,N_45278);
xnor UO_1210 (O_1210,N_45647,N_46119);
nand UO_1211 (O_1211,N_45103,N_46532);
or UO_1212 (O_1212,N_48492,N_45215);
nor UO_1213 (O_1213,N_48709,N_45005);
and UO_1214 (O_1214,N_48124,N_46817);
xor UO_1215 (O_1215,N_49284,N_46371);
nor UO_1216 (O_1216,N_48097,N_48725);
and UO_1217 (O_1217,N_45126,N_46591);
nand UO_1218 (O_1218,N_45281,N_47277);
nor UO_1219 (O_1219,N_46247,N_45917);
and UO_1220 (O_1220,N_46131,N_46715);
xnor UO_1221 (O_1221,N_47451,N_49487);
or UO_1222 (O_1222,N_46067,N_45387);
xnor UO_1223 (O_1223,N_49290,N_49909);
or UO_1224 (O_1224,N_48653,N_47320);
and UO_1225 (O_1225,N_47170,N_46413);
and UO_1226 (O_1226,N_48370,N_46699);
xnor UO_1227 (O_1227,N_49165,N_48093);
nor UO_1228 (O_1228,N_47667,N_49368);
and UO_1229 (O_1229,N_49299,N_48106);
xnor UO_1230 (O_1230,N_46147,N_48295);
xor UO_1231 (O_1231,N_45641,N_48955);
nor UO_1232 (O_1232,N_45697,N_45308);
xnor UO_1233 (O_1233,N_48055,N_45992);
nor UO_1234 (O_1234,N_48432,N_49236);
nand UO_1235 (O_1235,N_46354,N_48937);
or UO_1236 (O_1236,N_49736,N_49101);
xnor UO_1237 (O_1237,N_49554,N_48520);
nor UO_1238 (O_1238,N_46567,N_45100);
or UO_1239 (O_1239,N_45991,N_48204);
nor UO_1240 (O_1240,N_45980,N_46933);
xor UO_1241 (O_1241,N_46751,N_48166);
nor UO_1242 (O_1242,N_48019,N_49094);
nand UO_1243 (O_1243,N_49687,N_46303);
nand UO_1244 (O_1244,N_47961,N_45513);
or UO_1245 (O_1245,N_46643,N_48038);
nand UO_1246 (O_1246,N_45270,N_45337);
nor UO_1247 (O_1247,N_45377,N_48161);
xor UO_1248 (O_1248,N_46091,N_45826);
and UO_1249 (O_1249,N_45288,N_48525);
or UO_1250 (O_1250,N_45827,N_47065);
xor UO_1251 (O_1251,N_46265,N_47622);
xnor UO_1252 (O_1252,N_47003,N_49679);
nand UO_1253 (O_1253,N_46193,N_46032);
or UO_1254 (O_1254,N_45439,N_47630);
nor UO_1255 (O_1255,N_48863,N_48129);
or UO_1256 (O_1256,N_46257,N_46875);
xnor UO_1257 (O_1257,N_48310,N_46126);
xor UO_1258 (O_1258,N_45575,N_49818);
xnor UO_1259 (O_1259,N_49010,N_49828);
and UO_1260 (O_1260,N_45179,N_48414);
and UO_1261 (O_1261,N_46235,N_45644);
and UO_1262 (O_1262,N_46185,N_49494);
nand UO_1263 (O_1263,N_47388,N_48073);
nor UO_1264 (O_1264,N_46558,N_49635);
nand UO_1265 (O_1265,N_45012,N_45471);
or UO_1266 (O_1266,N_47428,N_47225);
nor UO_1267 (O_1267,N_45581,N_48629);
or UO_1268 (O_1268,N_47381,N_49731);
and UO_1269 (O_1269,N_45089,N_49190);
nand UO_1270 (O_1270,N_48746,N_48907);
and UO_1271 (O_1271,N_46705,N_46288);
and UO_1272 (O_1272,N_46077,N_47331);
nand UO_1273 (O_1273,N_47853,N_46755);
and UO_1274 (O_1274,N_49700,N_46673);
nor UO_1275 (O_1275,N_47968,N_48710);
nand UO_1276 (O_1276,N_48328,N_46574);
xnor UO_1277 (O_1277,N_47724,N_48230);
and UO_1278 (O_1278,N_46811,N_46992);
and UO_1279 (O_1279,N_48635,N_46309);
nand UO_1280 (O_1280,N_46612,N_45563);
or UO_1281 (O_1281,N_45756,N_46871);
nand UO_1282 (O_1282,N_49673,N_45453);
nand UO_1283 (O_1283,N_45472,N_49241);
and UO_1284 (O_1284,N_46890,N_46372);
and UO_1285 (O_1285,N_45492,N_47783);
xnor UO_1286 (O_1286,N_45709,N_49617);
and UO_1287 (O_1287,N_47595,N_48341);
or UO_1288 (O_1288,N_45117,N_49378);
nand UO_1289 (O_1289,N_49964,N_46236);
nor UO_1290 (O_1290,N_48506,N_46997);
nand UO_1291 (O_1291,N_46547,N_46674);
or UO_1292 (O_1292,N_47441,N_49571);
and UO_1293 (O_1293,N_47429,N_49681);
or UO_1294 (O_1294,N_46610,N_49366);
xor UO_1295 (O_1295,N_48864,N_45169);
nor UO_1296 (O_1296,N_47978,N_47519);
nor UO_1297 (O_1297,N_46930,N_45510);
and UO_1298 (O_1298,N_49191,N_47977);
or UO_1299 (O_1299,N_49396,N_45445);
or UO_1300 (O_1300,N_46774,N_49207);
nand UO_1301 (O_1301,N_48030,N_49029);
or UO_1302 (O_1302,N_49077,N_46688);
and UO_1303 (O_1303,N_49823,N_45912);
xor UO_1304 (O_1304,N_48732,N_46127);
nand UO_1305 (O_1305,N_47465,N_48882);
xor UO_1306 (O_1306,N_45873,N_46860);
nor UO_1307 (O_1307,N_49495,N_48567);
or UO_1308 (O_1308,N_47504,N_49533);
nand UO_1309 (O_1309,N_45481,N_47217);
or UO_1310 (O_1310,N_48006,N_47385);
nor UO_1311 (O_1311,N_49037,N_47808);
nor UO_1312 (O_1312,N_49886,N_46941);
xor UO_1313 (O_1313,N_46810,N_46456);
nor UO_1314 (O_1314,N_47096,N_47150);
xor UO_1315 (O_1315,N_47964,N_45250);
nor UO_1316 (O_1316,N_49867,N_48369);
and UO_1317 (O_1317,N_47048,N_48724);
xnor UO_1318 (O_1318,N_46025,N_49642);
nand UO_1319 (O_1319,N_46198,N_48013);
xnor UO_1320 (O_1320,N_45435,N_45017);
and UO_1321 (O_1321,N_46689,N_47922);
or UO_1322 (O_1322,N_47249,N_49111);
or UO_1323 (O_1323,N_49842,N_46486);
xnor UO_1324 (O_1324,N_47013,N_46790);
xnor UO_1325 (O_1325,N_45370,N_47555);
nor UO_1326 (O_1326,N_49247,N_45091);
xnor UO_1327 (O_1327,N_49669,N_49066);
nor UO_1328 (O_1328,N_49135,N_45940);
nand UO_1329 (O_1329,N_48500,N_49000);
nor UO_1330 (O_1330,N_45749,N_48600);
xnor UO_1331 (O_1331,N_48659,N_46280);
or UO_1332 (O_1332,N_45965,N_49525);
and UO_1333 (O_1333,N_48431,N_49118);
and UO_1334 (O_1334,N_47616,N_48897);
and UO_1335 (O_1335,N_47841,N_48548);
or UO_1336 (O_1336,N_45328,N_49980);
nor UO_1337 (O_1337,N_49825,N_45844);
and UO_1338 (O_1338,N_47257,N_45779);
nor UO_1339 (O_1339,N_49293,N_49231);
nand UO_1340 (O_1340,N_48080,N_46821);
nor UO_1341 (O_1341,N_45931,N_46451);
nand UO_1342 (O_1342,N_47345,N_49443);
xor UO_1343 (O_1343,N_48208,N_45415);
xnor UO_1344 (O_1344,N_47876,N_47740);
xor UO_1345 (O_1345,N_47892,N_48602);
nand UO_1346 (O_1346,N_48946,N_49325);
nor UO_1347 (O_1347,N_46924,N_46693);
and UO_1348 (O_1348,N_45380,N_47747);
and UO_1349 (O_1349,N_46759,N_48832);
nand UO_1350 (O_1350,N_48234,N_45177);
xnor UO_1351 (O_1351,N_48976,N_48831);
nand UO_1352 (O_1352,N_45000,N_47121);
xnor UO_1353 (O_1353,N_48049,N_47597);
and UO_1354 (O_1354,N_47021,N_49400);
or UO_1355 (O_1355,N_47732,N_48365);
nand UO_1356 (O_1356,N_46343,N_48562);
or UO_1357 (O_1357,N_49920,N_45889);
and UO_1358 (O_1358,N_49466,N_45767);
nand UO_1359 (O_1359,N_46100,N_46919);
nand UO_1360 (O_1360,N_47574,N_49171);
or UO_1361 (O_1361,N_49321,N_45358);
nand UO_1362 (O_1362,N_45261,N_48041);
nand UO_1363 (O_1363,N_49160,N_49199);
or UO_1364 (O_1364,N_49537,N_45832);
xor UO_1365 (O_1365,N_47640,N_45588);
nand UO_1366 (O_1366,N_49791,N_46746);
nor UO_1367 (O_1367,N_45128,N_45801);
and UO_1368 (O_1368,N_47989,N_45032);
nor UO_1369 (O_1369,N_45618,N_47959);
nor UO_1370 (O_1370,N_49155,N_46016);
xor UO_1371 (O_1371,N_48881,N_47030);
or UO_1372 (O_1372,N_49224,N_48531);
nor UO_1373 (O_1373,N_47319,N_45010);
nand UO_1374 (O_1374,N_47505,N_47719);
nand UO_1375 (O_1375,N_46267,N_46064);
nor UO_1376 (O_1376,N_45247,N_45847);
xnor UO_1377 (O_1377,N_45146,N_45711);
xor UO_1378 (O_1378,N_48178,N_46324);
xor UO_1379 (O_1379,N_49306,N_48088);
nor UO_1380 (O_1380,N_46268,N_48541);
nor UO_1381 (O_1381,N_45776,N_48744);
nor UO_1382 (O_1382,N_47672,N_47884);
nand UO_1383 (O_1383,N_47147,N_49727);
nor UO_1384 (O_1384,N_45321,N_49868);
nand UO_1385 (O_1385,N_48979,N_47931);
nand UO_1386 (O_1386,N_45698,N_46390);
or UO_1387 (O_1387,N_49133,N_48802);
and UO_1388 (O_1388,N_45573,N_46639);
and UO_1389 (O_1389,N_46915,N_48760);
or UO_1390 (O_1390,N_46270,N_48105);
nand UO_1391 (O_1391,N_46722,N_48586);
nand UO_1392 (O_1392,N_49363,N_47040);
nand UO_1393 (O_1393,N_47368,N_48403);
or UO_1394 (O_1394,N_47798,N_45452);
nand UO_1395 (O_1395,N_48641,N_48128);
nor UO_1396 (O_1396,N_48214,N_47780);
or UO_1397 (O_1397,N_47731,N_47714);
nor UO_1398 (O_1398,N_49139,N_46431);
nor UO_1399 (O_1399,N_49858,N_47980);
nand UO_1400 (O_1400,N_47784,N_45907);
xor UO_1401 (O_1401,N_47386,N_48340);
or UO_1402 (O_1402,N_46835,N_46905);
and UO_1403 (O_1403,N_46473,N_47326);
or UO_1404 (O_1404,N_49553,N_47313);
or UO_1405 (O_1405,N_47287,N_49479);
nor UO_1406 (O_1406,N_49015,N_47303);
or UO_1407 (O_1407,N_45044,N_47378);
nand UO_1408 (O_1408,N_46392,N_48048);
nor UO_1409 (O_1409,N_48203,N_49021);
and UO_1410 (O_1410,N_48575,N_46748);
and UO_1411 (O_1411,N_47674,N_49840);
xor UO_1412 (O_1412,N_48786,N_45643);
and UO_1413 (O_1413,N_45214,N_47439);
nand UO_1414 (O_1414,N_49142,N_47494);
nor UO_1415 (O_1415,N_48062,N_49816);
nand UO_1416 (O_1416,N_46174,N_46531);
and UO_1417 (O_1417,N_45631,N_49083);
nor UO_1418 (O_1418,N_49796,N_46123);
nor UO_1419 (O_1419,N_47341,N_45406);
xor UO_1420 (O_1420,N_48618,N_46357);
or UO_1421 (O_1421,N_48687,N_47468);
or UO_1422 (O_1422,N_46793,N_48235);
nand UO_1423 (O_1423,N_47258,N_48605);
or UO_1424 (O_1424,N_46651,N_47044);
xnor UO_1425 (O_1425,N_48058,N_47885);
and UO_1426 (O_1426,N_46508,N_49282);
and UO_1427 (O_1427,N_47189,N_49277);
nor UO_1428 (O_1428,N_49769,N_48164);
xor UO_1429 (O_1429,N_47697,N_46852);
nor UO_1430 (O_1430,N_46506,N_45168);
xnor UO_1431 (O_1431,N_49181,N_45879);
or UO_1432 (O_1432,N_45226,N_46154);
xor UO_1433 (O_1433,N_45152,N_49712);
nand UO_1434 (O_1434,N_47629,N_48435);
and UO_1435 (O_1435,N_45672,N_45778);
nor UO_1436 (O_1436,N_47137,N_46692);
nor UO_1437 (O_1437,N_45638,N_45396);
nor UO_1438 (O_1438,N_49511,N_48346);
nor UO_1439 (O_1439,N_45113,N_46996);
and UO_1440 (O_1440,N_47657,N_49143);
nor UO_1441 (O_1441,N_48017,N_49729);
and UO_1442 (O_1442,N_49844,N_47839);
xor UO_1443 (O_1443,N_47399,N_45613);
nor UO_1444 (O_1444,N_45301,N_46459);
nand UO_1445 (O_1445,N_47444,N_47308);
nor UO_1446 (O_1446,N_49374,N_48406);
xor UO_1447 (O_1447,N_48503,N_48268);
xnor UO_1448 (O_1448,N_46399,N_47146);
or UO_1449 (O_1449,N_48461,N_48117);
xnor UO_1450 (O_1450,N_49052,N_49634);
nand UO_1451 (O_1451,N_45921,N_49944);
xor UO_1452 (O_1452,N_46656,N_45002);
and UO_1453 (O_1453,N_46142,N_48316);
or UO_1454 (O_1454,N_49038,N_48681);
xnor UO_1455 (O_1455,N_46326,N_47167);
or UO_1456 (O_1456,N_45366,N_47835);
nand UO_1457 (O_1457,N_45878,N_47843);
xor UO_1458 (O_1458,N_47186,N_48413);
nand UO_1459 (O_1459,N_46838,N_45969);
and UO_1460 (O_1460,N_45478,N_48303);
and UO_1461 (O_1461,N_49253,N_45540);
nand UO_1462 (O_1462,N_48045,N_45660);
or UO_1463 (O_1463,N_46422,N_46124);
and UO_1464 (O_1464,N_47082,N_48348);
nor UO_1465 (O_1465,N_46332,N_47056);
xor UO_1466 (O_1466,N_49024,N_48008);
xor UO_1467 (O_1467,N_47470,N_48800);
and UO_1468 (O_1468,N_49608,N_46057);
and UO_1469 (O_1469,N_49239,N_45038);
nand UO_1470 (O_1470,N_45342,N_48649);
and UO_1471 (O_1471,N_45124,N_48661);
xor UO_1472 (O_1472,N_48250,N_47144);
nand UO_1473 (O_1473,N_49567,N_49323);
nand UO_1474 (O_1474,N_48539,N_46552);
nand UO_1475 (O_1475,N_49777,N_48337);
and UO_1476 (O_1476,N_49522,N_49267);
and UO_1477 (O_1477,N_46191,N_45080);
xor UO_1478 (O_1478,N_48351,N_48173);
or UO_1479 (O_1479,N_48287,N_45930);
xnor UO_1480 (O_1480,N_47658,N_46232);
xnor UO_1481 (O_1481,N_49474,N_48418);
or UO_1482 (O_1482,N_46998,N_49214);
nor UO_1483 (O_1483,N_49312,N_45306);
nor UO_1484 (O_1484,N_47177,N_45655);
nor UO_1485 (O_1485,N_47483,N_46507);
or UO_1486 (O_1486,N_45166,N_49948);
xor UO_1487 (O_1487,N_48753,N_45413);
nor UO_1488 (O_1488,N_49929,N_45900);
or UO_1489 (O_1489,N_49034,N_48453);
nor UO_1490 (O_1490,N_47414,N_49517);
xor UO_1491 (O_1491,N_49429,N_47116);
nand UO_1492 (O_1492,N_46536,N_47899);
or UO_1493 (O_1493,N_46843,N_46735);
or UO_1494 (O_1494,N_45532,N_48611);
xor UO_1495 (O_1495,N_45357,N_46136);
nand UO_1496 (O_1496,N_47949,N_46942);
nand UO_1497 (O_1497,N_49856,N_45979);
xor UO_1498 (O_1498,N_47192,N_48741);
xnor UO_1499 (O_1499,N_49937,N_48162);
nor UO_1500 (O_1500,N_47098,N_48136);
or UO_1501 (O_1501,N_47979,N_45272);
and UO_1502 (O_1502,N_49776,N_46208);
or UO_1503 (O_1503,N_45649,N_47260);
and UO_1504 (O_1504,N_45011,N_48536);
xor UO_1505 (O_1505,N_49896,N_45935);
xor UO_1506 (O_1506,N_49211,N_49030);
xnor UO_1507 (O_1507,N_46186,N_46578);
and UO_1508 (O_1508,N_47543,N_45885);
nor UO_1509 (O_1509,N_48780,N_47312);
nand UO_1510 (O_1510,N_46340,N_48499);
nand UO_1511 (O_1511,N_47547,N_47426);
or UO_1512 (O_1512,N_47621,N_46054);
nand UO_1513 (O_1513,N_46988,N_47849);
nand UO_1514 (O_1514,N_46035,N_49672);
nand UO_1515 (O_1515,N_48343,N_45235);
and UO_1516 (O_1516,N_48160,N_49163);
or UO_1517 (O_1517,N_49979,N_47198);
nand UO_1518 (O_1518,N_47477,N_47450);
xnor UO_1519 (O_1519,N_49968,N_47881);
nor UO_1520 (O_1520,N_46667,N_46858);
and UO_1521 (O_1521,N_47817,N_47545);
or UO_1522 (O_1522,N_46987,N_49992);
or UO_1523 (O_1523,N_49202,N_48572);
xor UO_1524 (O_1524,N_47832,N_48362);
xor UO_1525 (O_1525,N_48487,N_45784);
or UO_1526 (O_1526,N_45943,N_48149);
and UO_1527 (O_1527,N_45718,N_46778);
nor UO_1528 (O_1528,N_48372,N_49448);
nor UO_1529 (O_1529,N_48032,N_45694);
xnor UO_1530 (O_1530,N_49369,N_45555);
xnor UO_1531 (O_1531,N_46093,N_48965);
xor UO_1532 (O_1532,N_49957,N_48834);
and UO_1533 (O_1533,N_47596,N_46434);
nor UO_1534 (O_1534,N_49463,N_47297);
nand UO_1535 (O_1535,N_46291,N_49063);
nor UO_1536 (O_1536,N_49348,N_47943);
nor UO_1537 (O_1537,N_48170,N_45374);
xnor UO_1538 (O_1538,N_46405,N_48034);
xor UO_1539 (O_1539,N_45651,N_49750);
and UO_1540 (O_1540,N_49342,N_49283);
or UO_1541 (O_1541,N_45771,N_46470);
nor UO_1542 (O_1542,N_46587,N_46713);
nand UO_1543 (O_1543,N_49972,N_49017);
nor UO_1544 (O_1544,N_49711,N_49053);
nor UO_1545 (O_1545,N_48949,N_45789);
or UO_1546 (O_1546,N_49792,N_48929);
nand UO_1547 (O_1547,N_45763,N_46081);
and UO_1548 (O_1548,N_49497,N_45818);
and UO_1549 (O_1549,N_47811,N_45437);
or UO_1550 (O_1550,N_46292,N_49728);
and UO_1551 (O_1551,N_46927,N_49411);
and UO_1552 (O_1552,N_49794,N_45066);
nor UO_1553 (O_1553,N_46166,N_48108);
nand UO_1554 (O_1554,N_47562,N_49162);
nor UO_1555 (O_1555,N_45248,N_46112);
nand UO_1556 (O_1556,N_48190,N_47689);
and UO_1557 (O_1557,N_46986,N_46346);
xor UO_1558 (O_1558,N_45356,N_47196);
or UO_1559 (O_1559,N_46469,N_48756);
nand UO_1560 (O_1560,N_45857,N_49907);
nor UO_1561 (O_1561,N_48835,N_48596);
xor UO_1562 (O_1562,N_47820,N_47057);
xnor UO_1563 (O_1563,N_49206,N_47210);
nor UO_1564 (O_1564,N_45482,N_47183);
and UO_1565 (O_1565,N_47050,N_48134);
nand UO_1566 (O_1566,N_47404,N_49189);
and UO_1567 (O_1567,N_48715,N_49651);
and UO_1568 (O_1568,N_49076,N_48241);
nand UO_1569 (O_1569,N_46704,N_46482);
and UO_1570 (O_1570,N_46658,N_48302);
nand UO_1571 (O_1571,N_48581,N_45074);
nor UO_1572 (O_1572,N_45034,N_46437);
nand UO_1573 (O_1573,N_45654,N_49658);
and UO_1574 (O_1574,N_48018,N_47735);
nor UO_1575 (O_1575,N_46522,N_48003);
xnor UO_1576 (O_1576,N_49988,N_49280);
nor UO_1577 (O_1577,N_49582,N_46800);
and UO_1578 (O_1578,N_45275,N_47999);
xor UO_1579 (O_1579,N_46275,N_46261);
xor UO_1580 (O_1580,N_47054,N_49647);
and UO_1581 (O_1581,N_45127,N_46066);
nor UO_1582 (O_1582,N_49300,N_49762);
nor UO_1583 (O_1583,N_45364,N_48766);
nand UO_1584 (O_1584,N_45855,N_48947);
or UO_1585 (O_1585,N_45386,N_47782);
and UO_1586 (O_1586,N_47259,N_46564);
nand UO_1587 (O_1587,N_47948,N_49829);
xnor UO_1588 (O_1588,N_49146,N_48678);
xor UO_1589 (O_1589,N_48433,N_47244);
nor UO_1590 (O_1590,N_45692,N_46990);
nand UO_1591 (O_1591,N_45371,N_46089);
nand UO_1592 (O_1592,N_48044,N_46965);
nand UO_1593 (O_1593,N_49041,N_49359);
or UO_1594 (O_1594,N_48441,N_49989);
and UO_1595 (O_1595,N_48112,N_45148);
nor UO_1596 (O_1596,N_45118,N_49855);
xnor UO_1597 (O_1597,N_46973,N_47764);
nor UO_1598 (O_1598,N_46520,N_45073);
xnor UO_1599 (O_1599,N_46636,N_46879);
nand UO_1600 (O_1600,N_45505,N_49468);
nor UO_1601 (O_1601,N_47626,N_48885);
and UO_1602 (O_1602,N_48980,N_47854);
nor UO_1603 (O_1603,N_49414,N_45192);
or UO_1604 (O_1604,N_45564,N_48374);
nor UO_1605 (O_1605,N_47591,N_47905);
xnor UO_1606 (O_1606,N_48071,N_48793);
xor UO_1607 (O_1607,N_48865,N_49483);
xnor UO_1608 (O_1608,N_48521,N_46954);
nand UO_1609 (O_1609,N_45213,N_49848);
xnor UO_1610 (O_1610,N_47769,N_45249);
nand UO_1611 (O_1611,N_47939,N_45765);
nand UO_1612 (O_1612,N_46825,N_46501);
or UO_1613 (O_1613,N_45122,N_45973);
and UO_1614 (O_1614,N_48014,N_47812);
nand UO_1615 (O_1615,N_45019,N_49158);
and UO_1616 (O_1616,N_49860,N_47091);
xnor UO_1617 (O_1617,N_47852,N_49866);
or UO_1618 (O_1618,N_49464,N_48513);
xnor UO_1619 (O_1619,N_46551,N_45950);
nor UO_1620 (O_1620,N_47396,N_47564);
nor UO_1621 (O_1621,N_46961,N_46917);
and UO_1622 (O_1622,N_48684,N_47850);
and UO_1623 (O_1623,N_48932,N_46448);
and UO_1624 (O_1624,N_45919,N_48631);
nand UO_1625 (O_1625,N_49242,N_46272);
nand UO_1626 (O_1626,N_49650,N_46597);
nor UO_1627 (O_1627,N_46277,N_45949);
xor UO_1628 (O_1628,N_48005,N_48765);
nor UO_1629 (O_1629,N_49597,N_48759);
nand UO_1630 (O_1630,N_49134,N_49042);
nor UO_1631 (O_1631,N_45535,N_46609);
xnor UO_1632 (O_1632,N_49346,N_47078);
nand UO_1633 (O_1633,N_47877,N_49813);
nand UO_1634 (O_1634,N_47327,N_45234);
nand UO_1635 (O_1635,N_48564,N_48550);
nor UO_1636 (O_1636,N_48415,N_46206);
nor UO_1637 (O_1637,N_46299,N_45924);
or UO_1638 (O_1638,N_47355,N_48010);
and UO_1639 (O_1639,N_48743,N_46315);
xnor UO_1640 (O_1640,N_46777,N_47042);
nor UO_1641 (O_1641,N_49088,N_47725);
and UO_1642 (O_1642,N_48095,N_49946);
nor UO_1643 (O_1643,N_49430,N_46940);
xnor UO_1644 (O_1644,N_47490,N_47530);
or UO_1645 (O_1645,N_45591,N_47126);
xnor UO_1646 (O_1646,N_48849,N_45811);
and UO_1647 (O_1647,N_45946,N_45512);
nor UO_1648 (O_1648,N_49412,N_47521);
xnor UO_1649 (O_1649,N_48700,N_48748);
or UO_1650 (O_1650,N_46959,N_48762);
or UO_1651 (O_1651,N_48854,N_45136);
and UO_1652 (O_1652,N_47981,N_45497);
or UO_1653 (O_1653,N_49385,N_46617);
and UO_1654 (O_1654,N_46121,N_47089);
nor UO_1655 (O_1655,N_48312,N_49586);
xnor UO_1656 (O_1656,N_46351,N_49578);
nand UO_1657 (O_1657,N_49407,N_46027);
nand UO_1658 (O_1658,N_48788,N_48070);
and UO_1659 (O_1659,N_48619,N_49150);
and UO_1660 (O_1660,N_46177,N_49604);
nand UO_1661 (O_1661,N_48692,N_45496);
or UO_1662 (O_1662,N_47193,N_49125);
or UO_1663 (O_1663,N_47615,N_45197);
or UO_1664 (O_1664,N_45544,N_48620);
nor UO_1665 (O_1665,N_46201,N_48868);
or UO_1666 (O_1666,N_47498,N_48033);
or UO_1667 (O_1667,N_45910,N_47156);
nand UO_1668 (O_1668,N_49447,N_49754);
or UO_1669 (O_1669,N_47588,N_46725);
nand UO_1670 (O_1670,N_49524,N_47075);
xnor UO_1671 (O_1671,N_45939,N_47495);
nor UO_1672 (O_1672,N_48754,N_46675);
or UO_1673 (O_1673,N_46754,N_46666);
nand UO_1674 (O_1674,N_49551,N_49351);
or UO_1675 (O_1675,N_47473,N_46107);
nand UO_1676 (O_1676,N_49912,N_47825);
and UO_1677 (O_1677,N_47335,N_48768);
xnor UO_1678 (O_1678,N_49630,N_48529);
nor UO_1679 (O_1679,N_49167,N_46168);
nand UO_1680 (O_1680,N_45317,N_48869);
and UO_1681 (O_1681,N_45023,N_46926);
xor UO_1682 (O_1682,N_46023,N_48969);
nand UO_1683 (O_1683,N_47087,N_49636);
or UO_1684 (O_1684,N_49717,N_49198);
nor UO_1685 (O_1685,N_45498,N_46906);
xor UO_1686 (O_1686,N_49410,N_47281);
or UO_1687 (O_1687,N_49723,N_46542);
nor UO_1688 (O_1688,N_48420,N_46471);
nand UO_1689 (O_1689,N_45774,N_47975);
nor UO_1690 (O_1690,N_48680,N_47284);
and UO_1691 (O_1691,N_48674,N_47268);
nor UO_1692 (O_1692,N_45897,N_46330);
xnor UO_1693 (O_1693,N_48767,N_49859);
xnor UO_1694 (O_1694,N_48200,N_46376);
or UO_1695 (O_1695,N_45985,N_48375);
or UO_1696 (O_1696,N_49390,N_47374);
and UO_1697 (O_1697,N_46841,N_46157);
and UO_1698 (O_1698,N_45759,N_46633);
and UO_1699 (O_1699,N_45421,N_49477);
and UO_1700 (O_1700,N_46345,N_46504);
nand UO_1701 (O_1701,N_45070,N_46515);
nor UO_1702 (O_1702,N_47807,N_46492);
nor UO_1703 (O_1703,N_46216,N_46059);
nand UO_1704 (O_1704,N_48126,N_47742);
nor UO_1705 (O_1705,N_47966,N_48354);
or UO_1706 (O_1706,N_49536,N_47409);
nor UO_1707 (O_1707,N_49327,N_46175);
or UO_1708 (O_1708,N_49564,N_48624);
xnor UO_1709 (O_1709,N_46053,N_46148);
nor UO_1710 (O_1710,N_47289,N_47926);
or UO_1711 (O_1711,N_49755,N_45495);
nor UO_1712 (O_1712,N_45476,N_49684);
xnor UO_1713 (O_1713,N_46873,N_47159);
nor UO_1714 (O_1714,N_45336,N_48495);
nand UO_1715 (O_1715,N_45730,N_49612);
nand UO_1716 (O_1716,N_46611,N_47848);
nand UO_1717 (O_1717,N_46806,N_49084);
xor UO_1718 (O_1718,N_49703,N_47377);
nor UO_1719 (O_1719,N_46553,N_47760);
nand UO_1720 (O_1720,N_48526,N_49128);
xor UO_1721 (O_1721,N_49692,N_46493);
and UO_1722 (O_1722,N_47814,N_49648);
or UO_1723 (O_1723,N_47768,N_48490);
or UO_1724 (O_1724,N_45241,N_47516);
or UO_1725 (O_1725,N_46184,N_45457);
or UO_1726 (O_1726,N_48293,N_47240);
xor UO_1727 (O_1727,N_46260,N_46069);
xnor UO_1728 (O_1728,N_46744,N_45009);
or UO_1729 (O_1729,N_49881,N_46139);
and UO_1730 (O_1730,N_48052,N_49804);
or UO_1731 (O_1731,N_49116,N_48507);
xor UO_1732 (O_1732,N_48844,N_49898);
nor UO_1733 (O_1733,N_47310,N_46104);
and UO_1734 (O_1734,N_45454,N_47509);
and UO_1735 (O_1735,N_46967,N_46903);
nand UO_1736 (O_1736,N_49109,N_45932);
nor UO_1737 (O_1737,N_49851,N_49958);
nand UO_1738 (O_1738,N_49297,N_48177);
nor UO_1739 (O_1739,N_48887,N_46097);
nand UO_1740 (O_1740,N_47920,N_49006);
and UO_1741 (O_1741,N_47449,N_47759);
nand UO_1742 (O_1742,N_49499,N_49747);
or UO_1743 (O_1743,N_45648,N_48153);
nand UO_1744 (O_1744,N_48350,N_46576);
and UO_1745 (O_1745,N_45865,N_46714);
and UO_1746 (O_1746,N_49936,N_45716);
nand UO_1747 (O_1747,N_47569,N_46338);
and UO_1748 (O_1748,N_46462,N_45547);
xor UO_1749 (O_1749,N_48333,N_49060);
and UO_1750 (O_1750,N_45348,N_46460);
xor UO_1751 (O_1751,N_46768,N_47413);
nand UO_1752 (O_1752,N_47751,N_48702);
or UO_1753 (O_1753,N_47894,N_46803);
nor UO_1754 (O_1754,N_45775,N_46847);
nand UO_1755 (O_1755,N_47253,N_45042);
nand UO_1756 (O_1756,N_46662,N_48469);
xnor UO_1757 (O_1757,N_49895,N_48028);
xnor UO_1758 (O_1758,N_48411,N_47794);
xnor UO_1759 (O_1759,N_47819,N_45193);
or UO_1760 (O_1760,N_46702,N_48774);
nor UO_1761 (O_1761,N_48990,N_46668);
xor UO_1762 (O_1762,N_47941,N_45743);
and UO_1763 (O_1763,N_49677,N_48662);
and UO_1764 (O_1764,N_48465,N_49460);
or UO_1765 (O_1765,N_47553,N_49402);
nand UO_1766 (O_1766,N_49319,N_46152);
and UO_1767 (O_1767,N_47134,N_45603);
nor UO_1768 (O_1768,N_48496,N_48429);
and UO_1769 (O_1769,N_47334,N_48542);
and UO_1770 (O_1770,N_49073,N_48084);
nor UO_1771 (O_1771,N_45817,N_47831);
or UO_1772 (O_1772,N_49392,N_49872);
or UO_1773 (O_1773,N_46846,N_45948);
xor UO_1774 (O_1774,N_49626,N_48280);
or UO_1775 (O_1775,N_47531,N_45731);
nand UO_1776 (O_1776,N_45171,N_48847);
nor UO_1777 (O_1777,N_45424,N_46887);
nand UO_1778 (O_1778,N_46829,N_45056);
and UO_1779 (O_1779,N_49204,N_46913);
or UO_1780 (O_1780,N_45624,N_47775);
nand UO_1781 (O_1781,N_47373,N_48067);
or UO_1782 (O_1782,N_47371,N_46555);
xnor UO_1783 (O_1783,N_45752,N_45277);
or UO_1784 (O_1784,N_47309,N_48260);
or UO_1785 (O_1785,N_45751,N_47049);
xnor UO_1786 (O_1786,N_47489,N_48385);
xnor UO_1787 (O_1787,N_48669,N_45210);
nand UO_1788 (O_1788,N_49670,N_49710);
and UO_1789 (O_1789,N_47912,N_49997);
nor UO_1790 (O_1790,N_48894,N_47727);
xor UO_1791 (O_1791,N_48591,N_47556);
nor UO_1792 (O_1792,N_46683,N_49873);
and UO_1793 (O_1793,N_49465,N_45686);
or UO_1794 (O_1794,N_49914,N_49329);
nand UO_1795 (O_1795,N_49237,N_49645);
xor UO_1796 (O_1796,N_46313,N_45684);
xnor UO_1797 (O_1797,N_45204,N_46211);
xor UO_1798 (O_1798,N_45286,N_47106);
and UO_1799 (O_1799,N_46494,N_47383);
nor UO_1800 (O_1800,N_45998,N_47332);
or UO_1801 (O_1801,N_46910,N_48410);
nand UO_1802 (O_1802,N_47646,N_46540);
and UO_1803 (O_1803,N_48271,N_46876);
nand UO_1804 (O_1804,N_47737,N_45096);
and UO_1805 (O_1805,N_49622,N_45078);
and UO_1806 (O_1806,N_47333,N_48360);
and UO_1807 (O_1807,N_48850,N_45504);
xnor UO_1808 (O_1808,N_47938,N_49078);
xnor UO_1809 (O_1809,N_46640,N_47039);
or UO_1810 (O_1810,N_47898,N_47763);
nor UO_1811 (O_1811,N_46297,N_46215);
and UO_1812 (O_1812,N_49803,N_49424);
nand UO_1813 (O_1813,N_49485,N_48278);
nand UO_1814 (O_1814,N_49493,N_47111);
nand UO_1815 (O_1815,N_46868,N_46949);
xor UO_1816 (O_1816,N_46481,N_47190);
or UO_1817 (O_1817,N_49119,N_49773);
or UO_1818 (O_1818,N_46647,N_46173);
and UO_1819 (O_1819,N_47499,N_49272);
and UO_1820 (O_1820,N_48554,N_46401);
and UO_1821 (O_1821,N_46436,N_49740);
nand UO_1822 (O_1822,N_48900,N_47023);
or UO_1823 (O_1823,N_48113,N_47002);
nand UO_1824 (O_1824,N_49849,N_49718);
nand UO_1825 (O_1825,N_48749,N_45975);
xnor UO_1826 (O_1826,N_47581,N_49174);
nor UO_1827 (O_1827,N_45584,N_47799);
xor UO_1828 (O_1828,N_47802,N_46429);
nand UO_1829 (O_1829,N_47700,N_45381);
xor UO_1830 (O_1830,N_46706,N_45628);
or UO_1831 (O_1831,N_48491,N_48035);
and UO_1832 (O_1832,N_47464,N_45587);
xnor UO_1833 (O_1833,N_45156,N_46252);
or UO_1834 (O_1834,N_46017,N_49800);
xor UO_1835 (O_1835,N_49205,N_47954);
nor UO_1836 (O_1836,N_45183,N_46775);
xor UO_1837 (O_1837,N_45517,N_48356);
nor UO_1838 (O_1838,N_49573,N_45065);
and UO_1839 (O_1839,N_48655,N_48311);
nand UO_1840 (O_1840,N_48630,N_45344);
or UO_1841 (O_1841,N_49331,N_47008);
or UO_1842 (O_1842,N_45546,N_49364);
and UO_1843 (O_1843,N_48860,N_48644);
or UO_1844 (O_1844,N_49721,N_49436);
or UO_1845 (O_1845,N_47860,N_48473);
nand UO_1846 (O_1846,N_45553,N_45205);
xor UO_1847 (O_1847,N_47143,N_47349);
or UO_1848 (O_1848,N_47503,N_49307);
xnor UO_1849 (O_1849,N_46690,N_45449);
nand UO_1850 (O_1850,N_47515,N_47776);
xnor UO_1851 (O_1851,N_45706,N_49874);
and UO_1852 (O_1852,N_45369,N_47638);
nor UO_1853 (O_1853,N_48519,N_46442);
nor UO_1854 (O_1854,N_45236,N_49081);
or UO_1855 (O_1855,N_49179,N_45058);
nand UO_1856 (O_1856,N_48183,N_49059);
or UO_1857 (O_1857,N_48713,N_47120);
xor UO_1858 (O_1858,N_45047,N_47247);
nand UO_1859 (O_1859,N_45063,N_47570);
xor UO_1860 (O_1860,N_47712,N_47364);
and UO_1861 (O_1861,N_46389,N_47558);
xor UO_1862 (O_1862,N_49295,N_48273);
nor UO_1863 (O_1863,N_45090,N_46809);
nor UO_1864 (O_1864,N_48607,N_47726);
or UO_1865 (O_1865,N_48031,N_45787);
nor UO_1866 (O_1866,N_46220,N_47908);
nand UO_1867 (O_1867,N_45994,N_45137);
or UO_1868 (O_1868,N_49580,N_45882);
xor UO_1869 (O_1869,N_47965,N_47986);
xor UO_1870 (O_1870,N_45914,N_49610);
or UO_1871 (O_1871,N_49380,N_46655);
nor UO_1872 (O_1872,N_46956,N_45703);
and UO_1873 (O_1873,N_46427,N_46637);
or UO_1874 (O_1874,N_45440,N_46888);
or UO_1875 (O_1875,N_46602,N_48665);
nand UO_1876 (O_1876,N_48846,N_48557);
and UO_1877 (O_1877,N_46537,N_45303);
xor UO_1878 (O_1878,N_47176,N_45656);
xor UO_1879 (O_1879,N_47084,N_47256);
nand UO_1880 (O_1880,N_46195,N_46311);
nor UO_1881 (O_1881,N_46969,N_45960);
or UO_1882 (O_1882,N_47580,N_49252);
and UO_1883 (O_1883,N_46629,N_48686);
xor UO_1884 (O_1884,N_46914,N_47466);
nor UO_1885 (O_1885,N_49001,N_45500);
or UO_1886 (O_1886,N_49383,N_48471);
xnor UO_1887 (O_1887,N_45175,N_47346);
or UO_1888 (O_1888,N_46440,N_48434);
or UO_1889 (O_1889,N_46172,N_48902);
and UO_1890 (O_1890,N_49595,N_47269);
and UO_1891 (O_1891,N_46262,N_46600);
or UO_1892 (O_1892,N_45259,N_48840);
xor UO_1893 (O_1893,N_47706,N_47081);
nor UO_1894 (O_1894,N_47406,N_47059);
nor UO_1895 (O_1895,N_49137,N_45460);
nand UO_1896 (O_1896,N_49890,N_48472);
xor UO_1897 (O_1897,N_48922,N_49845);
nand UO_1898 (O_1898,N_46348,N_48909);
nand UO_1899 (O_1899,N_47919,N_45571);
xor UO_1900 (O_1900,N_49271,N_46935);
or UO_1901 (O_1901,N_46736,N_46740);
nand UO_1902 (O_1902,N_47627,N_46770);
and UO_1903 (O_1903,N_46328,N_47437);
nor UO_1904 (O_1904,N_49281,N_46141);
and UO_1905 (O_1905,N_47010,N_49945);
or UO_1906 (O_1906,N_46070,N_46971);
nand UO_1907 (O_1907,N_48478,N_47866);
nor UO_1908 (O_1908,N_49107,N_48751);
nor UO_1909 (O_1909,N_48829,N_49852);
xnor UO_1910 (O_1910,N_47438,N_49627);
nand UO_1911 (O_1911,N_45726,N_46258);
nor UO_1912 (O_1912,N_47178,N_48805);
nand UO_1913 (O_1913,N_48967,N_47722);
or UO_1914 (O_1914,N_47248,N_47035);
or UO_1915 (O_1915,N_46741,N_48074);
xnor UO_1916 (O_1916,N_45937,N_47921);
and UO_1917 (O_1917,N_49949,N_46495);
nand UO_1918 (O_1918,N_45622,N_48442);
xnor UO_1919 (O_1919,N_47928,N_45850);
nor UO_1920 (O_1920,N_46550,N_46294);
nand UO_1921 (O_1921,N_49333,N_45595);
xnor UO_1922 (O_1922,N_45562,N_49292);
or UO_1923 (O_1923,N_48368,N_47017);
nor UO_1924 (O_1924,N_46018,N_49500);
or UO_1925 (O_1925,N_45576,N_45401);
and UO_1926 (O_1926,N_46319,N_48000);
or UO_1927 (O_1927,N_49426,N_46820);
and UO_1928 (O_1928,N_45465,N_49229);
or UO_1929 (O_1929,N_48683,N_48169);
or UO_1930 (O_1930,N_46078,N_45224);
xor UO_1931 (O_1931,N_46339,N_47745);
nand UO_1932 (O_1932,N_45757,N_48167);
nand UO_1933 (O_1933,N_45029,N_47918);
xnor UO_1934 (O_1934,N_48672,N_45922);
and UO_1935 (O_1935,N_48993,N_48598);
nand UO_1936 (O_1936,N_45444,N_45798);
nand UO_1937 (O_1937,N_45174,N_48216);
nand UO_1938 (O_1938,N_45961,N_46533);
or UO_1939 (O_1939,N_49433,N_46881);
xnor UO_1940 (O_1940,N_45954,N_47419);
or UO_1941 (O_1941,N_46248,N_45003);
and UO_1942 (O_1942,N_48628,N_48763);
nor UO_1943 (O_1943,N_46752,N_49857);
nor UO_1944 (O_1944,N_47614,N_46449);
nand UO_1945 (O_1945,N_49188,N_46970);
nand UO_1946 (O_1946,N_48740,N_48770);
xor UO_1947 (O_1947,N_47584,N_48825);
nor UO_1948 (O_1948,N_46253,N_45041);
or UO_1949 (O_1949,N_47756,N_47347);
and UO_1950 (O_1950,N_48436,N_47456);
and UO_1951 (O_1951,N_47316,N_49766);
xnor UO_1952 (O_1952,N_47130,N_46525);
and UO_1953 (O_1953,N_48803,N_45284);
and UO_1954 (O_1954,N_46190,N_47510);
xor UO_1955 (O_1955,N_45745,N_49962);
xnor UO_1956 (O_1956,N_46948,N_47935);
nand UO_1957 (O_1957,N_49209,N_49884);
xnor UO_1958 (O_1958,N_47753,N_48229);
and UO_1959 (O_1959,N_49061,N_48159);
xor UO_1960 (O_1960,N_45446,N_47401);
xnor UO_1961 (O_1961,N_47422,N_46463);
nand UO_1962 (O_1962,N_49372,N_47323);
xnor UO_1963 (O_1963,N_46958,N_49258);
nor UO_1964 (O_1964,N_46943,N_48020);
xor UO_1965 (O_1965,N_48582,N_49212);
xor UO_1966 (O_1966,N_45736,N_49811);
or UO_1967 (O_1967,N_48546,N_45123);
or UO_1968 (O_1968,N_45320,N_47179);
xnor UO_1969 (O_1969,N_48439,N_48184);
nor UO_1970 (O_1970,N_48298,N_49324);
nand UO_1971 (O_1971,N_49805,N_47293);
or UO_1972 (O_1972,N_45981,N_49486);
or UO_1973 (O_1973,N_49735,N_48493);
nand UO_1974 (O_1974,N_46132,N_48623);
xor UO_1975 (O_1975,N_49725,N_45502);
and UO_1976 (O_1976,N_46762,N_48022);
or UO_1977 (O_1977,N_49771,N_45892);
nand UO_1978 (O_1978,N_47618,N_47122);
nor UO_1979 (O_1979,N_49963,N_45326);
or UO_1980 (O_1980,N_48387,N_47924);
xor UO_1981 (O_1981,N_48404,N_48677);
or UO_1982 (O_1982,N_48078,N_45052);
nand UO_1983 (O_1983,N_47583,N_45809);
xor UO_1984 (O_1984,N_47324,N_45345);
and UO_1985 (O_1985,N_48806,N_45075);
and UO_1986 (O_1986,N_49355,N_47946);
xor UO_1987 (O_1987,N_46771,N_47229);
xnor UO_1988 (O_1988,N_47613,N_48553);
xor UO_1989 (O_1989,N_46010,N_47561);
xnor UO_1990 (O_1990,N_45266,N_45203);
xor UO_1991 (O_1991,N_47290,N_48043);
nand UO_1992 (O_1992,N_46374,N_45178);
or UO_1993 (O_1993,N_47806,N_47461);
xnor UO_1994 (O_1994,N_47910,N_49476);
and UO_1995 (O_1995,N_45470,N_45830);
or UO_1996 (O_1996,N_49540,N_46052);
xnor UO_1997 (O_1997,N_45129,N_47132);
and UO_1998 (O_1998,N_46323,N_49427);
xnor UO_1999 (O_1999,N_48001,N_47455);
xnor UO_2000 (O_2000,N_47100,N_45959);
or UO_2001 (O_2001,N_45480,N_46659);
nor UO_2002 (O_2002,N_47771,N_46369);
and UO_2003 (O_2003,N_47578,N_48590);
nor UO_2004 (O_2004,N_47110,N_47141);
nand UO_2005 (O_2005,N_47713,N_46758);
or UO_2006 (O_2006,N_49715,N_48555);
or UO_2007 (O_2007,N_46644,N_46642);
and UO_2008 (O_2008,N_46749,N_46952);
nand UO_2009 (O_2009,N_45501,N_47518);
and UO_2010 (O_2010,N_48928,N_47104);
and UO_2011 (O_2011,N_45223,N_49423);
or UO_2012 (O_2012,N_47551,N_45856);
nand UO_2013 (O_2013,N_49698,N_49117);
and UO_2014 (O_2014,N_46020,N_47534);
nor UO_2015 (O_2015,N_48267,N_47278);
or UO_2016 (O_2016,N_47984,N_45483);
nor UO_2017 (O_2017,N_45157,N_48363);
and UO_2018 (O_2018,N_48731,N_46563);
nand UO_2019 (O_2019,N_49226,N_48408);
nand UO_2020 (O_2020,N_47034,N_48790);
or UO_2021 (O_2021,N_47343,N_45828);
or UO_2022 (O_2022,N_45972,N_49770);
and UO_2023 (O_2023,N_47650,N_48459);
and UO_2024 (O_2024,N_48059,N_49469);
nand UO_2025 (O_2025,N_45848,N_46403);
or UO_2026 (O_2026,N_47188,N_49164);
xor UO_2027 (O_2027,N_47433,N_45120);
nand UO_2028 (O_2028,N_47684,N_45908);
or UO_2029 (O_2029,N_45925,N_49971);
or UO_2030 (O_2030,N_46695,N_48638);
and UO_2031 (O_2031,N_48364,N_49942);
nor UO_2032 (O_2032,N_47874,N_46194);
nand UO_2033 (O_2033,N_49871,N_48040);
nor UO_2034 (O_2034,N_49876,N_45229);
or UO_2035 (O_2035,N_45184,N_46844);
xnor UO_2036 (O_2036,N_48855,N_46548);
and UO_2037 (O_2037,N_49384,N_45378);
nand UO_2038 (O_2038,N_45255,N_47652);
xnor UO_2039 (O_2039,N_48960,N_45389);
nand UO_2040 (O_2040,N_47655,N_46737);
or UO_2041 (O_2041,N_47901,N_49686);
nand UO_2042 (O_2042,N_48249,N_47214);
nor UO_2043 (O_2043,N_47200,N_48982);
xnor UO_2044 (O_2044,N_45812,N_47307);
nor UO_2045 (O_2045,N_48537,N_49025);
and UO_2046 (O_2046,N_49821,N_49161);
or UO_2047 (O_2047,N_45629,N_47185);
nand UO_2048 (O_2048,N_49761,N_49588);
and UO_2049 (O_2049,N_46231,N_49489);
nor UO_2050 (O_2050,N_46854,N_48822);
xnor UO_2051 (O_2051,N_48530,N_45596);
xor UO_2052 (O_2052,N_49505,N_48092);
nand UO_2053 (O_2053,N_49688,N_48107);
xnor UO_2054 (O_2054,N_46165,N_46669);
nor UO_2055 (O_2055,N_45589,N_47610);
and UO_2056 (O_2056,N_49352,N_46151);
nand UO_2057 (O_2057,N_48180,N_48389);
nor UO_2058 (O_2058,N_46383,N_46344);
and UO_2059 (O_2059,N_45777,N_47991);
xor UO_2060 (O_2060,N_48509,N_46341);
nor UO_2061 (O_2061,N_48899,N_49353);
nand UO_2062 (O_2062,N_49541,N_49313);
or UO_2063 (O_2063,N_46266,N_49607);
nor UO_2064 (O_2064,N_45738,N_47246);
or UO_2065 (O_2065,N_46210,N_45271);
xor UO_2066 (O_2066,N_49437,N_49733);
nand UO_2067 (O_2067,N_47649,N_47379);
nand UO_2068 (O_2068,N_45143,N_49734);
nor UO_2069 (O_2069,N_45158,N_47085);
xnor UO_2070 (O_2070,N_49720,N_48309);
and UO_2071 (O_2071,N_48532,N_45185);
nor UO_2072 (O_2072,N_45475,N_46932);
and UO_2073 (O_2073,N_47393,N_49013);
or UO_2074 (O_2074,N_47917,N_49632);
xnor UO_2075 (O_2075,N_49709,N_45138);
or UO_2076 (O_2076,N_47475,N_47254);
and UO_2077 (O_2077,N_45679,N_46407);
and UO_2078 (O_2078,N_49689,N_48151);
nor UO_2079 (O_2079,N_46250,N_46189);
xnor UO_2080 (O_2080,N_46135,N_47694);
xor UO_2081 (O_2081,N_46634,N_48131);
xnor UO_2082 (O_2082,N_47430,N_46812);
and UO_2083 (O_2083,N_48288,N_46622);
xnor UO_2084 (O_2084,N_48053,N_45824);
nor UO_2085 (O_2085,N_46757,N_48339);
or UO_2086 (O_2086,N_49705,N_45704);
and UO_2087 (O_2087,N_47940,N_49022);
nor UO_2088 (O_2088,N_48036,N_45913);
or UO_2089 (O_2089,N_45508,N_45462);
or UO_2090 (O_2090,N_48331,N_48256);
and UO_2091 (O_2091,N_49919,N_48875);
nand UO_2092 (O_2092,N_49827,N_46137);
nand UO_2093 (O_2093,N_49977,N_47142);
nand UO_2094 (O_2094,N_49954,N_47243);
or UO_2095 (O_2095,N_47590,N_49763);
nor UO_2096 (O_2096,N_46832,N_49056);
and UO_2097 (O_2097,N_49863,N_48383);
and UO_2098 (O_2098,N_48154,N_49320);
nand UO_2099 (O_2099,N_46570,N_46334);
nand UO_2100 (O_2100,N_48460,N_49264);
xor UO_2101 (O_2101,N_48578,N_46024);
xnor UO_2102 (O_2102,N_47895,N_49585);
nand UO_2103 (O_2103,N_47118,N_48977);
xor UO_2104 (O_2104,N_49593,N_45604);
nor UO_2105 (O_2105,N_49737,N_46568);
xnor UO_2106 (O_2106,N_49193,N_46769);
xnor UO_2107 (O_2107,N_46404,N_47864);
nand UO_2108 (O_2108,N_45803,N_45133);
or UO_2109 (O_2109,N_48029,N_49132);
nand UO_2110 (O_2110,N_49515,N_49218);
nand UO_2111 (O_2111,N_47028,N_45323);
nor UO_2112 (O_2112,N_47202,N_49080);
xnor UO_2113 (O_2113,N_45274,N_49555);
and UO_2114 (O_2114,N_45538,N_49371);
xnor UO_2115 (O_2115,N_47479,N_49488);
xor UO_2116 (O_2116,N_47528,N_48599);
xor UO_2117 (O_2117,N_49157,N_47911);
nor UO_2118 (O_2118,N_45536,N_47020);
and UO_2119 (O_2119,N_45792,N_49238);
nor UO_2120 (O_2120,N_48597,N_47241);
or UO_2121 (O_2121,N_46982,N_48515);
and UO_2122 (O_2122,N_47702,N_45450);
or UO_2123 (O_2123,N_49004,N_48918);
nand UO_2124 (O_2124,N_45657,N_49824);
nor UO_2125 (O_2125,N_46797,N_45590);
xor UO_2126 (O_2126,N_49011,N_47862);
nand UO_2127 (O_2127,N_48601,N_47803);
nor UO_2128 (O_2128,N_48026,N_45635);
xor UO_2129 (O_2129,N_48535,N_48077);
nor UO_2130 (O_2130,N_46764,N_48220);
nor UO_2131 (O_2131,N_48544,N_47856);
xor UO_2132 (O_2132,N_47716,N_48475);
or UO_2133 (O_2133,N_47741,N_48371);
and UO_2134 (O_2134,N_49902,N_48853);
nand UO_2135 (O_2135,N_48064,N_49459);
nor UO_2136 (O_2136,N_47191,N_48547);
or UO_2137 (O_2137,N_47787,N_45208);
xor UO_2138 (O_2138,N_49055,N_45582);
or UO_2139 (O_2139,N_48114,N_47804);
nor UO_2140 (O_2140,N_46981,N_47224);
or UO_2141 (O_2141,N_48175,N_45212);
nor UO_2142 (O_2142,N_46814,N_45062);
nand UO_2143 (O_2143,N_46496,N_48314);
or UO_2144 (O_2144,N_49802,N_47762);
or UO_2145 (O_2145,N_49354,N_45665);
and UO_2146 (O_2146,N_45293,N_47897);
or UO_2147 (O_2147,N_49836,N_48787);
xnor UO_2148 (O_2148,N_47589,N_48925);
and UO_2149 (O_2149,N_49491,N_45695);
nand UO_2150 (O_2150,N_49560,N_48194);
nor UO_2151 (O_2151,N_46005,N_46701);
and UO_2152 (O_2152,N_46953,N_48336);
nor UO_2153 (O_2153,N_46955,N_49708);
xor UO_2154 (O_2154,N_49606,N_47969);
nand UO_2155 (O_2155,N_49559,N_46824);
or UO_2156 (O_2156,N_45418,N_47482);
nand UO_2157 (O_2157,N_46004,N_45625);
or UO_2158 (O_2158,N_46509,N_45067);
nor UO_2159 (O_2159,N_45490,N_49322);
or UO_2160 (O_2160,N_47822,N_49916);
and UO_2161 (O_2161,N_45674,N_45267);
xnor UO_2162 (O_2162,N_48127,N_49245);
and UO_2163 (O_2163,N_46060,N_46134);
xnor UO_2164 (O_2164,N_49397,N_49123);
or UO_2165 (O_2165,N_48690,N_49966);
and UO_2166 (O_2166,N_47937,N_46355);
nor UO_2167 (O_2167,N_47094,N_48663);
nor UO_2168 (O_2168,N_46857,N_46301);
or UO_2169 (O_2169,N_46006,N_47585);
or UO_2170 (O_2170,N_49753,N_49765);
and UO_2171 (O_2171,N_49249,N_48327);
and UO_2172 (O_2172,N_48450,N_48913);
nand UO_2173 (O_2173,N_49693,N_46664);
nor UO_2174 (O_2174,N_46118,N_48494);
and UO_2175 (O_2175,N_46040,N_49404);
nor UO_2176 (O_2176,N_45996,N_49917);
xnor UO_2177 (O_2177,N_48262,N_49121);
and UO_2178 (O_2178,N_48116,N_48466);
nand UO_2179 (O_2179,N_49343,N_48171);
nand UO_2180 (O_2180,N_49590,N_46951);
xor UO_2181 (O_2181,N_45280,N_49798);
or UO_2182 (O_2182,N_46447,N_45227);
nand UO_2183 (O_2183,N_47434,N_49900);
nor UO_2184 (O_2184,N_49548,N_45976);
xnor UO_2185 (O_2185,N_47005,N_48257);
nor UO_2186 (O_2186,N_46892,N_45040);
nor UO_2187 (O_2187,N_49965,N_46363);
and UO_2188 (O_2188,N_48660,N_45407);
and UO_2189 (O_2189,N_49934,N_45400);
nand UO_2190 (O_2190,N_49233,N_45594);
nor UO_2191 (O_2191,N_48988,N_45173);
nand UO_2192 (O_2192,N_46273,N_46613);
nand UO_2193 (O_2193,N_48480,N_49058);
xnor UO_2194 (O_2194,N_45051,N_49955);
nor UO_2195 (O_2195,N_46146,N_47292);
and UO_2196 (O_2196,N_46728,N_49439);
xor UO_2197 (O_2197,N_49678,N_48225);
nand UO_2198 (O_2198,N_49719,N_48701);
xor UO_2199 (O_2199,N_48065,N_45291);
or UO_2200 (O_2200,N_45448,N_49918);
nor UO_2201 (O_2201,N_46037,N_48323);
and UO_2202 (O_2202,N_47046,N_46336);
and UO_2203 (O_2203,N_47701,N_48320);
xor UO_2204 (O_2204,N_48745,N_47376);
and UO_2205 (O_2205,N_46475,N_46604);
nor UO_2206 (O_2206,N_45349,N_46652);
nor UO_2207 (O_2207,N_49775,N_47868);
and UO_2208 (O_2208,N_47408,N_45305);
and UO_2209 (O_2209,N_47103,N_47019);
or UO_2210 (O_2210,N_47549,N_49159);
xnor UO_2211 (O_2211,N_46335,N_47548);
nor UO_2212 (O_2212,N_47024,N_47619);
and UO_2213 (O_2213,N_46072,N_45727);
xnor UO_2214 (O_2214,N_46034,N_47460);
nand UO_2215 (O_2215,N_45620,N_45499);
nor UO_2216 (O_2216,N_45509,N_45549);
or UO_2217 (O_2217,N_47314,N_48144);
and UO_2218 (O_2218,N_47815,N_45690);
xor UO_2219 (O_2219,N_47425,N_48321);
or UO_2220 (O_2220,N_48437,N_47353);
nor UO_2221 (O_2221,N_46900,N_48266);
nor UO_2222 (O_2222,N_48386,N_49953);
xnor UO_2223 (O_2223,N_47337,N_47678);
nor UO_2224 (O_2224,N_45795,N_45714);
or UO_2225 (O_2225,N_45202,N_49951);
or UO_2226 (O_2226,N_45506,N_47967);
nor UO_2227 (O_2227,N_46918,N_45866);
or UO_2228 (O_2228,N_49360,N_46947);
or UO_2229 (O_2229,N_49288,N_47679);
xnor UO_2230 (O_2230,N_48063,N_47442);
nor UO_2231 (O_2231,N_45135,N_47366);
nand UO_2232 (O_2232,N_45906,N_48637);
nand UO_2233 (O_2233,N_45565,N_46075);
nor UO_2234 (O_2234,N_47197,N_49393);
nor UO_2235 (O_2235,N_45155,N_47125);
nand UO_2236 (O_2236,N_45033,N_48963);
or UO_2237 (O_2237,N_49939,N_47174);
nand UO_2238 (O_2238,N_46709,N_45612);
nand UO_2239 (O_2239,N_47600,N_46993);
or UO_2240 (O_2240,N_47093,N_47446);
xnor UO_2241 (O_2241,N_46225,N_45382);
nor UO_2242 (O_2242,N_45069,N_45639);
nor UO_2243 (O_2243,N_48534,N_49943);
or UO_2244 (O_2244,N_46488,N_49579);
or UO_2245 (O_2245,N_47514,N_48876);
or UO_2246 (O_2246,N_45956,N_45084);
and UO_2247 (O_2247,N_45619,N_47230);
and UO_2248 (O_2248,N_49062,N_47263);
nand UO_2249 (O_2249,N_46589,N_48817);
nand UO_2250 (O_2250,N_47501,N_46946);
xnor UO_2251 (O_2251,N_49223,N_47963);
nor UO_2252 (O_2252,N_45099,N_46085);
xnor UO_2253 (O_2253,N_45217,N_45430);
nor UO_2254 (O_2254,N_48579,N_45516);
xnor UO_2255 (O_2255,N_48231,N_47536);
nor UO_2256 (O_2256,N_48987,N_45253);
xnor UO_2257 (O_2257,N_45634,N_49683);
xor UO_2258 (O_2258,N_48898,N_48023);
and UO_2259 (O_2259,N_49420,N_48671);
and UO_2260 (O_2260,N_48142,N_47397);
nor UO_2261 (O_2261,N_46571,N_45725);
nand UO_2262 (O_2262,N_48722,N_49026);
nand UO_2263 (O_2263,N_45923,N_45015);
nand UO_2264 (O_2264,N_46605,N_48587);
and UO_2265 (O_2265,N_48202,N_49510);
or UO_2266 (O_2266,N_45021,N_49473);
xnor UO_2267 (O_2267,N_46897,N_46271);
and UO_2268 (O_2268,N_47457,N_46785);
or UO_2269 (O_2269,N_49706,N_49339);
nand UO_2270 (O_2270,N_46598,N_45108);
xor UO_2271 (O_2271,N_46278,N_46087);
and UO_2272 (O_2272,N_45645,N_45968);
and UO_2273 (O_2273,N_45869,N_46697);
or UO_2274 (O_2274,N_45872,N_49637);
and UO_2275 (O_2275,N_49478,N_47846);
nand UO_2276 (O_2276,N_49428,N_47872);
xnor UO_2277 (O_2277,N_49869,N_48397);
xnor UO_2278 (O_2278,N_46180,N_49539);
xnor UO_2279 (O_2279,N_46415,N_47194);
or UO_2280 (O_2280,N_46022,N_49047);
nand UO_2281 (O_2281,N_45542,N_49496);
nor UO_2282 (O_2282,N_47541,N_49005);
or UO_2283 (O_2283,N_48226,N_48322);
xnor UO_2284 (O_2284,N_46781,N_48099);
or UO_2285 (O_2285,N_49441,N_48301);
or UO_2286 (O_2286,N_46128,N_47889);
xnor UO_2287 (O_2287,N_45409,N_46109);
nand UO_2288 (O_2288,N_45276,N_46444);
nand UO_2289 (O_2289,N_49330,N_49788);
or UO_2290 (O_2290,N_45769,N_47805);
xor UO_2291 (O_2291,N_47793,N_46856);
and UO_2292 (O_2292,N_49086,N_45240);
nand UO_2293 (O_2293,N_45035,N_45007);
and UO_2294 (O_2294,N_45834,N_45487);
and UO_2295 (O_2295,N_49534,N_48254);
nor UO_2296 (O_2296,N_46579,N_47577);
and UO_2297 (O_2297,N_47887,N_49071);
nor UO_2298 (O_2298,N_47836,N_49983);
or UO_2299 (O_2299,N_47539,N_45037);
xnor UO_2300 (O_2300,N_48566,N_47272);
or UO_2301 (O_2301,N_47688,N_49244);
xor UO_2302 (O_2302,N_46245,N_45394);
xor UO_2303 (O_2303,N_48353,N_45928);
nor UO_2304 (O_2304,N_47491,N_46030);
and UO_2305 (O_2305,N_46880,N_49504);
or UO_2306 (O_2306,N_49639,N_48501);
and UO_2307 (O_2307,N_48959,N_48879);
xor UO_2308 (O_2308,N_49526,N_46145);
or UO_2309 (O_2309,N_46703,N_45086);
nand UO_2310 (O_2310,N_49991,N_47575);
nor UO_2311 (O_2311,N_48265,N_45592);
nand UO_2312 (O_2312,N_46813,N_47435);
nor UO_2313 (O_2313,N_48956,N_47973);
and UO_2314 (O_2314,N_45952,N_48081);
nand UO_2315 (O_2315,N_49089,N_46003);
and UO_2316 (O_2316,N_45898,N_47022);
nor UO_2317 (O_2317,N_46869,N_45433);
or UO_2318 (O_2318,N_49455,N_48347);
or UO_2319 (O_2319,N_49309,N_48211);
nor UO_2320 (O_2320,N_47014,N_45083);
nor UO_2321 (O_2321,N_47136,N_46327);
nand UO_2322 (O_2322,N_48761,N_48082);
xnor UO_2323 (O_2323,N_48248,N_46776);
or UO_2324 (O_2324,N_49618,N_49724);
nand UO_2325 (O_2325,N_45761,N_46889);
xor UO_2326 (O_2326,N_45423,N_49051);
xnor UO_2327 (O_2327,N_45028,N_49370);
xnor UO_2328 (O_2328,N_46259,N_45340);
xnor UO_2329 (O_2329,N_49260,N_46199);
nor UO_2330 (O_2330,N_49931,N_45132);
nand UO_2331 (O_2331,N_49240,N_49546);
xor UO_2332 (O_2332,N_45712,N_48926);
nor UO_2333 (O_2333,N_48626,N_49982);
or UO_2334 (O_2334,N_47069,N_45974);
and UO_2335 (O_2335,N_47691,N_49350);
xnor UO_2336 (O_2336,N_47469,N_47016);
nand UO_2337 (O_2337,N_45300,N_47522);
and UO_2338 (O_2338,N_45963,N_46529);
nor UO_2339 (O_2339,N_48446,N_48815);
xnor UO_2340 (O_2340,N_48516,N_48285);
xor UO_2341 (O_2341,N_49654,N_49379);
and UO_2342 (O_2342,N_47723,N_46646);
and UO_2343 (O_2343,N_47083,N_47821);
nand UO_2344 (O_2344,N_47275,N_45140);
xnor UO_2345 (O_2345,N_46541,N_49367);
xnor UO_2346 (O_2346,N_46864,N_48056);
nor UO_2347 (O_2347,N_45493,N_47440);
and UO_2348 (O_2348,N_47267,N_49998);
nand UO_2349 (O_2349,N_46050,N_46632);
or UO_2350 (O_2350,N_46830,N_45206);
nor UO_2351 (O_2351,N_45523,N_48921);
or UO_2352 (O_2352,N_48196,N_49472);
xnor UO_2353 (O_2353,N_45836,N_45671);
or UO_2354 (O_2354,N_48984,N_48719);
xor UO_2355 (O_2355,N_45361,N_45397);
xor UO_2356 (O_2356,N_48255,N_48935);
xnor UO_2357 (O_2357,N_49875,N_49879);
and UO_2358 (O_2358,N_46872,N_49255);
and UO_2359 (O_2359,N_47097,N_45043);
and UO_2360 (O_2360,N_47301,N_48870);
or UO_2361 (O_2361,N_49467,N_47133);
and UO_2362 (O_2362,N_47209,N_49503);
and UO_2363 (O_2363,N_46439,N_46562);
xnor UO_2364 (O_2364,N_48352,N_47205);
and UO_2365 (O_2365,N_46083,N_48381);
or UO_2366 (O_2366,N_48218,N_46445);
or UO_2367 (O_2367,N_47592,N_48294);
xnor UO_2368 (O_2368,N_47101,N_47165);
or UO_2369 (O_2369,N_49596,N_47571);
and UO_2370 (O_2370,N_47612,N_45689);
and UO_2371 (O_2371,N_47237,N_47659);
xnor UO_2372 (O_2372,N_49136,N_46143);
nand UO_2373 (O_2373,N_49154,N_48104);
xor UO_2374 (O_2374,N_46362,N_49722);
and UO_2375 (O_2375,N_49341,N_47294);
nand UO_2376 (O_2376,N_48236,N_49043);
nand UO_2377 (O_2377,N_48275,N_49561);
nand UO_2378 (O_2378,N_48569,N_45748);
nand UO_2379 (O_2379,N_45050,N_47796);
nor UO_2380 (O_2380,N_49356,N_47184);
xor UO_2381 (O_2381,N_46836,N_48227);
or UO_2382 (O_2382,N_49605,N_47026);
xor UO_2383 (O_2383,N_46098,N_45355);
and UO_2384 (O_2384,N_45785,N_48514);
nand UO_2385 (O_2385,N_48342,N_45520);
and UO_2386 (O_2386,N_45814,N_45883);
or UO_2387 (O_2387,N_47448,N_45800);
nand UO_2388 (O_2388,N_49337,N_47311);
xor UO_2389 (O_2389,N_49888,N_45983);
and UO_2390 (O_2390,N_48239,N_45997);
nor UO_2391 (O_2391,N_48614,N_46453);
or UO_2392 (O_2392,N_49864,N_45221);
xor UO_2393 (O_2393,N_49475,N_45554);
xor UO_2394 (O_2394,N_48484,N_47829);
xnor UO_2395 (O_2395,N_49599,N_45938);
and UO_2396 (O_2396,N_49274,N_49248);
nor UO_2397 (O_2397,N_45292,N_45094);
nor UO_2398 (O_2398,N_47800,N_47252);
xor UO_2399 (O_2399,N_48884,N_46938);
and UO_2400 (O_2400,N_45416,N_47306);
and UO_2401 (O_2401,N_49978,N_47606);
or UO_2402 (O_2402,N_48593,N_46976);
and UO_2403 (O_2403,N_47392,N_47983);
or UO_2404 (O_2404,N_48423,N_47790);
nand UO_2405 (O_2405,N_47361,N_46414);
xor UO_2406 (O_2406,N_45605,N_48836);
or UO_2407 (O_2407,N_46823,N_46007);
or UO_2408 (O_2408,N_46479,N_47507);
xnor UO_2409 (O_2409,N_48781,N_48561);
or UO_2410 (O_2410,N_49820,N_45893);
or UO_2411 (O_2411,N_46499,N_45755);
and UO_2412 (O_2412,N_49365,N_47053);
nor UO_2413 (O_2413,N_49878,N_45327);
nor UO_2414 (O_2414,N_45405,N_46842);
nand UO_2415 (O_2415,N_49894,N_47634);
nand UO_2416 (O_2416,N_49941,N_45560);
nand UO_2417 (O_2417,N_46557,N_46183);
xnor UO_2418 (O_2418,N_46885,N_48736);
nand UO_2419 (O_2419,N_46805,N_47029);
nand UO_2420 (O_2420,N_45319,N_48563);
nor UO_2421 (O_2421,N_45428,N_47352);
nor UO_2422 (O_2422,N_46630,N_45843);
xnor UO_2423 (O_2423,N_46983,N_45802);
xnor UO_2424 (O_2424,N_49927,N_47739);
and UO_2425 (O_2425,N_49925,N_49103);
or UO_2426 (O_2426,N_47389,N_46373);
nand UO_2427 (O_2427,N_48359,N_45393);
nand UO_2428 (O_2428,N_48176,N_49178);
and UO_2429 (O_2429,N_48016,N_45388);
or UO_2430 (O_2430,N_49075,N_49175);
xnor UO_2431 (O_2431,N_48801,N_47598);
xnor UO_2432 (O_2432,N_48886,N_48939);
xnor UO_2433 (O_2433,N_48750,N_49195);
or UO_2434 (O_2434,N_45314,N_45162);
xor UO_2435 (O_2435,N_46994,N_46588);
and UO_2436 (O_2436,N_48215,N_45309);
nor UO_2437 (O_2437,N_48289,N_49808);
xnor UO_2438 (O_2438,N_47559,N_49131);
nor UO_2439 (O_2439,N_45139,N_45567);
nor UO_2440 (O_2440,N_49780,N_46461);
nor UO_2441 (O_2441,N_48366,N_48185);
or UO_2442 (O_2442,N_48609,N_48361);
xor UO_2443 (O_2443,N_46282,N_47060);
xor UO_2444 (O_2444,N_45720,N_48533);
and UO_2445 (O_2445,N_49817,N_46158);
nor UO_2446 (O_2446,N_49358,N_46419);
nand UO_2447 (O_2447,N_47481,N_46304);
and UO_2448 (O_2448,N_48568,N_48708);
nand UO_2449 (O_2449,N_48524,N_45055);
and UO_2450 (O_2450,N_49967,N_49314);
nand UO_2451 (O_2451,N_49401,N_45851);
or UO_2452 (O_2452,N_45947,N_45682);
nor UO_2453 (O_2453,N_45190,N_46546);
nor UO_2454 (O_2454,N_49666,N_47410);
nand UO_2455 (O_2455,N_48705,N_49304);
or UO_2456 (O_2456,N_49413,N_49148);
and UO_2457 (O_2457,N_45282,N_48538);
and UO_2458 (O_2458,N_48284,N_45429);
nand UO_2459 (O_2459,N_48952,N_46944);
nor UO_2460 (O_2460,N_45461,N_48205);
nand UO_2461 (O_2461,N_45601,N_48193);
nor UO_2462 (O_2462,N_47362,N_47683);
nand UO_2463 (O_2463,N_45621,N_46129);
xnor UO_2464 (O_2464,N_45678,N_45165);
or UO_2465 (O_2465,N_45728,N_48570);
xnor UO_2466 (O_2466,N_48941,N_46931);
nor UO_2467 (O_2467,N_49122,N_48667);
and UO_2468 (O_2468,N_48813,N_49587);
or UO_2469 (O_2469,N_46595,N_45228);
nor UO_2470 (O_2470,N_48699,N_48462);
xor UO_2471 (O_2471,N_49613,N_49243);
nor UO_2472 (O_2472,N_46753,N_47238);
nor UO_2473 (O_2473,N_45046,N_45237);
nor UO_2474 (O_2474,N_46110,N_45102);
or UO_2475 (O_2475,N_47262,N_47797);
xnor UO_2476 (O_2476,N_46791,N_48334);
xnor UO_2477 (O_2477,N_45521,N_45700);
xor UO_2478 (O_2478,N_47890,N_49257);
xor UO_2479 (O_2479,N_47813,N_49032);
nand UO_2480 (O_2480,N_46628,N_49124);
and UO_2481 (O_2481,N_49096,N_48181);
nor UO_2482 (O_2482,N_45561,N_47744);
xnor UO_2483 (O_2483,N_48338,N_48880);
xor UO_2484 (O_2484,N_48652,N_49482);
or UO_2485 (O_2485,N_48079,N_46734);
or UO_2486 (O_2486,N_46092,N_47673);
or UO_2487 (O_2487,N_45026,N_45001);
nor UO_2488 (O_2488,N_46594,N_48098);
xnor UO_2489 (O_2489,N_47158,N_47711);
or UO_2490 (O_2490,N_48615,N_48706);
and UO_2491 (O_2491,N_45806,N_47052);
xnor UO_2492 (O_2492,N_49373,N_48015);
and UO_2493 (O_2493,N_46580,N_46421);
xnor UO_2494 (O_2494,N_45172,N_47893);
nor UO_2495 (O_2495,N_48775,N_48816);
and UO_2496 (O_2496,N_49023,N_45363);
or UO_2497 (O_2497,N_48682,N_49809);
and UO_2498 (O_2498,N_47761,N_45330);
and UO_2499 (O_2499,N_47166,N_49675);
and UO_2500 (O_2500,N_48326,N_49729);
nand UO_2501 (O_2501,N_46320,N_48722);
xor UO_2502 (O_2502,N_45273,N_45323);
xnor UO_2503 (O_2503,N_45573,N_46783);
or UO_2504 (O_2504,N_45514,N_47491);
and UO_2505 (O_2505,N_48214,N_48185);
or UO_2506 (O_2506,N_46424,N_49006);
nand UO_2507 (O_2507,N_48215,N_46368);
nor UO_2508 (O_2508,N_48795,N_46423);
nor UO_2509 (O_2509,N_45174,N_47255);
xnor UO_2510 (O_2510,N_45818,N_49409);
and UO_2511 (O_2511,N_47620,N_47484);
and UO_2512 (O_2512,N_49674,N_49916);
and UO_2513 (O_2513,N_49595,N_46175);
nand UO_2514 (O_2514,N_47069,N_45822);
and UO_2515 (O_2515,N_48626,N_47944);
nor UO_2516 (O_2516,N_49550,N_47106);
or UO_2517 (O_2517,N_47473,N_46402);
and UO_2518 (O_2518,N_49237,N_47147);
or UO_2519 (O_2519,N_45006,N_48965);
and UO_2520 (O_2520,N_45968,N_48141);
nand UO_2521 (O_2521,N_46609,N_48849);
and UO_2522 (O_2522,N_49595,N_47117);
xor UO_2523 (O_2523,N_47480,N_46528);
and UO_2524 (O_2524,N_48381,N_49576);
or UO_2525 (O_2525,N_47382,N_46128);
nor UO_2526 (O_2526,N_49987,N_47693);
nor UO_2527 (O_2527,N_49396,N_46417);
xnor UO_2528 (O_2528,N_47773,N_48857);
or UO_2529 (O_2529,N_46520,N_46791);
or UO_2530 (O_2530,N_45253,N_48637);
nand UO_2531 (O_2531,N_48346,N_45156);
or UO_2532 (O_2532,N_47123,N_47892);
nor UO_2533 (O_2533,N_48351,N_46016);
xnor UO_2534 (O_2534,N_49274,N_46260);
and UO_2535 (O_2535,N_46032,N_47015);
or UO_2536 (O_2536,N_46325,N_46436);
or UO_2537 (O_2537,N_49343,N_45122);
nor UO_2538 (O_2538,N_46866,N_46088);
or UO_2539 (O_2539,N_49583,N_45388);
xor UO_2540 (O_2540,N_47074,N_47315);
nor UO_2541 (O_2541,N_46618,N_46755);
or UO_2542 (O_2542,N_49764,N_48626);
or UO_2543 (O_2543,N_49271,N_47583);
and UO_2544 (O_2544,N_45956,N_45820);
nor UO_2545 (O_2545,N_48613,N_47080);
nor UO_2546 (O_2546,N_47800,N_46868);
nor UO_2547 (O_2547,N_47353,N_45620);
nor UO_2548 (O_2548,N_48757,N_49516);
or UO_2549 (O_2549,N_47693,N_49297);
xor UO_2550 (O_2550,N_49003,N_46182);
nor UO_2551 (O_2551,N_45374,N_49142);
or UO_2552 (O_2552,N_49246,N_46161);
nor UO_2553 (O_2553,N_47241,N_47616);
nand UO_2554 (O_2554,N_47286,N_47822);
xor UO_2555 (O_2555,N_46105,N_45969);
xnor UO_2556 (O_2556,N_49988,N_48716);
or UO_2557 (O_2557,N_48200,N_46175);
or UO_2558 (O_2558,N_48119,N_48159);
nor UO_2559 (O_2559,N_45440,N_46130);
and UO_2560 (O_2560,N_45799,N_47314);
nand UO_2561 (O_2561,N_48142,N_47186);
xnor UO_2562 (O_2562,N_49854,N_48015);
or UO_2563 (O_2563,N_47663,N_49002);
nor UO_2564 (O_2564,N_47087,N_46606);
nor UO_2565 (O_2565,N_45904,N_47779);
or UO_2566 (O_2566,N_49595,N_49955);
nor UO_2567 (O_2567,N_48775,N_46278);
nor UO_2568 (O_2568,N_47985,N_49235);
and UO_2569 (O_2569,N_49138,N_46980);
nand UO_2570 (O_2570,N_46283,N_49095);
and UO_2571 (O_2571,N_46451,N_47999);
or UO_2572 (O_2572,N_45000,N_48892);
or UO_2573 (O_2573,N_47443,N_49335);
xor UO_2574 (O_2574,N_46706,N_45711);
xnor UO_2575 (O_2575,N_49977,N_45930);
or UO_2576 (O_2576,N_48526,N_48365);
nand UO_2577 (O_2577,N_49952,N_49093);
and UO_2578 (O_2578,N_47063,N_48324);
xor UO_2579 (O_2579,N_48599,N_45780);
xor UO_2580 (O_2580,N_45154,N_49025);
xor UO_2581 (O_2581,N_47369,N_47352);
xnor UO_2582 (O_2582,N_49822,N_49949);
or UO_2583 (O_2583,N_46829,N_46529);
or UO_2584 (O_2584,N_46773,N_49117);
xor UO_2585 (O_2585,N_47713,N_47557);
nor UO_2586 (O_2586,N_46145,N_45624);
nand UO_2587 (O_2587,N_47164,N_47382);
or UO_2588 (O_2588,N_45664,N_48368);
nand UO_2589 (O_2589,N_48404,N_48871);
nor UO_2590 (O_2590,N_49146,N_45934);
and UO_2591 (O_2591,N_46729,N_49261);
nor UO_2592 (O_2592,N_46283,N_46061);
nand UO_2593 (O_2593,N_48017,N_49640);
and UO_2594 (O_2594,N_47182,N_49753);
nor UO_2595 (O_2595,N_49532,N_46098);
or UO_2596 (O_2596,N_46471,N_47225);
nand UO_2597 (O_2597,N_45410,N_47228);
nand UO_2598 (O_2598,N_45402,N_48750);
xor UO_2599 (O_2599,N_47831,N_45498);
nor UO_2600 (O_2600,N_45570,N_45431);
nor UO_2601 (O_2601,N_47621,N_48622);
nand UO_2602 (O_2602,N_47934,N_45640);
or UO_2603 (O_2603,N_46953,N_49460);
nand UO_2604 (O_2604,N_46378,N_49454);
nor UO_2605 (O_2605,N_47554,N_48025);
nor UO_2606 (O_2606,N_47735,N_48714);
nor UO_2607 (O_2607,N_45746,N_49183);
nand UO_2608 (O_2608,N_47403,N_49143);
nor UO_2609 (O_2609,N_45252,N_47013);
or UO_2610 (O_2610,N_47320,N_47804);
xor UO_2611 (O_2611,N_45356,N_45914);
or UO_2612 (O_2612,N_49913,N_46218);
or UO_2613 (O_2613,N_49866,N_45220);
nor UO_2614 (O_2614,N_46276,N_45789);
or UO_2615 (O_2615,N_45207,N_49270);
xnor UO_2616 (O_2616,N_47381,N_47548);
or UO_2617 (O_2617,N_47924,N_48272);
xor UO_2618 (O_2618,N_47766,N_46225);
xnor UO_2619 (O_2619,N_48933,N_45421);
nor UO_2620 (O_2620,N_49771,N_48251);
or UO_2621 (O_2621,N_47257,N_47234);
nor UO_2622 (O_2622,N_46833,N_46138);
nand UO_2623 (O_2623,N_46767,N_48234);
xnor UO_2624 (O_2624,N_46724,N_45364);
and UO_2625 (O_2625,N_49961,N_45706);
nor UO_2626 (O_2626,N_45605,N_45206);
xnor UO_2627 (O_2627,N_49118,N_48124);
xnor UO_2628 (O_2628,N_47668,N_46305);
nor UO_2629 (O_2629,N_46545,N_46345);
xor UO_2630 (O_2630,N_48744,N_47644);
or UO_2631 (O_2631,N_45795,N_48598);
and UO_2632 (O_2632,N_47643,N_49441);
and UO_2633 (O_2633,N_48992,N_48095);
nor UO_2634 (O_2634,N_47126,N_46970);
xnor UO_2635 (O_2635,N_45868,N_49999);
nor UO_2636 (O_2636,N_46428,N_48193);
nand UO_2637 (O_2637,N_49756,N_45673);
or UO_2638 (O_2638,N_46563,N_48779);
xnor UO_2639 (O_2639,N_49166,N_45467);
nand UO_2640 (O_2640,N_49940,N_49413);
and UO_2641 (O_2641,N_48223,N_48968);
or UO_2642 (O_2642,N_46587,N_49385);
nand UO_2643 (O_2643,N_45790,N_49206);
xnor UO_2644 (O_2644,N_46127,N_45219);
nor UO_2645 (O_2645,N_49576,N_47832);
and UO_2646 (O_2646,N_45733,N_48634);
and UO_2647 (O_2647,N_45315,N_46783);
nor UO_2648 (O_2648,N_48748,N_45128);
or UO_2649 (O_2649,N_45416,N_49863);
xor UO_2650 (O_2650,N_45280,N_49257);
and UO_2651 (O_2651,N_47810,N_45950);
nor UO_2652 (O_2652,N_48791,N_45540);
and UO_2653 (O_2653,N_45689,N_45250);
nand UO_2654 (O_2654,N_48191,N_45928);
nor UO_2655 (O_2655,N_49754,N_45154);
and UO_2656 (O_2656,N_49662,N_45921);
and UO_2657 (O_2657,N_48519,N_45424);
nor UO_2658 (O_2658,N_48570,N_46952);
xor UO_2659 (O_2659,N_46116,N_49388);
nor UO_2660 (O_2660,N_46307,N_49892);
or UO_2661 (O_2661,N_49269,N_45977);
nor UO_2662 (O_2662,N_48731,N_49819);
or UO_2663 (O_2663,N_49228,N_46108);
nand UO_2664 (O_2664,N_48388,N_48995);
nor UO_2665 (O_2665,N_49213,N_45956);
xnor UO_2666 (O_2666,N_46335,N_49608);
nand UO_2667 (O_2667,N_48194,N_48008);
nor UO_2668 (O_2668,N_45962,N_45717);
nand UO_2669 (O_2669,N_48975,N_48101);
xnor UO_2670 (O_2670,N_48851,N_46686);
xor UO_2671 (O_2671,N_47383,N_45038);
nor UO_2672 (O_2672,N_47490,N_49389);
xnor UO_2673 (O_2673,N_47767,N_47891);
and UO_2674 (O_2674,N_48446,N_47866);
nand UO_2675 (O_2675,N_45250,N_46662);
nand UO_2676 (O_2676,N_47760,N_46517);
nor UO_2677 (O_2677,N_49744,N_46714);
and UO_2678 (O_2678,N_48847,N_46808);
nand UO_2679 (O_2679,N_45184,N_46285);
nand UO_2680 (O_2680,N_49582,N_46661);
xnor UO_2681 (O_2681,N_47524,N_49453);
nand UO_2682 (O_2682,N_49334,N_48652);
nand UO_2683 (O_2683,N_46360,N_47741);
nand UO_2684 (O_2684,N_45711,N_47927);
or UO_2685 (O_2685,N_47305,N_47115);
or UO_2686 (O_2686,N_46604,N_47564);
or UO_2687 (O_2687,N_46752,N_46333);
or UO_2688 (O_2688,N_48260,N_47957);
nor UO_2689 (O_2689,N_46170,N_48925);
and UO_2690 (O_2690,N_47989,N_47371);
and UO_2691 (O_2691,N_49278,N_48466);
nand UO_2692 (O_2692,N_49751,N_46727);
and UO_2693 (O_2693,N_48732,N_46521);
nand UO_2694 (O_2694,N_46198,N_49225);
nand UO_2695 (O_2695,N_46340,N_45876);
or UO_2696 (O_2696,N_48317,N_46887);
nand UO_2697 (O_2697,N_48378,N_49519);
nand UO_2698 (O_2698,N_45772,N_45768);
xor UO_2699 (O_2699,N_46367,N_47911);
nor UO_2700 (O_2700,N_46121,N_46786);
nor UO_2701 (O_2701,N_48361,N_45207);
xor UO_2702 (O_2702,N_45031,N_47227);
and UO_2703 (O_2703,N_47009,N_46652);
nor UO_2704 (O_2704,N_48999,N_46633);
and UO_2705 (O_2705,N_46635,N_45203);
nor UO_2706 (O_2706,N_46074,N_45701);
and UO_2707 (O_2707,N_45505,N_48102);
xnor UO_2708 (O_2708,N_46355,N_49088);
xor UO_2709 (O_2709,N_49531,N_47559);
or UO_2710 (O_2710,N_45521,N_47881);
and UO_2711 (O_2711,N_45513,N_48079);
or UO_2712 (O_2712,N_46042,N_48419);
or UO_2713 (O_2713,N_46992,N_48792);
nor UO_2714 (O_2714,N_48216,N_46275);
nand UO_2715 (O_2715,N_45483,N_46921);
nor UO_2716 (O_2716,N_46719,N_49819);
and UO_2717 (O_2717,N_49827,N_49392);
xor UO_2718 (O_2718,N_45878,N_45479);
or UO_2719 (O_2719,N_47558,N_46912);
nand UO_2720 (O_2720,N_49271,N_46623);
xor UO_2721 (O_2721,N_45061,N_48517);
or UO_2722 (O_2722,N_46463,N_48032);
or UO_2723 (O_2723,N_48083,N_45260);
or UO_2724 (O_2724,N_47332,N_45672);
nand UO_2725 (O_2725,N_49000,N_48890);
nor UO_2726 (O_2726,N_47751,N_48411);
or UO_2727 (O_2727,N_48903,N_48126);
or UO_2728 (O_2728,N_49221,N_45262);
xnor UO_2729 (O_2729,N_49303,N_47738);
and UO_2730 (O_2730,N_47654,N_49765);
or UO_2731 (O_2731,N_46826,N_47402);
or UO_2732 (O_2732,N_46861,N_48120);
nor UO_2733 (O_2733,N_49621,N_48408);
xor UO_2734 (O_2734,N_45603,N_48869);
nand UO_2735 (O_2735,N_48436,N_45040);
nand UO_2736 (O_2736,N_47237,N_48905);
nor UO_2737 (O_2737,N_49942,N_48483);
or UO_2738 (O_2738,N_47730,N_45803);
nor UO_2739 (O_2739,N_45521,N_48788);
and UO_2740 (O_2740,N_49958,N_48150);
xor UO_2741 (O_2741,N_46328,N_48770);
nand UO_2742 (O_2742,N_45550,N_49678);
nand UO_2743 (O_2743,N_46299,N_46236);
nor UO_2744 (O_2744,N_47857,N_47793);
xor UO_2745 (O_2745,N_47266,N_48799);
nand UO_2746 (O_2746,N_49938,N_47352);
nand UO_2747 (O_2747,N_45840,N_47212);
or UO_2748 (O_2748,N_45274,N_48450);
nand UO_2749 (O_2749,N_47236,N_49568);
xor UO_2750 (O_2750,N_45410,N_48520);
or UO_2751 (O_2751,N_49184,N_49352);
nor UO_2752 (O_2752,N_45000,N_46094);
or UO_2753 (O_2753,N_49898,N_48960);
xor UO_2754 (O_2754,N_49605,N_45520);
xor UO_2755 (O_2755,N_47551,N_49915);
and UO_2756 (O_2756,N_49686,N_49348);
or UO_2757 (O_2757,N_45905,N_46746);
and UO_2758 (O_2758,N_49106,N_46469);
and UO_2759 (O_2759,N_45298,N_49561);
and UO_2760 (O_2760,N_48039,N_48916);
and UO_2761 (O_2761,N_47418,N_48674);
nor UO_2762 (O_2762,N_48559,N_46004);
nand UO_2763 (O_2763,N_47051,N_45413);
nand UO_2764 (O_2764,N_49041,N_49605);
nand UO_2765 (O_2765,N_47868,N_47517);
xor UO_2766 (O_2766,N_48573,N_45171);
xor UO_2767 (O_2767,N_47112,N_49124);
xor UO_2768 (O_2768,N_46224,N_46103);
and UO_2769 (O_2769,N_45831,N_45991);
xnor UO_2770 (O_2770,N_45795,N_45168);
and UO_2771 (O_2771,N_48561,N_46010);
nor UO_2772 (O_2772,N_46120,N_47109);
nor UO_2773 (O_2773,N_47486,N_48336);
or UO_2774 (O_2774,N_48800,N_45622);
xnor UO_2775 (O_2775,N_45066,N_48418);
nor UO_2776 (O_2776,N_47126,N_46120);
or UO_2777 (O_2777,N_49368,N_48869);
xnor UO_2778 (O_2778,N_48708,N_45452);
or UO_2779 (O_2779,N_48265,N_47231);
or UO_2780 (O_2780,N_47066,N_45223);
nor UO_2781 (O_2781,N_49443,N_46049);
nand UO_2782 (O_2782,N_49407,N_45989);
and UO_2783 (O_2783,N_46901,N_46677);
nor UO_2784 (O_2784,N_46641,N_46627);
nor UO_2785 (O_2785,N_45206,N_45293);
nand UO_2786 (O_2786,N_46103,N_49535);
or UO_2787 (O_2787,N_48482,N_45780);
or UO_2788 (O_2788,N_45441,N_47299);
and UO_2789 (O_2789,N_47760,N_46687);
and UO_2790 (O_2790,N_49721,N_49093);
or UO_2791 (O_2791,N_48212,N_49512);
and UO_2792 (O_2792,N_46006,N_49831);
and UO_2793 (O_2793,N_45460,N_48640);
xor UO_2794 (O_2794,N_47911,N_46408);
nor UO_2795 (O_2795,N_46334,N_47061);
or UO_2796 (O_2796,N_49807,N_46627);
xnor UO_2797 (O_2797,N_45162,N_49553);
and UO_2798 (O_2798,N_47240,N_48798);
xnor UO_2799 (O_2799,N_49719,N_49955);
and UO_2800 (O_2800,N_46166,N_49333);
or UO_2801 (O_2801,N_47916,N_48362);
nor UO_2802 (O_2802,N_49939,N_47689);
xor UO_2803 (O_2803,N_46013,N_46231);
nand UO_2804 (O_2804,N_49075,N_49702);
and UO_2805 (O_2805,N_47732,N_48625);
xor UO_2806 (O_2806,N_46314,N_46807);
nand UO_2807 (O_2807,N_45819,N_48055);
or UO_2808 (O_2808,N_47017,N_45447);
and UO_2809 (O_2809,N_47080,N_46534);
nor UO_2810 (O_2810,N_47149,N_47810);
nand UO_2811 (O_2811,N_45775,N_49055);
and UO_2812 (O_2812,N_47416,N_46699);
xnor UO_2813 (O_2813,N_45098,N_46533);
and UO_2814 (O_2814,N_48541,N_49603);
or UO_2815 (O_2815,N_49795,N_45962);
nand UO_2816 (O_2816,N_46281,N_49971);
nor UO_2817 (O_2817,N_45828,N_47006);
nand UO_2818 (O_2818,N_47583,N_46206);
or UO_2819 (O_2819,N_48239,N_48331);
xor UO_2820 (O_2820,N_45044,N_47939);
nor UO_2821 (O_2821,N_45881,N_48558);
nor UO_2822 (O_2822,N_46722,N_49081);
and UO_2823 (O_2823,N_47066,N_49674);
or UO_2824 (O_2824,N_46691,N_49622);
and UO_2825 (O_2825,N_45446,N_45488);
nand UO_2826 (O_2826,N_48866,N_49401);
nor UO_2827 (O_2827,N_47808,N_46044);
nand UO_2828 (O_2828,N_45218,N_49524);
or UO_2829 (O_2829,N_46365,N_49270);
xor UO_2830 (O_2830,N_45951,N_45708);
nand UO_2831 (O_2831,N_47563,N_47089);
and UO_2832 (O_2832,N_46067,N_45176);
and UO_2833 (O_2833,N_47137,N_45707);
and UO_2834 (O_2834,N_45532,N_48098);
and UO_2835 (O_2835,N_47405,N_45491);
nor UO_2836 (O_2836,N_49480,N_48646);
xnor UO_2837 (O_2837,N_48398,N_46028);
and UO_2838 (O_2838,N_49236,N_45988);
nor UO_2839 (O_2839,N_48882,N_46156);
nand UO_2840 (O_2840,N_49878,N_46278);
or UO_2841 (O_2841,N_49828,N_49346);
xor UO_2842 (O_2842,N_48825,N_46327);
nand UO_2843 (O_2843,N_48368,N_49486);
xnor UO_2844 (O_2844,N_46748,N_46219);
and UO_2845 (O_2845,N_46044,N_47851);
nand UO_2846 (O_2846,N_47033,N_46095);
nand UO_2847 (O_2847,N_48751,N_45658);
nor UO_2848 (O_2848,N_49788,N_49297);
xor UO_2849 (O_2849,N_47039,N_45711);
and UO_2850 (O_2850,N_49525,N_46923);
or UO_2851 (O_2851,N_49449,N_45637);
nor UO_2852 (O_2852,N_49778,N_49374);
or UO_2853 (O_2853,N_46593,N_48111);
or UO_2854 (O_2854,N_48103,N_48555);
or UO_2855 (O_2855,N_46852,N_46690);
and UO_2856 (O_2856,N_49171,N_49513);
nor UO_2857 (O_2857,N_47147,N_45718);
nand UO_2858 (O_2858,N_49833,N_48194);
and UO_2859 (O_2859,N_47234,N_46688);
or UO_2860 (O_2860,N_49362,N_47916);
nand UO_2861 (O_2861,N_45626,N_48102);
or UO_2862 (O_2862,N_49334,N_45263);
xnor UO_2863 (O_2863,N_48463,N_47135);
nand UO_2864 (O_2864,N_45982,N_49228);
and UO_2865 (O_2865,N_46149,N_47618);
or UO_2866 (O_2866,N_47014,N_48981);
nand UO_2867 (O_2867,N_48159,N_47219);
and UO_2868 (O_2868,N_48245,N_47739);
nand UO_2869 (O_2869,N_46899,N_45020);
or UO_2870 (O_2870,N_49933,N_48553);
and UO_2871 (O_2871,N_48092,N_46821);
xor UO_2872 (O_2872,N_49667,N_47165);
xnor UO_2873 (O_2873,N_48049,N_47509);
xor UO_2874 (O_2874,N_47161,N_46204);
nor UO_2875 (O_2875,N_48411,N_48444);
xnor UO_2876 (O_2876,N_46860,N_46203);
and UO_2877 (O_2877,N_45057,N_47303);
or UO_2878 (O_2878,N_49667,N_49802);
nand UO_2879 (O_2879,N_47181,N_45077);
nand UO_2880 (O_2880,N_47124,N_45712);
nor UO_2881 (O_2881,N_48101,N_49728);
xor UO_2882 (O_2882,N_49539,N_45696);
nand UO_2883 (O_2883,N_49887,N_49917);
or UO_2884 (O_2884,N_47436,N_45592);
nand UO_2885 (O_2885,N_47796,N_46261);
xor UO_2886 (O_2886,N_49237,N_45706);
nand UO_2887 (O_2887,N_46967,N_48347);
xor UO_2888 (O_2888,N_49280,N_49123);
xor UO_2889 (O_2889,N_47693,N_46109);
nand UO_2890 (O_2890,N_47040,N_46178);
or UO_2891 (O_2891,N_47359,N_47638);
or UO_2892 (O_2892,N_49047,N_46162);
xor UO_2893 (O_2893,N_48214,N_46182);
nor UO_2894 (O_2894,N_47301,N_46694);
nand UO_2895 (O_2895,N_48718,N_46296);
and UO_2896 (O_2896,N_47035,N_45036);
and UO_2897 (O_2897,N_49999,N_48625);
or UO_2898 (O_2898,N_49949,N_45034);
nand UO_2899 (O_2899,N_48813,N_49033);
nor UO_2900 (O_2900,N_48733,N_47647);
or UO_2901 (O_2901,N_49568,N_45082);
xor UO_2902 (O_2902,N_49078,N_45447);
and UO_2903 (O_2903,N_48479,N_46700);
nand UO_2904 (O_2904,N_45805,N_48969);
and UO_2905 (O_2905,N_49856,N_45169);
and UO_2906 (O_2906,N_49700,N_49311);
xor UO_2907 (O_2907,N_47352,N_48815);
nor UO_2908 (O_2908,N_49688,N_49577);
and UO_2909 (O_2909,N_48476,N_46653);
xnor UO_2910 (O_2910,N_48757,N_47142);
or UO_2911 (O_2911,N_45677,N_45303);
xor UO_2912 (O_2912,N_45726,N_46529);
nand UO_2913 (O_2913,N_48677,N_46493);
or UO_2914 (O_2914,N_49081,N_45504);
and UO_2915 (O_2915,N_45216,N_48541);
nand UO_2916 (O_2916,N_46700,N_48692);
nor UO_2917 (O_2917,N_49904,N_47187);
and UO_2918 (O_2918,N_47953,N_46397);
nand UO_2919 (O_2919,N_47088,N_47391);
nand UO_2920 (O_2920,N_46536,N_49242);
xnor UO_2921 (O_2921,N_49191,N_48146);
xnor UO_2922 (O_2922,N_47342,N_47417);
xnor UO_2923 (O_2923,N_47424,N_45159);
or UO_2924 (O_2924,N_47170,N_45415);
nand UO_2925 (O_2925,N_45064,N_48213);
nor UO_2926 (O_2926,N_49654,N_46619);
nand UO_2927 (O_2927,N_47759,N_46713);
and UO_2928 (O_2928,N_47290,N_45630);
or UO_2929 (O_2929,N_45804,N_47747);
xor UO_2930 (O_2930,N_46950,N_46518);
xor UO_2931 (O_2931,N_49506,N_47181);
and UO_2932 (O_2932,N_46139,N_48671);
or UO_2933 (O_2933,N_48199,N_47224);
and UO_2934 (O_2934,N_46063,N_49735);
or UO_2935 (O_2935,N_45812,N_45201);
xor UO_2936 (O_2936,N_49176,N_45779);
nand UO_2937 (O_2937,N_48588,N_49870);
nor UO_2938 (O_2938,N_45041,N_48179);
or UO_2939 (O_2939,N_45017,N_48952);
nor UO_2940 (O_2940,N_48491,N_45842);
and UO_2941 (O_2941,N_45346,N_49320);
or UO_2942 (O_2942,N_48182,N_49553);
nand UO_2943 (O_2943,N_48984,N_49878);
xor UO_2944 (O_2944,N_47410,N_48104);
and UO_2945 (O_2945,N_46172,N_48977);
nand UO_2946 (O_2946,N_47496,N_48016);
nand UO_2947 (O_2947,N_46936,N_49476);
and UO_2948 (O_2948,N_47069,N_47047);
or UO_2949 (O_2949,N_48848,N_48562);
and UO_2950 (O_2950,N_46573,N_47801);
or UO_2951 (O_2951,N_47460,N_47745);
and UO_2952 (O_2952,N_49839,N_49336);
and UO_2953 (O_2953,N_46040,N_48581);
and UO_2954 (O_2954,N_47059,N_46811);
xor UO_2955 (O_2955,N_46261,N_47544);
or UO_2956 (O_2956,N_49021,N_47060);
xnor UO_2957 (O_2957,N_48464,N_47298);
nor UO_2958 (O_2958,N_47739,N_49194);
or UO_2959 (O_2959,N_45576,N_46616);
xor UO_2960 (O_2960,N_45068,N_48434);
nand UO_2961 (O_2961,N_46643,N_48045);
or UO_2962 (O_2962,N_47546,N_46366);
xnor UO_2963 (O_2963,N_48027,N_45165);
or UO_2964 (O_2964,N_49004,N_45560);
nand UO_2965 (O_2965,N_47095,N_45188);
and UO_2966 (O_2966,N_48929,N_49465);
nand UO_2967 (O_2967,N_48543,N_48582);
nor UO_2968 (O_2968,N_45490,N_48900);
nand UO_2969 (O_2969,N_47524,N_45615);
xnor UO_2970 (O_2970,N_45185,N_49284);
xnor UO_2971 (O_2971,N_45736,N_48747);
and UO_2972 (O_2972,N_46210,N_46397);
xor UO_2973 (O_2973,N_45266,N_47762);
xnor UO_2974 (O_2974,N_46727,N_45369);
nor UO_2975 (O_2975,N_49624,N_46131);
nor UO_2976 (O_2976,N_46672,N_49048);
xor UO_2977 (O_2977,N_45401,N_46522);
xnor UO_2978 (O_2978,N_46992,N_46595);
nor UO_2979 (O_2979,N_49475,N_47304);
xor UO_2980 (O_2980,N_46649,N_49672);
and UO_2981 (O_2981,N_49429,N_49853);
and UO_2982 (O_2982,N_48268,N_47219);
nor UO_2983 (O_2983,N_48322,N_47656);
xnor UO_2984 (O_2984,N_45935,N_45722);
xnor UO_2985 (O_2985,N_46164,N_45516);
or UO_2986 (O_2986,N_46404,N_49703);
nand UO_2987 (O_2987,N_45252,N_48296);
nand UO_2988 (O_2988,N_49252,N_45052);
or UO_2989 (O_2989,N_47059,N_48190);
nand UO_2990 (O_2990,N_49645,N_48828);
nand UO_2991 (O_2991,N_49975,N_49083);
nand UO_2992 (O_2992,N_46903,N_47449);
nor UO_2993 (O_2993,N_48729,N_46071);
nand UO_2994 (O_2994,N_47755,N_49215);
and UO_2995 (O_2995,N_45193,N_49429);
xor UO_2996 (O_2996,N_49092,N_45712);
or UO_2997 (O_2997,N_47973,N_46861);
xor UO_2998 (O_2998,N_48741,N_48701);
nor UO_2999 (O_2999,N_48832,N_45072);
or UO_3000 (O_3000,N_45516,N_49458);
xnor UO_3001 (O_3001,N_46438,N_46552);
xnor UO_3002 (O_3002,N_46777,N_48047);
and UO_3003 (O_3003,N_45498,N_46315);
or UO_3004 (O_3004,N_47903,N_48941);
and UO_3005 (O_3005,N_47867,N_45544);
or UO_3006 (O_3006,N_48761,N_49103);
nor UO_3007 (O_3007,N_45642,N_48562);
xor UO_3008 (O_3008,N_49994,N_47310);
xnor UO_3009 (O_3009,N_45620,N_48209);
xnor UO_3010 (O_3010,N_48247,N_48794);
nand UO_3011 (O_3011,N_45824,N_47406);
or UO_3012 (O_3012,N_47223,N_46836);
or UO_3013 (O_3013,N_47274,N_48217);
xor UO_3014 (O_3014,N_46728,N_48382);
or UO_3015 (O_3015,N_47814,N_49417);
or UO_3016 (O_3016,N_45774,N_45103);
xor UO_3017 (O_3017,N_49766,N_46900);
xnor UO_3018 (O_3018,N_49681,N_48485);
and UO_3019 (O_3019,N_45283,N_45144);
and UO_3020 (O_3020,N_46994,N_49206);
nor UO_3021 (O_3021,N_49536,N_45147);
or UO_3022 (O_3022,N_46683,N_46007);
nor UO_3023 (O_3023,N_46803,N_47631);
nor UO_3024 (O_3024,N_49447,N_45342);
nor UO_3025 (O_3025,N_45909,N_49715);
or UO_3026 (O_3026,N_47010,N_48338);
and UO_3027 (O_3027,N_49348,N_48962);
xnor UO_3028 (O_3028,N_47097,N_48769);
xnor UO_3029 (O_3029,N_45307,N_46535);
xor UO_3030 (O_3030,N_49039,N_48981);
xor UO_3031 (O_3031,N_46775,N_45166);
nand UO_3032 (O_3032,N_46649,N_46995);
xnor UO_3033 (O_3033,N_49429,N_47473);
or UO_3034 (O_3034,N_47817,N_49777);
nor UO_3035 (O_3035,N_49234,N_49615);
nand UO_3036 (O_3036,N_46744,N_49430);
xor UO_3037 (O_3037,N_48891,N_49468);
nand UO_3038 (O_3038,N_47848,N_48561);
and UO_3039 (O_3039,N_47385,N_49043);
and UO_3040 (O_3040,N_46508,N_49130);
nor UO_3041 (O_3041,N_48103,N_49409);
and UO_3042 (O_3042,N_46865,N_45014);
and UO_3043 (O_3043,N_45312,N_48097);
or UO_3044 (O_3044,N_46823,N_49817);
nand UO_3045 (O_3045,N_48996,N_46609);
and UO_3046 (O_3046,N_48142,N_49574);
nor UO_3047 (O_3047,N_47059,N_49751);
nand UO_3048 (O_3048,N_45958,N_45240);
nand UO_3049 (O_3049,N_49964,N_49232);
nor UO_3050 (O_3050,N_45421,N_45334);
nor UO_3051 (O_3051,N_47509,N_45164);
and UO_3052 (O_3052,N_45678,N_46821);
and UO_3053 (O_3053,N_48731,N_45456);
and UO_3054 (O_3054,N_46523,N_47996);
nor UO_3055 (O_3055,N_45754,N_49035);
nand UO_3056 (O_3056,N_49151,N_47835);
or UO_3057 (O_3057,N_45295,N_45774);
and UO_3058 (O_3058,N_48815,N_46064);
or UO_3059 (O_3059,N_49453,N_46057);
and UO_3060 (O_3060,N_49379,N_48195);
nor UO_3061 (O_3061,N_49719,N_47813);
xnor UO_3062 (O_3062,N_45009,N_46882);
or UO_3063 (O_3063,N_46326,N_49812);
xor UO_3064 (O_3064,N_48907,N_46501);
xor UO_3065 (O_3065,N_48973,N_46379);
or UO_3066 (O_3066,N_46433,N_46990);
or UO_3067 (O_3067,N_45042,N_49918);
xor UO_3068 (O_3068,N_47447,N_47244);
nand UO_3069 (O_3069,N_47274,N_48018);
nand UO_3070 (O_3070,N_45598,N_47856);
or UO_3071 (O_3071,N_49108,N_49163);
and UO_3072 (O_3072,N_47981,N_49506);
and UO_3073 (O_3073,N_46779,N_47872);
nand UO_3074 (O_3074,N_46499,N_49060);
or UO_3075 (O_3075,N_49950,N_49177);
xnor UO_3076 (O_3076,N_46916,N_48854);
nor UO_3077 (O_3077,N_46732,N_49810);
and UO_3078 (O_3078,N_49481,N_45279);
xor UO_3079 (O_3079,N_49253,N_45341);
nor UO_3080 (O_3080,N_49512,N_49788);
nand UO_3081 (O_3081,N_48839,N_46650);
xor UO_3082 (O_3082,N_48180,N_48691);
xnor UO_3083 (O_3083,N_45691,N_49656);
nor UO_3084 (O_3084,N_49409,N_47394);
xor UO_3085 (O_3085,N_48125,N_45163);
nor UO_3086 (O_3086,N_48664,N_47988);
xnor UO_3087 (O_3087,N_46267,N_46701);
nor UO_3088 (O_3088,N_48521,N_48669);
nor UO_3089 (O_3089,N_47089,N_49253);
and UO_3090 (O_3090,N_49706,N_48887);
and UO_3091 (O_3091,N_46710,N_46428);
or UO_3092 (O_3092,N_47636,N_49613);
or UO_3093 (O_3093,N_46217,N_47192);
nor UO_3094 (O_3094,N_45259,N_46285);
or UO_3095 (O_3095,N_47527,N_46305);
xor UO_3096 (O_3096,N_47775,N_49466);
nor UO_3097 (O_3097,N_46121,N_47891);
nand UO_3098 (O_3098,N_47356,N_46525);
xnor UO_3099 (O_3099,N_48144,N_47935);
and UO_3100 (O_3100,N_47395,N_46172);
or UO_3101 (O_3101,N_47198,N_47576);
nor UO_3102 (O_3102,N_49748,N_48309);
xnor UO_3103 (O_3103,N_48305,N_45256);
nand UO_3104 (O_3104,N_48936,N_48804);
xnor UO_3105 (O_3105,N_46215,N_46984);
nor UO_3106 (O_3106,N_48725,N_48348);
xnor UO_3107 (O_3107,N_49177,N_47548);
and UO_3108 (O_3108,N_45893,N_47604);
nor UO_3109 (O_3109,N_49103,N_49617);
nor UO_3110 (O_3110,N_47999,N_48370);
or UO_3111 (O_3111,N_48686,N_45913);
xnor UO_3112 (O_3112,N_46041,N_49319);
and UO_3113 (O_3113,N_49051,N_46334);
xnor UO_3114 (O_3114,N_47919,N_47687);
xor UO_3115 (O_3115,N_47612,N_46965);
or UO_3116 (O_3116,N_48366,N_47444);
nor UO_3117 (O_3117,N_49301,N_49734);
nor UO_3118 (O_3118,N_49219,N_47598);
or UO_3119 (O_3119,N_48597,N_49247);
or UO_3120 (O_3120,N_46048,N_46775);
or UO_3121 (O_3121,N_48510,N_47902);
and UO_3122 (O_3122,N_47955,N_46941);
nor UO_3123 (O_3123,N_49725,N_49780);
nand UO_3124 (O_3124,N_46540,N_46949);
nand UO_3125 (O_3125,N_48971,N_46033);
nand UO_3126 (O_3126,N_49340,N_46410);
or UO_3127 (O_3127,N_49802,N_47993);
nand UO_3128 (O_3128,N_45028,N_46069);
nor UO_3129 (O_3129,N_47650,N_45411);
or UO_3130 (O_3130,N_45909,N_46647);
nand UO_3131 (O_3131,N_46587,N_48771);
or UO_3132 (O_3132,N_47737,N_45144);
and UO_3133 (O_3133,N_48827,N_47839);
or UO_3134 (O_3134,N_48316,N_47913);
or UO_3135 (O_3135,N_46790,N_47588);
or UO_3136 (O_3136,N_47622,N_45172);
and UO_3137 (O_3137,N_46650,N_49641);
nor UO_3138 (O_3138,N_47836,N_49575);
xnor UO_3139 (O_3139,N_49304,N_47072);
nor UO_3140 (O_3140,N_48004,N_46996);
and UO_3141 (O_3141,N_46080,N_47182);
nand UO_3142 (O_3142,N_49739,N_46507);
xor UO_3143 (O_3143,N_46487,N_48516);
and UO_3144 (O_3144,N_47955,N_47927);
nand UO_3145 (O_3145,N_47142,N_45158);
xnor UO_3146 (O_3146,N_47309,N_45481);
nor UO_3147 (O_3147,N_49745,N_49900);
and UO_3148 (O_3148,N_49973,N_48993);
or UO_3149 (O_3149,N_48910,N_45573);
nand UO_3150 (O_3150,N_46742,N_49861);
and UO_3151 (O_3151,N_48209,N_49822);
or UO_3152 (O_3152,N_49386,N_45098);
xor UO_3153 (O_3153,N_45545,N_46031);
and UO_3154 (O_3154,N_47441,N_45937);
or UO_3155 (O_3155,N_45765,N_46775);
xnor UO_3156 (O_3156,N_47735,N_47730);
and UO_3157 (O_3157,N_49354,N_49867);
nand UO_3158 (O_3158,N_47666,N_48208);
and UO_3159 (O_3159,N_45321,N_47902);
and UO_3160 (O_3160,N_49562,N_45479);
or UO_3161 (O_3161,N_45031,N_45183);
or UO_3162 (O_3162,N_47988,N_45209);
and UO_3163 (O_3163,N_49194,N_47942);
nor UO_3164 (O_3164,N_47378,N_46458);
and UO_3165 (O_3165,N_47321,N_45847);
and UO_3166 (O_3166,N_45316,N_45394);
or UO_3167 (O_3167,N_46666,N_46611);
nand UO_3168 (O_3168,N_46956,N_47447);
nor UO_3169 (O_3169,N_49366,N_49454);
and UO_3170 (O_3170,N_48864,N_49335);
nand UO_3171 (O_3171,N_48201,N_46327);
and UO_3172 (O_3172,N_47967,N_45106);
or UO_3173 (O_3173,N_48693,N_48816);
xnor UO_3174 (O_3174,N_45493,N_45654);
or UO_3175 (O_3175,N_47228,N_45863);
nor UO_3176 (O_3176,N_48988,N_49711);
nand UO_3177 (O_3177,N_46844,N_46994);
or UO_3178 (O_3178,N_46862,N_47897);
xor UO_3179 (O_3179,N_49084,N_45234);
xnor UO_3180 (O_3180,N_48198,N_48155);
nor UO_3181 (O_3181,N_49865,N_46678);
nand UO_3182 (O_3182,N_48923,N_45960);
nor UO_3183 (O_3183,N_45401,N_48746);
nand UO_3184 (O_3184,N_48708,N_48939);
or UO_3185 (O_3185,N_48123,N_49335);
xor UO_3186 (O_3186,N_45099,N_49714);
xnor UO_3187 (O_3187,N_49063,N_45723);
nand UO_3188 (O_3188,N_49700,N_46290);
xnor UO_3189 (O_3189,N_47937,N_48175);
nand UO_3190 (O_3190,N_48218,N_46181);
nor UO_3191 (O_3191,N_46525,N_46649);
xor UO_3192 (O_3192,N_48775,N_47538);
nand UO_3193 (O_3193,N_45527,N_48317);
and UO_3194 (O_3194,N_47030,N_49424);
or UO_3195 (O_3195,N_48926,N_46260);
and UO_3196 (O_3196,N_47292,N_45827);
xor UO_3197 (O_3197,N_46753,N_49516);
nand UO_3198 (O_3198,N_49432,N_48548);
nand UO_3199 (O_3199,N_47720,N_46048);
nor UO_3200 (O_3200,N_48524,N_48860);
and UO_3201 (O_3201,N_46275,N_48845);
or UO_3202 (O_3202,N_47928,N_47911);
or UO_3203 (O_3203,N_46319,N_47866);
nor UO_3204 (O_3204,N_48735,N_46296);
or UO_3205 (O_3205,N_49217,N_48901);
nor UO_3206 (O_3206,N_45695,N_48153);
nand UO_3207 (O_3207,N_45674,N_48237);
nand UO_3208 (O_3208,N_49844,N_47443);
nand UO_3209 (O_3209,N_48079,N_49580);
or UO_3210 (O_3210,N_45029,N_49792);
and UO_3211 (O_3211,N_48770,N_49999);
nor UO_3212 (O_3212,N_48806,N_49379);
or UO_3213 (O_3213,N_49800,N_47863);
and UO_3214 (O_3214,N_47349,N_49271);
nor UO_3215 (O_3215,N_47159,N_49363);
nor UO_3216 (O_3216,N_49472,N_46477);
or UO_3217 (O_3217,N_49607,N_48934);
nor UO_3218 (O_3218,N_45034,N_48342);
nand UO_3219 (O_3219,N_47545,N_49700);
or UO_3220 (O_3220,N_49253,N_46206);
and UO_3221 (O_3221,N_45232,N_48474);
nand UO_3222 (O_3222,N_47256,N_47167);
nand UO_3223 (O_3223,N_46155,N_47298);
xor UO_3224 (O_3224,N_49105,N_49274);
nor UO_3225 (O_3225,N_48044,N_48342);
nand UO_3226 (O_3226,N_48947,N_47719);
nor UO_3227 (O_3227,N_48480,N_45755);
nand UO_3228 (O_3228,N_46575,N_48224);
nand UO_3229 (O_3229,N_48866,N_48864);
xnor UO_3230 (O_3230,N_47141,N_48345);
nor UO_3231 (O_3231,N_45561,N_47082);
nor UO_3232 (O_3232,N_47171,N_48677);
or UO_3233 (O_3233,N_46809,N_47711);
nand UO_3234 (O_3234,N_47726,N_46672);
or UO_3235 (O_3235,N_45316,N_46285);
nand UO_3236 (O_3236,N_48642,N_45494);
and UO_3237 (O_3237,N_49303,N_45456);
or UO_3238 (O_3238,N_47945,N_49116);
nor UO_3239 (O_3239,N_49515,N_46600);
nand UO_3240 (O_3240,N_47663,N_46629);
nor UO_3241 (O_3241,N_48142,N_49458);
nand UO_3242 (O_3242,N_45010,N_48234);
nand UO_3243 (O_3243,N_49934,N_46926);
and UO_3244 (O_3244,N_48494,N_45964);
xor UO_3245 (O_3245,N_49124,N_45561);
nor UO_3246 (O_3246,N_46671,N_48995);
nand UO_3247 (O_3247,N_48536,N_47919);
and UO_3248 (O_3248,N_48281,N_48238);
nand UO_3249 (O_3249,N_46954,N_48220);
or UO_3250 (O_3250,N_49049,N_49998);
nand UO_3251 (O_3251,N_49030,N_48792);
nand UO_3252 (O_3252,N_45723,N_49609);
nand UO_3253 (O_3253,N_49030,N_45303);
nor UO_3254 (O_3254,N_48627,N_47137);
or UO_3255 (O_3255,N_46513,N_46163);
nand UO_3256 (O_3256,N_46141,N_48466);
xnor UO_3257 (O_3257,N_47214,N_48232);
nor UO_3258 (O_3258,N_45637,N_48784);
nand UO_3259 (O_3259,N_45195,N_46160);
nand UO_3260 (O_3260,N_49293,N_45365);
xor UO_3261 (O_3261,N_47644,N_45565);
xnor UO_3262 (O_3262,N_48002,N_48758);
nand UO_3263 (O_3263,N_47106,N_46829);
nand UO_3264 (O_3264,N_49885,N_46960);
nand UO_3265 (O_3265,N_45141,N_47212);
or UO_3266 (O_3266,N_49618,N_49346);
nand UO_3267 (O_3267,N_45347,N_48784);
or UO_3268 (O_3268,N_49263,N_45312);
xor UO_3269 (O_3269,N_47005,N_49429);
xnor UO_3270 (O_3270,N_49050,N_46404);
nand UO_3271 (O_3271,N_47922,N_47294);
nand UO_3272 (O_3272,N_49074,N_49210);
or UO_3273 (O_3273,N_47560,N_49920);
and UO_3274 (O_3274,N_47831,N_45448);
xor UO_3275 (O_3275,N_45366,N_49792);
or UO_3276 (O_3276,N_49362,N_45362);
or UO_3277 (O_3277,N_49933,N_48659);
or UO_3278 (O_3278,N_45546,N_47566);
and UO_3279 (O_3279,N_46466,N_46406);
and UO_3280 (O_3280,N_47109,N_48726);
nand UO_3281 (O_3281,N_49227,N_45787);
xor UO_3282 (O_3282,N_45585,N_47143);
and UO_3283 (O_3283,N_45503,N_46757);
nor UO_3284 (O_3284,N_47559,N_45585);
nand UO_3285 (O_3285,N_45228,N_45762);
nor UO_3286 (O_3286,N_47105,N_46710);
or UO_3287 (O_3287,N_47759,N_45948);
nand UO_3288 (O_3288,N_49235,N_45121);
xnor UO_3289 (O_3289,N_48484,N_48950);
nor UO_3290 (O_3290,N_48726,N_47415);
or UO_3291 (O_3291,N_49953,N_47010);
and UO_3292 (O_3292,N_49810,N_49498);
xor UO_3293 (O_3293,N_45843,N_49321);
nand UO_3294 (O_3294,N_46904,N_49068);
nand UO_3295 (O_3295,N_49238,N_48036);
xor UO_3296 (O_3296,N_49570,N_46687);
xor UO_3297 (O_3297,N_47285,N_47022);
and UO_3298 (O_3298,N_46621,N_46860);
xor UO_3299 (O_3299,N_45963,N_49292);
nor UO_3300 (O_3300,N_46489,N_49607);
and UO_3301 (O_3301,N_45325,N_47669);
nor UO_3302 (O_3302,N_48882,N_49031);
and UO_3303 (O_3303,N_46780,N_48914);
nand UO_3304 (O_3304,N_47339,N_46342);
or UO_3305 (O_3305,N_47028,N_49947);
nand UO_3306 (O_3306,N_45448,N_46245);
xnor UO_3307 (O_3307,N_49178,N_46271);
and UO_3308 (O_3308,N_46398,N_46406);
or UO_3309 (O_3309,N_45260,N_47946);
xnor UO_3310 (O_3310,N_48001,N_46868);
or UO_3311 (O_3311,N_48100,N_48815);
or UO_3312 (O_3312,N_48137,N_49721);
or UO_3313 (O_3313,N_48409,N_46254);
nor UO_3314 (O_3314,N_46246,N_47561);
or UO_3315 (O_3315,N_46805,N_49588);
and UO_3316 (O_3316,N_48539,N_49334);
xor UO_3317 (O_3317,N_47356,N_47667);
nand UO_3318 (O_3318,N_46859,N_47248);
nor UO_3319 (O_3319,N_48881,N_45298);
or UO_3320 (O_3320,N_45543,N_46237);
or UO_3321 (O_3321,N_46019,N_47033);
nand UO_3322 (O_3322,N_48835,N_49171);
or UO_3323 (O_3323,N_46689,N_46922);
nor UO_3324 (O_3324,N_49661,N_49548);
xnor UO_3325 (O_3325,N_47616,N_45762);
nor UO_3326 (O_3326,N_46227,N_48024);
nor UO_3327 (O_3327,N_45937,N_49633);
and UO_3328 (O_3328,N_48978,N_46689);
xnor UO_3329 (O_3329,N_45207,N_45451);
xor UO_3330 (O_3330,N_46908,N_46031);
nand UO_3331 (O_3331,N_48648,N_45183);
and UO_3332 (O_3332,N_48406,N_49451);
and UO_3333 (O_3333,N_49855,N_49382);
nor UO_3334 (O_3334,N_46896,N_46539);
nand UO_3335 (O_3335,N_46593,N_47829);
nand UO_3336 (O_3336,N_48770,N_47768);
and UO_3337 (O_3337,N_47536,N_46404);
or UO_3338 (O_3338,N_45600,N_45001);
xnor UO_3339 (O_3339,N_47081,N_46178);
nand UO_3340 (O_3340,N_45039,N_48221);
and UO_3341 (O_3341,N_45285,N_49949);
nand UO_3342 (O_3342,N_47326,N_45031);
and UO_3343 (O_3343,N_48755,N_46414);
nand UO_3344 (O_3344,N_49412,N_46501);
xnor UO_3345 (O_3345,N_47868,N_47576);
and UO_3346 (O_3346,N_48985,N_46884);
nand UO_3347 (O_3347,N_45183,N_47999);
xnor UO_3348 (O_3348,N_48082,N_47304);
xnor UO_3349 (O_3349,N_45644,N_48492);
or UO_3350 (O_3350,N_47654,N_46322);
nand UO_3351 (O_3351,N_47582,N_46616);
xor UO_3352 (O_3352,N_49633,N_46806);
xor UO_3353 (O_3353,N_49724,N_46538);
xor UO_3354 (O_3354,N_49309,N_47007);
and UO_3355 (O_3355,N_47234,N_47241);
nand UO_3356 (O_3356,N_49710,N_45760);
xor UO_3357 (O_3357,N_49737,N_45007);
or UO_3358 (O_3358,N_48427,N_49309);
nor UO_3359 (O_3359,N_48576,N_47644);
nand UO_3360 (O_3360,N_49024,N_46837);
or UO_3361 (O_3361,N_49061,N_49528);
xor UO_3362 (O_3362,N_45880,N_48583);
and UO_3363 (O_3363,N_48027,N_48077);
nand UO_3364 (O_3364,N_49515,N_47672);
and UO_3365 (O_3365,N_49149,N_48897);
nor UO_3366 (O_3366,N_46999,N_49018);
or UO_3367 (O_3367,N_45712,N_47822);
nand UO_3368 (O_3368,N_48911,N_45095);
or UO_3369 (O_3369,N_49807,N_45614);
or UO_3370 (O_3370,N_48684,N_49756);
and UO_3371 (O_3371,N_49727,N_48560);
xnor UO_3372 (O_3372,N_47613,N_46737);
xnor UO_3373 (O_3373,N_48227,N_45393);
nand UO_3374 (O_3374,N_48870,N_49339);
xor UO_3375 (O_3375,N_49390,N_49317);
or UO_3376 (O_3376,N_49078,N_46113);
or UO_3377 (O_3377,N_46218,N_47577);
nor UO_3378 (O_3378,N_48263,N_48094);
nand UO_3379 (O_3379,N_49794,N_45958);
xnor UO_3380 (O_3380,N_45464,N_47584);
and UO_3381 (O_3381,N_46278,N_47422);
or UO_3382 (O_3382,N_47645,N_47586);
and UO_3383 (O_3383,N_46190,N_48441);
nand UO_3384 (O_3384,N_45026,N_46190);
and UO_3385 (O_3385,N_45055,N_45185);
nor UO_3386 (O_3386,N_49784,N_46803);
or UO_3387 (O_3387,N_47489,N_49091);
and UO_3388 (O_3388,N_46496,N_46651);
nand UO_3389 (O_3389,N_47402,N_49275);
nor UO_3390 (O_3390,N_47870,N_48105);
nand UO_3391 (O_3391,N_46173,N_46298);
and UO_3392 (O_3392,N_49292,N_45622);
nand UO_3393 (O_3393,N_46591,N_46062);
xnor UO_3394 (O_3394,N_47403,N_46886);
xor UO_3395 (O_3395,N_46145,N_45345);
xnor UO_3396 (O_3396,N_45547,N_47193);
xor UO_3397 (O_3397,N_47945,N_49205);
or UO_3398 (O_3398,N_47346,N_45728);
xor UO_3399 (O_3399,N_49926,N_45558);
or UO_3400 (O_3400,N_46561,N_47438);
and UO_3401 (O_3401,N_47233,N_47597);
or UO_3402 (O_3402,N_49386,N_46552);
or UO_3403 (O_3403,N_48901,N_48010);
nor UO_3404 (O_3404,N_47292,N_49605);
nor UO_3405 (O_3405,N_46255,N_45590);
nand UO_3406 (O_3406,N_49186,N_46362);
nor UO_3407 (O_3407,N_48676,N_49652);
or UO_3408 (O_3408,N_49118,N_47097);
xnor UO_3409 (O_3409,N_48957,N_48344);
or UO_3410 (O_3410,N_49080,N_46586);
or UO_3411 (O_3411,N_49867,N_46463);
xor UO_3412 (O_3412,N_49694,N_45488);
xor UO_3413 (O_3413,N_48037,N_45957);
nor UO_3414 (O_3414,N_48260,N_46811);
or UO_3415 (O_3415,N_45668,N_49131);
xor UO_3416 (O_3416,N_49925,N_48434);
xor UO_3417 (O_3417,N_45785,N_48943);
xnor UO_3418 (O_3418,N_48029,N_49295);
nor UO_3419 (O_3419,N_49931,N_48751);
nand UO_3420 (O_3420,N_47752,N_49966);
nand UO_3421 (O_3421,N_46914,N_48023);
and UO_3422 (O_3422,N_45639,N_45118);
nor UO_3423 (O_3423,N_48443,N_49702);
or UO_3424 (O_3424,N_49469,N_46885);
nand UO_3425 (O_3425,N_45548,N_47126);
nor UO_3426 (O_3426,N_47194,N_49189);
and UO_3427 (O_3427,N_49637,N_47691);
nand UO_3428 (O_3428,N_48578,N_45807);
or UO_3429 (O_3429,N_47934,N_46581);
nand UO_3430 (O_3430,N_45176,N_48213);
or UO_3431 (O_3431,N_46563,N_46896);
nor UO_3432 (O_3432,N_48722,N_46927);
xor UO_3433 (O_3433,N_47519,N_46092);
and UO_3434 (O_3434,N_45190,N_48552);
or UO_3435 (O_3435,N_47476,N_49745);
xor UO_3436 (O_3436,N_47801,N_48186);
nand UO_3437 (O_3437,N_46287,N_48246);
and UO_3438 (O_3438,N_47235,N_46420);
nand UO_3439 (O_3439,N_46217,N_46195);
nand UO_3440 (O_3440,N_47589,N_49704);
and UO_3441 (O_3441,N_46827,N_48246);
xor UO_3442 (O_3442,N_47028,N_46249);
or UO_3443 (O_3443,N_48422,N_46083);
nand UO_3444 (O_3444,N_47559,N_46461);
or UO_3445 (O_3445,N_47904,N_46306);
nand UO_3446 (O_3446,N_47353,N_46997);
or UO_3447 (O_3447,N_48278,N_48479);
nand UO_3448 (O_3448,N_47265,N_46202);
xor UO_3449 (O_3449,N_47341,N_49091);
and UO_3450 (O_3450,N_49162,N_49464);
or UO_3451 (O_3451,N_45107,N_47594);
nor UO_3452 (O_3452,N_49848,N_48060);
and UO_3453 (O_3453,N_49248,N_49422);
nand UO_3454 (O_3454,N_46375,N_48760);
xnor UO_3455 (O_3455,N_48043,N_46768);
nand UO_3456 (O_3456,N_48094,N_47323);
and UO_3457 (O_3457,N_47153,N_45668);
nor UO_3458 (O_3458,N_45103,N_49469);
nor UO_3459 (O_3459,N_48343,N_45559);
nor UO_3460 (O_3460,N_46666,N_46079);
xor UO_3461 (O_3461,N_49155,N_46105);
or UO_3462 (O_3462,N_45005,N_47908);
and UO_3463 (O_3463,N_49936,N_47917);
nand UO_3464 (O_3464,N_49698,N_48464);
and UO_3465 (O_3465,N_47269,N_49029);
and UO_3466 (O_3466,N_47634,N_47867);
nand UO_3467 (O_3467,N_45045,N_46557);
or UO_3468 (O_3468,N_49088,N_45800);
nand UO_3469 (O_3469,N_45406,N_49942);
nor UO_3470 (O_3470,N_47605,N_45017);
xnor UO_3471 (O_3471,N_45193,N_48423);
and UO_3472 (O_3472,N_48483,N_48500);
nand UO_3473 (O_3473,N_49819,N_46011);
xor UO_3474 (O_3474,N_49551,N_45079);
nor UO_3475 (O_3475,N_45574,N_46535);
xnor UO_3476 (O_3476,N_45293,N_47969);
nor UO_3477 (O_3477,N_47659,N_45565);
nand UO_3478 (O_3478,N_48949,N_49628);
and UO_3479 (O_3479,N_49062,N_45730);
nand UO_3480 (O_3480,N_48381,N_47706);
nor UO_3481 (O_3481,N_47136,N_49001);
xor UO_3482 (O_3482,N_49998,N_46588);
or UO_3483 (O_3483,N_47215,N_47088);
nor UO_3484 (O_3484,N_47389,N_46278);
and UO_3485 (O_3485,N_49767,N_45337);
nand UO_3486 (O_3486,N_47090,N_45475);
xnor UO_3487 (O_3487,N_49213,N_46219);
xnor UO_3488 (O_3488,N_49875,N_48175);
nand UO_3489 (O_3489,N_47013,N_46728);
and UO_3490 (O_3490,N_49703,N_46668);
nor UO_3491 (O_3491,N_49360,N_48339);
nand UO_3492 (O_3492,N_45871,N_45364);
or UO_3493 (O_3493,N_45162,N_47755);
and UO_3494 (O_3494,N_46338,N_45490);
or UO_3495 (O_3495,N_49965,N_49841);
nor UO_3496 (O_3496,N_45405,N_49847);
or UO_3497 (O_3497,N_49794,N_46753);
nor UO_3498 (O_3498,N_48002,N_46475);
nand UO_3499 (O_3499,N_45096,N_49637);
and UO_3500 (O_3500,N_48523,N_45167);
and UO_3501 (O_3501,N_49934,N_47637);
or UO_3502 (O_3502,N_45171,N_46125);
and UO_3503 (O_3503,N_46854,N_47319);
or UO_3504 (O_3504,N_46845,N_49268);
or UO_3505 (O_3505,N_46350,N_46050);
nand UO_3506 (O_3506,N_48726,N_45870);
and UO_3507 (O_3507,N_45772,N_45675);
xnor UO_3508 (O_3508,N_45745,N_47457);
or UO_3509 (O_3509,N_45538,N_46527);
or UO_3510 (O_3510,N_48989,N_47348);
nor UO_3511 (O_3511,N_45151,N_46726);
and UO_3512 (O_3512,N_47104,N_48381);
or UO_3513 (O_3513,N_46537,N_49690);
and UO_3514 (O_3514,N_49352,N_45532);
xnor UO_3515 (O_3515,N_47089,N_46648);
nor UO_3516 (O_3516,N_48145,N_45196);
and UO_3517 (O_3517,N_47080,N_45500);
xnor UO_3518 (O_3518,N_49116,N_46673);
or UO_3519 (O_3519,N_47050,N_48112);
xor UO_3520 (O_3520,N_45359,N_49328);
nor UO_3521 (O_3521,N_47683,N_45983);
xor UO_3522 (O_3522,N_47297,N_46995);
or UO_3523 (O_3523,N_45294,N_49375);
nand UO_3524 (O_3524,N_46590,N_45460);
or UO_3525 (O_3525,N_48030,N_47077);
nor UO_3526 (O_3526,N_45984,N_47467);
xor UO_3527 (O_3527,N_49722,N_46775);
nor UO_3528 (O_3528,N_49887,N_49397);
xnor UO_3529 (O_3529,N_49269,N_46012);
nor UO_3530 (O_3530,N_49731,N_46963);
and UO_3531 (O_3531,N_48586,N_49967);
and UO_3532 (O_3532,N_49145,N_49689);
nor UO_3533 (O_3533,N_47136,N_49906);
or UO_3534 (O_3534,N_46547,N_47491);
xnor UO_3535 (O_3535,N_49717,N_45105);
or UO_3536 (O_3536,N_48628,N_46941);
xor UO_3537 (O_3537,N_46111,N_48181);
nand UO_3538 (O_3538,N_49492,N_48486);
nand UO_3539 (O_3539,N_48331,N_45043);
or UO_3540 (O_3540,N_49064,N_48312);
xor UO_3541 (O_3541,N_47073,N_47263);
nor UO_3542 (O_3542,N_47524,N_47488);
xor UO_3543 (O_3543,N_45612,N_48434);
nand UO_3544 (O_3544,N_46069,N_48104);
and UO_3545 (O_3545,N_46310,N_48080);
nand UO_3546 (O_3546,N_47249,N_45156);
nor UO_3547 (O_3547,N_45723,N_48344);
nand UO_3548 (O_3548,N_47398,N_49811);
and UO_3549 (O_3549,N_45550,N_45755);
or UO_3550 (O_3550,N_48959,N_49391);
or UO_3551 (O_3551,N_46153,N_45951);
and UO_3552 (O_3552,N_48880,N_46142);
or UO_3553 (O_3553,N_47435,N_45891);
nor UO_3554 (O_3554,N_48273,N_46116);
or UO_3555 (O_3555,N_45764,N_46449);
and UO_3556 (O_3556,N_46558,N_47926);
or UO_3557 (O_3557,N_48146,N_48869);
and UO_3558 (O_3558,N_47397,N_46489);
nor UO_3559 (O_3559,N_45947,N_45911);
nand UO_3560 (O_3560,N_45971,N_49433);
or UO_3561 (O_3561,N_47979,N_48803);
nand UO_3562 (O_3562,N_45155,N_49795);
and UO_3563 (O_3563,N_48282,N_47499);
or UO_3564 (O_3564,N_49293,N_48987);
or UO_3565 (O_3565,N_45365,N_46026);
or UO_3566 (O_3566,N_46378,N_49820);
and UO_3567 (O_3567,N_46069,N_49339);
or UO_3568 (O_3568,N_46763,N_46495);
and UO_3569 (O_3569,N_48498,N_45248);
nand UO_3570 (O_3570,N_49509,N_47845);
xnor UO_3571 (O_3571,N_47060,N_47812);
and UO_3572 (O_3572,N_48551,N_49365);
nor UO_3573 (O_3573,N_46918,N_49251);
and UO_3574 (O_3574,N_48573,N_45891);
or UO_3575 (O_3575,N_46025,N_48237);
nand UO_3576 (O_3576,N_48259,N_47451);
nor UO_3577 (O_3577,N_47003,N_47997);
or UO_3578 (O_3578,N_47686,N_46104);
nand UO_3579 (O_3579,N_49231,N_45888);
or UO_3580 (O_3580,N_46896,N_47371);
xnor UO_3581 (O_3581,N_48125,N_49163);
nand UO_3582 (O_3582,N_48644,N_48902);
or UO_3583 (O_3583,N_47281,N_46279);
or UO_3584 (O_3584,N_46350,N_46726);
and UO_3585 (O_3585,N_45049,N_49651);
nor UO_3586 (O_3586,N_47183,N_47794);
xnor UO_3587 (O_3587,N_45453,N_48583);
and UO_3588 (O_3588,N_46334,N_47514);
xnor UO_3589 (O_3589,N_49185,N_47138);
and UO_3590 (O_3590,N_47161,N_46499);
or UO_3591 (O_3591,N_46918,N_46364);
nand UO_3592 (O_3592,N_47414,N_46847);
nor UO_3593 (O_3593,N_48105,N_49705);
and UO_3594 (O_3594,N_46872,N_48325);
or UO_3595 (O_3595,N_49002,N_47969);
and UO_3596 (O_3596,N_45150,N_49926);
and UO_3597 (O_3597,N_47873,N_47088);
or UO_3598 (O_3598,N_48498,N_48365);
nand UO_3599 (O_3599,N_49769,N_46395);
nand UO_3600 (O_3600,N_48691,N_48553);
xnor UO_3601 (O_3601,N_48402,N_46360);
or UO_3602 (O_3602,N_45347,N_47777);
or UO_3603 (O_3603,N_48058,N_47041);
and UO_3604 (O_3604,N_48634,N_46907);
nand UO_3605 (O_3605,N_46507,N_46588);
xor UO_3606 (O_3606,N_46476,N_48222);
nor UO_3607 (O_3607,N_47545,N_48896);
and UO_3608 (O_3608,N_49769,N_49597);
nor UO_3609 (O_3609,N_49582,N_46424);
nor UO_3610 (O_3610,N_45597,N_49061);
xor UO_3611 (O_3611,N_45564,N_46292);
or UO_3612 (O_3612,N_45567,N_45998);
xor UO_3613 (O_3613,N_47140,N_49173);
nor UO_3614 (O_3614,N_47609,N_46324);
nor UO_3615 (O_3615,N_45098,N_49714);
or UO_3616 (O_3616,N_49895,N_45478);
and UO_3617 (O_3617,N_45518,N_48821);
xor UO_3618 (O_3618,N_47176,N_45610);
xnor UO_3619 (O_3619,N_46727,N_46219);
xnor UO_3620 (O_3620,N_45013,N_47842);
xnor UO_3621 (O_3621,N_48298,N_47441);
nand UO_3622 (O_3622,N_49585,N_48050);
or UO_3623 (O_3623,N_49015,N_46115);
or UO_3624 (O_3624,N_49791,N_48232);
xnor UO_3625 (O_3625,N_46883,N_49795);
and UO_3626 (O_3626,N_46447,N_48261);
xnor UO_3627 (O_3627,N_46628,N_47776);
nand UO_3628 (O_3628,N_48861,N_48473);
nand UO_3629 (O_3629,N_48875,N_49245);
xor UO_3630 (O_3630,N_49832,N_46873);
and UO_3631 (O_3631,N_47486,N_46888);
nor UO_3632 (O_3632,N_46420,N_46739);
nand UO_3633 (O_3633,N_48852,N_48831);
and UO_3634 (O_3634,N_48027,N_45006);
and UO_3635 (O_3635,N_48649,N_48220);
nor UO_3636 (O_3636,N_45150,N_49234);
and UO_3637 (O_3637,N_45579,N_45169);
xor UO_3638 (O_3638,N_49659,N_49100);
xor UO_3639 (O_3639,N_49601,N_45737);
and UO_3640 (O_3640,N_46299,N_48431);
or UO_3641 (O_3641,N_48120,N_49015);
or UO_3642 (O_3642,N_45252,N_47023);
or UO_3643 (O_3643,N_46745,N_48564);
or UO_3644 (O_3644,N_46703,N_45501);
nand UO_3645 (O_3645,N_48706,N_47178);
nor UO_3646 (O_3646,N_48864,N_47124);
nor UO_3647 (O_3647,N_45890,N_48809);
or UO_3648 (O_3648,N_45780,N_48981);
xnor UO_3649 (O_3649,N_47389,N_48500);
or UO_3650 (O_3650,N_45870,N_47406);
xor UO_3651 (O_3651,N_46827,N_49702);
nor UO_3652 (O_3652,N_46077,N_45754);
xnor UO_3653 (O_3653,N_46907,N_46604);
and UO_3654 (O_3654,N_47772,N_45753);
or UO_3655 (O_3655,N_47096,N_49731);
and UO_3656 (O_3656,N_45665,N_46375);
or UO_3657 (O_3657,N_48941,N_48647);
and UO_3658 (O_3658,N_47062,N_45021);
or UO_3659 (O_3659,N_49631,N_46766);
and UO_3660 (O_3660,N_46880,N_47429);
xor UO_3661 (O_3661,N_48491,N_47086);
nand UO_3662 (O_3662,N_48427,N_47261);
or UO_3663 (O_3663,N_45189,N_48168);
xor UO_3664 (O_3664,N_49700,N_45075);
nand UO_3665 (O_3665,N_48973,N_46820);
and UO_3666 (O_3666,N_47174,N_46239);
and UO_3667 (O_3667,N_45029,N_48917);
or UO_3668 (O_3668,N_49763,N_45181);
nand UO_3669 (O_3669,N_48910,N_48949);
nor UO_3670 (O_3670,N_45903,N_47188);
nor UO_3671 (O_3671,N_49983,N_47566);
xor UO_3672 (O_3672,N_46910,N_46857);
nor UO_3673 (O_3673,N_47549,N_48378);
or UO_3674 (O_3674,N_49445,N_48446);
nand UO_3675 (O_3675,N_46248,N_46936);
nand UO_3676 (O_3676,N_48089,N_49640);
nand UO_3677 (O_3677,N_47859,N_46212);
nor UO_3678 (O_3678,N_47729,N_47118);
and UO_3679 (O_3679,N_46376,N_46189);
nand UO_3680 (O_3680,N_45045,N_45716);
or UO_3681 (O_3681,N_47803,N_46136);
or UO_3682 (O_3682,N_48474,N_45018);
xor UO_3683 (O_3683,N_45755,N_49577);
or UO_3684 (O_3684,N_49393,N_45217);
and UO_3685 (O_3685,N_47067,N_49782);
and UO_3686 (O_3686,N_47211,N_48014);
or UO_3687 (O_3687,N_45176,N_46581);
and UO_3688 (O_3688,N_48524,N_46962);
nor UO_3689 (O_3689,N_45363,N_45871);
and UO_3690 (O_3690,N_45604,N_45530);
or UO_3691 (O_3691,N_47368,N_47715);
nand UO_3692 (O_3692,N_49211,N_47598);
and UO_3693 (O_3693,N_46968,N_49523);
or UO_3694 (O_3694,N_46407,N_46655);
and UO_3695 (O_3695,N_47860,N_47859);
and UO_3696 (O_3696,N_47447,N_49006);
and UO_3697 (O_3697,N_46783,N_47168);
or UO_3698 (O_3698,N_48423,N_47671);
nor UO_3699 (O_3699,N_45906,N_48100);
nand UO_3700 (O_3700,N_46712,N_45492);
or UO_3701 (O_3701,N_45969,N_45886);
xnor UO_3702 (O_3702,N_45855,N_45628);
xor UO_3703 (O_3703,N_49689,N_46076);
or UO_3704 (O_3704,N_48893,N_47996);
and UO_3705 (O_3705,N_46432,N_49887);
or UO_3706 (O_3706,N_45377,N_46953);
xnor UO_3707 (O_3707,N_46166,N_45713);
nor UO_3708 (O_3708,N_45075,N_46206);
and UO_3709 (O_3709,N_49619,N_45876);
or UO_3710 (O_3710,N_45593,N_45632);
nor UO_3711 (O_3711,N_45114,N_45966);
nor UO_3712 (O_3712,N_46808,N_49913);
nand UO_3713 (O_3713,N_46514,N_46406);
nor UO_3714 (O_3714,N_49109,N_47426);
and UO_3715 (O_3715,N_48693,N_46608);
xnor UO_3716 (O_3716,N_45908,N_46694);
and UO_3717 (O_3717,N_47461,N_49157);
xor UO_3718 (O_3718,N_48082,N_47467);
xor UO_3719 (O_3719,N_48966,N_47908);
or UO_3720 (O_3720,N_47271,N_47241);
nor UO_3721 (O_3721,N_45219,N_49223);
nand UO_3722 (O_3722,N_45839,N_46812);
or UO_3723 (O_3723,N_48808,N_45983);
nor UO_3724 (O_3724,N_47502,N_49605);
and UO_3725 (O_3725,N_46218,N_48839);
nor UO_3726 (O_3726,N_45644,N_49280);
nand UO_3727 (O_3727,N_48845,N_49590);
nor UO_3728 (O_3728,N_45470,N_46309);
nor UO_3729 (O_3729,N_48455,N_45820);
nor UO_3730 (O_3730,N_49039,N_45881);
nand UO_3731 (O_3731,N_45824,N_48853);
and UO_3732 (O_3732,N_45658,N_45672);
nand UO_3733 (O_3733,N_47393,N_48326);
nor UO_3734 (O_3734,N_45800,N_48462);
and UO_3735 (O_3735,N_46932,N_47748);
nand UO_3736 (O_3736,N_46893,N_49933);
nor UO_3737 (O_3737,N_46613,N_47378);
or UO_3738 (O_3738,N_49570,N_49813);
or UO_3739 (O_3739,N_48203,N_49771);
nand UO_3740 (O_3740,N_45913,N_46868);
or UO_3741 (O_3741,N_46691,N_45648);
or UO_3742 (O_3742,N_49736,N_46950);
xor UO_3743 (O_3743,N_45608,N_48582);
or UO_3744 (O_3744,N_48319,N_47432);
or UO_3745 (O_3745,N_48759,N_46840);
xnor UO_3746 (O_3746,N_48185,N_47251);
xnor UO_3747 (O_3747,N_47867,N_49975);
nor UO_3748 (O_3748,N_48182,N_47416);
and UO_3749 (O_3749,N_48999,N_45627);
nor UO_3750 (O_3750,N_47478,N_49235);
and UO_3751 (O_3751,N_45442,N_45172);
or UO_3752 (O_3752,N_49009,N_48060);
nor UO_3753 (O_3753,N_47963,N_45794);
nor UO_3754 (O_3754,N_49012,N_46790);
xor UO_3755 (O_3755,N_49336,N_48303);
xor UO_3756 (O_3756,N_45126,N_48492);
nor UO_3757 (O_3757,N_49810,N_46481);
nand UO_3758 (O_3758,N_47271,N_47667);
or UO_3759 (O_3759,N_49857,N_47767);
nor UO_3760 (O_3760,N_49928,N_45956);
or UO_3761 (O_3761,N_47552,N_45874);
nand UO_3762 (O_3762,N_45778,N_47669);
and UO_3763 (O_3763,N_49968,N_49964);
nand UO_3764 (O_3764,N_46493,N_47408);
and UO_3765 (O_3765,N_48481,N_46945);
xnor UO_3766 (O_3766,N_48819,N_46660);
xor UO_3767 (O_3767,N_47251,N_49424);
or UO_3768 (O_3768,N_46156,N_48790);
xnor UO_3769 (O_3769,N_48129,N_49576);
nand UO_3770 (O_3770,N_49779,N_47542);
xnor UO_3771 (O_3771,N_46206,N_49992);
or UO_3772 (O_3772,N_49885,N_45902);
xor UO_3773 (O_3773,N_48973,N_48082);
and UO_3774 (O_3774,N_45394,N_47003);
nor UO_3775 (O_3775,N_46040,N_48083);
xnor UO_3776 (O_3776,N_49471,N_46228);
xor UO_3777 (O_3777,N_47910,N_45490);
xor UO_3778 (O_3778,N_47581,N_46905);
nand UO_3779 (O_3779,N_49266,N_46065);
nor UO_3780 (O_3780,N_48030,N_49237);
and UO_3781 (O_3781,N_47171,N_49249);
and UO_3782 (O_3782,N_45958,N_47101);
xor UO_3783 (O_3783,N_45525,N_47756);
nor UO_3784 (O_3784,N_46091,N_48046);
xor UO_3785 (O_3785,N_49996,N_48575);
and UO_3786 (O_3786,N_47978,N_46255);
xnor UO_3787 (O_3787,N_47539,N_49022);
nor UO_3788 (O_3788,N_45414,N_46809);
xnor UO_3789 (O_3789,N_45609,N_45393);
and UO_3790 (O_3790,N_45786,N_46621);
xor UO_3791 (O_3791,N_49533,N_46212);
xnor UO_3792 (O_3792,N_48466,N_49327);
or UO_3793 (O_3793,N_46416,N_45767);
and UO_3794 (O_3794,N_45126,N_48625);
nand UO_3795 (O_3795,N_47972,N_49356);
nor UO_3796 (O_3796,N_49064,N_45456);
nand UO_3797 (O_3797,N_47065,N_46382);
or UO_3798 (O_3798,N_48076,N_47365);
and UO_3799 (O_3799,N_49083,N_45352);
xnor UO_3800 (O_3800,N_47395,N_46987);
xnor UO_3801 (O_3801,N_49548,N_47215);
xor UO_3802 (O_3802,N_48597,N_48367);
or UO_3803 (O_3803,N_46064,N_45607);
xor UO_3804 (O_3804,N_46894,N_48879);
nor UO_3805 (O_3805,N_49518,N_47592);
nor UO_3806 (O_3806,N_48025,N_46252);
and UO_3807 (O_3807,N_45393,N_47174);
or UO_3808 (O_3808,N_48349,N_46909);
nand UO_3809 (O_3809,N_49269,N_48630);
xnor UO_3810 (O_3810,N_48688,N_46553);
nor UO_3811 (O_3811,N_45286,N_48051);
or UO_3812 (O_3812,N_48601,N_46067);
nand UO_3813 (O_3813,N_47008,N_48641);
and UO_3814 (O_3814,N_48224,N_47582);
nor UO_3815 (O_3815,N_48102,N_48830);
nand UO_3816 (O_3816,N_47989,N_47814);
and UO_3817 (O_3817,N_45320,N_49543);
xnor UO_3818 (O_3818,N_49017,N_47154);
or UO_3819 (O_3819,N_46371,N_49207);
or UO_3820 (O_3820,N_49322,N_45540);
or UO_3821 (O_3821,N_49579,N_45769);
and UO_3822 (O_3822,N_48671,N_49007);
nand UO_3823 (O_3823,N_46392,N_48339);
nor UO_3824 (O_3824,N_46404,N_45808);
xnor UO_3825 (O_3825,N_46658,N_49734);
nand UO_3826 (O_3826,N_49374,N_49257);
nor UO_3827 (O_3827,N_45375,N_48969);
and UO_3828 (O_3828,N_49293,N_47803);
xor UO_3829 (O_3829,N_49966,N_49782);
and UO_3830 (O_3830,N_47723,N_47711);
nor UO_3831 (O_3831,N_49874,N_49712);
xnor UO_3832 (O_3832,N_49103,N_45479);
nor UO_3833 (O_3833,N_45379,N_46548);
or UO_3834 (O_3834,N_45404,N_45396);
xor UO_3835 (O_3835,N_45444,N_45224);
nand UO_3836 (O_3836,N_46588,N_45164);
nor UO_3837 (O_3837,N_45167,N_48984);
and UO_3838 (O_3838,N_45505,N_45897);
and UO_3839 (O_3839,N_47119,N_47673);
or UO_3840 (O_3840,N_48981,N_48109);
or UO_3841 (O_3841,N_49755,N_46337);
and UO_3842 (O_3842,N_45385,N_48736);
and UO_3843 (O_3843,N_46961,N_48327);
xnor UO_3844 (O_3844,N_45674,N_48098);
and UO_3845 (O_3845,N_48219,N_45324);
and UO_3846 (O_3846,N_46931,N_46255);
xor UO_3847 (O_3847,N_48429,N_48864);
xor UO_3848 (O_3848,N_45249,N_47861);
nor UO_3849 (O_3849,N_45508,N_45553);
nand UO_3850 (O_3850,N_48969,N_47496);
nand UO_3851 (O_3851,N_49961,N_47378);
and UO_3852 (O_3852,N_45561,N_47793);
and UO_3853 (O_3853,N_48918,N_46843);
xor UO_3854 (O_3854,N_49371,N_49715);
nor UO_3855 (O_3855,N_45997,N_45488);
or UO_3856 (O_3856,N_45803,N_46099);
or UO_3857 (O_3857,N_47541,N_46450);
or UO_3858 (O_3858,N_49959,N_47945);
and UO_3859 (O_3859,N_48214,N_47160);
or UO_3860 (O_3860,N_45768,N_47955);
nor UO_3861 (O_3861,N_48668,N_46164);
nor UO_3862 (O_3862,N_48202,N_48971);
nand UO_3863 (O_3863,N_47070,N_47824);
nand UO_3864 (O_3864,N_45941,N_48900);
xor UO_3865 (O_3865,N_48486,N_45108);
or UO_3866 (O_3866,N_45102,N_49202);
and UO_3867 (O_3867,N_49856,N_46344);
and UO_3868 (O_3868,N_47777,N_48492);
or UO_3869 (O_3869,N_49491,N_45437);
nand UO_3870 (O_3870,N_46724,N_48842);
nor UO_3871 (O_3871,N_46691,N_49511);
nor UO_3872 (O_3872,N_45225,N_48862);
nand UO_3873 (O_3873,N_45141,N_48371);
nand UO_3874 (O_3874,N_49082,N_45011);
nand UO_3875 (O_3875,N_48724,N_47281);
or UO_3876 (O_3876,N_48288,N_45239);
and UO_3877 (O_3877,N_46192,N_45640);
nand UO_3878 (O_3878,N_45574,N_48565);
nor UO_3879 (O_3879,N_47536,N_47309);
nand UO_3880 (O_3880,N_45042,N_47013);
and UO_3881 (O_3881,N_45280,N_49592);
and UO_3882 (O_3882,N_45876,N_45117);
or UO_3883 (O_3883,N_49619,N_47193);
nor UO_3884 (O_3884,N_48906,N_45415);
and UO_3885 (O_3885,N_45783,N_48841);
nor UO_3886 (O_3886,N_49619,N_48310);
nor UO_3887 (O_3887,N_48849,N_49542);
nand UO_3888 (O_3888,N_48524,N_48289);
and UO_3889 (O_3889,N_48896,N_46203);
and UO_3890 (O_3890,N_49509,N_48067);
or UO_3891 (O_3891,N_47238,N_49881);
or UO_3892 (O_3892,N_45172,N_49483);
and UO_3893 (O_3893,N_47578,N_46009);
and UO_3894 (O_3894,N_48656,N_47394);
or UO_3895 (O_3895,N_47782,N_49585);
xor UO_3896 (O_3896,N_45592,N_47137);
xor UO_3897 (O_3897,N_48978,N_49017);
and UO_3898 (O_3898,N_45322,N_47165);
nor UO_3899 (O_3899,N_48839,N_46493);
nor UO_3900 (O_3900,N_48855,N_48715);
nand UO_3901 (O_3901,N_45790,N_47537);
and UO_3902 (O_3902,N_45808,N_48512);
nor UO_3903 (O_3903,N_46335,N_45735);
or UO_3904 (O_3904,N_48620,N_46217);
nand UO_3905 (O_3905,N_46247,N_48710);
nor UO_3906 (O_3906,N_48522,N_49681);
xnor UO_3907 (O_3907,N_46724,N_45439);
or UO_3908 (O_3908,N_45847,N_45639);
nor UO_3909 (O_3909,N_48240,N_47795);
or UO_3910 (O_3910,N_46385,N_47922);
xnor UO_3911 (O_3911,N_45991,N_46328);
nor UO_3912 (O_3912,N_45734,N_47899);
and UO_3913 (O_3913,N_47985,N_49284);
nand UO_3914 (O_3914,N_49748,N_49086);
or UO_3915 (O_3915,N_47305,N_48697);
xnor UO_3916 (O_3916,N_45010,N_46634);
nand UO_3917 (O_3917,N_47227,N_48747);
and UO_3918 (O_3918,N_48037,N_46701);
or UO_3919 (O_3919,N_46555,N_46854);
nand UO_3920 (O_3920,N_49338,N_48933);
nor UO_3921 (O_3921,N_45090,N_45467);
or UO_3922 (O_3922,N_47530,N_49923);
and UO_3923 (O_3923,N_49151,N_46668);
and UO_3924 (O_3924,N_49389,N_49917);
xor UO_3925 (O_3925,N_47310,N_48907);
nand UO_3926 (O_3926,N_46883,N_47609);
xnor UO_3927 (O_3927,N_48391,N_45869);
xor UO_3928 (O_3928,N_49757,N_48592);
or UO_3929 (O_3929,N_48458,N_47593);
nand UO_3930 (O_3930,N_48181,N_46839);
xor UO_3931 (O_3931,N_47429,N_46285);
nor UO_3932 (O_3932,N_45927,N_46166);
nand UO_3933 (O_3933,N_48902,N_48647);
nor UO_3934 (O_3934,N_45565,N_47635);
nor UO_3935 (O_3935,N_49067,N_49823);
nor UO_3936 (O_3936,N_46498,N_48394);
nor UO_3937 (O_3937,N_45703,N_46055);
xor UO_3938 (O_3938,N_45462,N_47350);
or UO_3939 (O_3939,N_47055,N_45701);
nand UO_3940 (O_3940,N_47208,N_45926);
or UO_3941 (O_3941,N_45276,N_46595);
nand UO_3942 (O_3942,N_45345,N_48496);
or UO_3943 (O_3943,N_45963,N_49419);
or UO_3944 (O_3944,N_49687,N_46929);
xnor UO_3945 (O_3945,N_46336,N_45148);
nand UO_3946 (O_3946,N_48314,N_46377);
or UO_3947 (O_3947,N_45634,N_47175);
nand UO_3948 (O_3948,N_46459,N_47305);
xor UO_3949 (O_3949,N_46303,N_48404);
or UO_3950 (O_3950,N_47052,N_47643);
and UO_3951 (O_3951,N_49742,N_49180);
xnor UO_3952 (O_3952,N_47730,N_46041);
xor UO_3953 (O_3953,N_47051,N_46565);
and UO_3954 (O_3954,N_48275,N_46993);
and UO_3955 (O_3955,N_47192,N_47482);
xnor UO_3956 (O_3956,N_47001,N_46693);
or UO_3957 (O_3957,N_46761,N_45441);
nor UO_3958 (O_3958,N_46786,N_45523);
or UO_3959 (O_3959,N_46093,N_45768);
or UO_3960 (O_3960,N_47403,N_48870);
or UO_3961 (O_3961,N_48080,N_49670);
nand UO_3962 (O_3962,N_45390,N_46418);
xor UO_3963 (O_3963,N_48059,N_45216);
or UO_3964 (O_3964,N_48271,N_46922);
and UO_3965 (O_3965,N_45816,N_47890);
nor UO_3966 (O_3966,N_48397,N_48105);
nand UO_3967 (O_3967,N_48149,N_45520);
nor UO_3968 (O_3968,N_46051,N_46343);
or UO_3969 (O_3969,N_49074,N_47034);
nand UO_3970 (O_3970,N_45864,N_47547);
nor UO_3971 (O_3971,N_49341,N_49042);
or UO_3972 (O_3972,N_46918,N_47980);
nor UO_3973 (O_3973,N_45993,N_49345);
nor UO_3974 (O_3974,N_47539,N_48809);
and UO_3975 (O_3975,N_48907,N_46488);
nor UO_3976 (O_3976,N_49214,N_45203);
nor UO_3977 (O_3977,N_48614,N_48270);
and UO_3978 (O_3978,N_49808,N_46124);
or UO_3979 (O_3979,N_48920,N_45256);
nand UO_3980 (O_3980,N_45802,N_47957);
or UO_3981 (O_3981,N_45626,N_45796);
nor UO_3982 (O_3982,N_47636,N_48925);
nor UO_3983 (O_3983,N_45462,N_45945);
and UO_3984 (O_3984,N_45961,N_48515);
nand UO_3985 (O_3985,N_46214,N_46812);
xor UO_3986 (O_3986,N_47790,N_46386);
xor UO_3987 (O_3987,N_48901,N_48702);
xnor UO_3988 (O_3988,N_45354,N_46484);
and UO_3989 (O_3989,N_46570,N_45430);
and UO_3990 (O_3990,N_48474,N_45418);
xnor UO_3991 (O_3991,N_46492,N_48684);
or UO_3992 (O_3992,N_48488,N_48365);
nor UO_3993 (O_3993,N_47556,N_45045);
xnor UO_3994 (O_3994,N_49486,N_49120);
nor UO_3995 (O_3995,N_49795,N_49035);
nor UO_3996 (O_3996,N_47925,N_47217);
or UO_3997 (O_3997,N_49973,N_45926);
xnor UO_3998 (O_3998,N_45056,N_47204);
nor UO_3999 (O_3999,N_45985,N_47505);
or UO_4000 (O_4000,N_48536,N_45850);
nor UO_4001 (O_4001,N_46576,N_45077);
xor UO_4002 (O_4002,N_48056,N_46588);
or UO_4003 (O_4003,N_45252,N_46890);
nand UO_4004 (O_4004,N_47112,N_49740);
nand UO_4005 (O_4005,N_48792,N_49874);
or UO_4006 (O_4006,N_49372,N_46562);
and UO_4007 (O_4007,N_48644,N_45232);
nand UO_4008 (O_4008,N_48092,N_47119);
nor UO_4009 (O_4009,N_45522,N_46243);
nand UO_4010 (O_4010,N_47919,N_46857);
and UO_4011 (O_4011,N_48457,N_45470);
xnor UO_4012 (O_4012,N_49876,N_45913);
nor UO_4013 (O_4013,N_48980,N_47038);
xor UO_4014 (O_4014,N_47845,N_49912);
xnor UO_4015 (O_4015,N_49146,N_45436);
and UO_4016 (O_4016,N_48372,N_46806);
and UO_4017 (O_4017,N_48038,N_46765);
and UO_4018 (O_4018,N_45278,N_46122);
nor UO_4019 (O_4019,N_45140,N_48502);
and UO_4020 (O_4020,N_48643,N_48133);
or UO_4021 (O_4021,N_45253,N_45329);
nor UO_4022 (O_4022,N_45098,N_45867);
xnor UO_4023 (O_4023,N_48348,N_46424);
or UO_4024 (O_4024,N_49863,N_48804);
xnor UO_4025 (O_4025,N_47964,N_48835);
nand UO_4026 (O_4026,N_46396,N_45537);
xor UO_4027 (O_4027,N_46659,N_47282);
nand UO_4028 (O_4028,N_49503,N_45827);
xnor UO_4029 (O_4029,N_48944,N_46910);
nand UO_4030 (O_4030,N_49843,N_45263);
nor UO_4031 (O_4031,N_48183,N_49993);
and UO_4032 (O_4032,N_49228,N_47201);
nor UO_4033 (O_4033,N_45981,N_49813);
xnor UO_4034 (O_4034,N_47747,N_46449);
nand UO_4035 (O_4035,N_46039,N_47392);
and UO_4036 (O_4036,N_46109,N_45576);
nand UO_4037 (O_4037,N_45017,N_45931);
nand UO_4038 (O_4038,N_47083,N_46683);
nor UO_4039 (O_4039,N_45627,N_46444);
xnor UO_4040 (O_4040,N_48201,N_47879);
xor UO_4041 (O_4041,N_47447,N_46177);
nor UO_4042 (O_4042,N_47110,N_47486);
xor UO_4043 (O_4043,N_45817,N_45573);
xor UO_4044 (O_4044,N_47065,N_46975);
nand UO_4045 (O_4045,N_49370,N_47782);
and UO_4046 (O_4046,N_49125,N_49576);
nor UO_4047 (O_4047,N_47237,N_49055);
and UO_4048 (O_4048,N_48379,N_45763);
or UO_4049 (O_4049,N_47052,N_49410);
nand UO_4050 (O_4050,N_47047,N_45280);
or UO_4051 (O_4051,N_45726,N_48551);
xor UO_4052 (O_4052,N_46929,N_49062);
xnor UO_4053 (O_4053,N_45626,N_48950);
or UO_4054 (O_4054,N_47651,N_47776);
xnor UO_4055 (O_4055,N_48102,N_48221);
or UO_4056 (O_4056,N_48756,N_45838);
nand UO_4057 (O_4057,N_46945,N_47747);
or UO_4058 (O_4058,N_48217,N_47898);
nor UO_4059 (O_4059,N_45536,N_49445);
xnor UO_4060 (O_4060,N_46403,N_49901);
xnor UO_4061 (O_4061,N_46459,N_45183);
nor UO_4062 (O_4062,N_45640,N_48590);
and UO_4063 (O_4063,N_45214,N_45649);
nand UO_4064 (O_4064,N_49222,N_49264);
nand UO_4065 (O_4065,N_48476,N_46810);
or UO_4066 (O_4066,N_48175,N_45121);
nand UO_4067 (O_4067,N_46613,N_48313);
xor UO_4068 (O_4068,N_49833,N_45663);
and UO_4069 (O_4069,N_46825,N_46510);
nor UO_4070 (O_4070,N_49076,N_48056);
xnor UO_4071 (O_4071,N_45710,N_46199);
and UO_4072 (O_4072,N_45168,N_46998);
nor UO_4073 (O_4073,N_47114,N_48844);
nand UO_4074 (O_4074,N_49107,N_49473);
xor UO_4075 (O_4075,N_47013,N_46519);
and UO_4076 (O_4076,N_47181,N_48079);
and UO_4077 (O_4077,N_48623,N_48446);
and UO_4078 (O_4078,N_48656,N_48009);
xor UO_4079 (O_4079,N_47780,N_49726);
and UO_4080 (O_4080,N_48155,N_49123);
or UO_4081 (O_4081,N_49872,N_45057);
and UO_4082 (O_4082,N_46528,N_47375);
xor UO_4083 (O_4083,N_47295,N_46340);
nor UO_4084 (O_4084,N_48992,N_48610);
and UO_4085 (O_4085,N_49717,N_46233);
nand UO_4086 (O_4086,N_45339,N_45042);
xnor UO_4087 (O_4087,N_47762,N_48246);
or UO_4088 (O_4088,N_49622,N_45919);
nand UO_4089 (O_4089,N_45147,N_46980);
or UO_4090 (O_4090,N_48442,N_47473);
and UO_4091 (O_4091,N_46376,N_49690);
nor UO_4092 (O_4092,N_46132,N_49256);
and UO_4093 (O_4093,N_48972,N_48382);
nand UO_4094 (O_4094,N_46878,N_47311);
or UO_4095 (O_4095,N_46593,N_49650);
or UO_4096 (O_4096,N_47264,N_47880);
nor UO_4097 (O_4097,N_45766,N_47136);
nand UO_4098 (O_4098,N_45113,N_46995);
nand UO_4099 (O_4099,N_49426,N_48175);
and UO_4100 (O_4100,N_49959,N_48037);
nor UO_4101 (O_4101,N_46205,N_45813);
nand UO_4102 (O_4102,N_46163,N_48294);
nand UO_4103 (O_4103,N_46405,N_45257);
xor UO_4104 (O_4104,N_47387,N_46145);
xor UO_4105 (O_4105,N_49033,N_49685);
nor UO_4106 (O_4106,N_48210,N_48865);
or UO_4107 (O_4107,N_47616,N_49007);
or UO_4108 (O_4108,N_45981,N_47798);
xnor UO_4109 (O_4109,N_48004,N_47278);
or UO_4110 (O_4110,N_45888,N_46213);
nand UO_4111 (O_4111,N_45963,N_48878);
nand UO_4112 (O_4112,N_46251,N_46237);
nor UO_4113 (O_4113,N_45406,N_45134);
and UO_4114 (O_4114,N_47251,N_45538);
xor UO_4115 (O_4115,N_45306,N_49650);
and UO_4116 (O_4116,N_48566,N_47080);
nor UO_4117 (O_4117,N_49632,N_49067);
nand UO_4118 (O_4118,N_45267,N_45513);
nand UO_4119 (O_4119,N_45778,N_49999);
xnor UO_4120 (O_4120,N_48294,N_49357);
nand UO_4121 (O_4121,N_47401,N_46691);
or UO_4122 (O_4122,N_46057,N_48978);
and UO_4123 (O_4123,N_46414,N_46468);
and UO_4124 (O_4124,N_45941,N_48861);
or UO_4125 (O_4125,N_46843,N_48182);
xnor UO_4126 (O_4126,N_47238,N_46712);
xor UO_4127 (O_4127,N_45608,N_49279);
nand UO_4128 (O_4128,N_45301,N_46540);
nor UO_4129 (O_4129,N_46025,N_46521);
and UO_4130 (O_4130,N_46076,N_46027);
and UO_4131 (O_4131,N_48954,N_46584);
nor UO_4132 (O_4132,N_49220,N_47866);
nor UO_4133 (O_4133,N_46599,N_46094);
and UO_4134 (O_4134,N_46974,N_46663);
or UO_4135 (O_4135,N_45909,N_45080);
xnor UO_4136 (O_4136,N_45104,N_48559);
and UO_4137 (O_4137,N_45078,N_45736);
xor UO_4138 (O_4138,N_48211,N_49739);
or UO_4139 (O_4139,N_48594,N_47032);
nand UO_4140 (O_4140,N_49779,N_45256);
xor UO_4141 (O_4141,N_46735,N_46390);
or UO_4142 (O_4142,N_45009,N_46381);
and UO_4143 (O_4143,N_48256,N_45788);
nand UO_4144 (O_4144,N_48579,N_48163);
nor UO_4145 (O_4145,N_48322,N_48762);
and UO_4146 (O_4146,N_47507,N_49191);
nor UO_4147 (O_4147,N_46839,N_49678);
nand UO_4148 (O_4148,N_47713,N_46625);
or UO_4149 (O_4149,N_48009,N_47335);
or UO_4150 (O_4150,N_49027,N_48965);
and UO_4151 (O_4151,N_46156,N_46019);
and UO_4152 (O_4152,N_49354,N_48137);
or UO_4153 (O_4153,N_46292,N_47100);
and UO_4154 (O_4154,N_48771,N_49311);
and UO_4155 (O_4155,N_49110,N_48077);
or UO_4156 (O_4156,N_49998,N_45201);
or UO_4157 (O_4157,N_45442,N_48267);
xor UO_4158 (O_4158,N_48227,N_45681);
or UO_4159 (O_4159,N_46490,N_49474);
nor UO_4160 (O_4160,N_49751,N_45743);
or UO_4161 (O_4161,N_46733,N_49917);
and UO_4162 (O_4162,N_47559,N_46686);
nand UO_4163 (O_4163,N_47583,N_45548);
nor UO_4164 (O_4164,N_45001,N_49295);
or UO_4165 (O_4165,N_49198,N_45659);
nor UO_4166 (O_4166,N_48580,N_45361);
or UO_4167 (O_4167,N_47964,N_45033);
xor UO_4168 (O_4168,N_48666,N_46971);
xor UO_4169 (O_4169,N_49471,N_49184);
or UO_4170 (O_4170,N_45151,N_47810);
or UO_4171 (O_4171,N_45299,N_45218);
or UO_4172 (O_4172,N_47820,N_47626);
and UO_4173 (O_4173,N_48201,N_46551);
nand UO_4174 (O_4174,N_46484,N_48938);
and UO_4175 (O_4175,N_45634,N_47365);
nand UO_4176 (O_4176,N_47779,N_48159);
or UO_4177 (O_4177,N_46168,N_48149);
or UO_4178 (O_4178,N_48271,N_49182);
xnor UO_4179 (O_4179,N_47169,N_49952);
and UO_4180 (O_4180,N_45682,N_45462);
and UO_4181 (O_4181,N_47173,N_46839);
and UO_4182 (O_4182,N_45651,N_47350);
nor UO_4183 (O_4183,N_47192,N_45203);
xor UO_4184 (O_4184,N_49809,N_49117);
xor UO_4185 (O_4185,N_48946,N_49076);
and UO_4186 (O_4186,N_48888,N_48042);
nor UO_4187 (O_4187,N_47829,N_48223);
or UO_4188 (O_4188,N_45011,N_47778);
nand UO_4189 (O_4189,N_45175,N_47219);
nor UO_4190 (O_4190,N_46245,N_48787);
or UO_4191 (O_4191,N_49410,N_48885);
nor UO_4192 (O_4192,N_49343,N_49834);
or UO_4193 (O_4193,N_48075,N_47956);
and UO_4194 (O_4194,N_48301,N_45212);
nand UO_4195 (O_4195,N_46078,N_49042);
and UO_4196 (O_4196,N_46829,N_47808);
nor UO_4197 (O_4197,N_49150,N_49951);
nor UO_4198 (O_4198,N_48427,N_47670);
nor UO_4199 (O_4199,N_45728,N_48110);
nand UO_4200 (O_4200,N_45823,N_45519);
xor UO_4201 (O_4201,N_48465,N_49068);
nand UO_4202 (O_4202,N_45867,N_45857);
xnor UO_4203 (O_4203,N_47461,N_47879);
xnor UO_4204 (O_4204,N_48152,N_45433);
nor UO_4205 (O_4205,N_49403,N_47434);
nor UO_4206 (O_4206,N_48804,N_49891);
and UO_4207 (O_4207,N_48958,N_49831);
nand UO_4208 (O_4208,N_49809,N_49619);
and UO_4209 (O_4209,N_45238,N_48705);
and UO_4210 (O_4210,N_45880,N_47948);
or UO_4211 (O_4211,N_45082,N_48104);
nand UO_4212 (O_4212,N_48220,N_46157);
xnor UO_4213 (O_4213,N_47258,N_45943);
and UO_4214 (O_4214,N_46086,N_47065);
nand UO_4215 (O_4215,N_45590,N_45632);
nand UO_4216 (O_4216,N_49802,N_47433);
nor UO_4217 (O_4217,N_46953,N_48500);
or UO_4218 (O_4218,N_45921,N_46396);
nor UO_4219 (O_4219,N_47981,N_45323);
nor UO_4220 (O_4220,N_47577,N_49586);
and UO_4221 (O_4221,N_46979,N_48505);
nor UO_4222 (O_4222,N_45838,N_45712);
nor UO_4223 (O_4223,N_49489,N_46284);
nor UO_4224 (O_4224,N_48909,N_45352);
or UO_4225 (O_4225,N_48074,N_48216);
or UO_4226 (O_4226,N_47450,N_49632);
nand UO_4227 (O_4227,N_49167,N_47959);
nor UO_4228 (O_4228,N_48880,N_49621);
nor UO_4229 (O_4229,N_49430,N_47313);
or UO_4230 (O_4230,N_46097,N_49999);
or UO_4231 (O_4231,N_45998,N_46233);
xnor UO_4232 (O_4232,N_47205,N_45559);
or UO_4233 (O_4233,N_47161,N_46269);
xnor UO_4234 (O_4234,N_48059,N_47368);
and UO_4235 (O_4235,N_48094,N_47275);
nor UO_4236 (O_4236,N_49897,N_48683);
or UO_4237 (O_4237,N_48824,N_48908);
xor UO_4238 (O_4238,N_46751,N_46973);
or UO_4239 (O_4239,N_45170,N_47900);
nand UO_4240 (O_4240,N_45256,N_45512);
and UO_4241 (O_4241,N_45400,N_49980);
xnor UO_4242 (O_4242,N_48248,N_49562);
xnor UO_4243 (O_4243,N_49921,N_46294);
or UO_4244 (O_4244,N_48402,N_49097);
or UO_4245 (O_4245,N_47775,N_45876);
nor UO_4246 (O_4246,N_49574,N_49733);
xor UO_4247 (O_4247,N_49317,N_48396);
nor UO_4248 (O_4248,N_46811,N_45641);
or UO_4249 (O_4249,N_47099,N_46833);
xnor UO_4250 (O_4250,N_49751,N_45326);
and UO_4251 (O_4251,N_45050,N_45450);
xor UO_4252 (O_4252,N_49611,N_46896);
or UO_4253 (O_4253,N_45734,N_45908);
or UO_4254 (O_4254,N_47299,N_47081);
nand UO_4255 (O_4255,N_48622,N_48187);
or UO_4256 (O_4256,N_48922,N_47143);
or UO_4257 (O_4257,N_46690,N_47108);
or UO_4258 (O_4258,N_46073,N_46550);
nand UO_4259 (O_4259,N_47211,N_47766);
and UO_4260 (O_4260,N_48031,N_49851);
and UO_4261 (O_4261,N_45591,N_49804);
nor UO_4262 (O_4262,N_47933,N_48920);
and UO_4263 (O_4263,N_47186,N_47087);
nand UO_4264 (O_4264,N_46851,N_47803);
or UO_4265 (O_4265,N_47239,N_45362);
nand UO_4266 (O_4266,N_49923,N_48462);
xor UO_4267 (O_4267,N_46626,N_48894);
xnor UO_4268 (O_4268,N_48959,N_47984);
nor UO_4269 (O_4269,N_49053,N_46477);
nand UO_4270 (O_4270,N_46347,N_48788);
or UO_4271 (O_4271,N_48952,N_46907);
xnor UO_4272 (O_4272,N_47547,N_47657);
nand UO_4273 (O_4273,N_47717,N_47249);
nor UO_4274 (O_4274,N_45847,N_46724);
nor UO_4275 (O_4275,N_47307,N_47425);
and UO_4276 (O_4276,N_49747,N_46043);
or UO_4277 (O_4277,N_46286,N_47453);
or UO_4278 (O_4278,N_47448,N_47891);
and UO_4279 (O_4279,N_49945,N_48744);
or UO_4280 (O_4280,N_46983,N_48599);
or UO_4281 (O_4281,N_45090,N_48577);
or UO_4282 (O_4282,N_48077,N_45636);
and UO_4283 (O_4283,N_45267,N_49215);
or UO_4284 (O_4284,N_49698,N_49662);
or UO_4285 (O_4285,N_45726,N_45100);
xor UO_4286 (O_4286,N_47332,N_47670);
and UO_4287 (O_4287,N_48604,N_47232);
or UO_4288 (O_4288,N_46823,N_49533);
and UO_4289 (O_4289,N_48290,N_49906);
nor UO_4290 (O_4290,N_49837,N_45780);
and UO_4291 (O_4291,N_46427,N_46794);
nor UO_4292 (O_4292,N_46461,N_47815);
nand UO_4293 (O_4293,N_49628,N_45453);
or UO_4294 (O_4294,N_46456,N_46423);
nor UO_4295 (O_4295,N_49661,N_49697);
and UO_4296 (O_4296,N_47830,N_47251);
nand UO_4297 (O_4297,N_46387,N_45445);
and UO_4298 (O_4298,N_49056,N_47634);
xor UO_4299 (O_4299,N_48338,N_49700);
xnor UO_4300 (O_4300,N_46330,N_46562);
and UO_4301 (O_4301,N_46941,N_46653);
and UO_4302 (O_4302,N_47897,N_48341);
nor UO_4303 (O_4303,N_48240,N_47242);
xnor UO_4304 (O_4304,N_47684,N_45703);
xor UO_4305 (O_4305,N_49078,N_49322);
nand UO_4306 (O_4306,N_47474,N_48293);
or UO_4307 (O_4307,N_49817,N_49135);
and UO_4308 (O_4308,N_45382,N_45697);
xor UO_4309 (O_4309,N_48043,N_47624);
nor UO_4310 (O_4310,N_45624,N_47346);
xnor UO_4311 (O_4311,N_45833,N_49586);
and UO_4312 (O_4312,N_47905,N_48433);
and UO_4313 (O_4313,N_49059,N_47973);
xor UO_4314 (O_4314,N_49292,N_49677);
xnor UO_4315 (O_4315,N_49033,N_47277);
nor UO_4316 (O_4316,N_48903,N_48351);
or UO_4317 (O_4317,N_49830,N_46532);
and UO_4318 (O_4318,N_46724,N_49206);
xor UO_4319 (O_4319,N_45618,N_45420);
or UO_4320 (O_4320,N_47444,N_46651);
nand UO_4321 (O_4321,N_48895,N_47742);
nand UO_4322 (O_4322,N_49276,N_47326);
nor UO_4323 (O_4323,N_49269,N_48873);
nand UO_4324 (O_4324,N_49245,N_48982);
nand UO_4325 (O_4325,N_49022,N_49770);
nor UO_4326 (O_4326,N_46624,N_46347);
and UO_4327 (O_4327,N_47932,N_47232);
and UO_4328 (O_4328,N_45584,N_47837);
nor UO_4329 (O_4329,N_46593,N_49744);
nor UO_4330 (O_4330,N_49690,N_48551);
or UO_4331 (O_4331,N_46002,N_45493);
xor UO_4332 (O_4332,N_46918,N_47848);
nor UO_4333 (O_4333,N_48986,N_46147);
or UO_4334 (O_4334,N_47180,N_47317);
or UO_4335 (O_4335,N_46278,N_47601);
nand UO_4336 (O_4336,N_45664,N_47351);
nor UO_4337 (O_4337,N_48976,N_47599);
xnor UO_4338 (O_4338,N_47038,N_46135);
and UO_4339 (O_4339,N_48364,N_45505);
or UO_4340 (O_4340,N_46886,N_47710);
xor UO_4341 (O_4341,N_49205,N_49047);
or UO_4342 (O_4342,N_48390,N_45869);
nor UO_4343 (O_4343,N_46206,N_49910);
and UO_4344 (O_4344,N_46156,N_48405);
or UO_4345 (O_4345,N_48451,N_47306);
or UO_4346 (O_4346,N_49882,N_46242);
or UO_4347 (O_4347,N_46127,N_48832);
or UO_4348 (O_4348,N_46556,N_47354);
nand UO_4349 (O_4349,N_45900,N_48672);
and UO_4350 (O_4350,N_47473,N_47842);
or UO_4351 (O_4351,N_46592,N_49291);
or UO_4352 (O_4352,N_47785,N_48306);
nor UO_4353 (O_4353,N_46443,N_47084);
and UO_4354 (O_4354,N_48072,N_45356);
nor UO_4355 (O_4355,N_49079,N_46458);
nor UO_4356 (O_4356,N_48676,N_45764);
nand UO_4357 (O_4357,N_49066,N_48745);
or UO_4358 (O_4358,N_48739,N_48444);
and UO_4359 (O_4359,N_47351,N_45569);
nor UO_4360 (O_4360,N_46622,N_45798);
nand UO_4361 (O_4361,N_45731,N_49747);
xnor UO_4362 (O_4362,N_46975,N_46262);
or UO_4363 (O_4363,N_49518,N_45990);
and UO_4364 (O_4364,N_47138,N_47703);
nor UO_4365 (O_4365,N_48793,N_47004);
nand UO_4366 (O_4366,N_47054,N_45857);
nand UO_4367 (O_4367,N_47332,N_46672);
nand UO_4368 (O_4368,N_48513,N_49432);
nor UO_4369 (O_4369,N_49929,N_48141);
nor UO_4370 (O_4370,N_47704,N_48318);
or UO_4371 (O_4371,N_49021,N_46543);
or UO_4372 (O_4372,N_47866,N_46124);
xor UO_4373 (O_4373,N_48419,N_46154);
or UO_4374 (O_4374,N_45359,N_49771);
xor UO_4375 (O_4375,N_45872,N_46540);
or UO_4376 (O_4376,N_45366,N_45646);
xnor UO_4377 (O_4377,N_49137,N_47058);
nor UO_4378 (O_4378,N_46818,N_45704);
xnor UO_4379 (O_4379,N_47701,N_45558);
nor UO_4380 (O_4380,N_49913,N_46675);
nand UO_4381 (O_4381,N_48068,N_46612);
and UO_4382 (O_4382,N_48024,N_45675);
xnor UO_4383 (O_4383,N_49608,N_49136);
xnor UO_4384 (O_4384,N_48193,N_45757);
and UO_4385 (O_4385,N_47728,N_45031);
xor UO_4386 (O_4386,N_46481,N_49797);
xor UO_4387 (O_4387,N_49627,N_45900);
and UO_4388 (O_4388,N_45354,N_48166);
and UO_4389 (O_4389,N_46969,N_46975);
or UO_4390 (O_4390,N_45634,N_48867);
and UO_4391 (O_4391,N_45863,N_49474);
nor UO_4392 (O_4392,N_48411,N_49328);
nor UO_4393 (O_4393,N_45659,N_49069);
and UO_4394 (O_4394,N_49632,N_46280);
or UO_4395 (O_4395,N_48864,N_48185);
or UO_4396 (O_4396,N_47752,N_47732);
and UO_4397 (O_4397,N_47568,N_48565);
nor UO_4398 (O_4398,N_46763,N_46225);
xor UO_4399 (O_4399,N_47509,N_47426);
nand UO_4400 (O_4400,N_45983,N_49320);
xor UO_4401 (O_4401,N_45935,N_47391);
or UO_4402 (O_4402,N_47875,N_49958);
nor UO_4403 (O_4403,N_49175,N_46839);
nor UO_4404 (O_4404,N_47293,N_45373);
and UO_4405 (O_4405,N_45372,N_49003);
nand UO_4406 (O_4406,N_47895,N_48077);
nor UO_4407 (O_4407,N_47955,N_45803);
or UO_4408 (O_4408,N_47541,N_49939);
or UO_4409 (O_4409,N_48593,N_48624);
or UO_4410 (O_4410,N_48112,N_48861);
or UO_4411 (O_4411,N_46847,N_48613);
nor UO_4412 (O_4412,N_49736,N_47583);
or UO_4413 (O_4413,N_47454,N_47717);
xnor UO_4414 (O_4414,N_45435,N_49881);
nor UO_4415 (O_4415,N_49750,N_47476);
nor UO_4416 (O_4416,N_48866,N_47124);
or UO_4417 (O_4417,N_49555,N_49332);
nand UO_4418 (O_4418,N_47404,N_49846);
xnor UO_4419 (O_4419,N_49341,N_46252);
or UO_4420 (O_4420,N_47627,N_45412);
and UO_4421 (O_4421,N_45892,N_45415);
or UO_4422 (O_4422,N_46658,N_47307);
nor UO_4423 (O_4423,N_45848,N_46130);
or UO_4424 (O_4424,N_49210,N_47253);
xor UO_4425 (O_4425,N_48094,N_46542);
nor UO_4426 (O_4426,N_47287,N_47543);
nand UO_4427 (O_4427,N_48888,N_49899);
nor UO_4428 (O_4428,N_47910,N_47935);
nor UO_4429 (O_4429,N_45414,N_45756);
xnor UO_4430 (O_4430,N_46591,N_49918);
or UO_4431 (O_4431,N_48024,N_46255);
nand UO_4432 (O_4432,N_46689,N_47319);
and UO_4433 (O_4433,N_48149,N_47753);
nor UO_4434 (O_4434,N_46079,N_45309);
and UO_4435 (O_4435,N_46133,N_45378);
xnor UO_4436 (O_4436,N_48617,N_46598);
nor UO_4437 (O_4437,N_49590,N_45597);
nand UO_4438 (O_4438,N_46123,N_47920);
nor UO_4439 (O_4439,N_49599,N_46094);
nand UO_4440 (O_4440,N_45983,N_47250);
and UO_4441 (O_4441,N_48716,N_49541);
or UO_4442 (O_4442,N_49890,N_46644);
or UO_4443 (O_4443,N_46021,N_47812);
nor UO_4444 (O_4444,N_45340,N_48511);
and UO_4445 (O_4445,N_45700,N_47725);
nor UO_4446 (O_4446,N_48876,N_48544);
or UO_4447 (O_4447,N_47476,N_49692);
xor UO_4448 (O_4448,N_45716,N_46132);
nor UO_4449 (O_4449,N_49722,N_47573);
and UO_4450 (O_4450,N_45654,N_45843);
nand UO_4451 (O_4451,N_48367,N_48512);
or UO_4452 (O_4452,N_48258,N_48149);
nor UO_4453 (O_4453,N_45336,N_46619);
xnor UO_4454 (O_4454,N_49483,N_47226);
nor UO_4455 (O_4455,N_46538,N_49393);
nor UO_4456 (O_4456,N_49922,N_49506);
and UO_4457 (O_4457,N_47944,N_47193);
nand UO_4458 (O_4458,N_48673,N_47373);
nand UO_4459 (O_4459,N_49907,N_46417);
nor UO_4460 (O_4460,N_45747,N_47644);
or UO_4461 (O_4461,N_49592,N_46172);
nor UO_4462 (O_4462,N_49995,N_46193);
and UO_4463 (O_4463,N_49220,N_45732);
or UO_4464 (O_4464,N_47392,N_48419);
nand UO_4465 (O_4465,N_49080,N_46354);
nor UO_4466 (O_4466,N_47547,N_49911);
nand UO_4467 (O_4467,N_46939,N_46616);
nor UO_4468 (O_4468,N_48901,N_47419);
and UO_4469 (O_4469,N_48182,N_45196);
xor UO_4470 (O_4470,N_45439,N_49679);
nor UO_4471 (O_4471,N_46877,N_45369);
nand UO_4472 (O_4472,N_48927,N_46229);
xnor UO_4473 (O_4473,N_47575,N_49308);
or UO_4474 (O_4474,N_48310,N_49091);
nor UO_4475 (O_4475,N_48029,N_46091);
xor UO_4476 (O_4476,N_47984,N_47167);
or UO_4477 (O_4477,N_49979,N_49908);
xor UO_4478 (O_4478,N_47631,N_46052);
xnor UO_4479 (O_4479,N_46564,N_46545);
nor UO_4480 (O_4480,N_47181,N_45349);
xnor UO_4481 (O_4481,N_45143,N_46529);
or UO_4482 (O_4482,N_48234,N_47634);
or UO_4483 (O_4483,N_47690,N_45411);
xnor UO_4484 (O_4484,N_49115,N_48170);
xnor UO_4485 (O_4485,N_45596,N_48981);
and UO_4486 (O_4486,N_46007,N_46395);
and UO_4487 (O_4487,N_45474,N_47843);
nor UO_4488 (O_4488,N_48145,N_47229);
nand UO_4489 (O_4489,N_48615,N_46507);
and UO_4490 (O_4490,N_49579,N_45851);
and UO_4491 (O_4491,N_45220,N_45711);
nand UO_4492 (O_4492,N_49403,N_45948);
or UO_4493 (O_4493,N_46284,N_45901);
xnor UO_4494 (O_4494,N_46412,N_47109);
xnor UO_4495 (O_4495,N_49358,N_49598);
xnor UO_4496 (O_4496,N_46841,N_48734);
xor UO_4497 (O_4497,N_49627,N_49266);
nand UO_4498 (O_4498,N_49273,N_45133);
and UO_4499 (O_4499,N_48052,N_49122);
or UO_4500 (O_4500,N_48159,N_45248);
xor UO_4501 (O_4501,N_48213,N_49122);
xor UO_4502 (O_4502,N_46335,N_46465);
nor UO_4503 (O_4503,N_48444,N_46031);
and UO_4504 (O_4504,N_49577,N_49639);
nor UO_4505 (O_4505,N_47198,N_46969);
nor UO_4506 (O_4506,N_48431,N_48483);
nor UO_4507 (O_4507,N_45012,N_48176);
xnor UO_4508 (O_4508,N_45336,N_48767);
nor UO_4509 (O_4509,N_46059,N_45992);
xor UO_4510 (O_4510,N_47737,N_48741);
or UO_4511 (O_4511,N_45391,N_48664);
and UO_4512 (O_4512,N_47468,N_48939);
and UO_4513 (O_4513,N_49725,N_45452);
nand UO_4514 (O_4514,N_45609,N_46179);
or UO_4515 (O_4515,N_47408,N_47406);
and UO_4516 (O_4516,N_49312,N_47101);
nor UO_4517 (O_4517,N_46946,N_45804);
nand UO_4518 (O_4518,N_46045,N_49971);
or UO_4519 (O_4519,N_48992,N_47652);
or UO_4520 (O_4520,N_47799,N_49042);
and UO_4521 (O_4521,N_45999,N_46443);
nand UO_4522 (O_4522,N_48353,N_46501);
and UO_4523 (O_4523,N_46635,N_49865);
xor UO_4524 (O_4524,N_49885,N_45685);
xor UO_4525 (O_4525,N_49102,N_47825);
or UO_4526 (O_4526,N_46213,N_47000);
xnor UO_4527 (O_4527,N_49420,N_49653);
or UO_4528 (O_4528,N_47682,N_49477);
xor UO_4529 (O_4529,N_45311,N_45786);
xnor UO_4530 (O_4530,N_46000,N_46844);
and UO_4531 (O_4531,N_45117,N_45103);
or UO_4532 (O_4532,N_45422,N_49630);
and UO_4533 (O_4533,N_48493,N_45040);
and UO_4534 (O_4534,N_45803,N_48869);
or UO_4535 (O_4535,N_49703,N_46344);
xor UO_4536 (O_4536,N_45913,N_49331);
or UO_4537 (O_4537,N_45262,N_48709);
or UO_4538 (O_4538,N_48902,N_45815);
nand UO_4539 (O_4539,N_47259,N_47732);
xnor UO_4540 (O_4540,N_48460,N_47692);
or UO_4541 (O_4541,N_49843,N_45942);
xnor UO_4542 (O_4542,N_47755,N_47645);
nor UO_4543 (O_4543,N_47540,N_49768);
nand UO_4544 (O_4544,N_49608,N_46029);
nand UO_4545 (O_4545,N_45977,N_47502);
or UO_4546 (O_4546,N_46553,N_45274);
nand UO_4547 (O_4547,N_47789,N_49274);
nand UO_4548 (O_4548,N_47105,N_46522);
and UO_4549 (O_4549,N_45209,N_48908);
or UO_4550 (O_4550,N_47458,N_49503);
xor UO_4551 (O_4551,N_45275,N_47582);
or UO_4552 (O_4552,N_46242,N_47023);
xor UO_4553 (O_4553,N_49819,N_46365);
xnor UO_4554 (O_4554,N_47879,N_48506);
nand UO_4555 (O_4555,N_47413,N_46211);
and UO_4556 (O_4556,N_49222,N_45480);
and UO_4557 (O_4557,N_46041,N_47075);
and UO_4558 (O_4558,N_46075,N_46664);
nor UO_4559 (O_4559,N_46042,N_47968);
nor UO_4560 (O_4560,N_47701,N_48797);
and UO_4561 (O_4561,N_46738,N_48351);
nor UO_4562 (O_4562,N_49259,N_45028);
nand UO_4563 (O_4563,N_48677,N_45109);
xor UO_4564 (O_4564,N_49042,N_47276);
nand UO_4565 (O_4565,N_47183,N_46961);
nand UO_4566 (O_4566,N_45294,N_49444);
or UO_4567 (O_4567,N_46276,N_49654);
nand UO_4568 (O_4568,N_45262,N_48692);
xnor UO_4569 (O_4569,N_48159,N_49124);
xor UO_4570 (O_4570,N_46516,N_48136);
xnor UO_4571 (O_4571,N_46244,N_46078);
xor UO_4572 (O_4572,N_47564,N_46035);
and UO_4573 (O_4573,N_49713,N_49746);
or UO_4574 (O_4574,N_49075,N_45538);
and UO_4575 (O_4575,N_48962,N_45710);
nand UO_4576 (O_4576,N_45737,N_45922);
or UO_4577 (O_4577,N_48458,N_49483);
and UO_4578 (O_4578,N_47071,N_48247);
xor UO_4579 (O_4579,N_49863,N_45968);
nand UO_4580 (O_4580,N_49974,N_47963);
nor UO_4581 (O_4581,N_46359,N_46536);
or UO_4582 (O_4582,N_48299,N_47719);
and UO_4583 (O_4583,N_47369,N_48006);
nor UO_4584 (O_4584,N_48799,N_49257);
xnor UO_4585 (O_4585,N_45707,N_46514);
or UO_4586 (O_4586,N_46915,N_46611);
nor UO_4587 (O_4587,N_46202,N_46797);
nand UO_4588 (O_4588,N_49020,N_46589);
and UO_4589 (O_4589,N_46954,N_45333);
and UO_4590 (O_4590,N_45172,N_47069);
or UO_4591 (O_4591,N_46813,N_48309);
xnor UO_4592 (O_4592,N_49377,N_45897);
nor UO_4593 (O_4593,N_45802,N_46971);
nor UO_4594 (O_4594,N_48049,N_49383);
or UO_4595 (O_4595,N_46810,N_48046);
xor UO_4596 (O_4596,N_47755,N_47609);
and UO_4597 (O_4597,N_49215,N_46471);
nor UO_4598 (O_4598,N_46691,N_48659);
nor UO_4599 (O_4599,N_47769,N_47833);
nor UO_4600 (O_4600,N_49588,N_47427);
and UO_4601 (O_4601,N_47539,N_48602);
xor UO_4602 (O_4602,N_49536,N_45650);
nand UO_4603 (O_4603,N_47037,N_49633);
nor UO_4604 (O_4604,N_47164,N_49938);
or UO_4605 (O_4605,N_47521,N_45220);
or UO_4606 (O_4606,N_49892,N_46139);
and UO_4607 (O_4607,N_45071,N_49562);
nand UO_4608 (O_4608,N_47236,N_49159);
nand UO_4609 (O_4609,N_47247,N_45751);
and UO_4610 (O_4610,N_46889,N_47458);
nand UO_4611 (O_4611,N_49407,N_45286);
or UO_4612 (O_4612,N_46787,N_47566);
nand UO_4613 (O_4613,N_48624,N_45790);
nand UO_4614 (O_4614,N_49489,N_48597);
or UO_4615 (O_4615,N_46277,N_46462);
or UO_4616 (O_4616,N_47903,N_48735);
nor UO_4617 (O_4617,N_46210,N_46357);
and UO_4618 (O_4618,N_46168,N_45158);
nand UO_4619 (O_4619,N_45215,N_46205);
xnor UO_4620 (O_4620,N_46890,N_48929);
nor UO_4621 (O_4621,N_48921,N_47734);
or UO_4622 (O_4622,N_47971,N_48774);
nor UO_4623 (O_4623,N_49695,N_48040);
or UO_4624 (O_4624,N_49373,N_45893);
xnor UO_4625 (O_4625,N_47005,N_47954);
xnor UO_4626 (O_4626,N_45431,N_49246);
nor UO_4627 (O_4627,N_46617,N_46230);
or UO_4628 (O_4628,N_47198,N_46794);
nor UO_4629 (O_4629,N_46222,N_49192);
or UO_4630 (O_4630,N_49655,N_46653);
or UO_4631 (O_4631,N_47032,N_45930);
xor UO_4632 (O_4632,N_47516,N_47151);
and UO_4633 (O_4633,N_46993,N_48424);
nor UO_4634 (O_4634,N_47257,N_47366);
and UO_4635 (O_4635,N_46142,N_48885);
or UO_4636 (O_4636,N_49259,N_47570);
or UO_4637 (O_4637,N_48994,N_48114);
nand UO_4638 (O_4638,N_49513,N_49819);
and UO_4639 (O_4639,N_49796,N_46300);
nand UO_4640 (O_4640,N_46237,N_46896);
nand UO_4641 (O_4641,N_46577,N_47611);
and UO_4642 (O_4642,N_45899,N_49320);
and UO_4643 (O_4643,N_47168,N_49950);
or UO_4644 (O_4644,N_48757,N_48328);
nand UO_4645 (O_4645,N_48201,N_47320);
xor UO_4646 (O_4646,N_46676,N_46831);
xnor UO_4647 (O_4647,N_47624,N_47299);
xnor UO_4648 (O_4648,N_49940,N_47834);
or UO_4649 (O_4649,N_49398,N_45463);
xnor UO_4650 (O_4650,N_47114,N_46249);
xor UO_4651 (O_4651,N_48202,N_48876);
nand UO_4652 (O_4652,N_48646,N_48604);
or UO_4653 (O_4653,N_49806,N_49292);
xor UO_4654 (O_4654,N_49002,N_47060);
xnor UO_4655 (O_4655,N_48493,N_46080);
xor UO_4656 (O_4656,N_48797,N_48014);
nor UO_4657 (O_4657,N_45832,N_46111);
or UO_4658 (O_4658,N_49502,N_47831);
xor UO_4659 (O_4659,N_49977,N_48330);
xor UO_4660 (O_4660,N_47454,N_47452);
nand UO_4661 (O_4661,N_48850,N_45652);
or UO_4662 (O_4662,N_47095,N_46867);
nand UO_4663 (O_4663,N_46163,N_49739);
and UO_4664 (O_4664,N_48631,N_48514);
nor UO_4665 (O_4665,N_46432,N_47167);
xor UO_4666 (O_4666,N_45634,N_48858);
or UO_4667 (O_4667,N_49184,N_46705);
nor UO_4668 (O_4668,N_48660,N_47161);
or UO_4669 (O_4669,N_48796,N_45740);
nor UO_4670 (O_4670,N_45759,N_49933);
nand UO_4671 (O_4671,N_45399,N_48120);
or UO_4672 (O_4672,N_49402,N_47568);
nand UO_4673 (O_4673,N_49448,N_47656);
xor UO_4674 (O_4674,N_47174,N_49860);
nand UO_4675 (O_4675,N_49481,N_46817);
nand UO_4676 (O_4676,N_48779,N_47519);
nand UO_4677 (O_4677,N_45024,N_46431);
and UO_4678 (O_4678,N_46904,N_48475);
nand UO_4679 (O_4679,N_46279,N_49445);
or UO_4680 (O_4680,N_45502,N_47617);
xnor UO_4681 (O_4681,N_47160,N_49399);
nand UO_4682 (O_4682,N_45604,N_45625);
xnor UO_4683 (O_4683,N_46485,N_48313);
nand UO_4684 (O_4684,N_46025,N_49439);
nand UO_4685 (O_4685,N_45132,N_47334);
and UO_4686 (O_4686,N_49434,N_49569);
nand UO_4687 (O_4687,N_48711,N_48072);
xnor UO_4688 (O_4688,N_46782,N_47637);
nor UO_4689 (O_4689,N_48172,N_46011);
xnor UO_4690 (O_4690,N_49954,N_47377);
nor UO_4691 (O_4691,N_49420,N_49519);
nand UO_4692 (O_4692,N_47183,N_46496);
and UO_4693 (O_4693,N_46581,N_48354);
nand UO_4694 (O_4694,N_48396,N_46724);
and UO_4695 (O_4695,N_47301,N_47116);
nand UO_4696 (O_4696,N_45068,N_47467);
or UO_4697 (O_4697,N_47486,N_47862);
and UO_4698 (O_4698,N_46508,N_48376);
or UO_4699 (O_4699,N_48422,N_45271);
nand UO_4700 (O_4700,N_49274,N_49755);
xor UO_4701 (O_4701,N_48279,N_48261);
xor UO_4702 (O_4702,N_47313,N_46377);
xor UO_4703 (O_4703,N_48014,N_49250);
xor UO_4704 (O_4704,N_45411,N_47550);
and UO_4705 (O_4705,N_46434,N_48543);
xor UO_4706 (O_4706,N_48207,N_46292);
or UO_4707 (O_4707,N_46864,N_49875);
or UO_4708 (O_4708,N_45910,N_45625);
nand UO_4709 (O_4709,N_48861,N_48806);
xor UO_4710 (O_4710,N_47085,N_49670);
xor UO_4711 (O_4711,N_49896,N_49517);
or UO_4712 (O_4712,N_48627,N_46890);
nand UO_4713 (O_4713,N_47886,N_48190);
nand UO_4714 (O_4714,N_49452,N_45470);
and UO_4715 (O_4715,N_47539,N_47646);
xnor UO_4716 (O_4716,N_49202,N_47710);
nand UO_4717 (O_4717,N_47792,N_45861);
and UO_4718 (O_4718,N_49515,N_49536);
and UO_4719 (O_4719,N_45538,N_45968);
and UO_4720 (O_4720,N_49733,N_45483);
nor UO_4721 (O_4721,N_48149,N_46165);
and UO_4722 (O_4722,N_47513,N_48521);
xnor UO_4723 (O_4723,N_49025,N_45019);
and UO_4724 (O_4724,N_47585,N_49183);
nor UO_4725 (O_4725,N_46974,N_47371);
or UO_4726 (O_4726,N_48497,N_46617);
and UO_4727 (O_4727,N_45094,N_45731);
nor UO_4728 (O_4728,N_45740,N_46374);
nand UO_4729 (O_4729,N_45968,N_46888);
and UO_4730 (O_4730,N_48739,N_45706);
and UO_4731 (O_4731,N_45370,N_49356);
and UO_4732 (O_4732,N_45103,N_45844);
nor UO_4733 (O_4733,N_47440,N_46284);
and UO_4734 (O_4734,N_47765,N_46958);
nor UO_4735 (O_4735,N_47668,N_48494);
xor UO_4736 (O_4736,N_45994,N_49357);
and UO_4737 (O_4737,N_47698,N_49385);
nor UO_4738 (O_4738,N_45742,N_46035);
nor UO_4739 (O_4739,N_49295,N_47613);
and UO_4740 (O_4740,N_49423,N_49910);
and UO_4741 (O_4741,N_48195,N_47429);
xor UO_4742 (O_4742,N_45408,N_47022);
xor UO_4743 (O_4743,N_49722,N_46015);
nand UO_4744 (O_4744,N_47213,N_48721);
xor UO_4745 (O_4745,N_48547,N_48419);
and UO_4746 (O_4746,N_49138,N_46825);
xnor UO_4747 (O_4747,N_47940,N_46510);
or UO_4748 (O_4748,N_45343,N_46125);
or UO_4749 (O_4749,N_47707,N_45036);
nor UO_4750 (O_4750,N_49672,N_49398);
and UO_4751 (O_4751,N_47395,N_48762);
nor UO_4752 (O_4752,N_48583,N_46822);
nand UO_4753 (O_4753,N_47035,N_47197);
or UO_4754 (O_4754,N_47031,N_47230);
nand UO_4755 (O_4755,N_46313,N_48220);
and UO_4756 (O_4756,N_45661,N_49850);
and UO_4757 (O_4757,N_49631,N_46783);
nor UO_4758 (O_4758,N_47140,N_45361);
xor UO_4759 (O_4759,N_45074,N_46084);
and UO_4760 (O_4760,N_48358,N_45296);
or UO_4761 (O_4761,N_47479,N_45869);
xor UO_4762 (O_4762,N_49571,N_45174);
xnor UO_4763 (O_4763,N_47301,N_48472);
or UO_4764 (O_4764,N_45218,N_49223);
or UO_4765 (O_4765,N_48590,N_49560);
xnor UO_4766 (O_4766,N_46120,N_45782);
or UO_4767 (O_4767,N_46613,N_49429);
nand UO_4768 (O_4768,N_48891,N_48660);
nand UO_4769 (O_4769,N_46794,N_46139);
nor UO_4770 (O_4770,N_48931,N_46728);
or UO_4771 (O_4771,N_48748,N_48903);
xnor UO_4772 (O_4772,N_47003,N_46113);
or UO_4773 (O_4773,N_45912,N_46591);
xor UO_4774 (O_4774,N_49136,N_48117);
and UO_4775 (O_4775,N_49917,N_48099);
xnor UO_4776 (O_4776,N_47400,N_46522);
or UO_4777 (O_4777,N_48904,N_45152);
and UO_4778 (O_4778,N_45993,N_49520);
and UO_4779 (O_4779,N_46515,N_46395);
or UO_4780 (O_4780,N_47232,N_45950);
or UO_4781 (O_4781,N_48273,N_48841);
nand UO_4782 (O_4782,N_45650,N_47872);
xor UO_4783 (O_4783,N_45135,N_45651);
xnor UO_4784 (O_4784,N_48301,N_47851);
nor UO_4785 (O_4785,N_47490,N_47409);
xor UO_4786 (O_4786,N_49615,N_47263);
or UO_4787 (O_4787,N_48993,N_48193);
or UO_4788 (O_4788,N_46369,N_49065);
nand UO_4789 (O_4789,N_45832,N_47584);
nand UO_4790 (O_4790,N_47472,N_46592);
nand UO_4791 (O_4791,N_49868,N_48715);
xnor UO_4792 (O_4792,N_46120,N_46224);
or UO_4793 (O_4793,N_49961,N_47687);
xor UO_4794 (O_4794,N_45566,N_49396);
nor UO_4795 (O_4795,N_47270,N_49692);
nand UO_4796 (O_4796,N_48086,N_47027);
nand UO_4797 (O_4797,N_49312,N_46191);
and UO_4798 (O_4798,N_46017,N_45184);
nor UO_4799 (O_4799,N_46490,N_49895);
nor UO_4800 (O_4800,N_45271,N_48506);
or UO_4801 (O_4801,N_47822,N_49562);
and UO_4802 (O_4802,N_45649,N_49330);
nand UO_4803 (O_4803,N_46574,N_48022);
xor UO_4804 (O_4804,N_45451,N_48186);
xor UO_4805 (O_4805,N_48502,N_47167);
nand UO_4806 (O_4806,N_45810,N_47537);
nor UO_4807 (O_4807,N_46507,N_47931);
nor UO_4808 (O_4808,N_46234,N_48199);
and UO_4809 (O_4809,N_47573,N_48199);
xnor UO_4810 (O_4810,N_48115,N_49932);
and UO_4811 (O_4811,N_48516,N_48884);
and UO_4812 (O_4812,N_47482,N_49023);
and UO_4813 (O_4813,N_49260,N_49383);
nand UO_4814 (O_4814,N_49167,N_49554);
or UO_4815 (O_4815,N_45960,N_45254);
nand UO_4816 (O_4816,N_49944,N_49290);
or UO_4817 (O_4817,N_46532,N_47692);
xnor UO_4818 (O_4818,N_45577,N_45411);
nor UO_4819 (O_4819,N_48296,N_47354);
or UO_4820 (O_4820,N_49082,N_45183);
nor UO_4821 (O_4821,N_47472,N_48520);
or UO_4822 (O_4822,N_47686,N_45302);
and UO_4823 (O_4823,N_48433,N_49874);
or UO_4824 (O_4824,N_47178,N_46242);
nor UO_4825 (O_4825,N_47482,N_46082);
nor UO_4826 (O_4826,N_47309,N_47778);
or UO_4827 (O_4827,N_45142,N_49047);
nor UO_4828 (O_4828,N_49819,N_49667);
or UO_4829 (O_4829,N_49558,N_49503);
or UO_4830 (O_4830,N_45624,N_49850);
nor UO_4831 (O_4831,N_45252,N_48845);
xor UO_4832 (O_4832,N_49682,N_49108);
and UO_4833 (O_4833,N_45019,N_46252);
or UO_4834 (O_4834,N_49541,N_49927);
nand UO_4835 (O_4835,N_45445,N_45320);
nand UO_4836 (O_4836,N_45765,N_49061);
xnor UO_4837 (O_4837,N_45254,N_49321);
or UO_4838 (O_4838,N_45258,N_46632);
or UO_4839 (O_4839,N_46394,N_46308);
and UO_4840 (O_4840,N_48820,N_48485);
nand UO_4841 (O_4841,N_47957,N_49489);
and UO_4842 (O_4842,N_47781,N_46676);
or UO_4843 (O_4843,N_48591,N_48144);
xnor UO_4844 (O_4844,N_46538,N_48114);
xnor UO_4845 (O_4845,N_45216,N_48294);
or UO_4846 (O_4846,N_45108,N_47698);
nor UO_4847 (O_4847,N_46919,N_47581);
xor UO_4848 (O_4848,N_45747,N_45953);
xnor UO_4849 (O_4849,N_46880,N_48829);
or UO_4850 (O_4850,N_45171,N_46457);
xor UO_4851 (O_4851,N_45686,N_47882);
or UO_4852 (O_4852,N_45457,N_46303);
and UO_4853 (O_4853,N_47731,N_49599);
nand UO_4854 (O_4854,N_45429,N_47136);
xor UO_4855 (O_4855,N_48777,N_49825);
nor UO_4856 (O_4856,N_45006,N_47020);
xor UO_4857 (O_4857,N_48327,N_49802);
nor UO_4858 (O_4858,N_45234,N_48719);
xnor UO_4859 (O_4859,N_46751,N_49022);
nor UO_4860 (O_4860,N_45696,N_48437);
nor UO_4861 (O_4861,N_48801,N_47978);
nor UO_4862 (O_4862,N_48796,N_46898);
or UO_4863 (O_4863,N_48909,N_46611);
and UO_4864 (O_4864,N_47303,N_49261);
and UO_4865 (O_4865,N_46644,N_46533);
or UO_4866 (O_4866,N_45995,N_47592);
nand UO_4867 (O_4867,N_46263,N_49307);
nand UO_4868 (O_4868,N_47250,N_48264);
and UO_4869 (O_4869,N_45970,N_47525);
nor UO_4870 (O_4870,N_47961,N_47051);
xor UO_4871 (O_4871,N_46498,N_49613);
and UO_4872 (O_4872,N_45043,N_47644);
or UO_4873 (O_4873,N_45891,N_49504);
nor UO_4874 (O_4874,N_47775,N_47567);
nand UO_4875 (O_4875,N_49668,N_45198);
nor UO_4876 (O_4876,N_46571,N_48770);
nor UO_4877 (O_4877,N_46352,N_45690);
or UO_4878 (O_4878,N_48552,N_46844);
xnor UO_4879 (O_4879,N_49187,N_48568);
or UO_4880 (O_4880,N_49456,N_45781);
nor UO_4881 (O_4881,N_45334,N_48476);
xor UO_4882 (O_4882,N_47699,N_48134);
nor UO_4883 (O_4883,N_47602,N_49415);
or UO_4884 (O_4884,N_47275,N_46874);
xor UO_4885 (O_4885,N_45873,N_48074);
or UO_4886 (O_4886,N_49420,N_45018);
nor UO_4887 (O_4887,N_46564,N_49743);
nor UO_4888 (O_4888,N_48911,N_46105);
nor UO_4889 (O_4889,N_49270,N_47002);
nand UO_4890 (O_4890,N_46322,N_49769);
or UO_4891 (O_4891,N_47386,N_46225);
nor UO_4892 (O_4892,N_48812,N_49090);
and UO_4893 (O_4893,N_46506,N_49916);
or UO_4894 (O_4894,N_47873,N_46092);
xor UO_4895 (O_4895,N_47260,N_49698);
xor UO_4896 (O_4896,N_46411,N_47724);
and UO_4897 (O_4897,N_47572,N_46622);
or UO_4898 (O_4898,N_46937,N_49511);
nor UO_4899 (O_4899,N_47158,N_49657);
xnor UO_4900 (O_4900,N_49707,N_49036);
xor UO_4901 (O_4901,N_49212,N_48933);
xnor UO_4902 (O_4902,N_46502,N_47500);
and UO_4903 (O_4903,N_46769,N_45804);
nor UO_4904 (O_4904,N_46740,N_46088);
nand UO_4905 (O_4905,N_47541,N_48105);
or UO_4906 (O_4906,N_45460,N_47845);
nor UO_4907 (O_4907,N_48014,N_48865);
nor UO_4908 (O_4908,N_46955,N_48312);
and UO_4909 (O_4909,N_47291,N_45848);
xnor UO_4910 (O_4910,N_46996,N_45916);
nor UO_4911 (O_4911,N_49120,N_49638);
and UO_4912 (O_4912,N_46605,N_48184);
nand UO_4913 (O_4913,N_47254,N_45802);
and UO_4914 (O_4914,N_46988,N_49275);
or UO_4915 (O_4915,N_45695,N_48707);
and UO_4916 (O_4916,N_47902,N_48134);
and UO_4917 (O_4917,N_45178,N_48319);
xnor UO_4918 (O_4918,N_49234,N_48827);
nor UO_4919 (O_4919,N_49317,N_45153);
nor UO_4920 (O_4920,N_49086,N_46638);
and UO_4921 (O_4921,N_48734,N_49370);
nand UO_4922 (O_4922,N_47061,N_48064);
nand UO_4923 (O_4923,N_47553,N_49117);
nand UO_4924 (O_4924,N_45771,N_46873);
or UO_4925 (O_4925,N_46034,N_49671);
nand UO_4926 (O_4926,N_47355,N_46337);
nand UO_4927 (O_4927,N_45559,N_46712);
nor UO_4928 (O_4928,N_48300,N_48386);
and UO_4929 (O_4929,N_46536,N_48882);
or UO_4930 (O_4930,N_49853,N_46966);
xor UO_4931 (O_4931,N_46635,N_45053);
or UO_4932 (O_4932,N_49926,N_48284);
nand UO_4933 (O_4933,N_48593,N_45170);
and UO_4934 (O_4934,N_45874,N_45079);
nand UO_4935 (O_4935,N_45493,N_46448);
or UO_4936 (O_4936,N_49206,N_49168);
xnor UO_4937 (O_4937,N_49761,N_46278);
and UO_4938 (O_4938,N_47632,N_47612);
and UO_4939 (O_4939,N_48204,N_47409);
or UO_4940 (O_4940,N_48039,N_48473);
or UO_4941 (O_4941,N_46278,N_45927);
nand UO_4942 (O_4942,N_45718,N_45582);
xnor UO_4943 (O_4943,N_48826,N_45327);
nor UO_4944 (O_4944,N_47231,N_47436);
xnor UO_4945 (O_4945,N_47189,N_46207);
or UO_4946 (O_4946,N_49992,N_47197);
or UO_4947 (O_4947,N_49904,N_46504);
xor UO_4948 (O_4948,N_48120,N_48067);
nor UO_4949 (O_4949,N_45529,N_48969);
xnor UO_4950 (O_4950,N_49103,N_49106);
nor UO_4951 (O_4951,N_47629,N_47526);
xor UO_4952 (O_4952,N_48793,N_46188);
xor UO_4953 (O_4953,N_47257,N_48134);
and UO_4954 (O_4954,N_46240,N_45429);
xnor UO_4955 (O_4955,N_48455,N_48062);
and UO_4956 (O_4956,N_48779,N_49773);
and UO_4957 (O_4957,N_49368,N_45636);
nor UO_4958 (O_4958,N_48031,N_45287);
xnor UO_4959 (O_4959,N_45507,N_47889);
and UO_4960 (O_4960,N_46930,N_46024);
nand UO_4961 (O_4961,N_46135,N_47395);
and UO_4962 (O_4962,N_49007,N_49518);
xnor UO_4963 (O_4963,N_47773,N_49402);
and UO_4964 (O_4964,N_49617,N_45058);
or UO_4965 (O_4965,N_46206,N_49367);
and UO_4966 (O_4966,N_48330,N_49765);
or UO_4967 (O_4967,N_46431,N_45455);
and UO_4968 (O_4968,N_47186,N_45436);
nor UO_4969 (O_4969,N_49514,N_45437);
nor UO_4970 (O_4970,N_47686,N_46982);
nand UO_4971 (O_4971,N_45390,N_47724);
and UO_4972 (O_4972,N_45915,N_49746);
xor UO_4973 (O_4973,N_48784,N_48134);
xnor UO_4974 (O_4974,N_47244,N_45830);
nand UO_4975 (O_4975,N_46758,N_48600);
nor UO_4976 (O_4976,N_46096,N_45604);
xor UO_4977 (O_4977,N_49231,N_48083);
and UO_4978 (O_4978,N_46823,N_45132);
and UO_4979 (O_4979,N_45692,N_47305);
or UO_4980 (O_4980,N_45346,N_45837);
nor UO_4981 (O_4981,N_48234,N_46333);
or UO_4982 (O_4982,N_47757,N_46340);
or UO_4983 (O_4983,N_48142,N_48532);
and UO_4984 (O_4984,N_46236,N_48035);
and UO_4985 (O_4985,N_48998,N_48582);
nand UO_4986 (O_4986,N_48328,N_46774);
nand UO_4987 (O_4987,N_47918,N_45074);
or UO_4988 (O_4988,N_46448,N_47346);
and UO_4989 (O_4989,N_49208,N_49318);
nand UO_4990 (O_4990,N_47061,N_47636);
nor UO_4991 (O_4991,N_47598,N_47639);
or UO_4992 (O_4992,N_46029,N_46314);
nand UO_4993 (O_4993,N_47645,N_48675);
and UO_4994 (O_4994,N_49725,N_45495);
or UO_4995 (O_4995,N_47239,N_45084);
nand UO_4996 (O_4996,N_48437,N_48895);
nor UO_4997 (O_4997,N_45934,N_49984);
xor UO_4998 (O_4998,N_45382,N_46123);
nand UO_4999 (O_4999,N_47597,N_46131);
endmodule