module basic_1000_10000_1500_10_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_767,In_170);
or U1 (N_1,In_111,In_143);
and U2 (N_2,In_747,In_238);
and U3 (N_3,In_66,In_862);
and U4 (N_4,In_242,In_24);
and U5 (N_5,In_799,In_563);
nor U6 (N_6,In_17,In_813);
nor U7 (N_7,In_212,In_416);
nand U8 (N_8,In_524,In_785);
nor U9 (N_9,In_616,In_795);
nor U10 (N_10,In_678,In_570);
or U11 (N_11,In_84,In_966);
nor U12 (N_12,In_661,In_203);
nand U13 (N_13,In_939,In_816);
or U14 (N_14,In_147,In_422);
or U15 (N_15,In_546,In_145);
or U16 (N_16,In_204,In_451);
or U17 (N_17,In_362,In_133);
nor U18 (N_18,In_405,In_632);
or U19 (N_19,In_403,In_595);
nor U20 (N_20,In_149,In_964);
nand U21 (N_21,In_831,In_116);
nand U22 (N_22,In_664,In_509);
nor U23 (N_23,In_114,In_357);
nor U24 (N_24,In_499,In_274);
and U25 (N_25,In_902,In_513);
or U26 (N_26,In_586,In_764);
or U27 (N_27,In_339,In_373);
nor U28 (N_28,In_787,In_968);
or U29 (N_29,In_257,In_463);
or U30 (N_30,In_762,In_47);
and U31 (N_31,In_783,In_383);
or U32 (N_32,In_943,In_683);
and U33 (N_33,In_11,In_584);
or U34 (N_34,In_548,In_708);
nor U35 (N_35,In_697,In_140);
nand U36 (N_36,In_142,In_930);
nand U37 (N_37,In_67,In_520);
nand U38 (N_38,In_781,In_115);
or U39 (N_39,In_555,In_447);
and U40 (N_40,In_270,In_456);
nand U41 (N_41,In_231,In_453);
and U42 (N_42,In_603,In_209);
and U43 (N_43,In_316,In_495);
nor U44 (N_44,In_190,In_109);
nor U45 (N_45,In_228,In_27);
xnor U46 (N_46,In_809,In_164);
and U47 (N_47,In_892,In_248);
nand U48 (N_48,In_60,In_984);
nor U49 (N_49,In_71,In_359);
and U50 (N_50,In_467,In_155);
nor U51 (N_51,In_946,In_618);
nor U52 (N_52,In_569,In_861);
nor U53 (N_53,In_670,In_778);
and U54 (N_54,In_870,In_773);
or U55 (N_55,In_458,In_927);
nand U56 (N_56,In_737,In_374);
nor U57 (N_57,In_356,In_776);
and U58 (N_58,In_835,In_286);
or U59 (N_59,In_536,In_293);
or U60 (N_60,In_343,In_470);
and U61 (N_61,In_667,In_239);
or U62 (N_62,In_977,In_527);
and U63 (N_63,In_597,In_825);
nor U64 (N_64,In_541,In_904);
or U65 (N_65,In_972,In_175);
nand U66 (N_66,In_103,In_262);
or U67 (N_67,In_250,In_395);
nor U68 (N_68,In_188,In_77);
nand U69 (N_69,In_211,In_918);
and U70 (N_70,In_69,In_913);
and U71 (N_71,In_675,In_868);
xnor U72 (N_72,In_672,In_402);
nand U73 (N_73,In_642,In_766);
and U74 (N_74,In_874,In_397);
or U75 (N_75,In_622,In_582);
nor U76 (N_76,In_480,In_611);
or U77 (N_77,In_971,In_985);
and U78 (N_78,In_755,In_104);
or U79 (N_79,In_756,In_179);
nor U80 (N_80,In_804,In_987);
or U81 (N_81,In_596,In_759);
nor U82 (N_82,In_330,In_376);
nand U83 (N_83,In_612,In_245);
nand U84 (N_84,In_812,In_478);
or U85 (N_85,In_853,In_765);
nand U86 (N_86,In_699,In_976);
or U87 (N_87,In_78,In_566);
or U88 (N_88,In_425,In_464);
nand U89 (N_89,In_259,In_493);
nand U90 (N_90,In_620,In_284);
and U91 (N_91,In_910,In_556);
nand U92 (N_92,In_899,In_342);
or U93 (N_93,In_588,In_543);
or U94 (N_94,In_518,In_191);
nand U95 (N_95,In_154,In_430);
nand U96 (N_96,In_466,In_194);
or U97 (N_97,In_540,In_68);
and U98 (N_98,In_76,In_750);
and U99 (N_99,In_221,In_802);
nor U100 (N_100,In_95,In_647);
and U101 (N_101,In_235,In_629);
nor U102 (N_102,In_208,In_117);
or U103 (N_103,In_656,In_973);
nand U104 (N_104,In_936,In_347);
nand U105 (N_105,In_681,In_217);
nand U106 (N_106,In_137,In_229);
and U107 (N_107,In_55,In_720);
or U108 (N_108,In_653,In_233);
or U109 (N_109,In_858,In_948);
or U110 (N_110,In_991,In_791);
nand U111 (N_111,In_637,In_933);
or U112 (N_112,In_352,In_907);
or U113 (N_113,In_298,In_167);
or U114 (N_114,In_153,In_805);
nor U115 (N_115,In_282,In_743);
or U116 (N_116,In_871,In_303);
nand U117 (N_117,In_657,In_215);
or U118 (N_118,In_334,In_200);
and U119 (N_119,In_21,In_23);
nand U120 (N_120,In_702,In_389);
and U121 (N_121,In_626,In_161);
nor U122 (N_122,In_901,In_539);
nor U123 (N_123,In_733,In_407);
or U124 (N_124,In_729,In_431);
and U125 (N_125,In_885,In_59);
nand U126 (N_126,In_947,In_85);
or U127 (N_127,In_158,In_57);
nand U128 (N_128,In_4,In_598);
nand U129 (N_129,In_741,In_655);
nor U130 (N_130,In_36,In_953);
nor U131 (N_131,In_591,In_328);
nand U132 (N_132,In_682,In_829);
xnor U133 (N_133,In_950,In_314);
or U134 (N_134,In_843,In_940);
nand U135 (N_135,In_94,In_487);
nor U136 (N_136,In_138,In_954);
and U137 (N_137,In_344,In_684);
or U138 (N_138,In_609,In_817);
or U139 (N_139,In_834,In_435);
and U140 (N_140,In_818,In_875);
and U141 (N_141,In_864,In_39);
nor U142 (N_142,In_792,In_491);
nor U143 (N_143,In_724,In_760);
or U144 (N_144,In_833,In_232);
nand U145 (N_145,In_725,In_998);
or U146 (N_146,In_20,In_735);
nand U147 (N_147,In_510,In_605);
and U148 (N_148,In_247,In_320);
nor U149 (N_149,In_5,In_291);
nor U150 (N_150,In_769,In_234);
or U151 (N_151,In_960,In_763);
nand U152 (N_152,In_341,In_227);
or U153 (N_153,In_925,In_294);
or U154 (N_154,In_528,In_450);
nor U155 (N_155,In_457,In_704);
or U156 (N_156,In_723,In_124);
nand U157 (N_157,In_183,In_44);
and U158 (N_158,In_160,In_614);
nor U159 (N_159,In_580,In_434);
or U160 (N_160,In_654,In_492);
nor U161 (N_161,In_599,In_700);
and U162 (N_162,In_623,In_346);
nor U163 (N_163,In_338,In_471);
nand U164 (N_164,In_989,In_884);
nor U165 (N_165,In_426,In_919);
nor U166 (N_166,In_610,In_449);
and U167 (N_167,In_419,In_577);
and U168 (N_168,In_676,In_353);
nor U169 (N_169,In_857,In_354);
or U170 (N_170,In_842,In_433);
or U171 (N_171,In_553,In_301);
nand U172 (N_172,In_881,In_942);
nor U173 (N_173,In_648,In_852);
nor U174 (N_174,In_443,In_886);
nand U175 (N_175,In_323,In_43);
or U176 (N_176,In_639,In_916);
nor U177 (N_177,In_460,In_367);
nand U178 (N_178,In_996,In_61);
and U179 (N_179,In_830,In_391);
or U180 (N_180,In_736,In_406);
nand U181 (N_181,In_928,In_428);
nor U182 (N_182,In_392,In_150);
nor U183 (N_183,In_779,In_172);
nor U184 (N_184,In_8,In_538);
nor U185 (N_185,In_982,In_462);
nand U186 (N_186,In_784,In_823);
nor U187 (N_187,In_519,In_967);
or U188 (N_188,In_978,In_269);
or U189 (N_189,In_777,In_472);
or U190 (N_190,In_437,In_613);
nor U191 (N_191,In_937,In_573);
nor U192 (N_192,In_366,In_220);
or U193 (N_193,In_712,In_315);
and U194 (N_194,In_171,In_912);
or U195 (N_195,In_63,In_876);
nand U196 (N_196,In_398,In_93);
nand U197 (N_197,In_692,In_299);
or U198 (N_198,In_267,In_788);
and U199 (N_199,In_707,In_680);
and U200 (N_200,In_485,In_836);
and U201 (N_201,In_333,In_459);
nor U202 (N_202,In_638,In_979);
nand U203 (N_203,In_6,In_304);
nor U204 (N_204,In_424,In_163);
nand U205 (N_205,In_689,In_839);
nand U206 (N_206,In_174,In_411);
nand U207 (N_207,In_926,In_896);
and U208 (N_208,In_752,In_13);
and U209 (N_209,In_14,In_698);
nand U210 (N_210,In_650,In_748);
xnor U211 (N_211,In_106,In_845);
nand U212 (N_212,In_285,In_202);
nor U213 (N_213,In_721,In_130);
and U214 (N_214,In_1,In_29);
nand U215 (N_215,In_815,In_685);
nor U216 (N_216,In_530,In_131);
and U217 (N_217,In_914,In_311);
nand U218 (N_218,In_761,In_955);
nor U219 (N_219,In_423,In_123);
or U220 (N_220,In_551,In_641);
nand U221 (N_221,In_414,In_542);
nor U222 (N_222,In_758,In_112);
nand U223 (N_223,In_474,In_452);
nor U224 (N_224,In_941,In_797);
or U225 (N_225,In_869,In_903);
and U226 (N_226,In_554,In_264);
xnor U227 (N_227,In_590,In_826);
nand U228 (N_228,In_992,In_585);
nor U229 (N_229,In_266,In_283);
xnor U230 (N_230,In_32,In_969);
nor U231 (N_231,In_477,In_52);
and U232 (N_232,In_935,In_281);
nand U233 (N_233,In_693,In_952);
nor U234 (N_234,In_562,In_889);
nor U235 (N_235,In_574,In_120);
nand U236 (N_236,In_306,In_921);
nor U237 (N_237,In_90,In_900);
or U238 (N_238,In_498,In_793);
and U239 (N_239,In_325,In_465);
nand U240 (N_240,In_73,In_807);
or U241 (N_241,In_128,In_951);
or U242 (N_242,In_475,In_532);
or U243 (N_243,In_81,In_385);
or U244 (N_244,In_75,In_295);
nand U245 (N_245,In_859,In_631);
nor U246 (N_246,In_418,In_380);
or U247 (N_247,In_62,In_489);
nor U248 (N_248,In_803,In_922);
and U249 (N_249,In_348,In_317);
nand U250 (N_250,In_565,In_658);
nand U251 (N_251,In_694,In_571);
or U252 (N_252,In_253,In_265);
nor U253 (N_253,In_810,In_696);
and U254 (N_254,In_48,In_560);
and U255 (N_255,In_272,In_624);
nand U256 (N_256,In_177,In_230);
or U257 (N_257,In_91,In_82);
and U258 (N_258,In_728,In_401);
and U259 (N_259,In_218,In_408);
nand U260 (N_260,In_387,In_3);
nand U261 (N_261,In_768,In_866);
or U262 (N_262,In_994,In_999);
or U263 (N_263,In_965,In_959);
nand U264 (N_264,In_302,In_744);
and U265 (N_265,In_51,In_181);
or U266 (N_266,In_162,In_193);
and U267 (N_267,In_278,In_438);
or U268 (N_268,In_975,In_717);
and U269 (N_269,In_319,In_80);
nor U270 (N_270,In_931,In_890);
nand U271 (N_271,In_848,In_860);
nor U272 (N_272,In_640,In_219);
or U273 (N_273,In_600,In_129);
and U274 (N_274,In_687,In_545);
nor U275 (N_275,In_820,In_96);
or U276 (N_276,In_275,In_932);
nor U277 (N_277,In_7,In_558);
and U278 (N_278,In_832,In_236);
or U279 (N_279,In_970,In_714);
nor U280 (N_280,In_87,In_50);
nand U281 (N_281,In_962,In_898);
nand U282 (N_282,In_742,In_608);
nor U283 (N_283,In_659,In_386);
nand U284 (N_284,In_119,In_308);
nand U285 (N_285,In_572,In_872);
nand U286 (N_286,In_615,In_806);
nand U287 (N_287,In_351,In_427);
xor U288 (N_288,In_621,In_350);
nand U289 (N_289,In_691,In_363);
nand U290 (N_290,In_86,In_243);
xor U291 (N_291,In_65,In_814);
nor U292 (N_292,In_30,In_327);
nor U293 (N_293,In_924,In_404);
nor U294 (N_294,In_677,In_176);
or U295 (N_295,In_448,In_732);
or U296 (N_296,In_100,In_393);
nor U297 (N_297,In_645,In_808);
nor U298 (N_298,In_186,In_662);
or U299 (N_299,In_440,In_709);
nor U300 (N_300,In_101,In_533);
nand U301 (N_301,In_811,In_607);
nand U302 (N_302,In_372,In_309);
and U303 (N_303,In_54,In_557);
nand U304 (N_304,In_148,In_390);
nor U305 (N_305,In_455,In_476);
and U306 (N_306,In_649,In_535);
and U307 (N_307,In_906,In_934);
or U308 (N_308,In_944,In_517);
and U309 (N_309,In_226,In_774);
and U310 (N_310,In_706,In_751);
nor U311 (N_311,In_534,In_679);
nand U312 (N_312,In_122,In_719);
and U313 (N_313,In_297,In_507);
or U314 (N_314,In_625,In_838);
nand U315 (N_315,In_144,In_289);
or U316 (N_316,In_216,In_695);
and U317 (N_317,In_141,In_963);
nor U318 (N_318,In_192,In_500);
or U319 (N_319,In_856,In_337);
or U320 (N_320,In_444,In_324);
and U321 (N_321,In_974,In_439);
nor U322 (N_322,In_713,In_486);
xnor U323 (N_323,In_636,In_56);
nand U324 (N_324,In_801,In_31);
or U325 (N_325,In_410,In_606);
or U326 (N_326,In_375,In_671);
and U327 (N_327,In_980,In_617);
or U328 (N_328,In_552,In_846);
nand U329 (N_329,In_479,In_360);
nand U330 (N_330,In_197,In_469);
and U331 (N_331,In_521,In_627);
and U332 (N_332,In_877,In_644);
nand U333 (N_333,In_537,In_296);
nand U334 (N_334,In_506,In_79);
or U335 (N_335,In_318,In_993);
and U336 (N_336,In_515,In_578);
xor U337 (N_337,In_646,In_201);
nor U338 (N_338,In_290,In_490);
nand U339 (N_339,In_261,In_74);
or U340 (N_340,In_746,In_997);
or U341 (N_341,In_102,In_849);
or U342 (N_342,In_446,In_41);
nor U343 (N_343,In_2,In_166);
nand U344 (N_344,In_911,In_409);
and U345 (N_345,In_173,In_757);
and U346 (N_346,In_878,In_824);
nand U347 (N_347,In_895,In_731);
nor U348 (N_348,In_529,In_722);
nor U349 (N_349,In_847,In_504);
nor U350 (N_350,In_432,In_628);
nor U351 (N_351,In_961,In_800);
or U352 (N_352,In_798,In_589);
or U353 (N_353,In_442,In_454);
or U354 (N_354,In_165,In_593);
or U355 (N_355,In_156,In_771);
nand U356 (N_356,In_42,In_958);
or U357 (N_357,In_983,In_920);
nand U358 (N_358,In_753,In_651);
nand U359 (N_359,In_503,In_635);
or U360 (N_360,In_822,In_688);
or U361 (N_361,In_381,In_894);
or U362 (N_362,In_483,In_118);
or U363 (N_363,In_279,In_770);
nor U364 (N_364,In_841,In_726);
or U365 (N_365,In_224,In_643);
nor U366 (N_366,In_300,In_844);
nand U367 (N_367,In_429,In_206);
nand U368 (N_368,In_923,In_880);
nor U369 (N_369,In_497,In_157);
and U370 (N_370,In_738,In_796);
nand U371 (N_371,In_18,In_837);
and U372 (N_372,In_310,In_196);
or U373 (N_373,In_718,In_957);
nand U374 (N_374,In_33,In_34);
nor U375 (N_375,In_601,In_15);
or U376 (N_376,In_98,In_855);
xnor U377 (N_377,In_252,In_255);
nand U378 (N_378,In_413,In_369);
or U379 (N_379,In_134,In_995);
nor U380 (N_380,In_187,In_564);
and U381 (N_381,In_136,In_16);
nor U382 (N_382,In_775,In_180);
or U383 (N_383,In_749,In_97);
or U384 (N_384,In_633,In_305);
nand U385 (N_385,In_468,In_436);
or U386 (N_386,In_547,In_909);
and U387 (N_387,In_505,In_139);
nand U388 (N_388,In_790,In_258);
nor U389 (N_389,In_592,In_888);
nand U390 (N_390,In_496,In_905);
nor U391 (N_391,In_365,In_113);
and U392 (N_392,In_125,In_9);
nand U393 (N_393,In_127,In_384);
nand U394 (N_394,In_669,In_727);
nor U395 (N_395,In_739,In_169);
nor U396 (N_396,In_579,In_508);
or U397 (N_397,In_45,In_168);
or U398 (N_398,In_531,In_581);
and U399 (N_399,In_195,In_867);
nand U400 (N_400,In_72,In_135);
or U401 (N_401,In_371,In_287);
nand U402 (N_402,In_364,In_850);
or U403 (N_403,In_663,In_151);
nor U404 (N_404,In_604,In_38);
nor U405 (N_405,In_312,In_666);
or U406 (N_406,In_28,In_559);
or U407 (N_407,In_891,In_249);
nor U408 (N_408,In_225,In_701);
and U409 (N_409,In_544,In_335);
or U410 (N_410,In_893,In_522);
nand U411 (N_411,In_786,In_981);
nor U412 (N_412,In_879,In_64);
nor U413 (N_413,In_561,In_481);
and U414 (N_414,In_821,In_88);
nor U415 (N_415,In_210,In_715);
nor U416 (N_416,In_273,In_441);
nor U417 (N_417,In_819,In_378);
nor U418 (N_418,In_349,In_782);
and U419 (N_419,In_205,In_263);
or U420 (N_420,In_594,In_986);
nor U421 (N_421,In_126,In_58);
nand U422 (N_422,In_794,In_35);
or U423 (N_423,In_494,In_370);
and U424 (N_424,In_332,In_198);
nand U425 (N_425,In_827,In_105);
and U426 (N_426,In_619,In_673);
nand U427 (N_427,In_549,In_251);
and U428 (N_428,In_634,In_237);
and U429 (N_429,In_244,In_587);
nor U430 (N_430,In_240,In_887);
nor U431 (N_431,In_89,In_184);
and U432 (N_432,In_883,In_576);
nand U433 (N_433,In_182,In_83);
and U434 (N_434,In_568,In_882);
nand U435 (N_435,In_990,In_525);
or U436 (N_436,In_417,In_711);
nand U437 (N_437,In_630,In_789);
or U438 (N_438,In_575,In_851);
nor U439 (N_439,In_754,In_512);
or U440 (N_440,In_665,In_214);
nor U441 (N_441,In_660,In_567);
nand U442 (N_442,In_189,In_377);
and U443 (N_443,In_132,In_674);
nor U444 (N_444,In_268,In_917);
nand U445 (N_445,In_780,In_396);
and U446 (N_446,In_358,In_92);
nand U447 (N_447,In_690,In_99);
or U448 (N_448,In_863,In_828);
nand U449 (N_449,In_178,In_482);
or U450 (N_450,In_772,In_12);
and U451 (N_451,In_716,In_705);
nand U452 (N_452,In_915,In_945);
nand U453 (N_453,In_415,In_445);
nand U454 (N_454,In_288,In_361);
or U455 (N_455,In_400,In_207);
or U456 (N_456,In_355,In_313);
and U457 (N_457,In_345,In_271);
nor U458 (N_458,In_421,In_213);
nor U459 (N_459,In_260,In_46);
and U460 (N_460,In_668,In_908);
nand U461 (N_461,In_340,In_514);
and U462 (N_462,In_107,In_246);
and U463 (N_463,In_473,In_159);
nand U464 (N_464,In_152,In_897);
xor U465 (N_465,In_929,In_10);
and U466 (N_466,In_526,In_292);
and U467 (N_467,In_256,In_110);
nor U468 (N_468,In_0,In_516);
nor U469 (N_469,In_70,In_730);
nand U470 (N_470,In_501,In_956);
or U471 (N_471,In_710,In_22);
and U472 (N_472,In_988,In_502);
or U473 (N_473,In_379,In_840);
nor U474 (N_474,In_523,In_949);
and U475 (N_475,In_331,In_461);
nand U476 (N_476,In_703,In_329);
nand U477 (N_477,In_399,In_185);
and U478 (N_478,In_873,In_25);
nor U479 (N_479,In_108,In_488);
nand U480 (N_480,In_412,In_652);
or U481 (N_481,In_550,In_734);
and U482 (N_482,In_280,In_321);
and U483 (N_483,In_484,In_336);
nor U484 (N_484,In_394,In_37);
or U485 (N_485,In_254,In_740);
or U486 (N_486,In_602,In_511);
or U487 (N_487,In_199,In_854);
and U488 (N_488,In_277,In_322);
and U489 (N_489,In_222,In_53);
nand U490 (N_490,In_146,In_223);
or U491 (N_491,In_938,In_745);
nor U492 (N_492,In_326,In_583);
and U493 (N_493,In_19,In_865);
nor U494 (N_494,In_241,In_382);
nor U495 (N_495,In_40,In_276);
and U496 (N_496,In_388,In_307);
nor U497 (N_497,In_121,In_49);
or U498 (N_498,In_686,In_26);
and U499 (N_499,In_420,In_368);
and U500 (N_500,In_634,In_583);
or U501 (N_501,In_232,In_839);
and U502 (N_502,In_29,In_477);
or U503 (N_503,In_957,In_426);
or U504 (N_504,In_247,In_638);
and U505 (N_505,In_587,In_271);
nor U506 (N_506,In_238,In_653);
nand U507 (N_507,In_340,In_461);
or U508 (N_508,In_816,In_678);
nand U509 (N_509,In_652,In_555);
or U510 (N_510,In_637,In_403);
or U511 (N_511,In_372,In_563);
nand U512 (N_512,In_706,In_540);
and U513 (N_513,In_977,In_447);
or U514 (N_514,In_238,In_525);
nand U515 (N_515,In_201,In_276);
nor U516 (N_516,In_91,In_71);
nor U517 (N_517,In_953,In_363);
and U518 (N_518,In_353,In_673);
nor U519 (N_519,In_967,In_922);
and U520 (N_520,In_459,In_473);
nor U521 (N_521,In_721,In_914);
or U522 (N_522,In_136,In_188);
nor U523 (N_523,In_814,In_446);
or U524 (N_524,In_992,In_833);
nand U525 (N_525,In_551,In_380);
and U526 (N_526,In_742,In_202);
nor U527 (N_527,In_903,In_410);
or U528 (N_528,In_664,In_953);
or U529 (N_529,In_943,In_759);
and U530 (N_530,In_503,In_127);
or U531 (N_531,In_53,In_708);
nand U532 (N_532,In_104,In_943);
or U533 (N_533,In_227,In_683);
and U534 (N_534,In_851,In_713);
nand U535 (N_535,In_191,In_512);
or U536 (N_536,In_34,In_922);
nand U537 (N_537,In_920,In_862);
or U538 (N_538,In_736,In_654);
nor U539 (N_539,In_645,In_562);
nand U540 (N_540,In_560,In_998);
nand U541 (N_541,In_421,In_324);
nor U542 (N_542,In_553,In_338);
nor U543 (N_543,In_452,In_421);
nand U544 (N_544,In_285,In_515);
nor U545 (N_545,In_967,In_384);
nand U546 (N_546,In_499,In_106);
and U547 (N_547,In_697,In_67);
nand U548 (N_548,In_383,In_941);
nand U549 (N_549,In_230,In_911);
and U550 (N_550,In_895,In_353);
nand U551 (N_551,In_401,In_770);
and U552 (N_552,In_556,In_963);
or U553 (N_553,In_208,In_602);
or U554 (N_554,In_623,In_394);
or U555 (N_555,In_359,In_979);
nand U556 (N_556,In_5,In_448);
nor U557 (N_557,In_648,In_392);
nand U558 (N_558,In_582,In_966);
nor U559 (N_559,In_454,In_300);
and U560 (N_560,In_219,In_954);
or U561 (N_561,In_29,In_96);
nor U562 (N_562,In_205,In_909);
or U563 (N_563,In_794,In_178);
and U564 (N_564,In_724,In_694);
and U565 (N_565,In_664,In_663);
nor U566 (N_566,In_694,In_506);
or U567 (N_567,In_797,In_469);
nand U568 (N_568,In_389,In_955);
or U569 (N_569,In_759,In_121);
or U570 (N_570,In_694,In_400);
nand U571 (N_571,In_518,In_864);
nor U572 (N_572,In_968,In_538);
or U573 (N_573,In_586,In_663);
and U574 (N_574,In_382,In_970);
and U575 (N_575,In_56,In_741);
or U576 (N_576,In_428,In_660);
nand U577 (N_577,In_679,In_574);
nand U578 (N_578,In_757,In_480);
and U579 (N_579,In_570,In_328);
nor U580 (N_580,In_55,In_93);
or U581 (N_581,In_245,In_483);
nand U582 (N_582,In_649,In_230);
and U583 (N_583,In_980,In_175);
or U584 (N_584,In_891,In_753);
nor U585 (N_585,In_409,In_539);
nand U586 (N_586,In_45,In_360);
and U587 (N_587,In_597,In_43);
nor U588 (N_588,In_618,In_328);
nand U589 (N_589,In_710,In_856);
nand U590 (N_590,In_540,In_557);
nand U591 (N_591,In_175,In_644);
nor U592 (N_592,In_874,In_318);
nand U593 (N_593,In_489,In_156);
or U594 (N_594,In_999,In_822);
and U595 (N_595,In_952,In_694);
or U596 (N_596,In_280,In_629);
xor U597 (N_597,In_523,In_77);
nand U598 (N_598,In_808,In_334);
or U599 (N_599,In_958,In_284);
nor U600 (N_600,In_596,In_538);
nor U601 (N_601,In_716,In_33);
nand U602 (N_602,In_767,In_798);
nor U603 (N_603,In_159,In_485);
or U604 (N_604,In_379,In_720);
nor U605 (N_605,In_309,In_434);
and U606 (N_606,In_637,In_467);
nand U607 (N_607,In_98,In_15);
nand U608 (N_608,In_567,In_382);
nor U609 (N_609,In_485,In_83);
nor U610 (N_610,In_950,In_129);
or U611 (N_611,In_182,In_377);
and U612 (N_612,In_961,In_307);
nor U613 (N_613,In_902,In_944);
or U614 (N_614,In_309,In_769);
nand U615 (N_615,In_148,In_712);
nand U616 (N_616,In_103,In_246);
or U617 (N_617,In_337,In_410);
and U618 (N_618,In_832,In_47);
nor U619 (N_619,In_943,In_232);
nor U620 (N_620,In_498,In_706);
nor U621 (N_621,In_300,In_104);
and U622 (N_622,In_323,In_421);
nand U623 (N_623,In_426,In_386);
nand U624 (N_624,In_11,In_34);
nor U625 (N_625,In_72,In_292);
nor U626 (N_626,In_337,In_345);
nand U627 (N_627,In_944,In_314);
nand U628 (N_628,In_195,In_920);
nor U629 (N_629,In_320,In_805);
nand U630 (N_630,In_630,In_584);
and U631 (N_631,In_31,In_604);
and U632 (N_632,In_780,In_90);
or U633 (N_633,In_547,In_899);
and U634 (N_634,In_391,In_490);
or U635 (N_635,In_10,In_736);
and U636 (N_636,In_311,In_751);
nand U637 (N_637,In_859,In_863);
or U638 (N_638,In_829,In_307);
or U639 (N_639,In_606,In_101);
or U640 (N_640,In_785,In_142);
and U641 (N_641,In_911,In_269);
nand U642 (N_642,In_187,In_317);
nand U643 (N_643,In_876,In_921);
and U644 (N_644,In_223,In_842);
nor U645 (N_645,In_883,In_302);
or U646 (N_646,In_983,In_953);
or U647 (N_647,In_109,In_980);
or U648 (N_648,In_899,In_969);
and U649 (N_649,In_951,In_407);
and U650 (N_650,In_79,In_335);
nand U651 (N_651,In_330,In_995);
nand U652 (N_652,In_946,In_227);
nand U653 (N_653,In_529,In_995);
and U654 (N_654,In_85,In_666);
or U655 (N_655,In_887,In_792);
or U656 (N_656,In_55,In_262);
and U657 (N_657,In_563,In_223);
or U658 (N_658,In_468,In_68);
nor U659 (N_659,In_171,In_54);
nand U660 (N_660,In_282,In_440);
nor U661 (N_661,In_956,In_308);
nor U662 (N_662,In_104,In_516);
nand U663 (N_663,In_858,In_445);
and U664 (N_664,In_606,In_165);
and U665 (N_665,In_315,In_640);
nand U666 (N_666,In_108,In_180);
and U667 (N_667,In_708,In_116);
nand U668 (N_668,In_27,In_402);
and U669 (N_669,In_251,In_611);
nor U670 (N_670,In_609,In_152);
nand U671 (N_671,In_859,In_451);
nand U672 (N_672,In_130,In_862);
nor U673 (N_673,In_3,In_431);
xor U674 (N_674,In_511,In_355);
or U675 (N_675,In_260,In_75);
nand U676 (N_676,In_86,In_235);
nor U677 (N_677,In_531,In_889);
and U678 (N_678,In_788,In_423);
or U679 (N_679,In_897,In_424);
nand U680 (N_680,In_592,In_340);
nand U681 (N_681,In_248,In_977);
and U682 (N_682,In_913,In_852);
nor U683 (N_683,In_68,In_639);
nand U684 (N_684,In_707,In_163);
nand U685 (N_685,In_477,In_779);
or U686 (N_686,In_296,In_522);
and U687 (N_687,In_193,In_510);
or U688 (N_688,In_142,In_344);
and U689 (N_689,In_769,In_478);
nand U690 (N_690,In_373,In_557);
or U691 (N_691,In_537,In_131);
nor U692 (N_692,In_669,In_93);
and U693 (N_693,In_878,In_462);
and U694 (N_694,In_338,In_557);
and U695 (N_695,In_644,In_688);
or U696 (N_696,In_485,In_317);
and U697 (N_697,In_743,In_906);
nor U698 (N_698,In_167,In_559);
and U699 (N_699,In_116,In_323);
nand U700 (N_700,In_354,In_93);
or U701 (N_701,In_62,In_284);
nor U702 (N_702,In_953,In_154);
or U703 (N_703,In_570,In_333);
and U704 (N_704,In_836,In_852);
and U705 (N_705,In_304,In_657);
and U706 (N_706,In_208,In_840);
nor U707 (N_707,In_430,In_467);
nand U708 (N_708,In_84,In_696);
nand U709 (N_709,In_936,In_463);
nand U710 (N_710,In_941,In_555);
or U711 (N_711,In_454,In_725);
nand U712 (N_712,In_533,In_238);
and U713 (N_713,In_376,In_451);
nand U714 (N_714,In_751,In_580);
or U715 (N_715,In_383,In_513);
or U716 (N_716,In_617,In_645);
nor U717 (N_717,In_144,In_501);
xnor U718 (N_718,In_831,In_22);
and U719 (N_719,In_258,In_788);
nor U720 (N_720,In_848,In_86);
nand U721 (N_721,In_956,In_605);
nand U722 (N_722,In_591,In_876);
nor U723 (N_723,In_440,In_670);
and U724 (N_724,In_434,In_57);
nand U725 (N_725,In_305,In_538);
nor U726 (N_726,In_885,In_950);
nor U727 (N_727,In_207,In_276);
and U728 (N_728,In_933,In_222);
nor U729 (N_729,In_440,In_224);
and U730 (N_730,In_982,In_681);
or U731 (N_731,In_517,In_98);
and U732 (N_732,In_357,In_220);
nor U733 (N_733,In_711,In_114);
nand U734 (N_734,In_886,In_544);
and U735 (N_735,In_771,In_297);
nor U736 (N_736,In_849,In_827);
and U737 (N_737,In_243,In_869);
or U738 (N_738,In_678,In_209);
and U739 (N_739,In_450,In_799);
nor U740 (N_740,In_3,In_149);
nand U741 (N_741,In_403,In_506);
or U742 (N_742,In_494,In_375);
or U743 (N_743,In_535,In_580);
xnor U744 (N_744,In_726,In_262);
and U745 (N_745,In_774,In_579);
and U746 (N_746,In_5,In_724);
and U747 (N_747,In_467,In_432);
nand U748 (N_748,In_385,In_959);
nand U749 (N_749,In_215,In_249);
or U750 (N_750,In_878,In_690);
and U751 (N_751,In_365,In_224);
or U752 (N_752,In_210,In_875);
nand U753 (N_753,In_592,In_232);
or U754 (N_754,In_715,In_579);
or U755 (N_755,In_561,In_962);
nand U756 (N_756,In_947,In_16);
and U757 (N_757,In_983,In_127);
and U758 (N_758,In_603,In_880);
or U759 (N_759,In_699,In_285);
xor U760 (N_760,In_815,In_401);
or U761 (N_761,In_909,In_362);
nand U762 (N_762,In_780,In_543);
nor U763 (N_763,In_373,In_351);
or U764 (N_764,In_488,In_999);
nor U765 (N_765,In_973,In_362);
nor U766 (N_766,In_220,In_212);
or U767 (N_767,In_397,In_504);
or U768 (N_768,In_871,In_532);
and U769 (N_769,In_943,In_25);
nand U770 (N_770,In_754,In_542);
and U771 (N_771,In_678,In_829);
nand U772 (N_772,In_13,In_913);
or U773 (N_773,In_844,In_904);
or U774 (N_774,In_308,In_99);
or U775 (N_775,In_262,In_130);
and U776 (N_776,In_914,In_841);
or U777 (N_777,In_223,In_934);
or U778 (N_778,In_536,In_721);
or U779 (N_779,In_234,In_184);
nand U780 (N_780,In_432,In_648);
nand U781 (N_781,In_609,In_219);
or U782 (N_782,In_590,In_820);
nor U783 (N_783,In_525,In_970);
and U784 (N_784,In_254,In_752);
and U785 (N_785,In_157,In_491);
and U786 (N_786,In_605,In_766);
nand U787 (N_787,In_289,In_676);
nor U788 (N_788,In_755,In_768);
or U789 (N_789,In_342,In_635);
or U790 (N_790,In_206,In_546);
nor U791 (N_791,In_837,In_90);
nand U792 (N_792,In_825,In_983);
nor U793 (N_793,In_405,In_636);
or U794 (N_794,In_672,In_808);
or U795 (N_795,In_846,In_476);
nand U796 (N_796,In_552,In_67);
and U797 (N_797,In_302,In_703);
and U798 (N_798,In_524,In_252);
nor U799 (N_799,In_511,In_593);
or U800 (N_800,In_921,In_48);
nor U801 (N_801,In_504,In_655);
nand U802 (N_802,In_632,In_568);
and U803 (N_803,In_938,In_165);
nand U804 (N_804,In_923,In_877);
nor U805 (N_805,In_672,In_800);
or U806 (N_806,In_42,In_867);
nor U807 (N_807,In_756,In_337);
nand U808 (N_808,In_848,In_474);
nand U809 (N_809,In_922,In_442);
and U810 (N_810,In_10,In_238);
and U811 (N_811,In_393,In_893);
nor U812 (N_812,In_168,In_376);
nand U813 (N_813,In_839,In_43);
or U814 (N_814,In_474,In_110);
nor U815 (N_815,In_753,In_737);
nand U816 (N_816,In_178,In_0);
or U817 (N_817,In_785,In_923);
and U818 (N_818,In_5,In_692);
or U819 (N_819,In_656,In_401);
nand U820 (N_820,In_901,In_868);
nor U821 (N_821,In_993,In_21);
and U822 (N_822,In_960,In_210);
nand U823 (N_823,In_391,In_470);
nand U824 (N_824,In_830,In_650);
nand U825 (N_825,In_22,In_987);
and U826 (N_826,In_310,In_215);
nor U827 (N_827,In_320,In_20);
nand U828 (N_828,In_524,In_480);
nand U829 (N_829,In_711,In_959);
and U830 (N_830,In_896,In_738);
or U831 (N_831,In_477,In_799);
nand U832 (N_832,In_316,In_407);
nand U833 (N_833,In_616,In_259);
nor U834 (N_834,In_428,In_789);
and U835 (N_835,In_416,In_313);
or U836 (N_836,In_758,In_795);
or U837 (N_837,In_710,In_362);
nand U838 (N_838,In_500,In_779);
nor U839 (N_839,In_120,In_244);
or U840 (N_840,In_324,In_570);
or U841 (N_841,In_887,In_966);
nand U842 (N_842,In_83,In_624);
nor U843 (N_843,In_9,In_454);
nand U844 (N_844,In_250,In_36);
nor U845 (N_845,In_646,In_381);
and U846 (N_846,In_875,In_700);
and U847 (N_847,In_99,In_207);
or U848 (N_848,In_95,In_870);
nor U849 (N_849,In_817,In_340);
or U850 (N_850,In_496,In_807);
or U851 (N_851,In_331,In_218);
and U852 (N_852,In_435,In_966);
and U853 (N_853,In_293,In_680);
and U854 (N_854,In_204,In_313);
nor U855 (N_855,In_401,In_275);
nand U856 (N_856,In_358,In_531);
nand U857 (N_857,In_506,In_482);
nor U858 (N_858,In_260,In_986);
nor U859 (N_859,In_320,In_87);
nor U860 (N_860,In_939,In_66);
nor U861 (N_861,In_757,In_747);
nand U862 (N_862,In_485,In_74);
or U863 (N_863,In_474,In_156);
and U864 (N_864,In_440,In_969);
or U865 (N_865,In_162,In_535);
nand U866 (N_866,In_796,In_834);
and U867 (N_867,In_959,In_747);
or U868 (N_868,In_981,In_575);
nand U869 (N_869,In_895,In_727);
nor U870 (N_870,In_890,In_54);
nand U871 (N_871,In_762,In_192);
or U872 (N_872,In_998,In_907);
nor U873 (N_873,In_835,In_977);
and U874 (N_874,In_719,In_104);
and U875 (N_875,In_310,In_606);
nand U876 (N_876,In_761,In_503);
and U877 (N_877,In_17,In_123);
or U878 (N_878,In_878,In_700);
or U879 (N_879,In_605,In_406);
nor U880 (N_880,In_32,In_844);
and U881 (N_881,In_141,In_398);
or U882 (N_882,In_218,In_393);
and U883 (N_883,In_404,In_187);
nand U884 (N_884,In_735,In_77);
nand U885 (N_885,In_739,In_935);
nand U886 (N_886,In_716,In_706);
or U887 (N_887,In_882,In_991);
nand U888 (N_888,In_340,In_32);
nor U889 (N_889,In_339,In_771);
and U890 (N_890,In_627,In_929);
nor U891 (N_891,In_331,In_854);
or U892 (N_892,In_523,In_705);
or U893 (N_893,In_616,In_260);
or U894 (N_894,In_570,In_772);
or U895 (N_895,In_729,In_140);
nor U896 (N_896,In_869,In_146);
and U897 (N_897,In_751,In_673);
and U898 (N_898,In_731,In_681);
and U899 (N_899,In_685,In_111);
nor U900 (N_900,In_216,In_986);
or U901 (N_901,In_545,In_417);
or U902 (N_902,In_28,In_770);
nor U903 (N_903,In_679,In_876);
nor U904 (N_904,In_286,In_775);
and U905 (N_905,In_283,In_680);
nor U906 (N_906,In_658,In_24);
or U907 (N_907,In_675,In_478);
and U908 (N_908,In_855,In_548);
nor U909 (N_909,In_849,In_461);
and U910 (N_910,In_697,In_179);
nand U911 (N_911,In_374,In_473);
or U912 (N_912,In_137,In_688);
or U913 (N_913,In_23,In_655);
nand U914 (N_914,In_410,In_213);
and U915 (N_915,In_763,In_974);
and U916 (N_916,In_607,In_522);
nor U917 (N_917,In_165,In_272);
and U918 (N_918,In_372,In_512);
nor U919 (N_919,In_256,In_460);
and U920 (N_920,In_527,In_786);
and U921 (N_921,In_999,In_919);
and U922 (N_922,In_596,In_859);
nor U923 (N_923,In_650,In_339);
or U924 (N_924,In_418,In_561);
nand U925 (N_925,In_95,In_345);
or U926 (N_926,In_633,In_721);
or U927 (N_927,In_756,In_914);
and U928 (N_928,In_256,In_960);
nor U929 (N_929,In_403,In_631);
nor U930 (N_930,In_409,In_138);
nand U931 (N_931,In_517,In_952);
and U932 (N_932,In_904,In_741);
nor U933 (N_933,In_297,In_275);
nor U934 (N_934,In_830,In_786);
or U935 (N_935,In_987,In_980);
nor U936 (N_936,In_494,In_768);
or U937 (N_937,In_849,In_151);
nand U938 (N_938,In_382,In_61);
and U939 (N_939,In_42,In_643);
nand U940 (N_940,In_600,In_914);
and U941 (N_941,In_620,In_671);
and U942 (N_942,In_12,In_550);
xor U943 (N_943,In_211,In_937);
and U944 (N_944,In_54,In_340);
nand U945 (N_945,In_600,In_652);
nand U946 (N_946,In_203,In_697);
or U947 (N_947,In_545,In_517);
and U948 (N_948,In_390,In_848);
or U949 (N_949,In_786,In_388);
or U950 (N_950,In_213,In_107);
and U951 (N_951,In_954,In_579);
nand U952 (N_952,In_976,In_50);
nor U953 (N_953,In_312,In_81);
nor U954 (N_954,In_671,In_723);
and U955 (N_955,In_831,In_852);
nor U956 (N_956,In_425,In_549);
and U957 (N_957,In_412,In_704);
xor U958 (N_958,In_365,In_999);
and U959 (N_959,In_398,In_341);
or U960 (N_960,In_830,In_792);
or U961 (N_961,In_893,In_184);
nand U962 (N_962,In_264,In_213);
nand U963 (N_963,In_45,In_432);
and U964 (N_964,In_718,In_211);
or U965 (N_965,In_391,In_715);
nor U966 (N_966,In_277,In_85);
nand U967 (N_967,In_203,In_946);
xnor U968 (N_968,In_514,In_728);
and U969 (N_969,In_919,In_51);
nand U970 (N_970,In_576,In_385);
or U971 (N_971,In_412,In_333);
or U972 (N_972,In_747,In_795);
nand U973 (N_973,In_385,In_66);
and U974 (N_974,In_654,In_443);
nand U975 (N_975,In_546,In_73);
nor U976 (N_976,In_342,In_190);
and U977 (N_977,In_6,In_585);
and U978 (N_978,In_981,In_467);
or U979 (N_979,In_9,In_294);
xor U980 (N_980,In_439,In_733);
or U981 (N_981,In_96,In_588);
or U982 (N_982,In_988,In_534);
nand U983 (N_983,In_399,In_88);
or U984 (N_984,In_111,In_329);
and U985 (N_985,In_375,In_881);
or U986 (N_986,In_959,In_124);
or U987 (N_987,In_405,In_979);
nand U988 (N_988,In_326,In_594);
or U989 (N_989,In_432,In_515);
nand U990 (N_990,In_84,In_697);
or U991 (N_991,In_953,In_932);
nand U992 (N_992,In_791,In_379);
nand U993 (N_993,In_677,In_472);
nand U994 (N_994,In_137,In_798);
nand U995 (N_995,In_442,In_78);
or U996 (N_996,In_109,In_335);
or U997 (N_997,In_374,In_878);
or U998 (N_998,In_444,In_809);
and U999 (N_999,In_425,In_156);
or U1000 (N_1000,N_715,N_511);
nand U1001 (N_1001,N_143,N_431);
nand U1002 (N_1002,N_301,N_16);
nand U1003 (N_1003,N_841,N_187);
nand U1004 (N_1004,N_25,N_525);
nor U1005 (N_1005,N_632,N_738);
or U1006 (N_1006,N_953,N_843);
nand U1007 (N_1007,N_427,N_188);
or U1008 (N_1008,N_647,N_332);
nand U1009 (N_1009,N_777,N_215);
nor U1010 (N_1010,N_813,N_896);
and U1011 (N_1011,N_91,N_461);
nand U1012 (N_1012,N_331,N_552);
and U1013 (N_1013,N_384,N_442);
nand U1014 (N_1014,N_463,N_283);
nor U1015 (N_1015,N_992,N_691);
or U1016 (N_1016,N_577,N_959);
nor U1017 (N_1017,N_54,N_419);
nor U1018 (N_1018,N_564,N_704);
nand U1019 (N_1019,N_29,N_53);
nor U1020 (N_1020,N_151,N_327);
or U1021 (N_1021,N_558,N_836);
and U1022 (N_1022,N_127,N_14);
nand U1023 (N_1023,N_369,N_263);
or U1024 (N_1024,N_454,N_993);
nor U1025 (N_1025,N_687,N_723);
nand U1026 (N_1026,N_638,N_167);
nor U1027 (N_1027,N_351,N_917);
nand U1028 (N_1028,N_951,N_858);
and U1029 (N_1029,N_627,N_550);
nand U1030 (N_1030,N_132,N_923);
xnor U1031 (N_1031,N_926,N_866);
nand U1032 (N_1032,N_815,N_329);
nand U1033 (N_1033,N_981,N_854);
nand U1034 (N_1034,N_977,N_678);
nor U1035 (N_1035,N_533,N_878);
or U1036 (N_1036,N_804,N_877);
nor U1037 (N_1037,N_223,N_174);
nand U1038 (N_1038,N_747,N_855);
nand U1039 (N_1039,N_293,N_278);
nand U1040 (N_1040,N_520,N_319);
nand U1041 (N_1041,N_537,N_938);
nor U1042 (N_1042,N_267,N_801);
and U1043 (N_1043,N_749,N_139);
or U1044 (N_1044,N_249,N_527);
or U1045 (N_1045,N_238,N_985);
and U1046 (N_1046,N_549,N_844);
or U1047 (N_1047,N_48,N_580);
or U1048 (N_1048,N_184,N_288);
or U1049 (N_1049,N_501,N_640);
or U1050 (N_1050,N_496,N_244);
nand U1051 (N_1051,N_446,N_780);
nor U1052 (N_1052,N_897,N_826);
nand U1053 (N_1053,N_927,N_483);
or U1054 (N_1054,N_593,N_879);
nor U1055 (N_1055,N_333,N_444);
and U1056 (N_1056,N_769,N_544);
nor U1057 (N_1057,N_756,N_845);
or U1058 (N_1058,N_27,N_388);
nor U1059 (N_1059,N_375,N_448);
nand U1060 (N_1060,N_712,N_925);
nor U1061 (N_1061,N_366,N_596);
nand U1062 (N_1062,N_141,N_659);
nor U1063 (N_1063,N_860,N_8);
or U1064 (N_1064,N_373,N_420);
nand U1065 (N_1065,N_401,N_553);
nand U1066 (N_1066,N_386,N_318);
nand U1067 (N_1067,N_284,N_277);
or U1068 (N_1068,N_831,N_493);
nand U1069 (N_1069,N_563,N_618);
and U1070 (N_1070,N_65,N_983);
nor U1071 (N_1071,N_44,N_107);
nor U1072 (N_1072,N_68,N_603);
and U1073 (N_1073,N_814,N_526);
and U1074 (N_1074,N_701,N_908);
or U1075 (N_1075,N_458,N_965);
or U1076 (N_1076,N_958,N_498);
and U1077 (N_1077,N_195,N_246);
or U1078 (N_1078,N_689,N_730);
or U1079 (N_1079,N_272,N_51);
or U1080 (N_1080,N_692,N_741);
nor U1081 (N_1081,N_688,N_186);
nand U1082 (N_1082,N_613,N_385);
or U1083 (N_1083,N_79,N_297);
or U1084 (N_1084,N_534,N_954);
or U1085 (N_1085,N_700,N_341);
nand U1086 (N_1086,N_9,N_115);
and U1087 (N_1087,N_674,N_616);
and U1088 (N_1088,N_709,N_473);
nor U1089 (N_1089,N_846,N_735);
nor U1090 (N_1090,N_821,N_683);
and U1091 (N_1091,N_979,N_905);
nand U1092 (N_1092,N_262,N_323);
nor U1093 (N_1093,N_468,N_380);
nor U1094 (N_1094,N_149,N_309);
nor U1095 (N_1095,N_58,N_538);
nor U1096 (N_1096,N_285,N_911);
nand U1097 (N_1097,N_716,N_52);
xor U1098 (N_1098,N_212,N_121);
or U1099 (N_1099,N_337,N_59);
nand U1100 (N_1100,N_984,N_447);
nand U1101 (N_1101,N_727,N_806);
nand U1102 (N_1102,N_834,N_276);
nor U1103 (N_1103,N_104,N_820);
nand U1104 (N_1104,N_363,N_376);
or U1105 (N_1105,N_529,N_587);
nand U1106 (N_1106,N_731,N_695);
nor U1107 (N_1107,N_898,N_205);
nor U1108 (N_1108,N_494,N_887);
or U1109 (N_1109,N_637,N_766);
nor U1110 (N_1110,N_795,N_807);
nand U1111 (N_1111,N_377,N_528);
nand U1112 (N_1112,N_560,N_429);
and U1113 (N_1113,N_606,N_98);
and U1114 (N_1114,N_340,N_764);
nand U1115 (N_1115,N_11,N_699);
nand U1116 (N_1116,N_290,N_97);
nor U1117 (N_1117,N_171,N_93);
nand U1118 (N_1118,N_698,N_559);
nor U1119 (N_1119,N_455,N_912);
or U1120 (N_1120,N_609,N_464);
nand U1121 (N_1121,N_907,N_33);
and U1122 (N_1122,N_909,N_517);
nor U1123 (N_1123,N_971,N_502);
nor U1124 (N_1124,N_681,N_658);
nor U1125 (N_1125,N_867,N_610);
and U1126 (N_1126,N_15,N_325);
and U1127 (N_1127,N_418,N_236);
nor U1128 (N_1128,N_177,N_729);
or U1129 (N_1129,N_936,N_734);
or U1130 (N_1130,N_405,N_686);
nor U1131 (N_1131,N_160,N_862);
nor U1132 (N_1132,N_356,N_438);
and U1133 (N_1133,N_191,N_57);
or U1134 (N_1134,N_792,N_144);
nor U1135 (N_1135,N_379,N_824);
nor U1136 (N_1136,N_955,N_154);
nand U1137 (N_1137,N_176,N_428);
and U1138 (N_1138,N_714,N_449);
nor U1139 (N_1139,N_671,N_287);
nor U1140 (N_1140,N_55,N_200);
nand U1141 (N_1141,N_583,N_956);
or U1142 (N_1142,N_503,N_805);
nor U1143 (N_1143,N_443,N_932);
and U1144 (N_1144,N_126,N_226);
nor U1145 (N_1145,N_181,N_588);
and U1146 (N_1146,N_988,N_778);
or U1147 (N_1147,N_417,N_653);
nand U1148 (N_1148,N_894,N_88);
nor U1149 (N_1149,N_865,N_743);
nand U1150 (N_1150,N_888,N_291);
nor U1151 (N_1151,N_515,N_651);
nor U1152 (N_1152,N_684,N_321);
nor U1153 (N_1153,N_83,N_962);
nand U1154 (N_1154,N_702,N_122);
or U1155 (N_1155,N_994,N_668);
nand U1156 (N_1156,N_343,N_763);
or U1157 (N_1157,N_775,N_541);
nand U1158 (N_1158,N_219,N_934);
nand U1159 (N_1159,N_545,N_625);
nor U1160 (N_1160,N_895,N_620);
or U1161 (N_1161,N_378,N_940);
nor U1162 (N_1162,N_270,N_239);
nand U1163 (N_1163,N_724,N_316);
nor U1164 (N_1164,N_679,N_64);
and U1165 (N_1165,N_46,N_335);
nand U1166 (N_1166,N_793,N_250);
nand U1167 (N_1167,N_75,N_95);
nor U1168 (N_1168,N_818,N_995);
nor U1169 (N_1169,N_31,N_211);
or U1170 (N_1170,N_462,N_737);
and U1171 (N_1171,N_361,N_488);
nor U1172 (N_1172,N_235,N_966);
and U1173 (N_1173,N_368,N_148);
and U1174 (N_1174,N_485,N_367);
and U1175 (N_1175,N_382,N_797);
and U1176 (N_1176,N_978,N_903);
nand U1177 (N_1177,N_633,N_299);
and U1178 (N_1178,N_773,N_359);
nor U1179 (N_1179,N_790,N_904);
nor U1180 (N_1180,N_974,N_507);
and U1181 (N_1181,N_519,N_875);
or U1182 (N_1182,N_601,N_915);
nand U1183 (N_1183,N_562,N_352);
nand U1184 (N_1184,N_812,N_74);
or U1185 (N_1185,N_592,N_349);
nand U1186 (N_1186,N_849,N_931);
nor U1187 (N_1187,N_696,N_120);
or U1188 (N_1188,N_292,N_47);
nor U1189 (N_1189,N_883,N_134);
and U1190 (N_1190,N_540,N_221);
or U1191 (N_1191,N_358,N_21);
and U1192 (N_1192,N_664,N_848);
or U1193 (N_1193,N_391,N_989);
or U1194 (N_1194,N_271,N_576);
and U1195 (N_1195,N_232,N_430);
nand U1196 (N_1196,N_961,N_713);
and U1197 (N_1197,N_476,N_662);
nand U1198 (N_1198,N_5,N_639);
or U1199 (N_1199,N_796,N_156);
and U1200 (N_1200,N_789,N_542);
nand U1201 (N_1201,N_510,N_178);
and U1202 (N_1202,N_452,N_300);
or U1203 (N_1203,N_35,N_539);
nand U1204 (N_1204,N_157,N_784);
and U1205 (N_1205,N_666,N_179);
and U1206 (N_1206,N_705,N_106);
and U1207 (N_1207,N_586,N_536);
or U1208 (N_1208,N_776,N_948);
nand U1209 (N_1209,N_920,N_767);
and U1210 (N_1210,N_269,N_350);
and U1211 (N_1211,N_924,N_108);
nor U1212 (N_1212,N_117,N_102);
nor U1213 (N_1213,N_234,N_437);
or U1214 (N_1214,N_611,N_18);
and U1215 (N_1215,N_116,N_851);
nor U1216 (N_1216,N_261,N_310);
nor U1217 (N_1217,N_61,N_968);
nor U1218 (N_1218,N_275,N_175);
nand U1219 (N_1219,N_644,N_779);
or U1220 (N_1220,N_710,N_402);
and U1221 (N_1221,N_312,N_508);
and U1222 (N_1222,N_86,N_92);
and U1223 (N_1223,N_227,N_937);
nand U1224 (N_1224,N_248,N_198);
or U1225 (N_1225,N_395,N_868);
nor U1226 (N_1226,N_78,N_311);
nor U1227 (N_1227,N_600,N_880);
or U1228 (N_1228,N_711,N_213);
nand U1229 (N_1229,N_146,N_233);
or U1230 (N_1230,N_921,N_825);
nand U1231 (N_1231,N_757,N_914);
nor U1232 (N_1232,N_80,N_646);
nor U1233 (N_1233,N_125,N_857);
nand U1234 (N_1234,N_902,N_336);
and U1235 (N_1235,N_969,N_750);
nor U1236 (N_1236,N_876,N_303);
nand U1237 (N_1237,N_885,N_130);
or U1238 (N_1238,N_295,N_416);
nand U1239 (N_1239,N_282,N_216);
nand U1240 (N_1240,N_669,N_803);
or U1241 (N_1241,N_393,N_946);
nand U1242 (N_1242,N_241,N_166);
nor U1243 (N_1243,N_390,N_572);
and U1244 (N_1244,N_830,N_354);
and U1245 (N_1245,N_294,N_403);
or U1246 (N_1246,N_870,N_414);
nor U1247 (N_1247,N_650,N_101);
or U1248 (N_1248,N_459,N_60);
nor U1249 (N_1249,N_231,N_218);
nand U1250 (N_1250,N_251,N_739);
nand U1251 (N_1251,N_694,N_582);
nor U1252 (N_1252,N_162,N_131);
nand U1253 (N_1253,N_168,N_242);
or U1254 (N_1254,N_863,N_87);
nand U1255 (N_1255,N_163,N_800);
and U1256 (N_1256,N_736,N_900);
and U1257 (N_1257,N_569,N_113);
nand U1258 (N_1258,N_40,N_94);
or U1259 (N_1259,N_258,N_947);
nand U1260 (N_1260,N_45,N_706);
or U1261 (N_1261,N_364,N_4);
nand U1262 (N_1262,N_348,N_257);
nand U1263 (N_1263,N_513,N_150);
nor U1264 (N_1264,N_7,N_518);
or U1265 (N_1265,N_543,N_661);
nor U1266 (N_1266,N_822,N_85);
or U1267 (N_1267,N_135,N_584);
nand U1268 (N_1268,N_567,N_114);
nand U1269 (N_1269,N_49,N_383);
or U1270 (N_1270,N_708,N_998);
or U1271 (N_1271,N_305,N_636);
or U1272 (N_1272,N_774,N_982);
or U1273 (N_1273,N_434,N_964);
nand U1274 (N_1274,N_794,N_893);
or U1275 (N_1275,N_480,N_71);
or U1276 (N_1276,N_635,N_392);
nor U1277 (N_1277,N_328,N_207);
nor U1278 (N_1278,N_289,N_952);
or U1279 (N_1279,N_859,N_3);
nand U1280 (N_1280,N_471,N_758);
and U1281 (N_1281,N_524,N_838);
or U1282 (N_1282,N_703,N_34);
nand U1283 (N_1283,N_62,N_939);
or U1284 (N_1284,N_585,N_128);
nor U1285 (N_1285,N_980,N_594);
nor U1286 (N_1286,N_597,N_387);
or U1287 (N_1287,N_381,N_274);
or U1288 (N_1288,N_612,N_406);
or U1289 (N_1289,N_889,N_628);
or U1290 (N_1290,N_630,N_619);
nor U1291 (N_1291,N_840,N_864);
nand U1292 (N_1292,N_762,N_677);
nor U1293 (N_1293,N_673,N_499);
nor U1294 (N_1294,N_718,N_882);
nor U1295 (N_1295,N_6,N_753);
and U1296 (N_1296,N_22,N_259);
and U1297 (N_1297,N_665,N_930);
and U1298 (N_1298,N_667,N_960);
nand U1299 (N_1299,N_30,N_590);
and U1300 (N_1300,N_260,N_90);
or U1301 (N_1301,N_365,N_73);
nor U1302 (N_1302,N_802,N_173);
or U1303 (N_1303,N_422,N_547);
and U1304 (N_1304,N_41,N_76);
nor U1305 (N_1305,N_591,N_672);
or U1306 (N_1306,N_469,N_353);
xor U1307 (N_1307,N_23,N_436);
nor U1308 (N_1308,N_362,N_599);
and U1309 (N_1309,N_505,N_771);
or U1310 (N_1310,N_786,N_404);
and U1311 (N_1311,N_514,N_396);
nand U1312 (N_1312,N_225,N_133);
nor U1313 (N_1313,N_0,N_214);
nor U1314 (N_1314,N_70,N_754);
or U1315 (N_1315,N_782,N_629);
nand U1316 (N_1316,N_910,N_622);
nor U1317 (N_1317,N_342,N_69);
or U1318 (N_1318,N_975,N_506);
and U1319 (N_1319,N_147,N_761);
or U1320 (N_1320,N_624,N_256);
nor U1321 (N_1321,N_660,N_929);
nor U1322 (N_1322,N_949,N_861);
or U1323 (N_1323,N_690,N_19);
nand U1324 (N_1324,N_206,N_987);
or U1325 (N_1325,N_602,N_685);
and U1326 (N_1326,N_566,N_732);
nor U1327 (N_1327,N_280,N_509);
nand U1328 (N_1328,N_138,N_752);
nand U1329 (N_1329,N_663,N_435);
nor U1330 (N_1330,N_265,N_605);
or U1331 (N_1331,N_322,N_886);
or U1332 (N_1332,N_424,N_273);
nor U1333 (N_1333,N_770,N_648);
nor U1334 (N_1334,N_913,N_823);
and U1335 (N_1335,N_456,N_159);
nor U1336 (N_1336,N_398,N_66);
or U1337 (N_1337,N_571,N_719);
or U1338 (N_1338,N_82,N_111);
nand U1339 (N_1339,N_581,N_313);
or U1340 (N_1340,N_495,N_783);
nor U1341 (N_1341,N_266,N_772);
nand U1342 (N_1342,N_12,N_453);
nand U1343 (N_1343,N_56,N_475);
or U1344 (N_1344,N_728,N_941);
and U1345 (N_1345,N_415,N_306);
and U1346 (N_1346,N_467,N_155);
or U1347 (N_1347,N_872,N_986);
and U1348 (N_1348,N_140,N_145);
or U1349 (N_1349,N_472,N_720);
nor U1350 (N_1350,N_43,N_487);
nor U1351 (N_1351,N_199,N_268);
nor U1352 (N_1352,N_871,N_680);
and U1353 (N_1353,N_649,N_707);
or U1354 (N_1354,N_445,N_615);
and U1355 (N_1355,N_193,N_555);
nand U1356 (N_1356,N_996,N_89);
nor U1357 (N_1357,N_165,N_370);
nor U1358 (N_1358,N_497,N_972);
nand U1359 (N_1359,N_810,N_164);
nor U1360 (N_1360,N_847,N_99);
or U1361 (N_1361,N_486,N_474);
and U1362 (N_1362,N_412,N_570);
and U1363 (N_1363,N_439,N_787);
or U1364 (N_1364,N_109,N_976);
nand U1365 (N_1365,N_411,N_400);
nor U1366 (N_1366,N_643,N_255);
nand U1367 (N_1367,N_24,N_748);
and U1368 (N_1368,N_899,N_264);
nand U1369 (N_1369,N_489,N_183);
nand U1370 (N_1370,N_110,N_809);
nand U1371 (N_1371,N_788,N_389);
or U1372 (N_1372,N_522,N_891);
and U1373 (N_1373,N_245,N_355);
or U1374 (N_1374,N_153,N_169);
and U1375 (N_1375,N_433,N_642);
nand U1376 (N_1376,N_478,N_614);
nand U1377 (N_1377,N_657,N_170);
nand U1378 (N_1378,N_32,N_217);
and U1379 (N_1379,N_161,N_338);
nand U1380 (N_1380,N_450,N_967);
or U1381 (N_1381,N_1,N_50);
nor U1382 (N_1382,N_394,N_717);
nor U1383 (N_1383,N_408,N_39);
nand U1384 (N_1384,N_320,N_196);
and U1385 (N_1385,N_799,N_465);
or U1386 (N_1386,N_816,N_237);
nor U1387 (N_1387,N_315,N_837);
or U1388 (N_1388,N_204,N_565);
nor U1389 (N_1389,N_791,N_693);
nor U1390 (N_1390,N_928,N_421);
and U1391 (N_1391,N_733,N_742);
nand U1392 (N_1392,N_656,N_304);
nor U1393 (N_1393,N_568,N_308);
nand U1394 (N_1394,N_96,N_890);
and U1395 (N_1395,N_374,N_504);
and U1396 (N_1396,N_197,N_781);
or U1397 (N_1397,N_675,N_247);
nor U1398 (N_1398,N_722,N_38);
nand U1399 (N_1399,N_477,N_189);
and U1400 (N_1400,N_479,N_918);
nor U1401 (N_1401,N_842,N_230);
nand U1402 (N_1402,N_484,N_314);
nor U1403 (N_1403,N_142,N_210);
nor U1404 (N_1404,N_228,N_641);
nand U1405 (N_1405,N_835,N_595);
nor U1406 (N_1406,N_626,N_10);
or U1407 (N_1407,N_935,N_281);
or U1408 (N_1408,N_347,N_129);
nand U1409 (N_1409,N_252,N_943);
nand U1410 (N_1410,N_209,N_426);
or U1411 (N_1411,N_745,N_828);
nand U1412 (N_1412,N_37,N_2);
nand U1413 (N_1413,N_185,N_551);
or U1414 (N_1414,N_17,N_645);
or U1415 (N_1415,N_670,N_208);
nand U1416 (N_1416,N_158,N_326);
or U1417 (N_1417,N_42,N_973);
nand U1418 (N_1418,N_654,N_922);
nand U1419 (N_1419,N_919,N_617);
or U1420 (N_1420,N_123,N_224);
or U1421 (N_1421,N_811,N_124);
nor U1422 (N_1422,N_202,N_873);
or U1423 (N_1423,N_697,N_324);
nor U1424 (N_1424,N_192,N_970);
nor U1425 (N_1425,N_77,N_357);
nand U1426 (N_1426,N_521,N_36);
nand U1427 (N_1427,N_317,N_118);
nor U1428 (N_1428,N_407,N_307);
nor U1429 (N_1429,N_190,N_460);
nand U1430 (N_1430,N_604,N_286);
and U1431 (N_1431,N_578,N_765);
or U1432 (N_1432,N_573,N_491);
or U1433 (N_1433,N_523,N_254);
or U1434 (N_1434,N_399,N_152);
nand U1435 (N_1435,N_901,N_512);
nand U1436 (N_1436,N_997,N_798);
nand U1437 (N_1437,N_833,N_634);
and U1438 (N_1438,N_759,N_302);
nand U1439 (N_1439,N_817,N_751);
nand U1440 (N_1440,N_829,N_916);
or U1441 (N_1441,N_874,N_410);
nand U1442 (N_1442,N_105,N_345);
nand U1443 (N_1443,N_999,N_253);
and U1444 (N_1444,N_852,N_746);
or U1445 (N_1445,N_136,N_72);
or U1446 (N_1446,N_548,N_906);
nand U1447 (N_1447,N_740,N_84);
or U1448 (N_1448,N_963,N_853);
or U1449 (N_1449,N_330,N_516);
and U1450 (N_1450,N_631,N_482);
xnor U1451 (N_1451,N_298,N_81);
and U1452 (N_1452,N_682,N_676);
nand U1453 (N_1453,N_220,N_623);
nor U1454 (N_1454,N_579,N_608);
nor U1455 (N_1455,N_850,N_112);
nand U1456 (N_1456,N_856,N_194);
nor U1457 (N_1457,N_532,N_334);
nand U1458 (N_1458,N_607,N_432);
and U1459 (N_1459,N_457,N_103);
nand U1460 (N_1460,N_137,N_481);
or U1461 (N_1461,N_466,N_832);
nor U1462 (N_1462,N_20,N_409);
nor U1463 (N_1463,N_933,N_827);
xnor U1464 (N_1464,N_279,N_892);
and U1465 (N_1465,N_13,N_425);
or U1466 (N_1466,N_222,N_451);
nand U1467 (N_1467,N_768,N_755);
nor U1468 (N_1468,N_182,N_945);
or U1469 (N_1469,N_490,N_839);
or U1470 (N_1470,N_990,N_371);
nand U1471 (N_1471,N_575,N_63);
nand U1472 (N_1472,N_808,N_535);
nor U1473 (N_1473,N_621,N_869);
nand U1474 (N_1474,N_589,N_26);
and U1475 (N_1475,N_172,N_561);
and U1476 (N_1476,N_470,N_944);
or U1477 (N_1477,N_881,N_652);
nor U1478 (N_1478,N_554,N_203);
and U1479 (N_1479,N_721,N_229);
or U1480 (N_1480,N_397,N_574);
nand U1481 (N_1481,N_957,N_344);
and U1482 (N_1482,N_557,N_726);
nand U1483 (N_1483,N_500,N_785);
and U1484 (N_1484,N_546,N_760);
nor U1485 (N_1485,N_942,N_655);
or U1486 (N_1486,N_180,N_492);
nand U1487 (N_1487,N_372,N_819);
nor U1488 (N_1488,N_360,N_413);
nand U1489 (N_1489,N_530,N_744);
nand U1490 (N_1490,N_991,N_725);
nand U1491 (N_1491,N_440,N_67);
xnor U1492 (N_1492,N_531,N_296);
nand U1493 (N_1493,N_201,N_28);
nand U1494 (N_1494,N_950,N_100);
and U1495 (N_1495,N_346,N_119);
nor U1496 (N_1496,N_884,N_243);
nor U1497 (N_1497,N_598,N_556);
and U1498 (N_1498,N_339,N_441);
nor U1499 (N_1499,N_240,N_423);
or U1500 (N_1500,N_241,N_434);
and U1501 (N_1501,N_458,N_634);
nor U1502 (N_1502,N_72,N_355);
or U1503 (N_1503,N_173,N_497);
or U1504 (N_1504,N_781,N_72);
or U1505 (N_1505,N_64,N_636);
and U1506 (N_1506,N_361,N_420);
nand U1507 (N_1507,N_906,N_318);
or U1508 (N_1508,N_427,N_623);
nand U1509 (N_1509,N_628,N_259);
nor U1510 (N_1510,N_215,N_437);
xnor U1511 (N_1511,N_531,N_33);
or U1512 (N_1512,N_688,N_602);
nand U1513 (N_1513,N_394,N_64);
nor U1514 (N_1514,N_711,N_607);
or U1515 (N_1515,N_228,N_542);
nand U1516 (N_1516,N_859,N_279);
nand U1517 (N_1517,N_585,N_729);
nor U1518 (N_1518,N_254,N_252);
nor U1519 (N_1519,N_41,N_23);
nor U1520 (N_1520,N_556,N_827);
nor U1521 (N_1521,N_868,N_816);
nand U1522 (N_1522,N_336,N_137);
or U1523 (N_1523,N_470,N_340);
and U1524 (N_1524,N_538,N_454);
and U1525 (N_1525,N_76,N_173);
and U1526 (N_1526,N_583,N_298);
nand U1527 (N_1527,N_225,N_122);
nor U1528 (N_1528,N_881,N_670);
or U1529 (N_1529,N_154,N_496);
and U1530 (N_1530,N_925,N_33);
and U1531 (N_1531,N_748,N_539);
nand U1532 (N_1532,N_876,N_669);
or U1533 (N_1533,N_201,N_263);
nand U1534 (N_1534,N_560,N_278);
nor U1535 (N_1535,N_715,N_33);
or U1536 (N_1536,N_702,N_16);
and U1537 (N_1537,N_844,N_664);
or U1538 (N_1538,N_869,N_866);
and U1539 (N_1539,N_608,N_755);
and U1540 (N_1540,N_375,N_326);
nor U1541 (N_1541,N_832,N_545);
nor U1542 (N_1542,N_564,N_964);
nor U1543 (N_1543,N_443,N_43);
nand U1544 (N_1544,N_965,N_439);
nor U1545 (N_1545,N_175,N_880);
nor U1546 (N_1546,N_109,N_739);
or U1547 (N_1547,N_887,N_256);
nor U1548 (N_1548,N_942,N_244);
or U1549 (N_1549,N_696,N_798);
and U1550 (N_1550,N_793,N_91);
nand U1551 (N_1551,N_671,N_946);
nor U1552 (N_1552,N_986,N_607);
and U1553 (N_1553,N_695,N_908);
nand U1554 (N_1554,N_146,N_345);
nand U1555 (N_1555,N_869,N_257);
nor U1556 (N_1556,N_33,N_181);
and U1557 (N_1557,N_404,N_356);
and U1558 (N_1558,N_71,N_208);
and U1559 (N_1559,N_500,N_882);
or U1560 (N_1560,N_109,N_289);
or U1561 (N_1561,N_713,N_244);
nand U1562 (N_1562,N_808,N_330);
nor U1563 (N_1563,N_731,N_285);
nand U1564 (N_1564,N_415,N_470);
nand U1565 (N_1565,N_440,N_380);
nand U1566 (N_1566,N_758,N_425);
and U1567 (N_1567,N_936,N_367);
or U1568 (N_1568,N_349,N_781);
nand U1569 (N_1569,N_714,N_112);
nand U1570 (N_1570,N_183,N_314);
or U1571 (N_1571,N_658,N_348);
or U1572 (N_1572,N_642,N_128);
nor U1573 (N_1573,N_862,N_122);
nand U1574 (N_1574,N_561,N_86);
nor U1575 (N_1575,N_913,N_279);
and U1576 (N_1576,N_870,N_221);
and U1577 (N_1577,N_919,N_912);
nor U1578 (N_1578,N_863,N_212);
nor U1579 (N_1579,N_841,N_206);
nand U1580 (N_1580,N_287,N_780);
and U1581 (N_1581,N_821,N_713);
nand U1582 (N_1582,N_118,N_376);
nor U1583 (N_1583,N_56,N_124);
nand U1584 (N_1584,N_355,N_728);
nor U1585 (N_1585,N_936,N_754);
nand U1586 (N_1586,N_133,N_355);
or U1587 (N_1587,N_380,N_613);
nand U1588 (N_1588,N_526,N_569);
or U1589 (N_1589,N_749,N_285);
and U1590 (N_1590,N_580,N_762);
and U1591 (N_1591,N_954,N_578);
nor U1592 (N_1592,N_860,N_999);
or U1593 (N_1593,N_121,N_317);
or U1594 (N_1594,N_360,N_870);
or U1595 (N_1595,N_776,N_848);
or U1596 (N_1596,N_632,N_837);
nand U1597 (N_1597,N_661,N_953);
nor U1598 (N_1598,N_646,N_884);
nor U1599 (N_1599,N_714,N_611);
nand U1600 (N_1600,N_698,N_232);
nor U1601 (N_1601,N_755,N_157);
or U1602 (N_1602,N_829,N_421);
nand U1603 (N_1603,N_39,N_957);
and U1604 (N_1604,N_967,N_729);
nand U1605 (N_1605,N_686,N_296);
nand U1606 (N_1606,N_935,N_99);
xnor U1607 (N_1607,N_484,N_758);
nand U1608 (N_1608,N_703,N_62);
nor U1609 (N_1609,N_439,N_220);
or U1610 (N_1610,N_486,N_257);
or U1611 (N_1611,N_294,N_82);
nor U1612 (N_1612,N_135,N_82);
nand U1613 (N_1613,N_49,N_864);
nand U1614 (N_1614,N_647,N_711);
and U1615 (N_1615,N_333,N_843);
nand U1616 (N_1616,N_14,N_840);
or U1617 (N_1617,N_566,N_24);
and U1618 (N_1618,N_979,N_663);
nor U1619 (N_1619,N_230,N_764);
nand U1620 (N_1620,N_85,N_27);
and U1621 (N_1621,N_638,N_106);
and U1622 (N_1622,N_545,N_343);
nand U1623 (N_1623,N_112,N_485);
nor U1624 (N_1624,N_600,N_117);
or U1625 (N_1625,N_437,N_871);
nand U1626 (N_1626,N_616,N_345);
and U1627 (N_1627,N_828,N_496);
or U1628 (N_1628,N_545,N_962);
or U1629 (N_1629,N_753,N_217);
and U1630 (N_1630,N_206,N_695);
nor U1631 (N_1631,N_893,N_95);
or U1632 (N_1632,N_18,N_550);
nand U1633 (N_1633,N_314,N_828);
nand U1634 (N_1634,N_145,N_841);
or U1635 (N_1635,N_42,N_340);
or U1636 (N_1636,N_577,N_674);
nor U1637 (N_1637,N_437,N_851);
nor U1638 (N_1638,N_855,N_320);
nand U1639 (N_1639,N_875,N_329);
and U1640 (N_1640,N_723,N_915);
nor U1641 (N_1641,N_977,N_651);
nand U1642 (N_1642,N_190,N_255);
nor U1643 (N_1643,N_392,N_856);
nand U1644 (N_1644,N_226,N_667);
and U1645 (N_1645,N_534,N_880);
or U1646 (N_1646,N_713,N_947);
and U1647 (N_1647,N_27,N_911);
nand U1648 (N_1648,N_738,N_936);
nor U1649 (N_1649,N_784,N_438);
and U1650 (N_1650,N_215,N_371);
or U1651 (N_1651,N_712,N_114);
and U1652 (N_1652,N_728,N_279);
nand U1653 (N_1653,N_605,N_46);
nand U1654 (N_1654,N_211,N_151);
or U1655 (N_1655,N_819,N_417);
nor U1656 (N_1656,N_436,N_740);
and U1657 (N_1657,N_428,N_61);
nand U1658 (N_1658,N_687,N_475);
nor U1659 (N_1659,N_149,N_487);
nor U1660 (N_1660,N_9,N_910);
or U1661 (N_1661,N_294,N_459);
or U1662 (N_1662,N_575,N_882);
or U1663 (N_1663,N_969,N_590);
nor U1664 (N_1664,N_292,N_376);
or U1665 (N_1665,N_426,N_921);
and U1666 (N_1666,N_936,N_398);
or U1667 (N_1667,N_765,N_881);
and U1668 (N_1668,N_165,N_586);
and U1669 (N_1669,N_352,N_346);
or U1670 (N_1670,N_483,N_226);
nand U1671 (N_1671,N_697,N_453);
nand U1672 (N_1672,N_370,N_679);
and U1673 (N_1673,N_566,N_113);
or U1674 (N_1674,N_517,N_598);
nand U1675 (N_1675,N_511,N_203);
nand U1676 (N_1676,N_814,N_229);
xnor U1677 (N_1677,N_351,N_289);
nand U1678 (N_1678,N_888,N_791);
and U1679 (N_1679,N_152,N_976);
and U1680 (N_1680,N_903,N_243);
nand U1681 (N_1681,N_443,N_650);
and U1682 (N_1682,N_45,N_684);
nor U1683 (N_1683,N_808,N_466);
and U1684 (N_1684,N_840,N_781);
xnor U1685 (N_1685,N_558,N_220);
nand U1686 (N_1686,N_603,N_738);
or U1687 (N_1687,N_476,N_928);
or U1688 (N_1688,N_855,N_4);
nor U1689 (N_1689,N_957,N_44);
nand U1690 (N_1690,N_816,N_60);
and U1691 (N_1691,N_765,N_572);
nand U1692 (N_1692,N_6,N_677);
or U1693 (N_1693,N_257,N_179);
or U1694 (N_1694,N_607,N_11);
nand U1695 (N_1695,N_804,N_912);
and U1696 (N_1696,N_824,N_25);
nand U1697 (N_1697,N_449,N_875);
and U1698 (N_1698,N_172,N_86);
nand U1699 (N_1699,N_480,N_37);
and U1700 (N_1700,N_483,N_96);
nand U1701 (N_1701,N_320,N_642);
and U1702 (N_1702,N_311,N_626);
nand U1703 (N_1703,N_416,N_697);
nor U1704 (N_1704,N_535,N_170);
nand U1705 (N_1705,N_963,N_162);
nand U1706 (N_1706,N_636,N_108);
nor U1707 (N_1707,N_195,N_599);
nand U1708 (N_1708,N_125,N_681);
or U1709 (N_1709,N_226,N_477);
nand U1710 (N_1710,N_511,N_147);
or U1711 (N_1711,N_656,N_786);
xnor U1712 (N_1712,N_540,N_718);
nor U1713 (N_1713,N_402,N_174);
nand U1714 (N_1714,N_535,N_171);
and U1715 (N_1715,N_348,N_340);
and U1716 (N_1716,N_313,N_673);
nand U1717 (N_1717,N_843,N_385);
nor U1718 (N_1718,N_934,N_537);
and U1719 (N_1719,N_12,N_130);
nand U1720 (N_1720,N_896,N_110);
nor U1721 (N_1721,N_546,N_692);
or U1722 (N_1722,N_106,N_891);
nand U1723 (N_1723,N_605,N_11);
and U1724 (N_1724,N_671,N_803);
or U1725 (N_1725,N_424,N_822);
and U1726 (N_1726,N_143,N_831);
and U1727 (N_1727,N_623,N_471);
nor U1728 (N_1728,N_989,N_599);
nor U1729 (N_1729,N_724,N_436);
xnor U1730 (N_1730,N_286,N_601);
nor U1731 (N_1731,N_72,N_737);
and U1732 (N_1732,N_568,N_251);
and U1733 (N_1733,N_579,N_458);
or U1734 (N_1734,N_2,N_113);
and U1735 (N_1735,N_458,N_125);
nand U1736 (N_1736,N_946,N_77);
and U1737 (N_1737,N_969,N_822);
nand U1738 (N_1738,N_349,N_472);
and U1739 (N_1739,N_905,N_581);
and U1740 (N_1740,N_346,N_579);
or U1741 (N_1741,N_231,N_608);
or U1742 (N_1742,N_352,N_446);
and U1743 (N_1743,N_466,N_880);
and U1744 (N_1744,N_213,N_236);
nor U1745 (N_1745,N_213,N_52);
nor U1746 (N_1746,N_434,N_979);
nor U1747 (N_1747,N_992,N_930);
and U1748 (N_1748,N_162,N_330);
nand U1749 (N_1749,N_480,N_905);
nand U1750 (N_1750,N_799,N_262);
nor U1751 (N_1751,N_132,N_189);
nor U1752 (N_1752,N_727,N_913);
or U1753 (N_1753,N_194,N_641);
or U1754 (N_1754,N_668,N_634);
nor U1755 (N_1755,N_594,N_984);
nand U1756 (N_1756,N_40,N_463);
nor U1757 (N_1757,N_472,N_360);
or U1758 (N_1758,N_381,N_172);
and U1759 (N_1759,N_530,N_228);
and U1760 (N_1760,N_331,N_200);
nand U1761 (N_1761,N_249,N_843);
or U1762 (N_1762,N_911,N_806);
or U1763 (N_1763,N_952,N_215);
or U1764 (N_1764,N_162,N_299);
and U1765 (N_1765,N_181,N_916);
nor U1766 (N_1766,N_375,N_745);
or U1767 (N_1767,N_356,N_13);
nand U1768 (N_1768,N_558,N_967);
nor U1769 (N_1769,N_914,N_415);
nor U1770 (N_1770,N_182,N_672);
or U1771 (N_1771,N_744,N_585);
nand U1772 (N_1772,N_998,N_880);
nand U1773 (N_1773,N_596,N_37);
and U1774 (N_1774,N_269,N_371);
and U1775 (N_1775,N_550,N_637);
or U1776 (N_1776,N_539,N_869);
or U1777 (N_1777,N_572,N_66);
nand U1778 (N_1778,N_617,N_568);
or U1779 (N_1779,N_766,N_957);
and U1780 (N_1780,N_394,N_7);
and U1781 (N_1781,N_9,N_209);
and U1782 (N_1782,N_592,N_22);
or U1783 (N_1783,N_62,N_540);
nor U1784 (N_1784,N_599,N_409);
and U1785 (N_1785,N_409,N_960);
or U1786 (N_1786,N_968,N_122);
nor U1787 (N_1787,N_571,N_484);
nor U1788 (N_1788,N_734,N_532);
nor U1789 (N_1789,N_117,N_661);
nand U1790 (N_1790,N_955,N_202);
or U1791 (N_1791,N_358,N_637);
nor U1792 (N_1792,N_768,N_282);
or U1793 (N_1793,N_502,N_422);
and U1794 (N_1794,N_858,N_573);
nor U1795 (N_1795,N_331,N_304);
and U1796 (N_1796,N_884,N_814);
nand U1797 (N_1797,N_688,N_794);
nand U1798 (N_1798,N_26,N_397);
nand U1799 (N_1799,N_345,N_370);
nand U1800 (N_1800,N_761,N_461);
nor U1801 (N_1801,N_779,N_182);
or U1802 (N_1802,N_396,N_68);
and U1803 (N_1803,N_784,N_59);
or U1804 (N_1804,N_455,N_521);
and U1805 (N_1805,N_4,N_97);
nand U1806 (N_1806,N_765,N_975);
or U1807 (N_1807,N_817,N_218);
nand U1808 (N_1808,N_770,N_793);
and U1809 (N_1809,N_721,N_460);
nor U1810 (N_1810,N_686,N_105);
and U1811 (N_1811,N_816,N_715);
nor U1812 (N_1812,N_201,N_842);
and U1813 (N_1813,N_542,N_993);
or U1814 (N_1814,N_247,N_129);
nand U1815 (N_1815,N_143,N_674);
nor U1816 (N_1816,N_714,N_431);
or U1817 (N_1817,N_430,N_720);
or U1818 (N_1818,N_118,N_378);
and U1819 (N_1819,N_54,N_200);
or U1820 (N_1820,N_875,N_453);
or U1821 (N_1821,N_833,N_800);
and U1822 (N_1822,N_799,N_121);
nand U1823 (N_1823,N_322,N_274);
or U1824 (N_1824,N_174,N_680);
nand U1825 (N_1825,N_892,N_747);
nor U1826 (N_1826,N_273,N_226);
or U1827 (N_1827,N_556,N_840);
and U1828 (N_1828,N_991,N_584);
nor U1829 (N_1829,N_510,N_241);
nor U1830 (N_1830,N_721,N_561);
or U1831 (N_1831,N_387,N_684);
or U1832 (N_1832,N_98,N_367);
or U1833 (N_1833,N_510,N_571);
and U1834 (N_1834,N_220,N_226);
nand U1835 (N_1835,N_251,N_431);
nor U1836 (N_1836,N_20,N_734);
and U1837 (N_1837,N_309,N_743);
nor U1838 (N_1838,N_964,N_384);
and U1839 (N_1839,N_516,N_115);
nor U1840 (N_1840,N_16,N_837);
or U1841 (N_1841,N_245,N_87);
or U1842 (N_1842,N_315,N_300);
or U1843 (N_1843,N_346,N_510);
nor U1844 (N_1844,N_415,N_662);
nor U1845 (N_1845,N_858,N_231);
nand U1846 (N_1846,N_328,N_919);
and U1847 (N_1847,N_611,N_26);
nor U1848 (N_1848,N_338,N_991);
nor U1849 (N_1849,N_322,N_224);
nand U1850 (N_1850,N_24,N_227);
nand U1851 (N_1851,N_226,N_413);
or U1852 (N_1852,N_856,N_502);
and U1853 (N_1853,N_516,N_688);
nand U1854 (N_1854,N_692,N_645);
nand U1855 (N_1855,N_310,N_742);
or U1856 (N_1856,N_317,N_447);
or U1857 (N_1857,N_699,N_588);
nor U1858 (N_1858,N_791,N_968);
nor U1859 (N_1859,N_198,N_433);
or U1860 (N_1860,N_969,N_402);
nor U1861 (N_1861,N_321,N_747);
nor U1862 (N_1862,N_671,N_968);
or U1863 (N_1863,N_943,N_762);
nand U1864 (N_1864,N_395,N_965);
nor U1865 (N_1865,N_847,N_38);
nand U1866 (N_1866,N_303,N_291);
nor U1867 (N_1867,N_453,N_212);
nor U1868 (N_1868,N_44,N_740);
nand U1869 (N_1869,N_282,N_860);
or U1870 (N_1870,N_520,N_879);
and U1871 (N_1871,N_152,N_938);
nor U1872 (N_1872,N_522,N_895);
or U1873 (N_1873,N_984,N_755);
and U1874 (N_1874,N_944,N_499);
or U1875 (N_1875,N_773,N_816);
or U1876 (N_1876,N_502,N_108);
nand U1877 (N_1877,N_176,N_98);
nand U1878 (N_1878,N_369,N_301);
and U1879 (N_1879,N_575,N_50);
nand U1880 (N_1880,N_133,N_820);
or U1881 (N_1881,N_544,N_134);
or U1882 (N_1882,N_796,N_212);
or U1883 (N_1883,N_28,N_997);
or U1884 (N_1884,N_15,N_849);
or U1885 (N_1885,N_386,N_201);
nand U1886 (N_1886,N_146,N_238);
nor U1887 (N_1887,N_242,N_433);
and U1888 (N_1888,N_856,N_63);
or U1889 (N_1889,N_350,N_611);
nor U1890 (N_1890,N_115,N_991);
and U1891 (N_1891,N_768,N_588);
or U1892 (N_1892,N_586,N_428);
nand U1893 (N_1893,N_91,N_735);
nand U1894 (N_1894,N_981,N_168);
nor U1895 (N_1895,N_919,N_51);
and U1896 (N_1896,N_807,N_9);
and U1897 (N_1897,N_165,N_895);
and U1898 (N_1898,N_234,N_762);
and U1899 (N_1899,N_912,N_340);
nand U1900 (N_1900,N_233,N_105);
nor U1901 (N_1901,N_264,N_774);
and U1902 (N_1902,N_901,N_179);
or U1903 (N_1903,N_326,N_790);
nor U1904 (N_1904,N_710,N_625);
or U1905 (N_1905,N_64,N_302);
or U1906 (N_1906,N_573,N_650);
nand U1907 (N_1907,N_686,N_320);
nand U1908 (N_1908,N_352,N_918);
or U1909 (N_1909,N_770,N_622);
or U1910 (N_1910,N_814,N_502);
and U1911 (N_1911,N_563,N_39);
or U1912 (N_1912,N_934,N_116);
nor U1913 (N_1913,N_373,N_450);
and U1914 (N_1914,N_939,N_583);
nor U1915 (N_1915,N_157,N_139);
or U1916 (N_1916,N_325,N_160);
nor U1917 (N_1917,N_357,N_628);
nand U1918 (N_1918,N_347,N_92);
or U1919 (N_1919,N_508,N_126);
or U1920 (N_1920,N_114,N_348);
and U1921 (N_1921,N_987,N_605);
nand U1922 (N_1922,N_41,N_139);
or U1923 (N_1923,N_86,N_814);
nand U1924 (N_1924,N_931,N_835);
nor U1925 (N_1925,N_224,N_697);
or U1926 (N_1926,N_304,N_251);
or U1927 (N_1927,N_498,N_442);
nor U1928 (N_1928,N_737,N_639);
and U1929 (N_1929,N_131,N_836);
nand U1930 (N_1930,N_488,N_438);
or U1931 (N_1931,N_514,N_803);
and U1932 (N_1932,N_846,N_894);
and U1933 (N_1933,N_997,N_523);
nor U1934 (N_1934,N_48,N_164);
or U1935 (N_1935,N_826,N_713);
and U1936 (N_1936,N_975,N_949);
and U1937 (N_1937,N_695,N_860);
nor U1938 (N_1938,N_860,N_633);
or U1939 (N_1939,N_837,N_447);
and U1940 (N_1940,N_862,N_269);
nor U1941 (N_1941,N_853,N_414);
or U1942 (N_1942,N_320,N_165);
nand U1943 (N_1943,N_631,N_260);
or U1944 (N_1944,N_802,N_561);
or U1945 (N_1945,N_799,N_81);
nand U1946 (N_1946,N_705,N_977);
nand U1947 (N_1947,N_522,N_49);
nand U1948 (N_1948,N_34,N_573);
nor U1949 (N_1949,N_292,N_430);
or U1950 (N_1950,N_951,N_846);
or U1951 (N_1951,N_367,N_938);
nor U1952 (N_1952,N_593,N_525);
and U1953 (N_1953,N_629,N_222);
nor U1954 (N_1954,N_250,N_740);
or U1955 (N_1955,N_747,N_214);
nand U1956 (N_1956,N_977,N_332);
nor U1957 (N_1957,N_168,N_333);
nand U1958 (N_1958,N_722,N_32);
and U1959 (N_1959,N_559,N_469);
nand U1960 (N_1960,N_626,N_257);
or U1961 (N_1961,N_981,N_719);
nor U1962 (N_1962,N_29,N_416);
and U1963 (N_1963,N_967,N_925);
nand U1964 (N_1964,N_942,N_230);
nand U1965 (N_1965,N_142,N_343);
or U1966 (N_1966,N_852,N_4);
and U1967 (N_1967,N_957,N_387);
xnor U1968 (N_1968,N_674,N_828);
or U1969 (N_1969,N_716,N_940);
nand U1970 (N_1970,N_128,N_546);
nand U1971 (N_1971,N_106,N_654);
or U1972 (N_1972,N_374,N_994);
or U1973 (N_1973,N_577,N_950);
nor U1974 (N_1974,N_908,N_267);
nand U1975 (N_1975,N_405,N_331);
nor U1976 (N_1976,N_566,N_462);
nor U1977 (N_1977,N_625,N_188);
or U1978 (N_1978,N_786,N_365);
nand U1979 (N_1979,N_651,N_506);
nand U1980 (N_1980,N_422,N_178);
and U1981 (N_1981,N_355,N_428);
nand U1982 (N_1982,N_934,N_998);
nand U1983 (N_1983,N_833,N_557);
and U1984 (N_1984,N_669,N_277);
and U1985 (N_1985,N_630,N_906);
or U1986 (N_1986,N_699,N_562);
or U1987 (N_1987,N_904,N_192);
nand U1988 (N_1988,N_408,N_63);
or U1989 (N_1989,N_519,N_459);
or U1990 (N_1990,N_595,N_952);
nor U1991 (N_1991,N_320,N_680);
nor U1992 (N_1992,N_247,N_108);
and U1993 (N_1993,N_544,N_759);
and U1994 (N_1994,N_860,N_606);
or U1995 (N_1995,N_407,N_927);
nor U1996 (N_1996,N_230,N_947);
nor U1997 (N_1997,N_231,N_775);
nand U1998 (N_1998,N_897,N_621);
xnor U1999 (N_1999,N_621,N_195);
nand U2000 (N_2000,N_1878,N_1656);
nand U2001 (N_2001,N_1196,N_1508);
xor U2002 (N_2002,N_1359,N_1502);
or U2003 (N_2003,N_1651,N_1608);
and U2004 (N_2004,N_1420,N_1436);
and U2005 (N_2005,N_1860,N_1473);
or U2006 (N_2006,N_1496,N_1354);
nor U2007 (N_2007,N_1298,N_1648);
and U2008 (N_2008,N_1754,N_1184);
or U2009 (N_2009,N_1564,N_1636);
and U2010 (N_2010,N_1816,N_1692);
nor U2011 (N_2011,N_1060,N_1227);
or U2012 (N_2012,N_1598,N_1269);
and U2013 (N_2013,N_1264,N_1961);
and U2014 (N_2014,N_1852,N_1945);
nor U2015 (N_2015,N_1101,N_1193);
nand U2016 (N_2016,N_1325,N_1090);
nand U2017 (N_2017,N_1019,N_1405);
or U2018 (N_2018,N_1821,N_1875);
nand U2019 (N_2019,N_1952,N_1590);
nand U2020 (N_2020,N_1086,N_1803);
and U2021 (N_2021,N_1880,N_1288);
nor U2022 (N_2022,N_1503,N_1977);
nor U2023 (N_2023,N_1332,N_1638);
or U2024 (N_2024,N_1318,N_1383);
nor U2025 (N_2025,N_1888,N_1222);
or U2026 (N_2026,N_1963,N_1770);
nand U2027 (N_2027,N_1307,N_1218);
or U2028 (N_2028,N_1480,N_1046);
nand U2029 (N_2029,N_1825,N_1246);
and U2030 (N_2030,N_1725,N_1824);
nand U2031 (N_2031,N_1815,N_1080);
nand U2032 (N_2032,N_1478,N_1919);
or U2033 (N_2033,N_1204,N_1512);
nor U2034 (N_2034,N_1263,N_1698);
and U2035 (N_2035,N_1402,N_1516);
nand U2036 (N_2036,N_1882,N_1289);
nor U2037 (N_2037,N_1450,N_1347);
nand U2038 (N_2038,N_1615,N_1546);
and U2039 (N_2039,N_1886,N_1419);
nor U2040 (N_2040,N_1772,N_1645);
nor U2041 (N_2041,N_1905,N_1000);
nor U2042 (N_2042,N_1774,N_1364);
nand U2043 (N_2043,N_1790,N_1997);
or U2044 (N_2044,N_1274,N_1303);
nor U2045 (N_2045,N_1600,N_1804);
xnor U2046 (N_2046,N_1545,N_1317);
and U2047 (N_2047,N_1808,N_1858);
nor U2048 (N_2048,N_1538,N_1747);
or U2049 (N_2049,N_1655,N_1437);
or U2050 (N_2050,N_1262,N_1641);
or U2051 (N_2051,N_1105,N_1744);
or U2052 (N_2052,N_1896,N_1031);
nor U2053 (N_2053,N_1191,N_1443);
and U2054 (N_2054,N_1434,N_1849);
or U2055 (N_2055,N_1374,N_1211);
nor U2056 (N_2056,N_1843,N_1304);
or U2057 (N_2057,N_1520,N_1074);
nand U2058 (N_2058,N_1728,N_1707);
or U2059 (N_2059,N_1376,N_1687);
nor U2060 (N_2060,N_1397,N_1435);
and U2061 (N_2061,N_1678,N_1382);
and U2062 (N_2062,N_1036,N_1235);
nand U2063 (N_2063,N_1225,N_1577);
nand U2064 (N_2064,N_1894,N_1526);
nor U2065 (N_2065,N_1792,N_1776);
nand U2066 (N_2066,N_1509,N_1898);
nor U2067 (N_2067,N_1007,N_1933);
or U2068 (N_2068,N_1885,N_1216);
nor U2069 (N_2069,N_1938,N_1033);
and U2070 (N_2070,N_1669,N_1029);
nor U2071 (N_2071,N_1291,N_1257);
nor U2072 (N_2072,N_1159,N_1139);
and U2073 (N_2073,N_1275,N_1667);
or U2074 (N_2074,N_1987,N_1908);
and U2075 (N_2075,N_1411,N_1644);
and U2076 (N_2076,N_1985,N_1389);
and U2077 (N_2077,N_1693,N_1884);
or U2078 (N_2078,N_1788,N_1053);
nor U2079 (N_2079,N_1125,N_1926);
or U2080 (N_2080,N_1034,N_1699);
nor U2081 (N_2081,N_1702,N_1284);
nor U2082 (N_2082,N_1872,N_1056);
nand U2083 (N_2083,N_1642,N_1144);
nor U2084 (N_2084,N_1927,N_1628);
nor U2085 (N_2085,N_1170,N_1633);
nor U2086 (N_2086,N_1188,N_1988);
and U2087 (N_2087,N_1458,N_1990);
nand U2088 (N_2088,N_1481,N_1757);
and U2089 (N_2089,N_1614,N_1617);
nor U2090 (N_2090,N_1517,N_1783);
and U2091 (N_2091,N_1940,N_1260);
nand U2092 (N_2092,N_1521,N_1560);
nor U2093 (N_2093,N_1212,N_1616);
nor U2094 (N_2094,N_1850,N_1575);
nand U2095 (N_2095,N_1349,N_1070);
nand U2096 (N_2096,N_1603,N_1553);
nand U2097 (N_2097,N_1375,N_1114);
nand U2098 (N_2098,N_1008,N_1604);
and U2099 (N_2099,N_1394,N_1181);
nand U2100 (N_2100,N_1705,N_1043);
and U2101 (N_2101,N_1918,N_1812);
nor U2102 (N_2102,N_1021,N_1069);
nor U2103 (N_2103,N_1955,N_1336);
nand U2104 (N_2104,N_1365,N_1947);
nor U2105 (N_2105,N_1543,N_1594);
nor U2106 (N_2106,N_1838,N_1483);
nor U2107 (N_2107,N_1539,N_1513);
nand U2108 (N_2108,N_1555,N_1833);
nor U2109 (N_2109,N_1559,N_1097);
and U2110 (N_2110,N_1281,N_1240);
nor U2111 (N_2111,N_1809,N_1460);
or U2112 (N_2112,N_1567,N_1746);
and U2113 (N_2113,N_1388,N_1652);
xnor U2114 (N_2114,N_1675,N_1384);
and U2115 (N_2115,N_1495,N_1529);
and U2116 (N_2116,N_1499,N_1295);
nand U2117 (N_2117,N_1012,N_1883);
or U2118 (N_2118,N_1920,N_1206);
or U2119 (N_2119,N_1620,N_1253);
or U2120 (N_2120,N_1208,N_1826);
and U2121 (N_2121,N_1906,N_1874);
and U2122 (N_2122,N_1362,N_1452);
nand U2123 (N_2123,N_1367,N_1950);
or U2124 (N_2124,N_1528,N_1805);
or U2125 (N_2125,N_1445,N_1971);
and U2126 (N_2126,N_1418,N_1856);
nor U2127 (N_2127,N_1680,N_1148);
and U2128 (N_2128,N_1429,N_1924);
or U2129 (N_2129,N_1368,N_1041);
or U2130 (N_2130,N_1037,N_1022);
xor U2131 (N_2131,N_1581,N_1161);
and U2132 (N_2132,N_1976,N_1631);
and U2133 (N_2133,N_1504,N_1082);
and U2134 (N_2134,N_1271,N_1781);
and U2135 (N_2135,N_1200,N_1876);
or U2136 (N_2136,N_1864,N_1109);
or U2137 (N_2137,N_1845,N_1356);
nand U2138 (N_2138,N_1568,N_1634);
nand U2139 (N_2139,N_1166,N_1565);
nand U2140 (N_2140,N_1627,N_1203);
or U2141 (N_2141,N_1960,N_1015);
or U2142 (N_2142,N_1727,N_1459);
nor U2143 (N_2143,N_1255,N_1925);
or U2144 (N_2144,N_1083,N_1002);
or U2145 (N_2145,N_1348,N_1327);
xor U2146 (N_2146,N_1266,N_1709);
nor U2147 (N_2147,N_1602,N_1914);
nor U2148 (N_2148,N_1563,N_1811);
nor U2149 (N_2149,N_1039,N_1424);
nor U2150 (N_2150,N_1229,N_1004);
nor U2151 (N_2151,N_1593,N_1723);
nand U2152 (N_2152,N_1487,N_1629);
and U2153 (N_2153,N_1351,N_1357);
nor U2154 (N_2154,N_1731,N_1350);
or U2155 (N_2155,N_1448,N_1066);
nand U2156 (N_2156,N_1686,N_1237);
nor U2157 (N_2157,N_1476,N_1361);
or U2158 (N_2158,N_1238,N_1230);
or U2159 (N_2159,N_1055,N_1551);
nand U2160 (N_2160,N_1928,N_1154);
nor U2161 (N_2161,N_1179,N_1975);
nand U2162 (N_2162,N_1566,N_1574);
and U2163 (N_2163,N_1189,N_1653);
or U2164 (N_2164,N_1778,N_1959);
or U2165 (N_2165,N_1265,N_1329);
nor U2166 (N_2166,N_1016,N_1897);
nand U2167 (N_2167,N_1078,N_1991);
or U2168 (N_2168,N_1416,N_1130);
or U2169 (N_2169,N_1335,N_1044);
or U2170 (N_2170,N_1057,N_1978);
or U2171 (N_2171,N_1548,N_1916);
and U2172 (N_2172,N_1717,N_1659);
and U2173 (N_2173,N_1489,N_1939);
nand U2174 (N_2174,N_1252,N_1587);
or U2175 (N_2175,N_1254,N_1923);
nand U2176 (N_2176,N_1626,N_1311);
nand U2177 (N_2177,N_1020,N_1589);
nand U2178 (N_2178,N_1537,N_1672);
or U2179 (N_2179,N_1447,N_1197);
and U2180 (N_2180,N_1911,N_1092);
and U2181 (N_2181,N_1187,N_1358);
nor U2182 (N_2182,N_1535,N_1980);
or U2183 (N_2183,N_1115,N_1721);
nor U2184 (N_2184,N_1180,N_1391);
nand U2185 (N_2185,N_1554,N_1091);
nand U2186 (N_2186,N_1138,N_1312);
or U2187 (N_2187,N_1724,N_1276);
or U2188 (N_2188,N_1773,N_1970);
nor U2189 (N_2189,N_1839,N_1400);
or U2190 (N_2190,N_1323,N_1477);
nand U2191 (N_2191,N_1527,N_1640);
and U2192 (N_2192,N_1127,N_1456);
nand U2193 (N_2193,N_1423,N_1028);
nand U2194 (N_2194,N_1433,N_1734);
nor U2195 (N_2195,N_1088,N_1992);
and U2196 (N_2196,N_1832,N_1837);
nor U2197 (N_2197,N_1401,N_1396);
or U2198 (N_2198,N_1395,N_1155);
nand U2199 (N_2199,N_1026,N_1782);
or U2200 (N_2200,N_1474,N_1464);
nand U2201 (N_2201,N_1339,N_1689);
or U2202 (N_2202,N_1904,N_1344);
nand U2203 (N_2203,N_1279,N_1964);
or U2204 (N_2204,N_1226,N_1704);
nand U2205 (N_2205,N_1326,N_1547);
or U2206 (N_2206,N_1922,N_1099);
nand U2207 (N_2207,N_1870,N_1573);
nor U2208 (N_2208,N_1338,N_1612);
or U2209 (N_2209,N_1597,N_1160);
nor U2210 (N_2210,N_1169,N_1890);
and U2211 (N_2211,N_1643,N_1540);
nor U2212 (N_2212,N_1061,N_1588);
or U2213 (N_2213,N_1868,N_1544);
nor U2214 (N_2214,N_1111,N_1306);
and U2215 (N_2215,N_1340,N_1465);
and U2216 (N_2216,N_1277,N_1846);
nand U2217 (N_2217,N_1713,N_1469);
nand U2218 (N_2218,N_1741,N_1557);
nor U2219 (N_2219,N_1984,N_1194);
or U2220 (N_2220,N_1393,N_1468);
nor U2221 (N_2221,N_1231,N_1268);
nand U2222 (N_2222,N_1836,N_1664);
or U2223 (N_2223,N_1484,N_1714);
and U2224 (N_2224,N_1830,N_1671);
nor U2225 (N_2225,N_1045,N_1417);
and U2226 (N_2226,N_1979,N_1601);
or U2227 (N_2227,N_1135,N_1162);
nor U2228 (N_2228,N_1425,N_1488);
or U2229 (N_2229,N_1625,N_1822);
nand U2230 (N_2230,N_1446,N_1862);
nor U2231 (N_2231,N_1583,N_1690);
or U2232 (N_2232,N_1942,N_1766);
and U2233 (N_2233,N_1847,N_1570);
or U2234 (N_2234,N_1534,N_1851);
and U2235 (N_2235,N_1280,N_1228);
and U2236 (N_2236,N_1110,N_1415);
nor U2237 (N_2237,N_1639,N_1763);
nor U2238 (N_2238,N_1813,N_1635);
or U2239 (N_2239,N_1974,N_1657);
nand U2240 (N_2240,N_1827,N_1605);
and U2241 (N_2241,N_1380,N_1006);
nor U2242 (N_2242,N_1378,N_1879);
and U2243 (N_2243,N_1682,N_1047);
or U2244 (N_2244,N_1752,N_1571);
and U2245 (N_2245,N_1491,N_1059);
and U2246 (N_2246,N_1192,N_1100);
nor U2247 (N_2247,N_1030,N_1956);
or U2248 (N_2248,N_1715,N_1751);
or U2249 (N_2249,N_1261,N_1842);
and U2250 (N_2250,N_1243,N_1806);
nand U2251 (N_2251,N_1523,N_1462);
nand U2252 (N_2252,N_1595,N_1498);
nand U2253 (N_2253,N_1077,N_1024);
nor U2254 (N_2254,N_1996,N_1929);
and U2255 (N_2255,N_1305,N_1319);
and U2256 (N_2256,N_1172,N_1764);
nor U2257 (N_2257,N_1234,N_1067);
nand U2258 (N_2258,N_1322,N_1663);
nand U2259 (N_2259,N_1691,N_1129);
and U2260 (N_2260,N_1132,N_1103);
and U2261 (N_2261,N_1313,N_1820);
nand U2262 (N_2262,N_1013,N_1666);
nor U2263 (N_2263,N_1454,N_1869);
nor U2264 (N_2264,N_1893,N_1490);
nor U2265 (N_2265,N_1861,N_1748);
xnor U2266 (N_2266,N_1217,N_1958);
or U2267 (N_2267,N_1835,N_1081);
nor U2268 (N_2268,N_1387,N_1683);
nor U2269 (N_2269,N_1844,N_1133);
nor U2270 (N_2270,N_1178,N_1320);
nor U2271 (N_2271,N_1937,N_1579);
and U2272 (N_2272,N_1867,N_1301);
nand U2273 (N_2273,N_1592,N_1510);
or U2274 (N_2274,N_1729,N_1710);
nand U2275 (N_2275,N_1780,N_1439);
nor U2276 (N_2276,N_1983,N_1558);
nand U2277 (N_2277,N_1834,N_1493);
xnor U2278 (N_2278,N_1441,N_1141);
nand U2279 (N_2279,N_1749,N_1726);
and U2280 (N_2280,N_1104,N_1250);
nor U2281 (N_2281,N_1119,N_1001);
and U2282 (N_2282,N_1116,N_1973);
nor U2283 (N_2283,N_1241,N_1999);
nand U2284 (N_2284,N_1112,N_1599);
or U2285 (N_2285,N_1126,N_1471);
nor U2286 (N_2286,N_1063,N_1466);
or U2287 (N_2287,N_1084,N_1165);
nand U2288 (N_2288,N_1409,N_1118);
and U2289 (N_2289,N_1143,N_1913);
and U2290 (N_2290,N_1158,N_1944);
or U2291 (N_2291,N_1005,N_1174);
nand U2292 (N_2292,N_1124,N_1224);
and U2293 (N_2293,N_1505,N_1533);
or U2294 (N_2294,N_1106,N_1068);
nand U2295 (N_2295,N_1292,N_1333);
nor U2296 (N_2296,N_1814,N_1841);
and U2297 (N_2297,N_1765,N_1685);
nand U2298 (N_2298,N_1302,N_1343);
nor U2299 (N_2299,N_1981,N_1128);
nand U2300 (N_2300,N_1580,N_1379);
or U2301 (N_2301,N_1096,N_1398);
nor U2302 (N_2302,N_1661,N_1802);
or U2303 (N_2303,N_1982,N_1895);
or U2304 (N_2304,N_1223,N_1247);
nand U2305 (N_2305,N_1522,N_1799);
nand U2306 (N_2306,N_1995,N_1785);
nand U2307 (N_2307,N_1931,N_1900);
nand U2308 (N_2308,N_1968,N_1486);
nand U2309 (N_2309,N_1965,N_1541);
or U2310 (N_2310,N_1742,N_1048);
or U2311 (N_2311,N_1051,N_1524);
nand U2312 (N_2312,N_1854,N_1736);
nand U2313 (N_2313,N_1817,N_1737);
or U2314 (N_2314,N_1946,N_1278);
and U2315 (N_2315,N_1199,N_1768);
nor U2316 (N_2316,N_1531,N_1511);
nor U2317 (N_2317,N_1403,N_1113);
and U2318 (N_2318,N_1556,N_1810);
nand U2319 (N_2319,N_1695,N_1214);
nor U2320 (N_2320,N_1286,N_1801);
or U2321 (N_2321,N_1514,N_1346);
nor U2322 (N_2322,N_1136,N_1142);
nand U2323 (N_2323,N_1032,N_1360);
nand U2324 (N_2324,N_1621,N_1296);
nor U2325 (N_2325,N_1703,N_1102);
and U2326 (N_2326,N_1935,N_1903);
nand U2327 (N_2327,N_1094,N_1371);
and U2328 (N_2328,N_1892,N_1930);
and U2329 (N_2329,N_1315,N_1011);
and U2330 (N_2330,N_1795,N_1202);
and U2331 (N_2331,N_1290,N_1185);
and U2332 (N_2332,N_1316,N_1023);
and U2333 (N_2333,N_1245,N_1087);
nor U2334 (N_2334,N_1299,N_1168);
nand U2335 (N_2335,N_1233,N_1921);
nor U2336 (N_2336,N_1107,N_1966);
nand U2337 (N_2337,N_1532,N_1151);
or U2338 (N_2338,N_1025,N_1712);
nand U2339 (N_2339,N_1767,N_1406);
or U2340 (N_2340,N_1793,N_1248);
or U2341 (N_2341,N_1120,N_1584);
nand U2342 (N_2342,N_1507,N_1891);
or U2343 (N_2343,N_1700,N_1609);
nand U2344 (N_2344,N_1670,N_1515);
and U2345 (N_2345,N_1866,N_1071);
nor U2346 (N_2346,N_1632,N_1463);
and U2347 (N_2347,N_1221,N_1058);
nand U2348 (N_2348,N_1285,N_1807);
nor U2349 (N_2349,N_1085,N_1889);
or U2350 (N_2350,N_1732,N_1236);
or U2351 (N_2351,N_1831,N_1220);
and U2352 (N_2352,N_1542,N_1800);
or U2353 (N_2353,N_1986,N_1345);
nor U2354 (N_2354,N_1777,N_1967);
or U2355 (N_2355,N_1915,N_1475);
and U2356 (N_2356,N_1381,N_1887);
nand U2357 (N_2357,N_1328,N_1209);
or U2358 (N_2358,N_1840,N_1561);
nand U2359 (N_2359,N_1582,N_1146);
nor U2360 (N_2360,N_1989,N_1948);
or U2361 (N_2361,N_1485,N_1525);
and U2362 (N_2362,N_1720,N_1334);
and U2363 (N_2363,N_1342,N_1674);
and U2364 (N_2364,N_1569,N_1470);
nor U2365 (N_2365,N_1009,N_1073);
nor U2366 (N_2366,N_1941,N_1753);
or U2367 (N_2367,N_1062,N_1684);
nand U2368 (N_2368,N_1242,N_1038);
or U2369 (N_2369,N_1859,N_1137);
and U2370 (N_2370,N_1760,N_1372);
nand U2371 (N_2371,N_1994,N_1413);
nand U2372 (N_2372,N_1164,N_1273);
or U2373 (N_2373,N_1186,N_1064);
or U2374 (N_2374,N_1797,N_1075);
nor U2375 (N_2375,N_1630,N_1018);
nor U2376 (N_2376,N_1701,N_1606);
nor U2377 (N_2377,N_1738,N_1855);
or U2378 (N_2378,N_1530,N_1549);
nand U2379 (N_2379,N_1453,N_1457);
nor U2380 (N_2380,N_1121,N_1743);
and U2381 (N_2381,N_1877,N_1972);
nor U2382 (N_2382,N_1205,N_1618);
or U2383 (N_2383,N_1412,N_1562);
nand U2384 (N_2384,N_1596,N_1093);
and U2385 (N_2385,N_1818,N_1750);
or U2386 (N_2386,N_1198,N_1789);
nor U2387 (N_2387,N_1215,N_1494);
nand U2388 (N_2388,N_1210,N_1251);
or U2389 (N_2389,N_1873,N_1035);
or U2390 (N_2390,N_1761,N_1003);
nand U2391 (N_2391,N_1366,N_1676);
nand U2392 (N_2392,N_1385,N_1182);
nor U2393 (N_2393,N_1177,N_1798);
or U2394 (N_2394,N_1518,N_1871);
nor U2395 (N_2395,N_1969,N_1500);
nor U2396 (N_2396,N_1054,N_1607);
nand U2397 (N_2397,N_1149,N_1098);
nor U2398 (N_2398,N_1176,N_1730);
nor U2399 (N_2399,N_1014,N_1679);
or U2400 (N_2400,N_1167,N_1479);
or U2401 (N_2401,N_1771,N_1330);
and U2402 (N_2402,N_1267,N_1232);
or U2403 (N_2403,N_1190,N_1147);
or U2404 (N_2404,N_1951,N_1440);
or U2405 (N_2405,N_1455,N_1694);
nor U2406 (N_2406,N_1353,N_1272);
or U2407 (N_2407,N_1337,N_1932);
and U2408 (N_2408,N_1769,N_1213);
xor U2409 (N_2409,N_1936,N_1708);
and U2410 (N_2410,N_1668,N_1451);
nand U2411 (N_2411,N_1646,N_1623);
nand U2412 (N_2412,N_1404,N_1239);
or U2413 (N_2413,N_1585,N_1722);
and U2414 (N_2414,N_1718,N_1259);
or U2415 (N_2415,N_1786,N_1444);
and U2416 (N_2416,N_1917,N_1027);
or U2417 (N_2417,N_1076,N_1355);
and U2418 (N_2418,N_1909,N_1681);
or U2419 (N_2419,N_1943,N_1300);
nor U2420 (N_2420,N_1249,N_1195);
nand U2421 (N_2421,N_1576,N_1591);
nor U2422 (N_2422,N_1461,N_1962);
or U2423 (N_2423,N_1117,N_1331);
nor U2424 (N_2424,N_1369,N_1392);
nand U2425 (N_2425,N_1953,N_1497);
nand U2426 (N_2426,N_1658,N_1421);
nand U2427 (N_2427,N_1711,N_1550);
or U2428 (N_2428,N_1791,N_1153);
nor U2429 (N_2429,N_1156,N_1370);
or U2430 (N_2430,N_1430,N_1293);
and U2431 (N_2431,N_1706,N_1145);
nand U2432 (N_2432,N_1201,N_1183);
and U2433 (N_2433,N_1501,N_1449);
or U2434 (N_2434,N_1719,N_1716);
and U2435 (N_2435,N_1432,N_1673);
and U2436 (N_2436,N_1677,N_1899);
and U2437 (N_2437,N_1095,N_1175);
and U2438 (N_2438,N_1089,N_1779);
or U2439 (N_2439,N_1794,N_1775);
nor U2440 (N_2440,N_1324,N_1756);
nand U2441 (N_2441,N_1954,N_1442);
nand U2442 (N_2442,N_1613,N_1622);
nor U2443 (N_2443,N_1363,N_1050);
or U2444 (N_2444,N_1049,N_1310);
nor U2445 (N_2445,N_1649,N_1152);
nor U2446 (N_2446,N_1270,N_1482);
and U2447 (N_2447,N_1745,N_1377);
or U2448 (N_2448,N_1647,N_1863);
nor U2449 (N_2449,N_1157,N_1386);
nand U2450 (N_2450,N_1244,N_1637);
and U2451 (N_2451,N_1428,N_1438);
or U2452 (N_2452,N_1796,N_1578);
and U2453 (N_2453,N_1688,N_1910);
or U2454 (N_2454,N_1912,N_1163);
nand U2455 (N_2455,N_1065,N_1733);
nand U2456 (N_2456,N_1427,N_1407);
or U2457 (N_2457,N_1572,N_1173);
nor U2458 (N_2458,N_1399,N_1219);
and U2459 (N_2459,N_1762,N_1993);
and U2460 (N_2460,N_1823,N_1848);
nand U2461 (N_2461,N_1611,N_1901);
and U2462 (N_2462,N_1735,N_1258);
nand U2463 (N_2463,N_1373,N_1828);
nand U2464 (N_2464,N_1853,N_1294);
and U2465 (N_2465,N_1414,N_1739);
and U2466 (N_2466,N_1787,N_1408);
and U2467 (N_2467,N_1134,N_1536);
and U2468 (N_2468,N_1759,N_1662);
or U2469 (N_2469,N_1740,N_1131);
nor U2470 (N_2470,N_1431,N_1472);
nand U2471 (N_2471,N_1314,N_1697);
xnor U2472 (N_2472,N_1321,N_1422);
or U2473 (N_2473,N_1610,N_1410);
nor U2474 (N_2474,N_1052,N_1758);
nand U2475 (N_2475,N_1949,N_1857);
and U2476 (N_2476,N_1829,N_1506);
or U2477 (N_2477,N_1072,N_1308);
nand U2478 (N_2478,N_1123,N_1934);
and U2479 (N_2479,N_1171,N_1696);
or U2480 (N_2480,N_1309,N_1040);
nand U2481 (N_2481,N_1665,N_1819);
and U2482 (N_2482,N_1017,N_1957);
nand U2483 (N_2483,N_1755,N_1390);
nor U2484 (N_2484,N_1650,N_1624);
and U2485 (N_2485,N_1660,N_1492);
and U2486 (N_2486,N_1150,N_1256);
or U2487 (N_2487,N_1519,N_1207);
nor U2488 (N_2488,N_1654,N_1586);
or U2489 (N_2489,N_1140,N_1283);
nand U2490 (N_2490,N_1297,N_1865);
and U2491 (N_2491,N_1467,N_1122);
nand U2492 (N_2492,N_1010,N_1784);
and U2493 (N_2493,N_1282,N_1881);
or U2494 (N_2494,N_1108,N_1552);
nand U2495 (N_2495,N_1287,N_1998);
and U2496 (N_2496,N_1079,N_1902);
and U2497 (N_2497,N_1619,N_1042);
and U2498 (N_2498,N_1341,N_1352);
or U2499 (N_2499,N_1907,N_1426);
or U2500 (N_2500,N_1668,N_1918);
nand U2501 (N_2501,N_1823,N_1811);
and U2502 (N_2502,N_1268,N_1261);
nor U2503 (N_2503,N_1071,N_1321);
or U2504 (N_2504,N_1037,N_1964);
nand U2505 (N_2505,N_1954,N_1792);
nor U2506 (N_2506,N_1527,N_1849);
or U2507 (N_2507,N_1568,N_1435);
or U2508 (N_2508,N_1260,N_1724);
nor U2509 (N_2509,N_1291,N_1444);
or U2510 (N_2510,N_1512,N_1388);
nand U2511 (N_2511,N_1468,N_1016);
nor U2512 (N_2512,N_1014,N_1503);
or U2513 (N_2513,N_1506,N_1348);
or U2514 (N_2514,N_1924,N_1016);
xnor U2515 (N_2515,N_1908,N_1014);
and U2516 (N_2516,N_1378,N_1264);
nand U2517 (N_2517,N_1662,N_1520);
nand U2518 (N_2518,N_1150,N_1290);
and U2519 (N_2519,N_1320,N_1296);
nand U2520 (N_2520,N_1618,N_1299);
or U2521 (N_2521,N_1082,N_1045);
or U2522 (N_2522,N_1433,N_1798);
nor U2523 (N_2523,N_1421,N_1633);
and U2524 (N_2524,N_1965,N_1572);
and U2525 (N_2525,N_1604,N_1044);
nand U2526 (N_2526,N_1984,N_1384);
nand U2527 (N_2527,N_1807,N_1731);
and U2528 (N_2528,N_1066,N_1992);
nand U2529 (N_2529,N_1904,N_1974);
or U2530 (N_2530,N_1339,N_1892);
nand U2531 (N_2531,N_1320,N_1310);
nand U2532 (N_2532,N_1281,N_1742);
nor U2533 (N_2533,N_1605,N_1696);
or U2534 (N_2534,N_1987,N_1460);
nor U2535 (N_2535,N_1660,N_1292);
nand U2536 (N_2536,N_1113,N_1402);
or U2537 (N_2537,N_1528,N_1096);
and U2538 (N_2538,N_1864,N_1100);
or U2539 (N_2539,N_1660,N_1608);
nand U2540 (N_2540,N_1941,N_1310);
nand U2541 (N_2541,N_1198,N_1018);
nand U2542 (N_2542,N_1131,N_1400);
and U2543 (N_2543,N_1462,N_1855);
or U2544 (N_2544,N_1738,N_1453);
and U2545 (N_2545,N_1886,N_1855);
and U2546 (N_2546,N_1350,N_1347);
or U2547 (N_2547,N_1255,N_1199);
or U2548 (N_2548,N_1968,N_1477);
or U2549 (N_2549,N_1121,N_1816);
or U2550 (N_2550,N_1070,N_1438);
nor U2551 (N_2551,N_1970,N_1686);
nand U2552 (N_2552,N_1868,N_1852);
or U2553 (N_2553,N_1494,N_1834);
nor U2554 (N_2554,N_1082,N_1789);
or U2555 (N_2555,N_1475,N_1389);
or U2556 (N_2556,N_1940,N_1085);
nand U2557 (N_2557,N_1336,N_1886);
xnor U2558 (N_2558,N_1625,N_1366);
and U2559 (N_2559,N_1123,N_1755);
nor U2560 (N_2560,N_1846,N_1555);
and U2561 (N_2561,N_1421,N_1572);
xor U2562 (N_2562,N_1755,N_1776);
nor U2563 (N_2563,N_1172,N_1178);
or U2564 (N_2564,N_1013,N_1817);
nor U2565 (N_2565,N_1082,N_1447);
and U2566 (N_2566,N_1081,N_1441);
or U2567 (N_2567,N_1000,N_1550);
or U2568 (N_2568,N_1877,N_1815);
and U2569 (N_2569,N_1497,N_1060);
nor U2570 (N_2570,N_1331,N_1620);
nand U2571 (N_2571,N_1234,N_1435);
nand U2572 (N_2572,N_1798,N_1755);
nand U2573 (N_2573,N_1140,N_1377);
and U2574 (N_2574,N_1293,N_1756);
nor U2575 (N_2575,N_1392,N_1909);
and U2576 (N_2576,N_1871,N_1747);
and U2577 (N_2577,N_1220,N_1996);
and U2578 (N_2578,N_1334,N_1736);
or U2579 (N_2579,N_1178,N_1131);
and U2580 (N_2580,N_1502,N_1680);
nor U2581 (N_2581,N_1976,N_1441);
and U2582 (N_2582,N_1844,N_1663);
or U2583 (N_2583,N_1898,N_1769);
xnor U2584 (N_2584,N_1915,N_1467);
and U2585 (N_2585,N_1167,N_1800);
and U2586 (N_2586,N_1174,N_1483);
and U2587 (N_2587,N_1014,N_1238);
and U2588 (N_2588,N_1034,N_1921);
nor U2589 (N_2589,N_1939,N_1610);
nand U2590 (N_2590,N_1527,N_1853);
and U2591 (N_2591,N_1490,N_1952);
nor U2592 (N_2592,N_1841,N_1664);
or U2593 (N_2593,N_1950,N_1839);
and U2594 (N_2594,N_1051,N_1681);
nand U2595 (N_2595,N_1067,N_1091);
xnor U2596 (N_2596,N_1292,N_1607);
nand U2597 (N_2597,N_1565,N_1511);
and U2598 (N_2598,N_1926,N_1078);
and U2599 (N_2599,N_1524,N_1250);
or U2600 (N_2600,N_1022,N_1154);
or U2601 (N_2601,N_1111,N_1446);
nor U2602 (N_2602,N_1387,N_1900);
and U2603 (N_2603,N_1480,N_1785);
and U2604 (N_2604,N_1299,N_1791);
nor U2605 (N_2605,N_1491,N_1848);
nand U2606 (N_2606,N_1951,N_1551);
nor U2607 (N_2607,N_1922,N_1325);
nor U2608 (N_2608,N_1157,N_1265);
and U2609 (N_2609,N_1262,N_1705);
nand U2610 (N_2610,N_1425,N_1163);
or U2611 (N_2611,N_1255,N_1960);
and U2612 (N_2612,N_1053,N_1278);
and U2613 (N_2613,N_1854,N_1441);
or U2614 (N_2614,N_1596,N_1021);
nor U2615 (N_2615,N_1033,N_1623);
nand U2616 (N_2616,N_1215,N_1033);
or U2617 (N_2617,N_1344,N_1687);
or U2618 (N_2618,N_1649,N_1334);
or U2619 (N_2619,N_1410,N_1562);
nor U2620 (N_2620,N_1816,N_1549);
or U2621 (N_2621,N_1984,N_1581);
nor U2622 (N_2622,N_1232,N_1887);
nor U2623 (N_2623,N_1353,N_1766);
nor U2624 (N_2624,N_1718,N_1795);
nor U2625 (N_2625,N_1443,N_1860);
and U2626 (N_2626,N_1852,N_1231);
nor U2627 (N_2627,N_1710,N_1174);
and U2628 (N_2628,N_1365,N_1096);
or U2629 (N_2629,N_1195,N_1032);
nor U2630 (N_2630,N_1494,N_1903);
nor U2631 (N_2631,N_1573,N_1721);
nor U2632 (N_2632,N_1996,N_1600);
or U2633 (N_2633,N_1757,N_1919);
or U2634 (N_2634,N_1136,N_1030);
nor U2635 (N_2635,N_1506,N_1522);
and U2636 (N_2636,N_1999,N_1372);
and U2637 (N_2637,N_1905,N_1219);
nor U2638 (N_2638,N_1157,N_1120);
and U2639 (N_2639,N_1174,N_1168);
or U2640 (N_2640,N_1775,N_1160);
or U2641 (N_2641,N_1608,N_1825);
nor U2642 (N_2642,N_1422,N_1416);
and U2643 (N_2643,N_1408,N_1758);
or U2644 (N_2644,N_1263,N_1283);
and U2645 (N_2645,N_1168,N_1731);
or U2646 (N_2646,N_1097,N_1728);
nand U2647 (N_2647,N_1207,N_1358);
nor U2648 (N_2648,N_1097,N_1833);
nand U2649 (N_2649,N_1414,N_1530);
nand U2650 (N_2650,N_1764,N_1669);
nand U2651 (N_2651,N_1412,N_1349);
nor U2652 (N_2652,N_1210,N_1139);
and U2653 (N_2653,N_1025,N_1653);
and U2654 (N_2654,N_1805,N_1384);
or U2655 (N_2655,N_1813,N_1932);
nand U2656 (N_2656,N_1094,N_1492);
or U2657 (N_2657,N_1468,N_1603);
or U2658 (N_2658,N_1030,N_1374);
or U2659 (N_2659,N_1386,N_1927);
nand U2660 (N_2660,N_1417,N_1000);
nor U2661 (N_2661,N_1703,N_1181);
and U2662 (N_2662,N_1423,N_1170);
nand U2663 (N_2663,N_1129,N_1529);
or U2664 (N_2664,N_1378,N_1009);
or U2665 (N_2665,N_1417,N_1904);
xnor U2666 (N_2666,N_1667,N_1726);
and U2667 (N_2667,N_1648,N_1864);
or U2668 (N_2668,N_1627,N_1234);
or U2669 (N_2669,N_1676,N_1582);
nor U2670 (N_2670,N_1519,N_1924);
and U2671 (N_2671,N_1558,N_1769);
and U2672 (N_2672,N_1645,N_1855);
nor U2673 (N_2673,N_1649,N_1273);
nand U2674 (N_2674,N_1441,N_1970);
or U2675 (N_2675,N_1328,N_1444);
or U2676 (N_2676,N_1370,N_1618);
nand U2677 (N_2677,N_1288,N_1512);
nor U2678 (N_2678,N_1469,N_1847);
nand U2679 (N_2679,N_1713,N_1126);
xnor U2680 (N_2680,N_1990,N_1522);
nor U2681 (N_2681,N_1094,N_1681);
nand U2682 (N_2682,N_1812,N_1135);
and U2683 (N_2683,N_1941,N_1169);
or U2684 (N_2684,N_1074,N_1313);
nor U2685 (N_2685,N_1597,N_1603);
or U2686 (N_2686,N_1323,N_1507);
or U2687 (N_2687,N_1495,N_1564);
or U2688 (N_2688,N_1030,N_1854);
or U2689 (N_2689,N_1775,N_1384);
and U2690 (N_2690,N_1424,N_1752);
or U2691 (N_2691,N_1255,N_1204);
nor U2692 (N_2692,N_1394,N_1653);
and U2693 (N_2693,N_1094,N_1459);
nor U2694 (N_2694,N_1220,N_1264);
or U2695 (N_2695,N_1888,N_1549);
or U2696 (N_2696,N_1263,N_1836);
nor U2697 (N_2697,N_1411,N_1814);
nor U2698 (N_2698,N_1090,N_1569);
nand U2699 (N_2699,N_1563,N_1600);
nand U2700 (N_2700,N_1475,N_1580);
and U2701 (N_2701,N_1085,N_1574);
nor U2702 (N_2702,N_1789,N_1126);
or U2703 (N_2703,N_1339,N_1894);
nand U2704 (N_2704,N_1227,N_1287);
nor U2705 (N_2705,N_1000,N_1223);
nor U2706 (N_2706,N_1918,N_1958);
nor U2707 (N_2707,N_1136,N_1554);
nor U2708 (N_2708,N_1230,N_1374);
or U2709 (N_2709,N_1835,N_1323);
nor U2710 (N_2710,N_1902,N_1007);
nor U2711 (N_2711,N_1546,N_1289);
or U2712 (N_2712,N_1332,N_1853);
or U2713 (N_2713,N_1185,N_1798);
nand U2714 (N_2714,N_1633,N_1627);
nand U2715 (N_2715,N_1268,N_1686);
and U2716 (N_2716,N_1956,N_1261);
and U2717 (N_2717,N_1443,N_1942);
and U2718 (N_2718,N_1798,N_1204);
and U2719 (N_2719,N_1321,N_1803);
or U2720 (N_2720,N_1769,N_1986);
nand U2721 (N_2721,N_1999,N_1764);
or U2722 (N_2722,N_1514,N_1707);
and U2723 (N_2723,N_1324,N_1290);
and U2724 (N_2724,N_1176,N_1943);
or U2725 (N_2725,N_1521,N_1412);
nand U2726 (N_2726,N_1630,N_1931);
and U2727 (N_2727,N_1903,N_1604);
nand U2728 (N_2728,N_1179,N_1468);
or U2729 (N_2729,N_1072,N_1456);
nand U2730 (N_2730,N_1646,N_1261);
or U2731 (N_2731,N_1091,N_1459);
nor U2732 (N_2732,N_1920,N_1177);
and U2733 (N_2733,N_1348,N_1343);
nand U2734 (N_2734,N_1777,N_1751);
and U2735 (N_2735,N_1843,N_1298);
and U2736 (N_2736,N_1453,N_1121);
xnor U2737 (N_2737,N_1227,N_1467);
or U2738 (N_2738,N_1946,N_1811);
nor U2739 (N_2739,N_1429,N_1999);
nor U2740 (N_2740,N_1209,N_1020);
and U2741 (N_2741,N_1288,N_1009);
nand U2742 (N_2742,N_1657,N_1726);
nor U2743 (N_2743,N_1652,N_1058);
nor U2744 (N_2744,N_1709,N_1733);
nand U2745 (N_2745,N_1783,N_1342);
nand U2746 (N_2746,N_1587,N_1983);
or U2747 (N_2747,N_1105,N_1430);
nand U2748 (N_2748,N_1099,N_1679);
or U2749 (N_2749,N_1809,N_1589);
and U2750 (N_2750,N_1891,N_1837);
or U2751 (N_2751,N_1008,N_1249);
nand U2752 (N_2752,N_1781,N_1517);
nand U2753 (N_2753,N_1837,N_1381);
or U2754 (N_2754,N_1884,N_1244);
nor U2755 (N_2755,N_1588,N_1051);
or U2756 (N_2756,N_1489,N_1732);
nand U2757 (N_2757,N_1127,N_1598);
nand U2758 (N_2758,N_1795,N_1468);
nand U2759 (N_2759,N_1141,N_1714);
and U2760 (N_2760,N_1250,N_1672);
or U2761 (N_2761,N_1349,N_1805);
and U2762 (N_2762,N_1722,N_1200);
nor U2763 (N_2763,N_1531,N_1150);
nand U2764 (N_2764,N_1042,N_1654);
and U2765 (N_2765,N_1754,N_1800);
and U2766 (N_2766,N_1059,N_1877);
nor U2767 (N_2767,N_1214,N_1926);
or U2768 (N_2768,N_1954,N_1416);
or U2769 (N_2769,N_1488,N_1738);
nand U2770 (N_2770,N_1088,N_1940);
or U2771 (N_2771,N_1880,N_1036);
and U2772 (N_2772,N_1320,N_1509);
and U2773 (N_2773,N_1428,N_1667);
nor U2774 (N_2774,N_1324,N_1308);
nor U2775 (N_2775,N_1867,N_1655);
nor U2776 (N_2776,N_1440,N_1345);
nand U2777 (N_2777,N_1041,N_1140);
and U2778 (N_2778,N_1265,N_1649);
nor U2779 (N_2779,N_1468,N_1940);
nand U2780 (N_2780,N_1904,N_1307);
and U2781 (N_2781,N_1658,N_1577);
or U2782 (N_2782,N_1777,N_1214);
nand U2783 (N_2783,N_1883,N_1550);
nor U2784 (N_2784,N_1520,N_1596);
nand U2785 (N_2785,N_1368,N_1058);
nor U2786 (N_2786,N_1780,N_1027);
and U2787 (N_2787,N_1052,N_1647);
and U2788 (N_2788,N_1750,N_1848);
and U2789 (N_2789,N_1633,N_1058);
or U2790 (N_2790,N_1117,N_1800);
and U2791 (N_2791,N_1320,N_1215);
and U2792 (N_2792,N_1608,N_1402);
nor U2793 (N_2793,N_1929,N_1907);
or U2794 (N_2794,N_1467,N_1176);
or U2795 (N_2795,N_1664,N_1967);
nor U2796 (N_2796,N_1307,N_1456);
nor U2797 (N_2797,N_1422,N_1167);
or U2798 (N_2798,N_1727,N_1890);
and U2799 (N_2799,N_1320,N_1917);
and U2800 (N_2800,N_1978,N_1227);
nand U2801 (N_2801,N_1546,N_1327);
nand U2802 (N_2802,N_1468,N_1536);
nand U2803 (N_2803,N_1216,N_1552);
nand U2804 (N_2804,N_1145,N_1577);
nand U2805 (N_2805,N_1552,N_1000);
nor U2806 (N_2806,N_1572,N_1504);
and U2807 (N_2807,N_1031,N_1537);
nand U2808 (N_2808,N_1959,N_1119);
nand U2809 (N_2809,N_1353,N_1721);
and U2810 (N_2810,N_1581,N_1982);
and U2811 (N_2811,N_1142,N_1956);
nor U2812 (N_2812,N_1856,N_1315);
and U2813 (N_2813,N_1315,N_1920);
xnor U2814 (N_2814,N_1847,N_1439);
or U2815 (N_2815,N_1334,N_1261);
or U2816 (N_2816,N_1715,N_1108);
nor U2817 (N_2817,N_1040,N_1916);
or U2818 (N_2818,N_1415,N_1775);
and U2819 (N_2819,N_1221,N_1227);
nor U2820 (N_2820,N_1213,N_1888);
nand U2821 (N_2821,N_1804,N_1527);
nand U2822 (N_2822,N_1011,N_1427);
and U2823 (N_2823,N_1572,N_1730);
nor U2824 (N_2824,N_1798,N_1638);
nand U2825 (N_2825,N_1650,N_1932);
nand U2826 (N_2826,N_1284,N_1241);
nand U2827 (N_2827,N_1132,N_1154);
and U2828 (N_2828,N_1290,N_1981);
xor U2829 (N_2829,N_1520,N_1192);
and U2830 (N_2830,N_1351,N_1853);
nand U2831 (N_2831,N_1913,N_1849);
nor U2832 (N_2832,N_1598,N_1642);
and U2833 (N_2833,N_1304,N_1260);
nor U2834 (N_2834,N_1557,N_1817);
nand U2835 (N_2835,N_1874,N_1847);
or U2836 (N_2836,N_1260,N_1090);
and U2837 (N_2837,N_1958,N_1515);
and U2838 (N_2838,N_1073,N_1672);
or U2839 (N_2839,N_1259,N_1640);
or U2840 (N_2840,N_1873,N_1941);
or U2841 (N_2841,N_1117,N_1965);
xor U2842 (N_2842,N_1982,N_1840);
nor U2843 (N_2843,N_1248,N_1162);
and U2844 (N_2844,N_1587,N_1965);
nand U2845 (N_2845,N_1908,N_1045);
nor U2846 (N_2846,N_1838,N_1666);
or U2847 (N_2847,N_1112,N_1870);
and U2848 (N_2848,N_1158,N_1138);
nor U2849 (N_2849,N_1391,N_1951);
or U2850 (N_2850,N_1832,N_1575);
or U2851 (N_2851,N_1298,N_1961);
and U2852 (N_2852,N_1081,N_1573);
or U2853 (N_2853,N_1468,N_1957);
nand U2854 (N_2854,N_1251,N_1154);
nand U2855 (N_2855,N_1120,N_1144);
and U2856 (N_2856,N_1326,N_1266);
or U2857 (N_2857,N_1001,N_1553);
and U2858 (N_2858,N_1734,N_1012);
or U2859 (N_2859,N_1210,N_1052);
or U2860 (N_2860,N_1634,N_1754);
nand U2861 (N_2861,N_1139,N_1244);
or U2862 (N_2862,N_1830,N_1883);
nand U2863 (N_2863,N_1845,N_1852);
and U2864 (N_2864,N_1696,N_1313);
and U2865 (N_2865,N_1261,N_1440);
and U2866 (N_2866,N_1747,N_1824);
nand U2867 (N_2867,N_1637,N_1872);
and U2868 (N_2868,N_1898,N_1511);
or U2869 (N_2869,N_1046,N_1847);
or U2870 (N_2870,N_1473,N_1933);
or U2871 (N_2871,N_1019,N_1456);
nand U2872 (N_2872,N_1830,N_1329);
or U2873 (N_2873,N_1917,N_1266);
nor U2874 (N_2874,N_1363,N_1043);
nor U2875 (N_2875,N_1494,N_1040);
nor U2876 (N_2876,N_1682,N_1053);
nand U2877 (N_2877,N_1381,N_1267);
nor U2878 (N_2878,N_1471,N_1289);
nand U2879 (N_2879,N_1357,N_1072);
nor U2880 (N_2880,N_1637,N_1163);
nand U2881 (N_2881,N_1909,N_1186);
nand U2882 (N_2882,N_1009,N_1991);
and U2883 (N_2883,N_1963,N_1372);
and U2884 (N_2884,N_1734,N_1966);
and U2885 (N_2885,N_1814,N_1068);
nor U2886 (N_2886,N_1205,N_1166);
nand U2887 (N_2887,N_1200,N_1077);
nand U2888 (N_2888,N_1917,N_1452);
or U2889 (N_2889,N_1651,N_1568);
nand U2890 (N_2890,N_1723,N_1177);
and U2891 (N_2891,N_1214,N_1933);
or U2892 (N_2892,N_1219,N_1388);
or U2893 (N_2893,N_1248,N_1077);
nand U2894 (N_2894,N_1886,N_1327);
nand U2895 (N_2895,N_1565,N_1629);
nor U2896 (N_2896,N_1858,N_1021);
and U2897 (N_2897,N_1787,N_1946);
nand U2898 (N_2898,N_1043,N_1614);
nand U2899 (N_2899,N_1824,N_1132);
nand U2900 (N_2900,N_1293,N_1798);
and U2901 (N_2901,N_1701,N_1186);
nor U2902 (N_2902,N_1594,N_1158);
nand U2903 (N_2903,N_1458,N_1676);
nor U2904 (N_2904,N_1229,N_1390);
or U2905 (N_2905,N_1353,N_1112);
and U2906 (N_2906,N_1220,N_1081);
nor U2907 (N_2907,N_1123,N_1888);
nor U2908 (N_2908,N_1608,N_1036);
nor U2909 (N_2909,N_1967,N_1490);
nor U2910 (N_2910,N_1982,N_1175);
and U2911 (N_2911,N_1876,N_1164);
and U2912 (N_2912,N_1420,N_1892);
and U2913 (N_2913,N_1633,N_1093);
nand U2914 (N_2914,N_1331,N_1404);
nand U2915 (N_2915,N_1441,N_1028);
nor U2916 (N_2916,N_1550,N_1753);
nand U2917 (N_2917,N_1011,N_1549);
and U2918 (N_2918,N_1907,N_1327);
nor U2919 (N_2919,N_1644,N_1653);
or U2920 (N_2920,N_1826,N_1920);
nor U2921 (N_2921,N_1076,N_1413);
nand U2922 (N_2922,N_1382,N_1075);
or U2923 (N_2923,N_1399,N_1954);
and U2924 (N_2924,N_1005,N_1322);
nor U2925 (N_2925,N_1943,N_1880);
nand U2926 (N_2926,N_1200,N_1126);
or U2927 (N_2927,N_1172,N_1770);
or U2928 (N_2928,N_1447,N_1769);
nor U2929 (N_2929,N_1626,N_1831);
and U2930 (N_2930,N_1693,N_1216);
or U2931 (N_2931,N_1166,N_1948);
or U2932 (N_2932,N_1705,N_1300);
or U2933 (N_2933,N_1126,N_1807);
and U2934 (N_2934,N_1398,N_1436);
and U2935 (N_2935,N_1533,N_1175);
nand U2936 (N_2936,N_1679,N_1934);
nand U2937 (N_2937,N_1773,N_1757);
and U2938 (N_2938,N_1800,N_1931);
and U2939 (N_2939,N_1951,N_1296);
and U2940 (N_2940,N_1993,N_1125);
and U2941 (N_2941,N_1167,N_1444);
nand U2942 (N_2942,N_1020,N_1428);
and U2943 (N_2943,N_1139,N_1624);
or U2944 (N_2944,N_1474,N_1396);
nor U2945 (N_2945,N_1087,N_1440);
nor U2946 (N_2946,N_1799,N_1329);
nand U2947 (N_2947,N_1381,N_1633);
or U2948 (N_2948,N_1634,N_1431);
nand U2949 (N_2949,N_1492,N_1931);
nor U2950 (N_2950,N_1975,N_1367);
or U2951 (N_2951,N_1419,N_1309);
nand U2952 (N_2952,N_1078,N_1899);
and U2953 (N_2953,N_1868,N_1636);
nand U2954 (N_2954,N_1153,N_1884);
or U2955 (N_2955,N_1978,N_1973);
or U2956 (N_2956,N_1525,N_1713);
nand U2957 (N_2957,N_1052,N_1332);
nor U2958 (N_2958,N_1743,N_1839);
and U2959 (N_2959,N_1557,N_1481);
or U2960 (N_2960,N_1910,N_1119);
or U2961 (N_2961,N_1356,N_1043);
nand U2962 (N_2962,N_1034,N_1179);
and U2963 (N_2963,N_1771,N_1301);
and U2964 (N_2964,N_1104,N_1476);
and U2965 (N_2965,N_1686,N_1195);
nand U2966 (N_2966,N_1526,N_1967);
and U2967 (N_2967,N_1229,N_1965);
nor U2968 (N_2968,N_1829,N_1998);
nor U2969 (N_2969,N_1097,N_1283);
and U2970 (N_2970,N_1757,N_1907);
or U2971 (N_2971,N_1091,N_1902);
nand U2972 (N_2972,N_1528,N_1839);
nor U2973 (N_2973,N_1849,N_1241);
nor U2974 (N_2974,N_1235,N_1565);
nand U2975 (N_2975,N_1979,N_1784);
and U2976 (N_2976,N_1263,N_1392);
nor U2977 (N_2977,N_1229,N_1000);
nand U2978 (N_2978,N_1882,N_1337);
or U2979 (N_2979,N_1368,N_1462);
nor U2980 (N_2980,N_1593,N_1024);
or U2981 (N_2981,N_1348,N_1526);
or U2982 (N_2982,N_1138,N_1774);
and U2983 (N_2983,N_1690,N_1329);
nand U2984 (N_2984,N_1707,N_1701);
nand U2985 (N_2985,N_1365,N_1574);
or U2986 (N_2986,N_1749,N_1906);
nor U2987 (N_2987,N_1125,N_1355);
nor U2988 (N_2988,N_1335,N_1085);
nand U2989 (N_2989,N_1809,N_1351);
nand U2990 (N_2990,N_1010,N_1298);
or U2991 (N_2991,N_1417,N_1201);
and U2992 (N_2992,N_1725,N_1529);
and U2993 (N_2993,N_1464,N_1440);
or U2994 (N_2994,N_1574,N_1010);
nand U2995 (N_2995,N_1078,N_1458);
nand U2996 (N_2996,N_1533,N_1361);
nand U2997 (N_2997,N_1865,N_1600);
and U2998 (N_2998,N_1242,N_1761);
or U2999 (N_2999,N_1717,N_1105);
nand U3000 (N_3000,N_2534,N_2819);
and U3001 (N_3001,N_2555,N_2562);
or U3002 (N_3002,N_2724,N_2468);
or U3003 (N_3003,N_2360,N_2774);
nor U3004 (N_3004,N_2745,N_2307);
or U3005 (N_3005,N_2173,N_2149);
nand U3006 (N_3006,N_2813,N_2627);
nand U3007 (N_3007,N_2021,N_2142);
and U3008 (N_3008,N_2662,N_2341);
nor U3009 (N_3009,N_2020,N_2080);
nor U3010 (N_3010,N_2296,N_2891);
or U3011 (N_3011,N_2130,N_2369);
or U3012 (N_3012,N_2012,N_2211);
and U3013 (N_3013,N_2525,N_2685);
or U3014 (N_3014,N_2645,N_2568);
nor U3015 (N_3015,N_2664,N_2210);
nor U3016 (N_3016,N_2680,N_2167);
nor U3017 (N_3017,N_2415,N_2985);
nand U3018 (N_3018,N_2877,N_2359);
and U3019 (N_3019,N_2945,N_2900);
or U3020 (N_3020,N_2803,N_2839);
nor U3021 (N_3021,N_2515,N_2282);
nor U3022 (N_3022,N_2390,N_2110);
nand U3023 (N_3023,N_2125,N_2655);
or U3024 (N_3024,N_2159,N_2491);
nor U3025 (N_3025,N_2538,N_2286);
nor U3026 (N_3026,N_2629,N_2826);
or U3027 (N_3027,N_2416,N_2011);
nand U3028 (N_3028,N_2967,N_2482);
nor U3029 (N_3029,N_2725,N_2492);
nor U3030 (N_3030,N_2437,N_2545);
and U3031 (N_3031,N_2344,N_2205);
nor U3032 (N_3032,N_2141,N_2185);
nor U3033 (N_3033,N_2836,N_2753);
nor U3034 (N_3034,N_2219,N_2171);
nor U3035 (N_3035,N_2245,N_2094);
nor U3036 (N_3036,N_2593,N_2764);
or U3037 (N_3037,N_2871,N_2950);
nand U3038 (N_3038,N_2320,N_2081);
or U3039 (N_3039,N_2844,N_2413);
or U3040 (N_3040,N_2394,N_2448);
and U3041 (N_3041,N_2833,N_2016);
or U3042 (N_3042,N_2500,N_2420);
nand U3043 (N_3043,N_2968,N_2124);
nor U3044 (N_3044,N_2935,N_2951);
and U3045 (N_3045,N_2118,N_2178);
or U3046 (N_3046,N_2030,N_2035);
xnor U3047 (N_3047,N_2668,N_2630);
nor U3048 (N_3048,N_2331,N_2926);
or U3049 (N_3049,N_2481,N_2911);
and U3050 (N_3050,N_2697,N_2823);
nand U3051 (N_3051,N_2698,N_2719);
and U3052 (N_3052,N_2794,N_2550);
and U3053 (N_3053,N_2983,N_2103);
nor U3054 (N_3054,N_2250,N_2116);
nand U3055 (N_3055,N_2706,N_2350);
and U3056 (N_3056,N_2643,N_2625);
and U3057 (N_3057,N_2086,N_2298);
or U3058 (N_3058,N_2034,N_2854);
and U3059 (N_3059,N_2592,N_2838);
and U3060 (N_3060,N_2692,N_2654);
nand U3061 (N_3061,N_2339,N_2033);
nor U3062 (N_3062,N_2365,N_2485);
and U3063 (N_3063,N_2965,N_2942);
nand U3064 (N_3064,N_2280,N_2934);
nand U3065 (N_3065,N_2564,N_2106);
nor U3066 (N_3066,N_2189,N_2901);
or U3067 (N_3067,N_2535,N_2640);
and U3068 (N_3068,N_2793,N_2291);
or U3069 (N_3069,N_2781,N_2997);
or U3070 (N_3070,N_2139,N_2423);
nor U3071 (N_3071,N_2343,N_2284);
and U3072 (N_3072,N_2755,N_2237);
nor U3073 (N_3073,N_2288,N_2557);
nand U3074 (N_3074,N_2271,N_2203);
xnor U3075 (N_3075,N_2148,N_2522);
and U3076 (N_3076,N_2441,N_2954);
and U3077 (N_3077,N_2073,N_2665);
nand U3078 (N_3078,N_2795,N_2824);
nand U3079 (N_3079,N_2843,N_2999);
nor U3080 (N_3080,N_2032,N_2054);
and U3081 (N_3081,N_2299,N_2315);
nand U3082 (N_3082,N_2959,N_2537);
and U3083 (N_3083,N_2278,N_2509);
and U3084 (N_3084,N_2262,N_2244);
or U3085 (N_3085,N_2647,N_2742);
or U3086 (N_3086,N_2811,N_2329);
or U3087 (N_3087,N_2913,N_2184);
nor U3088 (N_3088,N_2372,N_2695);
and U3089 (N_3089,N_2650,N_2883);
or U3090 (N_3090,N_2792,N_2608);
or U3091 (N_3091,N_2111,N_2536);
nand U3092 (N_3092,N_2170,N_2504);
nor U3093 (N_3093,N_2932,N_2025);
and U3094 (N_3094,N_2421,N_2850);
or U3095 (N_3095,N_2101,N_2261);
nand U3096 (N_3096,N_2731,N_2347);
nand U3097 (N_3097,N_2231,N_2379);
and U3098 (N_3098,N_2346,N_2206);
and U3099 (N_3099,N_2841,N_2022);
and U3100 (N_3100,N_2642,N_2517);
and U3101 (N_3101,N_2580,N_2682);
and U3102 (N_3102,N_2160,N_2464);
and U3103 (N_3103,N_2085,N_2332);
and U3104 (N_3104,N_2163,N_2031);
nor U3105 (N_3105,N_2104,N_2723);
or U3106 (N_3106,N_2461,N_2079);
xor U3107 (N_3107,N_2358,N_2115);
nand U3108 (N_3108,N_2513,N_2514);
and U3109 (N_3109,N_2075,N_2552);
or U3110 (N_3110,N_2456,N_2646);
or U3111 (N_3111,N_2218,N_2671);
and U3112 (N_3112,N_2093,N_2191);
or U3113 (N_3113,N_2677,N_2038);
nand U3114 (N_3114,N_2200,N_2388);
or U3115 (N_3115,N_2739,N_2524);
nor U3116 (N_3116,N_2693,N_2947);
and U3117 (N_3117,N_2409,N_2077);
nor U3118 (N_3118,N_2626,N_2921);
nor U3119 (N_3119,N_2366,N_2966);
nand U3120 (N_3120,N_2145,N_2330);
and U3121 (N_3121,N_2806,N_2447);
nand U3122 (N_3122,N_2567,N_2019);
nor U3123 (N_3123,N_2336,N_2804);
nor U3124 (N_3124,N_2469,N_2912);
and U3125 (N_3125,N_2771,N_2785);
nand U3126 (N_3126,N_2544,N_2858);
nor U3127 (N_3127,N_2380,N_2573);
nand U3128 (N_3128,N_2026,N_2196);
nor U3129 (N_3129,N_2128,N_2931);
nand U3130 (N_3130,N_2099,N_2156);
nor U3131 (N_3131,N_2247,N_2754);
and U3132 (N_3132,N_2224,N_2418);
nand U3133 (N_3133,N_2475,N_2972);
nand U3134 (N_3134,N_2052,N_2316);
nor U3135 (N_3135,N_2182,N_2711);
or U3136 (N_3136,N_2228,N_2837);
and U3137 (N_3137,N_2601,N_2887);
nand U3138 (N_3138,N_2113,N_2266);
or U3139 (N_3139,N_2782,N_2240);
and U3140 (N_3140,N_2164,N_2051);
and U3141 (N_3141,N_2994,N_2119);
and U3142 (N_3142,N_2979,N_2598);
nor U3143 (N_3143,N_2187,N_2402);
and U3144 (N_3144,N_2632,N_2684);
nand U3145 (N_3145,N_2374,N_2832);
or U3146 (N_3146,N_2855,N_2808);
nor U3147 (N_3147,N_2090,N_2209);
and U3148 (N_3148,N_2340,N_2373);
or U3149 (N_3149,N_2758,N_2432);
and U3150 (N_3150,N_2749,N_2066);
nand U3151 (N_3151,N_2805,N_2830);
and U3152 (N_3152,N_2208,N_2820);
and U3153 (N_3153,N_2740,N_2107);
nand U3154 (N_3154,N_2064,N_2589);
nand U3155 (N_3155,N_2988,N_2575);
nand U3156 (N_3156,N_2455,N_2962);
nand U3157 (N_3157,N_2326,N_2914);
nor U3158 (N_3158,N_2700,N_2548);
or U3159 (N_3159,N_2272,N_2578);
or U3160 (N_3160,N_2560,N_2975);
or U3161 (N_3161,N_2197,N_2623);
nor U3162 (N_3162,N_2490,N_2579);
nand U3163 (N_3163,N_2338,N_2223);
and U3164 (N_3164,N_2070,N_2230);
or U3165 (N_3165,N_2186,N_2896);
or U3166 (N_3166,N_2165,N_2328);
nor U3167 (N_3167,N_2474,N_2401);
and U3168 (N_3168,N_2920,N_2131);
or U3169 (N_3169,N_2400,N_2306);
nand U3170 (N_3170,N_2227,N_2006);
or U3171 (N_3171,N_2003,N_2289);
and U3172 (N_3172,N_2909,N_2737);
or U3173 (N_3173,N_2880,N_2465);
nor U3174 (N_3174,N_2644,N_2129);
and U3175 (N_3175,N_2588,N_2614);
nor U3176 (N_3176,N_2114,N_2239);
and U3177 (N_3177,N_2748,N_2023);
and U3178 (N_3178,N_2007,N_2084);
nor U3179 (N_3179,N_2789,N_2870);
nand U3180 (N_3180,N_2087,N_2304);
nand U3181 (N_3181,N_2501,N_2483);
or U3182 (N_3182,N_2984,N_2342);
or U3183 (N_3183,N_2842,N_2799);
nand U3184 (N_3184,N_2605,N_2956);
nand U3185 (N_3185,N_2987,N_2056);
or U3186 (N_3186,N_2417,N_2181);
xor U3187 (N_3187,N_2046,N_2220);
and U3188 (N_3188,N_2277,N_2572);
nor U3189 (N_3189,N_2109,N_2786);
nor U3190 (N_3190,N_2251,N_2459);
and U3191 (N_3191,N_2260,N_2484);
or U3192 (N_3192,N_2948,N_2439);
and U3193 (N_3193,N_2990,N_2657);
nor U3194 (N_3194,N_2936,N_2587);
and U3195 (N_3195,N_2886,N_2777);
or U3196 (N_3196,N_2856,N_2773);
or U3197 (N_3197,N_2193,N_2807);
nand U3198 (N_3198,N_2551,N_2775);
nor U3199 (N_3199,N_2744,N_2467);
and U3200 (N_3200,N_2757,N_2728);
and U3201 (N_3201,N_2002,N_2566);
or U3202 (N_3202,N_2606,N_2403);
and U3203 (N_3203,N_2202,N_2683);
nor U3204 (N_3204,N_2769,N_2917);
and U3205 (N_3205,N_2057,N_2472);
nor U3206 (N_3206,N_2096,N_2958);
nand U3207 (N_3207,N_2776,N_2290);
and U3208 (N_3208,N_2690,N_2355);
nor U3209 (N_3209,N_2798,N_2177);
nand U3210 (N_3210,N_2878,N_2424);
and U3211 (N_3211,N_2628,N_2893);
and U3212 (N_3212,N_2584,N_2151);
nand U3213 (N_3213,N_2345,N_2553);
nand U3214 (N_3214,N_2443,N_2168);
or U3215 (N_3215,N_2506,N_2300);
and U3216 (N_3216,N_2408,N_2297);
and U3217 (N_3217,N_2001,N_2670);
nand U3218 (N_3218,N_2709,N_2631);
or U3219 (N_3219,N_2162,N_2619);
nor U3220 (N_3220,N_2076,N_2493);
nand U3221 (N_3221,N_2736,N_2371);
nor U3222 (N_3222,N_2215,N_2814);
and U3223 (N_3223,N_2554,N_2929);
or U3224 (N_3224,N_2586,N_2204);
and U3225 (N_3225,N_2922,N_2498);
nand U3226 (N_3226,N_2082,N_2473);
nor U3227 (N_3227,N_2865,N_2686);
or U3228 (N_3228,N_2879,N_2663);
and U3229 (N_3229,N_2221,N_2312);
or U3230 (N_3230,N_2067,N_2188);
nor U3231 (N_3231,N_2232,N_2072);
or U3232 (N_3232,N_2146,N_2367);
and U3233 (N_3233,N_2651,N_2790);
nand U3234 (N_3234,N_2859,N_2732);
and U3235 (N_3235,N_2676,N_2691);
nor U3236 (N_3236,N_2787,N_2302);
nand U3237 (N_3237,N_2477,N_2977);
or U3238 (N_3238,N_2255,N_2652);
or U3239 (N_3239,N_2039,N_2058);
or U3240 (N_3240,N_2800,N_2895);
and U3241 (N_3241,N_2581,N_2729);
and U3242 (N_3242,N_2989,N_2194);
and U3243 (N_3243,N_2180,N_2069);
and U3244 (N_3244,N_2916,N_2516);
nor U3245 (N_3245,N_2386,N_2829);
nor U3246 (N_3246,N_2674,N_2822);
or U3247 (N_3247,N_2241,N_2810);
or U3248 (N_3248,N_2253,N_2257);
nor U3249 (N_3249,N_2065,N_2137);
and U3250 (N_3250,N_2314,N_2705);
or U3251 (N_3251,N_2694,N_2480);
nand U3252 (N_3252,N_2411,N_2494);
nand U3253 (N_3253,N_2610,N_2885);
or U3254 (N_3254,N_2273,N_2641);
and U3255 (N_3255,N_2061,N_2635);
and U3256 (N_3256,N_2426,N_2852);
nor U3257 (N_3257,N_2570,N_2466);
nand U3258 (N_3258,N_2961,N_2334);
or U3259 (N_3259,N_2565,N_2395);
nor U3260 (N_3260,N_2802,N_2243);
nand U3261 (N_3261,N_2730,N_2201);
or U3262 (N_3262,N_2818,N_2720);
and U3263 (N_3263,N_2287,N_2122);
or U3264 (N_3264,N_2910,N_2496);
and U3265 (N_3265,N_2558,N_2688);
or U3266 (N_3266,N_2571,N_2337);
nand U3267 (N_3267,N_2140,N_2495);
or U3268 (N_3268,N_2527,N_2574);
and U3269 (N_3269,N_2134,N_2313);
or U3270 (N_3270,N_2095,N_2460);
or U3271 (N_3271,N_2866,N_2017);
nor U3272 (N_3272,N_2704,N_2591);
and U3273 (N_3273,N_2973,N_2752);
nand U3274 (N_3274,N_2258,N_2845);
nor U3275 (N_3275,N_2351,N_2874);
and U3276 (N_3276,N_2393,N_2040);
or U3277 (N_3277,N_2892,N_2797);
nor U3278 (N_3278,N_2721,N_2746);
or U3279 (N_3279,N_2091,N_2609);
nand U3280 (N_3280,N_2190,N_2349);
nand U3281 (N_3281,N_2324,N_2414);
or U3282 (N_3282,N_2108,N_2569);
nor U3283 (N_3283,N_2648,N_2812);
or U3284 (N_3284,N_2009,N_2249);
or U3285 (N_3285,N_2161,N_2270);
or U3286 (N_3286,N_2512,N_2970);
nor U3287 (N_3287,N_2169,N_2399);
and U3288 (N_3288,N_2303,N_2993);
and U3289 (N_3289,N_2179,N_2599);
nor U3290 (N_3290,N_2766,N_2707);
nand U3291 (N_3291,N_2276,N_2348);
or U3292 (N_3292,N_2463,N_2097);
nand U3293 (N_3293,N_2768,N_2659);
nor U3294 (N_3294,N_2907,N_2528);
and U3295 (N_3295,N_2649,N_2759);
and U3296 (N_3296,N_2633,N_2708);
nand U3297 (N_3297,N_2846,N_2442);
and U3298 (N_3298,N_2582,N_2577);
nor U3299 (N_3299,N_2612,N_2045);
nor U3300 (N_3300,N_2433,N_2430);
and U3301 (N_3301,N_2868,N_2899);
and U3302 (N_3302,N_2638,N_2378);
or U3303 (N_3303,N_2767,N_2600);
or U3304 (N_3304,N_2236,N_2996);
nand U3305 (N_3305,N_2317,N_2727);
and U3306 (N_3306,N_2960,N_2595);
or U3307 (N_3307,N_2364,N_2422);
nor U3308 (N_3308,N_2863,N_2703);
or U3309 (N_3309,N_2445,N_2295);
and U3310 (N_3310,N_2834,N_2634);
nor U3311 (N_3311,N_2860,N_2702);
nand U3312 (N_3312,N_2319,N_2849);
or U3313 (N_3313,N_2943,N_2898);
or U3314 (N_3314,N_2144,N_2888);
nand U3315 (N_3315,N_2998,N_2015);
and U3316 (N_3316,N_2894,N_2102);
nor U3317 (N_3317,N_2050,N_2222);
or U3318 (N_3318,N_2981,N_2964);
nand U3319 (N_3319,N_2831,N_2992);
and U3320 (N_3320,N_2532,N_2675);
nand U3321 (N_3321,N_2294,N_2059);
or U3322 (N_3322,N_2488,N_2269);
nor U3323 (N_3323,N_2602,N_2861);
nand U3324 (N_3324,N_2726,N_2449);
nand U3325 (N_3325,N_2252,N_2656);
nor U3326 (N_3326,N_2323,N_2621);
and U3327 (N_3327,N_2658,N_2809);
nor U3328 (N_3328,N_2428,N_2876);
or U3329 (N_3329,N_2696,N_2733);
nand U3330 (N_3330,N_2383,N_2487);
nand U3331 (N_3331,N_2068,N_2207);
or U3332 (N_3332,N_2949,N_2004);
and U3333 (N_3333,N_2505,N_2563);
or U3334 (N_3334,N_2559,N_2853);
nor U3335 (N_3335,N_2507,N_2583);
nand U3336 (N_3336,N_2225,N_2738);
nand U3337 (N_3337,N_2391,N_2311);
nand U3338 (N_3338,N_2840,N_2539);
and U3339 (N_3339,N_2783,N_2419);
and U3340 (N_3340,N_2940,N_2884);
nand U3341 (N_3341,N_2957,N_2440);
and U3342 (N_3342,N_2963,N_2429);
nor U3343 (N_3343,N_2828,N_2980);
and U3344 (N_3344,N_2214,N_2924);
nand U3345 (N_3345,N_2120,N_2955);
and U3346 (N_3346,N_2044,N_2174);
or U3347 (N_3347,N_2071,N_2361);
nor U3348 (N_3348,N_2235,N_2672);
nor U3349 (N_3349,N_2519,N_2157);
or U3350 (N_3350,N_2308,N_2412);
and U3351 (N_3351,N_2135,N_2370);
or U3352 (N_3352,N_2105,N_2607);
xnor U3353 (N_3353,N_2281,N_2238);
nor U3354 (N_3354,N_2166,N_2511);
or U3355 (N_3355,N_2398,N_2027);
or U3356 (N_3356,N_2112,N_2136);
nor U3357 (N_3357,N_2890,N_2760);
nor U3358 (N_3358,N_2037,N_2353);
nand U3359 (N_3359,N_2751,N_2041);
nor U3360 (N_3360,N_2048,N_2479);
nand U3361 (N_3361,N_2679,N_2476);
nor U3362 (N_3362,N_2049,N_2747);
or U3363 (N_3363,N_2974,N_2615);
nor U3364 (N_3364,N_2576,N_2407);
nand U3365 (N_3365,N_2590,N_2872);
nor U3366 (N_3366,N_2923,N_2715);
nor U3367 (N_3367,N_2042,N_2368);
or U3368 (N_3368,N_2750,N_2248);
xnor U3369 (N_3369,N_2499,N_2918);
or U3370 (N_3370,N_2763,N_2780);
nand U3371 (N_3371,N_2325,N_2620);
and U3372 (N_3372,N_2889,N_2435);
or U3373 (N_3373,N_2801,N_2976);
nor U3374 (N_3374,N_2716,N_2765);
nand U3375 (N_3375,N_2431,N_2903);
nor U3376 (N_3376,N_2543,N_2521);
or U3377 (N_3377,N_2024,N_2713);
nor U3378 (N_3378,N_2063,N_2510);
nor U3379 (N_3379,N_2436,N_2335);
or U3380 (N_3380,N_2667,N_2176);
nor U3381 (N_3381,N_2470,N_2978);
and U3382 (N_3382,N_2242,N_2089);
and U3383 (N_3383,N_2375,N_2927);
or U3384 (N_3384,N_2133,N_2217);
and U3385 (N_3385,N_2678,N_2305);
and U3386 (N_3386,N_2126,N_2387);
nand U3387 (N_3387,N_2734,N_2661);
and U3388 (N_3388,N_2952,N_2546);
or U3389 (N_3389,N_2489,N_2622);
and U3390 (N_3390,N_2259,N_2410);
nor U3391 (N_3391,N_2301,N_2318);
and U3392 (N_3392,N_2078,N_2636);
nor U3393 (N_3393,N_2233,N_2062);
xor U3394 (N_3394,N_2827,N_2396);
nand U3395 (N_3395,N_2778,N_2906);
nor U3396 (N_3396,N_2847,N_2928);
nand U3397 (N_3397,N_2018,N_2523);
and U3398 (N_3398,N_2497,N_2817);
or U3399 (N_3399,N_2542,N_2404);
and U3400 (N_3400,N_2138,N_2772);
nor U3401 (N_3401,N_2267,N_2309);
nor U3402 (N_3402,N_2478,N_2055);
or U3403 (N_3403,N_2444,N_2561);
nand U3404 (N_3404,N_2603,N_2618);
nor U3405 (N_3405,N_2547,N_2937);
nor U3406 (N_3406,N_2333,N_2761);
nand U3407 (N_3407,N_2875,N_2352);
or U3408 (N_3408,N_2784,N_2717);
or U3409 (N_3409,N_2123,N_2226);
or U3410 (N_3410,N_2639,N_2100);
nand U3411 (N_3411,N_2712,N_2882);
nor U3412 (N_3412,N_2533,N_2995);
and U3413 (N_3413,N_2285,N_2718);
nor U3414 (N_3414,N_2264,N_2283);
nand U3415 (N_3415,N_2153,N_2256);
nand U3416 (N_3416,N_2152,N_2092);
nand U3417 (N_3417,N_2933,N_2857);
and U3418 (N_3418,N_2556,N_2848);
or U3419 (N_3419,N_2377,N_2597);
or U3420 (N_3420,N_2938,N_2274);
and U3421 (N_3421,N_2919,N_2385);
xnor U3422 (N_3422,N_2982,N_2384);
or U3423 (N_3423,N_2915,N_2624);
nand U3424 (N_3424,N_2611,N_2014);
nand U3425 (N_3425,N_2321,N_2392);
and U3426 (N_3426,N_2944,N_2788);
nor U3427 (N_3427,N_2991,N_2825);
or U3428 (N_3428,N_2971,N_2779);
nand U3429 (N_3429,N_2389,N_2450);
nor U3430 (N_3430,N_2000,N_2310);
nor U3431 (N_3431,N_2681,N_2791);
nand U3432 (N_3432,N_2446,N_2756);
or U3433 (N_3433,N_2653,N_2939);
or U3434 (N_3434,N_2503,N_2074);
nor U3435 (N_3435,N_2457,N_2183);
or U3436 (N_3436,N_2229,N_2613);
nand U3437 (N_3437,N_2043,N_2835);
or U3438 (N_3438,N_2585,N_2908);
nand U3439 (N_3439,N_2673,N_2327);
or U3440 (N_3440,N_2212,N_2520);
and U3441 (N_3441,N_2425,N_2941);
or U3442 (N_3442,N_2434,N_2147);
nand U3443 (N_3443,N_2047,N_2234);
and U3444 (N_3444,N_2013,N_2452);
or U3445 (N_3445,N_2216,N_2770);
nor U3446 (N_3446,N_2925,N_2088);
and U3447 (N_3447,N_2540,N_2199);
or U3448 (N_3448,N_2098,N_2005);
nor U3449 (N_3449,N_2735,N_2053);
and U3450 (N_3450,N_2406,N_2529);
and U3451 (N_3451,N_2710,N_2117);
or U3452 (N_3452,N_2127,N_2815);
and U3453 (N_3453,N_2905,N_2198);
or U3454 (N_3454,N_2486,N_2508);
nand U3455 (N_3455,N_2268,N_2530);
or U3456 (N_3456,N_2549,N_2669);
and U3457 (N_3457,N_2873,N_2279);
or U3458 (N_3458,N_2864,N_2438);
or U3459 (N_3459,N_2897,N_2453);
and U3460 (N_3460,N_2172,N_2275);
and U3461 (N_3461,N_2953,N_2604);
and U3462 (N_3462,N_2132,N_2246);
nor U3463 (N_3463,N_2292,N_2451);
nor U3464 (N_3464,N_2660,N_2362);
and U3465 (N_3465,N_2743,N_2376);
nor U3466 (N_3466,N_2796,N_2969);
nor U3467 (N_3467,N_2028,N_2904);
nor U3468 (N_3468,N_2869,N_2356);
nor U3469 (N_3469,N_2060,N_2594);
nor U3470 (N_3470,N_2265,N_2010);
nand U3471 (N_3471,N_2616,N_2029);
nor U3472 (N_3472,N_2293,N_2902);
and U3473 (N_3473,N_2821,N_2526);
and U3474 (N_3474,N_2382,N_2036);
nand U3475 (N_3475,N_2531,N_2722);
or U3476 (N_3476,N_2462,N_2405);
xor U3477 (N_3477,N_2322,N_2637);
nor U3478 (N_3478,N_2666,N_2762);
or U3479 (N_3479,N_2143,N_2213);
or U3480 (N_3480,N_2150,N_2502);
and U3481 (N_3481,N_2175,N_2867);
and U3482 (N_3482,N_2714,N_2699);
nand U3483 (N_3483,N_2518,N_2816);
and U3484 (N_3484,N_2881,N_2541);
nand U3485 (N_3485,N_2458,N_2701);
nand U3486 (N_3486,N_2154,N_2946);
or U3487 (N_3487,N_2357,N_2263);
or U3488 (N_3488,N_2596,N_2454);
nand U3489 (N_3489,N_2986,N_2121);
nand U3490 (N_3490,N_2617,N_2381);
nor U3491 (N_3491,N_2930,N_2192);
or U3492 (N_3492,N_2254,N_2195);
nand U3493 (N_3493,N_2158,N_2689);
and U3494 (N_3494,N_2397,N_2155);
or U3495 (N_3495,N_2851,N_2427);
nor U3496 (N_3496,N_2862,N_2008);
xnor U3497 (N_3497,N_2363,N_2083);
nand U3498 (N_3498,N_2354,N_2741);
or U3499 (N_3499,N_2471,N_2687);
nand U3500 (N_3500,N_2882,N_2804);
and U3501 (N_3501,N_2145,N_2957);
nand U3502 (N_3502,N_2421,N_2697);
and U3503 (N_3503,N_2049,N_2617);
nand U3504 (N_3504,N_2024,N_2829);
and U3505 (N_3505,N_2429,N_2090);
nand U3506 (N_3506,N_2842,N_2595);
and U3507 (N_3507,N_2643,N_2738);
and U3508 (N_3508,N_2488,N_2619);
nand U3509 (N_3509,N_2568,N_2334);
or U3510 (N_3510,N_2929,N_2462);
nand U3511 (N_3511,N_2158,N_2548);
nand U3512 (N_3512,N_2608,N_2184);
or U3513 (N_3513,N_2801,N_2756);
or U3514 (N_3514,N_2568,N_2409);
nand U3515 (N_3515,N_2788,N_2961);
nor U3516 (N_3516,N_2179,N_2085);
and U3517 (N_3517,N_2452,N_2258);
nor U3518 (N_3518,N_2256,N_2247);
nand U3519 (N_3519,N_2667,N_2925);
or U3520 (N_3520,N_2734,N_2589);
nor U3521 (N_3521,N_2859,N_2912);
and U3522 (N_3522,N_2494,N_2207);
nor U3523 (N_3523,N_2423,N_2233);
nor U3524 (N_3524,N_2892,N_2819);
nor U3525 (N_3525,N_2820,N_2467);
or U3526 (N_3526,N_2754,N_2660);
and U3527 (N_3527,N_2933,N_2271);
or U3528 (N_3528,N_2821,N_2783);
or U3529 (N_3529,N_2229,N_2791);
or U3530 (N_3530,N_2662,N_2587);
xor U3531 (N_3531,N_2678,N_2416);
and U3532 (N_3532,N_2140,N_2795);
nor U3533 (N_3533,N_2471,N_2607);
nor U3534 (N_3534,N_2604,N_2687);
and U3535 (N_3535,N_2432,N_2752);
nand U3536 (N_3536,N_2043,N_2993);
nand U3537 (N_3537,N_2939,N_2429);
and U3538 (N_3538,N_2275,N_2647);
nand U3539 (N_3539,N_2332,N_2000);
or U3540 (N_3540,N_2665,N_2196);
or U3541 (N_3541,N_2297,N_2276);
and U3542 (N_3542,N_2106,N_2753);
nand U3543 (N_3543,N_2785,N_2374);
or U3544 (N_3544,N_2818,N_2162);
or U3545 (N_3545,N_2038,N_2843);
nor U3546 (N_3546,N_2845,N_2679);
or U3547 (N_3547,N_2443,N_2806);
and U3548 (N_3548,N_2835,N_2271);
and U3549 (N_3549,N_2451,N_2881);
nand U3550 (N_3550,N_2245,N_2329);
nand U3551 (N_3551,N_2867,N_2452);
xnor U3552 (N_3552,N_2883,N_2064);
nor U3553 (N_3553,N_2129,N_2178);
and U3554 (N_3554,N_2084,N_2925);
and U3555 (N_3555,N_2393,N_2394);
and U3556 (N_3556,N_2189,N_2771);
nand U3557 (N_3557,N_2593,N_2074);
or U3558 (N_3558,N_2832,N_2582);
or U3559 (N_3559,N_2618,N_2947);
nand U3560 (N_3560,N_2199,N_2740);
or U3561 (N_3561,N_2066,N_2840);
nand U3562 (N_3562,N_2679,N_2343);
nand U3563 (N_3563,N_2744,N_2861);
or U3564 (N_3564,N_2367,N_2279);
nor U3565 (N_3565,N_2197,N_2316);
and U3566 (N_3566,N_2006,N_2971);
nand U3567 (N_3567,N_2274,N_2927);
or U3568 (N_3568,N_2097,N_2616);
nor U3569 (N_3569,N_2334,N_2974);
nand U3570 (N_3570,N_2755,N_2777);
or U3571 (N_3571,N_2879,N_2911);
nand U3572 (N_3572,N_2026,N_2615);
and U3573 (N_3573,N_2487,N_2664);
nor U3574 (N_3574,N_2569,N_2331);
nor U3575 (N_3575,N_2167,N_2417);
nor U3576 (N_3576,N_2468,N_2580);
or U3577 (N_3577,N_2888,N_2869);
nand U3578 (N_3578,N_2096,N_2098);
or U3579 (N_3579,N_2722,N_2930);
nor U3580 (N_3580,N_2170,N_2972);
nand U3581 (N_3581,N_2852,N_2178);
nand U3582 (N_3582,N_2992,N_2040);
nor U3583 (N_3583,N_2007,N_2381);
and U3584 (N_3584,N_2349,N_2473);
and U3585 (N_3585,N_2268,N_2853);
nor U3586 (N_3586,N_2744,N_2919);
nor U3587 (N_3587,N_2827,N_2169);
or U3588 (N_3588,N_2397,N_2473);
nor U3589 (N_3589,N_2255,N_2144);
nand U3590 (N_3590,N_2075,N_2271);
and U3591 (N_3591,N_2466,N_2854);
nand U3592 (N_3592,N_2700,N_2788);
and U3593 (N_3593,N_2770,N_2585);
or U3594 (N_3594,N_2402,N_2237);
or U3595 (N_3595,N_2275,N_2361);
nand U3596 (N_3596,N_2434,N_2566);
nand U3597 (N_3597,N_2251,N_2815);
nor U3598 (N_3598,N_2970,N_2266);
or U3599 (N_3599,N_2290,N_2527);
or U3600 (N_3600,N_2954,N_2061);
nand U3601 (N_3601,N_2245,N_2420);
or U3602 (N_3602,N_2865,N_2695);
and U3603 (N_3603,N_2518,N_2697);
and U3604 (N_3604,N_2405,N_2213);
and U3605 (N_3605,N_2698,N_2692);
and U3606 (N_3606,N_2979,N_2495);
nand U3607 (N_3607,N_2839,N_2559);
nor U3608 (N_3608,N_2815,N_2736);
nor U3609 (N_3609,N_2196,N_2896);
or U3610 (N_3610,N_2450,N_2460);
or U3611 (N_3611,N_2217,N_2101);
nor U3612 (N_3612,N_2538,N_2292);
or U3613 (N_3613,N_2979,N_2504);
or U3614 (N_3614,N_2701,N_2443);
or U3615 (N_3615,N_2557,N_2416);
and U3616 (N_3616,N_2808,N_2829);
nand U3617 (N_3617,N_2322,N_2588);
or U3618 (N_3618,N_2537,N_2895);
and U3619 (N_3619,N_2295,N_2022);
or U3620 (N_3620,N_2213,N_2386);
nand U3621 (N_3621,N_2779,N_2303);
nor U3622 (N_3622,N_2224,N_2752);
nor U3623 (N_3623,N_2019,N_2081);
and U3624 (N_3624,N_2736,N_2838);
nand U3625 (N_3625,N_2077,N_2494);
or U3626 (N_3626,N_2956,N_2353);
or U3627 (N_3627,N_2396,N_2045);
and U3628 (N_3628,N_2467,N_2145);
or U3629 (N_3629,N_2244,N_2305);
or U3630 (N_3630,N_2437,N_2246);
and U3631 (N_3631,N_2681,N_2114);
nand U3632 (N_3632,N_2620,N_2274);
and U3633 (N_3633,N_2140,N_2272);
or U3634 (N_3634,N_2187,N_2076);
nor U3635 (N_3635,N_2963,N_2368);
and U3636 (N_3636,N_2841,N_2634);
and U3637 (N_3637,N_2882,N_2247);
and U3638 (N_3638,N_2525,N_2067);
nand U3639 (N_3639,N_2949,N_2198);
nand U3640 (N_3640,N_2104,N_2064);
nand U3641 (N_3641,N_2454,N_2284);
nand U3642 (N_3642,N_2576,N_2378);
nand U3643 (N_3643,N_2215,N_2753);
nand U3644 (N_3644,N_2423,N_2623);
nor U3645 (N_3645,N_2302,N_2729);
nand U3646 (N_3646,N_2965,N_2261);
nand U3647 (N_3647,N_2230,N_2977);
nor U3648 (N_3648,N_2913,N_2460);
and U3649 (N_3649,N_2154,N_2811);
nor U3650 (N_3650,N_2236,N_2691);
and U3651 (N_3651,N_2381,N_2261);
and U3652 (N_3652,N_2592,N_2692);
or U3653 (N_3653,N_2272,N_2422);
or U3654 (N_3654,N_2778,N_2128);
or U3655 (N_3655,N_2234,N_2106);
nand U3656 (N_3656,N_2204,N_2003);
nand U3657 (N_3657,N_2521,N_2286);
or U3658 (N_3658,N_2438,N_2480);
nand U3659 (N_3659,N_2298,N_2650);
nand U3660 (N_3660,N_2049,N_2858);
and U3661 (N_3661,N_2516,N_2417);
nor U3662 (N_3662,N_2357,N_2315);
and U3663 (N_3663,N_2608,N_2472);
and U3664 (N_3664,N_2976,N_2974);
nor U3665 (N_3665,N_2281,N_2672);
or U3666 (N_3666,N_2490,N_2572);
or U3667 (N_3667,N_2806,N_2298);
nand U3668 (N_3668,N_2559,N_2656);
nand U3669 (N_3669,N_2882,N_2332);
nand U3670 (N_3670,N_2948,N_2154);
and U3671 (N_3671,N_2806,N_2699);
or U3672 (N_3672,N_2790,N_2168);
nor U3673 (N_3673,N_2343,N_2805);
nand U3674 (N_3674,N_2261,N_2387);
or U3675 (N_3675,N_2016,N_2510);
nand U3676 (N_3676,N_2063,N_2918);
nor U3677 (N_3677,N_2475,N_2995);
nor U3678 (N_3678,N_2014,N_2881);
nand U3679 (N_3679,N_2526,N_2661);
or U3680 (N_3680,N_2199,N_2330);
nor U3681 (N_3681,N_2963,N_2097);
nor U3682 (N_3682,N_2285,N_2185);
nand U3683 (N_3683,N_2717,N_2044);
or U3684 (N_3684,N_2168,N_2735);
nor U3685 (N_3685,N_2654,N_2888);
and U3686 (N_3686,N_2171,N_2820);
or U3687 (N_3687,N_2519,N_2266);
and U3688 (N_3688,N_2665,N_2860);
and U3689 (N_3689,N_2002,N_2141);
nand U3690 (N_3690,N_2673,N_2871);
and U3691 (N_3691,N_2320,N_2475);
nor U3692 (N_3692,N_2498,N_2269);
and U3693 (N_3693,N_2253,N_2530);
or U3694 (N_3694,N_2631,N_2762);
nor U3695 (N_3695,N_2796,N_2702);
or U3696 (N_3696,N_2621,N_2541);
or U3697 (N_3697,N_2097,N_2580);
nand U3698 (N_3698,N_2235,N_2698);
or U3699 (N_3699,N_2542,N_2286);
and U3700 (N_3700,N_2281,N_2968);
nand U3701 (N_3701,N_2328,N_2022);
nor U3702 (N_3702,N_2187,N_2004);
nand U3703 (N_3703,N_2905,N_2243);
and U3704 (N_3704,N_2291,N_2423);
nor U3705 (N_3705,N_2103,N_2146);
and U3706 (N_3706,N_2485,N_2073);
nand U3707 (N_3707,N_2348,N_2384);
or U3708 (N_3708,N_2131,N_2452);
nand U3709 (N_3709,N_2825,N_2843);
and U3710 (N_3710,N_2150,N_2636);
nand U3711 (N_3711,N_2738,N_2866);
nand U3712 (N_3712,N_2978,N_2930);
nor U3713 (N_3713,N_2712,N_2332);
and U3714 (N_3714,N_2928,N_2403);
nand U3715 (N_3715,N_2711,N_2220);
nand U3716 (N_3716,N_2654,N_2955);
nor U3717 (N_3717,N_2432,N_2039);
nand U3718 (N_3718,N_2095,N_2579);
and U3719 (N_3719,N_2455,N_2359);
nand U3720 (N_3720,N_2672,N_2427);
and U3721 (N_3721,N_2882,N_2991);
nand U3722 (N_3722,N_2536,N_2825);
nor U3723 (N_3723,N_2350,N_2194);
nor U3724 (N_3724,N_2245,N_2443);
nor U3725 (N_3725,N_2793,N_2146);
and U3726 (N_3726,N_2230,N_2111);
nor U3727 (N_3727,N_2459,N_2639);
or U3728 (N_3728,N_2020,N_2693);
nor U3729 (N_3729,N_2821,N_2818);
and U3730 (N_3730,N_2806,N_2746);
nor U3731 (N_3731,N_2196,N_2207);
and U3732 (N_3732,N_2759,N_2501);
nand U3733 (N_3733,N_2376,N_2032);
and U3734 (N_3734,N_2862,N_2362);
nand U3735 (N_3735,N_2547,N_2320);
nor U3736 (N_3736,N_2706,N_2106);
nor U3737 (N_3737,N_2483,N_2835);
nor U3738 (N_3738,N_2699,N_2038);
and U3739 (N_3739,N_2854,N_2464);
and U3740 (N_3740,N_2486,N_2228);
nor U3741 (N_3741,N_2841,N_2891);
or U3742 (N_3742,N_2170,N_2471);
nor U3743 (N_3743,N_2070,N_2373);
nand U3744 (N_3744,N_2028,N_2065);
xor U3745 (N_3745,N_2254,N_2005);
nor U3746 (N_3746,N_2722,N_2173);
or U3747 (N_3747,N_2631,N_2630);
nor U3748 (N_3748,N_2922,N_2189);
or U3749 (N_3749,N_2505,N_2687);
nand U3750 (N_3750,N_2626,N_2262);
and U3751 (N_3751,N_2426,N_2957);
and U3752 (N_3752,N_2975,N_2931);
xnor U3753 (N_3753,N_2798,N_2781);
nor U3754 (N_3754,N_2841,N_2319);
or U3755 (N_3755,N_2036,N_2845);
nand U3756 (N_3756,N_2439,N_2357);
or U3757 (N_3757,N_2579,N_2553);
nand U3758 (N_3758,N_2907,N_2959);
or U3759 (N_3759,N_2759,N_2579);
and U3760 (N_3760,N_2611,N_2765);
nand U3761 (N_3761,N_2510,N_2379);
or U3762 (N_3762,N_2733,N_2513);
nor U3763 (N_3763,N_2373,N_2910);
nor U3764 (N_3764,N_2054,N_2400);
nand U3765 (N_3765,N_2706,N_2680);
and U3766 (N_3766,N_2470,N_2225);
nor U3767 (N_3767,N_2896,N_2914);
xnor U3768 (N_3768,N_2740,N_2246);
nand U3769 (N_3769,N_2265,N_2962);
nand U3770 (N_3770,N_2579,N_2975);
nand U3771 (N_3771,N_2368,N_2886);
xnor U3772 (N_3772,N_2201,N_2996);
and U3773 (N_3773,N_2593,N_2324);
nor U3774 (N_3774,N_2840,N_2461);
or U3775 (N_3775,N_2926,N_2920);
nand U3776 (N_3776,N_2188,N_2716);
nor U3777 (N_3777,N_2793,N_2987);
and U3778 (N_3778,N_2689,N_2222);
nand U3779 (N_3779,N_2031,N_2339);
and U3780 (N_3780,N_2219,N_2185);
nor U3781 (N_3781,N_2215,N_2601);
nor U3782 (N_3782,N_2999,N_2238);
nand U3783 (N_3783,N_2895,N_2352);
or U3784 (N_3784,N_2177,N_2176);
and U3785 (N_3785,N_2778,N_2956);
nor U3786 (N_3786,N_2207,N_2998);
and U3787 (N_3787,N_2492,N_2351);
and U3788 (N_3788,N_2582,N_2849);
nand U3789 (N_3789,N_2793,N_2734);
nor U3790 (N_3790,N_2658,N_2264);
and U3791 (N_3791,N_2963,N_2058);
or U3792 (N_3792,N_2181,N_2151);
nor U3793 (N_3793,N_2782,N_2061);
and U3794 (N_3794,N_2413,N_2127);
nor U3795 (N_3795,N_2277,N_2073);
or U3796 (N_3796,N_2277,N_2057);
and U3797 (N_3797,N_2480,N_2099);
or U3798 (N_3798,N_2438,N_2699);
and U3799 (N_3799,N_2751,N_2305);
and U3800 (N_3800,N_2248,N_2371);
nand U3801 (N_3801,N_2274,N_2626);
or U3802 (N_3802,N_2240,N_2995);
nand U3803 (N_3803,N_2624,N_2474);
nand U3804 (N_3804,N_2756,N_2917);
nor U3805 (N_3805,N_2150,N_2323);
or U3806 (N_3806,N_2476,N_2094);
or U3807 (N_3807,N_2713,N_2236);
nand U3808 (N_3808,N_2222,N_2526);
and U3809 (N_3809,N_2121,N_2832);
nor U3810 (N_3810,N_2095,N_2329);
and U3811 (N_3811,N_2696,N_2780);
nor U3812 (N_3812,N_2188,N_2220);
nor U3813 (N_3813,N_2478,N_2602);
and U3814 (N_3814,N_2115,N_2587);
nand U3815 (N_3815,N_2845,N_2144);
or U3816 (N_3816,N_2699,N_2792);
nor U3817 (N_3817,N_2843,N_2808);
or U3818 (N_3818,N_2523,N_2977);
nand U3819 (N_3819,N_2279,N_2572);
nand U3820 (N_3820,N_2993,N_2947);
nand U3821 (N_3821,N_2951,N_2118);
nand U3822 (N_3822,N_2318,N_2603);
nand U3823 (N_3823,N_2640,N_2561);
and U3824 (N_3824,N_2601,N_2859);
and U3825 (N_3825,N_2540,N_2964);
or U3826 (N_3826,N_2531,N_2822);
nand U3827 (N_3827,N_2475,N_2365);
nor U3828 (N_3828,N_2895,N_2060);
nand U3829 (N_3829,N_2710,N_2451);
and U3830 (N_3830,N_2262,N_2372);
nand U3831 (N_3831,N_2800,N_2600);
nand U3832 (N_3832,N_2087,N_2492);
nor U3833 (N_3833,N_2092,N_2928);
and U3834 (N_3834,N_2997,N_2319);
and U3835 (N_3835,N_2280,N_2008);
nor U3836 (N_3836,N_2673,N_2289);
nand U3837 (N_3837,N_2708,N_2574);
and U3838 (N_3838,N_2669,N_2819);
or U3839 (N_3839,N_2850,N_2884);
nand U3840 (N_3840,N_2004,N_2542);
and U3841 (N_3841,N_2950,N_2544);
or U3842 (N_3842,N_2093,N_2591);
nor U3843 (N_3843,N_2981,N_2533);
and U3844 (N_3844,N_2071,N_2703);
and U3845 (N_3845,N_2299,N_2561);
and U3846 (N_3846,N_2385,N_2978);
nor U3847 (N_3847,N_2892,N_2480);
or U3848 (N_3848,N_2586,N_2053);
nor U3849 (N_3849,N_2965,N_2204);
or U3850 (N_3850,N_2214,N_2366);
nor U3851 (N_3851,N_2644,N_2983);
nand U3852 (N_3852,N_2314,N_2214);
and U3853 (N_3853,N_2648,N_2534);
nor U3854 (N_3854,N_2042,N_2231);
and U3855 (N_3855,N_2702,N_2705);
nor U3856 (N_3856,N_2302,N_2867);
and U3857 (N_3857,N_2007,N_2207);
and U3858 (N_3858,N_2368,N_2992);
and U3859 (N_3859,N_2846,N_2719);
or U3860 (N_3860,N_2380,N_2296);
and U3861 (N_3861,N_2364,N_2165);
or U3862 (N_3862,N_2060,N_2852);
and U3863 (N_3863,N_2613,N_2456);
or U3864 (N_3864,N_2856,N_2376);
and U3865 (N_3865,N_2906,N_2530);
and U3866 (N_3866,N_2372,N_2632);
nand U3867 (N_3867,N_2552,N_2888);
and U3868 (N_3868,N_2712,N_2726);
nand U3869 (N_3869,N_2889,N_2728);
or U3870 (N_3870,N_2665,N_2993);
nand U3871 (N_3871,N_2757,N_2045);
or U3872 (N_3872,N_2524,N_2227);
nand U3873 (N_3873,N_2486,N_2295);
or U3874 (N_3874,N_2258,N_2966);
or U3875 (N_3875,N_2389,N_2031);
xor U3876 (N_3876,N_2780,N_2840);
nand U3877 (N_3877,N_2626,N_2811);
or U3878 (N_3878,N_2266,N_2368);
and U3879 (N_3879,N_2786,N_2640);
or U3880 (N_3880,N_2481,N_2388);
nor U3881 (N_3881,N_2259,N_2407);
nor U3882 (N_3882,N_2733,N_2325);
and U3883 (N_3883,N_2502,N_2080);
or U3884 (N_3884,N_2931,N_2775);
and U3885 (N_3885,N_2938,N_2966);
and U3886 (N_3886,N_2351,N_2200);
nand U3887 (N_3887,N_2331,N_2726);
nor U3888 (N_3888,N_2592,N_2617);
or U3889 (N_3889,N_2132,N_2585);
or U3890 (N_3890,N_2706,N_2809);
nand U3891 (N_3891,N_2202,N_2819);
nand U3892 (N_3892,N_2511,N_2708);
nor U3893 (N_3893,N_2325,N_2743);
and U3894 (N_3894,N_2574,N_2952);
and U3895 (N_3895,N_2916,N_2247);
or U3896 (N_3896,N_2246,N_2442);
nor U3897 (N_3897,N_2139,N_2398);
and U3898 (N_3898,N_2043,N_2099);
or U3899 (N_3899,N_2474,N_2564);
nand U3900 (N_3900,N_2623,N_2636);
and U3901 (N_3901,N_2632,N_2907);
or U3902 (N_3902,N_2189,N_2505);
nand U3903 (N_3903,N_2956,N_2780);
and U3904 (N_3904,N_2461,N_2126);
and U3905 (N_3905,N_2183,N_2740);
and U3906 (N_3906,N_2528,N_2591);
or U3907 (N_3907,N_2868,N_2531);
nand U3908 (N_3908,N_2244,N_2171);
nor U3909 (N_3909,N_2983,N_2441);
and U3910 (N_3910,N_2589,N_2036);
or U3911 (N_3911,N_2503,N_2698);
nor U3912 (N_3912,N_2201,N_2076);
or U3913 (N_3913,N_2673,N_2886);
nand U3914 (N_3914,N_2629,N_2696);
xnor U3915 (N_3915,N_2025,N_2959);
nand U3916 (N_3916,N_2296,N_2064);
and U3917 (N_3917,N_2914,N_2034);
nand U3918 (N_3918,N_2266,N_2270);
nand U3919 (N_3919,N_2539,N_2445);
and U3920 (N_3920,N_2494,N_2922);
and U3921 (N_3921,N_2048,N_2367);
nor U3922 (N_3922,N_2910,N_2825);
nand U3923 (N_3923,N_2390,N_2374);
nand U3924 (N_3924,N_2550,N_2033);
and U3925 (N_3925,N_2361,N_2006);
or U3926 (N_3926,N_2316,N_2372);
or U3927 (N_3927,N_2275,N_2235);
nand U3928 (N_3928,N_2434,N_2287);
nor U3929 (N_3929,N_2192,N_2381);
nand U3930 (N_3930,N_2866,N_2371);
or U3931 (N_3931,N_2614,N_2194);
or U3932 (N_3932,N_2889,N_2497);
nand U3933 (N_3933,N_2889,N_2273);
or U3934 (N_3934,N_2297,N_2676);
and U3935 (N_3935,N_2819,N_2227);
nand U3936 (N_3936,N_2418,N_2812);
nor U3937 (N_3937,N_2315,N_2866);
nand U3938 (N_3938,N_2741,N_2319);
and U3939 (N_3939,N_2105,N_2390);
nor U3940 (N_3940,N_2641,N_2665);
or U3941 (N_3941,N_2006,N_2783);
and U3942 (N_3942,N_2605,N_2337);
nor U3943 (N_3943,N_2029,N_2626);
nor U3944 (N_3944,N_2483,N_2038);
and U3945 (N_3945,N_2782,N_2896);
and U3946 (N_3946,N_2752,N_2935);
or U3947 (N_3947,N_2827,N_2908);
or U3948 (N_3948,N_2168,N_2521);
nand U3949 (N_3949,N_2569,N_2343);
nor U3950 (N_3950,N_2865,N_2698);
nor U3951 (N_3951,N_2439,N_2778);
nor U3952 (N_3952,N_2019,N_2796);
nand U3953 (N_3953,N_2814,N_2622);
and U3954 (N_3954,N_2405,N_2173);
or U3955 (N_3955,N_2541,N_2001);
nor U3956 (N_3956,N_2762,N_2249);
nand U3957 (N_3957,N_2909,N_2250);
or U3958 (N_3958,N_2835,N_2794);
nor U3959 (N_3959,N_2194,N_2770);
or U3960 (N_3960,N_2998,N_2241);
nor U3961 (N_3961,N_2335,N_2850);
and U3962 (N_3962,N_2637,N_2659);
and U3963 (N_3963,N_2624,N_2318);
or U3964 (N_3964,N_2551,N_2582);
and U3965 (N_3965,N_2429,N_2817);
or U3966 (N_3966,N_2588,N_2991);
nand U3967 (N_3967,N_2932,N_2697);
and U3968 (N_3968,N_2286,N_2662);
and U3969 (N_3969,N_2436,N_2736);
and U3970 (N_3970,N_2409,N_2543);
or U3971 (N_3971,N_2521,N_2214);
nor U3972 (N_3972,N_2733,N_2543);
or U3973 (N_3973,N_2551,N_2052);
and U3974 (N_3974,N_2146,N_2604);
nand U3975 (N_3975,N_2595,N_2745);
and U3976 (N_3976,N_2208,N_2926);
or U3977 (N_3977,N_2322,N_2968);
or U3978 (N_3978,N_2552,N_2317);
or U3979 (N_3979,N_2211,N_2059);
nor U3980 (N_3980,N_2148,N_2420);
nor U3981 (N_3981,N_2871,N_2247);
or U3982 (N_3982,N_2488,N_2853);
or U3983 (N_3983,N_2768,N_2463);
and U3984 (N_3984,N_2214,N_2892);
or U3985 (N_3985,N_2634,N_2972);
or U3986 (N_3986,N_2194,N_2258);
or U3987 (N_3987,N_2412,N_2435);
or U3988 (N_3988,N_2507,N_2813);
and U3989 (N_3989,N_2351,N_2955);
or U3990 (N_3990,N_2345,N_2260);
nand U3991 (N_3991,N_2941,N_2151);
and U3992 (N_3992,N_2309,N_2274);
nand U3993 (N_3993,N_2810,N_2237);
nor U3994 (N_3994,N_2921,N_2156);
or U3995 (N_3995,N_2721,N_2522);
and U3996 (N_3996,N_2488,N_2104);
nor U3997 (N_3997,N_2975,N_2725);
or U3998 (N_3998,N_2183,N_2513);
nand U3999 (N_3999,N_2963,N_2319);
and U4000 (N_4000,N_3176,N_3343);
nor U4001 (N_4001,N_3779,N_3399);
nor U4002 (N_4002,N_3152,N_3339);
nand U4003 (N_4003,N_3356,N_3693);
nand U4004 (N_4004,N_3467,N_3436);
nor U4005 (N_4005,N_3081,N_3409);
nand U4006 (N_4006,N_3417,N_3931);
and U4007 (N_4007,N_3868,N_3673);
nand U4008 (N_4008,N_3963,N_3287);
nand U4009 (N_4009,N_3443,N_3117);
and U4010 (N_4010,N_3752,N_3217);
nor U4011 (N_4011,N_3090,N_3428);
and U4012 (N_4012,N_3555,N_3880);
or U4013 (N_4013,N_3448,N_3233);
and U4014 (N_4014,N_3910,N_3114);
nor U4015 (N_4015,N_3122,N_3519);
nor U4016 (N_4016,N_3213,N_3145);
or U4017 (N_4017,N_3241,N_3645);
and U4018 (N_4018,N_3707,N_3008);
nand U4019 (N_4019,N_3030,N_3984);
nor U4020 (N_4020,N_3071,N_3049);
or U4021 (N_4021,N_3418,N_3192);
nor U4022 (N_4022,N_3067,N_3063);
and U4023 (N_4023,N_3115,N_3004);
nand U4024 (N_4024,N_3949,N_3198);
nand U4025 (N_4025,N_3991,N_3812);
nor U4026 (N_4026,N_3980,N_3825);
and U4027 (N_4027,N_3348,N_3832);
or U4028 (N_4028,N_3018,N_3043);
nor U4029 (N_4029,N_3225,N_3613);
or U4030 (N_4030,N_3912,N_3402);
and U4031 (N_4031,N_3531,N_3572);
nand U4032 (N_4032,N_3316,N_3829);
nand U4033 (N_4033,N_3777,N_3580);
or U4034 (N_4034,N_3332,N_3838);
or U4035 (N_4035,N_3655,N_3070);
or U4036 (N_4036,N_3657,N_3643);
nand U4037 (N_4037,N_3535,N_3794);
and U4038 (N_4038,N_3651,N_3710);
nand U4039 (N_4039,N_3729,N_3895);
nand U4040 (N_4040,N_3042,N_3826);
and U4041 (N_4041,N_3512,N_3843);
nor U4042 (N_4042,N_3987,N_3060);
or U4043 (N_4043,N_3038,N_3040);
nand U4044 (N_4044,N_3876,N_3334);
and U4045 (N_4045,N_3559,N_3622);
and U4046 (N_4046,N_3670,N_3249);
or U4047 (N_4047,N_3215,N_3956);
nor U4048 (N_4048,N_3692,N_3890);
nand U4049 (N_4049,N_3297,N_3301);
and U4050 (N_4050,N_3100,N_3412);
or U4051 (N_4051,N_3682,N_3022);
or U4052 (N_4052,N_3097,N_3032);
or U4053 (N_4053,N_3863,N_3222);
or U4054 (N_4054,N_3260,N_3716);
or U4055 (N_4055,N_3495,N_3755);
and U4056 (N_4056,N_3615,N_3545);
nand U4057 (N_4057,N_3474,N_3437);
nand U4058 (N_4058,N_3484,N_3477);
nor U4059 (N_4059,N_3274,N_3568);
nand U4060 (N_4060,N_3886,N_3885);
and U4061 (N_4061,N_3524,N_3556);
or U4062 (N_4062,N_3375,N_3034);
and U4063 (N_4063,N_3313,N_3468);
or U4064 (N_4064,N_3749,N_3363);
nand U4065 (N_4065,N_3259,N_3626);
nor U4066 (N_4066,N_3658,N_3244);
nor U4067 (N_4067,N_3093,N_3677);
nor U4068 (N_4068,N_3841,N_3862);
or U4069 (N_4069,N_3698,N_3456);
or U4070 (N_4070,N_3455,N_3216);
nor U4071 (N_4071,N_3857,N_3517);
and U4072 (N_4072,N_3754,N_3257);
or U4073 (N_4073,N_3158,N_3609);
and U4074 (N_4074,N_3684,N_3634);
nor U4075 (N_4075,N_3187,N_3449);
and U4076 (N_4076,N_3065,N_3667);
nor U4077 (N_4077,N_3662,N_3708);
and U4078 (N_4078,N_3939,N_3828);
or U4079 (N_4079,N_3785,N_3091);
nor U4080 (N_4080,N_3272,N_3028);
and U4081 (N_4081,N_3011,N_3324);
and U4082 (N_4082,N_3346,N_3033);
nand U4083 (N_4083,N_3240,N_3269);
nand U4084 (N_4084,N_3665,N_3689);
nor U4085 (N_4085,N_3413,N_3731);
or U4086 (N_4086,N_3041,N_3848);
or U4087 (N_4087,N_3523,N_3219);
nand U4088 (N_4088,N_3965,N_3566);
nand U4089 (N_4089,N_3958,N_3354);
nor U4090 (N_4090,N_3914,N_3702);
or U4091 (N_4091,N_3636,N_3864);
nand U4092 (N_4092,N_3239,N_3952);
or U4093 (N_4093,N_3232,N_3170);
and U4094 (N_4094,N_3440,N_3483);
nand U4095 (N_4095,N_3036,N_3954);
and U4096 (N_4096,N_3314,N_3600);
and U4097 (N_4097,N_3140,N_3015);
nand U4098 (N_4098,N_3288,N_3768);
and U4099 (N_4099,N_3327,N_3389);
nand U4100 (N_4100,N_3398,N_3770);
nand U4101 (N_4101,N_3979,N_3948);
nor U4102 (N_4102,N_3978,N_3167);
nand U4103 (N_4103,N_3128,N_3421);
nand U4104 (N_4104,N_3915,N_3195);
nand U4105 (N_4105,N_3641,N_3672);
nand U4106 (N_4106,N_3317,N_3501);
nand U4107 (N_4107,N_3019,N_3762);
nor U4108 (N_4108,N_3784,N_3905);
nand U4109 (N_4109,N_3967,N_3388);
and U4110 (N_4110,N_3407,N_3526);
nand U4111 (N_4111,N_3059,N_3942);
and U4112 (N_4112,N_3599,N_3154);
or U4113 (N_4113,N_3552,N_3510);
or U4114 (N_4114,N_3532,N_3514);
xor U4115 (N_4115,N_3722,N_3685);
nor U4116 (N_4116,N_3284,N_3300);
nor U4117 (N_4117,N_3189,N_3352);
nand U4118 (N_4118,N_3380,N_3183);
nor U4119 (N_4119,N_3224,N_3810);
nand U4120 (N_4120,N_3445,N_3344);
or U4121 (N_4121,N_3002,N_3659);
or U4122 (N_4122,N_3271,N_3452);
and U4123 (N_4123,N_3783,N_3386);
nand U4124 (N_4124,N_3226,N_3111);
nand U4125 (N_4125,N_3856,N_3404);
and U4126 (N_4126,N_3121,N_3738);
xor U4127 (N_4127,N_3598,N_3906);
nand U4128 (N_4128,N_3577,N_3267);
and U4129 (N_4129,N_3927,N_3372);
nor U4130 (N_4130,N_3441,N_3602);
and U4131 (N_4131,N_3899,N_3424);
or U4132 (N_4132,N_3887,N_3465);
nand U4133 (N_4133,N_3697,N_3660);
xor U4134 (N_4134,N_3020,N_3279);
or U4135 (N_4135,N_3747,N_3878);
or U4136 (N_4136,N_3462,N_3359);
nor U4137 (N_4137,N_3262,N_3891);
nand U4138 (N_4138,N_3291,N_3368);
nand U4139 (N_4139,N_3955,N_3370);
or U4140 (N_4140,N_3083,N_3335);
and U4141 (N_4141,N_3503,N_3540);
or U4142 (N_4142,N_3666,N_3023);
or U4143 (N_4143,N_3246,N_3801);
nand U4144 (N_4144,N_3454,N_3098);
nand U4145 (N_4145,N_3296,N_3108);
nor U4146 (N_4146,N_3661,N_3024);
nand U4147 (N_4147,N_3079,N_3029);
and U4148 (N_4148,N_3750,N_3678);
and U4149 (N_4149,N_3896,N_3254);
nand U4150 (N_4150,N_3096,N_3101);
and U4151 (N_4151,N_3706,N_3074);
and U4152 (N_4152,N_3649,N_3295);
and U4153 (N_4153,N_3076,N_3406);
nand U4154 (N_4154,N_3650,N_3574);
nand U4155 (N_4155,N_3051,N_3423);
or U4156 (N_4156,N_3203,N_3381);
nand U4157 (N_4157,N_3957,N_3793);
and U4158 (N_4158,N_3819,N_3557);
nor U4159 (N_4159,N_3582,N_3941);
nor U4160 (N_4160,N_3333,N_3099);
or U4161 (N_4161,N_3564,N_3875);
nand U4162 (N_4162,N_3165,N_3851);
nor U4163 (N_4163,N_3610,N_3797);
or U4164 (N_4164,N_3457,N_3476);
nor U4165 (N_4165,N_3720,N_3253);
nor U4166 (N_4166,N_3080,N_3827);
or U4167 (N_4167,N_3237,N_3990);
or U4168 (N_4168,N_3579,N_3005);
nor U4169 (N_4169,N_3328,N_3596);
nand U4170 (N_4170,N_3902,N_3498);
nand U4171 (N_4171,N_3881,N_3761);
nand U4172 (N_4172,N_3153,N_3811);
nand U4173 (N_4173,N_3379,N_3478);
nand U4174 (N_4174,N_3593,N_3844);
or U4175 (N_4175,N_3904,N_3713);
nand U4176 (N_4176,N_3143,N_3823);
or U4177 (N_4177,N_3178,N_3200);
or U4178 (N_4178,N_3017,N_3394);
nand U4179 (N_4179,N_3617,N_3936);
nor U4180 (N_4180,N_3620,N_3687);
nand U4181 (N_4181,N_3135,N_3860);
and U4182 (N_4182,N_3282,N_3161);
and U4183 (N_4183,N_3182,N_3491);
nand U4184 (N_4184,N_3934,N_3137);
or U4185 (N_4185,N_3681,N_3275);
or U4186 (N_4186,N_3603,N_3536);
or U4187 (N_4187,N_3383,N_3930);
xnor U4188 (N_4188,N_3345,N_3571);
nor U4189 (N_4189,N_3999,N_3387);
nand U4190 (N_4190,N_3543,N_3270);
and U4191 (N_4191,N_3884,N_3576);
or U4192 (N_4192,N_3839,N_3674);
nand U4193 (N_4193,N_3903,N_3125);
nand U4194 (N_4194,N_3351,N_3094);
or U4195 (N_4195,N_3741,N_3730);
nand U4196 (N_4196,N_3116,N_3278);
or U4197 (N_4197,N_3146,N_3765);
and U4198 (N_4198,N_3138,N_3385);
nor U4199 (N_4199,N_3767,N_3554);
or U4200 (N_4200,N_3846,N_3102);
or U4201 (N_4201,N_3181,N_3590);
nor U4202 (N_4202,N_3711,N_3416);
and U4203 (N_4203,N_3961,N_3236);
and U4204 (N_4204,N_3243,N_3330);
or U4205 (N_4205,N_3774,N_3302);
or U4206 (N_4206,N_3893,N_3326);
or U4207 (N_4207,N_3155,N_3037);
and U4208 (N_4208,N_3888,N_3364);
or U4209 (N_4209,N_3220,N_3366);
nor U4210 (N_4210,N_3671,N_3721);
and U4211 (N_4211,N_3814,N_3513);
and U4212 (N_4212,N_3923,N_3358);
and U4213 (N_4213,N_3276,N_3892);
nand U4214 (N_4214,N_3141,N_3522);
or U4215 (N_4215,N_3818,N_3917);
or U4216 (N_4216,N_3132,N_3601);
or U4217 (N_4217,N_3807,N_3401);
nand U4218 (N_4218,N_3901,N_3186);
nand U4219 (N_4219,N_3759,N_3969);
nand U4220 (N_4220,N_3305,N_3668);
nand U4221 (N_4221,N_3322,N_3573);
and U4222 (N_4222,N_3319,N_3231);
or U4223 (N_4223,N_3057,N_3450);
nand U4224 (N_4224,N_3430,N_3422);
nor U4225 (N_4225,N_3369,N_3427);
or U4226 (N_4226,N_3870,N_3073);
nand U4227 (N_4227,N_3644,N_3981);
and U4228 (N_4228,N_3908,N_3800);
or U4229 (N_4229,N_3494,N_3337);
nor U4230 (N_4230,N_3925,N_3792);
nor U4231 (N_4231,N_3039,N_3391);
and U4232 (N_4232,N_3197,N_3194);
nand U4233 (N_4233,N_3410,N_3320);
nand U4234 (N_4234,N_3932,N_3016);
or U4235 (N_4235,N_3873,N_3638);
or U4236 (N_4236,N_3069,N_3553);
nand U4237 (N_4237,N_3718,N_3632);
or U4238 (N_4238,N_3970,N_3791);
or U4239 (N_4239,N_3919,N_3624);
nor U4240 (N_4240,N_3775,N_3837);
nor U4241 (N_4241,N_3298,N_3946);
or U4242 (N_4242,N_3530,N_3469);
or U4243 (N_4243,N_3499,N_3355);
nand U4244 (N_4244,N_3458,N_3382);
nor U4245 (N_4245,N_3508,N_3653);
nand U4246 (N_4246,N_3971,N_3336);
and U4247 (N_4247,N_3118,N_3854);
nand U4248 (N_4248,N_3180,N_3778);
or U4249 (N_4249,N_3594,N_3373);
or U4250 (N_4250,N_3447,N_3196);
or U4251 (N_4251,N_3585,N_3120);
or U4252 (N_4252,N_3309,N_3432);
nor U4253 (N_4253,N_3694,N_3078);
nand U4254 (N_4254,N_3633,N_3238);
or U4255 (N_4255,N_3877,N_3086);
nand U4256 (N_4256,N_3497,N_3329);
nand U4257 (N_4257,N_3605,N_3547);
and U4258 (N_4258,N_3966,N_3907);
nand U4259 (N_4259,N_3312,N_3006);
or U4260 (N_4260,N_3273,N_3280);
nor U4261 (N_4261,N_3075,N_3975);
or U4262 (N_4262,N_3546,N_3533);
nor U4263 (N_4263,N_3157,N_3725);
or U4264 (N_4264,N_3227,N_3110);
or U4265 (N_4265,N_3266,N_3490);
and U4266 (N_4266,N_3538,N_3340);
or U4267 (N_4267,N_3177,N_3699);
nor U4268 (N_4268,N_3611,N_3371);
or U4269 (N_4269,N_3053,N_3799);
and U4270 (N_4270,N_3938,N_3010);
nand U4271 (N_4271,N_3124,N_3054);
or U4272 (N_4272,N_3511,N_3353);
and U4273 (N_4273,N_3940,N_3787);
nand U4274 (N_4274,N_3664,N_3365);
nor U4275 (N_4275,N_3813,N_3680);
and U4276 (N_4276,N_3719,N_3631);
and U4277 (N_4277,N_3935,N_3400);
or U4278 (N_4278,N_3728,N_3607);
or U4279 (N_4279,N_3518,N_3669);
nor U4280 (N_4280,N_3968,N_3460);
nor U4281 (N_4281,N_3026,N_3000);
or U4282 (N_4282,N_3520,N_3204);
nand U4283 (N_4283,N_3567,N_3616);
and U4284 (N_4284,N_3147,N_3342);
nor U4285 (N_4285,N_3926,N_3898);
or U4286 (N_4286,N_3207,N_3943);
or U4287 (N_4287,N_3816,N_3265);
and U4288 (N_4288,N_3129,N_3855);
nor U4289 (N_4289,N_3845,N_3835);
or U4290 (N_4290,N_3894,N_3909);
and U4291 (N_4291,N_3009,N_3804);
or U4292 (N_4292,N_3727,N_3690);
nand U4293 (N_4293,N_3321,N_3998);
and U4294 (N_4294,N_3255,N_3229);
and U4295 (N_4295,N_3127,N_3960);
and U4296 (N_4296,N_3031,N_3676);
nor U4297 (N_4297,N_3639,N_3209);
nand U4298 (N_4298,N_3548,N_3318);
and U4299 (N_4299,N_3056,N_3871);
or U4300 (N_4300,N_3534,N_3874);
nand U4301 (N_4301,N_3679,N_3842);
and U4302 (N_4302,N_3304,N_3426);
nor U4303 (N_4303,N_3922,N_3612);
or U4304 (N_4304,N_3072,N_3223);
or U4305 (N_4305,N_3867,N_3836);
or U4306 (N_4306,N_3789,N_3463);
nor U4307 (N_4307,N_3654,N_3743);
and U4308 (N_4308,N_3377,N_3766);
nor U4309 (N_4309,N_3084,N_3614);
nand U4310 (N_4310,N_3865,N_3390);
and U4311 (N_4311,N_3630,N_3431);
nand U4312 (N_4312,N_3989,N_3395);
nand U4313 (N_4313,N_3289,N_3502);
and U4314 (N_4314,N_3185,N_3840);
xnor U4315 (N_4315,N_3188,N_3994);
or U4316 (N_4316,N_3261,N_3481);
and U4317 (N_4317,N_3983,N_3055);
nor U4318 (N_4318,N_3361,N_3234);
nor U4319 (N_4319,N_3803,N_3723);
nor U4320 (N_4320,N_3809,N_3558);
nand U4321 (N_4321,N_3061,N_3944);
nand U4322 (N_4322,N_3853,N_3193);
nand U4323 (N_4323,N_3976,N_3263);
or U4324 (N_4324,N_3264,N_3347);
nor U4325 (N_4325,N_3753,N_3168);
and U4326 (N_4326,N_3806,N_3808);
nand U4327 (N_4327,N_3516,N_3166);
or U4328 (N_4328,N_3703,N_3866);
or U4329 (N_4329,N_3795,N_3734);
nor U4330 (N_4330,N_3001,N_3105);
or U4331 (N_4331,N_3190,N_3509);
nand U4332 (N_4332,N_3591,N_3306);
nor U4333 (N_4333,N_3924,N_3782);
and U4334 (N_4334,N_3788,N_3824);
nand U4335 (N_4335,N_3208,N_3648);
and U4336 (N_4336,N_3174,N_3357);
or U4337 (N_4337,N_3142,N_3500);
or U4338 (N_4338,N_3315,N_3565);
or U4339 (N_4339,N_3542,N_3737);
nand U4340 (N_4340,N_3821,N_3618);
and U4341 (N_4341,N_3982,N_3937);
and U4342 (N_4342,N_3663,N_3066);
nor U4343 (N_4343,N_3169,N_3014);
nand U4344 (N_4344,N_3858,N_3179);
and U4345 (N_4345,N_3106,N_3701);
nor U4346 (N_4346,N_3092,N_3763);
nor U4347 (N_4347,N_3488,N_3472);
nor U4348 (N_4348,N_3714,N_3696);
nand U4349 (N_4349,N_3833,N_3496);
nand U4350 (N_4350,N_3642,N_3506);
or U4351 (N_4351,N_3191,N_3505);
nand U4352 (N_4352,N_3581,N_3739);
and U4353 (N_4353,N_3012,N_3376);
nand U4354 (N_4354,N_3830,N_3726);
or U4355 (N_4355,N_3466,N_3139);
and U4356 (N_4356,N_3293,N_3977);
and U4357 (N_4357,N_3308,N_3485);
nor U4358 (N_4358,N_3992,N_3479);
nand U4359 (N_4359,N_3281,N_3433);
and U4360 (N_4360,N_3715,N_3974);
or U4361 (N_4361,N_3211,N_3815);
nand U4362 (N_4362,N_3805,N_3918);
nor U4363 (N_4363,N_3847,N_3349);
nand U4364 (N_4364,N_3640,N_3544);
nand U4365 (N_4365,N_3290,N_3521);
or U4366 (N_4366,N_3095,N_3088);
nand U4367 (N_4367,N_3882,N_3492);
nand U4368 (N_4368,N_3541,N_3341);
or U4369 (N_4369,N_3442,N_3212);
nor U4370 (N_4370,N_3995,N_3628);
nand U4371 (N_4371,N_3587,N_3251);
nand U4372 (N_4372,N_3798,N_3705);
nand U4373 (N_4373,N_3820,N_3772);
nor U4374 (N_4374,N_3951,N_3629);
nor U4375 (N_4375,N_3163,N_3563);
nor U4376 (N_4376,N_3068,N_3414);
nor U4377 (N_4377,N_3872,N_3786);
and U4378 (N_4378,N_3164,N_3757);
and U4379 (N_4379,N_3360,N_3688);
and U4380 (N_4380,N_3286,N_3586);
nand U4381 (N_4381,N_3046,N_3691);
or U4382 (N_4382,N_3746,N_3796);
and U4383 (N_4383,N_3735,N_3113);
nand U4384 (N_4384,N_3627,N_3461);
and U4385 (N_4385,N_3686,N_3635);
or U4386 (N_4386,N_3700,N_3712);
and U4387 (N_4387,N_3184,N_3338);
and U4388 (N_4388,N_3964,N_3972);
or U4389 (N_4389,N_3575,N_3742);
nand U4390 (N_4390,N_3569,N_3393);
or U4391 (N_4391,N_3199,N_3962);
nor U4392 (N_4392,N_3045,N_3578);
or U4393 (N_4393,N_3527,N_3003);
or U4394 (N_4394,N_3780,N_3210);
or U4395 (N_4395,N_3405,N_3048);
nand U4396 (N_4396,N_3583,N_3459);
and U4397 (N_4397,N_3299,N_3160);
and U4398 (N_4398,N_3378,N_3156);
nand U4399 (N_4399,N_3119,N_3294);
or U4400 (N_4400,N_3027,N_3256);
nor U4401 (N_4401,N_3126,N_3769);
nor U4402 (N_4402,N_3529,N_3159);
nor U4403 (N_4403,N_3362,N_3850);
or U4404 (N_4404,N_3717,N_3621);
nor U4405 (N_4405,N_3756,N_3250);
nand U4406 (N_4406,N_3745,N_3751);
or U4407 (N_4407,N_3062,N_3525);
or U4408 (N_4408,N_3570,N_3415);
and U4409 (N_4409,N_3050,N_3539);
or U4410 (N_4410,N_3367,N_3151);
nor U4411 (N_4411,N_3047,N_3471);
nand U4412 (N_4412,N_3764,N_3446);
or U4413 (N_4413,N_3709,N_3331);
or U4414 (N_4414,N_3451,N_3307);
nor U4415 (N_4415,N_3425,N_3150);
and U4416 (N_4416,N_3311,N_3285);
nor U4417 (N_4417,N_3384,N_3292);
nand U4418 (N_4418,N_3704,N_3869);
nand U4419 (N_4419,N_3453,N_3831);
and U4420 (N_4420,N_3760,N_3235);
nor U4421 (N_4421,N_3144,N_3439);
or U4422 (N_4422,N_3131,N_3724);
nand U4423 (N_4423,N_3549,N_3172);
nor U4424 (N_4424,N_3619,N_3584);
nor U4425 (N_4425,N_3148,N_3652);
or U4426 (N_4426,N_3077,N_3064);
nor U4427 (N_4427,N_3277,N_3776);
or U4428 (N_4428,N_3434,N_3646);
nor U4429 (N_4429,N_3112,N_3911);
and U4430 (N_4430,N_3171,N_3861);
nand U4431 (N_4431,N_3350,N_3258);
or U4432 (N_4432,N_3859,N_3419);
and U4433 (N_4433,N_3913,N_3104);
and U4434 (N_4434,N_3218,N_3675);
xnor U4435 (N_4435,N_3044,N_3996);
nor U4436 (N_4436,N_3493,N_3173);
or U4437 (N_4437,N_3201,N_3647);
nand U4438 (N_4438,N_3988,N_3900);
nand U4439 (N_4439,N_3597,N_3103);
nand U4440 (N_4440,N_3959,N_3397);
nand U4441 (N_4441,N_3849,N_3879);
nand U4442 (N_4442,N_3695,N_3515);
nor U4443 (N_4443,N_3561,N_3834);
nor U4444 (N_4444,N_3920,N_3758);
nand U4445 (N_4445,N_3637,N_3087);
or U4446 (N_4446,N_3162,N_3268);
nor U4447 (N_4447,N_3921,N_3134);
and U4448 (N_4448,N_3435,N_3058);
and U4449 (N_4449,N_3464,N_3592);
nor U4450 (N_4450,N_3656,N_3985);
or U4451 (N_4451,N_3802,N_3480);
nand U4452 (N_4452,N_3748,N_3623);
or U4453 (N_4453,N_3973,N_3403);
nand U4454 (N_4454,N_3470,N_3475);
nor U4455 (N_4455,N_3740,N_3408);
and U4456 (N_4456,N_3230,N_3916);
or U4457 (N_4457,N_3109,N_3773);
nand U4458 (N_4458,N_3429,N_3997);
and U4459 (N_4459,N_3252,N_3202);
and U4460 (N_4460,N_3551,N_3438);
nor U4461 (N_4461,N_3822,N_3007);
and U4462 (N_4462,N_3013,N_3929);
nor U4463 (N_4463,N_3221,N_3205);
and U4464 (N_4464,N_3283,N_3528);
or U4465 (N_4465,N_3325,N_3744);
and U4466 (N_4466,N_3487,N_3245);
and U4467 (N_4467,N_3130,N_3149);
xor U4468 (N_4468,N_3608,N_3242);
or U4469 (N_4469,N_3021,N_3247);
or U4470 (N_4470,N_3310,N_3136);
and U4471 (N_4471,N_3206,N_3817);
nor U4472 (N_4472,N_3133,N_3082);
and U4473 (N_4473,N_3486,N_3175);
nand U4474 (N_4474,N_3248,N_3323);
nor U4475 (N_4475,N_3214,N_3897);
and U4476 (N_4476,N_3482,N_3733);
nand U4477 (N_4477,N_3589,N_3562);
or U4478 (N_4478,N_3374,N_3052);
or U4479 (N_4479,N_3560,N_3889);
nor U4480 (N_4480,N_3781,N_3392);
and U4481 (N_4481,N_3411,N_3085);
nand U4482 (N_4482,N_3473,N_3035);
nand U4483 (N_4483,N_3993,N_3736);
and U4484 (N_4484,N_3606,N_3986);
nor U4485 (N_4485,N_3107,N_3945);
nor U4486 (N_4486,N_3025,N_3444);
and U4487 (N_4487,N_3595,N_3588);
nand U4488 (N_4488,N_3947,N_3123);
nand U4489 (N_4489,N_3228,N_3537);
and U4490 (N_4490,N_3489,N_3732);
nand U4491 (N_4491,N_3507,N_3683);
nor U4492 (N_4492,N_3089,N_3625);
nand U4493 (N_4493,N_3396,N_3303);
and U4494 (N_4494,N_3950,N_3953);
and U4495 (N_4495,N_3550,N_3790);
or U4496 (N_4496,N_3928,N_3933);
and U4497 (N_4497,N_3883,N_3771);
and U4498 (N_4498,N_3504,N_3604);
nor U4499 (N_4499,N_3852,N_3420);
or U4500 (N_4500,N_3978,N_3684);
nor U4501 (N_4501,N_3251,N_3483);
or U4502 (N_4502,N_3122,N_3527);
and U4503 (N_4503,N_3256,N_3248);
nor U4504 (N_4504,N_3297,N_3144);
nor U4505 (N_4505,N_3296,N_3983);
nor U4506 (N_4506,N_3870,N_3499);
or U4507 (N_4507,N_3412,N_3226);
and U4508 (N_4508,N_3280,N_3129);
and U4509 (N_4509,N_3888,N_3752);
nand U4510 (N_4510,N_3881,N_3541);
nand U4511 (N_4511,N_3936,N_3963);
nand U4512 (N_4512,N_3954,N_3942);
or U4513 (N_4513,N_3897,N_3457);
and U4514 (N_4514,N_3741,N_3825);
or U4515 (N_4515,N_3315,N_3600);
nand U4516 (N_4516,N_3265,N_3645);
nand U4517 (N_4517,N_3734,N_3612);
or U4518 (N_4518,N_3278,N_3807);
or U4519 (N_4519,N_3077,N_3436);
nand U4520 (N_4520,N_3217,N_3943);
and U4521 (N_4521,N_3069,N_3912);
nand U4522 (N_4522,N_3565,N_3983);
nand U4523 (N_4523,N_3982,N_3447);
and U4524 (N_4524,N_3192,N_3294);
nand U4525 (N_4525,N_3001,N_3801);
and U4526 (N_4526,N_3064,N_3203);
nand U4527 (N_4527,N_3387,N_3849);
nor U4528 (N_4528,N_3324,N_3960);
and U4529 (N_4529,N_3028,N_3517);
nand U4530 (N_4530,N_3206,N_3006);
or U4531 (N_4531,N_3958,N_3929);
nand U4532 (N_4532,N_3907,N_3743);
nand U4533 (N_4533,N_3889,N_3374);
nand U4534 (N_4534,N_3382,N_3908);
nor U4535 (N_4535,N_3042,N_3855);
and U4536 (N_4536,N_3170,N_3292);
nand U4537 (N_4537,N_3402,N_3480);
nand U4538 (N_4538,N_3204,N_3586);
nor U4539 (N_4539,N_3362,N_3749);
nand U4540 (N_4540,N_3022,N_3669);
and U4541 (N_4541,N_3707,N_3386);
nand U4542 (N_4542,N_3351,N_3854);
and U4543 (N_4543,N_3315,N_3162);
xor U4544 (N_4544,N_3360,N_3690);
nand U4545 (N_4545,N_3276,N_3774);
and U4546 (N_4546,N_3170,N_3102);
nor U4547 (N_4547,N_3076,N_3070);
nand U4548 (N_4548,N_3493,N_3527);
nor U4549 (N_4549,N_3043,N_3687);
nand U4550 (N_4550,N_3568,N_3141);
or U4551 (N_4551,N_3972,N_3119);
and U4552 (N_4552,N_3908,N_3184);
nor U4553 (N_4553,N_3504,N_3053);
or U4554 (N_4554,N_3160,N_3201);
nand U4555 (N_4555,N_3501,N_3477);
or U4556 (N_4556,N_3239,N_3904);
nand U4557 (N_4557,N_3931,N_3372);
or U4558 (N_4558,N_3226,N_3953);
and U4559 (N_4559,N_3139,N_3707);
nand U4560 (N_4560,N_3610,N_3973);
and U4561 (N_4561,N_3213,N_3416);
or U4562 (N_4562,N_3308,N_3240);
and U4563 (N_4563,N_3523,N_3920);
nand U4564 (N_4564,N_3402,N_3230);
nand U4565 (N_4565,N_3244,N_3020);
and U4566 (N_4566,N_3867,N_3393);
or U4567 (N_4567,N_3397,N_3731);
and U4568 (N_4568,N_3029,N_3530);
nand U4569 (N_4569,N_3599,N_3649);
nand U4570 (N_4570,N_3812,N_3488);
nor U4571 (N_4571,N_3153,N_3821);
nand U4572 (N_4572,N_3936,N_3781);
or U4573 (N_4573,N_3885,N_3593);
nand U4574 (N_4574,N_3350,N_3117);
nand U4575 (N_4575,N_3631,N_3008);
nor U4576 (N_4576,N_3882,N_3529);
or U4577 (N_4577,N_3076,N_3226);
nor U4578 (N_4578,N_3013,N_3531);
or U4579 (N_4579,N_3772,N_3608);
or U4580 (N_4580,N_3944,N_3979);
and U4581 (N_4581,N_3085,N_3911);
and U4582 (N_4582,N_3580,N_3473);
and U4583 (N_4583,N_3497,N_3710);
nand U4584 (N_4584,N_3884,N_3280);
nand U4585 (N_4585,N_3912,N_3300);
or U4586 (N_4586,N_3766,N_3957);
or U4587 (N_4587,N_3340,N_3189);
or U4588 (N_4588,N_3634,N_3164);
or U4589 (N_4589,N_3642,N_3074);
nand U4590 (N_4590,N_3633,N_3508);
nand U4591 (N_4591,N_3515,N_3101);
nand U4592 (N_4592,N_3729,N_3905);
and U4593 (N_4593,N_3381,N_3281);
nor U4594 (N_4594,N_3615,N_3018);
or U4595 (N_4595,N_3787,N_3801);
nand U4596 (N_4596,N_3321,N_3825);
and U4597 (N_4597,N_3639,N_3687);
or U4598 (N_4598,N_3732,N_3982);
nor U4599 (N_4599,N_3594,N_3003);
or U4600 (N_4600,N_3898,N_3619);
nand U4601 (N_4601,N_3898,N_3559);
nand U4602 (N_4602,N_3888,N_3381);
or U4603 (N_4603,N_3093,N_3954);
nor U4604 (N_4604,N_3507,N_3054);
and U4605 (N_4605,N_3972,N_3530);
nor U4606 (N_4606,N_3940,N_3594);
and U4607 (N_4607,N_3238,N_3339);
nand U4608 (N_4608,N_3219,N_3638);
and U4609 (N_4609,N_3087,N_3727);
nand U4610 (N_4610,N_3389,N_3380);
or U4611 (N_4611,N_3384,N_3293);
or U4612 (N_4612,N_3542,N_3849);
nand U4613 (N_4613,N_3994,N_3677);
nor U4614 (N_4614,N_3532,N_3429);
nand U4615 (N_4615,N_3027,N_3910);
or U4616 (N_4616,N_3553,N_3819);
and U4617 (N_4617,N_3106,N_3248);
nand U4618 (N_4618,N_3097,N_3871);
nand U4619 (N_4619,N_3396,N_3453);
and U4620 (N_4620,N_3696,N_3804);
and U4621 (N_4621,N_3642,N_3567);
nor U4622 (N_4622,N_3382,N_3897);
nand U4623 (N_4623,N_3397,N_3753);
or U4624 (N_4624,N_3943,N_3781);
or U4625 (N_4625,N_3774,N_3377);
or U4626 (N_4626,N_3100,N_3243);
nand U4627 (N_4627,N_3972,N_3582);
nor U4628 (N_4628,N_3629,N_3306);
and U4629 (N_4629,N_3472,N_3706);
nor U4630 (N_4630,N_3850,N_3675);
nand U4631 (N_4631,N_3064,N_3522);
or U4632 (N_4632,N_3155,N_3446);
or U4633 (N_4633,N_3628,N_3341);
and U4634 (N_4634,N_3826,N_3486);
and U4635 (N_4635,N_3681,N_3661);
nor U4636 (N_4636,N_3425,N_3248);
or U4637 (N_4637,N_3327,N_3530);
nand U4638 (N_4638,N_3707,N_3851);
nand U4639 (N_4639,N_3201,N_3838);
or U4640 (N_4640,N_3883,N_3312);
nand U4641 (N_4641,N_3096,N_3115);
nor U4642 (N_4642,N_3898,N_3311);
and U4643 (N_4643,N_3241,N_3473);
nand U4644 (N_4644,N_3816,N_3931);
or U4645 (N_4645,N_3834,N_3513);
nor U4646 (N_4646,N_3194,N_3039);
nor U4647 (N_4647,N_3067,N_3266);
or U4648 (N_4648,N_3247,N_3018);
nand U4649 (N_4649,N_3938,N_3276);
or U4650 (N_4650,N_3046,N_3401);
and U4651 (N_4651,N_3287,N_3810);
or U4652 (N_4652,N_3181,N_3837);
nor U4653 (N_4653,N_3066,N_3274);
or U4654 (N_4654,N_3257,N_3021);
and U4655 (N_4655,N_3855,N_3428);
or U4656 (N_4656,N_3659,N_3887);
nand U4657 (N_4657,N_3448,N_3267);
nand U4658 (N_4658,N_3567,N_3767);
nand U4659 (N_4659,N_3042,N_3020);
nand U4660 (N_4660,N_3080,N_3105);
or U4661 (N_4661,N_3765,N_3509);
or U4662 (N_4662,N_3079,N_3568);
nand U4663 (N_4663,N_3809,N_3285);
nor U4664 (N_4664,N_3044,N_3461);
or U4665 (N_4665,N_3455,N_3746);
nand U4666 (N_4666,N_3771,N_3725);
and U4667 (N_4667,N_3235,N_3748);
or U4668 (N_4668,N_3214,N_3423);
nand U4669 (N_4669,N_3029,N_3898);
nand U4670 (N_4670,N_3568,N_3273);
nand U4671 (N_4671,N_3084,N_3268);
and U4672 (N_4672,N_3798,N_3717);
or U4673 (N_4673,N_3753,N_3565);
nor U4674 (N_4674,N_3901,N_3362);
nand U4675 (N_4675,N_3529,N_3558);
or U4676 (N_4676,N_3563,N_3979);
nor U4677 (N_4677,N_3450,N_3581);
nor U4678 (N_4678,N_3185,N_3268);
nor U4679 (N_4679,N_3127,N_3866);
xor U4680 (N_4680,N_3638,N_3566);
nor U4681 (N_4681,N_3025,N_3367);
nor U4682 (N_4682,N_3906,N_3956);
nand U4683 (N_4683,N_3886,N_3494);
xor U4684 (N_4684,N_3612,N_3202);
nor U4685 (N_4685,N_3230,N_3982);
nor U4686 (N_4686,N_3453,N_3174);
or U4687 (N_4687,N_3652,N_3262);
nand U4688 (N_4688,N_3131,N_3333);
or U4689 (N_4689,N_3033,N_3432);
nor U4690 (N_4690,N_3810,N_3940);
nand U4691 (N_4691,N_3775,N_3779);
and U4692 (N_4692,N_3132,N_3992);
and U4693 (N_4693,N_3969,N_3319);
and U4694 (N_4694,N_3863,N_3724);
nor U4695 (N_4695,N_3634,N_3711);
and U4696 (N_4696,N_3349,N_3094);
and U4697 (N_4697,N_3755,N_3231);
and U4698 (N_4698,N_3656,N_3471);
and U4699 (N_4699,N_3158,N_3875);
nand U4700 (N_4700,N_3820,N_3903);
and U4701 (N_4701,N_3751,N_3900);
nor U4702 (N_4702,N_3657,N_3852);
nand U4703 (N_4703,N_3738,N_3090);
nor U4704 (N_4704,N_3263,N_3147);
nand U4705 (N_4705,N_3353,N_3461);
or U4706 (N_4706,N_3303,N_3000);
nor U4707 (N_4707,N_3639,N_3580);
nor U4708 (N_4708,N_3103,N_3894);
xor U4709 (N_4709,N_3881,N_3562);
nor U4710 (N_4710,N_3519,N_3904);
nand U4711 (N_4711,N_3062,N_3703);
and U4712 (N_4712,N_3906,N_3592);
nand U4713 (N_4713,N_3068,N_3031);
nor U4714 (N_4714,N_3384,N_3719);
or U4715 (N_4715,N_3219,N_3338);
nand U4716 (N_4716,N_3821,N_3089);
nand U4717 (N_4717,N_3551,N_3619);
xor U4718 (N_4718,N_3249,N_3262);
nand U4719 (N_4719,N_3964,N_3965);
and U4720 (N_4720,N_3185,N_3313);
and U4721 (N_4721,N_3935,N_3297);
nand U4722 (N_4722,N_3022,N_3413);
or U4723 (N_4723,N_3953,N_3614);
and U4724 (N_4724,N_3350,N_3627);
nand U4725 (N_4725,N_3242,N_3710);
nand U4726 (N_4726,N_3296,N_3541);
and U4727 (N_4727,N_3926,N_3618);
nand U4728 (N_4728,N_3079,N_3060);
nand U4729 (N_4729,N_3261,N_3709);
or U4730 (N_4730,N_3518,N_3845);
nor U4731 (N_4731,N_3347,N_3950);
and U4732 (N_4732,N_3036,N_3309);
nand U4733 (N_4733,N_3912,N_3858);
and U4734 (N_4734,N_3589,N_3948);
nor U4735 (N_4735,N_3433,N_3458);
nand U4736 (N_4736,N_3729,N_3634);
and U4737 (N_4737,N_3979,N_3968);
nand U4738 (N_4738,N_3586,N_3923);
nor U4739 (N_4739,N_3737,N_3433);
nor U4740 (N_4740,N_3779,N_3653);
and U4741 (N_4741,N_3524,N_3036);
and U4742 (N_4742,N_3607,N_3041);
and U4743 (N_4743,N_3691,N_3841);
nand U4744 (N_4744,N_3778,N_3440);
and U4745 (N_4745,N_3142,N_3005);
nor U4746 (N_4746,N_3074,N_3221);
and U4747 (N_4747,N_3919,N_3628);
or U4748 (N_4748,N_3714,N_3077);
and U4749 (N_4749,N_3012,N_3276);
and U4750 (N_4750,N_3562,N_3086);
or U4751 (N_4751,N_3428,N_3693);
or U4752 (N_4752,N_3817,N_3393);
or U4753 (N_4753,N_3529,N_3241);
or U4754 (N_4754,N_3155,N_3068);
nor U4755 (N_4755,N_3908,N_3696);
or U4756 (N_4756,N_3288,N_3229);
or U4757 (N_4757,N_3402,N_3514);
nand U4758 (N_4758,N_3905,N_3194);
nor U4759 (N_4759,N_3757,N_3358);
or U4760 (N_4760,N_3990,N_3723);
or U4761 (N_4761,N_3416,N_3978);
or U4762 (N_4762,N_3164,N_3563);
and U4763 (N_4763,N_3459,N_3737);
or U4764 (N_4764,N_3320,N_3556);
nor U4765 (N_4765,N_3261,N_3156);
and U4766 (N_4766,N_3188,N_3366);
nor U4767 (N_4767,N_3950,N_3696);
nor U4768 (N_4768,N_3107,N_3436);
or U4769 (N_4769,N_3822,N_3776);
nand U4770 (N_4770,N_3241,N_3851);
and U4771 (N_4771,N_3895,N_3090);
and U4772 (N_4772,N_3756,N_3154);
or U4773 (N_4773,N_3060,N_3763);
nor U4774 (N_4774,N_3225,N_3711);
or U4775 (N_4775,N_3875,N_3939);
nor U4776 (N_4776,N_3153,N_3674);
and U4777 (N_4777,N_3687,N_3420);
nand U4778 (N_4778,N_3839,N_3755);
and U4779 (N_4779,N_3875,N_3615);
nor U4780 (N_4780,N_3691,N_3257);
or U4781 (N_4781,N_3087,N_3775);
nand U4782 (N_4782,N_3444,N_3755);
xor U4783 (N_4783,N_3812,N_3574);
nand U4784 (N_4784,N_3967,N_3051);
nor U4785 (N_4785,N_3901,N_3892);
and U4786 (N_4786,N_3427,N_3231);
or U4787 (N_4787,N_3721,N_3984);
nand U4788 (N_4788,N_3391,N_3855);
nor U4789 (N_4789,N_3036,N_3567);
or U4790 (N_4790,N_3429,N_3457);
or U4791 (N_4791,N_3184,N_3031);
or U4792 (N_4792,N_3391,N_3950);
nor U4793 (N_4793,N_3613,N_3544);
or U4794 (N_4794,N_3037,N_3838);
and U4795 (N_4795,N_3610,N_3486);
nand U4796 (N_4796,N_3357,N_3738);
and U4797 (N_4797,N_3416,N_3843);
or U4798 (N_4798,N_3725,N_3012);
nor U4799 (N_4799,N_3427,N_3633);
nor U4800 (N_4800,N_3216,N_3079);
nand U4801 (N_4801,N_3401,N_3174);
and U4802 (N_4802,N_3384,N_3506);
and U4803 (N_4803,N_3716,N_3482);
nand U4804 (N_4804,N_3347,N_3779);
or U4805 (N_4805,N_3798,N_3637);
xnor U4806 (N_4806,N_3234,N_3575);
nor U4807 (N_4807,N_3892,N_3418);
or U4808 (N_4808,N_3359,N_3154);
or U4809 (N_4809,N_3824,N_3762);
nor U4810 (N_4810,N_3918,N_3984);
nor U4811 (N_4811,N_3991,N_3986);
or U4812 (N_4812,N_3917,N_3464);
nand U4813 (N_4813,N_3984,N_3516);
nor U4814 (N_4814,N_3185,N_3941);
and U4815 (N_4815,N_3300,N_3124);
and U4816 (N_4816,N_3426,N_3371);
nand U4817 (N_4817,N_3318,N_3806);
nor U4818 (N_4818,N_3960,N_3248);
nor U4819 (N_4819,N_3529,N_3174);
or U4820 (N_4820,N_3439,N_3994);
nand U4821 (N_4821,N_3744,N_3338);
or U4822 (N_4822,N_3753,N_3598);
nand U4823 (N_4823,N_3592,N_3176);
and U4824 (N_4824,N_3505,N_3378);
and U4825 (N_4825,N_3875,N_3853);
or U4826 (N_4826,N_3128,N_3923);
nand U4827 (N_4827,N_3058,N_3010);
nor U4828 (N_4828,N_3644,N_3858);
and U4829 (N_4829,N_3362,N_3280);
nor U4830 (N_4830,N_3033,N_3749);
and U4831 (N_4831,N_3364,N_3497);
nor U4832 (N_4832,N_3549,N_3331);
and U4833 (N_4833,N_3284,N_3359);
nand U4834 (N_4834,N_3203,N_3406);
and U4835 (N_4835,N_3541,N_3929);
or U4836 (N_4836,N_3387,N_3476);
nand U4837 (N_4837,N_3298,N_3686);
and U4838 (N_4838,N_3342,N_3152);
and U4839 (N_4839,N_3706,N_3905);
nor U4840 (N_4840,N_3764,N_3438);
nand U4841 (N_4841,N_3441,N_3769);
and U4842 (N_4842,N_3110,N_3262);
nor U4843 (N_4843,N_3567,N_3323);
nor U4844 (N_4844,N_3023,N_3249);
nor U4845 (N_4845,N_3282,N_3999);
nand U4846 (N_4846,N_3988,N_3859);
or U4847 (N_4847,N_3310,N_3182);
nand U4848 (N_4848,N_3343,N_3275);
nor U4849 (N_4849,N_3688,N_3863);
nand U4850 (N_4850,N_3109,N_3358);
nand U4851 (N_4851,N_3678,N_3427);
and U4852 (N_4852,N_3909,N_3389);
nor U4853 (N_4853,N_3092,N_3734);
nand U4854 (N_4854,N_3725,N_3222);
nor U4855 (N_4855,N_3522,N_3619);
and U4856 (N_4856,N_3984,N_3233);
nor U4857 (N_4857,N_3591,N_3773);
nor U4858 (N_4858,N_3505,N_3764);
nand U4859 (N_4859,N_3213,N_3399);
nor U4860 (N_4860,N_3691,N_3021);
and U4861 (N_4861,N_3846,N_3185);
and U4862 (N_4862,N_3848,N_3860);
nor U4863 (N_4863,N_3882,N_3287);
and U4864 (N_4864,N_3924,N_3795);
and U4865 (N_4865,N_3690,N_3149);
and U4866 (N_4866,N_3874,N_3200);
nor U4867 (N_4867,N_3261,N_3734);
nand U4868 (N_4868,N_3538,N_3230);
and U4869 (N_4869,N_3744,N_3153);
or U4870 (N_4870,N_3958,N_3362);
or U4871 (N_4871,N_3824,N_3766);
or U4872 (N_4872,N_3806,N_3046);
or U4873 (N_4873,N_3705,N_3020);
nand U4874 (N_4874,N_3831,N_3476);
nand U4875 (N_4875,N_3740,N_3849);
and U4876 (N_4876,N_3572,N_3563);
or U4877 (N_4877,N_3106,N_3902);
and U4878 (N_4878,N_3705,N_3472);
nand U4879 (N_4879,N_3201,N_3600);
or U4880 (N_4880,N_3355,N_3287);
nand U4881 (N_4881,N_3827,N_3394);
and U4882 (N_4882,N_3849,N_3167);
or U4883 (N_4883,N_3550,N_3064);
nor U4884 (N_4884,N_3922,N_3908);
nand U4885 (N_4885,N_3041,N_3770);
and U4886 (N_4886,N_3750,N_3295);
xor U4887 (N_4887,N_3678,N_3699);
nor U4888 (N_4888,N_3325,N_3908);
nor U4889 (N_4889,N_3889,N_3426);
and U4890 (N_4890,N_3845,N_3540);
and U4891 (N_4891,N_3948,N_3168);
and U4892 (N_4892,N_3924,N_3532);
and U4893 (N_4893,N_3924,N_3266);
or U4894 (N_4894,N_3480,N_3390);
nor U4895 (N_4895,N_3495,N_3735);
or U4896 (N_4896,N_3716,N_3383);
or U4897 (N_4897,N_3070,N_3685);
or U4898 (N_4898,N_3770,N_3579);
nand U4899 (N_4899,N_3066,N_3519);
and U4900 (N_4900,N_3777,N_3146);
or U4901 (N_4901,N_3712,N_3868);
nor U4902 (N_4902,N_3463,N_3097);
and U4903 (N_4903,N_3909,N_3840);
and U4904 (N_4904,N_3024,N_3632);
or U4905 (N_4905,N_3583,N_3337);
or U4906 (N_4906,N_3789,N_3141);
nor U4907 (N_4907,N_3396,N_3448);
nand U4908 (N_4908,N_3547,N_3430);
and U4909 (N_4909,N_3404,N_3410);
or U4910 (N_4910,N_3366,N_3666);
nand U4911 (N_4911,N_3811,N_3483);
and U4912 (N_4912,N_3263,N_3397);
nand U4913 (N_4913,N_3634,N_3878);
and U4914 (N_4914,N_3641,N_3244);
nand U4915 (N_4915,N_3417,N_3376);
and U4916 (N_4916,N_3591,N_3370);
nor U4917 (N_4917,N_3834,N_3489);
nand U4918 (N_4918,N_3301,N_3357);
nor U4919 (N_4919,N_3641,N_3242);
nor U4920 (N_4920,N_3783,N_3102);
or U4921 (N_4921,N_3716,N_3897);
and U4922 (N_4922,N_3957,N_3720);
nor U4923 (N_4923,N_3939,N_3142);
nand U4924 (N_4924,N_3814,N_3702);
and U4925 (N_4925,N_3033,N_3579);
nor U4926 (N_4926,N_3163,N_3301);
nor U4927 (N_4927,N_3744,N_3756);
and U4928 (N_4928,N_3791,N_3193);
nand U4929 (N_4929,N_3484,N_3794);
nor U4930 (N_4930,N_3841,N_3129);
xnor U4931 (N_4931,N_3064,N_3030);
or U4932 (N_4932,N_3096,N_3309);
or U4933 (N_4933,N_3458,N_3183);
nor U4934 (N_4934,N_3977,N_3647);
nand U4935 (N_4935,N_3547,N_3870);
and U4936 (N_4936,N_3710,N_3441);
nor U4937 (N_4937,N_3130,N_3345);
and U4938 (N_4938,N_3433,N_3995);
nor U4939 (N_4939,N_3820,N_3881);
xnor U4940 (N_4940,N_3122,N_3687);
nor U4941 (N_4941,N_3762,N_3775);
xnor U4942 (N_4942,N_3897,N_3822);
and U4943 (N_4943,N_3832,N_3097);
and U4944 (N_4944,N_3231,N_3129);
nand U4945 (N_4945,N_3414,N_3886);
and U4946 (N_4946,N_3316,N_3253);
nand U4947 (N_4947,N_3917,N_3551);
nor U4948 (N_4948,N_3549,N_3846);
nand U4949 (N_4949,N_3593,N_3610);
nor U4950 (N_4950,N_3505,N_3590);
nand U4951 (N_4951,N_3709,N_3252);
or U4952 (N_4952,N_3111,N_3818);
nor U4953 (N_4953,N_3268,N_3805);
or U4954 (N_4954,N_3895,N_3998);
nor U4955 (N_4955,N_3347,N_3432);
or U4956 (N_4956,N_3921,N_3716);
or U4957 (N_4957,N_3961,N_3728);
nand U4958 (N_4958,N_3723,N_3805);
or U4959 (N_4959,N_3958,N_3062);
nand U4960 (N_4960,N_3161,N_3370);
xnor U4961 (N_4961,N_3425,N_3016);
nor U4962 (N_4962,N_3867,N_3723);
nand U4963 (N_4963,N_3362,N_3738);
and U4964 (N_4964,N_3498,N_3436);
nor U4965 (N_4965,N_3429,N_3275);
nor U4966 (N_4966,N_3728,N_3981);
and U4967 (N_4967,N_3634,N_3691);
or U4968 (N_4968,N_3780,N_3655);
nand U4969 (N_4969,N_3545,N_3065);
and U4970 (N_4970,N_3853,N_3095);
nor U4971 (N_4971,N_3475,N_3776);
nand U4972 (N_4972,N_3599,N_3767);
and U4973 (N_4973,N_3162,N_3294);
and U4974 (N_4974,N_3626,N_3048);
and U4975 (N_4975,N_3280,N_3380);
nor U4976 (N_4976,N_3983,N_3998);
and U4977 (N_4977,N_3423,N_3487);
or U4978 (N_4978,N_3279,N_3528);
and U4979 (N_4979,N_3359,N_3845);
nand U4980 (N_4980,N_3554,N_3987);
or U4981 (N_4981,N_3307,N_3100);
or U4982 (N_4982,N_3090,N_3186);
nor U4983 (N_4983,N_3628,N_3552);
nor U4984 (N_4984,N_3531,N_3309);
and U4985 (N_4985,N_3738,N_3463);
and U4986 (N_4986,N_3279,N_3091);
nand U4987 (N_4987,N_3147,N_3629);
and U4988 (N_4988,N_3805,N_3816);
nor U4989 (N_4989,N_3205,N_3085);
and U4990 (N_4990,N_3649,N_3446);
or U4991 (N_4991,N_3615,N_3845);
nor U4992 (N_4992,N_3801,N_3536);
or U4993 (N_4993,N_3603,N_3906);
nor U4994 (N_4994,N_3224,N_3400);
nor U4995 (N_4995,N_3729,N_3077);
nand U4996 (N_4996,N_3065,N_3955);
or U4997 (N_4997,N_3227,N_3241);
nor U4998 (N_4998,N_3011,N_3395);
nor U4999 (N_4999,N_3279,N_3052);
nand U5000 (N_5000,N_4389,N_4331);
nand U5001 (N_5001,N_4538,N_4722);
and U5002 (N_5002,N_4823,N_4440);
nor U5003 (N_5003,N_4866,N_4103);
nand U5004 (N_5004,N_4643,N_4934);
or U5005 (N_5005,N_4749,N_4995);
and U5006 (N_5006,N_4859,N_4757);
and U5007 (N_5007,N_4210,N_4009);
nand U5008 (N_5008,N_4144,N_4745);
nand U5009 (N_5009,N_4892,N_4076);
nand U5010 (N_5010,N_4896,N_4290);
nor U5011 (N_5011,N_4758,N_4195);
nor U5012 (N_5012,N_4016,N_4809);
and U5013 (N_5013,N_4512,N_4420);
or U5014 (N_5014,N_4003,N_4747);
nand U5015 (N_5015,N_4278,N_4048);
or U5016 (N_5016,N_4034,N_4721);
and U5017 (N_5017,N_4352,N_4376);
nor U5018 (N_5018,N_4573,N_4702);
nand U5019 (N_5019,N_4148,N_4391);
or U5020 (N_5020,N_4614,N_4097);
and U5021 (N_5021,N_4407,N_4057);
and U5022 (N_5022,N_4616,N_4431);
and U5023 (N_5023,N_4160,N_4728);
nand U5024 (N_5024,N_4313,N_4200);
nor U5025 (N_5025,N_4143,N_4150);
or U5026 (N_5026,N_4243,N_4631);
nand U5027 (N_5027,N_4387,N_4026);
or U5028 (N_5028,N_4489,N_4190);
or U5029 (N_5029,N_4186,N_4116);
or U5030 (N_5030,N_4484,N_4342);
or U5031 (N_5031,N_4580,N_4030);
or U5032 (N_5032,N_4045,N_4867);
or U5033 (N_5033,N_4427,N_4818);
or U5034 (N_5034,N_4215,N_4838);
nand U5035 (N_5035,N_4385,N_4474);
nand U5036 (N_5036,N_4106,N_4002);
nor U5037 (N_5037,N_4032,N_4693);
nor U5038 (N_5038,N_4274,N_4323);
or U5039 (N_5039,N_4732,N_4434);
nor U5040 (N_5040,N_4320,N_4343);
nor U5041 (N_5041,N_4304,N_4824);
nor U5042 (N_5042,N_4107,N_4104);
or U5043 (N_5043,N_4166,N_4406);
and U5044 (N_5044,N_4065,N_4714);
and U5045 (N_5045,N_4888,N_4607);
or U5046 (N_5046,N_4084,N_4379);
nand U5047 (N_5047,N_4390,N_4445);
nor U5048 (N_5048,N_4428,N_4677);
nand U5049 (N_5049,N_4766,N_4925);
nor U5050 (N_5050,N_4014,N_4956);
and U5051 (N_5051,N_4327,N_4531);
nor U5052 (N_5052,N_4910,N_4754);
nand U5053 (N_5053,N_4444,N_4609);
or U5054 (N_5054,N_4613,N_4211);
nor U5055 (N_5055,N_4558,N_4288);
and U5056 (N_5056,N_4337,N_4124);
and U5057 (N_5057,N_4687,N_4546);
or U5058 (N_5058,N_4247,N_4472);
nand U5059 (N_5059,N_4040,N_4822);
and U5060 (N_5060,N_4173,N_4506);
nor U5061 (N_5061,N_4088,N_4534);
nand U5062 (N_5062,N_4830,N_4435);
or U5063 (N_5063,N_4375,N_4196);
or U5064 (N_5064,N_4547,N_4673);
and U5065 (N_5065,N_4311,N_4096);
nor U5066 (N_5066,N_4101,N_4697);
or U5067 (N_5067,N_4436,N_4539);
or U5068 (N_5068,N_4115,N_4933);
and U5069 (N_5069,N_4516,N_4615);
nor U5070 (N_5070,N_4363,N_4183);
or U5071 (N_5071,N_4479,N_4711);
or U5072 (N_5072,N_4502,N_4552);
or U5073 (N_5073,N_4370,N_4276);
or U5074 (N_5074,N_4907,N_4949);
and U5075 (N_5075,N_4495,N_4662);
nor U5076 (N_5076,N_4665,N_4362);
or U5077 (N_5077,N_4204,N_4081);
nand U5078 (N_5078,N_4828,N_4307);
and U5079 (N_5079,N_4620,N_4346);
and U5080 (N_5080,N_4131,N_4037);
and U5081 (N_5081,N_4686,N_4819);
and U5082 (N_5082,N_4821,N_4356);
nor U5083 (N_5083,N_4238,N_4837);
or U5084 (N_5084,N_4466,N_4943);
nand U5085 (N_5085,N_4227,N_4622);
nand U5086 (N_5086,N_4475,N_4685);
nand U5087 (N_5087,N_4449,N_4645);
or U5088 (N_5088,N_4796,N_4799);
or U5089 (N_5089,N_4091,N_4465);
or U5090 (N_5090,N_4717,N_4256);
nand U5091 (N_5091,N_4606,N_4325);
and U5092 (N_5092,N_4078,N_4712);
nor U5093 (N_5093,N_4043,N_4634);
nand U5094 (N_5094,N_4865,N_4366);
nand U5095 (N_5095,N_4197,N_4660);
nor U5096 (N_5096,N_4595,N_4666);
and U5097 (N_5097,N_4765,N_4062);
nand U5098 (N_5098,N_4726,N_4521);
or U5099 (N_5099,N_4561,N_4382);
nand U5100 (N_5100,N_4785,N_4813);
and U5101 (N_5101,N_4291,N_4586);
nor U5102 (N_5102,N_4938,N_4271);
and U5103 (N_5103,N_4090,N_4610);
or U5104 (N_5104,N_4075,N_4018);
nor U5105 (N_5105,N_4840,N_4638);
nand U5106 (N_5106,N_4921,N_4007);
nor U5107 (N_5107,N_4171,N_4876);
and U5108 (N_5108,N_4364,N_4680);
nand U5109 (N_5109,N_4013,N_4345);
and U5110 (N_5110,N_4470,N_4410);
nor U5111 (N_5111,N_4740,N_4229);
nand U5112 (N_5112,N_4053,N_4292);
nor U5113 (N_5113,N_4651,N_4361);
nand U5114 (N_5114,N_4804,N_4523);
or U5115 (N_5115,N_4825,N_4085);
xnor U5116 (N_5116,N_4155,N_4133);
nor U5117 (N_5117,N_4977,N_4532);
nor U5118 (N_5118,N_4808,N_4898);
and U5119 (N_5119,N_4241,N_4263);
nor U5120 (N_5120,N_4224,N_4504);
nor U5121 (N_5121,N_4460,N_4682);
or U5122 (N_5122,N_4033,N_4626);
and U5123 (N_5123,N_4782,N_4378);
or U5124 (N_5124,N_4242,N_4476);
and U5125 (N_5125,N_4168,N_4891);
and U5126 (N_5126,N_4773,N_4761);
nand U5127 (N_5127,N_4403,N_4841);
nand U5128 (N_5128,N_4494,N_4272);
or U5129 (N_5129,N_4082,N_4394);
and U5130 (N_5130,N_4914,N_4635);
nand U5131 (N_5131,N_4142,N_4365);
or U5132 (N_5132,N_4676,N_4718);
or U5133 (N_5133,N_4857,N_4354);
nor U5134 (N_5134,N_4054,N_4095);
or U5135 (N_5135,N_4854,N_4960);
nor U5136 (N_5136,N_4303,N_4768);
or U5137 (N_5137,N_4039,N_4945);
or U5138 (N_5138,N_4158,N_4480);
nand U5139 (N_5139,N_4679,N_4911);
or U5140 (N_5140,N_4151,N_4264);
nor U5141 (N_5141,N_4163,N_4912);
nand U5142 (N_5142,N_4762,N_4529);
or U5143 (N_5143,N_4126,N_4985);
or U5144 (N_5144,N_4301,N_4525);
nor U5145 (N_5145,N_4441,N_4738);
or U5146 (N_5146,N_4519,N_4652);
nand U5147 (N_5147,N_4931,N_4844);
and U5148 (N_5148,N_4087,N_4948);
or U5149 (N_5149,N_4257,N_4770);
nand U5150 (N_5150,N_4778,N_4261);
nand U5151 (N_5151,N_4100,N_4618);
nand U5152 (N_5152,N_4500,N_4259);
and U5153 (N_5153,N_4456,N_4672);
nor U5154 (N_5154,N_4791,N_4862);
nor U5155 (N_5155,N_4737,N_4513);
nor U5156 (N_5156,N_4417,N_4755);
nand U5157 (N_5157,N_4418,N_4027);
or U5158 (N_5158,N_4232,N_4649);
nor U5159 (N_5159,N_4395,N_4599);
nor U5160 (N_5160,N_4946,N_4498);
or U5161 (N_5161,N_4217,N_4357);
or U5162 (N_5162,N_4083,N_4192);
and U5163 (N_5163,N_4569,N_4992);
nor U5164 (N_5164,N_4180,N_4262);
and U5165 (N_5165,N_4909,N_4764);
nor U5166 (N_5166,N_4706,N_4939);
nor U5167 (N_5167,N_4942,N_4899);
or U5168 (N_5168,N_4459,N_4974);
nor U5169 (N_5169,N_4134,N_4863);
nor U5170 (N_5170,N_4073,N_4284);
and U5171 (N_5171,N_4986,N_4450);
or U5172 (N_5172,N_4371,N_4641);
nand U5173 (N_5173,N_4553,N_4172);
and U5174 (N_5174,N_4965,N_4113);
or U5175 (N_5175,N_4293,N_4596);
and U5176 (N_5176,N_4806,N_4267);
nor U5177 (N_5177,N_4887,N_4727);
nor U5178 (N_5178,N_4077,N_4692);
nand U5179 (N_5179,N_4924,N_4298);
nand U5180 (N_5180,N_4185,N_4833);
nor U5181 (N_5181,N_4976,N_4001);
and U5182 (N_5182,N_4266,N_4636);
and U5183 (N_5183,N_4571,N_4355);
or U5184 (N_5184,N_4683,N_4954);
nor U5185 (N_5185,N_4415,N_4878);
or U5186 (N_5186,N_4856,N_4592);
or U5187 (N_5187,N_4971,N_4492);
nand U5188 (N_5188,N_4182,N_4701);
and U5189 (N_5189,N_4581,N_4324);
nand U5190 (N_5190,N_4165,N_4880);
nor U5191 (N_5191,N_4556,N_4404);
nor U5192 (N_5192,N_4218,N_4326);
or U5193 (N_5193,N_4152,N_4296);
nand U5194 (N_5194,N_4287,N_4109);
or U5195 (N_5195,N_4852,N_4674);
or U5196 (N_5196,N_4594,N_4501);
and U5197 (N_5197,N_4932,N_4125);
nor U5198 (N_5198,N_4208,N_4756);
nand U5199 (N_5199,N_4829,N_4559);
nand U5200 (N_5200,N_4792,N_4164);
nor U5201 (N_5201,N_4663,N_4255);
or U5202 (N_5202,N_4386,N_4038);
nand U5203 (N_5203,N_4842,N_4917);
and U5204 (N_5204,N_4332,N_4093);
nor U5205 (N_5205,N_4451,N_4246);
and U5206 (N_5206,N_4877,N_4020);
or U5207 (N_5207,N_4112,N_4889);
nor U5208 (N_5208,N_4251,N_4120);
and U5209 (N_5209,N_4383,N_4279);
or U5210 (N_5210,N_4544,N_4514);
and U5211 (N_5211,N_4280,N_4029);
nor U5212 (N_5212,N_4788,N_4881);
or U5213 (N_5213,N_4870,N_4780);
nor U5214 (N_5214,N_4826,N_4079);
or U5215 (N_5215,N_4815,N_4597);
nand U5216 (N_5216,N_4589,N_4294);
nor U5217 (N_5217,N_4055,N_4381);
or U5218 (N_5218,N_4414,N_4194);
nor U5219 (N_5219,N_4805,N_4608);
or U5220 (N_5220,N_4950,N_4963);
or U5221 (N_5221,N_4537,N_4213);
nor U5222 (N_5222,N_4729,N_4012);
and U5223 (N_5223,N_4187,N_4179);
nand U5224 (N_5224,N_4214,N_4604);
or U5225 (N_5225,N_4836,N_4372);
nor U5226 (N_5226,N_4004,N_4353);
nor U5227 (N_5227,N_4904,N_4930);
nand U5228 (N_5228,N_4019,N_4318);
and U5229 (N_5229,N_4795,N_4817);
and U5230 (N_5230,N_4540,N_4154);
or U5231 (N_5231,N_4700,N_4511);
or U5232 (N_5232,N_4035,N_4858);
nor U5233 (N_5233,N_4868,N_4050);
and U5234 (N_5234,N_4999,N_4188);
nand U5235 (N_5235,N_4563,N_4072);
nand U5236 (N_5236,N_4042,N_4225);
or U5237 (N_5237,N_4774,N_4820);
and U5238 (N_5238,N_4181,N_4067);
and U5239 (N_5239,N_4136,N_4111);
nand U5240 (N_5240,N_4835,N_4433);
nor U5241 (N_5241,N_4300,N_4222);
nor U5242 (N_5242,N_4170,N_4250);
nand U5243 (N_5243,N_4810,N_4918);
nand U5244 (N_5244,N_4309,N_4753);
nand U5245 (N_5245,N_4786,N_4966);
or U5246 (N_5246,N_4659,N_4882);
or U5247 (N_5247,N_4691,N_4630);
nand U5248 (N_5248,N_4982,N_4270);
nand U5249 (N_5249,N_4527,N_4282);
nor U5250 (N_5250,N_4099,N_4056);
and U5251 (N_5251,N_4510,N_4330);
or U5252 (N_5252,N_4477,N_4123);
nor U5253 (N_5253,N_4647,N_4374);
and U5254 (N_5254,N_4191,N_4231);
nand U5255 (N_5255,N_4623,N_4807);
nor U5256 (N_5256,N_4396,N_4600);
nand U5257 (N_5257,N_4936,N_4890);
nand U5258 (N_5258,N_4781,N_4446);
and U5259 (N_5259,N_4074,N_4258);
nor U5260 (N_5260,N_4011,N_4743);
nand U5261 (N_5261,N_4421,N_4426);
nor U5262 (N_5262,N_4989,N_4046);
nand U5263 (N_5263,N_4260,N_4716);
nand U5264 (N_5264,N_4855,N_4802);
and U5265 (N_5265,N_4399,N_4159);
nor U5266 (N_5266,N_4310,N_4316);
nand U5267 (N_5267,N_4703,N_4025);
nor U5268 (N_5268,N_4582,N_4958);
nand U5269 (N_5269,N_4505,N_4707);
or U5270 (N_5270,N_4555,N_4696);
nor U5271 (N_5271,N_4071,N_4688);
and U5272 (N_5272,N_4234,N_4803);
or U5273 (N_5273,N_4927,N_4336);
nor U5274 (N_5274,N_4603,N_4681);
and U5275 (N_5275,N_4627,N_4709);
nor U5276 (N_5276,N_4520,N_4277);
or U5277 (N_5277,N_4964,N_4219);
or U5278 (N_5278,N_4708,N_4664);
nor U5279 (N_5279,N_4129,N_4605);
or U5280 (N_5280,N_4454,N_4734);
and U5281 (N_5281,N_4739,N_4657);
nand U5282 (N_5282,N_4130,N_4347);
nand U5283 (N_5283,N_4831,N_4548);
or U5284 (N_5284,N_4928,N_4968);
or U5285 (N_5285,N_4488,N_4061);
nand U5286 (N_5286,N_4102,N_4973);
nand U5287 (N_5287,N_4733,N_4886);
and U5288 (N_5288,N_4199,N_4457);
nand U5289 (N_5289,N_4189,N_4670);
and U5290 (N_5290,N_4463,N_4509);
and U5291 (N_5291,N_4860,N_4397);
nor U5292 (N_5292,N_4926,N_4408);
and U5293 (N_5293,N_4535,N_4658);
nand U5294 (N_5294,N_4351,N_4157);
or U5295 (N_5295,N_4269,N_4873);
nor U5296 (N_5296,N_4962,N_4167);
nor U5297 (N_5297,N_4128,N_4047);
and U5298 (N_5298,N_4064,N_4602);
or U5299 (N_5299,N_4223,N_4086);
or U5300 (N_5300,N_4874,N_4530);
or U5301 (N_5301,N_4028,N_4006);
nor U5302 (N_5302,N_4156,N_4314);
or U5303 (N_5303,N_4405,N_4240);
nand U5304 (N_5304,N_4834,N_4750);
nor U5305 (N_5305,N_4730,N_4575);
or U5306 (N_5306,N_4419,N_4467);
and U5307 (N_5307,N_4845,N_4360);
nor U5308 (N_5308,N_4646,N_4883);
nand U5309 (N_5309,N_4998,N_4338);
nand U5310 (N_5310,N_4335,N_4895);
nor U5311 (N_5311,N_4482,N_4975);
and U5312 (N_5312,N_4132,N_4060);
nand U5313 (N_5313,N_4341,N_4230);
or U5314 (N_5314,N_4632,N_4800);
nand U5315 (N_5315,N_4759,N_4972);
nor U5316 (N_5316,N_4894,N_4411);
or U5317 (N_5317,N_4127,N_4448);
nand U5318 (N_5318,N_4935,N_4846);
nor U5319 (N_5319,N_4432,N_4049);
or U5320 (N_5320,N_4611,N_4579);
nor U5321 (N_5321,N_4790,N_4369);
nor U5322 (N_5322,N_4562,N_4145);
and U5323 (N_5323,N_4748,N_4497);
nand U5324 (N_5324,N_4121,N_4508);
nand U5325 (N_5325,N_4207,N_4254);
or U5326 (N_5326,N_4902,N_4098);
and U5327 (N_5327,N_4578,N_4731);
or U5328 (N_5328,N_4485,N_4221);
or U5329 (N_5329,N_4216,N_4550);
nor U5330 (N_5330,N_4705,N_4625);
and U5331 (N_5331,N_4654,N_4528);
nand U5332 (N_5332,N_4741,N_4884);
nand U5333 (N_5333,N_4416,N_4010);
nor U5334 (N_5334,N_4572,N_4587);
and U5335 (N_5335,N_4349,N_4900);
or U5336 (N_5336,N_4358,N_4853);
or U5337 (N_5337,N_4851,N_4031);
nor U5338 (N_5338,N_4135,N_4312);
and U5339 (N_5339,N_4794,N_4667);
nor U5340 (N_5340,N_4486,N_4639);
nor U5341 (N_5341,N_4239,N_4308);
and U5342 (N_5342,N_4812,N_4468);
nand U5343 (N_5343,N_4490,N_4661);
or U5344 (N_5344,N_4235,N_4328);
and U5345 (N_5345,N_4483,N_4493);
or U5346 (N_5346,N_4265,N_4644);
or U5347 (N_5347,N_4574,N_4137);
nand U5348 (N_5348,N_4464,N_4499);
and U5349 (N_5349,N_4089,N_4036);
nand U5350 (N_5350,N_4793,N_4801);
or U5351 (N_5351,N_4299,N_4205);
or U5352 (N_5352,N_4704,N_4393);
and U5353 (N_5353,N_4913,N_4952);
and U5354 (N_5354,N_4699,N_4922);
nor U5355 (N_5355,N_4458,N_4777);
xor U5356 (N_5356,N_4720,N_4481);
and U5357 (N_5357,N_4984,N_4253);
nand U5358 (N_5358,N_4916,N_4567);
nand U5359 (N_5359,N_4901,N_4744);
or U5360 (N_5360,N_4690,N_4425);
and U5361 (N_5361,N_4348,N_4769);
or U5362 (N_5362,N_4684,N_4906);
nand U5363 (N_5363,N_4669,N_4487);
nand U5364 (N_5364,N_4775,N_4024);
or U5365 (N_5365,N_4437,N_4576);
nor U5366 (N_5366,N_4543,N_4044);
nor U5367 (N_5367,N_4161,N_4118);
nor U5368 (N_5368,N_4957,N_4245);
nor U5369 (N_5369,N_4967,N_4951);
and U5370 (N_5370,N_4503,N_4590);
and U5371 (N_5371,N_4248,N_4478);
or U5372 (N_5372,N_4373,N_4080);
nor U5373 (N_5373,N_4612,N_4429);
nor U5374 (N_5374,N_4066,N_4893);
nand U5375 (N_5375,N_4117,N_4092);
or U5376 (N_5376,N_4438,N_4713);
nor U5377 (N_5377,N_4455,N_4798);
nand U5378 (N_5378,N_4058,N_4496);
nor U5379 (N_5379,N_4864,N_4203);
nor U5380 (N_5380,N_4285,N_4996);
nand U5381 (N_5381,N_4771,N_4306);
or U5382 (N_5382,N_4175,N_4252);
and U5383 (N_5383,N_4069,N_4811);
or U5384 (N_5384,N_4052,N_4637);
nand U5385 (N_5385,N_4319,N_4668);
nand U5386 (N_5386,N_4871,N_4719);
or U5387 (N_5387,N_4153,N_4671);
and U5388 (N_5388,N_4797,N_4507);
nand U5389 (N_5389,N_4138,N_4551);
nand U5390 (N_5390,N_4752,N_4678);
and U5391 (N_5391,N_4443,N_4322);
nand U5392 (N_5392,N_4850,N_4461);
nor U5393 (N_5393,N_4923,N_4970);
or U5394 (N_5394,N_4198,N_4377);
nand U5395 (N_5395,N_4452,N_4491);
nand U5396 (N_5396,N_4340,N_4517);
nor U5397 (N_5397,N_4212,N_4776);
nor U5398 (N_5398,N_4545,N_4839);
nand U5399 (N_5399,N_4367,N_4929);
nor U5400 (N_5400,N_4695,N_4228);
nor U5401 (N_5401,N_4409,N_4430);
or U5402 (N_5402,N_4725,N_4903);
or U5403 (N_5403,N_4593,N_4783);
nand U5404 (N_5404,N_4640,N_4698);
and U5405 (N_5405,N_4233,N_4542);
or U5406 (N_5406,N_4619,N_4380);
nor U5407 (N_5407,N_4848,N_4827);
nand U5408 (N_5408,N_4447,N_4843);
and U5409 (N_5409,N_4779,N_4515);
and U5410 (N_5410,N_4629,N_4110);
nor U5411 (N_5411,N_4981,N_4384);
xor U5412 (N_5412,N_4915,N_4329);
nand U5413 (N_5413,N_4518,N_4206);
or U5414 (N_5414,N_4584,N_4140);
or U5415 (N_5415,N_4940,N_4177);
and U5416 (N_5416,N_4070,N_4969);
nand U5417 (N_5417,N_4295,N_4473);
nor U5418 (N_5418,N_4273,N_4286);
and U5419 (N_5419,N_4400,N_4368);
nand U5420 (N_5420,N_4655,N_4005);
and U5421 (N_5421,N_4522,N_4988);
nor U5422 (N_5422,N_4000,N_4315);
and U5423 (N_5423,N_4565,N_4959);
nor U5424 (N_5424,N_4178,N_4114);
nor U5425 (N_5425,N_4524,N_4226);
nor U5426 (N_5426,N_4816,N_4202);
nor U5427 (N_5427,N_4146,N_4119);
nand U5428 (N_5428,N_4401,N_4767);
nor U5429 (N_5429,N_4869,N_4236);
nand U5430 (N_5430,N_4947,N_4334);
nand U5431 (N_5431,N_4875,N_4621);
or U5432 (N_5432,N_4469,N_4022);
nor U5433 (N_5433,N_4321,N_4536);
nor U5434 (N_5434,N_4162,N_4879);
nor U5435 (N_5435,N_4861,N_4149);
and U5436 (N_5436,N_4289,N_4169);
nand U5437 (N_5437,N_4993,N_4566);
and U5438 (N_5438,N_4184,N_4051);
nor U5439 (N_5439,N_4832,N_4402);
or U5440 (N_5440,N_4656,N_4297);
or U5441 (N_5441,N_4344,N_4105);
and U5442 (N_5442,N_4068,N_4955);
or U5443 (N_5443,N_4350,N_4568);
or U5444 (N_5444,N_4742,N_4108);
and U5445 (N_5445,N_4275,N_4422);
and U5446 (N_5446,N_4598,N_4585);
nand U5447 (N_5447,N_4633,N_4139);
nor U5448 (N_5448,N_4642,N_4201);
or U5449 (N_5449,N_4564,N_4392);
or U5450 (N_5450,N_4591,N_4908);
and U5451 (N_5451,N_4023,N_4979);
or U5452 (N_5452,N_4937,N_4897);
nand U5453 (N_5453,N_4944,N_4953);
nor U5454 (N_5454,N_4570,N_4588);
or U5455 (N_5455,N_4388,N_4220);
nand U5456 (N_5456,N_4122,N_4735);
nor U5457 (N_5457,N_4359,N_4237);
and U5458 (N_5458,N_4008,N_4281);
and U5459 (N_5459,N_4885,N_4784);
nor U5460 (N_5460,N_4978,N_4994);
nor U5461 (N_5461,N_4059,N_4141);
nor U5462 (N_5462,N_4244,N_4021);
nor U5463 (N_5463,N_4715,N_4193);
nand U5464 (N_5464,N_4041,N_4624);
and U5465 (N_5465,N_4617,N_4987);
or U5466 (N_5466,N_4789,N_4560);
and U5467 (N_5467,N_4412,N_4577);
nand U5468 (N_5468,N_4919,N_4423);
and U5469 (N_5469,N_4814,N_4694);
and U5470 (N_5470,N_4847,N_4533);
nor U5471 (N_5471,N_4147,N_4990);
or U5472 (N_5472,N_4526,N_4648);
nand U5473 (N_5473,N_4094,N_4176);
or U5474 (N_5474,N_4941,N_4628);
nand U5475 (N_5475,N_4724,N_4991);
nand U5476 (N_5476,N_4209,N_4442);
and U5477 (N_5477,N_4905,N_4063);
nor U5478 (N_5478,N_4549,N_4174);
nor U5479 (N_5479,N_4283,N_4249);
nor U5480 (N_5480,N_4541,N_4710);
and U5481 (N_5481,N_4471,N_4557);
nand U5482 (N_5482,N_4983,N_4601);
xnor U5483 (N_5483,N_4763,N_4736);
nor U5484 (N_5484,N_4583,N_4017);
xnor U5485 (N_5485,N_4872,N_4333);
and U5486 (N_5486,N_4723,N_4268);
or U5487 (N_5487,N_4751,N_4760);
nor U5488 (N_5488,N_4980,N_4689);
or U5489 (N_5489,N_4453,N_4650);
and U5490 (N_5490,N_4772,N_4439);
and U5491 (N_5491,N_4787,N_4317);
xnor U5492 (N_5492,N_4413,N_4339);
nand U5493 (N_5493,N_4554,N_4462);
nor U5494 (N_5494,N_4849,N_4398);
nor U5495 (N_5495,N_4015,N_4997);
or U5496 (N_5496,N_4305,N_4746);
nor U5497 (N_5497,N_4302,N_4961);
nand U5498 (N_5498,N_4653,N_4675);
and U5499 (N_5499,N_4920,N_4424);
or U5500 (N_5500,N_4034,N_4002);
or U5501 (N_5501,N_4377,N_4923);
nand U5502 (N_5502,N_4723,N_4618);
nand U5503 (N_5503,N_4794,N_4792);
and U5504 (N_5504,N_4303,N_4793);
or U5505 (N_5505,N_4586,N_4126);
nand U5506 (N_5506,N_4529,N_4543);
nor U5507 (N_5507,N_4152,N_4351);
and U5508 (N_5508,N_4083,N_4368);
or U5509 (N_5509,N_4707,N_4343);
and U5510 (N_5510,N_4955,N_4977);
nor U5511 (N_5511,N_4036,N_4001);
nand U5512 (N_5512,N_4630,N_4641);
nand U5513 (N_5513,N_4970,N_4190);
and U5514 (N_5514,N_4726,N_4357);
nand U5515 (N_5515,N_4851,N_4810);
nand U5516 (N_5516,N_4766,N_4098);
and U5517 (N_5517,N_4174,N_4031);
or U5518 (N_5518,N_4911,N_4790);
nor U5519 (N_5519,N_4483,N_4401);
and U5520 (N_5520,N_4385,N_4116);
nor U5521 (N_5521,N_4947,N_4641);
and U5522 (N_5522,N_4252,N_4664);
or U5523 (N_5523,N_4162,N_4634);
or U5524 (N_5524,N_4727,N_4171);
nand U5525 (N_5525,N_4936,N_4688);
and U5526 (N_5526,N_4921,N_4654);
nand U5527 (N_5527,N_4325,N_4062);
and U5528 (N_5528,N_4913,N_4452);
nand U5529 (N_5529,N_4900,N_4426);
and U5530 (N_5530,N_4925,N_4547);
and U5531 (N_5531,N_4236,N_4317);
nor U5532 (N_5532,N_4227,N_4913);
nor U5533 (N_5533,N_4898,N_4755);
nand U5534 (N_5534,N_4058,N_4540);
nor U5535 (N_5535,N_4584,N_4275);
nand U5536 (N_5536,N_4178,N_4492);
nor U5537 (N_5537,N_4029,N_4165);
and U5538 (N_5538,N_4030,N_4208);
xor U5539 (N_5539,N_4564,N_4888);
nand U5540 (N_5540,N_4534,N_4652);
nand U5541 (N_5541,N_4756,N_4148);
nor U5542 (N_5542,N_4926,N_4586);
or U5543 (N_5543,N_4251,N_4959);
nor U5544 (N_5544,N_4729,N_4140);
and U5545 (N_5545,N_4544,N_4088);
nand U5546 (N_5546,N_4727,N_4078);
or U5547 (N_5547,N_4741,N_4987);
and U5548 (N_5548,N_4572,N_4972);
nor U5549 (N_5549,N_4624,N_4574);
nand U5550 (N_5550,N_4987,N_4044);
nor U5551 (N_5551,N_4784,N_4795);
and U5552 (N_5552,N_4151,N_4085);
nor U5553 (N_5553,N_4788,N_4327);
nand U5554 (N_5554,N_4194,N_4632);
nand U5555 (N_5555,N_4705,N_4803);
nand U5556 (N_5556,N_4020,N_4445);
or U5557 (N_5557,N_4715,N_4496);
nand U5558 (N_5558,N_4764,N_4186);
and U5559 (N_5559,N_4858,N_4955);
and U5560 (N_5560,N_4145,N_4402);
and U5561 (N_5561,N_4652,N_4948);
and U5562 (N_5562,N_4449,N_4515);
and U5563 (N_5563,N_4025,N_4099);
nor U5564 (N_5564,N_4266,N_4737);
nand U5565 (N_5565,N_4661,N_4906);
nor U5566 (N_5566,N_4419,N_4483);
nand U5567 (N_5567,N_4512,N_4898);
or U5568 (N_5568,N_4696,N_4161);
nand U5569 (N_5569,N_4271,N_4747);
or U5570 (N_5570,N_4919,N_4582);
nor U5571 (N_5571,N_4579,N_4303);
or U5572 (N_5572,N_4327,N_4039);
or U5573 (N_5573,N_4041,N_4742);
nor U5574 (N_5574,N_4321,N_4619);
and U5575 (N_5575,N_4676,N_4062);
nand U5576 (N_5576,N_4199,N_4437);
and U5577 (N_5577,N_4586,N_4594);
nand U5578 (N_5578,N_4655,N_4695);
nand U5579 (N_5579,N_4080,N_4638);
nand U5580 (N_5580,N_4357,N_4093);
nand U5581 (N_5581,N_4684,N_4099);
or U5582 (N_5582,N_4916,N_4468);
nor U5583 (N_5583,N_4058,N_4843);
and U5584 (N_5584,N_4608,N_4084);
and U5585 (N_5585,N_4191,N_4161);
or U5586 (N_5586,N_4806,N_4087);
nor U5587 (N_5587,N_4040,N_4274);
or U5588 (N_5588,N_4607,N_4733);
nor U5589 (N_5589,N_4146,N_4268);
nor U5590 (N_5590,N_4413,N_4959);
or U5591 (N_5591,N_4540,N_4135);
and U5592 (N_5592,N_4299,N_4018);
nand U5593 (N_5593,N_4412,N_4564);
and U5594 (N_5594,N_4255,N_4848);
nor U5595 (N_5595,N_4952,N_4981);
nor U5596 (N_5596,N_4188,N_4929);
or U5597 (N_5597,N_4947,N_4280);
or U5598 (N_5598,N_4307,N_4478);
nor U5599 (N_5599,N_4336,N_4218);
or U5600 (N_5600,N_4889,N_4119);
nand U5601 (N_5601,N_4816,N_4243);
nand U5602 (N_5602,N_4411,N_4353);
and U5603 (N_5603,N_4255,N_4100);
nand U5604 (N_5604,N_4238,N_4688);
and U5605 (N_5605,N_4928,N_4783);
nand U5606 (N_5606,N_4375,N_4808);
nand U5607 (N_5607,N_4816,N_4985);
nor U5608 (N_5608,N_4790,N_4607);
or U5609 (N_5609,N_4321,N_4382);
nand U5610 (N_5610,N_4535,N_4955);
nand U5611 (N_5611,N_4822,N_4044);
and U5612 (N_5612,N_4812,N_4103);
nand U5613 (N_5613,N_4659,N_4691);
and U5614 (N_5614,N_4995,N_4224);
and U5615 (N_5615,N_4271,N_4609);
nand U5616 (N_5616,N_4532,N_4714);
nand U5617 (N_5617,N_4545,N_4326);
nand U5618 (N_5618,N_4927,N_4964);
nor U5619 (N_5619,N_4904,N_4508);
or U5620 (N_5620,N_4154,N_4608);
and U5621 (N_5621,N_4400,N_4344);
and U5622 (N_5622,N_4248,N_4886);
and U5623 (N_5623,N_4957,N_4484);
nor U5624 (N_5624,N_4792,N_4673);
or U5625 (N_5625,N_4669,N_4476);
nand U5626 (N_5626,N_4579,N_4401);
nor U5627 (N_5627,N_4726,N_4825);
or U5628 (N_5628,N_4036,N_4226);
nor U5629 (N_5629,N_4464,N_4850);
or U5630 (N_5630,N_4907,N_4948);
or U5631 (N_5631,N_4878,N_4338);
nor U5632 (N_5632,N_4260,N_4608);
nor U5633 (N_5633,N_4949,N_4066);
or U5634 (N_5634,N_4047,N_4693);
nand U5635 (N_5635,N_4048,N_4119);
nand U5636 (N_5636,N_4543,N_4158);
and U5637 (N_5637,N_4483,N_4992);
nor U5638 (N_5638,N_4585,N_4871);
or U5639 (N_5639,N_4703,N_4054);
nor U5640 (N_5640,N_4643,N_4985);
or U5641 (N_5641,N_4620,N_4898);
nor U5642 (N_5642,N_4542,N_4393);
nor U5643 (N_5643,N_4383,N_4633);
nand U5644 (N_5644,N_4275,N_4158);
nand U5645 (N_5645,N_4716,N_4146);
nand U5646 (N_5646,N_4212,N_4228);
or U5647 (N_5647,N_4282,N_4636);
or U5648 (N_5648,N_4637,N_4041);
nor U5649 (N_5649,N_4966,N_4465);
nor U5650 (N_5650,N_4920,N_4209);
nor U5651 (N_5651,N_4446,N_4200);
nor U5652 (N_5652,N_4464,N_4049);
nand U5653 (N_5653,N_4968,N_4912);
and U5654 (N_5654,N_4136,N_4698);
nor U5655 (N_5655,N_4580,N_4354);
nand U5656 (N_5656,N_4205,N_4882);
nor U5657 (N_5657,N_4088,N_4704);
and U5658 (N_5658,N_4546,N_4338);
nor U5659 (N_5659,N_4920,N_4004);
and U5660 (N_5660,N_4052,N_4405);
and U5661 (N_5661,N_4296,N_4769);
xnor U5662 (N_5662,N_4101,N_4348);
nand U5663 (N_5663,N_4215,N_4784);
nand U5664 (N_5664,N_4026,N_4571);
and U5665 (N_5665,N_4353,N_4802);
and U5666 (N_5666,N_4909,N_4694);
or U5667 (N_5667,N_4994,N_4232);
and U5668 (N_5668,N_4028,N_4558);
or U5669 (N_5669,N_4697,N_4262);
and U5670 (N_5670,N_4284,N_4725);
or U5671 (N_5671,N_4181,N_4413);
nor U5672 (N_5672,N_4122,N_4010);
nand U5673 (N_5673,N_4907,N_4884);
and U5674 (N_5674,N_4777,N_4151);
or U5675 (N_5675,N_4292,N_4866);
or U5676 (N_5676,N_4336,N_4706);
nor U5677 (N_5677,N_4015,N_4702);
or U5678 (N_5678,N_4108,N_4924);
nand U5679 (N_5679,N_4932,N_4230);
or U5680 (N_5680,N_4669,N_4550);
and U5681 (N_5681,N_4313,N_4002);
or U5682 (N_5682,N_4799,N_4196);
nand U5683 (N_5683,N_4449,N_4399);
nor U5684 (N_5684,N_4493,N_4964);
or U5685 (N_5685,N_4353,N_4984);
xnor U5686 (N_5686,N_4133,N_4793);
or U5687 (N_5687,N_4839,N_4680);
or U5688 (N_5688,N_4072,N_4262);
or U5689 (N_5689,N_4815,N_4426);
and U5690 (N_5690,N_4242,N_4626);
or U5691 (N_5691,N_4193,N_4380);
or U5692 (N_5692,N_4416,N_4183);
nand U5693 (N_5693,N_4865,N_4501);
and U5694 (N_5694,N_4791,N_4802);
nand U5695 (N_5695,N_4213,N_4540);
nor U5696 (N_5696,N_4301,N_4483);
and U5697 (N_5697,N_4952,N_4341);
and U5698 (N_5698,N_4787,N_4018);
nand U5699 (N_5699,N_4325,N_4960);
nor U5700 (N_5700,N_4510,N_4706);
nor U5701 (N_5701,N_4305,N_4180);
and U5702 (N_5702,N_4719,N_4148);
nor U5703 (N_5703,N_4422,N_4486);
nor U5704 (N_5704,N_4266,N_4401);
nor U5705 (N_5705,N_4440,N_4800);
or U5706 (N_5706,N_4370,N_4299);
or U5707 (N_5707,N_4454,N_4498);
and U5708 (N_5708,N_4243,N_4419);
nor U5709 (N_5709,N_4794,N_4260);
nor U5710 (N_5710,N_4922,N_4875);
nor U5711 (N_5711,N_4173,N_4951);
nor U5712 (N_5712,N_4956,N_4543);
nand U5713 (N_5713,N_4980,N_4227);
and U5714 (N_5714,N_4922,N_4590);
nor U5715 (N_5715,N_4903,N_4067);
nor U5716 (N_5716,N_4977,N_4862);
xor U5717 (N_5717,N_4146,N_4025);
or U5718 (N_5718,N_4559,N_4718);
nor U5719 (N_5719,N_4179,N_4521);
nand U5720 (N_5720,N_4201,N_4765);
or U5721 (N_5721,N_4223,N_4025);
or U5722 (N_5722,N_4278,N_4123);
nand U5723 (N_5723,N_4648,N_4843);
and U5724 (N_5724,N_4621,N_4228);
nand U5725 (N_5725,N_4804,N_4703);
or U5726 (N_5726,N_4512,N_4393);
or U5727 (N_5727,N_4203,N_4259);
nor U5728 (N_5728,N_4253,N_4676);
and U5729 (N_5729,N_4023,N_4491);
nand U5730 (N_5730,N_4490,N_4196);
or U5731 (N_5731,N_4227,N_4856);
xor U5732 (N_5732,N_4963,N_4492);
and U5733 (N_5733,N_4218,N_4502);
or U5734 (N_5734,N_4221,N_4050);
nand U5735 (N_5735,N_4723,N_4653);
nor U5736 (N_5736,N_4050,N_4022);
and U5737 (N_5737,N_4753,N_4662);
or U5738 (N_5738,N_4292,N_4716);
nor U5739 (N_5739,N_4629,N_4182);
or U5740 (N_5740,N_4688,N_4043);
nor U5741 (N_5741,N_4796,N_4419);
or U5742 (N_5742,N_4783,N_4807);
nand U5743 (N_5743,N_4110,N_4711);
nand U5744 (N_5744,N_4049,N_4544);
or U5745 (N_5745,N_4802,N_4678);
nand U5746 (N_5746,N_4465,N_4053);
nand U5747 (N_5747,N_4752,N_4748);
nand U5748 (N_5748,N_4052,N_4310);
and U5749 (N_5749,N_4993,N_4513);
or U5750 (N_5750,N_4664,N_4901);
or U5751 (N_5751,N_4894,N_4936);
or U5752 (N_5752,N_4477,N_4532);
and U5753 (N_5753,N_4050,N_4403);
nand U5754 (N_5754,N_4826,N_4814);
and U5755 (N_5755,N_4550,N_4544);
nor U5756 (N_5756,N_4678,N_4044);
or U5757 (N_5757,N_4863,N_4908);
and U5758 (N_5758,N_4327,N_4772);
and U5759 (N_5759,N_4396,N_4874);
and U5760 (N_5760,N_4500,N_4514);
nor U5761 (N_5761,N_4599,N_4769);
and U5762 (N_5762,N_4952,N_4138);
and U5763 (N_5763,N_4614,N_4210);
or U5764 (N_5764,N_4230,N_4542);
or U5765 (N_5765,N_4595,N_4928);
nand U5766 (N_5766,N_4468,N_4923);
nor U5767 (N_5767,N_4663,N_4886);
and U5768 (N_5768,N_4214,N_4480);
and U5769 (N_5769,N_4617,N_4637);
nor U5770 (N_5770,N_4609,N_4769);
or U5771 (N_5771,N_4375,N_4835);
and U5772 (N_5772,N_4481,N_4595);
nand U5773 (N_5773,N_4609,N_4489);
and U5774 (N_5774,N_4298,N_4665);
nor U5775 (N_5775,N_4520,N_4300);
and U5776 (N_5776,N_4047,N_4940);
and U5777 (N_5777,N_4053,N_4441);
and U5778 (N_5778,N_4274,N_4596);
nor U5779 (N_5779,N_4272,N_4253);
or U5780 (N_5780,N_4192,N_4507);
or U5781 (N_5781,N_4755,N_4513);
or U5782 (N_5782,N_4304,N_4882);
nor U5783 (N_5783,N_4261,N_4162);
and U5784 (N_5784,N_4996,N_4213);
nand U5785 (N_5785,N_4249,N_4221);
or U5786 (N_5786,N_4697,N_4805);
nand U5787 (N_5787,N_4376,N_4037);
or U5788 (N_5788,N_4532,N_4758);
xor U5789 (N_5789,N_4293,N_4664);
or U5790 (N_5790,N_4873,N_4795);
nor U5791 (N_5791,N_4777,N_4597);
or U5792 (N_5792,N_4315,N_4152);
xor U5793 (N_5793,N_4934,N_4583);
nor U5794 (N_5794,N_4721,N_4363);
nand U5795 (N_5795,N_4097,N_4236);
and U5796 (N_5796,N_4714,N_4682);
nand U5797 (N_5797,N_4597,N_4316);
nor U5798 (N_5798,N_4494,N_4337);
and U5799 (N_5799,N_4967,N_4506);
nand U5800 (N_5800,N_4862,N_4404);
or U5801 (N_5801,N_4854,N_4197);
nand U5802 (N_5802,N_4835,N_4877);
and U5803 (N_5803,N_4187,N_4608);
and U5804 (N_5804,N_4823,N_4152);
or U5805 (N_5805,N_4587,N_4559);
or U5806 (N_5806,N_4916,N_4923);
or U5807 (N_5807,N_4970,N_4030);
nor U5808 (N_5808,N_4970,N_4247);
nand U5809 (N_5809,N_4840,N_4693);
nor U5810 (N_5810,N_4612,N_4104);
nand U5811 (N_5811,N_4847,N_4139);
nor U5812 (N_5812,N_4550,N_4054);
nor U5813 (N_5813,N_4552,N_4152);
or U5814 (N_5814,N_4876,N_4616);
and U5815 (N_5815,N_4157,N_4193);
and U5816 (N_5816,N_4305,N_4327);
or U5817 (N_5817,N_4172,N_4648);
and U5818 (N_5818,N_4921,N_4807);
nand U5819 (N_5819,N_4541,N_4784);
nand U5820 (N_5820,N_4286,N_4519);
nor U5821 (N_5821,N_4508,N_4429);
and U5822 (N_5822,N_4222,N_4565);
nand U5823 (N_5823,N_4609,N_4918);
or U5824 (N_5824,N_4304,N_4911);
or U5825 (N_5825,N_4102,N_4974);
and U5826 (N_5826,N_4707,N_4286);
or U5827 (N_5827,N_4641,N_4170);
or U5828 (N_5828,N_4363,N_4113);
nand U5829 (N_5829,N_4222,N_4487);
and U5830 (N_5830,N_4670,N_4356);
nand U5831 (N_5831,N_4757,N_4835);
nor U5832 (N_5832,N_4846,N_4143);
nand U5833 (N_5833,N_4165,N_4095);
and U5834 (N_5834,N_4484,N_4520);
nand U5835 (N_5835,N_4781,N_4171);
nor U5836 (N_5836,N_4977,N_4882);
and U5837 (N_5837,N_4086,N_4072);
nand U5838 (N_5838,N_4308,N_4192);
nor U5839 (N_5839,N_4655,N_4056);
and U5840 (N_5840,N_4456,N_4514);
nand U5841 (N_5841,N_4989,N_4291);
nor U5842 (N_5842,N_4938,N_4972);
nor U5843 (N_5843,N_4539,N_4955);
or U5844 (N_5844,N_4244,N_4246);
nand U5845 (N_5845,N_4914,N_4868);
nand U5846 (N_5846,N_4867,N_4424);
or U5847 (N_5847,N_4172,N_4427);
nand U5848 (N_5848,N_4045,N_4018);
and U5849 (N_5849,N_4729,N_4438);
nor U5850 (N_5850,N_4269,N_4638);
nor U5851 (N_5851,N_4785,N_4554);
nor U5852 (N_5852,N_4100,N_4175);
and U5853 (N_5853,N_4791,N_4514);
and U5854 (N_5854,N_4781,N_4609);
nand U5855 (N_5855,N_4494,N_4647);
nand U5856 (N_5856,N_4666,N_4736);
and U5857 (N_5857,N_4331,N_4240);
and U5858 (N_5858,N_4351,N_4729);
or U5859 (N_5859,N_4875,N_4414);
and U5860 (N_5860,N_4712,N_4423);
and U5861 (N_5861,N_4760,N_4051);
or U5862 (N_5862,N_4163,N_4782);
and U5863 (N_5863,N_4048,N_4353);
or U5864 (N_5864,N_4176,N_4891);
nor U5865 (N_5865,N_4332,N_4148);
and U5866 (N_5866,N_4783,N_4224);
and U5867 (N_5867,N_4583,N_4637);
nor U5868 (N_5868,N_4935,N_4555);
and U5869 (N_5869,N_4751,N_4205);
and U5870 (N_5870,N_4907,N_4151);
and U5871 (N_5871,N_4775,N_4675);
nor U5872 (N_5872,N_4533,N_4080);
or U5873 (N_5873,N_4832,N_4257);
nand U5874 (N_5874,N_4067,N_4095);
nor U5875 (N_5875,N_4332,N_4843);
nand U5876 (N_5876,N_4075,N_4772);
nand U5877 (N_5877,N_4171,N_4178);
or U5878 (N_5878,N_4782,N_4109);
nand U5879 (N_5879,N_4899,N_4731);
nand U5880 (N_5880,N_4508,N_4326);
nand U5881 (N_5881,N_4373,N_4868);
and U5882 (N_5882,N_4371,N_4581);
nor U5883 (N_5883,N_4030,N_4960);
or U5884 (N_5884,N_4416,N_4618);
or U5885 (N_5885,N_4422,N_4835);
and U5886 (N_5886,N_4225,N_4224);
nor U5887 (N_5887,N_4865,N_4058);
nand U5888 (N_5888,N_4496,N_4464);
nand U5889 (N_5889,N_4426,N_4872);
and U5890 (N_5890,N_4447,N_4520);
and U5891 (N_5891,N_4140,N_4840);
or U5892 (N_5892,N_4926,N_4078);
and U5893 (N_5893,N_4980,N_4041);
and U5894 (N_5894,N_4382,N_4004);
nand U5895 (N_5895,N_4387,N_4823);
nor U5896 (N_5896,N_4141,N_4758);
and U5897 (N_5897,N_4982,N_4376);
nand U5898 (N_5898,N_4239,N_4243);
or U5899 (N_5899,N_4376,N_4086);
and U5900 (N_5900,N_4238,N_4513);
and U5901 (N_5901,N_4410,N_4752);
and U5902 (N_5902,N_4959,N_4816);
and U5903 (N_5903,N_4376,N_4323);
nor U5904 (N_5904,N_4217,N_4376);
nand U5905 (N_5905,N_4144,N_4924);
or U5906 (N_5906,N_4667,N_4087);
nand U5907 (N_5907,N_4176,N_4544);
or U5908 (N_5908,N_4126,N_4958);
nand U5909 (N_5909,N_4550,N_4422);
or U5910 (N_5910,N_4317,N_4704);
nor U5911 (N_5911,N_4394,N_4840);
or U5912 (N_5912,N_4052,N_4691);
nand U5913 (N_5913,N_4049,N_4495);
nand U5914 (N_5914,N_4914,N_4503);
or U5915 (N_5915,N_4992,N_4740);
and U5916 (N_5916,N_4163,N_4461);
or U5917 (N_5917,N_4303,N_4311);
or U5918 (N_5918,N_4051,N_4958);
or U5919 (N_5919,N_4155,N_4550);
or U5920 (N_5920,N_4840,N_4223);
nand U5921 (N_5921,N_4061,N_4602);
nor U5922 (N_5922,N_4405,N_4313);
nand U5923 (N_5923,N_4324,N_4779);
and U5924 (N_5924,N_4434,N_4246);
or U5925 (N_5925,N_4430,N_4959);
and U5926 (N_5926,N_4130,N_4171);
nand U5927 (N_5927,N_4705,N_4161);
xor U5928 (N_5928,N_4852,N_4023);
nor U5929 (N_5929,N_4870,N_4173);
nor U5930 (N_5930,N_4260,N_4467);
nand U5931 (N_5931,N_4332,N_4462);
and U5932 (N_5932,N_4531,N_4320);
or U5933 (N_5933,N_4261,N_4347);
and U5934 (N_5934,N_4319,N_4637);
nand U5935 (N_5935,N_4552,N_4140);
and U5936 (N_5936,N_4830,N_4932);
nor U5937 (N_5937,N_4060,N_4421);
or U5938 (N_5938,N_4056,N_4093);
nor U5939 (N_5939,N_4412,N_4112);
and U5940 (N_5940,N_4879,N_4257);
and U5941 (N_5941,N_4667,N_4695);
or U5942 (N_5942,N_4729,N_4770);
nand U5943 (N_5943,N_4005,N_4987);
or U5944 (N_5944,N_4383,N_4737);
and U5945 (N_5945,N_4982,N_4842);
nand U5946 (N_5946,N_4354,N_4606);
or U5947 (N_5947,N_4492,N_4914);
nand U5948 (N_5948,N_4422,N_4459);
and U5949 (N_5949,N_4179,N_4670);
nand U5950 (N_5950,N_4234,N_4270);
or U5951 (N_5951,N_4852,N_4651);
nand U5952 (N_5952,N_4702,N_4001);
or U5953 (N_5953,N_4257,N_4404);
or U5954 (N_5954,N_4851,N_4939);
nor U5955 (N_5955,N_4018,N_4228);
or U5956 (N_5956,N_4313,N_4844);
or U5957 (N_5957,N_4033,N_4412);
and U5958 (N_5958,N_4161,N_4570);
nor U5959 (N_5959,N_4537,N_4139);
nor U5960 (N_5960,N_4195,N_4897);
or U5961 (N_5961,N_4080,N_4464);
nor U5962 (N_5962,N_4205,N_4811);
nand U5963 (N_5963,N_4116,N_4749);
and U5964 (N_5964,N_4599,N_4479);
nand U5965 (N_5965,N_4256,N_4400);
or U5966 (N_5966,N_4295,N_4889);
or U5967 (N_5967,N_4881,N_4549);
nor U5968 (N_5968,N_4230,N_4570);
and U5969 (N_5969,N_4573,N_4965);
or U5970 (N_5970,N_4191,N_4818);
nor U5971 (N_5971,N_4633,N_4173);
nand U5972 (N_5972,N_4489,N_4029);
and U5973 (N_5973,N_4685,N_4958);
nor U5974 (N_5974,N_4031,N_4221);
nand U5975 (N_5975,N_4452,N_4498);
or U5976 (N_5976,N_4685,N_4590);
or U5977 (N_5977,N_4782,N_4445);
or U5978 (N_5978,N_4664,N_4693);
nor U5979 (N_5979,N_4373,N_4019);
nand U5980 (N_5980,N_4873,N_4826);
nor U5981 (N_5981,N_4095,N_4061);
nand U5982 (N_5982,N_4977,N_4060);
or U5983 (N_5983,N_4797,N_4049);
nand U5984 (N_5984,N_4661,N_4351);
nor U5985 (N_5985,N_4109,N_4310);
nand U5986 (N_5986,N_4730,N_4767);
or U5987 (N_5987,N_4190,N_4475);
nand U5988 (N_5988,N_4133,N_4794);
nand U5989 (N_5989,N_4439,N_4188);
nand U5990 (N_5990,N_4077,N_4141);
nor U5991 (N_5991,N_4174,N_4252);
and U5992 (N_5992,N_4377,N_4826);
and U5993 (N_5993,N_4958,N_4687);
and U5994 (N_5994,N_4667,N_4029);
nor U5995 (N_5995,N_4427,N_4924);
or U5996 (N_5996,N_4020,N_4696);
nor U5997 (N_5997,N_4656,N_4709);
nor U5998 (N_5998,N_4715,N_4189);
or U5999 (N_5999,N_4416,N_4313);
nand U6000 (N_6000,N_5004,N_5421);
or U6001 (N_6001,N_5966,N_5057);
nand U6002 (N_6002,N_5969,N_5326);
nor U6003 (N_6003,N_5587,N_5566);
nor U6004 (N_6004,N_5740,N_5558);
and U6005 (N_6005,N_5138,N_5096);
and U6006 (N_6006,N_5839,N_5881);
and U6007 (N_6007,N_5619,N_5127);
nor U6008 (N_6008,N_5997,N_5649);
or U6009 (N_6009,N_5202,N_5098);
and U6010 (N_6010,N_5122,N_5471);
xor U6011 (N_6011,N_5840,N_5778);
and U6012 (N_6012,N_5808,N_5699);
nor U6013 (N_6013,N_5894,N_5938);
nand U6014 (N_6014,N_5199,N_5152);
and U6015 (N_6015,N_5119,N_5251);
or U6016 (N_6016,N_5815,N_5963);
nor U6017 (N_6017,N_5356,N_5504);
nand U6018 (N_6018,N_5606,N_5920);
xnor U6019 (N_6019,N_5351,N_5091);
nand U6020 (N_6020,N_5018,N_5427);
xor U6021 (N_6021,N_5424,N_5365);
or U6022 (N_6022,N_5375,N_5035);
or U6023 (N_6023,N_5039,N_5784);
xor U6024 (N_6024,N_5249,N_5209);
nor U6025 (N_6025,N_5716,N_5368);
or U6026 (N_6026,N_5385,N_5491);
or U6027 (N_6027,N_5232,N_5627);
nor U6028 (N_6028,N_5506,N_5306);
nand U6029 (N_6029,N_5450,N_5792);
and U6030 (N_6030,N_5156,N_5182);
or U6031 (N_6031,N_5392,N_5257);
nor U6032 (N_6032,N_5522,N_5547);
nor U6033 (N_6033,N_5794,N_5694);
nand U6034 (N_6034,N_5975,N_5541);
or U6035 (N_6035,N_5618,N_5086);
nor U6036 (N_6036,N_5419,N_5610);
nor U6037 (N_6037,N_5540,N_5790);
or U6038 (N_6038,N_5067,N_5492);
or U6039 (N_6039,N_5988,N_5551);
and U6040 (N_6040,N_5171,N_5296);
or U6041 (N_6041,N_5775,N_5494);
and U6042 (N_6042,N_5561,N_5668);
and U6043 (N_6043,N_5638,N_5343);
or U6044 (N_6044,N_5193,N_5749);
nor U6045 (N_6045,N_5016,N_5274);
and U6046 (N_6046,N_5115,N_5885);
nor U6047 (N_6047,N_5639,N_5810);
nor U6048 (N_6048,N_5349,N_5761);
and U6049 (N_6049,N_5032,N_5484);
nand U6050 (N_6050,N_5361,N_5636);
nor U6051 (N_6051,N_5594,N_5940);
or U6052 (N_6052,N_5855,N_5329);
xor U6053 (N_6053,N_5560,N_5283);
or U6054 (N_6054,N_5178,N_5173);
nor U6055 (N_6055,N_5085,N_5876);
nor U6056 (N_6056,N_5317,N_5160);
or U6057 (N_6057,N_5137,N_5764);
and U6058 (N_6058,N_5889,N_5516);
and U6059 (N_6059,N_5316,N_5493);
nand U6060 (N_6060,N_5413,N_5222);
nor U6061 (N_6061,N_5254,N_5913);
or U6062 (N_6062,N_5422,N_5463);
or U6063 (N_6063,N_5981,N_5549);
nand U6064 (N_6064,N_5847,N_5212);
xnor U6065 (N_6065,N_5866,N_5366);
and U6066 (N_6066,N_5322,N_5256);
nor U6067 (N_6067,N_5056,N_5060);
and U6068 (N_6068,N_5945,N_5025);
or U6069 (N_6069,N_5809,N_5722);
nor U6070 (N_6070,N_5169,N_5744);
or U6071 (N_6071,N_5403,N_5191);
and U6072 (N_6072,N_5844,N_5872);
or U6073 (N_6073,N_5243,N_5724);
nand U6074 (N_6074,N_5479,N_5539);
or U6075 (N_6075,N_5512,N_5175);
nand U6076 (N_6076,N_5336,N_5405);
and U6077 (N_6077,N_5933,N_5011);
nor U6078 (N_6078,N_5519,N_5475);
or U6079 (N_6079,N_5782,N_5674);
nand U6080 (N_6080,N_5497,N_5428);
nand U6081 (N_6081,N_5581,N_5298);
nor U6082 (N_6082,N_5440,N_5962);
and U6083 (N_6083,N_5164,N_5895);
nand U6084 (N_6084,N_5373,N_5412);
nor U6085 (N_6085,N_5576,N_5635);
nor U6086 (N_6086,N_5134,N_5604);
or U6087 (N_6087,N_5629,N_5667);
and U6088 (N_6088,N_5457,N_5353);
or U6089 (N_6089,N_5906,N_5888);
and U6090 (N_6090,N_5672,N_5731);
nand U6091 (N_6091,N_5118,N_5991);
nor U6092 (N_6092,N_5605,N_5686);
or U6093 (N_6093,N_5609,N_5733);
and U6094 (N_6094,N_5781,N_5632);
nor U6095 (N_6095,N_5684,N_5009);
or U6096 (N_6096,N_5931,N_5341);
and U6097 (N_6097,N_5281,N_5544);
nor U6098 (N_6098,N_5350,N_5758);
and U6099 (N_6099,N_5460,N_5130);
nand U6100 (N_6100,N_5150,N_5853);
nor U6101 (N_6101,N_5584,N_5472);
nor U6102 (N_6102,N_5346,N_5532);
nand U6103 (N_6103,N_5564,N_5569);
or U6104 (N_6104,N_5364,N_5452);
or U6105 (N_6105,N_5950,N_5803);
nor U6106 (N_6106,N_5624,N_5465);
and U6107 (N_6107,N_5528,N_5650);
nor U6108 (N_6108,N_5395,N_5340);
and U6109 (N_6109,N_5029,N_5290);
nand U6110 (N_6110,N_5603,N_5299);
nand U6111 (N_6111,N_5633,N_5867);
nand U6112 (N_6112,N_5661,N_5623);
or U6113 (N_6113,N_5978,N_5214);
or U6114 (N_6114,N_5687,N_5344);
nand U6115 (N_6115,N_5875,N_5683);
or U6116 (N_6116,N_5148,N_5613);
nand U6117 (N_6117,N_5843,N_5027);
or U6118 (N_6118,N_5158,N_5240);
nand U6119 (N_6119,N_5197,N_5359);
or U6120 (N_6120,N_5964,N_5830);
nand U6121 (N_6121,N_5458,N_5703);
nand U6122 (N_6122,N_5741,N_5402);
nor U6123 (N_6123,N_5267,N_5262);
nand U6124 (N_6124,N_5600,N_5088);
and U6125 (N_6125,N_5985,N_5655);
nand U6126 (N_6126,N_5320,N_5024);
nand U6127 (N_6127,N_5126,N_5878);
or U6128 (N_6128,N_5147,N_5410);
nand U6129 (N_6129,N_5313,N_5841);
and U6130 (N_6130,N_5498,N_5729);
nand U6131 (N_6131,N_5480,N_5332);
nor U6132 (N_6132,N_5300,N_5064);
nand U6133 (N_6133,N_5101,N_5012);
nor U6134 (N_6134,N_5242,N_5297);
and U6135 (N_6135,N_5534,N_5080);
and U6136 (N_6136,N_5562,N_5223);
and U6137 (N_6137,N_5614,N_5951);
nor U6138 (N_6138,N_5189,N_5932);
or U6139 (N_6139,N_5074,N_5508);
nor U6140 (N_6140,N_5928,N_5415);
nand U6141 (N_6141,N_5241,N_5244);
nor U6142 (N_6142,N_5631,N_5800);
or U6143 (N_6143,N_5078,N_5165);
and U6144 (N_6144,N_5153,N_5593);
nand U6145 (N_6145,N_5167,N_5184);
or U6146 (N_6146,N_5280,N_5807);
or U6147 (N_6147,N_5858,N_5213);
xor U6148 (N_6148,N_5176,N_5545);
nor U6149 (N_6149,N_5579,N_5974);
nor U6150 (N_6150,N_5260,N_5909);
and U6151 (N_6151,N_5680,N_5899);
and U6152 (N_6152,N_5367,N_5669);
and U6153 (N_6153,N_5082,N_5575);
and U6154 (N_6154,N_5112,N_5712);
nor U6155 (N_6155,N_5651,N_5166);
nand U6156 (N_6156,N_5771,N_5658);
and U6157 (N_6157,N_5537,N_5058);
and U6158 (N_6158,N_5221,N_5620);
and U6159 (N_6159,N_5690,N_5521);
and U6160 (N_6160,N_5210,N_5907);
or U6161 (N_6161,N_5665,N_5128);
nor U6162 (N_6162,N_5753,N_5666);
nand U6163 (N_6163,N_5510,N_5076);
or U6164 (N_6164,N_5959,N_5507);
or U6165 (N_6165,N_5026,N_5826);
nand U6166 (N_6166,N_5580,N_5999);
and U6167 (N_6167,N_5490,N_5805);
or U6168 (N_6168,N_5760,N_5338);
and U6169 (N_6169,N_5929,N_5161);
or U6170 (N_6170,N_5124,N_5235);
or U6171 (N_6171,N_5390,N_5796);
xor U6172 (N_6172,N_5116,N_5383);
nor U6173 (N_6173,N_5070,N_5588);
or U6174 (N_6174,N_5864,N_5530);
nand U6175 (N_6175,N_5533,N_5892);
nand U6176 (N_6176,N_5890,N_5113);
and U6177 (N_6177,N_5149,N_5391);
nand U6178 (N_6178,N_5984,N_5615);
nand U6179 (N_6179,N_5005,N_5045);
nor U6180 (N_6180,N_5469,N_5496);
nand U6181 (N_6181,N_5372,N_5400);
nor U6182 (N_6182,N_5114,N_5611);
or U6183 (N_6183,N_5990,N_5279);
or U6184 (N_6184,N_5308,N_5448);
nor U6185 (N_6185,N_5947,N_5718);
and U6186 (N_6186,N_5312,N_5411);
nand U6187 (N_6187,N_5259,N_5717);
and U6188 (N_6188,N_5220,N_5766);
nand U6189 (N_6189,N_5965,N_5157);
or U6190 (N_6190,N_5132,N_5047);
and U6191 (N_6191,N_5289,N_5218);
nand U6192 (N_6192,N_5812,N_5386);
nor U6193 (N_6193,N_5704,N_5677);
and U6194 (N_6194,N_5832,N_5739);
and U6195 (N_6195,N_5897,N_5466);
nor U6196 (N_6196,N_5068,N_5430);
and U6197 (N_6197,N_5468,N_5657);
nor U6198 (N_6198,N_5154,N_5676);
and U6199 (N_6199,N_5902,N_5179);
nand U6200 (N_6200,N_5871,N_5816);
or U6201 (N_6201,N_5905,N_5592);
nor U6202 (N_6202,N_5865,N_5567);
nand U6203 (N_6203,N_5354,N_5204);
or U6204 (N_6204,N_5886,N_5162);
nor U6205 (N_6205,N_5662,N_5488);
and U6206 (N_6206,N_5002,N_5489);
or U6207 (N_6207,N_5084,N_5535);
or U6208 (N_6208,N_5526,N_5735);
nand U6209 (N_6209,N_5310,N_5224);
or U6210 (N_6210,N_5315,N_5713);
and U6211 (N_6211,N_5925,N_5837);
and U6212 (N_6212,N_5813,N_5461);
and U6213 (N_6213,N_5656,N_5647);
or U6214 (N_6214,N_5783,N_5467);
and U6215 (N_6215,N_5319,N_5525);
nand U6216 (N_6216,N_5277,N_5327);
nor U6217 (N_6217,N_5337,N_5598);
or U6218 (N_6218,N_5125,N_5763);
and U6219 (N_6219,N_5013,N_5948);
or U6220 (N_6220,N_5958,N_5845);
nand U6221 (N_6221,N_5887,N_5833);
or U6222 (N_6222,N_5986,N_5660);
nand U6223 (N_6223,N_5325,N_5989);
nand U6224 (N_6224,N_5836,N_5087);
or U6225 (N_6225,N_5955,N_5170);
and U6226 (N_6226,N_5123,N_5314);
or U6227 (N_6227,N_5001,N_5630);
and U6228 (N_6228,N_5198,N_5095);
nand U6229 (N_6229,N_5725,N_5228);
and U6230 (N_6230,N_5755,N_5896);
nand U6231 (N_6231,N_5653,N_5707);
nand U6232 (N_6232,N_5245,N_5416);
nor U6233 (N_6233,N_5053,N_5303);
and U6234 (N_6234,N_5476,N_5563);
or U6235 (N_6235,N_5520,N_5767);
nor U6236 (N_6236,N_5486,N_5384);
or U6237 (N_6237,N_5565,N_5092);
nand U6238 (N_6238,N_5120,N_5229);
or U6239 (N_6239,N_5916,N_5028);
or U6240 (N_6240,N_5689,N_5834);
nand U6241 (N_6241,N_5608,N_5922);
nor U6242 (N_6242,N_5456,N_5570);
or U6243 (N_6243,N_5140,N_5040);
and U6244 (N_6244,N_5518,N_5443);
and U6245 (N_6245,N_5023,N_5720);
nand U6246 (N_6246,N_5206,N_5129);
nor U6247 (N_6247,N_5473,N_5747);
nand U6248 (N_6248,N_5451,N_5436);
nand U6249 (N_6249,N_5139,N_5874);
nor U6250 (N_6250,N_5652,N_5555);
or U6251 (N_6251,N_5578,N_5190);
or U6252 (N_6252,N_5856,N_5706);
nor U6253 (N_6253,N_5641,N_5482);
or U6254 (N_6254,N_5301,N_5972);
and U6255 (N_6255,N_5982,N_5524);
and U6256 (N_6256,N_5953,N_5265);
or U6257 (N_6257,N_5770,N_5993);
and U6258 (N_6258,N_5247,N_5216);
nand U6259 (N_6259,N_5726,N_5441);
nand U6260 (N_6260,N_5513,N_5234);
nor U6261 (N_6261,N_5681,N_5846);
or U6262 (N_6262,N_5934,N_5601);
nor U6263 (N_6263,N_5709,N_5659);
or U6264 (N_6264,N_5015,N_5215);
nor U6265 (N_6265,N_5069,N_5898);
nor U6266 (N_6266,N_5924,N_5585);
nor U6267 (N_6267,N_5671,N_5302);
or U6268 (N_6268,N_5106,N_5250);
or U6269 (N_6269,N_5330,N_5284);
and U6270 (N_6270,N_5935,N_5414);
or U6271 (N_6271,N_5995,N_5737);
nand U6272 (N_6272,N_5939,N_5263);
nand U6273 (N_6273,N_5347,N_5177);
or U6274 (N_6274,N_5432,N_5180);
nor U6275 (N_6275,N_5599,N_5102);
and U6276 (N_6276,N_5970,N_5863);
nor U6277 (N_6277,N_5799,N_5976);
nor U6278 (N_6278,N_5750,N_5646);
nor U6279 (N_6279,N_5501,N_5577);
and U6280 (N_6280,N_5062,N_5246);
nor U6281 (N_6281,N_5051,N_5702);
nand U6282 (N_6282,N_5675,N_5954);
nand U6283 (N_6283,N_5044,N_5318);
or U6284 (N_6284,N_5854,N_5517);
nor U6285 (N_6285,N_5882,N_5200);
and U6286 (N_6286,N_5333,N_5374);
nor U6287 (N_6287,N_5762,N_5968);
or U6288 (N_6288,N_5961,N_5435);
or U6289 (N_6289,N_5582,N_5503);
nor U6290 (N_6290,N_5207,N_5185);
or U6291 (N_6291,N_5055,N_5802);
or U6292 (N_6292,N_5362,N_5879);
xnor U6293 (N_6293,N_5914,N_5117);
nor U6294 (N_6294,N_5977,N_5335);
and U6295 (N_6295,N_5369,N_5742);
and U6296 (N_6296,N_5143,N_5957);
nand U6297 (N_6297,N_5678,N_5546);
and U6298 (N_6298,N_5930,N_5100);
nor U6299 (N_6299,N_5192,N_5291);
or U6300 (N_6300,N_5110,N_5926);
or U6301 (N_6301,N_5891,N_5514);
nand U6302 (N_6302,N_5828,N_5328);
and U6303 (N_6303,N_5033,N_5688);
nand U6304 (N_6304,N_5304,N_5278);
nor U6305 (N_6305,N_5168,N_5949);
or U6306 (N_6306,N_5942,N_5048);
nor U6307 (N_6307,N_5000,N_5648);
or U6308 (N_6308,N_5772,N_5459);
nand U6309 (N_6309,N_5987,N_5081);
and U6310 (N_6310,N_5380,N_5208);
and U6311 (N_6311,N_5034,N_5342);
nor U6312 (N_6312,N_5821,N_5073);
or U6313 (N_6313,N_5923,N_5746);
nor U6314 (N_6314,N_5483,N_5823);
nor U6315 (N_6315,N_5321,N_5072);
and U6316 (N_6316,N_5527,N_5019);
and U6317 (N_6317,N_5556,N_5714);
and U6318 (N_6318,N_5869,N_5880);
and U6319 (N_6319,N_5022,N_5231);
nand U6320 (N_6320,N_5543,N_5103);
and U6321 (N_6321,N_5111,N_5937);
or U6322 (N_6322,N_5941,N_5612);
nor U6323 (N_6323,N_5785,N_5352);
or U6324 (N_6324,N_5911,N_5804);
nor U6325 (N_6325,N_5695,N_5787);
nand U6326 (N_6326,N_5754,N_5418);
or U6327 (N_6327,N_5253,N_5901);
nor U6328 (N_6328,N_5734,N_5685);
or U6329 (N_6329,N_5701,N_5270);
and U6330 (N_6330,N_5589,N_5423);
or U6331 (N_6331,N_5759,N_5919);
nor U6332 (N_6332,N_5258,N_5574);
and U6333 (N_6333,N_5046,N_5960);
nor U6334 (N_6334,N_5756,N_5305);
or U6335 (N_6335,N_5236,N_5288);
or U6336 (N_6336,N_5286,N_5883);
and U6337 (N_6337,N_5765,N_5174);
and U6338 (N_6338,N_5181,N_5811);
nand U6339 (N_6339,N_5697,N_5531);
nand U6340 (N_6340,N_5339,N_5786);
or U6341 (N_6341,N_5425,N_5670);
or U6342 (N_6342,N_5625,N_5696);
and U6343 (N_6343,N_5644,N_5155);
and U6344 (N_6344,N_5041,N_5773);
nand U6345 (N_6345,N_5806,N_5239);
and U6346 (N_6346,N_5237,N_5264);
nor U6347 (N_6347,N_5568,N_5455);
or U6348 (N_6348,N_5017,N_5912);
nor U6349 (N_6349,N_5692,N_5276);
or U6350 (N_6350,N_5509,N_5877);
nand U6351 (N_6351,N_5820,N_5370);
or U6352 (N_6352,N_5822,N_5089);
nand U6353 (N_6353,N_5107,N_5728);
nand U6354 (N_6354,N_5851,N_5634);
or U6355 (N_6355,N_5723,N_5227);
and U6356 (N_6356,N_5529,N_5602);
and U6357 (N_6357,N_5159,N_5271);
nor U6358 (N_6358,N_5075,N_5131);
nand U6359 (N_6359,N_5203,N_5377);
nand U6360 (N_6360,N_5038,N_5586);
nor U6361 (N_6361,N_5389,N_5133);
nor U6362 (N_6362,N_5745,N_5571);
nor U6363 (N_6363,N_5827,N_5408);
or U6364 (N_6364,N_5590,N_5282);
nor U6365 (N_6365,N_5861,N_5393);
and U6366 (N_6366,N_5992,N_5252);
or U6367 (N_6367,N_5542,N_5010);
or U6368 (N_6368,N_5487,N_5943);
or U6369 (N_6369,N_5730,N_5442);
nand U6370 (N_6370,N_5495,N_5797);
or U6371 (N_6371,N_5275,N_5622);
and U6372 (N_6372,N_5505,N_5287);
and U6373 (N_6373,N_5708,N_5921);
and U6374 (N_6374,N_5550,N_5768);
xnor U6375 (N_6375,N_5788,N_5397);
nor U6376 (N_6376,N_5626,N_5003);
nand U6377 (N_6377,N_5779,N_5061);
xor U6378 (N_6378,N_5453,N_5617);
nand U6379 (N_6379,N_5093,N_5438);
and U6380 (N_6380,N_5936,N_5751);
or U6381 (N_6381,N_5272,N_5141);
or U6382 (N_6382,N_5417,N_5973);
or U6383 (N_6383,N_5715,N_5363);
nor U6384 (N_6384,N_5769,N_5066);
and U6385 (N_6385,N_5640,N_5036);
or U6386 (N_6386,N_5020,N_5944);
nor U6387 (N_6387,N_5268,N_5201);
nand U6388 (N_6388,N_5211,N_5536);
and U6389 (N_6389,N_5842,N_5083);
nor U6390 (N_6390,N_5396,N_5572);
or U6391 (N_6391,N_5721,N_5835);
and U6392 (N_6392,N_5382,N_5292);
xor U6393 (N_6393,N_5559,N_5952);
nand U6394 (N_6394,N_5979,N_5791);
nand U6395 (N_6395,N_5360,N_5870);
nand U6396 (N_6396,N_5829,N_5927);
or U6397 (N_6397,N_5682,N_5474);
nor U6398 (N_6398,N_5444,N_5818);
nor U6399 (N_6399,N_5109,N_5387);
nor U6400 (N_6400,N_5918,N_5523);
nand U6401 (N_6401,N_5777,N_5183);
and U6402 (N_6402,N_5309,N_5050);
nor U6403 (N_6403,N_5401,N_5371);
or U6404 (N_6404,N_5700,N_5433);
or U6405 (N_6405,N_5054,N_5552);
nand U6406 (N_6406,N_5596,N_5908);
and U6407 (N_6407,N_5357,N_5679);
nor U6408 (N_6408,N_5477,N_5285);
nor U6409 (N_6409,N_5711,N_5151);
and U6410 (N_6410,N_5324,N_5621);
and U6411 (N_6411,N_5736,N_5266);
and U6412 (N_6412,N_5063,N_5429);
and U6413 (N_6413,N_5860,N_5780);
nor U6414 (N_6414,N_5219,N_5323);
nand U6415 (N_6415,N_5743,N_5121);
nor U6416 (N_6416,N_5814,N_5037);
or U6417 (N_6417,N_5698,N_5994);
nand U6418 (N_6418,N_5049,N_5643);
nand U6419 (N_6419,N_5233,N_5030);
nand U6420 (N_6420,N_5014,N_5789);
nor U6421 (N_6421,N_5008,N_5859);
and U6422 (N_6422,N_5104,N_5031);
nor U6423 (N_6423,N_5850,N_5378);
nand U6424 (N_6424,N_5398,N_5499);
and U6425 (N_6425,N_5376,N_5021);
and U6426 (N_6426,N_5097,N_5293);
and U6427 (N_6427,N_5163,N_5255);
and U6428 (N_6428,N_5294,N_5426);
nor U6429 (N_6429,N_5295,N_5757);
nand U6430 (N_6430,N_5849,N_5334);
nor U6431 (N_6431,N_5485,N_5470);
nand U6432 (N_6432,N_5217,N_5573);
or U6433 (N_6433,N_5446,N_5515);
and U6434 (N_6434,N_5998,N_5857);
nand U6435 (N_6435,N_5597,N_5910);
nor U6436 (N_6436,N_5079,N_5595);
or U6437 (N_6437,N_5077,N_5238);
and U6438 (N_6438,N_5663,N_5172);
and U6439 (N_6439,N_5144,N_5205);
and U6440 (N_6440,N_5848,N_5195);
and U6441 (N_6441,N_5394,N_5500);
nand U6442 (N_6442,N_5065,N_5637);
nor U6443 (N_6443,N_5345,N_5431);
or U6444 (N_6444,N_5188,N_5187);
nand U6445 (N_6445,N_5868,N_5226);
nor U6446 (N_6446,N_5554,N_5404);
nand U6447 (N_6447,N_5454,N_5798);
nand U6448 (N_6448,N_5381,N_5852);
or U6449 (N_6449,N_5645,N_5135);
nor U6450 (N_6450,N_5654,N_5331);
or U6451 (N_6451,N_5946,N_5090);
or U6452 (N_6452,N_5915,N_5439);
nand U6453 (N_6453,N_5186,N_5399);
nand U6454 (N_6454,N_5538,N_5752);
nand U6455 (N_6455,N_5591,N_5824);
nand U6456 (N_6456,N_5094,N_5557);
or U6457 (N_6457,N_5511,N_5248);
nand U6458 (N_6458,N_5348,N_5956);
or U6459 (N_6459,N_5194,N_5732);
xnor U6460 (N_6460,N_5502,N_5838);
nand U6461 (N_6461,N_5307,N_5379);
and U6462 (N_6462,N_5136,N_5642);
or U6463 (N_6463,N_5793,N_5719);
nand U6464 (N_6464,N_5738,N_5893);
or U6465 (N_6465,N_5043,N_5776);
or U6466 (N_6466,N_5971,N_5447);
or U6467 (N_6467,N_5434,N_5071);
nand U6468 (N_6468,N_5007,N_5705);
nor U6469 (N_6469,N_5710,N_5406);
and U6470 (N_6470,N_5462,N_5727);
or U6471 (N_6471,N_5388,N_5983);
nor U6472 (N_6472,N_5917,N_5445);
or U6473 (N_6473,N_5873,N_5825);
and U6474 (N_6474,N_5693,N_5225);
and U6475 (N_6475,N_5553,N_5616);
xor U6476 (N_6476,N_5437,N_5481);
or U6477 (N_6477,N_5464,N_5059);
nand U6478 (N_6478,N_5831,N_5358);
or U6479 (N_6479,N_5230,N_5099);
or U6480 (N_6480,N_5261,N_5145);
nand U6481 (N_6481,N_5409,N_5273);
nand U6482 (N_6482,N_5142,N_5801);
nand U6483 (N_6483,N_5052,N_5691);
and U6484 (N_6484,N_5583,N_5105);
nand U6485 (N_6485,N_5006,N_5884);
or U6486 (N_6486,N_5407,N_5673);
and U6487 (N_6487,N_5196,N_5146);
or U6488 (N_6488,N_5996,N_5980);
or U6489 (N_6489,N_5108,N_5628);
and U6490 (N_6490,N_5607,N_5795);
nor U6491 (N_6491,N_5817,N_5355);
nor U6492 (N_6492,N_5862,N_5900);
or U6493 (N_6493,N_5819,N_5664);
and U6494 (N_6494,N_5449,N_5748);
and U6495 (N_6495,N_5478,N_5774);
or U6496 (N_6496,N_5904,N_5269);
and U6497 (N_6497,N_5420,N_5042);
or U6498 (N_6498,N_5967,N_5311);
nor U6499 (N_6499,N_5903,N_5548);
nor U6500 (N_6500,N_5064,N_5292);
and U6501 (N_6501,N_5126,N_5474);
or U6502 (N_6502,N_5339,N_5883);
and U6503 (N_6503,N_5005,N_5754);
and U6504 (N_6504,N_5520,N_5467);
or U6505 (N_6505,N_5888,N_5955);
or U6506 (N_6506,N_5254,N_5842);
nor U6507 (N_6507,N_5603,N_5587);
and U6508 (N_6508,N_5277,N_5485);
and U6509 (N_6509,N_5383,N_5640);
nand U6510 (N_6510,N_5580,N_5672);
nand U6511 (N_6511,N_5582,N_5515);
and U6512 (N_6512,N_5034,N_5700);
or U6513 (N_6513,N_5658,N_5409);
and U6514 (N_6514,N_5582,N_5872);
or U6515 (N_6515,N_5106,N_5335);
or U6516 (N_6516,N_5429,N_5038);
or U6517 (N_6517,N_5354,N_5876);
and U6518 (N_6518,N_5807,N_5924);
nor U6519 (N_6519,N_5218,N_5324);
nand U6520 (N_6520,N_5526,N_5489);
and U6521 (N_6521,N_5634,N_5783);
or U6522 (N_6522,N_5486,N_5736);
or U6523 (N_6523,N_5558,N_5024);
or U6524 (N_6524,N_5151,N_5956);
or U6525 (N_6525,N_5475,N_5091);
and U6526 (N_6526,N_5399,N_5322);
and U6527 (N_6527,N_5619,N_5125);
xor U6528 (N_6528,N_5916,N_5944);
nand U6529 (N_6529,N_5177,N_5857);
and U6530 (N_6530,N_5707,N_5427);
or U6531 (N_6531,N_5313,N_5865);
nand U6532 (N_6532,N_5647,N_5048);
and U6533 (N_6533,N_5322,N_5186);
or U6534 (N_6534,N_5170,N_5897);
and U6535 (N_6535,N_5085,N_5666);
or U6536 (N_6536,N_5130,N_5912);
nor U6537 (N_6537,N_5941,N_5446);
nand U6538 (N_6538,N_5520,N_5371);
nor U6539 (N_6539,N_5543,N_5511);
nor U6540 (N_6540,N_5946,N_5278);
nand U6541 (N_6541,N_5002,N_5849);
or U6542 (N_6542,N_5191,N_5937);
nand U6543 (N_6543,N_5077,N_5632);
and U6544 (N_6544,N_5924,N_5203);
or U6545 (N_6545,N_5611,N_5495);
or U6546 (N_6546,N_5894,N_5889);
and U6547 (N_6547,N_5698,N_5028);
nor U6548 (N_6548,N_5598,N_5286);
and U6549 (N_6549,N_5091,N_5632);
nor U6550 (N_6550,N_5760,N_5813);
nand U6551 (N_6551,N_5531,N_5514);
and U6552 (N_6552,N_5010,N_5848);
nor U6553 (N_6553,N_5918,N_5382);
nand U6554 (N_6554,N_5527,N_5272);
or U6555 (N_6555,N_5834,N_5290);
nor U6556 (N_6556,N_5677,N_5814);
nand U6557 (N_6557,N_5990,N_5402);
and U6558 (N_6558,N_5665,N_5259);
nand U6559 (N_6559,N_5260,N_5804);
nand U6560 (N_6560,N_5050,N_5731);
nor U6561 (N_6561,N_5207,N_5587);
nand U6562 (N_6562,N_5141,N_5348);
or U6563 (N_6563,N_5569,N_5492);
and U6564 (N_6564,N_5122,N_5495);
nand U6565 (N_6565,N_5123,N_5446);
nor U6566 (N_6566,N_5822,N_5759);
or U6567 (N_6567,N_5235,N_5933);
nand U6568 (N_6568,N_5519,N_5810);
or U6569 (N_6569,N_5942,N_5229);
and U6570 (N_6570,N_5527,N_5991);
or U6571 (N_6571,N_5752,N_5879);
or U6572 (N_6572,N_5594,N_5345);
nand U6573 (N_6573,N_5880,N_5550);
or U6574 (N_6574,N_5787,N_5289);
and U6575 (N_6575,N_5183,N_5372);
and U6576 (N_6576,N_5779,N_5485);
nor U6577 (N_6577,N_5504,N_5429);
nor U6578 (N_6578,N_5242,N_5160);
nand U6579 (N_6579,N_5827,N_5422);
and U6580 (N_6580,N_5063,N_5846);
nand U6581 (N_6581,N_5408,N_5775);
nor U6582 (N_6582,N_5425,N_5997);
nor U6583 (N_6583,N_5282,N_5131);
nor U6584 (N_6584,N_5490,N_5886);
nand U6585 (N_6585,N_5667,N_5434);
or U6586 (N_6586,N_5896,N_5548);
nor U6587 (N_6587,N_5540,N_5682);
nor U6588 (N_6588,N_5814,N_5034);
nand U6589 (N_6589,N_5057,N_5787);
nand U6590 (N_6590,N_5097,N_5083);
nor U6591 (N_6591,N_5437,N_5358);
nand U6592 (N_6592,N_5623,N_5176);
nor U6593 (N_6593,N_5341,N_5206);
nand U6594 (N_6594,N_5244,N_5072);
nor U6595 (N_6595,N_5063,N_5457);
nor U6596 (N_6596,N_5675,N_5186);
and U6597 (N_6597,N_5741,N_5086);
xor U6598 (N_6598,N_5181,N_5322);
and U6599 (N_6599,N_5385,N_5005);
and U6600 (N_6600,N_5908,N_5157);
or U6601 (N_6601,N_5771,N_5960);
nor U6602 (N_6602,N_5002,N_5587);
nand U6603 (N_6603,N_5619,N_5717);
and U6604 (N_6604,N_5579,N_5928);
nand U6605 (N_6605,N_5651,N_5185);
nand U6606 (N_6606,N_5209,N_5689);
nand U6607 (N_6607,N_5432,N_5864);
nor U6608 (N_6608,N_5033,N_5821);
and U6609 (N_6609,N_5515,N_5887);
nand U6610 (N_6610,N_5036,N_5167);
nand U6611 (N_6611,N_5806,N_5197);
nand U6612 (N_6612,N_5117,N_5894);
and U6613 (N_6613,N_5337,N_5059);
nand U6614 (N_6614,N_5524,N_5958);
or U6615 (N_6615,N_5489,N_5399);
or U6616 (N_6616,N_5242,N_5944);
and U6617 (N_6617,N_5135,N_5410);
and U6618 (N_6618,N_5425,N_5873);
nor U6619 (N_6619,N_5275,N_5335);
xor U6620 (N_6620,N_5634,N_5007);
and U6621 (N_6621,N_5260,N_5074);
and U6622 (N_6622,N_5636,N_5680);
or U6623 (N_6623,N_5886,N_5321);
nor U6624 (N_6624,N_5801,N_5591);
and U6625 (N_6625,N_5933,N_5748);
and U6626 (N_6626,N_5906,N_5907);
nor U6627 (N_6627,N_5550,N_5970);
nand U6628 (N_6628,N_5174,N_5537);
and U6629 (N_6629,N_5760,N_5117);
nand U6630 (N_6630,N_5160,N_5985);
nand U6631 (N_6631,N_5885,N_5864);
or U6632 (N_6632,N_5846,N_5612);
nand U6633 (N_6633,N_5654,N_5987);
and U6634 (N_6634,N_5853,N_5906);
or U6635 (N_6635,N_5777,N_5733);
and U6636 (N_6636,N_5002,N_5468);
nor U6637 (N_6637,N_5788,N_5210);
nand U6638 (N_6638,N_5505,N_5040);
or U6639 (N_6639,N_5108,N_5409);
or U6640 (N_6640,N_5027,N_5139);
and U6641 (N_6641,N_5334,N_5578);
nand U6642 (N_6642,N_5522,N_5494);
nand U6643 (N_6643,N_5389,N_5884);
nand U6644 (N_6644,N_5156,N_5072);
nor U6645 (N_6645,N_5828,N_5841);
or U6646 (N_6646,N_5679,N_5719);
or U6647 (N_6647,N_5327,N_5697);
nand U6648 (N_6648,N_5191,N_5751);
and U6649 (N_6649,N_5883,N_5560);
nor U6650 (N_6650,N_5680,N_5206);
or U6651 (N_6651,N_5382,N_5594);
and U6652 (N_6652,N_5675,N_5170);
or U6653 (N_6653,N_5502,N_5836);
nor U6654 (N_6654,N_5912,N_5722);
nand U6655 (N_6655,N_5988,N_5507);
nand U6656 (N_6656,N_5867,N_5253);
and U6657 (N_6657,N_5909,N_5542);
and U6658 (N_6658,N_5349,N_5686);
and U6659 (N_6659,N_5505,N_5639);
and U6660 (N_6660,N_5000,N_5165);
and U6661 (N_6661,N_5485,N_5460);
nor U6662 (N_6662,N_5774,N_5949);
or U6663 (N_6663,N_5597,N_5566);
nand U6664 (N_6664,N_5446,N_5859);
nand U6665 (N_6665,N_5062,N_5919);
nor U6666 (N_6666,N_5269,N_5241);
nor U6667 (N_6667,N_5129,N_5613);
xor U6668 (N_6668,N_5907,N_5202);
and U6669 (N_6669,N_5064,N_5937);
or U6670 (N_6670,N_5692,N_5070);
and U6671 (N_6671,N_5277,N_5063);
xor U6672 (N_6672,N_5616,N_5169);
and U6673 (N_6673,N_5821,N_5976);
nand U6674 (N_6674,N_5758,N_5803);
and U6675 (N_6675,N_5566,N_5264);
or U6676 (N_6676,N_5856,N_5988);
nor U6677 (N_6677,N_5487,N_5318);
nor U6678 (N_6678,N_5219,N_5734);
and U6679 (N_6679,N_5624,N_5058);
and U6680 (N_6680,N_5231,N_5265);
or U6681 (N_6681,N_5165,N_5228);
and U6682 (N_6682,N_5839,N_5512);
nand U6683 (N_6683,N_5285,N_5620);
xor U6684 (N_6684,N_5773,N_5983);
and U6685 (N_6685,N_5429,N_5678);
or U6686 (N_6686,N_5084,N_5368);
nand U6687 (N_6687,N_5828,N_5135);
nor U6688 (N_6688,N_5806,N_5817);
nand U6689 (N_6689,N_5804,N_5232);
and U6690 (N_6690,N_5068,N_5189);
nor U6691 (N_6691,N_5025,N_5792);
nor U6692 (N_6692,N_5337,N_5285);
nor U6693 (N_6693,N_5140,N_5168);
nand U6694 (N_6694,N_5944,N_5926);
nand U6695 (N_6695,N_5473,N_5696);
nand U6696 (N_6696,N_5623,N_5808);
nor U6697 (N_6697,N_5320,N_5682);
or U6698 (N_6698,N_5243,N_5902);
and U6699 (N_6699,N_5269,N_5534);
or U6700 (N_6700,N_5386,N_5179);
nand U6701 (N_6701,N_5552,N_5775);
and U6702 (N_6702,N_5092,N_5973);
nor U6703 (N_6703,N_5757,N_5656);
nor U6704 (N_6704,N_5035,N_5406);
nand U6705 (N_6705,N_5634,N_5559);
or U6706 (N_6706,N_5110,N_5185);
nand U6707 (N_6707,N_5744,N_5736);
or U6708 (N_6708,N_5328,N_5628);
and U6709 (N_6709,N_5632,N_5059);
nor U6710 (N_6710,N_5727,N_5782);
nor U6711 (N_6711,N_5933,N_5095);
nor U6712 (N_6712,N_5918,N_5771);
nor U6713 (N_6713,N_5729,N_5697);
or U6714 (N_6714,N_5810,N_5376);
or U6715 (N_6715,N_5504,N_5164);
and U6716 (N_6716,N_5043,N_5981);
nor U6717 (N_6717,N_5983,N_5219);
or U6718 (N_6718,N_5666,N_5529);
and U6719 (N_6719,N_5861,N_5638);
or U6720 (N_6720,N_5399,N_5926);
nor U6721 (N_6721,N_5693,N_5912);
and U6722 (N_6722,N_5176,N_5403);
or U6723 (N_6723,N_5078,N_5565);
nand U6724 (N_6724,N_5979,N_5439);
nor U6725 (N_6725,N_5091,N_5603);
nand U6726 (N_6726,N_5114,N_5207);
nand U6727 (N_6727,N_5079,N_5504);
nor U6728 (N_6728,N_5281,N_5982);
nand U6729 (N_6729,N_5960,N_5655);
nand U6730 (N_6730,N_5253,N_5910);
nor U6731 (N_6731,N_5048,N_5440);
nand U6732 (N_6732,N_5266,N_5024);
and U6733 (N_6733,N_5704,N_5640);
and U6734 (N_6734,N_5085,N_5863);
nand U6735 (N_6735,N_5303,N_5445);
xor U6736 (N_6736,N_5720,N_5132);
or U6737 (N_6737,N_5591,N_5884);
or U6738 (N_6738,N_5275,N_5492);
nand U6739 (N_6739,N_5767,N_5251);
nor U6740 (N_6740,N_5625,N_5894);
nor U6741 (N_6741,N_5478,N_5762);
and U6742 (N_6742,N_5357,N_5664);
or U6743 (N_6743,N_5769,N_5084);
and U6744 (N_6744,N_5308,N_5857);
or U6745 (N_6745,N_5640,N_5115);
nand U6746 (N_6746,N_5331,N_5032);
or U6747 (N_6747,N_5296,N_5355);
nor U6748 (N_6748,N_5196,N_5062);
nand U6749 (N_6749,N_5682,N_5600);
nor U6750 (N_6750,N_5138,N_5701);
nand U6751 (N_6751,N_5656,N_5908);
or U6752 (N_6752,N_5821,N_5241);
or U6753 (N_6753,N_5341,N_5403);
or U6754 (N_6754,N_5250,N_5471);
nand U6755 (N_6755,N_5507,N_5728);
or U6756 (N_6756,N_5684,N_5739);
or U6757 (N_6757,N_5955,N_5527);
nand U6758 (N_6758,N_5227,N_5196);
nand U6759 (N_6759,N_5675,N_5451);
nor U6760 (N_6760,N_5278,N_5493);
nand U6761 (N_6761,N_5543,N_5721);
and U6762 (N_6762,N_5066,N_5503);
and U6763 (N_6763,N_5138,N_5357);
nor U6764 (N_6764,N_5091,N_5097);
nand U6765 (N_6765,N_5847,N_5171);
nor U6766 (N_6766,N_5018,N_5139);
and U6767 (N_6767,N_5554,N_5652);
or U6768 (N_6768,N_5664,N_5651);
or U6769 (N_6769,N_5166,N_5431);
nor U6770 (N_6770,N_5017,N_5233);
nor U6771 (N_6771,N_5320,N_5498);
nand U6772 (N_6772,N_5972,N_5996);
or U6773 (N_6773,N_5296,N_5903);
or U6774 (N_6774,N_5968,N_5267);
nor U6775 (N_6775,N_5563,N_5784);
nor U6776 (N_6776,N_5714,N_5577);
nor U6777 (N_6777,N_5887,N_5952);
and U6778 (N_6778,N_5041,N_5309);
nand U6779 (N_6779,N_5293,N_5203);
and U6780 (N_6780,N_5105,N_5940);
nand U6781 (N_6781,N_5183,N_5319);
or U6782 (N_6782,N_5750,N_5509);
or U6783 (N_6783,N_5843,N_5572);
or U6784 (N_6784,N_5997,N_5972);
or U6785 (N_6785,N_5033,N_5999);
xor U6786 (N_6786,N_5059,N_5812);
nor U6787 (N_6787,N_5110,N_5512);
and U6788 (N_6788,N_5112,N_5471);
nand U6789 (N_6789,N_5269,N_5184);
and U6790 (N_6790,N_5209,N_5238);
nand U6791 (N_6791,N_5613,N_5546);
nor U6792 (N_6792,N_5544,N_5225);
nand U6793 (N_6793,N_5007,N_5621);
or U6794 (N_6794,N_5544,N_5628);
nand U6795 (N_6795,N_5351,N_5111);
nor U6796 (N_6796,N_5175,N_5869);
and U6797 (N_6797,N_5876,N_5047);
or U6798 (N_6798,N_5243,N_5366);
and U6799 (N_6799,N_5146,N_5252);
nand U6800 (N_6800,N_5366,N_5302);
nand U6801 (N_6801,N_5587,N_5024);
nor U6802 (N_6802,N_5029,N_5577);
nand U6803 (N_6803,N_5618,N_5382);
or U6804 (N_6804,N_5147,N_5961);
or U6805 (N_6805,N_5820,N_5243);
xnor U6806 (N_6806,N_5708,N_5809);
nand U6807 (N_6807,N_5505,N_5870);
or U6808 (N_6808,N_5148,N_5378);
nor U6809 (N_6809,N_5365,N_5843);
nand U6810 (N_6810,N_5080,N_5316);
nor U6811 (N_6811,N_5329,N_5619);
and U6812 (N_6812,N_5710,N_5781);
nand U6813 (N_6813,N_5253,N_5970);
and U6814 (N_6814,N_5678,N_5424);
nor U6815 (N_6815,N_5598,N_5740);
nand U6816 (N_6816,N_5771,N_5273);
nor U6817 (N_6817,N_5990,N_5377);
nand U6818 (N_6818,N_5557,N_5276);
and U6819 (N_6819,N_5487,N_5645);
nand U6820 (N_6820,N_5835,N_5333);
or U6821 (N_6821,N_5235,N_5106);
nor U6822 (N_6822,N_5164,N_5917);
and U6823 (N_6823,N_5747,N_5671);
and U6824 (N_6824,N_5648,N_5504);
nor U6825 (N_6825,N_5448,N_5849);
or U6826 (N_6826,N_5640,N_5736);
and U6827 (N_6827,N_5607,N_5071);
or U6828 (N_6828,N_5466,N_5006);
nor U6829 (N_6829,N_5852,N_5140);
nand U6830 (N_6830,N_5199,N_5346);
nand U6831 (N_6831,N_5358,N_5544);
nor U6832 (N_6832,N_5795,N_5210);
nor U6833 (N_6833,N_5303,N_5160);
or U6834 (N_6834,N_5668,N_5630);
and U6835 (N_6835,N_5415,N_5500);
and U6836 (N_6836,N_5610,N_5051);
nor U6837 (N_6837,N_5377,N_5936);
and U6838 (N_6838,N_5891,N_5027);
and U6839 (N_6839,N_5128,N_5221);
or U6840 (N_6840,N_5817,N_5426);
nand U6841 (N_6841,N_5116,N_5596);
nor U6842 (N_6842,N_5291,N_5379);
or U6843 (N_6843,N_5310,N_5782);
or U6844 (N_6844,N_5717,N_5352);
nand U6845 (N_6845,N_5181,N_5491);
and U6846 (N_6846,N_5220,N_5621);
or U6847 (N_6847,N_5864,N_5418);
and U6848 (N_6848,N_5330,N_5238);
nand U6849 (N_6849,N_5548,N_5053);
nand U6850 (N_6850,N_5499,N_5472);
and U6851 (N_6851,N_5717,N_5858);
nand U6852 (N_6852,N_5146,N_5391);
nand U6853 (N_6853,N_5363,N_5948);
or U6854 (N_6854,N_5963,N_5393);
nand U6855 (N_6855,N_5215,N_5898);
nor U6856 (N_6856,N_5292,N_5582);
or U6857 (N_6857,N_5880,N_5299);
nor U6858 (N_6858,N_5727,N_5670);
or U6859 (N_6859,N_5431,N_5747);
nand U6860 (N_6860,N_5228,N_5520);
and U6861 (N_6861,N_5449,N_5239);
and U6862 (N_6862,N_5164,N_5831);
and U6863 (N_6863,N_5210,N_5196);
nand U6864 (N_6864,N_5900,N_5430);
or U6865 (N_6865,N_5923,N_5403);
xnor U6866 (N_6866,N_5997,N_5179);
or U6867 (N_6867,N_5199,N_5420);
nand U6868 (N_6868,N_5517,N_5834);
and U6869 (N_6869,N_5836,N_5443);
nand U6870 (N_6870,N_5967,N_5480);
nor U6871 (N_6871,N_5975,N_5808);
and U6872 (N_6872,N_5300,N_5976);
nand U6873 (N_6873,N_5959,N_5575);
nor U6874 (N_6874,N_5261,N_5175);
or U6875 (N_6875,N_5609,N_5070);
or U6876 (N_6876,N_5074,N_5443);
and U6877 (N_6877,N_5102,N_5719);
and U6878 (N_6878,N_5464,N_5762);
or U6879 (N_6879,N_5937,N_5205);
nor U6880 (N_6880,N_5333,N_5780);
xor U6881 (N_6881,N_5700,N_5537);
or U6882 (N_6882,N_5922,N_5519);
nand U6883 (N_6883,N_5457,N_5450);
or U6884 (N_6884,N_5303,N_5677);
nand U6885 (N_6885,N_5496,N_5338);
and U6886 (N_6886,N_5927,N_5130);
nor U6887 (N_6887,N_5894,N_5291);
and U6888 (N_6888,N_5946,N_5448);
or U6889 (N_6889,N_5078,N_5101);
nor U6890 (N_6890,N_5963,N_5639);
or U6891 (N_6891,N_5329,N_5799);
or U6892 (N_6892,N_5757,N_5671);
nor U6893 (N_6893,N_5658,N_5253);
nor U6894 (N_6894,N_5485,N_5015);
and U6895 (N_6895,N_5823,N_5959);
nor U6896 (N_6896,N_5723,N_5607);
nand U6897 (N_6897,N_5955,N_5819);
nand U6898 (N_6898,N_5878,N_5489);
and U6899 (N_6899,N_5285,N_5968);
or U6900 (N_6900,N_5975,N_5465);
or U6901 (N_6901,N_5371,N_5448);
and U6902 (N_6902,N_5585,N_5494);
or U6903 (N_6903,N_5395,N_5616);
nor U6904 (N_6904,N_5923,N_5119);
nand U6905 (N_6905,N_5427,N_5661);
or U6906 (N_6906,N_5595,N_5594);
and U6907 (N_6907,N_5974,N_5289);
nor U6908 (N_6908,N_5533,N_5444);
nand U6909 (N_6909,N_5506,N_5019);
nand U6910 (N_6910,N_5345,N_5619);
nand U6911 (N_6911,N_5839,N_5709);
nor U6912 (N_6912,N_5074,N_5152);
nor U6913 (N_6913,N_5864,N_5142);
nand U6914 (N_6914,N_5793,N_5256);
and U6915 (N_6915,N_5924,N_5569);
or U6916 (N_6916,N_5978,N_5075);
nand U6917 (N_6917,N_5346,N_5832);
or U6918 (N_6918,N_5828,N_5770);
and U6919 (N_6919,N_5193,N_5297);
nor U6920 (N_6920,N_5536,N_5720);
or U6921 (N_6921,N_5696,N_5828);
and U6922 (N_6922,N_5859,N_5306);
and U6923 (N_6923,N_5969,N_5663);
nand U6924 (N_6924,N_5173,N_5737);
nand U6925 (N_6925,N_5686,N_5848);
and U6926 (N_6926,N_5793,N_5589);
nand U6927 (N_6927,N_5626,N_5922);
nand U6928 (N_6928,N_5332,N_5265);
and U6929 (N_6929,N_5607,N_5263);
and U6930 (N_6930,N_5131,N_5624);
and U6931 (N_6931,N_5910,N_5239);
or U6932 (N_6932,N_5533,N_5329);
and U6933 (N_6933,N_5826,N_5218);
and U6934 (N_6934,N_5767,N_5141);
nor U6935 (N_6935,N_5935,N_5470);
nor U6936 (N_6936,N_5123,N_5241);
or U6937 (N_6937,N_5439,N_5735);
nand U6938 (N_6938,N_5499,N_5578);
and U6939 (N_6939,N_5388,N_5541);
nor U6940 (N_6940,N_5629,N_5600);
or U6941 (N_6941,N_5450,N_5080);
nor U6942 (N_6942,N_5920,N_5585);
nor U6943 (N_6943,N_5819,N_5061);
or U6944 (N_6944,N_5147,N_5985);
nand U6945 (N_6945,N_5484,N_5273);
and U6946 (N_6946,N_5221,N_5474);
and U6947 (N_6947,N_5755,N_5117);
nand U6948 (N_6948,N_5287,N_5369);
nand U6949 (N_6949,N_5238,N_5220);
nand U6950 (N_6950,N_5240,N_5418);
or U6951 (N_6951,N_5076,N_5890);
nor U6952 (N_6952,N_5250,N_5115);
or U6953 (N_6953,N_5379,N_5942);
nor U6954 (N_6954,N_5086,N_5647);
and U6955 (N_6955,N_5384,N_5912);
nand U6956 (N_6956,N_5339,N_5845);
nand U6957 (N_6957,N_5900,N_5200);
nand U6958 (N_6958,N_5421,N_5259);
nor U6959 (N_6959,N_5016,N_5235);
or U6960 (N_6960,N_5752,N_5313);
nor U6961 (N_6961,N_5320,N_5779);
nand U6962 (N_6962,N_5112,N_5948);
nand U6963 (N_6963,N_5877,N_5889);
nor U6964 (N_6964,N_5802,N_5036);
and U6965 (N_6965,N_5425,N_5765);
nor U6966 (N_6966,N_5649,N_5403);
nand U6967 (N_6967,N_5253,N_5782);
nand U6968 (N_6968,N_5268,N_5212);
or U6969 (N_6969,N_5316,N_5077);
and U6970 (N_6970,N_5081,N_5121);
nor U6971 (N_6971,N_5259,N_5662);
nor U6972 (N_6972,N_5810,N_5391);
nor U6973 (N_6973,N_5313,N_5104);
nand U6974 (N_6974,N_5537,N_5023);
or U6975 (N_6975,N_5756,N_5699);
or U6976 (N_6976,N_5974,N_5848);
or U6977 (N_6977,N_5586,N_5984);
nand U6978 (N_6978,N_5077,N_5225);
or U6979 (N_6979,N_5852,N_5911);
or U6980 (N_6980,N_5243,N_5259);
and U6981 (N_6981,N_5719,N_5081);
nand U6982 (N_6982,N_5233,N_5289);
and U6983 (N_6983,N_5248,N_5206);
and U6984 (N_6984,N_5762,N_5417);
or U6985 (N_6985,N_5015,N_5543);
or U6986 (N_6986,N_5764,N_5091);
nor U6987 (N_6987,N_5504,N_5755);
nand U6988 (N_6988,N_5715,N_5530);
xor U6989 (N_6989,N_5578,N_5183);
nand U6990 (N_6990,N_5192,N_5968);
or U6991 (N_6991,N_5869,N_5186);
or U6992 (N_6992,N_5745,N_5057);
nand U6993 (N_6993,N_5575,N_5558);
and U6994 (N_6994,N_5553,N_5861);
nand U6995 (N_6995,N_5579,N_5369);
and U6996 (N_6996,N_5887,N_5221);
and U6997 (N_6997,N_5226,N_5832);
nand U6998 (N_6998,N_5027,N_5349);
nand U6999 (N_6999,N_5041,N_5267);
nand U7000 (N_7000,N_6765,N_6198);
or U7001 (N_7001,N_6527,N_6111);
or U7002 (N_7002,N_6698,N_6138);
and U7003 (N_7003,N_6122,N_6908);
and U7004 (N_7004,N_6174,N_6975);
nand U7005 (N_7005,N_6465,N_6075);
or U7006 (N_7006,N_6031,N_6312);
or U7007 (N_7007,N_6674,N_6385);
and U7008 (N_7008,N_6723,N_6616);
nor U7009 (N_7009,N_6080,N_6968);
or U7010 (N_7010,N_6981,N_6913);
or U7011 (N_7011,N_6850,N_6023);
and U7012 (N_7012,N_6733,N_6716);
nand U7013 (N_7013,N_6855,N_6758);
nor U7014 (N_7014,N_6669,N_6889);
nor U7015 (N_7015,N_6757,N_6335);
or U7016 (N_7016,N_6717,N_6433);
and U7017 (N_7017,N_6618,N_6297);
and U7018 (N_7018,N_6989,N_6180);
or U7019 (N_7019,N_6193,N_6918);
nor U7020 (N_7020,N_6957,N_6689);
or U7021 (N_7021,N_6597,N_6730);
or U7022 (N_7022,N_6208,N_6960);
and U7023 (N_7023,N_6523,N_6234);
or U7024 (N_7024,N_6721,N_6376);
and U7025 (N_7025,N_6500,N_6749);
nor U7026 (N_7026,N_6593,N_6298);
nor U7027 (N_7027,N_6836,N_6192);
and U7028 (N_7028,N_6492,N_6745);
and U7029 (N_7029,N_6648,N_6403);
or U7030 (N_7030,N_6411,N_6040);
and U7031 (N_7031,N_6476,N_6951);
or U7032 (N_7032,N_6853,N_6175);
or U7033 (N_7033,N_6501,N_6947);
nor U7034 (N_7034,N_6462,N_6787);
nor U7035 (N_7035,N_6191,N_6041);
nor U7036 (N_7036,N_6553,N_6676);
and U7037 (N_7037,N_6109,N_6296);
or U7038 (N_7038,N_6228,N_6469);
and U7039 (N_7039,N_6262,N_6466);
nor U7040 (N_7040,N_6242,N_6516);
nor U7041 (N_7041,N_6678,N_6359);
nand U7042 (N_7042,N_6604,N_6831);
or U7043 (N_7043,N_6961,N_6509);
and U7044 (N_7044,N_6504,N_6290);
or U7045 (N_7045,N_6454,N_6368);
and U7046 (N_7046,N_6330,N_6531);
and U7047 (N_7047,N_6857,N_6423);
nor U7048 (N_7048,N_6598,N_6962);
nor U7049 (N_7049,N_6937,N_6496);
nand U7050 (N_7050,N_6770,N_6627);
nor U7051 (N_7051,N_6437,N_6768);
nand U7052 (N_7052,N_6356,N_6093);
nand U7053 (N_7053,N_6197,N_6780);
xnor U7054 (N_7054,N_6426,N_6060);
nand U7055 (N_7055,N_6868,N_6455);
nor U7056 (N_7056,N_6347,N_6893);
nor U7057 (N_7057,N_6588,N_6083);
nor U7058 (N_7058,N_6950,N_6609);
or U7059 (N_7059,N_6932,N_6828);
nand U7060 (N_7060,N_6364,N_6769);
and U7061 (N_7061,N_6566,N_6453);
or U7062 (N_7062,N_6752,N_6092);
nor U7063 (N_7063,N_6998,N_6892);
or U7064 (N_7064,N_6265,N_6329);
and U7065 (N_7065,N_6136,N_6910);
nand U7066 (N_7066,N_6503,N_6896);
nor U7067 (N_7067,N_6659,N_6846);
and U7068 (N_7068,N_6587,N_6771);
nor U7069 (N_7069,N_6570,N_6672);
nand U7070 (N_7070,N_6580,N_6547);
or U7071 (N_7071,N_6418,N_6762);
and U7072 (N_7072,N_6007,N_6240);
and U7073 (N_7073,N_6452,N_6131);
or U7074 (N_7074,N_6089,N_6431);
nor U7075 (N_7075,N_6322,N_6499);
or U7076 (N_7076,N_6379,N_6935);
nand U7077 (N_7077,N_6577,N_6059);
nor U7078 (N_7078,N_6984,N_6130);
or U7079 (N_7079,N_6076,N_6777);
nor U7080 (N_7080,N_6024,N_6849);
nand U7081 (N_7081,N_6515,N_6833);
or U7082 (N_7082,N_6339,N_6635);
or U7083 (N_7083,N_6800,N_6061);
and U7084 (N_7084,N_6782,N_6629);
nand U7085 (N_7085,N_6933,N_6562);
or U7086 (N_7086,N_6365,N_6994);
nor U7087 (N_7087,N_6390,N_6468);
nor U7088 (N_7088,N_6530,N_6837);
or U7089 (N_7089,N_6350,N_6249);
nor U7090 (N_7090,N_6393,N_6345);
nand U7091 (N_7091,N_6711,N_6812);
nand U7092 (N_7092,N_6605,N_6697);
or U7093 (N_7093,N_6840,N_6712);
nor U7094 (N_7094,N_6664,N_6544);
and U7095 (N_7095,N_6886,N_6569);
nand U7096 (N_7096,N_6299,N_6766);
nor U7097 (N_7097,N_6009,N_6282);
or U7098 (N_7098,N_6796,N_6128);
nand U7099 (N_7099,N_6263,N_6222);
or U7100 (N_7100,N_6978,N_6206);
nor U7101 (N_7101,N_6874,N_6891);
nor U7102 (N_7102,N_6255,N_6420);
or U7103 (N_7103,N_6946,N_6909);
nor U7104 (N_7104,N_6417,N_6829);
nand U7105 (N_7105,N_6253,N_6919);
nand U7106 (N_7106,N_6087,N_6145);
nand U7107 (N_7107,N_6344,N_6825);
nand U7108 (N_7108,N_6451,N_6668);
nor U7109 (N_7109,N_6890,N_6912);
nor U7110 (N_7110,N_6943,N_6907);
and U7111 (N_7111,N_6410,N_6311);
or U7112 (N_7112,N_6187,N_6900);
and U7113 (N_7113,N_6218,N_6475);
and U7114 (N_7114,N_6212,N_6854);
or U7115 (N_7115,N_6589,N_6223);
or U7116 (N_7116,N_6799,N_6068);
nand U7117 (N_7117,N_6980,N_6692);
nor U7118 (N_7118,N_6966,N_6600);
nor U7119 (N_7119,N_6326,N_6791);
or U7120 (N_7120,N_6005,N_6784);
nand U7121 (N_7121,N_6623,N_6338);
nor U7122 (N_7122,N_6818,N_6924);
and U7123 (N_7123,N_6883,N_6313);
and U7124 (N_7124,N_6018,N_6897);
nor U7125 (N_7125,N_6861,N_6824);
and U7126 (N_7126,N_6838,N_6642);
nor U7127 (N_7127,N_6902,N_6397);
nand U7128 (N_7128,N_6944,N_6184);
nor U7129 (N_7129,N_6622,N_6404);
and U7130 (N_7130,N_6217,N_6655);
nor U7131 (N_7131,N_6285,N_6781);
nor U7132 (N_7132,N_6823,N_6363);
or U7133 (N_7133,N_6077,N_6084);
nand U7134 (N_7134,N_6688,N_6295);
nor U7135 (N_7135,N_6244,N_6822);
or U7136 (N_7136,N_6091,N_6178);
nand U7137 (N_7137,N_6687,N_6232);
nand U7138 (N_7138,N_6351,N_6168);
nand U7139 (N_7139,N_6786,N_6540);
nand U7140 (N_7140,N_6614,N_6287);
xnor U7141 (N_7141,N_6596,N_6072);
nor U7142 (N_7142,N_6663,N_6159);
and U7143 (N_7143,N_6301,N_6794);
nand U7144 (N_7144,N_6537,N_6096);
nand U7145 (N_7145,N_6526,N_6308);
and U7146 (N_7146,N_6014,N_6449);
nand U7147 (N_7147,N_6247,N_6641);
nor U7148 (N_7148,N_6384,N_6288);
or U7149 (N_7149,N_6680,N_6394);
nand U7150 (N_7150,N_6971,N_6065);
nand U7151 (N_7151,N_6141,N_6133);
xor U7152 (N_7152,N_6051,N_6274);
or U7153 (N_7153,N_6209,N_6914);
or U7154 (N_7154,N_6033,N_6876);
nor U7155 (N_7155,N_6066,N_6134);
and U7156 (N_7156,N_6383,N_6895);
nor U7157 (N_7157,N_6923,N_6964);
nand U7158 (N_7158,N_6518,N_6603);
nand U7159 (N_7159,N_6006,N_6038);
or U7160 (N_7160,N_6508,N_6252);
nand U7161 (N_7161,N_6592,N_6165);
nand U7162 (N_7162,N_6992,N_6429);
or U7163 (N_7163,N_6583,N_6069);
nor U7164 (N_7164,N_6699,N_6319);
nand U7165 (N_7165,N_6754,N_6070);
and U7166 (N_7166,N_6948,N_6953);
or U7167 (N_7167,N_6665,N_6767);
or U7168 (N_7168,N_6507,N_6389);
nor U7169 (N_7169,N_6602,N_6158);
nor U7170 (N_7170,N_6990,N_6549);
nand U7171 (N_7171,N_6008,N_6485);
or U7172 (N_7172,N_6186,N_6053);
nand U7173 (N_7173,N_6559,N_6154);
or U7174 (N_7174,N_6422,N_6085);
and U7175 (N_7175,N_6027,N_6750);
and U7176 (N_7176,N_6866,N_6965);
or U7177 (N_7177,N_6243,N_6434);
nor U7178 (N_7178,N_6331,N_6458);
nor U7179 (N_7179,N_6214,N_6921);
nor U7180 (N_7180,N_6929,N_6682);
nand U7181 (N_7181,N_6694,N_6864);
and U7182 (N_7182,N_6310,N_6880);
nand U7183 (N_7183,N_6367,N_6114);
nor U7184 (N_7184,N_6764,N_6300);
or U7185 (N_7185,N_6022,N_6233);
or U7186 (N_7186,N_6149,N_6219);
nand U7187 (N_7187,N_6237,N_6400);
and U7188 (N_7188,N_6512,N_6976);
or U7189 (N_7189,N_6188,N_6955);
nand U7190 (N_7190,N_6925,N_6029);
nor U7191 (N_7191,N_6408,N_6432);
nor U7192 (N_7192,N_6425,N_6164);
nand U7193 (N_7193,N_6306,N_6064);
nor U7194 (N_7194,N_6567,N_6124);
or U7195 (N_7195,N_6147,N_6289);
nor U7196 (N_7196,N_6353,N_6621);
and U7197 (N_7197,N_6776,N_6732);
or U7198 (N_7198,N_6107,N_6905);
nor U7199 (N_7199,N_6806,N_6506);
nor U7200 (N_7200,N_6049,N_6294);
nor U7201 (N_7201,N_6775,N_6025);
nand U7202 (N_7202,N_6019,N_6701);
nor U7203 (N_7203,N_6557,N_6456);
nor U7204 (N_7204,N_6755,N_6182);
and U7205 (N_7205,N_6427,N_6004);
or U7206 (N_7206,N_6380,N_6554);
or U7207 (N_7207,N_6057,N_6620);
nor U7208 (N_7208,N_6239,N_6100);
or U7209 (N_7209,N_6123,N_6346);
nor U7210 (N_7210,N_6477,N_6584);
and U7211 (N_7211,N_6626,N_6035);
and U7212 (N_7212,N_6152,N_6738);
nor U7213 (N_7213,N_6284,N_6525);
and U7214 (N_7214,N_6773,N_6667);
nand U7215 (N_7215,N_6067,N_6143);
nand U7216 (N_7216,N_6714,N_6011);
nor U7217 (N_7217,N_6542,N_6280);
or U7218 (N_7218,N_6079,N_6472);
nor U7219 (N_7219,N_6207,N_6607);
nor U7220 (N_7220,N_6640,N_6724);
nand U7221 (N_7221,N_6481,N_6129);
or U7222 (N_7222,N_6785,N_6256);
nor U7223 (N_7223,N_6360,N_6858);
or U7224 (N_7224,N_6576,N_6625);
or U7225 (N_7225,N_6117,N_6113);
or U7226 (N_7226,N_6759,N_6538);
or U7227 (N_7227,N_6517,N_6705);
nor U7228 (N_7228,N_6443,N_6877);
and U7229 (N_7229,N_6120,N_6988);
or U7230 (N_7230,N_6643,N_6774);
and U7231 (N_7231,N_6644,N_6213);
and U7232 (N_7232,N_6421,N_6751);
nand U7233 (N_7233,N_6012,N_6445);
or U7234 (N_7234,N_6843,N_6591);
nand U7235 (N_7235,N_6438,N_6808);
nor U7236 (N_7236,N_6970,N_6302);
and U7237 (N_7237,N_6963,N_6082);
nor U7238 (N_7238,N_6078,N_6409);
nand U7239 (N_7239,N_6869,N_6804);
and U7240 (N_7240,N_6686,N_6928);
nor U7241 (N_7241,N_6863,N_6817);
nand U7242 (N_7242,N_6448,N_6888);
nand U7243 (N_7243,N_6690,N_6832);
or U7244 (N_7244,N_6718,N_6391);
nor U7245 (N_7245,N_6565,N_6327);
or U7246 (N_7246,N_6851,N_6987);
nor U7247 (N_7247,N_6741,N_6195);
and U7248 (N_7248,N_6495,N_6046);
nor U7249 (N_7249,N_6646,N_6558);
or U7250 (N_7250,N_6974,N_6899);
nor U7251 (N_7251,N_6702,N_6793);
nand U7252 (N_7252,N_6283,N_6094);
nand U7253 (N_7253,N_6572,N_6266);
nand U7254 (N_7254,N_6396,N_6706);
and U7255 (N_7255,N_6037,N_6634);
nor U7256 (N_7256,N_6163,N_6074);
and U7257 (N_7257,N_6997,N_6238);
or U7258 (N_7258,N_6939,N_6631);
nand U7259 (N_7259,N_6235,N_6709);
or U7260 (N_7260,N_6820,N_6304);
nand U7261 (N_7261,N_6166,N_6862);
nand U7262 (N_7262,N_6847,N_6071);
nor U7263 (N_7263,N_6673,N_6852);
xor U7264 (N_7264,N_6632,N_6802);
and U7265 (N_7265,N_6132,N_6952);
and U7266 (N_7266,N_6871,N_6653);
or U7267 (N_7267,N_6882,N_6073);
and U7268 (N_7268,N_6150,N_6743);
nor U7269 (N_7269,N_6349,N_6881);
nor U7270 (N_7270,N_6873,N_6548);
nand U7271 (N_7271,N_6205,N_6333);
and U7272 (N_7272,N_6999,N_6772);
nor U7273 (N_7273,N_6760,N_6315);
nand U7274 (N_7274,N_6906,N_6636);
nand U7275 (N_7275,N_6728,N_6292);
nor U7276 (N_7276,N_6148,N_6783);
and U7277 (N_7277,N_6413,N_6405);
or U7278 (N_7278,N_6834,N_6248);
or U7279 (N_7279,N_6585,N_6279);
and U7280 (N_7280,N_6259,N_6210);
nand U7281 (N_7281,N_6521,N_6606);
or U7282 (N_7282,N_6245,N_6654);
nand U7283 (N_7283,N_6720,N_6830);
nor U7284 (N_7284,N_6221,N_6028);
nand U7285 (N_7285,N_6484,N_6519);
and U7286 (N_7286,N_6352,N_6945);
nor U7287 (N_7287,N_6582,N_6169);
nand U7288 (N_7288,N_6662,N_6489);
or U7289 (N_7289,N_6461,N_6372);
nor U7290 (N_7290,N_6323,N_6798);
nand U7291 (N_7291,N_6194,N_6742);
nor U7292 (N_7292,N_6015,N_6696);
or U7293 (N_7293,N_6875,N_6348);
nand U7294 (N_7294,N_6727,N_6859);
or U7295 (N_7295,N_6551,N_6043);
nor U7296 (N_7296,N_6801,N_6457);
and U7297 (N_7297,N_6478,N_6270);
nand U7298 (N_7298,N_6419,N_6740);
nand U7299 (N_7299,N_6949,N_6993);
nor U7300 (N_7300,N_6860,N_6382);
and U7301 (N_7301,N_6552,N_6991);
nand U7302 (N_7302,N_6805,N_6246);
or U7303 (N_7303,N_6224,N_6870);
and U7304 (N_7304,N_6357,N_6707);
or U7305 (N_7305,N_6715,N_6328);
nand U7306 (N_7306,N_6303,N_6753);
and U7307 (N_7307,N_6286,N_6487);
nor U7308 (N_7308,N_6633,N_6550);
nand U7309 (N_7309,N_6325,N_6713);
nor U7310 (N_7310,N_6810,N_6336);
and U7311 (N_7311,N_6985,N_6139);
nand U7312 (N_7312,N_6324,N_6318);
nor U7313 (N_7313,N_6176,N_6691);
nor U7314 (N_7314,N_6435,N_6938);
and U7315 (N_7315,N_6402,N_6293);
or U7316 (N_7316,N_6258,N_6001);
or U7317 (N_7317,N_6872,N_6479);
and U7318 (N_7318,N_6995,N_6220);
or U7319 (N_7319,N_6230,N_6660);
nor U7320 (N_7320,N_6726,N_6695);
and U7321 (N_7321,N_6407,N_6528);
or U7322 (N_7322,N_6211,N_6278);
or U7323 (N_7323,N_6658,N_6520);
and U7324 (N_7324,N_6157,N_6160);
and U7325 (N_7325,N_6354,N_6568);
or U7326 (N_7326,N_6374,N_6493);
nand U7327 (N_7327,N_6267,N_6615);
nor U7328 (N_7328,N_6619,N_6056);
or U7329 (N_7329,N_6167,N_6108);
or U7330 (N_7330,N_6483,N_6047);
nor U7331 (N_7331,N_6748,N_6564);
nand U7332 (N_7332,N_6460,N_6839);
and U7333 (N_7333,N_6972,N_6617);
and U7334 (N_7334,N_6386,N_6739);
nor U7335 (N_7335,N_6579,N_6704);
or U7336 (N_7336,N_6013,N_6229);
and U7337 (N_7337,N_6556,N_6112);
or U7338 (N_7338,N_6098,N_6841);
or U7339 (N_7339,N_6126,N_6887);
and U7340 (N_7340,N_6725,N_6026);
nor U7341 (N_7341,N_6201,N_6594);
or U7342 (N_7342,N_6779,N_6459);
and U7343 (N_7343,N_6657,N_6366);
nor U7344 (N_7344,N_6102,N_6415);
and U7345 (N_7345,N_6442,N_6844);
nor U7346 (N_7346,N_6936,N_6398);
nor U7347 (N_7347,N_6700,N_6251);
or U7348 (N_7348,N_6444,N_6052);
or U7349 (N_7349,N_6610,N_6502);
nor U7350 (N_7350,N_6790,N_6464);
or U7351 (N_7351,N_6153,N_6722);
and U7352 (N_7352,N_6942,N_6155);
and U7353 (N_7353,N_6482,N_6827);
or U7354 (N_7354,N_6281,N_6369);
or U7355 (N_7355,N_6885,N_6135);
nand U7356 (N_7356,N_6081,N_6179);
and U7357 (N_7357,N_6639,N_6370);
nor U7358 (N_7358,N_6355,N_6560);
or U7359 (N_7359,N_6269,N_6819);
or U7360 (N_7360,N_6797,N_6671);
and U7361 (N_7361,N_6967,N_6291);
or U7362 (N_7362,N_6361,N_6125);
and U7363 (N_7363,N_6103,N_6388);
and U7364 (N_7364,N_6378,N_6309);
nand U7365 (N_7365,N_6036,N_6809);
nor U7366 (N_7366,N_6652,N_6529);
and U7367 (N_7367,N_6666,N_6826);
nor U7368 (N_7368,N_6463,N_6305);
and U7369 (N_7369,N_6095,N_6693);
and U7370 (N_7370,N_6171,N_6020);
or U7371 (N_7371,N_6044,N_6063);
and U7372 (N_7372,N_6162,N_6058);
nor U7373 (N_7373,N_6630,N_6439);
nand U7374 (N_7374,N_6473,N_6571);
xnor U7375 (N_7375,N_6231,N_6651);
nor U7376 (N_7376,N_6505,N_6561);
or U7377 (N_7377,N_6734,N_6941);
nand U7378 (N_7378,N_6110,N_6039);
nor U7379 (N_7379,N_6894,N_6744);
nand U7380 (N_7380,N_6227,N_6901);
or U7381 (N_7381,N_6811,N_6204);
nand U7382 (N_7382,N_6034,N_6983);
or U7383 (N_7383,N_6342,N_6532);
nand U7384 (N_7384,N_6010,N_6086);
nand U7385 (N_7385,N_6030,N_6471);
nor U7386 (N_7386,N_6954,N_6684);
or U7387 (N_7387,N_6277,N_6016);
or U7388 (N_7388,N_6645,N_6189);
nor U7389 (N_7389,N_6973,N_6151);
nand U7390 (N_7390,N_6513,N_6424);
or U7391 (N_7391,N_6414,N_6903);
nand U7392 (N_7392,N_6729,N_6737);
and U7393 (N_7393,N_6821,N_6399);
nor U7394 (N_7394,N_6467,N_6628);
or U7395 (N_7395,N_6446,N_6719);
or U7396 (N_7396,N_6835,N_6661);
nand U7397 (N_7397,N_6017,N_6275);
nand U7398 (N_7398,N_6703,N_6216);
nand U7399 (N_7399,N_6215,N_6264);
nand U7400 (N_7400,N_6795,N_6003);
nand U7401 (N_7401,N_6756,N_6054);
nand U7402 (N_7402,N_6430,N_6491);
xnor U7403 (N_7403,N_6930,N_6865);
nor U7404 (N_7404,N_6021,N_6146);
or U7405 (N_7405,N_6142,N_6273);
or U7406 (N_7406,N_6685,N_6681);
nor U7407 (N_7407,N_6498,N_6608);
nor U7408 (N_7408,N_6581,N_6276);
nor U7409 (N_7409,N_6170,N_6332);
and U7410 (N_7410,N_6916,N_6555);
nor U7411 (N_7411,N_6735,N_6226);
nand U7412 (N_7412,N_6497,N_6392);
and U7413 (N_7413,N_6000,N_6260);
nand U7414 (N_7414,N_6807,N_6116);
and U7415 (N_7415,N_6373,N_6969);
or U7416 (N_7416,N_6172,N_6708);
or U7417 (N_7417,N_6788,N_6371);
and U7418 (N_7418,N_6183,N_6524);
nand U7419 (N_7419,N_6927,N_6254);
nor U7420 (N_7420,N_6986,N_6778);
nand U7421 (N_7421,N_6341,N_6250);
and U7422 (N_7422,N_6546,N_6181);
nor U7423 (N_7423,N_6731,N_6316);
and U7424 (N_7424,N_6062,N_6241);
nor U7425 (N_7425,N_6563,N_6196);
nor U7426 (N_7426,N_6683,N_6578);
and U7427 (N_7427,N_6097,N_6173);
or U7428 (N_7428,N_6200,N_6271);
nand U7429 (N_7429,N_6099,N_6105);
nand U7430 (N_7430,N_6050,N_6958);
or U7431 (N_7431,N_6486,N_6115);
or U7432 (N_7432,N_6387,N_6911);
or U7433 (N_7433,N_6670,N_6814);
and U7434 (N_7434,N_6375,N_6118);
or U7435 (N_7435,N_6848,N_6590);
nor U7436 (N_7436,N_6002,N_6611);
nor U7437 (N_7437,N_6395,N_6956);
nand U7438 (N_7438,N_6494,N_6510);
nor U7439 (N_7439,N_6934,N_6815);
or U7440 (N_7440,N_6842,N_6320);
and U7441 (N_7441,N_6789,N_6048);
nor U7442 (N_7442,N_6104,N_6406);
and U7443 (N_7443,N_6803,N_6416);
nand U7444 (N_7444,N_6679,N_6595);
nand U7445 (N_7445,N_6314,N_6931);
nand U7446 (N_7446,N_6710,N_6340);
nand U7447 (N_7447,N_6474,N_6090);
nand U7448 (N_7448,N_6761,N_6447);
xnor U7449 (N_7449,N_6268,N_6736);
or U7450 (N_7450,N_6140,N_6792);
nor U7451 (N_7451,N_6337,N_6307);
nand U7452 (N_7452,N_6675,N_6982);
or U7453 (N_7453,N_6436,N_6533);
nand U7454 (N_7454,N_6979,N_6358);
or U7455 (N_7455,N_6647,N_6541);
nand U7456 (N_7456,N_6624,N_6156);
nand U7457 (N_7457,N_6601,N_6522);
nor U7458 (N_7458,N_6177,N_6878);
nand U7459 (N_7459,N_6088,N_6121);
and U7460 (N_7460,N_6650,N_6535);
nor U7461 (N_7461,N_6412,N_6032);
or U7462 (N_7462,N_6119,N_6536);
nor U7463 (N_7463,N_6763,N_6480);
nor U7464 (N_7464,N_6746,N_6813);
nand U7465 (N_7465,N_6490,N_6613);
nand U7466 (N_7466,N_6904,N_6450);
nand U7467 (N_7467,N_6185,N_6042);
and U7468 (N_7468,N_6202,N_6747);
or U7469 (N_7469,N_6867,N_6915);
xnor U7470 (N_7470,N_6441,N_6225);
nand U7471 (N_7471,N_6977,N_6381);
or U7472 (N_7472,N_6199,N_6677);
nor U7473 (N_7473,N_6045,N_6334);
nand U7474 (N_7474,N_6649,N_6101);
nor U7475 (N_7475,N_6377,N_6343);
nand U7476 (N_7476,N_6470,N_6190);
nand U7477 (N_7477,N_6856,N_6127);
and U7478 (N_7478,N_6656,N_6638);
nand U7479 (N_7479,N_6539,N_6612);
and U7480 (N_7480,N_6106,N_6321);
nand U7481 (N_7481,N_6514,N_6545);
nand U7482 (N_7482,N_6257,N_6959);
nand U7483 (N_7483,N_6599,N_6488);
nand U7484 (N_7484,N_6144,N_6534);
and U7485 (N_7485,N_6137,N_6261);
xor U7486 (N_7486,N_6511,N_6996);
and U7487 (N_7487,N_6926,N_6816);
xor U7488 (N_7488,N_6586,N_6317);
or U7489 (N_7489,N_6236,N_6440);
and U7490 (N_7490,N_6879,N_6574);
nand U7491 (N_7491,N_6940,N_6161);
and U7492 (N_7492,N_6917,N_6637);
nand U7493 (N_7493,N_6272,N_6543);
nor U7494 (N_7494,N_6845,N_6401);
or U7495 (N_7495,N_6203,N_6055);
and U7496 (N_7496,N_6362,N_6573);
and U7497 (N_7497,N_6428,N_6898);
or U7498 (N_7498,N_6922,N_6920);
and U7499 (N_7499,N_6575,N_6884);
or U7500 (N_7500,N_6169,N_6193);
nor U7501 (N_7501,N_6312,N_6170);
nor U7502 (N_7502,N_6378,N_6815);
and U7503 (N_7503,N_6569,N_6183);
nor U7504 (N_7504,N_6459,N_6238);
nand U7505 (N_7505,N_6335,N_6205);
nand U7506 (N_7506,N_6698,N_6135);
or U7507 (N_7507,N_6399,N_6902);
and U7508 (N_7508,N_6805,N_6921);
or U7509 (N_7509,N_6449,N_6975);
or U7510 (N_7510,N_6569,N_6253);
nor U7511 (N_7511,N_6454,N_6528);
nand U7512 (N_7512,N_6258,N_6445);
or U7513 (N_7513,N_6299,N_6823);
nand U7514 (N_7514,N_6401,N_6009);
or U7515 (N_7515,N_6996,N_6372);
nand U7516 (N_7516,N_6076,N_6131);
nand U7517 (N_7517,N_6869,N_6036);
nor U7518 (N_7518,N_6812,N_6106);
nand U7519 (N_7519,N_6230,N_6068);
and U7520 (N_7520,N_6828,N_6829);
nand U7521 (N_7521,N_6044,N_6754);
and U7522 (N_7522,N_6563,N_6167);
nor U7523 (N_7523,N_6339,N_6261);
nor U7524 (N_7524,N_6860,N_6690);
and U7525 (N_7525,N_6474,N_6511);
and U7526 (N_7526,N_6640,N_6858);
and U7527 (N_7527,N_6169,N_6952);
or U7528 (N_7528,N_6454,N_6815);
or U7529 (N_7529,N_6656,N_6342);
and U7530 (N_7530,N_6642,N_6420);
nand U7531 (N_7531,N_6276,N_6407);
nor U7532 (N_7532,N_6782,N_6238);
and U7533 (N_7533,N_6636,N_6090);
nor U7534 (N_7534,N_6673,N_6373);
nand U7535 (N_7535,N_6843,N_6771);
nor U7536 (N_7536,N_6786,N_6108);
or U7537 (N_7537,N_6738,N_6263);
or U7538 (N_7538,N_6649,N_6737);
and U7539 (N_7539,N_6902,N_6440);
or U7540 (N_7540,N_6797,N_6265);
or U7541 (N_7541,N_6540,N_6512);
and U7542 (N_7542,N_6824,N_6205);
and U7543 (N_7543,N_6916,N_6155);
nor U7544 (N_7544,N_6733,N_6509);
nor U7545 (N_7545,N_6228,N_6639);
and U7546 (N_7546,N_6018,N_6856);
nand U7547 (N_7547,N_6870,N_6497);
and U7548 (N_7548,N_6762,N_6620);
nand U7549 (N_7549,N_6820,N_6014);
and U7550 (N_7550,N_6519,N_6935);
or U7551 (N_7551,N_6884,N_6531);
nor U7552 (N_7552,N_6155,N_6274);
nor U7553 (N_7553,N_6697,N_6974);
nand U7554 (N_7554,N_6374,N_6394);
nor U7555 (N_7555,N_6864,N_6283);
xnor U7556 (N_7556,N_6746,N_6064);
nor U7557 (N_7557,N_6560,N_6450);
nand U7558 (N_7558,N_6644,N_6525);
nand U7559 (N_7559,N_6485,N_6641);
or U7560 (N_7560,N_6732,N_6327);
and U7561 (N_7561,N_6788,N_6177);
nand U7562 (N_7562,N_6889,N_6485);
and U7563 (N_7563,N_6681,N_6348);
nand U7564 (N_7564,N_6968,N_6991);
or U7565 (N_7565,N_6091,N_6222);
and U7566 (N_7566,N_6110,N_6210);
nand U7567 (N_7567,N_6785,N_6009);
or U7568 (N_7568,N_6204,N_6224);
nand U7569 (N_7569,N_6390,N_6394);
nand U7570 (N_7570,N_6154,N_6310);
nor U7571 (N_7571,N_6991,N_6391);
nand U7572 (N_7572,N_6291,N_6568);
or U7573 (N_7573,N_6927,N_6301);
or U7574 (N_7574,N_6926,N_6235);
nor U7575 (N_7575,N_6335,N_6695);
nand U7576 (N_7576,N_6046,N_6037);
or U7577 (N_7577,N_6822,N_6296);
nand U7578 (N_7578,N_6384,N_6388);
nand U7579 (N_7579,N_6249,N_6703);
nand U7580 (N_7580,N_6672,N_6290);
and U7581 (N_7581,N_6903,N_6847);
and U7582 (N_7582,N_6156,N_6190);
or U7583 (N_7583,N_6610,N_6141);
nand U7584 (N_7584,N_6843,N_6628);
or U7585 (N_7585,N_6119,N_6598);
nand U7586 (N_7586,N_6322,N_6476);
nor U7587 (N_7587,N_6418,N_6513);
nand U7588 (N_7588,N_6983,N_6085);
or U7589 (N_7589,N_6844,N_6904);
nor U7590 (N_7590,N_6116,N_6580);
nor U7591 (N_7591,N_6042,N_6326);
nor U7592 (N_7592,N_6411,N_6297);
and U7593 (N_7593,N_6639,N_6742);
or U7594 (N_7594,N_6356,N_6437);
nor U7595 (N_7595,N_6011,N_6155);
nor U7596 (N_7596,N_6818,N_6154);
nor U7597 (N_7597,N_6189,N_6035);
and U7598 (N_7598,N_6800,N_6123);
and U7599 (N_7599,N_6558,N_6104);
or U7600 (N_7600,N_6493,N_6641);
nand U7601 (N_7601,N_6396,N_6818);
nand U7602 (N_7602,N_6226,N_6703);
and U7603 (N_7603,N_6355,N_6383);
and U7604 (N_7604,N_6249,N_6098);
nand U7605 (N_7605,N_6085,N_6126);
nand U7606 (N_7606,N_6867,N_6552);
and U7607 (N_7607,N_6140,N_6039);
nand U7608 (N_7608,N_6374,N_6968);
and U7609 (N_7609,N_6943,N_6462);
nand U7610 (N_7610,N_6148,N_6808);
nand U7611 (N_7611,N_6025,N_6267);
nand U7612 (N_7612,N_6958,N_6677);
nand U7613 (N_7613,N_6575,N_6383);
and U7614 (N_7614,N_6387,N_6793);
or U7615 (N_7615,N_6670,N_6917);
nand U7616 (N_7616,N_6697,N_6222);
nand U7617 (N_7617,N_6031,N_6458);
nor U7618 (N_7618,N_6129,N_6461);
nor U7619 (N_7619,N_6636,N_6684);
nand U7620 (N_7620,N_6842,N_6032);
nor U7621 (N_7621,N_6397,N_6775);
nor U7622 (N_7622,N_6566,N_6741);
nand U7623 (N_7623,N_6945,N_6920);
or U7624 (N_7624,N_6366,N_6646);
and U7625 (N_7625,N_6806,N_6692);
and U7626 (N_7626,N_6800,N_6115);
nor U7627 (N_7627,N_6638,N_6031);
nand U7628 (N_7628,N_6488,N_6304);
nor U7629 (N_7629,N_6702,N_6990);
or U7630 (N_7630,N_6739,N_6714);
or U7631 (N_7631,N_6752,N_6104);
or U7632 (N_7632,N_6817,N_6047);
nand U7633 (N_7633,N_6886,N_6201);
nand U7634 (N_7634,N_6403,N_6563);
nor U7635 (N_7635,N_6945,N_6107);
or U7636 (N_7636,N_6528,N_6731);
and U7637 (N_7637,N_6893,N_6668);
and U7638 (N_7638,N_6093,N_6304);
or U7639 (N_7639,N_6541,N_6198);
or U7640 (N_7640,N_6779,N_6724);
nand U7641 (N_7641,N_6329,N_6940);
and U7642 (N_7642,N_6126,N_6975);
nand U7643 (N_7643,N_6850,N_6872);
nor U7644 (N_7644,N_6513,N_6083);
and U7645 (N_7645,N_6840,N_6225);
or U7646 (N_7646,N_6055,N_6569);
or U7647 (N_7647,N_6426,N_6851);
and U7648 (N_7648,N_6129,N_6720);
and U7649 (N_7649,N_6810,N_6515);
or U7650 (N_7650,N_6465,N_6513);
nand U7651 (N_7651,N_6504,N_6757);
nor U7652 (N_7652,N_6154,N_6007);
nor U7653 (N_7653,N_6925,N_6518);
nand U7654 (N_7654,N_6484,N_6680);
nand U7655 (N_7655,N_6130,N_6264);
nor U7656 (N_7656,N_6545,N_6138);
and U7657 (N_7657,N_6454,N_6788);
nand U7658 (N_7658,N_6849,N_6357);
or U7659 (N_7659,N_6991,N_6809);
nor U7660 (N_7660,N_6724,N_6548);
nand U7661 (N_7661,N_6148,N_6615);
nand U7662 (N_7662,N_6657,N_6819);
or U7663 (N_7663,N_6064,N_6958);
and U7664 (N_7664,N_6136,N_6689);
nand U7665 (N_7665,N_6114,N_6252);
nor U7666 (N_7666,N_6955,N_6596);
or U7667 (N_7667,N_6003,N_6282);
nor U7668 (N_7668,N_6327,N_6635);
or U7669 (N_7669,N_6347,N_6795);
nor U7670 (N_7670,N_6184,N_6826);
or U7671 (N_7671,N_6863,N_6086);
or U7672 (N_7672,N_6671,N_6965);
xnor U7673 (N_7673,N_6975,N_6713);
nand U7674 (N_7674,N_6342,N_6646);
and U7675 (N_7675,N_6871,N_6832);
and U7676 (N_7676,N_6923,N_6807);
nor U7677 (N_7677,N_6730,N_6111);
and U7678 (N_7678,N_6766,N_6339);
nor U7679 (N_7679,N_6798,N_6349);
or U7680 (N_7680,N_6872,N_6575);
nand U7681 (N_7681,N_6204,N_6595);
nand U7682 (N_7682,N_6683,N_6307);
nand U7683 (N_7683,N_6305,N_6995);
or U7684 (N_7684,N_6382,N_6734);
nand U7685 (N_7685,N_6775,N_6388);
nor U7686 (N_7686,N_6682,N_6863);
and U7687 (N_7687,N_6946,N_6517);
nand U7688 (N_7688,N_6078,N_6890);
nand U7689 (N_7689,N_6211,N_6217);
nand U7690 (N_7690,N_6517,N_6747);
or U7691 (N_7691,N_6704,N_6266);
nor U7692 (N_7692,N_6781,N_6938);
nand U7693 (N_7693,N_6551,N_6718);
nand U7694 (N_7694,N_6595,N_6467);
and U7695 (N_7695,N_6253,N_6540);
nand U7696 (N_7696,N_6480,N_6980);
nor U7697 (N_7697,N_6548,N_6736);
or U7698 (N_7698,N_6609,N_6499);
and U7699 (N_7699,N_6449,N_6316);
nand U7700 (N_7700,N_6371,N_6634);
nor U7701 (N_7701,N_6537,N_6655);
or U7702 (N_7702,N_6190,N_6276);
and U7703 (N_7703,N_6845,N_6176);
and U7704 (N_7704,N_6212,N_6825);
or U7705 (N_7705,N_6411,N_6918);
and U7706 (N_7706,N_6954,N_6432);
nor U7707 (N_7707,N_6652,N_6992);
or U7708 (N_7708,N_6422,N_6800);
nand U7709 (N_7709,N_6112,N_6594);
and U7710 (N_7710,N_6575,N_6316);
or U7711 (N_7711,N_6020,N_6711);
and U7712 (N_7712,N_6325,N_6723);
or U7713 (N_7713,N_6412,N_6415);
or U7714 (N_7714,N_6850,N_6199);
nor U7715 (N_7715,N_6167,N_6202);
xor U7716 (N_7716,N_6408,N_6469);
or U7717 (N_7717,N_6707,N_6377);
and U7718 (N_7718,N_6537,N_6936);
nand U7719 (N_7719,N_6034,N_6485);
or U7720 (N_7720,N_6979,N_6030);
nor U7721 (N_7721,N_6928,N_6751);
nor U7722 (N_7722,N_6049,N_6557);
or U7723 (N_7723,N_6974,N_6661);
or U7724 (N_7724,N_6635,N_6620);
nand U7725 (N_7725,N_6598,N_6329);
nor U7726 (N_7726,N_6325,N_6383);
nor U7727 (N_7727,N_6071,N_6984);
xor U7728 (N_7728,N_6386,N_6987);
or U7729 (N_7729,N_6645,N_6256);
and U7730 (N_7730,N_6427,N_6505);
nor U7731 (N_7731,N_6978,N_6687);
nand U7732 (N_7732,N_6056,N_6841);
nand U7733 (N_7733,N_6589,N_6104);
or U7734 (N_7734,N_6299,N_6755);
nor U7735 (N_7735,N_6454,N_6918);
nand U7736 (N_7736,N_6125,N_6751);
and U7737 (N_7737,N_6632,N_6084);
or U7738 (N_7738,N_6663,N_6340);
nor U7739 (N_7739,N_6069,N_6679);
nor U7740 (N_7740,N_6091,N_6473);
and U7741 (N_7741,N_6655,N_6469);
and U7742 (N_7742,N_6453,N_6964);
or U7743 (N_7743,N_6793,N_6467);
nor U7744 (N_7744,N_6756,N_6192);
nor U7745 (N_7745,N_6141,N_6425);
and U7746 (N_7746,N_6577,N_6952);
and U7747 (N_7747,N_6666,N_6298);
or U7748 (N_7748,N_6287,N_6433);
and U7749 (N_7749,N_6369,N_6228);
nor U7750 (N_7750,N_6633,N_6235);
and U7751 (N_7751,N_6619,N_6104);
or U7752 (N_7752,N_6709,N_6359);
or U7753 (N_7753,N_6305,N_6834);
nor U7754 (N_7754,N_6524,N_6202);
or U7755 (N_7755,N_6631,N_6751);
nor U7756 (N_7756,N_6645,N_6183);
nand U7757 (N_7757,N_6468,N_6248);
or U7758 (N_7758,N_6023,N_6417);
and U7759 (N_7759,N_6668,N_6299);
and U7760 (N_7760,N_6694,N_6505);
nand U7761 (N_7761,N_6072,N_6308);
nor U7762 (N_7762,N_6674,N_6461);
or U7763 (N_7763,N_6865,N_6876);
or U7764 (N_7764,N_6208,N_6673);
and U7765 (N_7765,N_6131,N_6520);
nand U7766 (N_7766,N_6870,N_6332);
nor U7767 (N_7767,N_6448,N_6076);
or U7768 (N_7768,N_6332,N_6025);
nor U7769 (N_7769,N_6016,N_6987);
or U7770 (N_7770,N_6330,N_6973);
and U7771 (N_7771,N_6108,N_6353);
nand U7772 (N_7772,N_6783,N_6288);
nand U7773 (N_7773,N_6470,N_6700);
or U7774 (N_7774,N_6309,N_6648);
and U7775 (N_7775,N_6826,N_6501);
and U7776 (N_7776,N_6568,N_6821);
and U7777 (N_7777,N_6165,N_6429);
and U7778 (N_7778,N_6883,N_6680);
nor U7779 (N_7779,N_6864,N_6865);
and U7780 (N_7780,N_6914,N_6819);
nor U7781 (N_7781,N_6767,N_6969);
xor U7782 (N_7782,N_6157,N_6930);
nor U7783 (N_7783,N_6881,N_6542);
and U7784 (N_7784,N_6081,N_6767);
or U7785 (N_7785,N_6605,N_6498);
nor U7786 (N_7786,N_6499,N_6863);
nand U7787 (N_7787,N_6789,N_6376);
or U7788 (N_7788,N_6471,N_6933);
nor U7789 (N_7789,N_6072,N_6451);
and U7790 (N_7790,N_6907,N_6925);
nand U7791 (N_7791,N_6479,N_6780);
and U7792 (N_7792,N_6219,N_6477);
or U7793 (N_7793,N_6735,N_6096);
and U7794 (N_7794,N_6380,N_6183);
or U7795 (N_7795,N_6575,N_6465);
nor U7796 (N_7796,N_6534,N_6929);
and U7797 (N_7797,N_6217,N_6024);
and U7798 (N_7798,N_6310,N_6637);
or U7799 (N_7799,N_6787,N_6539);
and U7800 (N_7800,N_6109,N_6617);
or U7801 (N_7801,N_6395,N_6659);
xor U7802 (N_7802,N_6869,N_6758);
nand U7803 (N_7803,N_6597,N_6371);
nand U7804 (N_7804,N_6728,N_6288);
and U7805 (N_7805,N_6707,N_6835);
nand U7806 (N_7806,N_6029,N_6325);
nand U7807 (N_7807,N_6097,N_6288);
nand U7808 (N_7808,N_6026,N_6038);
nor U7809 (N_7809,N_6494,N_6549);
or U7810 (N_7810,N_6418,N_6702);
and U7811 (N_7811,N_6213,N_6533);
nor U7812 (N_7812,N_6765,N_6775);
nand U7813 (N_7813,N_6095,N_6734);
or U7814 (N_7814,N_6420,N_6547);
nand U7815 (N_7815,N_6060,N_6717);
nor U7816 (N_7816,N_6232,N_6732);
nand U7817 (N_7817,N_6723,N_6209);
nor U7818 (N_7818,N_6614,N_6876);
nor U7819 (N_7819,N_6598,N_6024);
nor U7820 (N_7820,N_6606,N_6250);
nand U7821 (N_7821,N_6506,N_6393);
or U7822 (N_7822,N_6494,N_6835);
nor U7823 (N_7823,N_6636,N_6923);
and U7824 (N_7824,N_6508,N_6869);
nand U7825 (N_7825,N_6648,N_6676);
and U7826 (N_7826,N_6918,N_6111);
and U7827 (N_7827,N_6082,N_6401);
or U7828 (N_7828,N_6981,N_6082);
or U7829 (N_7829,N_6333,N_6451);
nor U7830 (N_7830,N_6021,N_6387);
or U7831 (N_7831,N_6514,N_6067);
nor U7832 (N_7832,N_6799,N_6699);
nand U7833 (N_7833,N_6308,N_6130);
nand U7834 (N_7834,N_6302,N_6907);
nor U7835 (N_7835,N_6534,N_6054);
and U7836 (N_7836,N_6879,N_6151);
or U7837 (N_7837,N_6748,N_6065);
nand U7838 (N_7838,N_6648,N_6307);
or U7839 (N_7839,N_6918,N_6913);
or U7840 (N_7840,N_6664,N_6907);
nor U7841 (N_7841,N_6299,N_6582);
or U7842 (N_7842,N_6305,N_6745);
nand U7843 (N_7843,N_6096,N_6566);
nor U7844 (N_7844,N_6845,N_6131);
nand U7845 (N_7845,N_6593,N_6675);
or U7846 (N_7846,N_6646,N_6753);
or U7847 (N_7847,N_6014,N_6257);
or U7848 (N_7848,N_6148,N_6562);
nor U7849 (N_7849,N_6631,N_6785);
nand U7850 (N_7850,N_6246,N_6248);
nand U7851 (N_7851,N_6518,N_6254);
or U7852 (N_7852,N_6558,N_6923);
nand U7853 (N_7853,N_6605,N_6339);
and U7854 (N_7854,N_6230,N_6522);
or U7855 (N_7855,N_6907,N_6485);
or U7856 (N_7856,N_6634,N_6914);
nor U7857 (N_7857,N_6010,N_6054);
nand U7858 (N_7858,N_6515,N_6441);
nor U7859 (N_7859,N_6699,N_6484);
nand U7860 (N_7860,N_6690,N_6478);
and U7861 (N_7861,N_6231,N_6998);
nand U7862 (N_7862,N_6577,N_6413);
nand U7863 (N_7863,N_6394,N_6497);
and U7864 (N_7864,N_6782,N_6883);
and U7865 (N_7865,N_6011,N_6934);
nand U7866 (N_7866,N_6636,N_6264);
nor U7867 (N_7867,N_6225,N_6299);
and U7868 (N_7868,N_6599,N_6669);
or U7869 (N_7869,N_6803,N_6105);
nor U7870 (N_7870,N_6526,N_6945);
nor U7871 (N_7871,N_6315,N_6574);
nor U7872 (N_7872,N_6773,N_6854);
and U7873 (N_7873,N_6283,N_6359);
nand U7874 (N_7874,N_6545,N_6785);
and U7875 (N_7875,N_6108,N_6114);
xnor U7876 (N_7876,N_6647,N_6136);
nor U7877 (N_7877,N_6743,N_6868);
and U7878 (N_7878,N_6518,N_6971);
nor U7879 (N_7879,N_6554,N_6420);
and U7880 (N_7880,N_6129,N_6451);
or U7881 (N_7881,N_6829,N_6206);
nand U7882 (N_7882,N_6953,N_6667);
and U7883 (N_7883,N_6793,N_6041);
and U7884 (N_7884,N_6705,N_6962);
nand U7885 (N_7885,N_6375,N_6047);
and U7886 (N_7886,N_6417,N_6321);
nor U7887 (N_7887,N_6570,N_6735);
and U7888 (N_7888,N_6408,N_6017);
or U7889 (N_7889,N_6158,N_6428);
or U7890 (N_7890,N_6507,N_6569);
or U7891 (N_7891,N_6863,N_6982);
or U7892 (N_7892,N_6648,N_6101);
nand U7893 (N_7893,N_6307,N_6185);
and U7894 (N_7894,N_6000,N_6578);
or U7895 (N_7895,N_6215,N_6306);
nor U7896 (N_7896,N_6489,N_6160);
and U7897 (N_7897,N_6411,N_6384);
nand U7898 (N_7898,N_6440,N_6318);
nor U7899 (N_7899,N_6867,N_6870);
nand U7900 (N_7900,N_6561,N_6718);
nand U7901 (N_7901,N_6812,N_6766);
nand U7902 (N_7902,N_6685,N_6935);
and U7903 (N_7903,N_6927,N_6690);
nand U7904 (N_7904,N_6441,N_6597);
or U7905 (N_7905,N_6530,N_6965);
nand U7906 (N_7906,N_6549,N_6682);
nor U7907 (N_7907,N_6337,N_6808);
nor U7908 (N_7908,N_6214,N_6676);
and U7909 (N_7909,N_6307,N_6177);
and U7910 (N_7910,N_6481,N_6828);
and U7911 (N_7911,N_6089,N_6895);
nand U7912 (N_7912,N_6298,N_6082);
and U7913 (N_7913,N_6638,N_6147);
and U7914 (N_7914,N_6939,N_6189);
nand U7915 (N_7915,N_6770,N_6827);
or U7916 (N_7916,N_6202,N_6187);
or U7917 (N_7917,N_6498,N_6389);
nand U7918 (N_7918,N_6736,N_6978);
or U7919 (N_7919,N_6525,N_6661);
and U7920 (N_7920,N_6229,N_6648);
or U7921 (N_7921,N_6402,N_6368);
nand U7922 (N_7922,N_6689,N_6994);
nand U7923 (N_7923,N_6595,N_6213);
nor U7924 (N_7924,N_6244,N_6918);
and U7925 (N_7925,N_6559,N_6090);
nor U7926 (N_7926,N_6971,N_6007);
nand U7927 (N_7927,N_6520,N_6262);
nor U7928 (N_7928,N_6945,N_6391);
and U7929 (N_7929,N_6606,N_6393);
or U7930 (N_7930,N_6014,N_6947);
and U7931 (N_7931,N_6234,N_6212);
nor U7932 (N_7932,N_6814,N_6201);
or U7933 (N_7933,N_6523,N_6605);
or U7934 (N_7934,N_6106,N_6686);
and U7935 (N_7935,N_6365,N_6087);
or U7936 (N_7936,N_6522,N_6789);
nor U7937 (N_7937,N_6845,N_6929);
nor U7938 (N_7938,N_6696,N_6248);
or U7939 (N_7939,N_6206,N_6651);
and U7940 (N_7940,N_6636,N_6017);
and U7941 (N_7941,N_6088,N_6822);
or U7942 (N_7942,N_6157,N_6446);
nand U7943 (N_7943,N_6183,N_6967);
or U7944 (N_7944,N_6135,N_6944);
or U7945 (N_7945,N_6089,N_6505);
or U7946 (N_7946,N_6545,N_6806);
and U7947 (N_7947,N_6066,N_6036);
or U7948 (N_7948,N_6969,N_6350);
nand U7949 (N_7949,N_6855,N_6703);
and U7950 (N_7950,N_6841,N_6736);
nand U7951 (N_7951,N_6438,N_6451);
nor U7952 (N_7952,N_6742,N_6848);
nand U7953 (N_7953,N_6016,N_6360);
nand U7954 (N_7954,N_6550,N_6245);
and U7955 (N_7955,N_6626,N_6020);
and U7956 (N_7956,N_6628,N_6788);
and U7957 (N_7957,N_6392,N_6510);
nor U7958 (N_7958,N_6403,N_6749);
or U7959 (N_7959,N_6239,N_6186);
nor U7960 (N_7960,N_6408,N_6368);
nand U7961 (N_7961,N_6756,N_6884);
nand U7962 (N_7962,N_6466,N_6120);
nand U7963 (N_7963,N_6272,N_6427);
or U7964 (N_7964,N_6283,N_6167);
nand U7965 (N_7965,N_6248,N_6018);
and U7966 (N_7966,N_6643,N_6491);
or U7967 (N_7967,N_6676,N_6373);
and U7968 (N_7968,N_6857,N_6136);
and U7969 (N_7969,N_6240,N_6755);
nand U7970 (N_7970,N_6668,N_6832);
nand U7971 (N_7971,N_6410,N_6247);
nor U7972 (N_7972,N_6194,N_6289);
and U7973 (N_7973,N_6831,N_6463);
nand U7974 (N_7974,N_6727,N_6648);
or U7975 (N_7975,N_6826,N_6736);
or U7976 (N_7976,N_6919,N_6766);
and U7977 (N_7977,N_6680,N_6863);
nor U7978 (N_7978,N_6149,N_6598);
or U7979 (N_7979,N_6911,N_6668);
or U7980 (N_7980,N_6938,N_6388);
nor U7981 (N_7981,N_6754,N_6193);
nand U7982 (N_7982,N_6915,N_6487);
nor U7983 (N_7983,N_6837,N_6689);
nor U7984 (N_7984,N_6448,N_6417);
and U7985 (N_7985,N_6924,N_6005);
nor U7986 (N_7986,N_6132,N_6184);
and U7987 (N_7987,N_6038,N_6662);
and U7988 (N_7988,N_6562,N_6099);
nand U7989 (N_7989,N_6828,N_6327);
nand U7990 (N_7990,N_6685,N_6650);
or U7991 (N_7991,N_6293,N_6523);
and U7992 (N_7992,N_6143,N_6053);
nand U7993 (N_7993,N_6041,N_6357);
nand U7994 (N_7994,N_6329,N_6862);
or U7995 (N_7995,N_6954,N_6349);
nor U7996 (N_7996,N_6928,N_6691);
and U7997 (N_7997,N_6317,N_6185);
and U7998 (N_7998,N_6881,N_6202);
nor U7999 (N_7999,N_6330,N_6483);
and U8000 (N_8000,N_7827,N_7971);
or U8001 (N_8001,N_7941,N_7497);
nor U8002 (N_8002,N_7984,N_7522);
nand U8003 (N_8003,N_7189,N_7348);
or U8004 (N_8004,N_7669,N_7034);
or U8005 (N_8005,N_7548,N_7791);
xor U8006 (N_8006,N_7302,N_7944);
or U8007 (N_8007,N_7903,N_7778);
and U8008 (N_8008,N_7081,N_7428);
and U8009 (N_8009,N_7256,N_7082);
or U8010 (N_8010,N_7992,N_7575);
and U8011 (N_8011,N_7614,N_7319);
nand U8012 (N_8012,N_7580,N_7641);
and U8013 (N_8013,N_7261,N_7927);
nor U8014 (N_8014,N_7070,N_7433);
or U8015 (N_8015,N_7775,N_7111);
or U8016 (N_8016,N_7964,N_7481);
or U8017 (N_8017,N_7878,N_7719);
nor U8018 (N_8018,N_7464,N_7780);
and U8019 (N_8019,N_7829,N_7867);
and U8020 (N_8020,N_7200,N_7924);
and U8021 (N_8021,N_7417,N_7682);
nor U8022 (N_8022,N_7132,N_7917);
nand U8023 (N_8023,N_7840,N_7347);
or U8024 (N_8024,N_7698,N_7598);
nand U8025 (N_8025,N_7394,N_7247);
and U8026 (N_8026,N_7879,N_7241);
and U8027 (N_8027,N_7080,N_7385);
or U8028 (N_8028,N_7202,N_7744);
nand U8029 (N_8029,N_7540,N_7676);
or U8030 (N_8030,N_7337,N_7090);
and U8031 (N_8031,N_7317,N_7496);
nor U8032 (N_8032,N_7229,N_7190);
nor U8033 (N_8033,N_7864,N_7471);
nand U8034 (N_8034,N_7239,N_7215);
and U8035 (N_8035,N_7187,N_7456);
nand U8036 (N_8036,N_7527,N_7224);
nor U8037 (N_8037,N_7503,N_7830);
xnor U8038 (N_8038,N_7367,N_7923);
and U8039 (N_8039,N_7759,N_7774);
nor U8040 (N_8040,N_7168,N_7834);
and U8041 (N_8041,N_7591,N_7243);
nand U8042 (N_8042,N_7270,N_7896);
and U8043 (N_8043,N_7662,N_7194);
and U8044 (N_8044,N_7642,N_7113);
nand U8045 (N_8045,N_7566,N_7981);
and U8046 (N_8046,N_7913,N_7396);
nand U8047 (N_8047,N_7868,N_7426);
and U8048 (N_8048,N_7369,N_7005);
or U8049 (N_8049,N_7060,N_7521);
nand U8050 (N_8050,N_7326,N_7714);
nand U8051 (N_8051,N_7545,N_7926);
nand U8052 (N_8052,N_7483,N_7723);
nor U8053 (N_8053,N_7335,N_7966);
nand U8054 (N_8054,N_7116,N_7814);
xnor U8055 (N_8055,N_7680,N_7089);
and U8056 (N_8056,N_7399,N_7360);
and U8057 (N_8057,N_7942,N_7516);
nor U8058 (N_8058,N_7318,N_7502);
nor U8059 (N_8059,N_7079,N_7799);
and U8060 (N_8060,N_7467,N_7782);
nand U8061 (N_8061,N_7169,N_7510);
nor U8062 (N_8062,N_7210,N_7410);
and U8063 (N_8063,N_7870,N_7478);
or U8064 (N_8064,N_7253,N_7732);
nand U8065 (N_8065,N_7010,N_7085);
or U8066 (N_8066,N_7972,N_7710);
or U8067 (N_8067,N_7826,N_7582);
and U8068 (N_8068,N_7308,N_7574);
or U8069 (N_8069,N_7726,N_7486);
nand U8070 (N_8070,N_7852,N_7245);
and U8071 (N_8071,N_7407,N_7693);
or U8072 (N_8072,N_7636,N_7570);
or U8073 (N_8073,N_7706,N_7024);
and U8074 (N_8074,N_7003,N_7828);
and U8075 (N_8075,N_7760,N_7841);
and U8076 (N_8076,N_7259,N_7808);
or U8077 (N_8077,N_7011,N_7249);
nand U8078 (N_8078,N_7139,N_7894);
or U8079 (N_8079,N_7753,N_7821);
or U8080 (N_8080,N_7498,N_7620);
and U8081 (N_8081,N_7431,N_7621);
or U8082 (N_8082,N_7465,N_7217);
nor U8083 (N_8083,N_7793,N_7763);
and U8084 (N_8084,N_7655,N_7755);
nor U8085 (N_8085,N_7400,N_7017);
nor U8086 (N_8086,N_7551,N_7330);
nand U8087 (N_8087,N_7746,N_7846);
or U8088 (N_8088,N_7482,N_7576);
or U8089 (N_8089,N_7520,N_7262);
or U8090 (N_8090,N_7184,N_7271);
nor U8091 (N_8091,N_7833,N_7815);
nand U8092 (N_8092,N_7051,N_7750);
nand U8093 (N_8093,N_7383,N_7543);
or U8094 (N_8094,N_7938,N_7107);
or U8095 (N_8095,N_7544,N_7386);
or U8096 (N_8096,N_7356,N_7102);
or U8097 (N_8097,N_7052,N_7514);
and U8098 (N_8098,N_7050,N_7104);
xnor U8099 (N_8099,N_7951,N_7606);
nand U8100 (N_8100,N_7579,N_7742);
nor U8101 (N_8101,N_7766,N_7473);
nor U8102 (N_8102,N_7556,N_7121);
and U8103 (N_8103,N_7268,N_7059);
or U8104 (N_8104,N_7028,N_7488);
and U8105 (N_8105,N_7316,N_7862);
nor U8106 (N_8106,N_7398,N_7860);
and U8107 (N_8107,N_7062,N_7092);
or U8108 (N_8108,N_7629,N_7696);
and U8109 (N_8109,N_7097,N_7390);
or U8110 (N_8110,N_7295,N_7177);
and U8111 (N_8111,N_7962,N_7118);
or U8112 (N_8112,N_7743,N_7352);
nor U8113 (N_8113,N_7195,N_7920);
nor U8114 (N_8114,N_7199,N_7949);
nand U8115 (N_8115,N_7203,N_7622);
nand U8116 (N_8116,N_7336,N_7320);
nor U8117 (N_8117,N_7847,N_7688);
nand U8118 (N_8118,N_7016,N_7979);
nand U8119 (N_8119,N_7954,N_7929);
nand U8120 (N_8120,N_7258,N_7376);
and U8121 (N_8121,N_7162,N_7377);
and U8122 (N_8122,N_7493,N_7880);
nor U8123 (N_8123,N_7310,N_7648);
and U8124 (N_8124,N_7930,N_7154);
nor U8125 (N_8125,N_7067,N_7875);
xnor U8126 (N_8126,N_7305,N_7240);
or U8127 (N_8127,N_7188,N_7466);
nor U8128 (N_8128,N_7468,N_7266);
nor U8129 (N_8129,N_7301,N_7639);
or U8130 (N_8130,N_7722,N_7299);
nand U8131 (N_8131,N_7842,N_7569);
nand U8132 (N_8132,N_7207,N_7150);
and U8133 (N_8133,N_7366,N_7756);
nor U8134 (N_8134,N_7103,N_7100);
nor U8135 (N_8135,N_7687,N_7141);
and U8136 (N_8136,N_7858,N_7106);
nor U8137 (N_8137,N_7932,N_7147);
nand U8138 (N_8138,N_7739,N_7487);
and U8139 (N_8139,N_7006,N_7234);
and U8140 (N_8140,N_7430,N_7695);
nor U8141 (N_8141,N_7991,N_7233);
or U8142 (N_8142,N_7853,N_7748);
or U8143 (N_8143,N_7128,N_7015);
nand U8144 (N_8144,N_7654,N_7174);
and U8145 (N_8145,N_7115,N_7628);
and U8146 (N_8146,N_7382,N_7123);
or U8147 (N_8147,N_7599,N_7442);
nand U8148 (N_8148,N_7035,N_7044);
nor U8149 (N_8149,N_7735,N_7640);
and U8150 (N_8150,N_7345,N_7952);
nand U8151 (N_8151,N_7637,N_7851);
or U8152 (N_8152,N_7577,N_7267);
and U8153 (N_8153,N_7029,N_7443);
nand U8154 (N_8154,N_7083,N_7357);
or U8155 (N_8155,N_7624,N_7623);
nor U8156 (N_8156,N_7532,N_7076);
nand U8157 (N_8157,N_7323,N_7408);
nand U8158 (N_8158,N_7149,N_7908);
nand U8159 (N_8159,N_7046,N_7988);
and U8160 (N_8160,N_7573,N_7800);
and U8161 (N_8161,N_7156,N_7402);
nor U8162 (N_8162,N_7368,N_7789);
and U8163 (N_8163,N_7562,N_7039);
nor U8164 (N_8164,N_7186,N_7762);
and U8165 (N_8165,N_7429,N_7893);
nor U8166 (N_8166,N_7772,N_7959);
and U8167 (N_8167,N_7370,N_7284);
nand U8168 (N_8168,N_7511,N_7794);
or U8169 (N_8169,N_7831,N_7453);
and U8170 (N_8170,N_7697,N_7343);
nor U8171 (N_8171,N_7304,N_7470);
nand U8172 (N_8172,N_7474,N_7086);
nand U8173 (N_8173,N_7885,N_7379);
nand U8174 (N_8174,N_7146,N_7784);
and U8175 (N_8175,N_7170,N_7524);
nand U8176 (N_8176,N_7578,N_7990);
or U8177 (N_8177,N_7823,N_7296);
and U8178 (N_8178,N_7285,N_7649);
or U8179 (N_8179,N_7022,N_7530);
or U8180 (N_8180,N_7440,N_7138);
nand U8181 (N_8181,N_7110,N_7288);
or U8182 (N_8182,N_7825,N_7886);
nand U8183 (N_8183,N_7925,N_7228);
nor U8184 (N_8184,N_7197,N_7978);
nand U8185 (N_8185,N_7378,N_7593);
or U8186 (N_8186,N_7069,N_7631);
nand U8187 (N_8187,N_7179,N_7787);
nor U8188 (N_8188,N_7372,N_7279);
and U8189 (N_8189,N_7164,N_7718);
nor U8190 (N_8190,N_7071,N_7950);
nor U8191 (N_8191,N_7845,N_7321);
and U8192 (N_8192,N_7617,N_7445);
or U8193 (N_8193,N_7452,N_7209);
nand U8194 (N_8194,N_7987,N_7747);
nand U8195 (N_8195,N_7447,N_7127);
nor U8196 (N_8196,N_7122,N_7955);
xnor U8197 (N_8197,N_7341,N_7713);
nor U8198 (N_8198,N_7283,N_7061);
or U8199 (N_8199,N_7246,N_7012);
and U8200 (N_8200,N_7707,N_7176);
nand U8201 (N_8201,N_7685,N_7783);
nor U8202 (N_8202,N_7597,N_7692);
or U8203 (N_8203,N_7008,N_7387);
nor U8204 (N_8204,N_7507,N_7651);
nand U8205 (N_8205,N_7644,N_7235);
or U8206 (N_8206,N_7451,N_7126);
nand U8207 (N_8207,N_7178,N_7415);
xor U8208 (N_8208,N_7472,N_7983);
nor U8209 (N_8209,N_7004,N_7725);
or U8210 (N_8210,N_7792,N_7492);
nor U8211 (N_8211,N_7460,N_7583);
nor U8212 (N_8212,N_7250,N_7358);
nand U8213 (N_8213,N_7094,N_7222);
nor U8214 (N_8214,N_7822,N_7936);
nand U8215 (N_8215,N_7934,N_7095);
nand U8216 (N_8216,N_7537,N_7663);
or U8217 (N_8217,N_7084,N_7119);
nand U8218 (N_8218,N_7730,N_7171);
nor U8219 (N_8219,N_7741,N_7324);
nor U8220 (N_8220,N_7869,N_7907);
and U8221 (N_8221,N_7584,N_7334);
nand U8222 (N_8222,N_7811,N_7674);
nor U8223 (N_8223,N_7679,N_7489);
and U8224 (N_8224,N_7018,N_7838);
or U8225 (N_8225,N_7340,N_7329);
nand U8226 (N_8226,N_7594,N_7785);
xnor U8227 (N_8227,N_7940,N_7225);
nor U8228 (N_8228,N_7384,N_7957);
and U8229 (N_8229,N_7803,N_7736);
and U8230 (N_8230,N_7098,N_7626);
nor U8231 (N_8231,N_7269,N_7715);
nor U8232 (N_8232,N_7088,N_7419);
nor U8233 (N_8233,N_7767,N_7625);
and U8234 (N_8234,N_7604,N_7975);
nand U8235 (N_8235,N_7839,N_7423);
or U8236 (N_8236,N_7563,N_7422);
nor U8237 (N_8237,N_7668,N_7727);
and U8238 (N_8238,N_7255,N_7882);
nand U8239 (N_8239,N_7592,N_7708);
nor U8240 (N_8240,N_7533,N_7916);
and U8241 (N_8241,N_7559,N_7133);
or U8242 (N_8242,N_7817,N_7509);
or U8243 (N_8243,N_7531,N_7884);
or U8244 (N_8244,N_7220,N_7777);
or U8245 (N_8245,N_7491,N_7998);
nor U8246 (N_8246,N_7557,N_7716);
and U8247 (N_8247,N_7657,N_7213);
or U8248 (N_8248,N_7776,N_7265);
nor U8249 (N_8249,N_7633,N_7684);
nor U8250 (N_8250,N_7993,N_7810);
nor U8251 (N_8251,N_7148,N_7311);
or U8252 (N_8252,N_7205,N_7325);
and U8253 (N_8253,N_7434,N_7589);
and U8254 (N_8254,N_7595,N_7131);
xnor U8255 (N_8255,N_7729,N_7538);
or U8256 (N_8256,N_7694,N_7105);
nand U8257 (N_8257,N_7395,N_7117);
nor U8258 (N_8258,N_7970,N_7292);
nand U8259 (N_8259,N_7182,N_7855);
and U8260 (N_8260,N_7495,N_7702);
nor U8261 (N_8261,N_7037,N_7602);
or U8262 (N_8262,N_7689,N_7137);
nor U8263 (N_8263,N_7192,N_7172);
and U8264 (N_8264,N_7824,N_7627);
nand U8265 (N_8265,N_7675,N_7152);
and U8266 (N_8266,N_7526,N_7036);
nand U8267 (N_8267,N_7032,N_7479);
nand U8268 (N_8268,N_7666,N_7953);
or U8269 (N_8269,N_7001,N_7312);
nor U8270 (N_8270,N_7346,N_7989);
nor U8271 (N_8271,N_7667,N_7159);
nor U8272 (N_8272,N_7596,N_7701);
nor U8273 (N_8273,N_7251,N_7534);
nor U8274 (N_8274,N_7307,N_7454);
and U8275 (N_8275,N_7281,N_7450);
nand U8276 (N_8276,N_7837,N_7500);
or U8277 (N_8277,N_7752,N_7705);
nand U8278 (N_8278,N_7091,N_7999);
or U8279 (N_8279,N_7153,N_7615);
or U8280 (N_8280,N_7731,N_7145);
or U8281 (N_8281,N_7699,N_7365);
or U8282 (N_8282,N_7173,N_7709);
nor U8283 (N_8283,N_7634,N_7891);
nor U8284 (N_8284,N_7077,N_7788);
or U8285 (N_8285,N_7931,N_7053);
and U8286 (N_8286,N_7065,N_7677);
and U8287 (N_8287,N_7733,N_7802);
nor U8288 (N_8288,N_7236,N_7529);
nand U8289 (N_8289,N_7055,N_7280);
or U8290 (N_8290,N_7818,N_7198);
and U8291 (N_8291,N_7000,N_7773);
nand U8292 (N_8292,N_7590,N_7298);
and U8293 (N_8293,N_7968,N_7294);
and U8294 (N_8294,N_7397,N_7919);
and U8295 (N_8295,N_7211,N_7734);
or U8296 (N_8296,N_7555,N_7751);
nand U8297 (N_8297,N_7322,N_7535);
nor U8298 (N_8298,N_7613,N_7135);
nor U8299 (N_8299,N_7045,N_7857);
nand U8300 (N_8300,N_7344,N_7260);
nor U8301 (N_8301,N_7561,N_7512);
or U8302 (N_8302,N_7448,N_7761);
and U8303 (N_8303,N_7638,N_7277);
and U8304 (N_8304,N_7165,N_7758);
nor U8305 (N_8305,N_7568,N_7175);
or U8306 (N_8306,N_7588,N_7911);
nor U8307 (N_8307,N_7519,N_7129);
and U8308 (N_8308,N_7796,N_7508);
nor U8309 (N_8309,N_7553,N_7373);
or U8310 (N_8310,N_7795,N_7994);
nor U8311 (N_8311,N_7063,N_7381);
or U8312 (N_8312,N_7947,N_7565);
nand U8313 (N_8313,N_7819,N_7158);
or U8314 (N_8314,N_7986,N_7338);
and U8315 (N_8315,N_7572,N_7567);
nand U8316 (N_8316,N_7401,N_7854);
or U8317 (N_8317,N_7303,N_7469);
nand U8318 (N_8318,N_7832,N_7193);
or U8319 (N_8319,N_7965,N_7518);
or U8320 (N_8320,N_7525,N_7242);
nand U8321 (N_8321,N_7887,N_7455);
nor U8322 (N_8322,N_7652,N_7900);
and U8323 (N_8323,N_7073,N_7134);
or U8324 (N_8324,N_7659,N_7672);
nor U8325 (N_8325,N_7608,N_7359);
or U8326 (N_8326,N_7112,N_7866);
and U8327 (N_8327,N_7485,N_7921);
nor U8328 (N_8328,N_7230,N_7332);
and U8329 (N_8329,N_7645,N_7363);
nand U8330 (N_8330,N_7350,N_7068);
and U8331 (N_8331,N_7915,N_7601);
nand U8332 (N_8332,N_7181,N_7391);
nor U8333 (N_8333,N_7309,N_7058);
or U8334 (N_8334,N_7995,N_7505);
nand U8335 (N_8335,N_7717,N_7700);
or U8336 (N_8336,N_7720,N_7208);
and U8337 (N_8337,N_7314,N_7124);
nand U8338 (N_8338,N_7013,N_7541);
nand U8339 (N_8339,N_7254,N_7064);
or U8340 (N_8340,N_7611,N_7937);
and U8341 (N_8341,N_7961,N_7724);
or U8342 (N_8342,N_7960,N_7874);
and U8343 (N_8343,N_7813,N_7221);
and U8344 (N_8344,N_7605,N_7361);
nand U8345 (N_8345,N_7420,N_7125);
and U8346 (N_8346,N_7779,N_7528);
or U8347 (N_8347,N_7997,N_7143);
and U8348 (N_8348,N_7843,N_7056);
nand U8349 (N_8349,N_7388,N_7586);
nor U8350 (N_8350,N_7109,N_7328);
nor U8351 (N_8351,N_7946,N_7413);
or U8352 (N_8352,N_7196,N_7754);
nand U8353 (N_8353,N_7002,N_7371);
nor U8354 (N_8354,N_7042,N_7740);
nand U8355 (N_8355,N_7339,N_7801);
nand U8356 (N_8356,N_7040,N_7030);
nand U8357 (N_8357,N_7290,N_7166);
and U8358 (N_8358,N_7928,N_7871);
nor U8359 (N_8359,N_7227,N_7272);
nor U8360 (N_8360,N_7093,N_7504);
nand U8361 (N_8361,N_7798,N_7151);
nand U8362 (N_8362,N_7216,N_7786);
nand U8363 (N_8363,N_7163,N_7665);
and U8364 (N_8364,N_7201,N_7996);
or U8365 (N_8365,N_7031,N_7041);
and U8366 (N_8366,N_7945,N_7416);
or U8367 (N_8367,N_7275,N_7905);
nand U8368 (N_8368,N_7764,N_7836);
nor U8369 (N_8369,N_7484,N_7405);
nand U8370 (N_8370,N_7252,N_7437);
and U8371 (N_8371,N_7120,N_7212);
and U8372 (N_8372,N_7411,N_7600);
nor U8373 (N_8373,N_7436,N_7691);
nand U8374 (N_8374,N_7412,N_7300);
nor U8375 (N_8375,N_7914,N_7231);
or U8376 (N_8376,N_7140,N_7043);
or U8377 (N_8377,N_7099,N_7237);
and U8378 (N_8378,N_7439,N_7306);
and U8379 (N_8379,N_7441,N_7546);
or U8380 (N_8380,N_7425,N_7155);
and U8381 (N_8381,N_7619,N_7681);
or U8382 (N_8382,N_7670,N_7297);
nor U8383 (N_8383,N_7342,N_7315);
nor U8384 (N_8384,N_7020,N_7585);
nand U8385 (N_8385,N_7671,N_7406);
and U8386 (N_8386,N_7806,N_7393);
nand U8387 (N_8387,N_7289,N_7797);
and U8388 (N_8388,N_7403,N_7844);
or U8389 (N_8389,N_7872,N_7895);
nand U8390 (N_8390,N_7282,N_7009);
nor U8391 (N_8391,N_7499,N_7849);
nand U8392 (N_8392,N_7523,N_7749);
or U8393 (N_8393,N_7087,N_7096);
nor U8394 (N_8394,N_7897,N_7144);
or U8395 (N_8395,N_7587,N_7809);
or U8396 (N_8396,N_7501,N_7618);
or U8397 (N_8397,N_7414,N_7912);
and U8398 (N_8398,N_7904,N_7883);
nor U8399 (N_8399,N_7835,N_7890);
or U8400 (N_8400,N_7812,N_7075);
nand U8401 (N_8401,N_7554,N_7223);
nor U8402 (N_8402,N_7160,N_7157);
or U8403 (N_8403,N_7049,N_7603);
nand U8404 (N_8404,N_7038,N_7130);
and U8405 (N_8405,N_7982,N_7683);
nand U8406 (N_8406,N_7446,N_7257);
nor U8407 (N_8407,N_7418,N_7461);
nor U8408 (N_8408,N_7161,N_7805);
or U8409 (N_8409,N_7362,N_7673);
or U8410 (N_8410,N_7313,N_7048);
nor U8411 (N_8411,N_7985,N_7459);
nor U8412 (N_8412,N_7770,N_7191);
nand U8413 (N_8413,N_7630,N_7392);
nor U8414 (N_8414,N_7263,N_7581);
nand U8415 (N_8415,N_7935,N_7078);
nand U8416 (N_8416,N_7517,N_7737);
or U8417 (N_8417,N_7542,N_7274);
nor U8418 (N_8418,N_7771,N_7910);
nand U8419 (N_8419,N_7876,N_7204);
nor U8420 (N_8420,N_7948,N_7494);
xnor U8421 (N_8421,N_7327,N_7353);
or U8422 (N_8422,N_7476,N_7656);
and U8423 (N_8423,N_7550,N_7881);
or U8424 (N_8424,N_7276,N_7026);
nand U8425 (N_8425,N_7536,N_7007);
nor U8426 (N_8426,N_7404,N_7539);
and U8427 (N_8427,N_7552,N_7114);
nor U8428 (N_8428,N_7607,N_7856);
or U8429 (N_8429,N_7653,N_7444);
or U8430 (N_8430,N_7980,N_7850);
nor U8431 (N_8431,N_7865,N_7728);
or U8432 (N_8432,N_7609,N_7790);
nand U8433 (N_8433,N_7477,N_7349);
and U8434 (N_8434,N_7214,N_7977);
nor U8435 (N_8435,N_7909,N_7650);
nand U8436 (N_8436,N_7863,N_7976);
and U8437 (N_8437,N_7351,N_7054);
nand U8438 (N_8438,N_7635,N_7218);
and U8439 (N_8439,N_7969,N_7183);
or U8440 (N_8440,N_7380,N_7560);
and U8441 (N_8441,N_7902,N_7421);
or U8442 (N_8442,N_7974,N_7463);
nand U8443 (N_8443,N_7564,N_7027);
nand U8444 (N_8444,N_7506,N_7632);
nand U8445 (N_8445,N_7232,N_7264);
nor U8446 (N_8446,N_7973,N_7244);
or U8447 (N_8447,N_7820,N_7690);
or U8448 (N_8448,N_7807,N_7859);
nor U8449 (N_8449,N_7286,N_7355);
nand U8450 (N_8450,N_7888,N_7738);
or U8451 (N_8451,N_7047,N_7658);
nand U8452 (N_8452,N_7704,N_7816);
nand U8453 (N_8453,N_7374,N_7956);
or U8454 (N_8454,N_7021,N_7432);
and U8455 (N_8455,N_7331,N_7848);
or U8456 (N_8456,N_7333,N_7643);
and U8457 (N_8457,N_7206,N_7646);
nor U8458 (N_8458,N_7057,N_7547);
nor U8459 (N_8459,N_7427,N_7515);
nor U8460 (N_8460,N_7967,N_7804);
or U8461 (N_8461,N_7661,N_7072);
or U8462 (N_8462,N_7943,N_7712);
nor U8463 (N_8463,N_7023,N_7906);
nor U8464 (N_8464,N_7703,N_7475);
nand U8465 (N_8465,N_7449,N_7273);
and U8466 (N_8466,N_7745,N_7480);
and U8467 (N_8467,N_7889,N_7033);
or U8468 (N_8468,N_7901,N_7074);
and U8469 (N_8469,N_7757,N_7877);
and U8470 (N_8470,N_7616,N_7678);
and U8471 (N_8471,N_7108,N_7424);
or U8472 (N_8472,N_7101,N_7219);
and U8473 (N_8473,N_7892,N_7765);
nand U8474 (N_8474,N_7409,N_7612);
nand U8475 (N_8475,N_7167,N_7293);
and U8476 (N_8476,N_7610,N_7066);
nor U8477 (N_8477,N_7549,N_7458);
and U8478 (N_8478,N_7873,N_7185);
xnor U8479 (N_8479,N_7922,N_7958);
nor U8480 (N_8480,N_7457,N_7899);
and U8481 (N_8481,N_7918,N_7933);
nor U8482 (N_8482,N_7019,N_7861);
nand U8483 (N_8483,N_7462,N_7238);
nor U8484 (N_8484,N_7664,N_7136);
and U8485 (N_8485,N_7248,N_7389);
nor U8486 (N_8486,N_7025,N_7438);
or U8487 (N_8487,N_7014,N_7647);
nand U8488 (N_8488,N_7768,N_7291);
and U8489 (N_8489,N_7963,N_7435);
nand U8490 (N_8490,N_7721,N_7287);
nand U8491 (N_8491,N_7781,N_7278);
nor U8492 (N_8492,N_7898,N_7180);
nor U8493 (N_8493,N_7354,N_7660);
nor U8494 (N_8494,N_7939,N_7142);
and U8495 (N_8495,N_7571,N_7375);
nand U8496 (N_8496,N_7711,N_7490);
or U8497 (N_8497,N_7686,N_7364);
and U8498 (N_8498,N_7513,N_7558);
nor U8499 (N_8499,N_7226,N_7769);
xor U8500 (N_8500,N_7570,N_7297);
nor U8501 (N_8501,N_7329,N_7360);
nor U8502 (N_8502,N_7865,N_7188);
nor U8503 (N_8503,N_7189,N_7022);
or U8504 (N_8504,N_7352,N_7171);
nor U8505 (N_8505,N_7037,N_7430);
nor U8506 (N_8506,N_7030,N_7693);
nor U8507 (N_8507,N_7540,N_7651);
and U8508 (N_8508,N_7488,N_7588);
nor U8509 (N_8509,N_7493,N_7634);
nand U8510 (N_8510,N_7794,N_7509);
or U8511 (N_8511,N_7011,N_7821);
and U8512 (N_8512,N_7566,N_7539);
and U8513 (N_8513,N_7537,N_7214);
nand U8514 (N_8514,N_7821,N_7690);
or U8515 (N_8515,N_7041,N_7952);
and U8516 (N_8516,N_7119,N_7528);
nand U8517 (N_8517,N_7593,N_7715);
and U8518 (N_8518,N_7810,N_7890);
or U8519 (N_8519,N_7132,N_7695);
or U8520 (N_8520,N_7184,N_7179);
nor U8521 (N_8521,N_7224,N_7700);
nor U8522 (N_8522,N_7381,N_7541);
nor U8523 (N_8523,N_7062,N_7225);
nand U8524 (N_8524,N_7282,N_7092);
nand U8525 (N_8525,N_7480,N_7380);
nand U8526 (N_8526,N_7541,N_7868);
xor U8527 (N_8527,N_7512,N_7353);
nor U8528 (N_8528,N_7628,N_7307);
and U8529 (N_8529,N_7883,N_7813);
or U8530 (N_8530,N_7334,N_7603);
or U8531 (N_8531,N_7130,N_7309);
nor U8532 (N_8532,N_7290,N_7057);
or U8533 (N_8533,N_7175,N_7015);
nand U8534 (N_8534,N_7730,N_7785);
nor U8535 (N_8535,N_7119,N_7258);
nor U8536 (N_8536,N_7101,N_7213);
nor U8537 (N_8537,N_7362,N_7818);
xor U8538 (N_8538,N_7813,N_7845);
nand U8539 (N_8539,N_7152,N_7305);
nor U8540 (N_8540,N_7379,N_7682);
or U8541 (N_8541,N_7887,N_7277);
or U8542 (N_8542,N_7599,N_7586);
xnor U8543 (N_8543,N_7032,N_7012);
or U8544 (N_8544,N_7976,N_7721);
or U8545 (N_8545,N_7794,N_7681);
nand U8546 (N_8546,N_7873,N_7897);
nand U8547 (N_8547,N_7018,N_7082);
and U8548 (N_8548,N_7234,N_7466);
or U8549 (N_8549,N_7465,N_7764);
nor U8550 (N_8550,N_7831,N_7615);
and U8551 (N_8551,N_7300,N_7522);
and U8552 (N_8552,N_7844,N_7078);
and U8553 (N_8553,N_7425,N_7641);
and U8554 (N_8554,N_7469,N_7232);
or U8555 (N_8555,N_7396,N_7276);
nor U8556 (N_8556,N_7850,N_7482);
and U8557 (N_8557,N_7012,N_7581);
and U8558 (N_8558,N_7106,N_7614);
or U8559 (N_8559,N_7841,N_7123);
or U8560 (N_8560,N_7965,N_7943);
or U8561 (N_8561,N_7293,N_7562);
or U8562 (N_8562,N_7652,N_7751);
and U8563 (N_8563,N_7309,N_7742);
and U8564 (N_8564,N_7427,N_7552);
nor U8565 (N_8565,N_7911,N_7450);
and U8566 (N_8566,N_7174,N_7506);
or U8567 (N_8567,N_7993,N_7905);
nor U8568 (N_8568,N_7006,N_7801);
or U8569 (N_8569,N_7518,N_7609);
and U8570 (N_8570,N_7921,N_7266);
or U8571 (N_8571,N_7800,N_7655);
or U8572 (N_8572,N_7751,N_7451);
nand U8573 (N_8573,N_7175,N_7713);
and U8574 (N_8574,N_7362,N_7393);
and U8575 (N_8575,N_7259,N_7512);
or U8576 (N_8576,N_7804,N_7798);
and U8577 (N_8577,N_7016,N_7148);
xor U8578 (N_8578,N_7851,N_7267);
nor U8579 (N_8579,N_7965,N_7162);
or U8580 (N_8580,N_7282,N_7209);
nor U8581 (N_8581,N_7257,N_7730);
nand U8582 (N_8582,N_7719,N_7908);
or U8583 (N_8583,N_7275,N_7282);
nor U8584 (N_8584,N_7110,N_7603);
xor U8585 (N_8585,N_7505,N_7949);
nor U8586 (N_8586,N_7946,N_7652);
or U8587 (N_8587,N_7451,N_7013);
and U8588 (N_8588,N_7892,N_7195);
and U8589 (N_8589,N_7445,N_7443);
or U8590 (N_8590,N_7546,N_7681);
and U8591 (N_8591,N_7250,N_7385);
nor U8592 (N_8592,N_7503,N_7430);
nor U8593 (N_8593,N_7980,N_7522);
nand U8594 (N_8594,N_7494,N_7832);
or U8595 (N_8595,N_7988,N_7549);
nand U8596 (N_8596,N_7681,N_7187);
nand U8597 (N_8597,N_7404,N_7375);
nand U8598 (N_8598,N_7162,N_7217);
nand U8599 (N_8599,N_7183,N_7099);
nand U8600 (N_8600,N_7042,N_7885);
or U8601 (N_8601,N_7541,N_7339);
nor U8602 (N_8602,N_7139,N_7740);
nand U8603 (N_8603,N_7485,N_7793);
and U8604 (N_8604,N_7461,N_7644);
nand U8605 (N_8605,N_7998,N_7826);
nand U8606 (N_8606,N_7332,N_7870);
and U8607 (N_8607,N_7654,N_7187);
nand U8608 (N_8608,N_7953,N_7182);
nand U8609 (N_8609,N_7661,N_7870);
xnor U8610 (N_8610,N_7534,N_7739);
nor U8611 (N_8611,N_7213,N_7195);
and U8612 (N_8612,N_7823,N_7648);
nor U8613 (N_8613,N_7443,N_7104);
or U8614 (N_8614,N_7493,N_7284);
nand U8615 (N_8615,N_7575,N_7143);
nand U8616 (N_8616,N_7605,N_7292);
and U8617 (N_8617,N_7789,N_7487);
and U8618 (N_8618,N_7297,N_7846);
or U8619 (N_8619,N_7694,N_7041);
nand U8620 (N_8620,N_7360,N_7657);
nand U8621 (N_8621,N_7406,N_7923);
or U8622 (N_8622,N_7833,N_7720);
or U8623 (N_8623,N_7137,N_7826);
or U8624 (N_8624,N_7460,N_7382);
nand U8625 (N_8625,N_7228,N_7631);
nor U8626 (N_8626,N_7317,N_7764);
nand U8627 (N_8627,N_7922,N_7753);
and U8628 (N_8628,N_7359,N_7066);
nand U8629 (N_8629,N_7432,N_7927);
or U8630 (N_8630,N_7586,N_7681);
and U8631 (N_8631,N_7461,N_7610);
xor U8632 (N_8632,N_7196,N_7809);
or U8633 (N_8633,N_7329,N_7153);
nand U8634 (N_8634,N_7370,N_7631);
nand U8635 (N_8635,N_7684,N_7751);
or U8636 (N_8636,N_7570,N_7994);
nand U8637 (N_8637,N_7749,N_7527);
or U8638 (N_8638,N_7406,N_7435);
and U8639 (N_8639,N_7145,N_7426);
nand U8640 (N_8640,N_7953,N_7306);
nor U8641 (N_8641,N_7970,N_7950);
and U8642 (N_8642,N_7895,N_7298);
nor U8643 (N_8643,N_7854,N_7621);
nor U8644 (N_8644,N_7789,N_7938);
and U8645 (N_8645,N_7142,N_7474);
or U8646 (N_8646,N_7665,N_7482);
nor U8647 (N_8647,N_7131,N_7845);
nor U8648 (N_8648,N_7414,N_7014);
or U8649 (N_8649,N_7826,N_7277);
and U8650 (N_8650,N_7012,N_7759);
nor U8651 (N_8651,N_7170,N_7971);
and U8652 (N_8652,N_7771,N_7646);
nand U8653 (N_8653,N_7456,N_7198);
and U8654 (N_8654,N_7490,N_7599);
or U8655 (N_8655,N_7010,N_7331);
and U8656 (N_8656,N_7690,N_7303);
nor U8657 (N_8657,N_7956,N_7690);
or U8658 (N_8658,N_7903,N_7234);
nor U8659 (N_8659,N_7600,N_7159);
and U8660 (N_8660,N_7694,N_7964);
nand U8661 (N_8661,N_7887,N_7722);
and U8662 (N_8662,N_7965,N_7517);
nand U8663 (N_8663,N_7657,N_7601);
or U8664 (N_8664,N_7371,N_7006);
nor U8665 (N_8665,N_7202,N_7934);
and U8666 (N_8666,N_7279,N_7499);
or U8667 (N_8667,N_7472,N_7829);
nand U8668 (N_8668,N_7039,N_7587);
xor U8669 (N_8669,N_7184,N_7174);
or U8670 (N_8670,N_7900,N_7651);
and U8671 (N_8671,N_7266,N_7403);
xor U8672 (N_8672,N_7807,N_7060);
and U8673 (N_8673,N_7677,N_7176);
and U8674 (N_8674,N_7923,N_7735);
nand U8675 (N_8675,N_7207,N_7136);
nor U8676 (N_8676,N_7283,N_7521);
nand U8677 (N_8677,N_7603,N_7830);
nand U8678 (N_8678,N_7076,N_7603);
nor U8679 (N_8679,N_7447,N_7639);
and U8680 (N_8680,N_7502,N_7669);
or U8681 (N_8681,N_7097,N_7354);
or U8682 (N_8682,N_7453,N_7500);
nor U8683 (N_8683,N_7970,N_7891);
or U8684 (N_8684,N_7378,N_7995);
nand U8685 (N_8685,N_7662,N_7786);
and U8686 (N_8686,N_7492,N_7015);
and U8687 (N_8687,N_7646,N_7663);
nor U8688 (N_8688,N_7550,N_7087);
xor U8689 (N_8689,N_7794,N_7354);
nand U8690 (N_8690,N_7717,N_7007);
and U8691 (N_8691,N_7053,N_7279);
and U8692 (N_8692,N_7741,N_7023);
or U8693 (N_8693,N_7903,N_7398);
and U8694 (N_8694,N_7195,N_7557);
nand U8695 (N_8695,N_7764,N_7840);
nand U8696 (N_8696,N_7202,N_7144);
nor U8697 (N_8697,N_7460,N_7631);
nand U8698 (N_8698,N_7446,N_7090);
or U8699 (N_8699,N_7367,N_7723);
nor U8700 (N_8700,N_7980,N_7391);
and U8701 (N_8701,N_7468,N_7616);
nor U8702 (N_8702,N_7987,N_7348);
nor U8703 (N_8703,N_7592,N_7140);
or U8704 (N_8704,N_7193,N_7370);
or U8705 (N_8705,N_7846,N_7176);
nor U8706 (N_8706,N_7760,N_7754);
or U8707 (N_8707,N_7434,N_7779);
nand U8708 (N_8708,N_7696,N_7321);
and U8709 (N_8709,N_7283,N_7838);
or U8710 (N_8710,N_7696,N_7035);
and U8711 (N_8711,N_7905,N_7843);
or U8712 (N_8712,N_7149,N_7854);
nand U8713 (N_8713,N_7670,N_7879);
nor U8714 (N_8714,N_7966,N_7823);
or U8715 (N_8715,N_7091,N_7246);
or U8716 (N_8716,N_7505,N_7245);
nand U8717 (N_8717,N_7056,N_7786);
nor U8718 (N_8718,N_7705,N_7042);
or U8719 (N_8719,N_7026,N_7514);
nand U8720 (N_8720,N_7062,N_7967);
nand U8721 (N_8721,N_7190,N_7012);
nand U8722 (N_8722,N_7983,N_7200);
and U8723 (N_8723,N_7065,N_7597);
and U8724 (N_8724,N_7482,N_7692);
or U8725 (N_8725,N_7888,N_7628);
and U8726 (N_8726,N_7163,N_7088);
or U8727 (N_8727,N_7487,N_7840);
nor U8728 (N_8728,N_7834,N_7996);
nand U8729 (N_8729,N_7953,N_7248);
or U8730 (N_8730,N_7504,N_7112);
nand U8731 (N_8731,N_7915,N_7059);
and U8732 (N_8732,N_7342,N_7012);
and U8733 (N_8733,N_7809,N_7618);
or U8734 (N_8734,N_7062,N_7016);
nand U8735 (N_8735,N_7263,N_7315);
or U8736 (N_8736,N_7628,N_7759);
and U8737 (N_8737,N_7691,N_7021);
or U8738 (N_8738,N_7005,N_7929);
xnor U8739 (N_8739,N_7775,N_7458);
nor U8740 (N_8740,N_7085,N_7176);
or U8741 (N_8741,N_7760,N_7925);
and U8742 (N_8742,N_7233,N_7957);
nand U8743 (N_8743,N_7267,N_7273);
and U8744 (N_8744,N_7677,N_7208);
nor U8745 (N_8745,N_7446,N_7625);
and U8746 (N_8746,N_7952,N_7506);
nand U8747 (N_8747,N_7468,N_7472);
or U8748 (N_8748,N_7595,N_7635);
and U8749 (N_8749,N_7465,N_7584);
and U8750 (N_8750,N_7768,N_7131);
nor U8751 (N_8751,N_7195,N_7705);
or U8752 (N_8752,N_7406,N_7162);
or U8753 (N_8753,N_7264,N_7792);
or U8754 (N_8754,N_7439,N_7541);
and U8755 (N_8755,N_7786,N_7420);
and U8756 (N_8756,N_7296,N_7562);
nor U8757 (N_8757,N_7441,N_7751);
xnor U8758 (N_8758,N_7239,N_7934);
nor U8759 (N_8759,N_7577,N_7005);
nor U8760 (N_8760,N_7725,N_7977);
or U8761 (N_8761,N_7985,N_7192);
nand U8762 (N_8762,N_7363,N_7275);
and U8763 (N_8763,N_7122,N_7847);
nor U8764 (N_8764,N_7777,N_7461);
nand U8765 (N_8765,N_7437,N_7143);
and U8766 (N_8766,N_7472,N_7553);
and U8767 (N_8767,N_7802,N_7046);
nor U8768 (N_8768,N_7103,N_7204);
nand U8769 (N_8769,N_7604,N_7101);
nand U8770 (N_8770,N_7046,N_7529);
or U8771 (N_8771,N_7709,N_7158);
nor U8772 (N_8772,N_7495,N_7083);
and U8773 (N_8773,N_7126,N_7006);
nor U8774 (N_8774,N_7527,N_7663);
and U8775 (N_8775,N_7366,N_7079);
nor U8776 (N_8776,N_7257,N_7483);
xor U8777 (N_8777,N_7670,N_7454);
and U8778 (N_8778,N_7776,N_7488);
nand U8779 (N_8779,N_7315,N_7656);
or U8780 (N_8780,N_7731,N_7250);
or U8781 (N_8781,N_7937,N_7332);
or U8782 (N_8782,N_7147,N_7037);
nand U8783 (N_8783,N_7960,N_7636);
nand U8784 (N_8784,N_7546,N_7727);
nand U8785 (N_8785,N_7211,N_7481);
nor U8786 (N_8786,N_7200,N_7205);
nand U8787 (N_8787,N_7279,N_7595);
or U8788 (N_8788,N_7847,N_7725);
nor U8789 (N_8789,N_7645,N_7818);
or U8790 (N_8790,N_7920,N_7528);
or U8791 (N_8791,N_7786,N_7911);
nand U8792 (N_8792,N_7837,N_7401);
nand U8793 (N_8793,N_7503,N_7256);
nor U8794 (N_8794,N_7522,N_7247);
nand U8795 (N_8795,N_7082,N_7289);
and U8796 (N_8796,N_7527,N_7406);
nand U8797 (N_8797,N_7163,N_7834);
and U8798 (N_8798,N_7695,N_7126);
nor U8799 (N_8799,N_7554,N_7792);
or U8800 (N_8800,N_7457,N_7334);
nand U8801 (N_8801,N_7782,N_7041);
nor U8802 (N_8802,N_7664,N_7264);
nand U8803 (N_8803,N_7477,N_7529);
nand U8804 (N_8804,N_7511,N_7279);
and U8805 (N_8805,N_7846,N_7364);
and U8806 (N_8806,N_7784,N_7086);
nand U8807 (N_8807,N_7876,N_7630);
nand U8808 (N_8808,N_7619,N_7886);
nor U8809 (N_8809,N_7237,N_7892);
nor U8810 (N_8810,N_7645,N_7314);
and U8811 (N_8811,N_7818,N_7063);
nor U8812 (N_8812,N_7505,N_7720);
or U8813 (N_8813,N_7585,N_7014);
nand U8814 (N_8814,N_7912,N_7024);
or U8815 (N_8815,N_7322,N_7951);
or U8816 (N_8816,N_7532,N_7149);
or U8817 (N_8817,N_7243,N_7104);
nand U8818 (N_8818,N_7771,N_7945);
or U8819 (N_8819,N_7747,N_7897);
or U8820 (N_8820,N_7643,N_7995);
nor U8821 (N_8821,N_7572,N_7268);
and U8822 (N_8822,N_7942,N_7190);
and U8823 (N_8823,N_7593,N_7603);
or U8824 (N_8824,N_7936,N_7518);
nand U8825 (N_8825,N_7187,N_7045);
nor U8826 (N_8826,N_7413,N_7476);
and U8827 (N_8827,N_7989,N_7854);
and U8828 (N_8828,N_7806,N_7519);
xnor U8829 (N_8829,N_7769,N_7475);
nand U8830 (N_8830,N_7982,N_7259);
nor U8831 (N_8831,N_7260,N_7819);
or U8832 (N_8832,N_7848,N_7814);
nor U8833 (N_8833,N_7498,N_7180);
nand U8834 (N_8834,N_7924,N_7848);
and U8835 (N_8835,N_7849,N_7673);
nor U8836 (N_8836,N_7811,N_7086);
nand U8837 (N_8837,N_7324,N_7027);
and U8838 (N_8838,N_7929,N_7718);
nor U8839 (N_8839,N_7596,N_7364);
and U8840 (N_8840,N_7244,N_7626);
or U8841 (N_8841,N_7805,N_7139);
nand U8842 (N_8842,N_7110,N_7109);
or U8843 (N_8843,N_7312,N_7194);
or U8844 (N_8844,N_7196,N_7663);
nand U8845 (N_8845,N_7815,N_7773);
or U8846 (N_8846,N_7074,N_7281);
and U8847 (N_8847,N_7413,N_7511);
nor U8848 (N_8848,N_7919,N_7468);
nand U8849 (N_8849,N_7115,N_7357);
nand U8850 (N_8850,N_7047,N_7504);
and U8851 (N_8851,N_7199,N_7577);
nand U8852 (N_8852,N_7156,N_7404);
and U8853 (N_8853,N_7285,N_7436);
nand U8854 (N_8854,N_7808,N_7901);
or U8855 (N_8855,N_7200,N_7195);
nand U8856 (N_8856,N_7014,N_7869);
nand U8857 (N_8857,N_7128,N_7123);
or U8858 (N_8858,N_7045,N_7152);
and U8859 (N_8859,N_7849,N_7943);
nand U8860 (N_8860,N_7974,N_7074);
or U8861 (N_8861,N_7438,N_7794);
nand U8862 (N_8862,N_7719,N_7937);
nor U8863 (N_8863,N_7256,N_7488);
or U8864 (N_8864,N_7344,N_7490);
or U8865 (N_8865,N_7528,N_7508);
nor U8866 (N_8866,N_7091,N_7174);
nand U8867 (N_8867,N_7669,N_7189);
or U8868 (N_8868,N_7376,N_7758);
nand U8869 (N_8869,N_7778,N_7549);
or U8870 (N_8870,N_7981,N_7823);
and U8871 (N_8871,N_7670,N_7739);
nand U8872 (N_8872,N_7752,N_7060);
or U8873 (N_8873,N_7874,N_7213);
and U8874 (N_8874,N_7128,N_7072);
xor U8875 (N_8875,N_7474,N_7814);
or U8876 (N_8876,N_7548,N_7098);
and U8877 (N_8877,N_7820,N_7049);
nand U8878 (N_8878,N_7094,N_7922);
and U8879 (N_8879,N_7927,N_7147);
nor U8880 (N_8880,N_7296,N_7732);
or U8881 (N_8881,N_7532,N_7840);
nor U8882 (N_8882,N_7763,N_7963);
nand U8883 (N_8883,N_7936,N_7197);
nand U8884 (N_8884,N_7986,N_7845);
nor U8885 (N_8885,N_7404,N_7989);
nand U8886 (N_8886,N_7771,N_7695);
nand U8887 (N_8887,N_7728,N_7966);
or U8888 (N_8888,N_7807,N_7044);
nor U8889 (N_8889,N_7607,N_7874);
or U8890 (N_8890,N_7226,N_7019);
nor U8891 (N_8891,N_7777,N_7891);
and U8892 (N_8892,N_7810,N_7673);
or U8893 (N_8893,N_7789,N_7982);
nor U8894 (N_8894,N_7685,N_7905);
and U8895 (N_8895,N_7224,N_7300);
nand U8896 (N_8896,N_7824,N_7711);
and U8897 (N_8897,N_7190,N_7968);
nor U8898 (N_8898,N_7652,N_7084);
nor U8899 (N_8899,N_7485,N_7528);
and U8900 (N_8900,N_7703,N_7932);
nor U8901 (N_8901,N_7868,N_7252);
nor U8902 (N_8902,N_7142,N_7982);
and U8903 (N_8903,N_7681,N_7010);
and U8904 (N_8904,N_7861,N_7061);
or U8905 (N_8905,N_7695,N_7324);
and U8906 (N_8906,N_7613,N_7254);
and U8907 (N_8907,N_7670,N_7883);
nor U8908 (N_8908,N_7813,N_7686);
and U8909 (N_8909,N_7866,N_7528);
or U8910 (N_8910,N_7552,N_7783);
or U8911 (N_8911,N_7286,N_7442);
and U8912 (N_8912,N_7930,N_7667);
and U8913 (N_8913,N_7836,N_7701);
nor U8914 (N_8914,N_7327,N_7836);
or U8915 (N_8915,N_7485,N_7239);
nand U8916 (N_8916,N_7578,N_7465);
or U8917 (N_8917,N_7515,N_7247);
nand U8918 (N_8918,N_7443,N_7230);
or U8919 (N_8919,N_7299,N_7684);
or U8920 (N_8920,N_7374,N_7629);
or U8921 (N_8921,N_7887,N_7582);
nor U8922 (N_8922,N_7513,N_7144);
nand U8923 (N_8923,N_7478,N_7078);
nor U8924 (N_8924,N_7672,N_7322);
nor U8925 (N_8925,N_7308,N_7946);
and U8926 (N_8926,N_7571,N_7569);
nor U8927 (N_8927,N_7487,N_7190);
or U8928 (N_8928,N_7504,N_7738);
nor U8929 (N_8929,N_7995,N_7452);
or U8930 (N_8930,N_7478,N_7538);
nand U8931 (N_8931,N_7331,N_7286);
or U8932 (N_8932,N_7041,N_7856);
and U8933 (N_8933,N_7389,N_7140);
nor U8934 (N_8934,N_7852,N_7243);
nor U8935 (N_8935,N_7071,N_7601);
nor U8936 (N_8936,N_7488,N_7865);
nand U8937 (N_8937,N_7778,N_7410);
or U8938 (N_8938,N_7312,N_7868);
or U8939 (N_8939,N_7930,N_7701);
nor U8940 (N_8940,N_7501,N_7176);
or U8941 (N_8941,N_7884,N_7225);
and U8942 (N_8942,N_7465,N_7199);
or U8943 (N_8943,N_7679,N_7012);
and U8944 (N_8944,N_7420,N_7964);
and U8945 (N_8945,N_7127,N_7248);
or U8946 (N_8946,N_7759,N_7298);
and U8947 (N_8947,N_7543,N_7996);
nor U8948 (N_8948,N_7105,N_7299);
nor U8949 (N_8949,N_7703,N_7819);
nand U8950 (N_8950,N_7209,N_7434);
nand U8951 (N_8951,N_7825,N_7758);
or U8952 (N_8952,N_7612,N_7597);
xnor U8953 (N_8953,N_7463,N_7792);
and U8954 (N_8954,N_7979,N_7145);
nand U8955 (N_8955,N_7507,N_7415);
nand U8956 (N_8956,N_7605,N_7268);
nor U8957 (N_8957,N_7956,N_7440);
nor U8958 (N_8958,N_7653,N_7583);
or U8959 (N_8959,N_7171,N_7170);
or U8960 (N_8960,N_7381,N_7978);
and U8961 (N_8961,N_7313,N_7212);
and U8962 (N_8962,N_7495,N_7605);
and U8963 (N_8963,N_7812,N_7312);
nand U8964 (N_8964,N_7013,N_7138);
nand U8965 (N_8965,N_7664,N_7938);
and U8966 (N_8966,N_7910,N_7306);
nand U8967 (N_8967,N_7653,N_7362);
nor U8968 (N_8968,N_7211,N_7868);
nor U8969 (N_8969,N_7011,N_7027);
nand U8970 (N_8970,N_7122,N_7079);
nor U8971 (N_8971,N_7540,N_7877);
nand U8972 (N_8972,N_7688,N_7698);
and U8973 (N_8973,N_7947,N_7476);
nand U8974 (N_8974,N_7994,N_7082);
nor U8975 (N_8975,N_7626,N_7394);
or U8976 (N_8976,N_7010,N_7128);
and U8977 (N_8977,N_7277,N_7326);
nor U8978 (N_8978,N_7211,N_7415);
nand U8979 (N_8979,N_7133,N_7938);
and U8980 (N_8980,N_7457,N_7163);
nand U8981 (N_8981,N_7227,N_7403);
nand U8982 (N_8982,N_7854,N_7679);
nand U8983 (N_8983,N_7202,N_7873);
or U8984 (N_8984,N_7104,N_7682);
nand U8985 (N_8985,N_7275,N_7107);
nor U8986 (N_8986,N_7713,N_7767);
and U8987 (N_8987,N_7481,N_7196);
nand U8988 (N_8988,N_7514,N_7995);
nor U8989 (N_8989,N_7167,N_7576);
or U8990 (N_8990,N_7517,N_7805);
nand U8991 (N_8991,N_7258,N_7774);
or U8992 (N_8992,N_7061,N_7338);
and U8993 (N_8993,N_7064,N_7172);
nor U8994 (N_8994,N_7057,N_7704);
nor U8995 (N_8995,N_7144,N_7196);
nand U8996 (N_8996,N_7654,N_7701);
or U8997 (N_8997,N_7933,N_7009);
or U8998 (N_8998,N_7038,N_7607);
nor U8999 (N_8999,N_7605,N_7895);
or U9000 (N_9000,N_8516,N_8017);
nand U9001 (N_9001,N_8337,N_8299);
and U9002 (N_9002,N_8548,N_8515);
and U9003 (N_9003,N_8882,N_8644);
nor U9004 (N_9004,N_8174,N_8962);
nand U9005 (N_9005,N_8471,N_8066);
or U9006 (N_9006,N_8592,N_8960);
or U9007 (N_9007,N_8406,N_8971);
and U9008 (N_9008,N_8306,N_8150);
nand U9009 (N_9009,N_8462,N_8772);
nand U9010 (N_9010,N_8566,N_8658);
or U9011 (N_9011,N_8062,N_8929);
nor U9012 (N_9012,N_8187,N_8199);
or U9013 (N_9013,N_8068,N_8395);
nand U9014 (N_9014,N_8727,N_8993);
nand U9015 (N_9015,N_8116,N_8864);
nand U9016 (N_9016,N_8156,N_8500);
nand U9017 (N_9017,N_8710,N_8538);
or U9018 (N_9018,N_8517,N_8753);
nor U9019 (N_9019,N_8442,N_8736);
or U9020 (N_9020,N_8280,N_8902);
and U9021 (N_9021,N_8126,N_8326);
and U9022 (N_9022,N_8135,N_8679);
nand U9023 (N_9023,N_8848,N_8943);
nor U9024 (N_9024,N_8480,N_8999);
nand U9025 (N_9025,N_8537,N_8610);
and U9026 (N_9026,N_8478,N_8869);
and U9027 (N_9027,N_8502,N_8122);
nand U9028 (N_9028,N_8323,N_8889);
nand U9029 (N_9029,N_8165,N_8413);
or U9030 (N_9030,N_8855,N_8910);
and U9031 (N_9031,N_8585,N_8856);
or U9032 (N_9032,N_8059,N_8191);
and U9033 (N_9033,N_8843,N_8955);
and U9034 (N_9034,N_8650,N_8005);
or U9035 (N_9035,N_8108,N_8268);
and U9036 (N_9036,N_8933,N_8540);
nor U9037 (N_9037,N_8805,N_8524);
nor U9038 (N_9038,N_8518,N_8798);
and U9039 (N_9039,N_8988,N_8481);
or U9040 (N_9040,N_8120,N_8714);
and U9041 (N_9041,N_8655,N_8691);
and U9042 (N_9042,N_8789,N_8594);
and U9043 (N_9043,N_8099,N_8737);
nor U9044 (N_9044,N_8035,N_8352);
and U9045 (N_9045,N_8436,N_8290);
nor U9046 (N_9046,N_8282,N_8899);
or U9047 (N_9047,N_8400,N_8200);
nand U9048 (N_9048,N_8508,N_8872);
nand U9049 (N_9049,N_8365,N_8275);
or U9050 (N_9050,N_8366,N_8942);
nand U9051 (N_9051,N_8241,N_8162);
nand U9052 (N_9052,N_8274,N_8204);
or U9053 (N_9053,N_8341,N_8130);
nand U9054 (N_9054,N_8056,N_8997);
nor U9055 (N_9055,N_8036,N_8243);
nand U9056 (N_9056,N_8473,N_8060);
nor U9057 (N_9057,N_8022,N_8852);
or U9058 (N_9058,N_8925,N_8778);
nand U9059 (N_9059,N_8101,N_8578);
or U9060 (N_9060,N_8901,N_8086);
nor U9061 (N_9061,N_8031,N_8945);
or U9062 (N_9062,N_8976,N_8892);
and U9063 (N_9063,N_8153,N_8475);
nor U9064 (N_9064,N_8819,N_8620);
nand U9065 (N_9065,N_8996,N_8820);
and U9066 (N_9066,N_8923,N_8982);
and U9067 (N_9067,N_8379,N_8277);
nand U9068 (N_9068,N_8513,N_8296);
or U9069 (N_9069,N_8761,N_8032);
nand U9070 (N_9070,N_8083,N_8407);
or U9071 (N_9071,N_8426,N_8968);
and U9072 (N_9072,N_8980,N_8535);
nand U9073 (N_9073,N_8951,N_8850);
nand U9074 (N_9074,N_8904,N_8432);
nand U9075 (N_9075,N_8707,N_8709);
nand U9076 (N_9076,N_8396,N_8956);
nand U9077 (N_9077,N_8703,N_8424);
nor U9078 (N_9078,N_8356,N_8970);
nor U9079 (N_9079,N_8453,N_8371);
nor U9080 (N_9080,N_8530,N_8809);
nor U9081 (N_9081,N_8950,N_8986);
or U9082 (N_9082,N_8417,N_8701);
nor U9083 (N_9083,N_8724,N_8105);
nand U9084 (N_9084,N_8281,N_8106);
or U9085 (N_9085,N_8653,N_8414);
or U9086 (N_9086,N_8219,N_8217);
nand U9087 (N_9087,N_8263,N_8713);
nand U9088 (N_9088,N_8776,N_8773);
nor U9089 (N_9089,N_8596,N_8561);
and U9090 (N_9090,N_8279,N_8912);
nand U9091 (N_9091,N_8770,N_8639);
or U9092 (N_9092,N_8472,N_8792);
or U9093 (N_9093,N_8553,N_8924);
or U9094 (N_9094,N_8868,N_8952);
nand U9095 (N_9095,N_8229,N_8160);
and U9096 (N_9096,N_8754,N_8532);
and U9097 (N_9097,N_8763,N_8900);
and U9098 (N_9098,N_8291,N_8208);
nor U9099 (N_9099,N_8370,N_8195);
and U9100 (N_9100,N_8214,N_8682);
nand U9101 (N_9101,N_8461,N_8368);
or U9102 (N_9102,N_8771,N_8452);
nand U9103 (N_9103,N_8427,N_8209);
and U9104 (N_9104,N_8460,N_8363);
or U9105 (N_9105,N_8410,N_8562);
nor U9106 (N_9106,N_8775,N_8690);
nor U9107 (N_9107,N_8227,N_8542);
nor U9108 (N_9108,N_8621,N_8939);
and U9109 (N_9109,N_8878,N_8359);
nor U9110 (N_9110,N_8874,N_8322);
and U9111 (N_9111,N_8249,N_8800);
nand U9112 (N_9112,N_8154,N_8786);
and U9113 (N_9113,N_8206,N_8894);
nor U9114 (N_9114,N_8766,N_8492);
or U9115 (N_9115,N_8293,N_8568);
and U9116 (N_9116,N_8705,N_8308);
or U9117 (N_9117,N_8725,N_8815);
and U9118 (N_9118,N_8300,N_8493);
and U9119 (N_9119,N_8087,N_8203);
nand U9120 (N_9120,N_8314,N_8015);
nand U9121 (N_9121,N_8842,N_8834);
nand U9122 (N_9122,N_8526,N_8425);
and U9123 (N_9123,N_8391,N_8448);
nor U9124 (N_9124,N_8270,N_8877);
nand U9125 (N_9125,N_8098,N_8258);
or U9126 (N_9126,N_8584,N_8088);
and U9127 (N_9127,N_8262,N_8930);
and U9128 (N_9128,N_8913,N_8218);
nand U9129 (N_9129,N_8334,N_8489);
or U9130 (N_9130,N_8089,N_8704);
nor U9131 (N_9131,N_8756,N_8392);
nand U9132 (N_9132,N_8601,N_8388);
nand U9133 (N_9133,N_8587,N_8459);
nor U9134 (N_9134,N_8885,N_8038);
nor U9135 (N_9135,N_8433,N_8260);
nor U9136 (N_9136,N_8879,N_8065);
and U9137 (N_9137,N_8267,N_8826);
and U9138 (N_9138,N_8495,N_8304);
and U9139 (N_9139,N_8543,N_8745);
and U9140 (N_9140,N_8932,N_8409);
or U9141 (N_9141,N_8579,N_8908);
and U9142 (N_9142,N_8733,N_8807);
nor U9143 (N_9143,N_8198,N_8115);
nor U9144 (N_9144,N_8905,N_8397);
or U9145 (N_9145,N_8257,N_8250);
nand U9146 (N_9146,N_8335,N_8081);
or U9147 (N_9147,N_8180,N_8687);
nor U9148 (N_9148,N_8172,N_8230);
or U9149 (N_9149,N_8264,N_8070);
and U9150 (N_9150,N_8317,N_8283);
and U9151 (N_9151,N_8236,N_8234);
or U9152 (N_9152,N_8688,N_8074);
nor U9153 (N_9153,N_8445,N_8696);
or U9154 (N_9154,N_8085,N_8567);
xnor U9155 (N_9155,N_8494,N_8097);
nor U9156 (N_9156,N_8129,N_8350);
or U9157 (N_9157,N_8643,N_8179);
nand U9158 (N_9158,N_8926,N_8576);
nor U9159 (N_9159,N_8469,N_8064);
and U9160 (N_9160,N_8928,N_8813);
nor U9161 (N_9161,N_8496,N_8573);
and U9162 (N_9162,N_8802,N_8019);
or U9163 (N_9163,N_8529,N_8752);
nand U9164 (N_9164,N_8716,N_8636);
and U9165 (N_9165,N_8810,N_8569);
nand U9166 (N_9166,N_8147,N_8865);
and U9167 (N_9167,N_8833,N_8630);
nand U9168 (N_9168,N_8666,N_8523);
and U9169 (N_9169,N_8975,N_8367);
or U9170 (N_9170,N_8665,N_8223);
and U9171 (N_9171,N_8828,N_8963);
or U9172 (N_9172,N_8791,N_8044);
nand U9173 (N_9173,N_8069,N_8830);
nor U9174 (N_9174,N_8215,N_8803);
nor U9175 (N_9175,N_8292,N_8261);
or U9176 (N_9176,N_8556,N_8186);
and U9177 (N_9177,N_8514,N_8284);
nand U9178 (N_9178,N_8190,N_8987);
or U9179 (N_9179,N_8605,N_8862);
nor U9180 (N_9180,N_8273,N_8033);
or U9181 (N_9181,N_8210,N_8266);
and U9182 (N_9182,N_8151,N_8028);
and U9183 (N_9183,N_8891,N_8607);
nor U9184 (N_9184,N_8053,N_8510);
nand U9185 (N_9185,N_8037,N_8712);
and U9186 (N_9186,N_8765,N_8245);
nor U9187 (N_9187,N_8112,N_8534);
nor U9188 (N_9188,N_8182,N_8618);
nand U9189 (N_9189,N_8123,N_8822);
nor U9190 (N_9190,N_8477,N_8663);
nand U9191 (N_9191,N_8132,N_8845);
nand U9192 (N_9192,N_8743,N_8564);
or U9193 (N_9193,N_8221,N_8231);
nor U9194 (N_9194,N_8507,N_8604);
nand U9195 (N_9195,N_8404,N_8042);
and U9196 (N_9196,N_8898,N_8434);
and U9197 (N_9197,N_8646,N_8829);
nor U9198 (N_9198,N_8411,N_8590);
and U9199 (N_9199,N_8840,N_8046);
nand U9200 (N_9200,N_8063,N_8779);
and U9201 (N_9201,N_8652,N_8398);
nor U9202 (N_9202,N_8144,N_8094);
or U9203 (N_9203,N_8415,N_8512);
nor U9204 (N_9204,N_8797,N_8353);
or U9205 (N_9205,N_8732,N_8806);
or U9206 (N_9206,N_8661,N_8740);
and U9207 (N_9207,N_8609,N_8985);
nand U9208 (N_9208,N_8207,N_8808);
and U9209 (N_9209,N_8787,N_8429);
nand U9210 (N_9210,N_8374,N_8004);
nand U9211 (N_9211,N_8138,N_8318);
and U9212 (N_9212,N_8811,N_8043);
and U9213 (N_9213,N_8121,N_8201);
nand U9214 (N_9214,N_8312,N_8909);
or U9215 (N_9215,N_8938,N_8100);
and U9216 (N_9216,N_8054,N_8265);
or U9217 (N_9217,N_8315,N_8936);
and U9218 (N_9218,N_8835,N_8795);
or U9219 (N_9219,N_8801,N_8384);
nand U9220 (N_9220,N_8405,N_8825);
or U9221 (N_9221,N_8305,N_8149);
nor U9222 (N_9222,N_8155,N_8672);
nand U9223 (N_9223,N_8657,N_8216);
nor U9224 (N_9224,N_8599,N_8248);
or U9225 (N_9225,N_8664,N_8464);
and U9226 (N_9226,N_8345,N_8611);
nand U9227 (N_9227,N_8757,N_8456);
and U9228 (N_9228,N_8339,N_8422);
and U9229 (N_9229,N_8947,N_8883);
or U9230 (N_9230,N_8915,N_8613);
and U9231 (N_9231,N_8272,N_8593);
nand U9232 (N_9232,N_8301,N_8252);
nand U9233 (N_9233,N_8159,N_8364);
and U9234 (N_9234,N_8637,N_8571);
nand U9235 (N_9235,N_8141,N_8550);
nand U9236 (N_9236,N_8555,N_8055);
nor U9237 (N_9237,N_8747,N_8259);
nor U9238 (N_9238,N_8602,N_8615);
and U9239 (N_9239,N_8648,N_8606);
and U9240 (N_9240,N_8981,N_8814);
and U9241 (N_9241,N_8220,N_8226);
or U9242 (N_9242,N_8953,N_8916);
and U9243 (N_9243,N_8598,N_8817);
nor U9244 (N_9244,N_8447,N_8642);
or U9245 (N_9245,N_8622,N_8333);
nor U9246 (N_9246,N_8104,N_8839);
xor U9247 (N_9247,N_8177,N_8362);
or U9248 (N_9248,N_8948,N_8027);
nor U9249 (N_9249,N_8026,N_8823);
nand U9250 (N_9250,N_8145,N_8175);
and U9251 (N_9251,N_8946,N_8832);
nor U9252 (N_9252,N_8237,N_8884);
and U9253 (N_9253,N_8706,N_8197);
nand U9254 (N_9254,N_8780,N_8441);
nand U9255 (N_9255,N_8790,N_8423);
xor U9256 (N_9256,N_8612,N_8390);
nand U9257 (N_9257,N_8498,N_8316);
or U9258 (N_9258,N_8194,N_8189);
nor U9259 (N_9259,N_8457,N_8491);
nand U9260 (N_9260,N_8146,N_8185);
and U9261 (N_9261,N_8233,N_8858);
nor U9262 (N_9262,N_8444,N_8139);
nand U9263 (N_9263,N_8533,N_8431);
nand U9264 (N_9264,N_8418,N_8010);
nor U9265 (N_9265,N_8559,N_8631);
and U9266 (N_9266,N_8821,N_8992);
or U9267 (N_9267,N_8769,N_8973);
nor U9268 (N_9268,N_8857,N_8096);
nor U9269 (N_9269,N_8040,N_8640);
nor U9270 (N_9270,N_8678,N_8689);
nand U9271 (N_9271,N_8846,N_8307);
or U9272 (N_9272,N_8718,N_8127);
and U9273 (N_9273,N_8369,N_8479);
nand U9274 (N_9274,N_8178,N_8880);
nor U9275 (N_9275,N_8624,N_8354);
or U9276 (N_9276,N_8079,N_8940);
and U9277 (N_9277,N_8298,N_8488);
nand U9278 (N_9278,N_8838,N_8034);
and U9279 (N_9279,N_8890,N_8991);
nand U9280 (N_9280,N_8294,N_8255);
and U9281 (N_9281,N_8668,N_8050);
nor U9282 (N_9282,N_8133,N_8377);
and U9283 (N_9283,N_8777,N_8399);
nand U9284 (N_9284,N_8171,N_8114);
or U9285 (N_9285,N_8860,N_8870);
or U9286 (N_9286,N_8157,N_8551);
nor U9287 (N_9287,N_8785,N_8443);
and U9288 (N_9288,N_8583,N_8387);
nand U9289 (N_9289,N_8673,N_8324);
nor U9290 (N_9290,N_8061,N_8376);
and U9291 (N_9291,N_8468,N_8343);
and U9292 (N_9292,N_8505,N_8107);
nor U9293 (N_9293,N_8325,N_8454);
and U9294 (N_9294,N_8007,N_8205);
and U9295 (N_9295,N_8254,N_8628);
and U9296 (N_9296,N_8289,N_8244);
and U9297 (N_9297,N_8438,N_8213);
and U9298 (N_9298,N_8692,N_8656);
or U9299 (N_9299,N_8541,N_8224);
nand U9300 (N_9300,N_8309,N_8449);
nor U9301 (N_9301,N_8483,N_8455);
nor U9302 (N_9302,N_8076,N_8119);
or U9303 (N_9303,N_8954,N_8173);
or U9304 (N_9304,N_8021,N_8558);
xnor U9305 (N_9305,N_8764,N_8378);
nor U9306 (N_9306,N_8949,N_8887);
or U9307 (N_9307,N_8546,N_8225);
or U9308 (N_9308,N_8020,N_8168);
nand U9309 (N_9309,N_8685,N_8793);
xor U9310 (N_9310,N_8781,N_8381);
nand U9311 (N_9311,N_8458,N_8684);
nand U9312 (N_9312,N_8974,N_8011);
or U9313 (N_9313,N_8729,N_8708);
and U9314 (N_9314,N_8519,N_8351);
and U9315 (N_9315,N_8577,N_8118);
nand U9316 (N_9316,N_8762,N_8389);
nand U9317 (N_9317,N_8202,N_8634);
nor U9318 (N_9318,N_8586,N_8827);
or U9319 (N_9319,N_8340,N_8499);
or U9320 (N_9320,N_8768,N_8163);
nand U9321 (N_9321,N_8674,N_8446);
nand U9322 (N_9322,N_8675,N_8049);
or U9323 (N_9323,N_8723,N_8193);
nand U9324 (N_9324,N_8600,N_8623);
or U9325 (N_9325,N_8329,N_8057);
xnor U9326 (N_9326,N_8931,N_8285);
nor U9327 (N_9327,N_8698,N_8419);
nor U9328 (N_9328,N_8385,N_8288);
nand U9329 (N_9329,N_8751,N_8730);
nand U9330 (N_9330,N_8603,N_8346);
and U9331 (N_9331,N_8873,N_8818);
nor U9332 (N_9332,N_8719,N_8092);
nor U9333 (N_9333,N_8563,N_8967);
nand U9334 (N_9334,N_8025,N_8886);
or U9335 (N_9335,N_8702,N_8450);
nand U9336 (N_9336,N_8103,N_8859);
or U9337 (N_9337,N_8965,N_8744);
nand U9338 (N_9338,N_8321,N_8750);
nor U9339 (N_9339,N_8009,N_8140);
or U9340 (N_9340,N_8520,N_8073);
nor U9341 (N_9341,N_8597,N_8242);
nor U9342 (N_9342,N_8582,N_8547);
and U9343 (N_9343,N_8632,N_8972);
and U9344 (N_9344,N_8522,N_8310);
nor U9345 (N_9345,N_8565,N_8161);
nor U9346 (N_9346,N_8721,N_8699);
nand U9347 (N_9347,N_8794,N_8503);
xnor U9348 (N_9348,N_8196,N_8013);
nand U9349 (N_9349,N_8918,N_8029);
or U9350 (N_9350,N_8188,N_8402);
or U9351 (N_9351,N_8041,N_8758);
nor U9352 (N_9352,N_8686,N_8357);
and U9353 (N_9353,N_8783,N_8654);
nor U9354 (N_9354,N_8552,N_8228);
nor U9355 (N_9355,N_8012,N_8907);
or U9356 (N_9356,N_8633,N_8428);
or U9357 (N_9357,N_8430,N_8176);
nor U9358 (N_9358,N_8774,N_8001);
and U9359 (N_9359,N_8003,N_8077);
or U9360 (N_9360,N_8626,N_8235);
or U9361 (N_9361,N_8647,N_8671);
nand U9362 (N_9362,N_8681,N_8591);
nand U9363 (N_9363,N_8403,N_8080);
or U9364 (N_9364,N_8896,N_8311);
or U9365 (N_9365,N_8170,N_8212);
or U9366 (N_9366,N_8536,N_8888);
or U9367 (N_9367,N_8058,N_8184);
nand U9368 (N_9368,N_8297,N_8934);
or U9369 (N_9369,N_8738,N_8903);
or U9370 (N_9370,N_8977,N_8328);
and U9371 (N_9371,N_8361,N_8358);
nor U9372 (N_9372,N_8372,N_8093);
nand U9373 (N_9373,N_8439,N_8589);
nand U9374 (N_9374,N_8386,N_8539);
and U9375 (N_9375,N_8711,N_8693);
and U9376 (N_9376,N_8421,N_8222);
nand U9377 (N_9377,N_8435,N_8670);
or U9378 (N_9378,N_8841,N_8669);
or U9379 (N_9379,N_8497,N_8167);
or U9380 (N_9380,N_8239,N_8651);
nor U9381 (N_9381,N_8731,N_8580);
and U9382 (N_9382,N_8662,N_8978);
and U9383 (N_9383,N_8572,N_8095);
nand U9384 (N_9384,N_8588,N_8240);
and U9385 (N_9385,N_8124,N_8554);
and U9386 (N_9386,N_8148,N_8330);
and U9387 (N_9387,N_8635,N_8990);
nand U9388 (N_9388,N_8128,N_8749);
and U9389 (N_9389,N_8917,N_8067);
nand U9390 (N_9390,N_8627,N_8232);
nand U9391 (N_9391,N_8320,N_8169);
and U9392 (N_9392,N_8109,N_8837);
or U9393 (N_9393,N_8608,N_8911);
nor U9394 (N_9394,N_8451,N_8741);
nand U9395 (N_9395,N_8984,N_8137);
and U9396 (N_9396,N_8720,N_8521);
or U9397 (N_9397,N_8166,N_8474);
or U9398 (N_9398,N_8158,N_8549);
nor U9399 (N_9399,N_8509,N_8957);
or U9400 (N_9400,N_8742,N_8935);
nor U9401 (N_9401,N_8286,N_8560);
and U9402 (N_9402,N_8111,N_8287);
nor U9403 (N_9403,N_8336,N_8920);
and U9404 (N_9404,N_8412,N_8238);
and U9405 (N_9405,N_8000,N_8966);
nor U9406 (N_9406,N_8861,N_8360);
nor U9407 (N_9407,N_8748,N_8348);
nor U9408 (N_9408,N_8824,N_8575);
nand U9409 (N_9409,N_8338,N_8767);
nand U9410 (N_9410,N_8875,N_8465);
or U9411 (N_9411,N_8484,N_8799);
or U9412 (N_9412,N_8511,N_8332);
nand U9413 (N_9413,N_8871,N_8504);
nor U9414 (N_9414,N_8486,N_8804);
or U9415 (N_9415,N_8849,N_8253);
nor U9416 (N_9416,N_8937,N_8969);
nor U9417 (N_9417,N_8619,N_8641);
or U9418 (N_9418,N_8866,N_8722);
nand U9419 (N_9419,N_8192,N_8078);
or U9420 (N_9420,N_8683,N_8760);
nor U9421 (N_9421,N_8476,N_8501);
nor U9422 (N_9422,N_8735,N_8844);
nand U9423 (N_9423,N_8256,N_8276);
and U9424 (N_9424,N_8964,N_8271);
nor U9425 (N_9425,N_8183,N_8544);
and U9426 (N_9426,N_8327,N_8893);
and U9427 (N_9427,N_8881,N_8788);
nand U9428 (N_9428,N_8347,N_8625);
nand U9429 (N_9429,N_8181,N_8303);
nor U9430 (N_9430,N_8581,N_8595);
or U9431 (N_9431,N_8863,N_8796);
nor U9432 (N_9432,N_8466,N_8921);
nor U9433 (N_9433,N_8437,N_8659);
nand U9434 (N_9434,N_8979,N_8812);
nor U9435 (N_9435,N_8616,N_8383);
nand U9436 (N_9436,N_8313,N_8629);
nor U9437 (N_9437,N_8463,N_8531);
nand U9438 (N_9438,N_8344,N_8676);
nand U9439 (N_9439,N_8331,N_8545);
nand U9440 (N_9440,N_8734,N_8998);
or U9441 (N_9441,N_8649,N_8867);
xnor U9442 (N_9442,N_8002,N_8487);
nand U9443 (N_9443,N_8071,N_8482);
nand U9444 (N_9444,N_8914,N_8574);
and U9445 (N_9445,N_8090,N_8251);
and U9446 (N_9446,N_8006,N_8164);
nor U9447 (N_9447,N_8091,N_8847);
nand U9448 (N_9448,N_8008,N_8051);
and U9449 (N_9449,N_8739,N_8667);
and U9450 (N_9450,N_8961,N_8490);
nand U9451 (N_9451,N_8102,N_8246);
nand U9452 (N_9452,N_8143,N_8697);
and U9453 (N_9453,N_8470,N_8876);
nand U9454 (N_9454,N_8728,N_8854);
nor U9455 (N_9455,N_8525,N_8994);
nor U9456 (N_9456,N_8922,N_8782);
and U9457 (N_9457,N_8125,N_8897);
or U9458 (N_9458,N_8831,N_8030);
or U9459 (N_9459,N_8117,N_8527);
or U9460 (N_9460,N_8680,N_8278);
nand U9461 (N_9461,N_8024,N_8506);
nand U9462 (N_9462,N_8382,N_8989);
nand U9463 (N_9463,N_8014,N_8113);
nor U9464 (N_9464,N_8557,N_8958);
nand U9465 (N_9465,N_8851,N_8072);
or U9466 (N_9466,N_8440,N_8420);
and U9467 (N_9467,N_8373,N_8467);
and U9468 (N_9468,N_8355,N_8836);
nand U9469 (N_9469,N_8131,N_8944);
nor U9470 (N_9470,N_8295,N_8759);
or U9471 (N_9471,N_8895,N_8142);
nor U9472 (N_9472,N_8152,N_8349);
nor U9473 (N_9473,N_8016,N_8408);
or U9474 (N_9474,N_8375,N_8717);
xor U9475 (N_9475,N_8906,N_8959);
nor U9476 (N_9476,N_8784,N_8302);
nand U9477 (N_9477,N_8816,N_8927);
nor U9478 (N_9478,N_8677,N_8048);
and U9479 (N_9479,N_8645,N_8394);
or U9480 (N_9480,N_8047,N_8995);
and U9481 (N_9481,N_8941,N_8018);
and U9482 (N_9482,N_8380,N_8638);
nor U9483 (N_9483,N_8023,N_8075);
and U9484 (N_9484,N_8660,N_8617);
nor U9485 (N_9485,N_8134,N_8700);
or U9486 (N_9486,N_8614,N_8211);
nor U9487 (N_9487,N_8528,N_8485);
and U9488 (N_9488,N_8052,N_8039);
nand U9489 (N_9489,N_8695,N_8269);
or U9490 (N_9490,N_8247,N_8726);
or U9491 (N_9491,N_8755,N_8694);
or U9492 (N_9492,N_8401,N_8082);
nor U9493 (N_9493,N_8715,N_8084);
or U9494 (N_9494,N_8319,N_8110);
and U9495 (N_9495,N_8416,N_8393);
nand U9496 (N_9496,N_8342,N_8919);
nand U9497 (N_9497,N_8853,N_8983);
nor U9498 (N_9498,N_8045,N_8136);
xor U9499 (N_9499,N_8570,N_8746);
or U9500 (N_9500,N_8090,N_8082);
and U9501 (N_9501,N_8414,N_8039);
or U9502 (N_9502,N_8397,N_8564);
nand U9503 (N_9503,N_8179,N_8621);
nor U9504 (N_9504,N_8673,N_8721);
and U9505 (N_9505,N_8646,N_8209);
or U9506 (N_9506,N_8290,N_8888);
and U9507 (N_9507,N_8444,N_8455);
or U9508 (N_9508,N_8449,N_8781);
and U9509 (N_9509,N_8453,N_8162);
nor U9510 (N_9510,N_8949,N_8537);
nand U9511 (N_9511,N_8377,N_8764);
and U9512 (N_9512,N_8792,N_8222);
or U9513 (N_9513,N_8291,N_8791);
or U9514 (N_9514,N_8976,N_8643);
and U9515 (N_9515,N_8388,N_8959);
or U9516 (N_9516,N_8114,N_8165);
nor U9517 (N_9517,N_8796,N_8103);
nand U9518 (N_9518,N_8658,N_8857);
or U9519 (N_9519,N_8872,N_8772);
nand U9520 (N_9520,N_8674,N_8076);
nor U9521 (N_9521,N_8393,N_8935);
and U9522 (N_9522,N_8618,N_8195);
or U9523 (N_9523,N_8650,N_8467);
nor U9524 (N_9524,N_8766,N_8158);
nor U9525 (N_9525,N_8454,N_8965);
or U9526 (N_9526,N_8360,N_8240);
or U9527 (N_9527,N_8210,N_8838);
or U9528 (N_9528,N_8343,N_8835);
nor U9529 (N_9529,N_8559,N_8317);
or U9530 (N_9530,N_8532,N_8962);
and U9531 (N_9531,N_8848,N_8011);
nor U9532 (N_9532,N_8812,N_8442);
nor U9533 (N_9533,N_8101,N_8209);
nor U9534 (N_9534,N_8031,N_8814);
nor U9535 (N_9535,N_8924,N_8219);
xnor U9536 (N_9536,N_8601,N_8158);
or U9537 (N_9537,N_8458,N_8158);
nand U9538 (N_9538,N_8417,N_8069);
or U9539 (N_9539,N_8633,N_8376);
and U9540 (N_9540,N_8976,N_8831);
nand U9541 (N_9541,N_8764,N_8191);
nor U9542 (N_9542,N_8646,N_8407);
and U9543 (N_9543,N_8048,N_8673);
or U9544 (N_9544,N_8020,N_8046);
nor U9545 (N_9545,N_8161,N_8685);
or U9546 (N_9546,N_8110,N_8495);
nand U9547 (N_9547,N_8477,N_8193);
nor U9548 (N_9548,N_8527,N_8001);
nor U9549 (N_9549,N_8508,N_8770);
and U9550 (N_9550,N_8827,N_8086);
nor U9551 (N_9551,N_8187,N_8649);
and U9552 (N_9552,N_8542,N_8854);
or U9553 (N_9553,N_8255,N_8480);
or U9554 (N_9554,N_8840,N_8811);
xor U9555 (N_9555,N_8029,N_8866);
nand U9556 (N_9556,N_8802,N_8806);
or U9557 (N_9557,N_8144,N_8100);
nor U9558 (N_9558,N_8683,N_8800);
or U9559 (N_9559,N_8482,N_8949);
nor U9560 (N_9560,N_8323,N_8667);
or U9561 (N_9561,N_8714,N_8648);
and U9562 (N_9562,N_8816,N_8711);
nand U9563 (N_9563,N_8215,N_8560);
nand U9564 (N_9564,N_8196,N_8176);
or U9565 (N_9565,N_8326,N_8190);
nor U9566 (N_9566,N_8998,N_8421);
nand U9567 (N_9567,N_8553,N_8857);
and U9568 (N_9568,N_8425,N_8727);
or U9569 (N_9569,N_8338,N_8412);
nor U9570 (N_9570,N_8369,N_8620);
nor U9571 (N_9571,N_8232,N_8136);
or U9572 (N_9572,N_8866,N_8445);
or U9573 (N_9573,N_8373,N_8110);
and U9574 (N_9574,N_8725,N_8603);
nor U9575 (N_9575,N_8044,N_8891);
and U9576 (N_9576,N_8233,N_8332);
and U9577 (N_9577,N_8666,N_8270);
nor U9578 (N_9578,N_8895,N_8180);
nand U9579 (N_9579,N_8881,N_8699);
nand U9580 (N_9580,N_8646,N_8427);
nand U9581 (N_9581,N_8593,N_8497);
nor U9582 (N_9582,N_8165,N_8007);
or U9583 (N_9583,N_8779,N_8712);
and U9584 (N_9584,N_8996,N_8519);
and U9585 (N_9585,N_8125,N_8903);
or U9586 (N_9586,N_8680,N_8852);
and U9587 (N_9587,N_8715,N_8586);
nor U9588 (N_9588,N_8683,N_8023);
and U9589 (N_9589,N_8945,N_8703);
nand U9590 (N_9590,N_8522,N_8295);
and U9591 (N_9591,N_8477,N_8504);
nand U9592 (N_9592,N_8460,N_8681);
nor U9593 (N_9593,N_8934,N_8457);
and U9594 (N_9594,N_8044,N_8246);
nor U9595 (N_9595,N_8388,N_8138);
and U9596 (N_9596,N_8657,N_8710);
or U9597 (N_9597,N_8241,N_8381);
and U9598 (N_9598,N_8051,N_8183);
and U9599 (N_9599,N_8490,N_8693);
and U9600 (N_9600,N_8895,N_8636);
nand U9601 (N_9601,N_8970,N_8558);
and U9602 (N_9602,N_8298,N_8650);
nand U9603 (N_9603,N_8801,N_8362);
and U9604 (N_9604,N_8320,N_8956);
nand U9605 (N_9605,N_8273,N_8472);
and U9606 (N_9606,N_8660,N_8843);
and U9607 (N_9607,N_8449,N_8896);
and U9608 (N_9608,N_8749,N_8517);
xnor U9609 (N_9609,N_8835,N_8022);
nor U9610 (N_9610,N_8522,N_8938);
and U9611 (N_9611,N_8777,N_8791);
nor U9612 (N_9612,N_8984,N_8696);
or U9613 (N_9613,N_8323,N_8805);
and U9614 (N_9614,N_8162,N_8600);
nor U9615 (N_9615,N_8224,N_8672);
nor U9616 (N_9616,N_8688,N_8026);
nor U9617 (N_9617,N_8484,N_8425);
or U9618 (N_9618,N_8952,N_8437);
nor U9619 (N_9619,N_8515,N_8773);
nor U9620 (N_9620,N_8963,N_8220);
and U9621 (N_9621,N_8287,N_8104);
and U9622 (N_9622,N_8201,N_8829);
or U9623 (N_9623,N_8323,N_8205);
nand U9624 (N_9624,N_8296,N_8570);
or U9625 (N_9625,N_8183,N_8590);
nand U9626 (N_9626,N_8234,N_8296);
or U9627 (N_9627,N_8588,N_8578);
nor U9628 (N_9628,N_8093,N_8706);
nor U9629 (N_9629,N_8668,N_8906);
and U9630 (N_9630,N_8429,N_8869);
or U9631 (N_9631,N_8825,N_8140);
nor U9632 (N_9632,N_8924,N_8666);
or U9633 (N_9633,N_8252,N_8782);
or U9634 (N_9634,N_8847,N_8815);
and U9635 (N_9635,N_8345,N_8213);
nor U9636 (N_9636,N_8528,N_8107);
nor U9637 (N_9637,N_8043,N_8736);
or U9638 (N_9638,N_8020,N_8605);
and U9639 (N_9639,N_8043,N_8363);
nor U9640 (N_9640,N_8492,N_8252);
or U9641 (N_9641,N_8005,N_8263);
and U9642 (N_9642,N_8681,N_8197);
and U9643 (N_9643,N_8037,N_8528);
nand U9644 (N_9644,N_8280,N_8231);
nor U9645 (N_9645,N_8930,N_8902);
nor U9646 (N_9646,N_8637,N_8527);
or U9647 (N_9647,N_8572,N_8416);
nor U9648 (N_9648,N_8532,N_8103);
nand U9649 (N_9649,N_8401,N_8597);
nor U9650 (N_9650,N_8022,N_8952);
nand U9651 (N_9651,N_8835,N_8294);
nor U9652 (N_9652,N_8749,N_8596);
or U9653 (N_9653,N_8748,N_8936);
nand U9654 (N_9654,N_8466,N_8830);
or U9655 (N_9655,N_8983,N_8397);
nand U9656 (N_9656,N_8281,N_8730);
nor U9657 (N_9657,N_8907,N_8269);
nand U9658 (N_9658,N_8393,N_8075);
and U9659 (N_9659,N_8583,N_8885);
nor U9660 (N_9660,N_8976,N_8886);
nor U9661 (N_9661,N_8193,N_8865);
and U9662 (N_9662,N_8112,N_8337);
or U9663 (N_9663,N_8265,N_8440);
and U9664 (N_9664,N_8238,N_8839);
nor U9665 (N_9665,N_8154,N_8248);
nor U9666 (N_9666,N_8466,N_8562);
xnor U9667 (N_9667,N_8102,N_8513);
or U9668 (N_9668,N_8582,N_8289);
and U9669 (N_9669,N_8510,N_8863);
or U9670 (N_9670,N_8085,N_8448);
nor U9671 (N_9671,N_8963,N_8274);
nor U9672 (N_9672,N_8016,N_8745);
nand U9673 (N_9673,N_8074,N_8734);
nor U9674 (N_9674,N_8862,N_8201);
or U9675 (N_9675,N_8296,N_8065);
nand U9676 (N_9676,N_8659,N_8274);
nor U9677 (N_9677,N_8805,N_8909);
nor U9678 (N_9678,N_8981,N_8546);
or U9679 (N_9679,N_8513,N_8526);
or U9680 (N_9680,N_8339,N_8486);
or U9681 (N_9681,N_8594,N_8916);
and U9682 (N_9682,N_8586,N_8662);
or U9683 (N_9683,N_8730,N_8859);
or U9684 (N_9684,N_8458,N_8234);
nor U9685 (N_9685,N_8278,N_8178);
nand U9686 (N_9686,N_8117,N_8354);
nor U9687 (N_9687,N_8356,N_8230);
nand U9688 (N_9688,N_8722,N_8404);
or U9689 (N_9689,N_8811,N_8897);
and U9690 (N_9690,N_8877,N_8429);
nor U9691 (N_9691,N_8870,N_8618);
or U9692 (N_9692,N_8396,N_8949);
nor U9693 (N_9693,N_8843,N_8978);
nand U9694 (N_9694,N_8886,N_8997);
and U9695 (N_9695,N_8150,N_8262);
and U9696 (N_9696,N_8996,N_8971);
or U9697 (N_9697,N_8729,N_8849);
or U9698 (N_9698,N_8282,N_8299);
nand U9699 (N_9699,N_8707,N_8764);
nand U9700 (N_9700,N_8159,N_8052);
nand U9701 (N_9701,N_8913,N_8489);
and U9702 (N_9702,N_8678,N_8699);
or U9703 (N_9703,N_8938,N_8452);
and U9704 (N_9704,N_8788,N_8457);
nor U9705 (N_9705,N_8126,N_8034);
and U9706 (N_9706,N_8209,N_8964);
and U9707 (N_9707,N_8840,N_8213);
and U9708 (N_9708,N_8330,N_8321);
and U9709 (N_9709,N_8420,N_8142);
nand U9710 (N_9710,N_8925,N_8879);
nor U9711 (N_9711,N_8261,N_8549);
and U9712 (N_9712,N_8731,N_8774);
or U9713 (N_9713,N_8990,N_8934);
and U9714 (N_9714,N_8291,N_8082);
nor U9715 (N_9715,N_8916,N_8249);
or U9716 (N_9716,N_8295,N_8094);
and U9717 (N_9717,N_8061,N_8522);
nor U9718 (N_9718,N_8663,N_8950);
and U9719 (N_9719,N_8285,N_8945);
xor U9720 (N_9720,N_8652,N_8123);
nor U9721 (N_9721,N_8014,N_8223);
and U9722 (N_9722,N_8156,N_8371);
or U9723 (N_9723,N_8707,N_8318);
or U9724 (N_9724,N_8582,N_8416);
nand U9725 (N_9725,N_8479,N_8569);
nor U9726 (N_9726,N_8868,N_8346);
nand U9727 (N_9727,N_8426,N_8232);
nor U9728 (N_9728,N_8786,N_8435);
or U9729 (N_9729,N_8328,N_8967);
nand U9730 (N_9730,N_8693,N_8632);
nor U9731 (N_9731,N_8573,N_8224);
or U9732 (N_9732,N_8616,N_8470);
and U9733 (N_9733,N_8858,N_8458);
nand U9734 (N_9734,N_8799,N_8606);
and U9735 (N_9735,N_8729,N_8140);
nor U9736 (N_9736,N_8441,N_8179);
or U9737 (N_9737,N_8438,N_8768);
and U9738 (N_9738,N_8449,N_8290);
and U9739 (N_9739,N_8376,N_8030);
and U9740 (N_9740,N_8244,N_8066);
or U9741 (N_9741,N_8406,N_8860);
or U9742 (N_9742,N_8821,N_8467);
xnor U9743 (N_9743,N_8801,N_8394);
and U9744 (N_9744,N_8833,N_8511);
nand U9745 (N_9745,N_8049,N_8683);
nand U9746 (N_9746,N_8344,N_8682);
nor U9747 (N_9747,N_8953,N_8566);
nand U9748 (N_9748,N_8608,N_8733);
nand U9749 (N_9749,N_8724,N_8645);
nor U9750 (N_9750,N_8142,N_8825);
nand U9751 (N_9751,N_8455,N_8203);
or U9752 (N_9752,N_8830,N_8789);
nor U9753 (N_9753,N_8047,N_8829);
nand U9754 (N_9754,N_8998,N_8513);
nand U9755 (N_9755,N_8433,N_8335);
and U9756 (N_9756,N_8885,N_8773);
nand U9757 (N_9757,N_8174,N_8511);
and U9758 (N_9758,N_8021,N_8398);
nand U9759 (N_9759,N_8067,N_8198);
nand U9760 (N_9760,N_8076,N_8582);
nand U9761 (N_9761,N_8393,N_8364);
and U9762 (N_9762,N_8248,N_8416);
nor U9763 (N_9763,N_8098,N_8815);
nor U9764 (N_9764,N_8484,N_8389);
nand U9765 (N_9765,N_8681,N_8250);
or U9766 (N_9766,N_8184,N_8703);
nand U9767 (N_9767,N_8571,N_8704);
or U9768 (N_9768,N_8688,N_8908);
or U9769 (N_9769,N_8562,N_8563);
nand U9770 (N_9770,N_8244,N_8331);
or U9771 (N_9771,N_8849,N_8956);
and U9772 (N_9772,N_8921,N_8834);
nor U9773 (N_9773,N_8136,N_8558);
and U9774 (N_9774,N_8573,N_8018);
nor U9775 (N_9775,N_8958,N_8887);
and U9776 (N_9776,N_8185,N_8559);
nand U9777 (N_9777,N_8992,N_8485);
and U9778 (N_9778,N_8791,N_8909);
or U9779 (N_9779,N_8302,N_8249);
nor U9780 (N_9780,N_8445,N_8054);
or U9781 (N_9781,N_8331,N_8055);
nand U9782 (N_9782,N_8243,N_8931);
nor U9783 (N_9783,N_8771,N_8115);
and U9784 (N_9784,N_8753,N_8486);
or U9785 (N_9785,N_8382,N_8613);
nor U9786 (N_9786,N_8498,N_8357);
or U9787 (N_9787,N_8913,N_8743);
nand U9788 (N_9788,N_8135,N_8988);
nor U9789 (N_9789,N_8168,N_8006);
nand U9790 (N_9790,N_8458,N_8499);
or U9791 (N_9791,N_8866,N_8840);
nand U9792 (N_9792,N_8857,N_8565);
and U9793 (N_9793,N_8589,N_8721);
nand U9794 (N_9794,N_8054,N_8695);
nand U9795 (N_9795,N_8437,N_8919);
nor U9796 (N_9796,N_8520,N_8472);
nand U9797 (N_9797,N_8339,N_8411);
nand U9798 (N_9798,N_8980,N_8808);
nand U9799 (N_9799,N_8857,N_8990);
nand U9800 (N_9800,N_8599,N_8103);
or U9801 (N_9801,N_8873,N_8682);
nand U9802 (N_9802,N_8191,N_8335);
and U9803 (N_9803,N_8708,N_8715);
nor U9804 (N_9804,N_8767,N_8602);
or U9805 (N_9805,N_8939,N_8937);
and U9806 (N_9806,N_8755,N_8329);
and U9807 (N_9807,N_8413,N_8843);
nor U9808 (N_9808,N_8337,N_8091);
and U9809 (N_9809,N_8330,N_8369);
nor U9810 (N_9810,N_8009,N_8969);
or U9811 (N_9811,N_8681,N_8689);
nand U9812 (N_9812,N_8094,N_8527);
or U9813 (N_9813,N_8615,N_8898);
and U9814 (N_9814,N_8377,N_8849);
nand U9815 (N_9815,N_8963,N_8087);
and U9816 (N_9816,N_8732,N_8687);
or U9817 (N_9817,N_8360,N_8661);
nor U9818 (N_9818,N_8166,N_8770);
and U9819 (N_9819,N_8999,N_8133);
nand U9820 (N_9820,N_8757,N_8103);
nand U9821 (N_9821,N_8879,N_8546);
and U9822 (N_9822,N_8537,N_8492);
nor U9823 (N_9823,N_8915,N_8891);
and U9824 (N_9824,N_8163,N_8239);
nand U9825 (N_9825,N_8184,N_8340);
nand U9826 (N_9826,N_8108,N_8590);
nor U9827 (N_9827,N_8987,N_8341);
and U9828 (N_9828,N_8943,N_8693);
and U9829 (N_9829,N_8812,N_8324);
nand U9830 (N_9830,N_8522,N_8001);
nor U9831 (N_9831,N_8490,N_8147);
xnor U9832 (N_9832,N_8866,N_8829);
nand U9833 (N_9833,N_8038,N_8009);
nand U9834 (N_9834,N_8332,N_8196);
or U9835 (N_9835,N_8940,N_8033);
nand U9836 (N_9836,N_8582,N_8902);
and U9837 (N_9837,N_8965,N_8833);
or U9838 (N_9838,N_8304,N_8052);
nor U9839 (N_9839,N_8052,N_8944);
or U9840 (N_9840,N_8221,N_8308);
or U9841 (N_9841,N_8261,N_8752);
or U9842 (N_9842,N_8075,N_8680);
or U9843 (N_9843,N_8270,N_8377);
and U9844 (N_9844,N_8101,N_8198);
nand U9845 (N_9845,N_8668,N_8508);
or U9846 (N_9846,N_8592,N_8775);
nand U9847 (N_9847,N_8084,N_8273);
or U9848 (N_9848,N_8454,N_8225);
and U9849 (N_9849,N_8088,N_8632);
and U9850 (N_9850,N_8812,N_8224);
or U9851 (N_9851,N_8282,N_8443);
and U9852 (N_9852,N_8293,N_8578);
nor U9853 (N_9853,N_8062,N_8692);
xnor U9854 (N_9854,N_8308,N_8933);
and U9855 (N_9855,N_8461,N_8965);
or U9856 (N_9856,N_8987,N_8532);
or U9857 (N_9857,N_8772,N_8427);
and U9858 (N_9858,N_8775,N_8358);
or U9859 (N_9859,N_8131,N_8504);
nand U9860 (N_9860,N_8844,N_8630);
or U9861 (N_9861,N_8084,N_8601);
and U9862 (N_9862,N_8698,N_8106);
nand U9863 (N_9863,N_8117,N_8442);
nor U9864 (N_9864,N_8025,N_8428);
xor U9865 (N_9865,N_8776,N_8944);
and U9866 (N_9866,N_8424,N_8024);
and U9867 (N_9867,N_8803,N_8323);
and U9868 (N_9868,N_8169,N_8108);
nand U9869 (N_9869,N_8242,N_8154);
or U9870 (N_9870,N_8947,N_8688);
nand U9871 (N_9871,N_8186,N_8900);
nand U9872 (N_9872,N_8845,N_8949);
or U9873 (N_9873,N_8343,N_8732);
nor U9874 (N_9874,N_8863,N_8939);
nand U9875 (N_9875,N_8442,N_8157);
nand U9876 (N_9876,N_8967,N_8953);
and U9877 (N_9877,N_8702,N_8036);
nor U9878 (N_9878,N_8405,N_8584);
and U9879 (N_9879,N_8291,N_8553);
nor U9880 (N_9880,N_8815,N_8535);
or U9881 (N_9881,N_8606,N_8377);
nand U9882 (N_9882,N_8613,N_8276);
nor U9883 (N_9883,N_8185,N_8369);
nand U9884 (N_9884,N_8898,N_8097);
or U9885 (N_9885,N_8457,N_8117);
or U9886 (N_9886,N_8700,N_8410);
nand U9887 (N_9887,N_8621,N_8230);
and U9888 (N_9888,N_8486,N_8179);
and U9889 (N_9889,N_8438,N_8307);
xnor U9890 (N_9890,N_8415,N_8900);
nor U9891 (N_9891,N_8258,N_8529);
and U9892 (N_9892,N_8231,N_8597);
xor U9893 (N_9893,N_8302,N_8176);
nand U9894 (N_9894,N_8339,N_8764);
and U9895 (N_9895,N_8069,N_8811);
and U9896 (N_9896,N_8666,N_8078);
nor U9897 (N_9897,N_8131,N_8457);
nand U9898 (N_9898,N_8127,N_8561);
and U9899 (N_9899,N_8957,N_8176);
or U9900 (N_9900,N_8644,N_8735);
xnor U9901 (N_9901,N_8868,N_8672);
nor U9902 (N_9902,N_8454,N_8390);
nand U9903 (N_9903,N_8562,N_8891);
or U9904 (N_9904,N_8643,N_8423);
nor U9905 (N_9905,N_8339,N_8587);
or U9906 (N_9906,N_8746,N_8820);
nand U9907 (N_9907,N_8430,N_8121);
or U9908 (N_9908,N_8431,N_8937);
and U9909 (N_9909,N_8470,N_8039);
nor U9910 (N_9910,N_8047,N_8754);
nor U9911 (N_9911,N_8217,N_8378);
or U9912 (N_9912,N_8720,N_8784);
and U9913 (N_9913,N_8724,N_8818);
and U9914 (N_9914,N_8963,N_8118);
nor U9915 (N_9915,N_8380,N_8834);
and U9916 (N_9916,N_8891,N_8643);
and U9917 (N_9917,N_8454,N_8805);
nor U9918 (N_9918,N_8665,N_8654);
nand U9919 (N_9919,N_8909,N_8300);
nand U9920 (N_9920,N_8240,N_8870);
or U9921 (N_9921,N_8461,N_8820);
and U9922 (N_9922,N_8043,N_8378);
or U9923 (N_9923,N_8408,N_8603);
nor U9924 (N_9924,N_8971,N_8659);
nor U9925 (N_9925,N_8362,N_8963);
and U9926 (N_9926,N_8662,N_8315);
nand U9927 (N_9927,N_8459,N_8772);
xnor U9928 (N_9928,N_8110,N_8920);
nor U9929 (N_9929,N_8098,N_8783);
xnor U9930 (N_9930,N_8987,N_8688);
and U9931 (N_9931,N_8691,N_8688);
nor U9932 (N_9932,N_8301,N_8917);
nor U9933 (N_9933,N_8166,N_8702);
nand U9934 (N_9934,N_8447,N_8760);
and U9935 (N_9935,N_8144,N_8633);
nand U9936 (N_9936,N_8226,N_8427);
or U9937 (N_9937,N_8616,N_8382);
nand U9938 (N_9938,N_8661,N_8312);
xor U9939 (N_9939,N_8134,N_8312);
nor U9940 (N_9940,N_8920,N_8038);
nor U9941 (N_9941,N_8729,N_8691);
xnor U9942 (N_9942,N_8598,N_8382);
nor U9943 (N_9943,N_8451,N_8715);
and U9944 (N_9944,N_8564,N_8631);
or U9945 (N_9945,N_8909,N_8990);
nand U9946 (N_9946,N_8628,N_8433);
nand U9947 (N_9947,N_8637,N_8522);
or U9948 (N_9948,N_8523,N_8421);
nand U9949 (N_9949,N_8853,N_8285);
and U9950 (N_9950,N_8935,N_8782);
nor U9951 (N_9951,N_8216,N_8919);
and U9952 (N_9952,N_8102,N_8742);
nand U9953 (N_9953,N_8631,N_8686);
and U9954 (N_9954,N_8092,N_8014);
or U9955 (N_9955,N_8322,N_8863);
nand U9956 (N_9956,N_8959,N_8103);
or U9957 (N_9957,N_8116,N_8411);
or U9958 (N_9958,N_8181,N_8313);
or U9959 (N_9959,N_8741,N_8544);
or U9960 (N_9960,N_8997,N_8324);
and U9961 (N_9961,N_8542,N_8023);
nand U9962 (N_9962,N_8848,N_8378);
or U9963 (N_9963,N_8246,N_8704);
and U9964 (N_9964,N_8036,N_8635);
nor U9965 (N_9965,N_8120,N_8872);
nand U9966 (N_9966,N_8740,N_8483);
or U9967 (N_9967,N_8444,N_8625);
and U9968 (N_9968,N_8878,N_8649);
nor U9969 (N_9969,N_8487,N_8625);
nand U9970 (N_9970,N_8233,N_8406);
or U9971 (N_9971,N_8370,N_8197);
nor U9972 (N_9972,N_8984,N_8145);
and U9973 (N_9973,N_8558,N_8777);
nor U9974 (N_9974,N_8283,N_8972);
nor U9975 (N_9975,N_8405,N_8696);
nor U9976 (N_9976,N_8491,N_8216);
and U9977 (N_9977,N_8533,N_8011);
and U9978 (N_9978,N_8845,N_8086);
nor U9979 (N_9979,N_8705,N_8323);
nand U9980 (N_9980,N_8981,N_8837);
or U9981 (N_9981,N_8713,N_8513);
and U9982 (N_9982,N_8404,N_8314);
and U9983 (N_9983,N_8436,N_8185);
nand U9984 (N_9984,N_8163,N_8014);
nor U9985 (N_9985,N_8881,N_8939);
nor U9986 (N_9986,N_8160,N_8239);
nand U9987 (N_9987,N_8599,N_8463);
nor U9988 (N_9988,N_8488,N_8645);
and U9989 (N_9989,N_8143,N_8233);
nor U9990 (N_9990,N_8208,N_8216);
nand U9991 (N_9991,N_8904,N_8200);
nand U9992 (N_9992,N_8041,N_8610);
and U9993 (N_9993,N_8125,N_8649);
or U9994 (N_9994,N_8708,N_8055);
and U9995 (N_9995,N_8413,N_8253);
and U9996 (N_9996,N_8194,N_8804);
and U9997 (N_9997,N_8936,N_8203);
nand U9998 (N_9998,N_8989,N_8047);
or U9999 (N_9999,N_8213,N_8759);
or UO_0 (O_0,N_9988,N_9272);
nor UO_1 (O_1,N_9424,N_9570);
xor UO_2 (O_2,N_9754,N_9886);
nand UO_3 (O_3,N_9611,N_9544);
nand UO_4 (O_4,N_9769,N_9857);
nand UO_5 (O_5,N_9014,N_9048);
nand UO_6 (O_6,N_9280,N_9294);
or UO_7 (O_7,N_9936,N_9697);
or UO_8 (O_8,N_9281,N_9352);
and UO_9 (O_9,N_9856,N_9070);
or UO_10 (O_10,N_9493,N_9121);
nand UO_11 (O_11,N_9358,N_9390);
or UO_12 (O_12,N_9053,N_9598);
nor UO_13 (O_13,N_9098,N_9238);
nor UO_14 (O_14,N_9533,N_9197);
and UO_15 (O_15,N_9976,N_9799);
or UO_16 (O_16,N_9711,N_9196);
or UO_17 (O_17,N_9442,N_9681);
and UO_18 (O_18,N_9163,N_9762);
and UO_19 (O_19,N_9554,N_9908);
or UO_20 (O_20,N_9470,N_9170);
or UO_21 (O_21,N_9339,N_9379);
and UO_22 (O_22,N_9334,N_9228);
nor UO_23 (O_23,N_9964,N_9518);
or UO_24 (O_24,N_9250,N_9046);
nand UO_25 (O_25,N_9993,N_9188);
nand UO_26 (O_26,N_9378,N_9991);
or UO_27 (O_27,N_9286,N_9017);
or UO_28 (O_28,N_9782,N_9589);
nor UO_29 (O_29,N_9372,N_9296);
and UO_30 (O_30,N_9135,N_9956);
and UO_31 (O_31,N_9109,N_9235);
nand UO_32 (O_32,N_9313,N_9282);
nand UO_33 (O_33,N_9445,N_9409);
or UO_34 (O_34,N_9467,N_9822);
and UO_35 (O_35,N_9316,N_9410);
nor UO_36 (O_36,N_9088,N_9577);
and UO_37 (O_37,N_9978,N_9021);
nand UO_38 (O_38,N_9726,N_9745);
and UO_39 (O_39,N_9325,N_9970);
or UO_40 (O_40,N_9877,N_9096);
and UO_41 (O_41,N_9116,N_9317);
nor UO_42 (O_42,N_9278,N_9226);
nand UO_43 (O_43,N_9860,N_9093);
nor UO_44 (O_44,N_9688,N_9568);
xor UO_45 (O_45,N_9214,N_9308);
nand UO_46 (O_46,N_9086,N_9350);
nand UO_47 (O_47,N_9547,N_9950);
nor UO_48 (O_48,N_9312,N_9175);
nor UO_49 (O_49,N_9905,N_9418);
nand UO_50 (O_50,N_9402,N_9172);
nand UO_51 (O_51,N_9451,N_9225);
nor UO_52 (O_52,N_9403,N_9232);
nand UO_53 (O_53,N_9985,N_9663);
or UO_54 (O_54,N_9536,N_9244);
nand UO_55 (O_55,N_9692,N_9671);
or UO_56 (O_56,N_9099,N_9884);
or UO_57 (O_57,N_9833,N_9474);
or UO_58 (O_58,N_9345,N_9842);
nor UO_59 (O_59,N_9038,N_9215);
nor UO_60 (O_60,N_9369,N_9731);
nor UO_61 (O_61,N_9505,N_9182);
nand UO_62 (O_62,N_9440,N_9847);
or UO_63 (O_63,N_9887,N_9254);
nor UO_64 (O_64,N_9443,N_9210);
and UO_65 (O_65,N_9789,N_9944);
and UO_66 (O_66,N_9179,N_9617);
nand UO_67 (O_67,N_9145,N_9699);
nand UO_68 (O_68,N_9000,N_9634);
xor UO_69 (O_69,N_9768,N_9954);
and UO_70 (O_70,N_9784,N_9728);
or UO_71 (O_71,N_9147,N_9411);
nand UO_72 (O_72,N_9625,N_9230);
nand UO_73 (O_73,N_9113,N_9817);
nand UO_74 (O_74,N_9690,N_9776);
or UO_75 (O_75,N_9723,N_9426);
and UO_76 (O_76,N_9185,N_9119);
or UO_77 (O_77,N_9716,N_9268);
nor UO_78 (O_78,N_9526,N_9169);
nand UO_79 (O_79,N_9330,N_9881);
or UO_80 (O_80,N_9868,N_9123);
and UO_81 (O_81,N_9669,N_9560);
or UO_82 (O_82,N_9340,N_9042);
xor UO_83 (O_83,N_9298,N_9024);
or UO_84 (O_84,N_9227,N_9851);
nor UO_85 (O_85,N_9320,N_9828);
or UO_86 (O_86,N_9090,N_9200);
nor UO_87 (O_87,N_9329,N_9331);
nor UO_88 (O_88,N_9208,N_9069);
and UO_89 (O_89,N_9551,N_9914);
nand UO_90 (O_90,N_9148,N_9387);
and UO_91 (O_91,N_9303,N_9391);
nand UO_92 (O_92,N_9456,N_9673);
nor UO_93 (O_93,N_9818,N_9190);
and UO_94 (O_94,N_9804,N_9894);
nand UO_95 (O_95,N_9134,N_9370);
or UO_96 (O_96,N_9261,N_9165);
nand UO_97 (O_97,N_9029,N_9622);
and UO_98 (O_98,N_9830,N_9381);
or UO_99 (O_99,N_9707,N_9650);
and UO_100 (O_100,N_9582,N_9623);
nor UO_101 (O_101,N_9873,N_9735);
and UO_102 (O_102,N_9428,N_9146);
nand UO_103 (O_103,N_9421,N_9010);
nand UO_104 (O_104,N_9118,N_9760);
nor UO_105 (O_105,N_9502,N_9785);
nor UO_106 (O_106,N_9160,N_9618);
and UO_107 (O_107,N_9449,N_9721);
and UO_108 (O_108,N_9981,N_9034);
nand UO_109 (O_109,N_9064,N_9327);
nor UO_110 (O_110,N_9620,N_9357);
nand UO_111 (O_111,N_9504,N_9246);
nor UO_112 (O_112,N_9880,N_9888);
and UO_113 (O_113,N_9071,N_9930);
nor UO_114 (O_114,N_9561,N_9571);
nor UO_115 (O_115,N_9394,N_9102);
nor UO_116 (O_116,N_9496,N_9239);
or UO_117 (O_117,N_9791,N_9766);
nor UO_118 (O_118,N_9904,N_9129);
or UO_119 (O_119,N_9051,N_9600);
nor UO_120 (O_120,N_9968,N_9380);
nor UO_121 (O_121,N_9565,N_9780);
or UO_122 (O_122,N_9104,N_9992);
and UO_123 (O_123,N_9212,N_9601);
or UO_124 (O_124,N_9987,N_9866);
nand UO_125 (O_125,N_9702,N_9872);
and UO_126 (O_126,N_9427,N_9157);
or UO_127 (O_127,N_9685,N_9986);
or UO_128 (O_128,N_9299,N_9657);
nand UO_129 (O_129,N_9967,N_9245);
nor UO_130 (O_130,N_9288,N_9243);
or UO_131 (O_131,N_9750,N_9095);
nand UO_132 (O_132,N_9293,N_9258);
nand UO_133 (O_133,N_9771,N_9656);
nor UO_134 (O_134,N_9259,N_9389);
nand UO_135 (O_135,N_9062,N_9265);
and UO_136 (O_136,N_9948,N_9942);
or UO_137 (O_137,N_9759,N_9337);
nor UO_138 (O_138,N_9018,N_9183);
and UO_139 (O_139,N_9709,N_9068);
nand UO_140 (O_140,N_9342,N_9525);
nor UO_141 (O_141,N_9187,N_9624);
nand UO_142 (O_142,N_9002,N_9036);
nand UO_143 (O_143,N_9945,N_9925);
nand UO_144 (O_144,N_9139,N_9162);
and UO_145 (O_145,N_9962,N_9315);
nor UO_146 (O_146,N_9635,N_9700);
nand UO_147 (O_147,N_9111,N_9028);
and UO_148 (O_148,N_9026,N_9097);
or UO_149 (O_149,N_9468,N_9471);
and UO_150 (O_150,N_9575,N_9608);
or UO_151 (O_151,N_9112,N_9736);
nand UO_152 (O_152,N_9066,N_9810);
nand UO_153 (O_153,N_9395,N_9220);
nand UO_154 (O_154,N_9501,N_9616);
nor UO_155 (O_155,N_9730,N_9740);
and UO_156 (O_156,N_9485,N_9779);
nor UO_157 (O_157,N_9016,N_9291);
nand UO_158 (O_158,N_9845,N_9943);
nor UO_159 (O_159,N_9841,N_9871);
and UO_160 (O_160,N_9934,N_9412);
or UO_161 (O_161,N_9264,N_9903);
and UO_162 (O_162,N_9453,N_9549);
nor UO_163 (O_163,N_9269,N_9285);
nand UO_164 (O_164,N_9605,N_9995);
and UO_165 (O_165,N_9676,N_9802);
and UO_166 (O_166,N_9240,N_9606);
nand UO_167 (O_167,N_9863,N_9492);
nor UO_168 (O_168,N_9741,N_9138);
or UO_169 (O_169,N_9081,N_9279);
nor UO_170 (O_170,N_9341,N_9400);
or UO_171 (O_171,N_9631,N_9940);
nand UO_172 (O_172,N_9130,N_9977);
nand UO_173 (O_173,N_9743,N_9592);
nor UO_174 (O_174,N_9870,N_9722);
nand UO_175 (O_175,N_9224,N_9167);
nor UO_176 (O_176,N_9216,N_9209);
nor UO_177 (O_177,N_9161,N_9717);
and UO_178 (O_178,N_9392,N_9824);
and UO_179 (O_179,N_9637,N_9475);
nand UO_180 (O_180,N_9057,N_9490);
nor UO_181 (O_181,N_9304,N_9798);
nor UO_182 (O_182,N_9698,N_9434);
and UO_183 (O_183,N_9647,N_9867);
nand UO_184 (O_184,N_9953,N_9457);
nor UO_185 (O_185,N_9022,N_9898);
nand UO_186 (O_186,N_9191,N_9301);
nand UO_187 (O_187,N_9194,N_9846);
and UO_188 (O_188,N_9030,N_9687);
or UO_189 (O_189,N_9719,N_9439);
and UO_190 (O_190,N_9176,N_9125);
nand UO_191 (O_191,N_9506,N_9251);
or UO_192 (O_192,N_9480,N_9488);
nand UO_193 (O_193,N_9660,N_9491);
or UO_194 (O_194,N_9843,N_9523);
nand UO_195 (O_195,N_9919,N_9832);
and UO_196 (O_196,N_9609,N_9563);
nand UO_197 (O_197,N_9039,N_9756);
or UO_198 (O_198,N_9466,N_9874);
or UO_199 (O_199,N_9052,N_9640);
and UO_200 (O_200,N_9537,N_9534);
nand UO_201 (O_201,N_9961,N_9423);
or UO_202 (O_202,N_9477,N_9154);
and UO_203 (O_203,N_9861,N_9420);
xor UO_204 (O_204,N_9626,N_9969);
nor UO_205 (O_205,N_9654,N_9393);
nor UO_206 (O_206,N_9614,N_9686);
and UO_207 (O_207,N_9141,N_9946);
nand UO_208 (O_208,N_9503,N_9899);
or UO_209 (O_209,N_9292,N_9748);
or UO_210 (O_210,N_9829,N_9432);
nand UO_211 (O_211,N_9831,N_9023);
nor UO_212 (O_212,N_9757,N_9926);
and UO_213 (O_213,N_9302,N_9584);
or UO_214 (O_214,N_9484,N_9371);
and UO_215 (O_215,N_9207,N_9579);
and UO_216 (O_216,N_9850,N_9783);
nand UO_217 (O_217,N_9438,N_9865);
nor UO_218 (O_218,N_9966,N_9181);
nor UO_219 (O_219,N_9581,N_9452);
nand UO_220 (O_220,N_9234,N_9001);
and UO_221 (O_221,N_9297,N_9939);
nand UO_222 (O_222,N_9083,N_9263);
nand UO_223 (O_223,N_9838,N_9694);
and UO_224 (O_224,N_9376,N_9364);
nand UO_225 (O_225,N_9295,N_9218);
and UO_226 (O_226,N_9255,N_9604);
nand UO_227 (O_227,N_9636,N_9100);
and UO_228 (O_228,N_9027,N_9260);
and UO_229 (O_229,N_9009,N_9419);
nand UO_230 (O_230,N_9662,N_9415);
nand UO_231 (O_231,N_9284,N_9174);
nor UO_232 (O_232,N_9487,N_9892);
nand UO_233 (O_233,N_9035,N_9907);
nand UO_234 (O_234,N_9947,N_9155);
nand UO_235 (O_235,N_9497,N_9429);
xor UO_236 (O_236,N_9924,N_9704);
or UO_237 (O_237,N_9007,N_9450);
nor UO_238 (O_238,N_9535,N_9511);
nand UO_239 (O_239,N_9204,N_9803);
nor UO_240 (O_240,N_9094,N_9222);
nand UO_241 (O_241,N_9374,N_9955);
nor UO_242 (O_242,N_9909,N_9596);
nor UO_243 (O_243,N_9540,N_9834);
nor UO_244 (O_244,N_9679,N_9971);
nand UO_245 (O_245,N_9712,N_9201);
or UO_246 (O_246,N_9463,N_9593);
nand UO_247 (O_247,N_9556,N_9347);
nor UO_248 (O_248,N_9151,N_9353);
nand UO_249 (O_249,N_9801,N_9765);
nand UO_250 (O_250,N_9580,N_9812);
and UO_251 (O_251,N_9965,N_9247);
nand UO_252 (O_252,N_9764,N_9854);
or UO_253 (O_253,N_9082,N_9911);
nand UO_254 (O_254,N_9217,N_9641);
and UO_255 (O_255,N_9266,N_9049);
nand UO_256 (O_256,N_9132,N_9011);
and UO_257 (O_257,N_9460,N_9495);
and UO_258 (O_258,N_9621,N_9823);
nand UO_259 (O_259,N_9963,N_9077);
nor UO_260 (O_260,N_9249,N_9890);
nor UO_261 (O_261,N_9314,N_9332);
or UO_262 (O_262,N_9852,N_9586);
and UO_263 (O_263,N_9032,N_9318);
nor UO_264 (O_264,N_9486,N_9328);
and UO_265 (O_265,N_9508,N_9569);
or UO_266 (O_266,N_9054,N_9629);
nor UO_267 (O_267,N_9793,N_9652);
or UO_268 (O_268,N_9043,N_9221);
nand UO_269 (O_269,N_9696,N_9891);
or UO_270 (O_270,N_9408,N_9105);
nand UO_271 (O_271,N_9058,N_9336);
nand UO_272 (O_272,N_9144,N_9464);
and UO_273 (O_273,N_9516,N_9814);
nor UO_274 (O_274,N_9072,N_9820);
and UO_275 (O_275,N_9189,N_9177);
and UO_276 (O_276,N_9562,N_9806);
and UO_277 (O_277,N_9404,N_9859);
nor UO_278 (O_278,N_9642,N_9733);
or UO_279 (O_279,N_9559,N_9273);
nand UO_280 (O_280,N_9658,N_9396);
xor UO_281 (O_281,N_9816,N_9128);
nand UO_282 (O_282,N_9758,N_9153);
nor UO_283 (O_283,N_9283,N_9896);
or UO_284 (O_284,N_9732,N_9665);
or UO_285 (O_285,N_9233,N_9931);
nand UO_286 (O_286,N_9725,N_9276);
nand UO_287 (O_287,N_9984,N_9373);
nor UO_288 (O_288,N_9786,N_9590);
nand UO_289 (O_289,N_9938,N_9045);
nand UO_290 (O_290,N_9897,N_9729);
or UO_291 (O_291,N_9761,N_9479);
nor UO_292 (O_292,N_9513,N_9689);
and UO_293 (O_293,N_9557,N_9158);
or UO_294 (O_294,N_9524,N_9869);
and UO_295 (O_295,N_9229,N_9517);
or UO_296 (O_296,N_9649,N_9444);
nor UO_297 (O_297,N_9693,N_9794);
nor UO_298 (O_298,N_9033,N_9499);
nand UO_299 (O_299,N_9792,N_9980);
and UO_300 (O_300,N_9242,N_9015);
and UO_301 (O_301,N_9753,N_9489);
and UO_302 (O_302,N_9110,N_9973);
nand UO_303 (O_303,N_9773,N_9781);
xor UO_304 (O_304,N_9431,N_9482);
nand UO_305 (O_305,N_9885,N_9815);
or UO_306 (O_306,N_9882,N_9531);
nand UO_307 (O_307,N_9257,N_9178);
nand UO_308 (O_308,N_9084,N_9414);
and UO_309 (O_309,N_9734,N_9025);
or UO_310 (O_310,N_9858,N_9742);
or UO_311 (O_311,N_9935,N_9691);
or UO_312 (O_312,N_9975,N_9136);
and UO_313 (O_313,N_9927,N_9458);
nand UO_314 (O_314,N_9277,N_9708);
and UO_315 (O_315,N_9576,N_9333);
and UO_316 (O_316,N_9840,N_9076);
or UO_317 (O_317,N_9448,N_9368);
or UO_318 (O_318,N_9682,N_9323);
and UO_319 (O_319,N_9120,N_9900);
nand UO_320 (O_320,N_9433,N_9951);
nand UO_321 (O_321,N_9117,N_9202);
or UO_322 (O_322,N_9115,N_9530);
nand UO_323 (O_323,N_9041,N_9529);
and UO_324 (O_324,N_9594,N_9603);
or UO_325 (O_325,N_9005,N_9008);
and UO_326 (O_326,N_9542,N_9122);
nor UO_327 (O_327,N_9630,N_9289);
and UO_328 (O_328,N_9720,N_9619);
nor UO_329 (O_329,N_9223,N_9338);
nand UO_330 (O_330,N_9349,N_9548);
and UO_331 (O_331,N_9566,N_9050);
nor UO_332 (O_332,N_9195,N_9319);
nand UO_333 (O_333,N_9979,N_9648);
nand UO_334 (O_334,N_9478,N_9455);
nand UO_335 (O_335,N_9821,N_9003);
nand UO_336 (O_336,N_9300,N_9994);
and UO_337 (O_337,N_9646,N_9500);
or UO_338 (O_338,N_9990,N_9365);
or UO_339 (O_339,N_9186,N_9004);
or UO_340 (O_340,N_9539,N_9958);
nand UO_341 (O_341,N_9055,N_9895);
and UO_342 (O_342,N_9510,N_9819);
nor UO_343 (O_343,N_9521,N_9211);
nand UO_344 (O_344,N_9628,N_9164);
xor UO_345 (O_345,N_9324,N_9080);
or UO_346 (O_346,N_9675,N_9737);
and UO_347 (O_347,N_9416,N_9695);
and UO_348 (O_348,N_9031,N_9775);
nand UO_349 (O_349,N_9913,N_9047);
nor UO_350 (O_350,N_9974,N_9362);
nor UO_351 (O_351,N_9344,N_9398);
or UO_352 (O_352,N_9447,N_9901);
and UO_353 (O_353,N_9929,N_9638);
and UO_354 (O_354,N_9063,N_9354);
and UO_355 (O_355,N_9126,N_9883);
or UO_356 (O_356,N_9715,N_9321);
nand UO_357 (O_357,N_9231,N_9836);
nand UO_358 (O_358,N_9399,N_9326);
nand UO_359 (O_359,N_9351,N_9275);
and UO_360 (O_360,N_9583,N_9013);
nor UO_361 (O_361,N_9875,N_9643);
and UO_362 (O_362,N_9797,N_9684);
or UO_363 (O_363,N_9385,N_9397);
or UO_364 (O_364,N_9808,N_9382);
and UO_365 (O_365,N_9607,N_9472);
nor UO_366 (O_366,N_9166,N_9952);
nand UO_367 (O_367,N_9714,N_9790);
nand UO_368 (O_368,N_9644,N_9476);
or UO_369 (O_369,N_9168,N_9366);
and UO_370 (O_370,N_9921,N_9307);
nand UO_371 (O_371,N_9853,N_9778);
nand UO_372 (O_372,N_9879,N_9989);
or UO_373 (O_373,N_9067,N_9912);
and UO_374 (O_374,N_9848,N_9527);
or UO_375 (O_375,N_9664,N_9079);
nand UO_376 (O_376,N_9384,N_9106);
or UO_377 (O_377,N_9772,N_9143);
or UO_378 (O_378,N_9546,N_9602);
and UO_379 (O_379,N_9550,N_9795);
or UO_380 (O_380,N_9668,N_9755);
nand UO_381 (O_381,N_9061,N_9928);
and UO_382 (O_382,N_9767,N_9587);
and UO_383 (O_383,N_9494,N_9206);
or UO_384 (O_384,N_9674,N_9599);
nor UO_385 (O_385,N_9091,N_9588);
nand UO_386 (O_386,N_9271,N_9441);
nand UO_387 (O_387,N_9078,N_9998);
and UO_388 (O_388,N_9407,N_9809);
nand UO_389 (O_389,N_9667,N_9902);
or UO_390 (O_390,N_9835,N_9290);
nor UO_391 (O_391,N_9763,N_9959);
and UO_392 (O_392,N_9555,N_9983);
or UO_393 (O_393,N_9459,N_9922);
nand UO_394 (O_394,N_9252,N_9519);
and UO_395 (O_395,N_9615,N_9469);
and UO_396 (O_396,N_9538,N_9101);
nor UO_397 (O_397,N_9972,N_9591);
and UO_398 (O_398,N_9683,N_9572);
and UO_399 (O_399,N_9124,N_9465);
nand UO_400 (O_400,N_9744,N_9253);
and UO_401 (O_401,N_9425,N_9149);
nor UO_402 (O_402,N_9788,N_9595);
nor UO_403 (O_403,N_9363,N_9670);
or UO_404 (O_404,N_9889,N_9906);
and UO_405 (O_405,N_9862,N_9713);
nor UO_406 (O_406,N_9661,N_9309);
and UO_407 (O_407,N_9114,N_9677);
nand UO_408 (O_408,N_9405,N_9545);
and UO_409 (O_409,N_9864,N_9335);
or UO_410 (O_410,N_9127,N_9205);
nand UO_411 (O_411,N_9567,N_9346);
nand UO_412 (O_412,N_9839,N_9982);
xnor UO_413 (O_413,N_9639,N_9180);
nand UO_414 (O_414,N_9270,N_9203);
nand UO_415 (O_415,N_9915,N_9150);
or UO_416 (O_416,N_9878,N_9483);
or UO_417 (O_417,N_9893,N_9311);
nor UO_418 (O_418,N_9219,N_9612);
or UO_419 (O_419,N_9171,N_9108);
nand UO_420 (O_420,N_9645,N_9937);
or UO_421 (O_421,N_9800,N_9193);
nor UO_422 (O_422,N_9932,N_9355);
and UO_423 (O_423,N_9241,N_9262);
and UO_424 (O_424,N_9655,N_9844);
or UO_425 (O_425,N_9553,N_9633);
and UO_426 (O_426,N_9107,N_9787);
or UO_427 (O_427,N_9543,N_9359);
nand UO_428 (O_428,N_9705,N_9564);
nor UO_429 (O_429,N_9876,N_9481);
or UO_430 (O_430,N_9274,N_9044);
nor UO_431 (O_431,N_9701,N_9627);
and UO_432 (O_432,N_9375,N_9739);
nand UO_433 (O_433,N_9040,N_9377);
and UO_434 (O_434,N_9306,N_9020);
nand UO_435 (O_435,N_9747,N_9159);
nor UO_436 (O_436,N_9059,N_9140);
and UO_437 (O_437,N_9446,N_9092);
and UO_438 (O_438,N_9383,N_9706);
xnor UO_439 (O_439,N_9672,N_9827);
nand UO_440 (O_440,N_9522,N_9916);
and UO_441 (O_441,N_9552,N_9461);
nor UO_442 (O_442,N_9388,N_9597);
or UO_443 (O_443,N_9436,N_9997);
or UO_444 (O_444,N_9498,N_9287);
or UO_445 (O_445,N_9703,N_9777);
nand UO_446 (O_446,N_9678,N_9198);
or UO_447 (O_447,N_9367,N_9343);
and UO_448 (O_448,N_9417,N_9413);
nor UO_449 (O_449,N_9152,N_9386);
and UO_450 (O_450,N_9360,N_9710);
and UO_451 (O_451,N_9133,N_9213);
and UO_452 (O_452,N_9019,N_9796);
and UO_453 (O_453,N_9653,N_9356);
and UO_454 (O_454,N_9949,N_9751);
nor UO_455 (O_455,N_9322,N_9430);
and UO_456 (O_456,N_9770,N_9060);
nor UO_457 (O_457,N_9941,N_9056);
nor UO_458 (O_458,N_9917,N_9541);
nand UO_459 (O_459,N_9087,N_9574);
nor UO_460 (O_460,N_9613,N_9923);
or UO_461 (O_461,N_9957,N_9462);
nor UO_462 (O_462,N_9825,N_9173);
nor UO_463 (O_463,N_9837,N_9573);
or UO_464 (O_464,N_9774,N_9738);
and UO_465 (O_465,N_9361,N_9437);
nand UO_466 (O_466,N_9142,N_9267);
nor UO_467 (O_467,N_9752,N_9131);
nand UO_468 (O_468,N_9507,N_9813);
nor UO_469 (O_469,N_9422,N_9960);
nor UO_470 (O_470,N_9718,N_9724);
and UO_471 (O_471,N_9920,N_9406);
or UO_472 (O_472,N_9727,N_9849);
nand UO_473 (O_473,N_9933,N_9305);
nor UO_474 (O_474,N_9085,N_9512);
or UO_475 (O_475,N_9666,N_9089);
or UO_476 (O_476,N_9012,N_9075);
or UO_477 (O_477,N_9509,N_9749);
nor UO_478 (O_478,N_9473,N_9074);
or UO_479 (O_479,N_9184,N_9918);
nor UO_480 (O_480,N_9401,N_9632);
or UO_481 (O_481,N_9558,N_9236);
nand UO_482 (O_482,N_9248,N_9585);
nor UO_483 (O_483,N_9192,N_9746);
or UO_484 (O_484,N_9256,N_9578);
nand UO_485 (O_485,N_9006,N_9999);
and UO_486 (O_486,N_9996,N_9680);
nand UO_487 (O_487,N_9520,N_9811);
or UO_488 (O_488,N_9310,N_9199);
and UO_489 (O_489,N_9037,N_9659);
nor UO_490 (O_490,N_9237,N_9454);
xnor UO_491 (O_491,N_9532,N_9137);
nor UO_492 (O_492,N_9103,N_9435);
nand UO_493 (O_493,N_9156,N_9348);
nor UO_494 (O_494,N_9610,N_9651);
or UO_495 (O_495,N_9805,N_9065);
nand UO_496 (O_496,N_9855,N_9073);
nor UO_497 (O_497,N_9515,N_9807);
and UO_498 (O_498,N_9528,N_9514);
nor UO_499 (O_499,N_9826,N_9910);
or UO_500 (O_500,N_9673,N_9051);
and UO_501 (O_501,N_9661,N_9489);
and UO_502 (O_502,N_9083,N_9519);
nor UO_503 (O_503,N_9752,N_9727);
or UO_504 (O_504,N_9490,N_9627);
or UO_505 (O_505,N_9422,N_9489);
nand UO_506 (O_506,N_9375,N_9107);
nor UO_507 (O_507,N_9769,N_9038);
and UO_508 (O_508,N_9754,N_9180);
nand UO_509 (O_509,N_9394,N_9165);
nand UO_510 (O_510,N_9886,N_9922);
nor UO_511 (O_511,N_9086,N_9912);
or UO_512 (O_512,N_9891,N_9494);
or UO_513 (O_513,N_9845,N_9062);
or UO_514 (O_514,N_9171,N_9718);
nand UO_515 (O_515,N_9539,N_9993);
and UO_516 (O_516,N_9069,N_9488);
nor UO_517 (O_517,N_9801,N_9011);
nand UO_518 (O_518,N_9456,N_9720);
nand UO_519 (O_519,N_9213,N_9963);
or UO_520 (O_520,N_9691,N_9630);
nor UO_521 (O_521,N_9282,N_9196);
nand UO_522 (O_522,N_9175,N_9090);
nand UO_523 (O_523,N_9571,N_9292);
or UO_524 (O_524,N_9034,N_9972);
nor UO_525 (O_525,N_9731,N_9043);
or UO_526 (O_526,N_9963,N_9740);
and UO_527 (O_527,N_9018,N_9126);
nand UO_528 (O_528,N_9771,N_9693);
nand UO_529 (O_529,N_9548,N_9772);
or UO_530 (O_530,N_9829,N_9803);
or UO_531 (O_531,N_9279,N_9558);
or UO_532 (O_532,N_9008,N_9929);
nand UO_533 (O_533,N_9464,N_9135);
nor UO_534 (O_534,N_9162,N_9030);
and UO_535 (O_535,N_9179,N_9839);
and UO_536 (O_536,N_9424,N_9681);
nor UO_537 (O_537,N_9485,N_9266);
and UO_538 (O_538,N_9470,N_9172);
nand UO_539 (O_539,N_9673,N_9049);
and UO_540 (O_540,N_9687,N_9678);
or UO_541 (O_541,N_9039,N_9818);
nor UO_542 (O_542,N_9896,N_9970);
or UO_543 (O_543,N_9385,N_9954);
nand UO_544 (O_544,N_9640,N_9554);
nand UO_545 (O_545,N_9361,N_9896);
or UO_546 (O_546,N_9013,N_9219);
nand UO_547 (O_547,N_9262,N_9822);
or UO_548 (O_548,N_9699,N_9029);
or UO_549 (O_549,N_9941,N_9470);
nor UO_550 (O_550,N_9522,N_9894);
and UO_551 (O_551,N_9072,N_9537);
and UO_552 (O_552,N_9613,N_9325);
nand UO_553 (O_553,N_9514,N_9607);
nand UO_554 (O_554,N_9199,N_9874);
or UO_555 (O_555,N_9755,N_9019);
and UO_556 (O_556,N_9272,N_9710);
nand UO_557 (O_557,N_9807,N_9130);
or UO_558 (O_558,N_9239,N_9816);
nor UO_559 (O_559,N_9874,N_9848);
or UO_560 (O_560,N_9356,N_9422);
nor UO_561 (O_561,N_9053,N_9436);
nor UO_562 (O_562,N_9685,N_9346);
or UO_563 (O_563,N_9623,N_9745);
or UO_564 (O_564,N_9000,N_9855);
and UO_565 (O_565,N_9146,N_9797);
nor UO_566 (O_566,N_9542,N_9696);
nand UO_567 (O_567,N_9439,N_9262);
or UO_568 (O_568,N_9803,N_9441);
or UO_569 (O_569,N_9979,N_9752);
and UO_570 (O_570,N_9660,N_9954);
and UO_571 (O_571,N_9069,N_9790);
nor UO_572 (O_572,N_9222,N_9497);
nor UO_573 (O_573,N_9884,N_9459);
nand UO_574 (O_574,N_9095,N_9224);
nand UO_575 (O_575,N_9754,N_9062);
nand UO_576 (O_576,N_9368,N_9540);
nand UO_577 (O_577,N_9366,N_9417);
and UO_578 (O_578,N_9418,N_9563);
or UO_579 (O_579,N_9341,N_9009);
nor UO_580 (O_580,N_9254,N_9051);
nand UO_581 (O_581,N_9946,N_9620);
nand UO_582 (O_582,N_9474,N_9487);
nand UO_583 (O_583,N_9782,N_9848);
and UO_584 (O_584,N_9682,N_9298);
nor UO_585 (O_585,N_9604,N_9179);
and UO_586 (O_586,N_9628,N_9796);
and UO_587 (O_587,N_9490,N_9958);
nor UO_588 (O_588,N_9882,N_9311);
or UO_589 (O_589,N_9251,N_9118);
or UO_590 (O_590,N_9586,N_9187);
and UO_591 (O_591,N_9167,N_9627);
nand UO_592 (O_592,N_9719,N_9180);
and UO_593 (O_593,N_9527,N_9014);
and UO_594 (O_594,N_9116,N_9830);
and UO_595 (O_595,N_9746,N_9634);
and UO_596 (O_596,N_9689,N_9725);
nand UO_597 (O_597,N_9017,N_9391);
and UO_598 (O_598,N_9207,N_9326);
and UO_599 (O_599,N_9563,N_9714);
and UO_600 (O_600,N_9727,N_9449);
nor UO_601 (O_601,N_9954,N_9612);
nand UO_602 (O_602,N_9584,N_9145);
or UO_603 (O_603,N_9563,N_9105);
nand UO_604 (O_604,N_9242,N_9582);
nor UO_605 (O_605,N_9471,N_9366);
and UO_606 (O_606,N_9208,N_9459);
nor UO_607 (O_607,N_9217,N_9631);
nor UO_608 (O_608,N_9276,N_9747);
nor UO_609 (O_609,N_9949,N_9215);
nand UO_610 (O_610,N_9876,N_9433);
or UO_611 (O_611,N_9376,N_9049);
nor UO_612 (O_612,N_9178,N_9471);
and UO_613 (O_613,N_9923,N_9504);
nor UO_614 (O_614,N_9401,N_9337);
nor UO_615 (O_615,N_9357,N_9537);
or UO_616 (O_616,N_9574,N_9318);
nand UO_617 (O_617,N_9535,N_9071);
or UO_618 (O_618,N_9472,N_9702);
or UO_619 (O_619,N_9239,N_9587);
or UO_620 (O_620,N_9335,N_9257);
and UO_621 (O_621,N_9888,N_9119);
nand UO_622 (O_622,N_9713,N_9468);
and UO_623 (O_623,N_9565,N_9595);
nor UO_624 (O_624,N_9999,N_9462);
or UO_625 (O_625,N_9461,N_9078);
and UO_626 (O_626,N_9283,N_9972);
or UO_627 (O_627,N_9713,N_9769);
nand UO_628 (O_628,N_9554,N_9090);
and UO_629 (O_629,N_9468,N_9647);
nand UO_630 (O_630,N_9107,N_9674);
or UO_631 (O_631,N_9102,N_9068);
nor UO_632 (O_632,N_9901,N_9557);
and UO_633 (O_633,N_9709,N_9115);
nand UO_634 (O_634,N_9764,N_9295);
and UO_635 (O_635,N_9689,N_9015);
nand UO_636 (O_636,N_9079,N_9208);
and UO_637 (O_637,N_9320,N_9415);
and UO_638 (O_638,N_9565,N_9452);
or UO_639 (O_639,N_9833,N_9660);
nor UO_640 (O_640,N_9699,N_9428);
nor UO_641 (O_641,N_9394,N_9602);
and UO_642 (O_642,N_9515,N_9405);
and UO_643 (O_643,N_9933,N_9396);
nand UO_644 (O_644,N_9053,N_9676);
xnor UO_645 (O_645,N_9563,N_9951);
nand UO_646 (O_646,N_9956,N_9280);
or UO_647 (O_647,N_9921,N_9952);
nor UO_648 (O_648,N_9750,N_9467);
nor UO_649 (O_649,N_9710,N_9668);
or UO_650 (O_650,N_9326,N_9372);
nor UO_651 (O_651,N_9350,N_9153);
nand UO_652 (O_652,N_9298,N_9930);
nand UO_653 (O_653,N_9413,N_9202);
nor UO_654 (O_654,N_9803,N_9493);
and UO_655 (O_655,N_9591,N_9586);
nor UO_656 (O_656,N_9971,N_9996);
and UO_657 (O_657,N_9645,N_9044);
nor UO_658 (O_658,N_9270,N_9399);
nand UO_659 (O_659,N_9705,N_9610);
or UO_660 (O_660,N_9281,N_9613);
nand UO_661 (O_661,N_9929,N_9047);
nor UO_662 (O_662,N_9360,N_9404);
and UO_663 (O_663,N_9128,N_9964);
nand UO_664 (O_664,N_9505,N_9863);
or UO_665 (O_665,N_9277,N_9360);
nand UO_666 (O_666,N_9261,N_9325);
or UO_667 (O_667,N_9751,N_9130);
or UO_668 (O_668,N_9317,N_9148);
and UO_669 (O_669,N_9768,N_9485);
or UO_670 (O_670,N_9303,N_9112);
or UO_671 (O_671,N_9509,N_9314);
nand UO_672 (O_672,N_9719,N_9853);
or UO_673 (O_673,N_9908,N_9470);
or UO_674 (O_674,N_9223,N_9827);
nand UO_675 (O_675,N_9669,N_9853);
and UO_676 (O_676,N_9483,N_9833);
and UO_677 (O_677,N_9330,N_9986);
nand UO_678 (O_678,N_9937,N_9807);
nor UO_679 (O_679,N_9800,N_9137);
nor UO_680 (O_680,N_9765,N_9448);
nor UO_681 (O_681,N_9627,N_9604);
and UO_682 (O_682,N_9322,N_9138);
or UO_683 (O_683,N_9946,N_9672);
and UO_684 (O_684,N_9599,N_9555);
nand UO_685 (O_685,N_9630,N_9061);
nand UO_686 (O_686,N_9984,N_9363);
xnor UO_687 (O_687,N_9905,N_9507);
nor UO_688 (O_688,N_9391,N_9663);
nand UO_689 (O_689,N_9752,N_9616);
and UO_690 (O_690,N_9729,N_9082);
and UO_691 (O_691,N_9781,N_9679);
nor UO_692 (O_692,N_9085,N_9880);
and UO_693 (O_693,N_9036,N_9516);
nand UO_694 (O_694,N_9667,N_9024);
nand UO_695 (O_695,N_9186,N_9472);
nand UO_696 (O_696,N_9794,N_9443);
nand UO_697 (O_697,N_9506,N_9801);
nor UO_698 (O_698,N_9103,N_9790);
or UO_699 (O_699,N_9495,N_9727);
or UO_700 (O_700,N_9545,N_9678);
nand UO_701 (O_701,N_9519,N_9541);
nand UO_702 (O_702,N_9978,N_9647);
or UO_703 (O_703,N_9824,N_9325);
or UO_704 (O_704,N_9284,N_9367);
nand UO_705 (O_705,N_9390,N_9154);
nor UO_706 (O_706,N_9376,N_9106);
nand UO_707 (O_707,N_9608,N_9991);
nand UO_708 (O_708,N_9789,N_9168);
or UO_709 (O_709,N_9318,N_9520);
xnor UO_710 (O_710,N_9050,N_9546);
nand UO_711 (O_711,N_9191,N_9347);
or UO_712 (O_712,N_9091,N_9828);
and UO_713 (O_713,N_9082,N_9039);
nand UO_714 (O_714,N_9355,N_9086);
and UO_715 (O_715,N_9077,N_9375);
and UO_716 (O_716,N_9286,N_9076);
or UO_717 (O_717,N_9767,N_9935);
or UO_718 (O_718,N_9106,N_9313);
nand UO_719 (O_719,N_9579,N_9349);
nor UO_720 (O_720,N_9106,N_9280);
nor UO_721 (O_721,N_9994,N_9082);
nand UO_722 (O_722,N_9894,N_9838);
nor UO_723 (O_723,N_9123,N_9259);
or UO_724 (O_724,N_9405,N_9444);
and UO_725 (O_725,N_9482,N_9774);
nand UO_726 (O_726,N_9496,N_9338);
or UO_727 (O_727,N_9537,N_9852);
nor UO_728 (O_728,N_9828,N_9748);
nand UO_729 (O_729,N_9288,N_9891);
nor UO_730 (O_730,N_9478,N_9933);
nand UO_731 (O_731,N_9120,N_9521);
nand UO_732 (O_732,N_9583,N_9069);
or UO_733 (O_733,N_9958,N_9399);
nand UO_734 (O_734,N_9591,N_9566);
nand UO_735 (O_735,N_9070,N_9188);
nand UO_736 (O_736,N_9772,N_9030);
nand UO_737 (O_737,N_9713,N_9957);
or UO_738 (O_738,N_9031,N_9888);
and UO_739 (O_739,N_9041,N_9312);
and UO_740 (O_740,N_9834,N_9048);
and UO_741 (O_741,N_9154,N_9530);
or UO_742 (O_742,N_9870,N_9973);
nor UO_743 (O_743,N_9232,N_9365);
and UO_744 (O_744,N_9598,N_9752);
nor UO_745 (O_745,N_9775,N_9306);
or UO_746 (O_746,N_9339,N_9804);
and UO_747 (O_747,N_9912,N_9663);
nand UO_748 (O_748,N_9431,N_9700);
nor UO_749 (O_749,N_9778,N_9697);
nand UO_750 (O_750,N_9680,N_9493);
and UO_751 (O_751,N_9271,N_9045);
or UO_752 (O_752,N_9087,N_9071);
nor UO_753 (O_753,N_9312,N_9648);
or UO_754 (O_754,N_9718,N_9926);
or UO_755 (O_755,N_9764,N_9668);
and UO_756 (O_756,N_9318,N_9837);
or UO_757 (O_757,N_9768,N_9418);
or UO_758 (O_758,N_9058,N_9288);
nand UO_759 (O_759,N_9712,N_9480);
nand UO_760 (O_760,N_9117,N_9453);
nor UO_761 (O_761,N_9626,N_9539);
nor UO_762 (O_762,N_9122,N_9029);
nor UO_763 (O_763,N_9869,N_9029);
nor UO_764 (O_764,N_9052,N_9834);
nand UO_765 (O_765,N_9530,N_9495);
nand UO_766 (O_766,N_9335,N_9128);
nor UO_767 (O_767,N_9190,N_9215);
nor UO_768 (O_768,N_9609,N_9197);
or UO_769 (O_769,N_9530,N_9248);
or UO_770 (O_770,N_9142,N_9788);
nor UO_771 (O_771,N_9248,N_9061);
or UO_772 (O_772,N_9644,N_9605);
nor UO_773 (O_773,N_9121,N_9250);
nand UO_774 (O_774,N_9563,N_9136);
nand UO_775 (O_775,N_9458,N_9335);
nand UO_776 (O_776,N_9279,N_9583);
nor UO_777 (O_777,N_9666,N_9902);
or UO_778 (O_778,N_9873,N_9023);
or UO_779 (O_779,N_9611,N_9637);
nand UO_780 (O_780,N_9947,N_9229);
and UO_781 (O_781,N_9555,N_9335);
nor UO_782 (O_782,N_9100,N_9586);
nor UO_783 (O_783,N_9377,N_9560);
nor UO_784 (O_784,N_9403,N_9520);
and UO_785 (O_785,N_9004,N_9155);
nor UO_786 (O_786,N_9419,N_9696);
and UO_787 (O_787,N_9499,N_9804);
nand UO_788 (O_788,N_9283,N_9503);
or UO_789 (O_789,N_9532,N_9927);
nor UO_790 (O_790,N_9506,N_9534);
or UO_791 (O_791,N_9451,N_9417);
nand UO_792 (O_792,N_9826,N_9682);
or UO_793 (O_793,N_9675,N_9611);
and UO_794 (O_794,N_9652,N_9566);
and UO_795 (O_795,N_9288,N_9813);
or UO_796 (O_796,N_9592,N_9266);
nand UO_797 (O_797,N_9612,N_9925);
or UO_798 (O_798,N_9131,N_9226);
nor UO_799 (O_799,N_9098,N_9973);
nand UO_800 (O_800,N_9911,N_9640);
nor UO_801 (O_801,N_9284,N_9132);
or UO_802 (O_802,N_9111,N_9883);
nand UO_803 (O_803,N_9069,N_9257);
nor UO_804 (O_804,N_9280,N_9683);
nor UO_805 (O_805,N_9886,N_9975);
nor UO_806 (O_806,N_9921,N_9205);
or UO_807 (O_807,N_9753,N_9240);
nor UO_808 (O_808,N_9226,N_9172);
nand UO_809 (O_809,N_9867,N_9363);
nor UO_810 (O_810,N_9939,N_9523);
nand UO_811 (O_811,N_9119,N_9305);
nand UO_812 (O_812,N_9234,N_9834);
nor UO_813 (O_813,N_9950,N_9202);
or UO_814 (O_814,N_9771,N_9367);
nand UO_815 (O_815,N_9562,N_9281);
or UO_816 (O_816,N_9041,N_9403);
nand UO_817 (O_817,N_9964,N_9458);
and UO_818 (O_818,N_9792,N_9076);
nand UO_819 (O_819,N_9578,N_9935);
nand UO_820 (O_820,N_9430,N_9189);
nand UO_821 (O_821,N_9696,N_9773);
and UO_822 (O_822,N_9455,N_9058);
nor UO_823 (O_823,N_9853,N_9017);
nand UO_824 (O_824,N_9919,N_9356);
and UO_825 (O_825,N_9394,N_9989);
nor UO_826 (O_826,N_9613,N_9245);
nand UO_827 (O_827,N_9122,N_9857);
nand UO_828 (O_828,N_9816,N_9668);
nor UO_829 (O_829,N_9092,N_9240);
nor UO_830 (O_830,N_9949,N_9279);
nand UO_831 (O_831,N_9138,N_9337);
nand UO_832 (O_832,N_9819,N_9037);
or UO_833 (O_833,N_9567,N_9167);
and UO_834 (O_834,N_9450,N_9651);
nor UO_835 (O_835,N_9032,N_9605);
or UO_836 (O_836,N_9381,N_9166);
or UO_837 (O_837,N_9015,N_9773);
or UO_838 (O_838,N_9845,N_9470);
or UO_839 (O_839,N_9601,N_9055);
or UO_840 (O_840,N_9183,N_9859);
and UO_841 (O_841,N_9670,N_9631);
or UO_842 (O_842,N_9780,N_9549);
and UO_843 (O_843,N_9271,N_9193);
or UO_844 (O_844,N_9125,N_9961);
nand UO_845 (O_845,N_9640,N_9978);
and UO_846 (O_846,N_9460,N_9718);
nor UO_847 (O_847,N_9101,N_9841);
nor UO_848 (O_848,N_9551,N_9339);
nand UO_849 (O_849,N_9675,N_9024);
or UO_850 (O_850,N_9830,N_9296);
and UO_851 (O_851,N_9083,N_9125);
nor UO_852 (O_852,N_9887,N_9823);
nand UO_853 (O_853,N_9219,N_9699);
and UO_854 (O_854,N_9982,N_9928);
nand UO_855 (O_855,N_9008,N_9954);
nand UO_856 (O_856,N_9361,N_9814);
and UO_857 (O_857,N_9413,N_9708);
nand UO_858 (O_858,N_9623,N_9696);
nor UO_859 (O_859,N_9000,N_9443);
or UO_860 (O_860,N_9557,N_9712);
nor UO_861 (O_861,N_9552,N_9522);
nand UO_862 (O_862,N_9053,N_9221);
nor UO_863 (O_863,N_9548,N_9983);
and UO_864 (O_864,N_9072,N_9232);
or UO_865 (O_865,N_9356,N_9270);
nand UO_866 (O_866,N_9494,N_9032);
and UO_867 (O_867,N_9020,N_9542);
nand UO_868 (O_868,N_9291,N_9809);
and UO_869 (O_869,N_9438,N_9214);
nand UO_870 (O_870,N_9291,N_9453);
and UO_871 (O_871,N_9409,N_9774);
and UO_872 (O_872,N_9344,N_9193);
and UO_873 (O_873,N_9984,N_9947);
and UO_874 (O_874,N_9089,N_9421);
nor UO_875 (O_875,N_9362,N_9970);
nand UO_876 (O_876,N_9329,N_9351);
and UO_877 (O_877,N_9299,N_9507);
nand UO_878 (O_878,N_9979,N_9750);
nor UO_879 (O_879,N_9697,N_9328);
nor UO_880 (O_880,N_9313,N_9377);
and UO_881 (O_881,N_9700,N_9815);
nand UO_882 (O_882,N_9694,N_9339);
nor UO_883 (O_883,N_9949,N_9381);
and UO_884 (O_884,N_9831,N_9752);
and UO_885 (O_885,N_9205,N_9389);
or UO_886 (O_886,N_9937,N_9375);
or UO_887 (O_887,N_9986,N_9546);
nand UO_888 (O_888,N_9860,N_9757);
or UO_889 (O_889,N_9528,N_9194);
and UO_890 (O_890,N_9607,N_9065);
nor UO_891 (O_891,N_9092,N_9890);
xnor UO_892 (O_892,N_9770,N_9520);
nand UO_893 (O_893,N_9911,N_9885);
nor UO_894 (O_894,N_9220,N_9054);
and UO_895 (O_895,N_9071,N_9056);
and UO_896 (O_896,N_9005,N_9942);
and UO_897 (O_897,N_9235,N_9234);
or UO_898 (O_898,N_9809,N_9915);
and UO_899 (O_899,N_9280,N_9637);
or UO_900 (O_900,N_9286,N_9172);
nor UO_901 (O_901,N_9411,N_9969);
nand UO_902 (O_902,N_9899,N_9179);
or UO_903 (O_903,N_9514,N_9116);
nor UO_904 (O_904,N_9749,N_9405);
and UO_905 (O_905,N_9239,N_9299);
nand UO_906 (O_906,N_9371,N_9593);
and UO_907 (O_907,N_9172,N_9837);
and UO_908 (O_908,N_9583,N_9998);
nor UO_909 (O_909,N_9660,N_9175);
nand UO_910 (O_910,N_9263,N_9091);
or UO_911 (O_911,N_9093,N_9391);
nor UO_912 (O_912,N_9460,N_9299);
nand UO_913 (O_913,N_9333,N_9760);
or UO_914 (O_914,N_9617,N_9926);
nor UO_915 (O_915,N_9004,N_9063);
and UO_916 (O_916,N_9393,N_9062);
nor UO_917 (O_917,N_9440,N_9808);
or UO_918 (O_918,N_9531,N_9116);
or UO_919 (O_919,N_9903,N_9879);
xnor UO_920 (O_920,N_9126,N_9415);
nor UO_921 (O_921,N_9359,N_9118);
nor UO_922 (O_922,N_9460,N_9780);
nand UO_923 (O_923,N_9679,N_9629);
nor UO_924 (O_924,N_9981,N_9331);
nor UO_925 (O_925,N_9860,N_9704);
or UO_926 (O_926,N_9508,N_9028);
nand UO_927 (O_927,N_9619,N_9692);
nor UO_928 (O_928,N_9340,N_9597);
nor UO_929 (O_929,N_9634,N_9731);
nor UO_930 (O_930,N_9977,N_9999);
or UO_931 (O_931,N_9353,N_9607);
and UO_932 (O_932,N_9660,N_9890);
or UO_933 (O_933,N_9277,N_9942);
nor UO_934 (O_934,N_9557,N_9490);
or UO_935 (O_935,N_9208,N_9440);
or UO_936 (O_936,N_9192,N_9087);
or UO_937 (O_937,N_9114,N_9269);
nor UO_938 (O_938,N_9256,N_9230);
and UO_939 (O_939,N_9789,N_9967);
nand UO_940 (O_940,N_9979,N_9969);
or UO_941 (O_941,N_9642,N_9388);
or UO_942 (O_942,N_9527,N_9424);
and UO_943 (O_943,N_9290,N_9568);
and UO_944 (O_944,N_9835,N_9001);
nand UO_945 (O_945,N_9595,N_9279);
nand UO_946 (O_946,N_9545,N_9533);
and UO_947 (O_947,N_9847,N_9933);
nand UO_948 (O_948,N_9105,N_9666);
or UO_949 (O_949,N_9819,N_9358);
and UO_950 (O_950,N_9796,N_9890);
nand UO_951 (O_951,N_9843,N_9946);
nand UO_952 (O_952,N_9102,N_9950);
or UO_953 (O_953,N_9336,N_9147);
nor UO_954 (O_954,N_9069,N_9532);
or UO_955 (O_955,N_9576,N_9063);
or UO_956 (O_956,N_9674,N_9888);
nor UO_957 (O_957,N_9939,N_9548);
nor UO_958 (O_958,N_9087,N_9358);
or UO_959 (O_959,N_9884,N_9551);
nor UO_960 (O_960,N_9850,N_9240);
nand UO_961 (O_961,N_9586,N_9122);
xor UO_962 (O_962,N_9929,N_9851);
nor UO_963 (O_963,N_9063,N_9912);
nor UO_964 (O_964,N_9681,N_9966);
nor UO_965 (O_965,N_9787,N_9553);
or UO_966 (O_966,N_9928,N_9612);
nand UO_967 (O_967,N_9136,N_9207);
or UO_968 (O_968,N_9429,N_9340);
and UO_969 (O_969,N_9656,N_9775);
nor UO_970 (O_970,N_9773,N_9338);
and UO_971 (O_971,N_9750,N_9182);
nor UO_972 (O_972,N_9543,N_9291);
and UO_973 (O_973,N_9136,N_9502);
nor UO_974 (O_974,N_9050,N_9854);
and UO_975 (O_975,N_9866,N_9589);
nand UO_976 (O_976,N_9475,N_9711);
or UO_977 (O_977,N_9254,N_9821);
nand UO_978 (O_978,N_9610,N_9117);
nand UO_979 (O_979,N_9760,N_9077);
and UO_980 (O_980,N_9852,N_9330);
nand UO_981 (O_981,N_9279,N_9791);
or UO_982 (O_982,N_9512,N_9881);
nand UO_983 (O_983,N_9077,N_9952);
nand UO_984 (O_984,N_9357,N_9390);
or UO_985 (O_985,N_9408,N_9686);
or UO_986 (O_986,N_9468,N_9721);
nand UO_987 (O_987,N_9712,N_9309);
nor UO_988 (O_988,N_9266,N_9166);
or UO_989 (O_989,N_9376,N_9240);
nor UO_990 (O_990,N_9709,N_9079);
and UO_991 (O_991,N_9886,N_9400);
nand UO_992 (O_992,N_9327,N_9422);
or UO_993 (O_993,N_9772,N_9745);
and UO_994 (O_994,N_9926,N_9138);
nand UO_995 (O_995,N_9910,N_9462);
and UO_996 (O_996,N_9542,N_9308);
nor UO_997 (O_997,N_9566,N_9241);
and UO_998 (O_998,N_9836,N_9222);
nor UO_999 (O_999,N_9971,N_9427);
and UO_1000 (O_1000,N_9998,N_9483);
nor UO_1001 (O_1001,N_9667,N_9097);
and UO_1002 (O_1002,N_9390,N_9526);
nor UO_1003 (O_1003,N_9837,N_9422);
or UO_1004 (O_1004,N_9142,N_9561);
and UO_1005 (O_1005,N_9164,N_9815);
nor UO_1006 (O_1006,N_9315,N_9084);
nor UO_1007 (O_1007,N_9296,N_9072);
nor UO_1008 (O_1008,N_9820,N_9851);
or UO_1009 (O_1009,N_9337,N_9753);
nor UO_1010 (O_1010,N_9878,N_9989);
nand UO_1011 (O_1011,N_9214,N_9607);
and UO_1012 (O_1012,N_9918,N_9953);
and UO_1013 (O_1013,N_9347,N_9374);
or UO_1014 (O_1014,N_9913,N_9373);
nor UO_1015 (O_1015,N_9995,N_9736);
xnor UO_1016 (O_1016,N_9818,N_9023);
nor UO_1017 (O_1017,N_9426,N_9983);
and UO_1018 (O_1018,N_9131,N_9069);
nor UO_1019 (O_1019,N_9694,N_9911);
or UO_1020 (O_1020,N_9553,N_9483);
nand UO_1021 (O_1021,N_9916,N_9440);
nor UO_1022 (O_1022,N_9410,N_9394);
nand UO_1023 (O_1023,N_9480,N_9542);
nor UO_1024 (O_1024,N_9190,N_9467);
nand UO_1025 (O_1025,N_9717,N_9959);
and UO_1026 (O_1026,N_9703,N_9235);
nand UO_1027 (O_1027,N_9038,N_9815);
nand UO_1028 (O_1028,N_9278,N_9149);
nor UO_1029 (O_1029,N_9773,N_9988);
or UO_1030 (O_1030,N_9257,N_9849);
and UO_1031 (O_1031,N_9997,N_9479);
and UO_1032 (O_1032,N_9922,N_9295);
and UO_1033 (O_1033,N_9105,N_9971);
nor UO_1034 (O_1034,N_9678,N_9109);
or UO_1035 (O_1035,N_9148,N_9491);
nor UO_1036 (O_1036,N_9427,N_9925);
and UO_1037 (O_1037,N_9186,N_9428);
nand UO_1038 (O_1038,N_9684,N_9832);
and UO_1039 (O_1039,N_9395,N_9458);
nor UO_1040 (O_1040,N_9156,N_9047);
and UO_1041 (O_1041,N_9053,N_9856);
and UO_1042 (O_1042,N_9274,N_9447);
nand UO_1043 (O_1043,N_9561,N_9414);
and UO_1044 (O_1044,N_9823,N_9734);
and UO_1045 (O_1045,N_9333,N_9038);
or UO_1046 (O_1046,N_9873,N_9806);
or UO_1047 (O_1047,N_9672,N_9434);
and UO_1048 (O_1048,N_9759,N_9933);
nand UO_1049 (O_1049,N_9381,N_9243);
nand UO_1050 (O_1050,N_9827,N_9195);
nand UO_1051 (O_1051,N_9190,N_9113);
nor UO_1052 (O_1052,N_9966,N_9660);
or UO_1053 (O_1053,N_9578,N_9336);
nor UO_1054 (O_1054,N_9502,N_9405);
nand UO_1055 (O_1055,N_9524,N_9831);
nand UO_1056 (O_1056,N_9458,N_9666);
or UO_1057 (O_1057,N_9489,N_9262);
nand UO_1058 (O_1058,N_9524,N_9392);
nor UO_1059 (O_1059,N_9273,N_9584);
nand UO_1060 (O_1060,N_9582,N_9671);
and UO_1061 (O_1061,N_9901,N_9642);
or UO_1062 (O_1062,N_9721,N_9978);
or UO_1063 (O_1063,N_9269,N_9427);
or UO_1064 (O_1064,N_9446,N_9507);
or UO_1065 (O_1065,N_9189,N_9827);
nor UO_1066 (O_1066,N_9317,N_9954);
or UO_1067 (O_1067,N_9716,N_9038);
nor UO_1068 (O_1068,N_9766,N_9384);
or UO_1069 (O_1069,N_9284,N_9938);
nor UO_1070 (O_1070,N_9140,N_9042);
nand UO_1071 (O_1071,N_9571,N_9585);
or UO_1072 (O_1072,N_9741,N_9452);
nand UO_1073 (O_1073,N_9508,N_9826);
and UO_1074 (O_1074,N_9977,N_9791);
or UO_1075 (O_1075,N_9424,N_9163);
and UO_1076 (O_1076,N_9558,N_9375);
nor UO_1077 (O_1077,N_9599,N_9355);
or UO_1078 (O_1078,N_9952,N_9318);
or UO_1079 (O_1079,N_9818,N_9688);
and UO_1080 (O_1080,N_9749,N_9913);
and UO_1081 (O_1081,N_9513,N_9992);
nor UO_1082 (O_1082,N_9527,N_9941);
or UO_1083 (O_1083,N_9719,N_9976);
nand UO_1084 (O_1084,N_9898,N_9131);
nand UO_1085 (O_1085,N_9646,N_9084);
nor UO_1086 (O_1086,N_9291,N_9128);
and UO_1087 (O_1087,N_9728,N_9247);
and UO_1088 (O_1088,N_9513,N_9152);
or UO_1089 (O_1089,N_9904,N_9242);
nand UO_1090 (O_1090,N_9276,N_9663);
or UO_1091 (O_1091,N_9537,N_9260);
nor UO_1092 (O_1092,N_9528,N_9493);
or UO_1093 (O_1093,N_9078,N_9513);
nor UO_1094 (O_1094,N_9467,N_9217);
and UO_1095 (O_1095,N_9972,N_9551);
and UO_1096 (O_1096,N_9109,N_9568);
nand UO_1097 (O_1097,N_9935,N_9553);
and UO_1098 (O_1098,N_9217,N_9052);
nand UO_1099 (O_1099,N_9835,N_9892);
and UO_1100 (O_1100,N_9693,N_9314);
or UO_1101 (O_1101,N_9514,N_9186);
nand UO_1102 (O_1102,N_9724,N_9013);
nand UO_1103 (O_1103,N_9769,N_9921);
and UO_1104 (O_1104,N_9426,N_9077);
nor UO_1105 (O_1105,N_9612,N_9207);
nand UO_1106 (O_1106,N_9772,N_9831);
nor UO_1107 (O_1107,N_9280,N_9484);
nand UO_1108 (O_1108,N_9131,N_9335);
and UO_1109 (O_1109,N_9175,N_9027);
or UO_1110 (O_1110,N_9097,N_9112);
and UO_1111 (O_1111,N_9074,N_9221);
xnor UO_1112 (O_1112,N_9821,N_9786);
or UO_1113 (O_1113,N_9463,N_9117);
nor UO_1114 (O_1114,N_9412,N_9229);
or UO_1115 (O_1115,N_9253,N_9981);
nand UO_1116 (O_1116,N_9004,N_9228);
and UO_1117 (O_1117,N_9067,N_9075);
nor UO_1118 (O_1118,N_9764,N_9940);
nand UO_1119 (O_1119,N_9808,N_9738);
nor UO_1120 (O_1120,N_9121,N_9602);
nor UO_1121 (O_1121,N_9892,N_9173);
and UO_1122 (O_1122,N_9398,N_9884);
nor UO_1123 (O_1123,N_9307,N_9845);
nand UO_1124 (O_1124,N_9874,N_9357);
nor UO_1125 (O_1125,N_9926,N_9018);
and UO_1126 (O_1126,N_9035,N_9964);
nor UO_1127 (O_1127,N_9818,N_9404);
nor UO_1128 (O_1128,N_9795,N_9066);
or UO_1129 (O_1129,N_9804,N_9513);
nand UO_1130 (O_1130,N_9198,N_9340);
nor UO_1131 (O_1131,N_9898,N_9691);
and UO_1132 (O_1132,N_9397,N_9897);
nor UO_1133 (O_1133,N_9397,N_9494);
nor UO_1134 (O_1134,N_9942,N_9885);
nand UO_1135 (O_1135,N_9503,N_9474);
nand UO_1136 (O_1136,N_9718,N_9028);
and UO_1137 (O_1137,N_9316,N_9947);
or UO_1138 (O_1138,N_9373,N_9225);
and UO_1139 (O_1139,N_9572,N_9102);
nand UO_1140 (O_1140,N_9729,N_9422);
and UO_1141 (O_1141,N_9986,N_9967);
or UO_1142 (O_1142,N_9743,N_9300);
and UO_1143 (O_1143,N_9256,N_9799);
or UO_1144 (O_1144,N_9778,N_9192);
or UO_1145 (O_1145,N_9526,N_9914);
and UO_1146 (O_1146,N_9817,N_9292);
nor UO_1147 (O_1147,N_9218,N_9933);
nand UO_1148 (O_1148,N_9913,N_9607);
or UO_1149 (O_1149,N_9323,N_9800);
nand UO_1150 (O_1150,N_9089,N_9177);
or UO_1151 (O_1151,N_9789,N_9002);
nor UO_1152 (O_1152,N_9329,N_9704);
nand UO_1153 (O_1153,N_9917,N_9670);
nor UO_1154 (O_1154,N_9031,N_9159);
or UO_1155 (O_1155,N_9766,N_9777);
or UO_1156 (O_1156,N_9682,N_9074);
and UO_1157 (O_1157,N_9234,N_9352);
nor UO_1158 (O_1158,N_9178,N_9371);
nand UO_1159 (O_1159,N_9885,N_9337);
and UO_1160 (O_1160,N_9164,N_9138);
or UO_1161 (O_1161,N_9435,N_9449);
nand UO_1162 (O_1162,N_9508,N_9924);
or UO_1163 (O_1163,N_9025,N_9259);
or UO_1164 (O_1164,N_9385,N_9720);
nand UO_1165 (O_1165,N_9997,N_9515);
nor UO_1166 (O_1166,N_9909,N_9539);
nand UO_1167 (O_1167,N_9403,N_9959);
nor UO_1168 (O_1168,N_9734,N_9492);
and UO_1169 (O_1169,N_9798,N_9191);
and UO_1170 (O_1170,N_9694,N_9671);
nor UO_1171 (O_1171,N_9190,N_9816);
nand UO_1172 (O_1172,N_9416,N_9982);
or UO_1173 (O_1173,N_9789,N_9344);
or UO_1174 (O_1174,N_9417,N_9426);
nand UO_1175 (O_1175,N_9754,N_9652);
or UO_1176 (O_1176,N_9618,N_9073);
nand UO_1177 (O_1177,N_9789,N_9454);
nor UO_1178 (O_1178,N_9052,N_9685);
and UO_1179 (O_1179,N_9348,N_9370);
and UO_1180 (O_1180,N_9429,N_9108);
nor UO_1181 (O_1181,N_9962,N_9997);
nor UO_1182 (O_1182,N_9756,N_9447);
nand UO_1183 (O_1183,N_9149,N_9212);
nand UO_1184 (O_1184,N_9255,N_9895);
nand UO_1185 (O_1185,N_9624,N_9710);
nor UO_1186 (O_1186,N_9513,N_9493);
and UO_1187 (O_1187,N_9195,N_9881);
or UO_1188 (O_1188,N_9646,N_9148);
or UO_1189 (O_1189,N_9449,N_9511);
nor UO_1190 (O_1190,N_9227,N_9173);
and UO_1191 (O_1191,N_9517,N_9379);
nand UO_1192 (O_1192,N_9923,N_9569);
and UO_1193 (O_1193,N_9284,N_9757);
nor UO_1194 (O_1194,N_9415,N_9555);
or UO_1195 (O_1195,N_9036,N_9753);
nand UO_1196 (O_1196,N_9725,N_9086);
nor UO_1197 (O_1197,N_9561,N_9295);
and UO_1198 (O_1198,N_9894,N_9282);
nor UO_1199 (O_1199,N_9827,N_9067);
nand UO_1200 (O_1200,N_9082,N_9058);
nand UO_1201 (O_1201,N_9682,N_9697);
or UO_1202 (O_1202,N_9058,N_9547);
nor UO_1203 (O_1203,N_9921,N_9882);
nand UO_1204 (O_1204,N_9653,N_9442);
and UO_1205 (O_1205,N_9166,N_9071);
and UO_1206 (O_1206,N_9703,N_9931);
nand UO_1207 (O_1207,N_9055,N_9558);
and UO_1208 (O_1208,N_9847,N_9259);
nand UO_1209 (O_1209,N_9478,N_9660);
nor UO_1210 (O_1210,N_9974,N_9158);
nand UO_1211 (O_1211,N_9643,N_9392);
nor UO_1212 (O_1212,N_9352,N_9607);
nand UO_1213 (O_1213,N_9748,N_9343);
nand UO_1214 (O_1214,N_9717,N_9155);
and UO_1215 (O_1215,N_9015,N_9468);
nor UO_1216 (O_1216,N_9602,N_9405);
nor UO_1217 (O_1217,N_9514,N_9746);
or UO_1218 (O_1218,N_9975,N_9658);
and UO_1219 (O_1219,N_9514,N_9282);
and UO_1220 (O_1220,N_9347,N_9827);
or UO_1221 (O_1221,N_9316,N_9990);
or UO_1222 (O_1222,N_9538,N_9342);
and UO_1223 (O_1223,N_9396,N_9958);
nand UO_1224 (O_1224,N_9794,N_9692);
nand UO_1225 (O_1225,N_9817,N_9940);
or UO_1226 (O_1226,N_9741,N_9385);
nand UO_1227 (O_1227,N_9806,N_9534);
nor UO_1228 (O_1228,N_9166,N_9041);
or UO_1229 (O_1229,N_9387,N_9735);
nand UO_1230 (O_1230,N_9970,N_9100);
or UO_1231 (O_1231,N_9933,N_9786);
and UO_1232 (O_1232,N_9476,N_9380);
nand UO_1233 (O_1233,N_9236,N_9183);
and UO_1234 (O_1234,N_9430,N_9013);
and UO_1235 (O_1235,N_9746,N_9181);
nor UO_1236 (O_1236,N_9404,N_9132);
and UO_1237 (O_1237,N_9426,N_9345);
and UO_1238 (O_1238,N_9079,N_9235);
and UO_1239 (O_1239,N_9890,N_9920);
nand UO_1240 (O_1240,N_9441,N_9622);
and UO_1241 (O_1241,N_9356,N_9318);
nand UO_1242 (O_1242,N_9027,N_9072);
and UO_1243 (O_1243,N_9007,N_9202);
nand UO_1244 (O_1244,N_9108,N_9600);
nor UO_1245 (O_1245,N_9610,N_9633);
nand UO_1246 (O_1246,N_9945,N_9757);
nand UO_1247 (O_1247,N_9883,N_9482);
and UO_1248 (O_1248,N_9754,N_9086);
nor UO_1249 (O_1249,N_9630,N_9346);
and UO_1250 (O_1250,N_9643,N_9798);
or UO_1251 (O_1251,N_9200,N_9616);
nand UO_1252 (O_1252,N_9161,N_9342);
nor UO_1253 (O_1253,N_9868,N_9754);
nor UO_1254 (O_1254,N_9774,N_9615);
or UO_1255 (O_1255,N_9461,N_9296);
nor UO_1256 (O_1256,N_9193,N_9501);
nor UO_1257 (O_1257,N_9086,N_9173);
or UO_1258 (O_1258,N_9629,N_9281);
and UO_1259 (O_1259,N_9443,N_9945);
or UO_1260 (O_1260,N_9265,N_9579);
nor UO_1261 (O_1261,N_9039,N_9028);
and UO_1262 (O_1262,N_9121,N_9520);
xor UO_1263 (O_1263,N_9816,N_9565);
nand UO_1264 (O_1264,N_9712,N_9903);
and UO_1265 (O_1265,N_9777,N_9528);
or UO_1266 (O_1266,N_9496,N_9311);
nor UO_1267 (O_1267,N_9969,N_9903);
and UO_1268 (O_1268,N_9266,N_9612);
nor UO_1269 (O_1269,N_9912,N_9098);
nand UO_1270 (O_1270,N_9995,N_9016);
nor UO_1271 (O_1271,N_9061,N_9566);
nand UO_1272 (O_1272,N_9561,N_9297);
and UO_1273 (O_1273,N_9118,N_9146);
nor UO_1274 (O_1274,N_9535,N_9255);
or UO_1275 (O_1275,N_9665,N_9729);
nand UO_1276 (O_1276,N_9956,N_9096);
nand UO_1277 (O_1277,N_9191,N_9757);
or UO_1278 (O_1278,N_9933,N_9049);
nand UO_1279 (O_1279,N_9178,N_9787);
or UO_1280 (O_1280,N_9464,N_9275);
and UO_1281 (O_1281,N_9882,N_9623);
nand UO_1282 (O_1282,N_9565,N_9420);
and UO_1283 (O_1283,N_9540,N_9606);
nor UO_1284 (O_1284,N_9573,N_9378);
nand UO_1285 (O_1285,N_9680,N_9723);
nand UO_1286 (O_1286,N_9613,N_9913);
and UO_1287 (O_1287,N_9236,N_9476);
and UO_1288 (O_1288,N_9451,N_9795);
and UO_1289 (O_1289,N_9132,N_9019);
nor UO_1290 (O_1290,N_9662,N_9896);
and UO_1291 (O_1291,N_9437,N_9499);
and UO_1292 (O_1292,N_9261,N_9625);
and UO_1293 (O_1293,N_9711,N_9646);
or UO_1294 (O_1294,N_9672,N_9104);
nand UO_1295 (O_1295,N_9786,N_9833);
nand UO_1296 (O_1296,N_9457,N_9492);
nor UO_1297 (O_1297,N_9261,N_9513);
or UO_1298 (O_1298,N_9000,N_9337);
or UO_1299 (O_1299,N_9048,N_9452);
nand UO_1300 (O_1300,N_9669,N_9462);
nand UO_1301 (O_1301,N_9543,N_9527);
nand UO_1302 (O_1302,N_9552,N_9379);
nor UO_1303 (O_1303,N_9339,N_9825);
and UO_1304 (O_1304,N_9287,N_9562);
or UO_1305 (O_1305,N_9625,N_9080);
or UO_1306 (O_1306,N_9629,N_9088);
and UO_1307 (O_1307,N_9505,N_9407);
nor UO_1308 (O_1308,N_9730,N_9688);
and UO_1309 (O_1309,N_9477,N_9709);
nand UO_1310 (O_1310,N_9861,N_9880);
nor UO_1311 (O_1311,N_9629,N_9814);
or UO_1312 (O_1312,N_9345,N_9665);
and UO_1313 (O_1313,N_9028,N_9531);
nor UO_1314 (O_1314,N_9733,N_9171);
nor UO_1315 (O_1315,N_9332,N_9313);
and UO_1316 (O_1316,N_9905,N_9351);
nand UO_1317 (O_1317,N_9936,N_9084);
nand UO_1318 (O_1318,N_9404,N_9456);
nor UO_1319 (O_1319,N_9441,N_9847);
nand UO_1320 (O_1320,N_9188,N_9141);
and UO_1321 (O_1321,N_9910,N_9908);
nor UO_1322 (O_1322,N_9026,N_9207);
or UO_1323 (O_1323,N_9327,N_9429);
nor UO_1324 (O_1324,N_9316,N_9574);
nor UO_1325 (O_1325,N_9618,N_9683);
nand UO_1326 (O_1326,N_9417,N_9043);
nor UO_1327 (O_1327,N_9644,N_9898);
or UO_1328 (O_1328,N_9533,N_9205);
nand UO_1329 (O_1329,N_9410,N_9814);
nor UO_1330 (O_1330,N_9394,N_9191);
and UO_1331 (O_1331,N_9541,N_9272);
and UO_1332 (O_1332,N_9301,N_9716);
nor UO_1333 (O_1333,N_9667,N_9640);
and UO_1334 (O_1334,N_9882,N_9643);
or UO_1335 (O_1335,N_9066,N_9380);
nand UO_1336 (O_1336,N_9456,N_9758);
nand UO_1337 (O_1337,N_9400,N_9264);
nand UO_1338 (O_1338,N_9441,N_9249);
nand UO_1339 (O_1339,N_9689,N_9125);
nand UO_1340 (O_1340,N_9950,N_9644);
nor UO_1341 (O_1341,N_9711,N_9854);
nand UO_1342 (O_1342,N_9678,N_9480);
and UO_1343 (O_1343,N_9511,N_9143);
and UO_1344 (O_1344,N_9143,N_9491);
and UO_1345 (O_1345,N_9132,N_9272);
nand UO_1346 (O_1346,N_9666,N_9359);
nor UO_1347 (O_1347,N_9405,N_9667);
nor UO_1348 (O_1348,N_9935,N_9918);
nor UO_1349 (O_1349,N_9048,N_9252);
and UO_1350 (O_1350,N_9485,N_9392);
nand UO_1351 (O_1351,N_9022,N_9777);
nand UO_1352 (O_1352,N_9478,N_9159);
or UO_1353 (O_1353,N_9757,N_9109);
nor UO_1354 (O_1354,N_9334,N_9515);
nor UO_1355 (O_1355,N_9099,N_9520);
nand UO_1356 (O_1356,N_9307,N_9676);
and UO_1357 (O_1357,N_9517,N_9221);
and UO_1358 (O_1358,N_9437,N_9388);
and UO_1359 (O_1359,N_9466,N_9224);
and UO_1360 (O_1360,N_9707,N_9902);
nand UO_1361 (O_1361,N_9302,N_9029);
or UO_1362 (O_1362,N_9764,N_9325);
xnor UO_1363 (O_1363,N_9683,N_9436);
nor UO_1364 (O_1364,N_9403,N_9785);
or UO_1365 (O_1365,N_9818,N_9168);
or UO_1366 (O_1366,N_9965,N_9366);
and UO_1367 (O_1367,N_9633,N_9996);
and UO_1368 (O_1368,N_9310,N_9174);
nor UO_1369 (O_1369,N_9733,N_9979);
and UO_1370 (O_1370,N_9132,N_9828);
or UO_1371 (O_1371,N_9275,N_9240);
nor UO_1372 (O_1372,N_9918,N_9655);
or UO_1373 (O_1373,N_9327,N_9744);
nand UO_1374 (O_1374,N_9039,N_9953);
or UO_1375 (O_1375,N_9888,N_9342);
and UO_1376 (O_1376,N_9423,N_9949);
nand UO_1377 (O_1377,N_9045,N_9704);
and UO_1378 (O_1378,N_9323,N_9082);
or UO_1379 (O_1379,N_9732,N_9227);
nand UO_1380 (O_1380,N_9009,N_9125);
and UO_1381 (O_1381,N_9561,N_9622);
or UO_1382 (O_1382,N_9090,N_9102);
nand UO_1383 (O_1383,N_9904,N_9279);
nor UO_1384 (O_1384,N_9399,N_9103);
or UO_1385 (O_1385,N_9446,N_9175);
nand UO_1386 (O_1386,N_9596,N_9541);
or UO_1387 (O_1387,N_9785,N_9033);
and UO_1388 (O_1388,N_9351,N_9450);
nor UO_1389 (O_1389,N_9444,N_9223);
nand UO_1390 (O_1390,N_9432,N_9070);
nor UO_1391 (O_1391,N_9415,N_9431);
nand UO_1392 (O_1392,N_9812,N_9879);
or UO_1393 (O_1393,N_9447,N_9153);
and UO_1394 (O_1394,N_9385,N_9009);
nand UO_1395 (O_1395,N_9954,N_9574);
nand UO_1396 (O_1396,N_9988,N_9149);
and UO_1397 (O_1397,N_9069,N_9810);
and UO_1398 (O_1398,N_9955,N_9738);
and UO_1399 (O_1399,N_9609,N_9621);
nand UO_1400 (O_1400,N_9868,N_9002);
and UO_1401 (O_1401,N_9654,N_9382);
and UO_1402 (O_1402,N_9018,N_9011);
nor UO_1403 (O_1403,N_9717,N_9098);
and UO_1404 (O_1404,N_9690,N_9514);
or UO_1405 (O_1405,N_9145,N_9091);
nor UO_1406 (O_1406,N_9198,N_9150);
nor UO_1407 (O_1407,N_9749,N_9475);
nor UO_1408 (O_1408,N_9966,N_9249);
nand UO_1409 (O_1409,N_9546,N_9282);
or UO_1410 (O_1410,N_9116,N_9708);
or UO_1411 (O_1411,N_9294,N_9320);
nor UO_1412 (O_1412,N_9241,N_9768);
and UO_1413 (O_1413,N_9609,N_9324);
nand UO_1414 (O_1414,N_9187,N_9675);
or UO_1415 (O_1415,N_9607,N_9185);
nor UO_1416 (O_1416,N_9571,N_9170);
or UO_1417 (O_1417,N_9739,N_9988);
nor UO_1418 (O_1418,N_9456,N_9839);
and UO_1419 (O_1419,N_9170,N_9794);
or UO_1420 (O_1420,N_9349,N_9247);
nor UO_1421 (O_1421,N_9534,N_9523);
and UO_1422 (O_1422,N_9918,N_9904);
nor UO_1423 (O_1423,N_9366,N_9649);
and UO_1424 (O_1424,N_9342,N_9874);
nand UO_1425 (O_1425,N_9055,N_9467);
nand UO_1426 (O_1426,N_9588,N_9064);
and UO_1427 (O_1427,N_9095,N_9447);
and UO_1428 (O_1428,N_9558,N_9848);
nor UO_1429 (O_1429,N_9707,N_9317);
nand UO_1430 (O_1430,N_9251,N_9861);
nand UO_1431 (O_1431,N_9527,N_9808);
or UO_1432 (O_1432,N_9541,N_9768);
nor UO_1433 (O_1433,N_9807,N_9761);
nor UO_1434 (O_1434,N_9364,N_9551);
nand UO_1435 (O_1435,N_9775,N_9608);
nor UO_1436 (O_1436,N_9190,N_9764);
and UO_1437 (O_1437,N_9233,N_9437);
and UO_1438 (O_1438,N_9929,N_9741);
nand UO_1439 (O_1439,N_9765,N_9940);
nand UO_1440 (O_1440,N_9880,N_9186);
or UO_1441 (O_1441,N_9833,N_9866);
xnor UO_1442 (O_1442,N_9626,N_9030);
nand UO_1443 (O_1443,N_9374,N_9183);
and UO_1444 (O_1444,N_9388,N_9008);
nand UO_1445 (O_1445,N_9502,N_9450);
and UO_1446 (O_1446,N_9080,N_9972);
nand UO_1447 (O_1447,N_9202,N_9752);
or UO_1448 (O_1448,N_9247,N_9578);
nor UO_1449 (O_1449,N_9661,N_9949);
nand UO_1450 (O_1450,N_9956,N_9572);
nand UO_1451 (O_1451,N_9629,N_9030);
nor UO_1452 (O_1452,N_9204,N_9798);
nand UO_1453 (O_1453,N_9852,N_9942);
and UO_1454 (O_1454,N_9982,N_9897);
nand UO_1455 (O_1455,N_9466,N_9292);
nand UO_1456 (O_1456,N_9052,N_9615);
and UO_1457 (O_1457,N_9972,N_9745);
or UO_1458 (O_1458,N_9306,N_9532);
nand UO_1459 (O_1459,N_9810,N_9190);
nand UO_1460 (O_1460,N_9380,N_9534);
nor UO_1461 (O_1461,N_9272,N_9363);
or UO_1462 (O_1462,N_9802,N_9913);
nor UO_1463 (O_1463,N_9440,N_9767);
or UO_1464 (O_1464,N_9541,N_9798);
nor UO_1465 (O_1465,N_9661,N_9556);
and UO_1466 (O_1466,N_9395,N_9287);
nor UO_1467 (O_1467,N_9394,N_9578);
nand UO_1468 (O_1468,N_9108,N_9157);
or UO_1469 (O_1469,N_9308,N_9273);
and UO_1470 (O_1470,N_9569,N_9717);
nor UO_1471 (O_1471,N_9375,N_9178);
and UO_1472 (O_1472,N_9245,N_9699);
and UO_1473 (O_1473,N_9774,N_9404);
or UO_1474 (O_1474,N_9405,N_9514);
or UO_1475 (O_1475,N_9988,N_9456);
nand UO_1476 (O_1476,N_9028,N_9886);
nor UO_1477 (O_1477,N_9355,N_9991);
or UO_1478 (O_1478,N_9446,N_9003);
nor UO_1479 (O_1479,N_9458,N_9055);
or UO_1480 (O_1480,N_9875,N_9511);
nor UO_1481 (O_1481,N_9463,N_9238);
or UO_1482 (O_1482,N_9082,N_9959);
and UO_1483 (O_1483,N_9729,N_9674);
and UO_1484 (O_1484,N_9436,N_9680);
xnor UO_1485 (O_1485,N_9627,N_9069);
nor UO_1486 (O_1486,N_9369,N_9555);
or UO_1487 (O_1487,N_9927,N_9939);
nor UO_1488 (O_1488,N_9422,N_9436);
nand UO_1489 (O_1489,N_9357,N_9981);
and UO_1490 (O_1490,N_9229,N_9221);
nor UO_1491 (O_1491,N_9544,N_9005);
or UO_1492 (O_1492,N_9683,N_9348);
nor UO_1493 (O_1493,N_9341,N_9835);
and UO_1494 (O_1494,N_9962,N_9158);
or UO_1495 (O_1495,N_9822,N_9963);
xor UO_1496 (O_1496,N_9611,N_9103);
or UO_1497 (O_1497,N_9951,N_9310);
nand UO_1498 (O_1498,N_9106,N_9277);
nand UO_1499 (O_1499,N_9038,N_9348);
endmodule