module basic_500_3000_500_50_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_90,In_147);
and U1 (N_1,In_347,In_283);
and U2 (N_2,In_414,In_493);
and U3 (N_3,In_419,In_161);
nor U4 (N_4,In_441,In_464);
nand U5 (N_5,In_253,In_416);
nor U6 (N_6,In_262,In_427);
nor U7 (N_7,In_418,In_462);
or U8 (N_8,In_412,In_48);
and U9 (N_9,In_240,In_49);
and U10 (N_10,In_233,In_120);
nand U11 (N_11,In_256,In_445);
nor U12 (N_12,In_465,In_26);
nor U13 (N_13,In_307,In_115);
and U14 (N_14,In_263,In_244);
or U15 (N_15,In_242,In_148);
or U16 (N_16,In_32,In_467);
or U17 (N_17,In_47,In_237);
and U18 (N_18,In_54,In_352);
and U19 (N_19,In_291,In_104);
nand U20 (N_20,In_353,In_274);
and U21 (N_21,In_431,In_391);
or U22 (N_22,In_371,In_20);
or U23 (N_23,In_411,In_152);
and U24 (N_24,In_284,In_174);
or U25 (N_25,In_209,In_436);
and U26 (N_26,In_144,In_325);
and U27 (N_27,In_33,In_278);
nand U28 (N_28,In_128,In_133);
and U29 (N_29,In_83,In_158);
and U30 (N_30,In_15,In_403);
and U31 (N_31,In_303,In_38);
nand U32 (N_32,In_215,In_27);
nor U33 (N_33,In_337,In_308);
and U34 (N_34,In_79,In_232);
nand U35 (N_35,In_390,In_169);
or U36 (N_36,In_107,In_134);
nand U37 (N_37,In_3,In_62);
nor U38 (N_38,In_276,In_488);
or U39 (N_39,In_135,In_175);
or U40 (N_40,In_167,In_499);
nand U41 (N_41,In_21,In_130);
nor U42 (N_42,In_199,In_282);
nand U43 (N_43,In_63,In_398);
and U44 (N_44,In_365,In_476);
and U45 (N_45,In_124,In_91);
and U46 (N_46,In_108,In_447);
nand U47 (N_47,In_397,In_59);
or U48 (N_48,In_45,In_340);
and U49 (N_49,In_245,In_203);
nand U50 (N_50,In_279,In_22);
nor U51 (N_51,In_320,In_331);
nand U52 (N_52,In_268,In_378);
nor U53 (N_53,In_40,In_487);
or U54 (N_54,In_28,In_463);
nor U55 (N_55,In_311,In_402);
or U56 (N_56,In_112,In_180);
nand U57 (N_57,In_294,In_344);
nor U58 (N_58,In_323,In_221);
nand U59 (N_59,In_10,In_142);
or U60 (N_60,N_17,In_188);
nor U61 (N_61,In_43,In_422);
and U62 (N_62,In_155,In_318);
nor U63 (N_63,In_299,In_35);
and U64 (N_64,In_78,In_216);
nand U65 (N_65,N_42,In_66);
xnor U66 (N_66,In_6,In_92);
nor U67 (N_67,In_448,In_80);
or U68 (N_68,N_5,In_7);
or U69 (N_69,In_251,In_145);
nand U70 (N_70,In_332,N_41);
nand U71 (N_71,N_0,In_410);
nand U72 (N_72,In_247,In_300);
and U73 (N_73,In_395,In_220);
nand U74 (N_74,In_129,In_154);
or U75 (N_75,N_30,In_290);
or U76 (N_76,In_490,In_457);
and U77 (N_77,In_305,In_351);
and U78 (N_78,In_29,In_428);
and U79 (N_79,In_179,In_470);
nor U80 (N_80,In_481,In_329);
or U81 (N_81,In_327,N_39);
or U82 (N_82,In_114,In_56);
nor U83 (N_83,In_460,In_342);
nor U84 (N_84,In_44,In_399);
nand U85 (N_85,In_304,N_48);
nand U86 (N_86,In_96,In_498);
xor U87 (N_87,In_440,In_408);
nand U88 (N_88,In_210,N_23);
and U89 (N_89,In_183,In_84);
and U90 (N_90,In_374,In_225);
nor U91 (N_91,In_37,In_100);
nand U92 (N_92,In_429,In_185);
and U93 (N_93,In_187,In_453);
or U94 (N_94,In_492,N_1);
nor U95 (N_95,In_361,N_21);
and U96 (N_96,In_444,In_286);
nand U97 (N_97,In_150,In_349);
and U98 (N_98,In_76,In_345);
nand U99 (N_99,In_302,In_25);
nor U100 (N_100,N_4,In_359);
nand U101 (N_101,In_275,In_5);
nand U102 (N_102,N_13,In_17);
and U103 (N_103,In_181,In_373);
nand U104 (N_104,In_370,In_341);
nand U105 (N_105,N_6,In_229);
and U106 (N_106,In_326,In_424);
and U107 (N_107,In_52,In_2);
nand U108 (N_108,In_354,N_31);
or U109 (N_109,In_136,In_228);
or U110 (N_110,In_99,In_170);
and U111 (N_111,In_451,N_56);
nor U112 (N_112,In_93,In_207);
nor U113 (N_113,In_118,N_40);
and U114 (N_114,In_11,In_479);
and U115 (N_115,In_392,In_313);
and U116 (N_116,In_23,In_211);
nand U117 (N_117,In_41,In_172);
or U118 (N_118,In_166,N_35);
or U119 (N_119,In_404,In_106);
or U120 (N_120,In_389,In_469);
and U121 (N_121,In_333,In_458);
nand U122 (N_122,In_420,In_423);
nand U123 (N_123,N_101,N_82);
or U124 (N_124,In_163,In_239);
nor U125 (N_125,In_64,In_36);
or U126 (N_126,In_330,In_149);
nor U127 (N_127,N_66,N_83);
nor U128 (N_128,In_277,In_139);
and U129 (N_129,In_9,In_461);
and U130 (N_130,In_312,In_393);
and U131 (N_131,N_3,In_213);
nand U132 (N_132,N_71,In_430);
or U133 (N_133,In_369,In_324);
nand U134 (N_134,N_108,In_18);
and U135 (N_135,In_443,N_58);
nor U136 (N_136,N_60,N_113);
or U137 (N_137,In_439,In_126);
nand U138 (N_138,In_71,N_117);
or U139 (N_139,In_226,In_189);
nand U140 (N_140,In_208,In_417);
and U141 (N_141,In_421,In_231);
or U142 (N_142,N_89,N_47);
and U143 (N_143,In_364,In_433);
and U144 (N_144,N_38,In_309);
nor U145 (N_145,In_75,In_259);
or U146 (N_146,In_217,In_4);
nand U147 (N_147,In_346,In_223);
nor U148 (N_148,In_362,In_317);
nor U149 (N_149,In_69,In_219);
or U150 (N_150,In_86,In_298);
nand U151 (N_151,In_474,In_413);
nand U152 (N_152,In_8,N_99);
and U153 (N_153,In_194,N_80);
and U154 (N_154,In_218,In_394);
or U155 (N_155,N_55,In_450);
or U156 (N_156,In_486,In_366);
nor U157 (N_157,In_57,In_103);
and U158 (N_158,In_125,In_68);
and U159 (N_159,In_319,In_200);
nor U160 (N_160,In_260,In_1);
nand U161 (N_161,In_292,In_385);
nor U162 (N_162,In_288,N_93);
or U163 (N_163,In_494,In_296);
and U164 (N_164,In_384,In_202);
and U165 (N_165,In_316,N_10);
and U166 (N_166,N_22,In_72);
or U167 (N_167,N_43,In_355);
nand U168 (N_168,N_61,In_388);
or U169 (N_169,In_137,In_272);
nand U170 (N_170,In_227,N_15);
or U171 (N_171,In_380,In_348);
nand U172 (N_172,In_249,N_52);
or U173 (N_173,In_254,In_101);
and U174 (N_174,In_238,In_98);
nand U175 (N_175,In_190,N_76);
nor U176 (N_176,In_24,In_281);
xnor U177 (N_177,N_59,In_97);
and U178 (N_178,N_72,N_19);
and U179 (N_179,In_236,N_94);
nor U180 (N_180,In_42,In_335);
and U181 (N_181,In_265,In_122);
nor U182 (N_182,N_104,In_471);
and U183 (N_183,N_63,N_166);
nand U184 (N_184,N_128,N_119);
and U185 (N_185,N_86,In_34);
and U186 (N_186,N_7,N_107);
and U187 (N_187,In_400,In_252);
and U188 (N_188,In_77,In_382);
nor U189 (N_189,In_426,In_153);
nor U190 (N_190,In_468,In_141);
or U191 (N_191,In_375,In_271);
nand U192 (N_192,N_148,In_295);
nor U193 (N_193,N_161,In_297);
nand U194 (N_194,In_198,N_169);
nand U195 (N_195,In_165,N_28);
or U196 (N_196,In_73,In_88);
nor U197 (N_197,In_482,In_178);
and U198 (N_198,In_123,In_435);
and U199 (N_199,N_74,N_154);
and U200 (N_200,In_39,In_127);
or U201 (N_201,In_350,N_162);
or U202 (N_202,N_65,In_478);
and U203 (N_203,In_119,In_480);
or U204 (N_204,In_168,In_206);
or U205 (N_205,N_45,N_173);
nor U206 (N_206,In_287,N_179);
nand U207 (N_207,N_159,In_184);
nor U208 (N_208,In_368,In_338);
and U209 (N_209,In_437,N_122);
nor U210 (N_210,In_89,N_88);
nand U211 (N_211,In_65,N_33);
and U212 (N_212,N_165,In_182);
and U213 (N_213,In_315,In_405);
nor U214 (N_214,In_314,In_201);
nor U215 (N_215,In_111,N_37);
and U216 (N_216,In_246,N_100);
nand U217 (N_217,N_120,In_310);
nor U218 (N_218,In_489,In_192);
nor U219 (N_219,In_248,N_106);
or U220 (N_220,In_13,In_459);
or U221 (N_221,N_95,N_115);
nand U222 (N_222,In_205,In_46);
nor U223 (N_223,In_51,In_379);
nor U224 (N_224,In_496,N_78);
nor U225 (N_225,In_406,In_306);
nand U226 (N_226,In_138,N_57);
and U227 (N_227,In_255,N_34);
nand U228 (N_228,In_53,In_257);
nor U229 (N_229,In_339,In_195);
or U230 (N_230,N_97,N_75);
and U231 (N_231,N_46,N_51);
or U232 (N_232,In_270,In_381);
nor U233 (N_233,N_24,N_150);
nor U234 (N_234,N_171,In_241);
or U235 (N_235,In_377,In_157);
or U236 (N_236,N_145,In_343);
or U237 (N_237,N_79,In_367);
nand U238 (N_238,N_32,N_11);
nand U239 (N_239,N_70,N_27);
and U240 (N_240,In_162,N_193);
or U241 (N_241,In_131,N_110);
and U242 (N_242,In_267,In_70);
nand U243 (N_243,N_232,N_164);
and U244 (N_244,N_50,N_233);
or U245 (N_245,In_105,In_109);
or U246 (N_246,In_243,N_160);
nor U247 (N_247,In_358,In_407);
nor U248 (N_248,N_139,In_197);
nor U249 (N_249,In_82,N_91);
and U250 (N_250,In_55,N_53);
or U251 (N_251,N_217,N_133);
nand U252 (N_252,N_174,N_90);
and U253 (N_253,In_477,N_235);
nor U254 (N_254,N_67,In_269);
and U255 (N_255,In_396,N_223);
nand U256 (N_256,In_164,N_111);
nor U257 (N_257,N_228,In_280);
or U258 (N_258,In_376,In_87);
or U259 (N_259,N_195,N_141);
or U260 (N_260,N_188,In_85);
nand U261 (N_261,In_386,N_182);
and U262 (N_262,In_483,N_134);
nor U263 (N_263,In_143,In_456);
and U264 (N_264,In_322,N_54);
and U265 (N_265,N_202,In_222);
and U266 (N_266,N_87,N_14);
and U267 (N_267,In_475,N_234);
and U268 (N_268,In_334,N_156);
and U269 (N_269,In_383,N_92);
and U270 (N_270,In_425,N_214);
nand U271 (N_271,In_363,N_219);
and U272 (N_272,N_125,N_138);
nor U273 (N_273,N_123,In_473);
nand U274 (N_274,N_98,In_357);
and U275 (N_275,In_193,N_26);
or U276 (N_276,In_485,N_18);
and U277 (N_277,N_168,In_146);
or U278 (N_278,In_176,In_264);
nor U279 (N_279,N_102,N_216);
nand U280 (N_280,In_454,N_62);
or U281 (N_281,N_142,N_158);
or U282 (N_282,In_273,In_360);
and U283 (N_283,N_212,In_434);
nor U284 (N_284,N_226,In_61);
nor U285 (N_285,N_203,N_170);
nand U286 (N_286,In_113,In_497);
and U287 (N_287,In_14,In_234);
nand U288 (N_288,N_121,N_178);
and U289 (N_289,N_105,In_12);
nor U290 (N_290,In_31,N_44);
and U291 (N_291,N_231,In_160);
nor U292 (N_292,N_25,N_49);
and U293 (N_293,In_121,N_124);
or U294 (N_294,N_143,N_176);
nor U295 (N_295,N_172,N_213);
nand U296 (N_296,In_102,N_207);
nand U297 (N_297,N_200,N_192);
or U298 (N_298,N_152,In_409);
nand U299 (N_299,N_84,N_191);
nor U300 (N_300,N_177,N_283);
or U301 (N_301,N_180,N_183);
and U302 (N_302,In_495,In_372);
and U303 (N_303,N_103,N_68);
nand U304 (N_304,In_293,In_186);
or U305 (N_305,In_387,N_272);
or U306 (N_306,N_282,In_438);
nand U307 (N_307,N_224,N_175);
nor U308 (N_308,N_238,N_208);
nand U309 (N_309,In_117,N_276);
nand U310 (N_310,N_215,In_16);
nor U311 (N_311,N_255,In_230);
and U312 (N_312,N_137,N_132);
and U313 (N_313,In_235,N_250);
nand U314 (N_314,N_151,In_401);
or U315 (N_315,N_278,In_442);
nor U316 (N_316,N_144,In_261);
or U317 (N_317,N_277,N_240);
and U318 (N_318,In_156,N_227);
nor U319 (N_319,In_484,N_273);
and U320 (N_320,N_96,N_64);
nor U321 (N_321,N_130,N_270);
or U322 (N_322,N_284,N_221);
or U323 (N_323,N_73,N_126);
nand U324 (N_324,N_146,N_299);
nor U325 (N_325,N_69,In_266);
nand U326 (N_326,N_112,N_243);
nand U327 (N_327,N_210,N_298);
and U328 (N_328,In_212,N_263);
or U329 (N_329,N_265,N_292);
and U330 (N_330,In_19,N_258);
or U331 (N_331,N_274,In_116);
and U332 (N_332,In_285,In_250);
and U333 (N_333,In_446,N_254);
nor U334 (N_334,N_225,N_262);
nand U335 (N_335,N_181,N_293);
nand U336 (N_336,In_336,N_194);
nand U337 (N_337,In_58,N_157);
or U338 (N_338,In_67,N_184);
nand U339 (N_339,In_455,N_187);
or U340 (N_340,In_95,N_163);
or U341 (N_341,N_189,In_140);
nor U342 (N_342,In_159,N_136);
nor U343 (N_343,N_186,N_241);
and U344 (N_344,In_171,N_260);
nor U345 (N_345,In_224,N_85);
nand U346 (N_346,In_466,N_155);
or U347 (N_347,In_258,N_256);
xor U348 (N_348,In_356,N_269);
and U349 (N_349,N_257,N_114);
or U350 (N_350,N_129,In_74);
and U351 (N_351,N_209,N_204);
nor U352 (N_352,N_9,In_81);
or U353 (N_353,N_252,N_237);
and U354 (N_354,N_239,N_109);
and U355 (N_355,N_266,N_294);
nor U356 (N_356,In_328,N_127);
or U357 (N_357,In_301,N_140);
and U358 (N_358,N_199,N_201);
and U359 (N_359,In_289,N_153);
or U360 (N_360,N_275,N_353);
nor U361 (N_361,N_334,N_147);
nor U362 (N_362,N_268,N_211);
and U363 (N_363,N_355,N_345);
or U364 (N_364,In_60,N_347);
or U365 (N_365,N_328,N_341);
and U366 (N_366,N_229,N_230);
and U367 (N_367,N_338,N_340);
nor U368 (N_368,N_354,N_196);
and U369 (N_369,N_8,N_306);
and U370 (N_370,N_346,N_322);
and U371 (N_371,In_449,N_245);
nor U372 (N_372,N_236,In_191);
nand U373 (N_373,N_330,N_327);
or U374 (N_374,N_323,N_185);
nand U375 (N_375,N_36,N_167);
nand U376 (N_376,N_206,N_296);
nor U377 (N_377,N_244,N_291);
or U378 (N_378,In_452,In_110);
and U379 (N_379,N_286,N_198);
nand U380 (N_380,N_319,In_0);
or U381 (N_381,In_50,N_12);
or U382 (N_382,N_310,N_29);
nand U383 (N_383,N_348,N_289);
and U384 (N_384,N_344,N_197);
or U385 (N_385,N_261,N_290);
and U386 (N_386,In_30,N_281);
or U387 (N_387,N_331,N_303);
or U388 (N_388,N_336,N_335);
nand U389 (N_389,N_343,N_300);
nor U390 (N_390,N_337,N_325);
and U391 (N_391,In_151,N_116);
and U392 (N_392,N_246,N_295);
and U393 (N_393,N_149,N_312);
or U394 (N_394,N_320,N_318);
and U395 (N_395,N_20,N_316);
nor U396 (N_396,N_324,N_287);
nand U397 (N_397,In_132,N_242);
or U398 (N_398,N_314,N_309);
nor U399 (N_399,N_259,N_81);
nand U400 (N_400,N_297,N_248);
or U401 (N_401,N_251,N_302);
nor U402 (N_402,N_288,N_222);
and U403 (N_403,N_220,N_205);
or U404 (N_404,In_173,N_247);
nand U405 (N_405,N_357,In_491);
nor U406 (N_406,In_321,N_350);
or U407 (N_407,N_333,N_131);
and U408 (N_408,N_317,N_315);
nand U409 (N_409,N_16,N_342);
nor U410 (N_410,N_305,N_321);
and U411 (N_411,N_339,In_432);
nand U412 (N_412,N_285,N_279);
nand U413 (N_413,N_271,N_359);
and U414 (N_414,N_349,N_307);
nand U415 (N_415,N_301,In_94);
and U416 (N_416,N_358,N_352);
nor U417 (N_417,N_264,N_135);
nand U418 (N_418,N_267,N_118);
and U419 (N_419,N_313,N_280);
or U420 (N_420,N_412,N_401);
nor U421 (N_421,N_400,N_409);
nand U422 (N_422,N_386,N_367);
or U423 (N_423,N_385,N_407);
or U424 (N_424,N_363,N_373);
nor U425 (N_425,N_402,N_408);
or U426 (N_426,N_395,N_404);
nor U427 (N_427,N_378,N_365);
or U428 (N_428,N_397,N_253);
or U429 (N_429,N_362,N_388);
and U430 (N_430,N_329,N_405);
and U431 (N_431,N_410,N_375);
or U432 (N_432,N_406,N_411);
and U433 (N_433,N_384,N_304);
nand U434 (N_434,N_391,N_332);
and U435 (N_435,N_379,N_380);
or U436 (N_436,In_204,In_415);
nor U437 (N_437,N_418,N_308);
and U438 (N_438,N_368,In_177);
nor U439 (N_439,N_311,N_416);
and U440 (N_440,N_413,N_415);
nor U441 (N_441,N_190,N_394);
or U442 (N_442,N_326,N_387);
nor U443 (N_443,N_389,In_472);
or U444 (N_444,N_351,N_377);
and U445 (N_445,N_399,N_356);
or U446 (N_446,In_214,N_218);
nand U447 (N_447,N_376,N_382);
and U448 (N_448,N_360,N_419);
nor U449 (N_449,N_403,N_390);
and U450 (N_450,N_417,N_396);
nand U451 (N_451,N_372,N_77);
or U452 (N_452,N_374,N_381);
nand U453 (N_453,N_2,N_398);
nor U454 (N_454,N_414,N_249);
nand U455 (N_455,N_370,N_392);
nor U456 (N_456,N_383,N_366);
or U457 (N_457,N_371,In_196);
nor U458 (N_458,N_369,N_393);
nand U459 (N_459,N_364,N_361);
nor U460 (N_460,N_329,N_397);
nand U461 (N_461,N_351,N_395);
or U462 (N_462,N_332,N_362);
and U463 (N_463,N_402,N_367);
nand U464 (N_464,N_408,N_382);
nor U465 (N_465,N_411,N_416);
or U466 (N_466,In_214,N_403);
nand U467 (N_467,N_218,N_404);
nand U468 (N_468,N_190,N_380);
nor U469 (N_469,N_332,N_372);
nand U470 (N_470,N_416,N_218);
nor U471 (N_471,N_410,N_408);
or U472 (N_472,N_404,N_329);
or U473 (N_473,N_411,N_385);
nor U474 (N_474,N_332,N_398);
nor U475 (N_475,In_196,N_253);
nand U476 (N_476,N_393,N_385);
nor U477 (N_477,N_249,N_403);
nand U478 (N_478,N_370,N_412);
or U479 (N_479,N_77,N_365);
and U480 (N_480,N_424,N_425);
nor U481 (N_481,N_470,N_459);
nor U482 (N_482,N_450,N_447);
or U483 (N_483,N_475,N_432);
nand U484 (N_484,N_448,N_439);
nand U485 (N_485,N_430,N_458);
and U486 (N_486,N_463,N_438);
nand U487 (N_487,N_465,N_473);
nor U488 (N_488,N_454,N_420);
nor U489 (N_489,N_443,N_440);
and U490 (N_490,N_474,N_423);
nor U491 (N_491,N_464,N_469);
or U492 (N_492,N_456,N_433);
nand U493 (N_493,N_446,N_452);
nor U494 (N_494,N_467,N_428);
and U495 (N_495,N_422,N_426);
nor U496 (N_496,N_476,N_427);
xnor U497 (N_497,N_442,N_479);
nand U498 (N_498,N_431,N_461);
nand U499 (N_499,N_444,N_421);
nand U500 (N_500,N_466,N_445);
or U501 (N_501,N_441,N_477);
nor U502 (N_502,N_449,N_429);
nand U503 (N_503,N_457,N_468);
nor U504 (N_504,N_460,N_437);
nor U505 (N_505,N_451,N_453);
nor U506 (N_506,N_462,N_471);
nor U507 (N_507,N_436,N_434);
nand U508 (N_508,N_455,N_435);
nor U509 (N_509,N_472,N_478);
or U510 (N_510,N_426,N_443);
and U511 (N_511,N_463,N_430);
or U512 (N_512,N_479,N_452);
nor U513 (N_513,N_430,N_438);
nand U514 (N_514,N_470,N_439);
nand U515 (N_515,N_425,N_444);
nor U516 (N_516,N_441,N_456);
nand U517 (N_517,N_437,N_479);
and U518 (N_518,N_469,N_461);
nand U519 (N_519,N_433,N_462);
nor U520 (N_520,N_463,N_478);
and U521 (N_521,N_471,N_428);
nor U522 (N_522,N_447,N_442);
nand U523 (N_523,N_476,N_435);
and U524 (N_524,N_428,N_459);
nand U525 (N_525,N_474,N_478);
and U526 (N_526,N_439,N_426);
and U527 (N_527,N_479,N_463);
nor U528 (N_528,N_435,N_421);
and U529 (N_529,N_430,N_462);
nor U530 (N_530,N_462,N_441);
nor U531 (N_531,N_476,N_458);
and U532 (N_532,N_439,N_453);
nor U533 (N_533,N_429,N_430);
or U534 (N_534,N_443,N_425);
nand U535 (N_535,N_451,N_478);
and U536 (N_536,N_451,N_455);
nor U537 (N_537,N_462,N_420);
and U538 (N_538,N_461,N_433);
or U539 (N_539,N_477,N_465);
or U540 (N_540,N_486,N_502);
or U541 (N_541,N_537,N_520);
nor U542 (N_542,N_485,N_529);
and U543 (N_543,N_507,N_501);
and U544 (N_544,N_500,N_492);
or U545 (N_545,N_512,N_498);
nand U546 (N_546,N_505,N_523);
and U547 (N_547,N_503,N_535);
or U548 (N_548,N_511,N_524);
nand U549 (N_549,N_532,N_496);
or U550 (N_550,N_488,N_521);
nand U551 (N_551,N_517,N_493);
nor U552 (N_552,N_515,N_489);
nor U553 (N_553,N_483,N_504);
and U554 (N_554,N_530,N_538);
or U555 (N_555,N_484,N_518);
nand U556 (N_556,N_527,N_522);
nor U557 (N_557,N_508,N_533);
or U558 (N_558,N_480,N_506);
or U559 (N_559,N_539,N_536);
nand U560 (N_560,N_490,N_516);
nand U561 (N_561,N_526,N_482);
or U562 (N_562,N_534,N_531);
and U563 (N_563,N_514,N_513);
nor U564 (N_564,N_494,N_491);
nor U565 (N_565,N_519,N_481);
nand U566 (N_566,N_487,N_497);
nand U567 (N_567,N_528,N_499);
or U568 (N_568,N_510,N_495);
nand U569 (N_569,N_525,N_509);
xor U570 (N_570,N_496,N_492);
nor U571 (N_571,N_512,N_501);
nand U572 (N_572,N_536,N_535);
or U573 (N_573,N_516,N_498);
and U574 (N_574,N_486,N_531);
nand U575 (N_575,N_502,N_525);
nor U576 (N_576,N_536,N_500);
and U577 (N_577,N_529,N_490);
nand U578 (N_578,N_504,N_503);
nor U579 (N_579,N_484,N_496);
and U580 (N_580,N_512,N_500);
nand U581 (N_581,N_531,N_509);
and U582 (N_582,N_482,N_514);
nand U583 (N_583,N_497,N_514);
and U584 (N_584,N_524,N_497);
nand U585 (N_585,N_493,N_524);
or U586 (N_586,N_485,N_533);
or U587 (N_587,N_513,N_502);
nand U588 (N_588,N_531,N_490);
nor U589 (N_589,N_517,N_528);
nand U590 (N_590,N_526,N_493);
and U591 (N_591,N_487,N_533);
and U592 (N_592,N_501,N_534);
nand U593 (N_593,N_511,N_525);
nor U594 (N_594,N_507,N_534);
nor U595 (N_595,N_489,N_525);
and U596 (N_596,N_533,N_500);
nor U597 (N_597,N_536,N_480);
nor U598 (N_598,N_489,N_491);
or U599 (N_599,N_518,N_485);
nand U600 (N_600,N_572,N_551);
nand U601 (N_601,N_552,N_595);
nand U602 (N_602,N_593,N_588);
or U603 (N_603,N_574,N_582);
nor U604 (N_604,N_556,N_550);
and U605 (N_605,N_585,N_583);
nand U606 (N_606,N_561,N_569);
and U607 (N_607,N_553,N_554);
or U608 (N_608,N_562,N_565);
nand U609 (N_609,N_568,N_558);
and U610 (N_610,N_559,N_541);
nand U611 (N_611,N_589,N_560);
nor U612 (N_612,N_548,N_540);
nor U613 (N_613,N_557,N_543);
nor U614 (N_614,N_587,N_546);
nor U615 (N_615,N_597,N_584);
or U616 (N_616,N_575,N_599);
nand U617 (N_617,N_547,N_567);
nand U618 (N_618,N_570,N_598);
nor U619 (N_619,N_590,N_579);
nand U620 (N_620,N_573,N_544);
or U621 (N_621,N_591,N_586);
nand U622 (N_622,N_577,N_592);
nand U623 (N_623,N_566,N_576);
and U624 (N_624,N_594,N_596);
nor U625 (N_625,N_564,N_578);
nor U626 (N_626,N_545,N_563);
nor U627 (N_627,N_571,N_555);
and U628 (N_628,N_549,N_580);
nand U629 (N_629,N_581,N_542);
or U630 (N_630,N_568,N_559);
nand U631 (N_631,N_570,N_581);
or U632 (N_632,N_582,N_570);
nand U633 (N_633,N_560,N_567);
or U634 (N_634,N_579,N_596);
nand U635 (N_635,N_584,N_575);
nor U636 (N_636,N_592,N_554);
or U637 (N_637,N_544,N_597);
and U638 (N_638,N_540,N_562);
or U639 (N_639,N_595,N_583);
nor U640 (N_640,N_597,N_554);
nand U641 (N_641,N_592,N_548);
nand U642 (N_642,N_563,N_544);
or U643 (N_643,N_583,N_587);
and U644 (N_644,N_557,N_583);
or U645 (N_645,N_585,N_590);
and U646 (N_646,N_555,N_576);
or U647 (N_647,N_568,N_595);
nor U648 (N_648,N_552,N_576);
or U649 (N_649,N_567,N_566);
nor U650 (N_650,N_551,N_598);
nand U651 (N_651,N_586,N_575);
nor U652 (N_652,N_597,N_596);
nor U653 (N_653,N_552,N_555);
nand U654 (N_654,N_559,N_588);
nor U655 (N_655,N_584,N_588);
nand U656 (N_656,N_549,N_561);
or U657 (N_657,N_542,N_566);
and U658 (N_658,N_589,N_583);
nand U659 (N_659,N_564,N_559);
or U660 (N_660,N_645,N_608);
and U661 (N_661,N_635,N_619);
or U662 (N_662,N_607,N_637);
nand U663 (N_663,N_600,N_625);
nor U664 (N_664,N_640,N_659);
nor U665 (N_665,N_605,N_615);
nand U666 (N_666,N_638,N_631);
nor U667 (N_667,N_653,N_606);
and U668 (N_668,N_610,N_626);
or U669 (N_669,N_627,N_618);
or U670 (N_670,N_646,N_658);
and U671 (N_671,N_629,N_655);
nand U672 (N_672,N_654,N_623);
nor U673 (N_673,N_632,N_642);
or U674 (N_674,N_603,N_641);
or U675 (N_675,N_620,N_647);
and U676 (N_676,N_630,N_652);
or U677 (N_677,N_611,N_639);
nor U678 (N_678,N_621,N_609);
nand U679 (N_679,N_601,N_657);
and U680 (N_680,N_613,N_633);
and U681 (N_681,N_602,N_644);
nand U682 (N_682,N_616,N_634);
nand U683 (N_683,N_650,N_617);
or U684 (N_684,N_612,N_614);
nand U685 (N_685,N_648,N_628);
nand U686 (N_686,N_636,N_649);
and U687 (N_687,N_643,N_656);
and U688 (N_688,N_624,N_604);
and U689 (N_689,N_622,N_651);
and U690 (N_690,N_657,N_658);
and U691 (N_691,N_656,N_620);
nand U692 (N_692,N_613,N_604);
or U693 (N_693,N_616,N_603);
or U694 (N_694,N_601,N_631);
and U695 (N_695,N_629,N_620);
nor U696 (N_696,N_645,N_605);
nand U697 (N_697,N_633,N_636);
nor U698 (N_698,N_624,N_646);
or U699 (N_699,N_659,N_645);
and U700 (N_700,N_648,N_653);
nor U701 (N_701,N_625,N_623);
nand U702 (N_702,N_648,N_651);
nand U703 (N_703,N_635,N_604);
or U704 (N_704,N_612,N_600);
nand U705 (N_705,N_649,N_630);
nor U706 (N_706,N_640,N_631);
nor U707 (N_707,N_641,N_613);
nor U708 (N_708,N_619,N_606);
nor U709 (N_709,N_606,N_602);
or U710 (N_710,N_600,N_628);
nor U711 (N_711,N_603,N_628);
nor U712 (N_712,N_600,N_630);
and U713 (N_713,N_602,N_638);
xor U714 (N_714,N_656,N_609);
or U715 (N_715,N_656,N_644);
or U716 (N_716,N_610,N_619);
nor U717 (N_717,N_655,N_640);
or U718 (N_718,N_627,N_603);
or U719 (N_719,N_620,N_615);
or U720 (N_720,N_668,N_700);
nor U721 (N_721,N_679,N_713);
nand U722 (N_722,N_663,N_660);
nand U723 (N_723,N_695,N_669);
and U724 (N_724,N_705,N_677);
or U725 (N_725,N_692,N_662);
nand U726 (N_726,N_698,N_707);
nor U727 (N_727,N_687,N_672);
and U728 (N_728,N_680,N_682);
and U729 (N_729,N_708,N_703);
nor U730 (N_730,N_702,N_673);
and U731 (N_731,N_696,N_694);
and U732 (N_732,N_709,N_719);
and U733 (N_733,N_685,N_710);
or U734 (N_734,N_717,N_714);
and U735 (N_735,N_661,N_718);
nor U736 (N_736,N_715,N_674);
nand U737 (N_737,N_666,N_684);
or U738 (N_738,N_688,N_678);
and U739 (N_739,N_689,N_670);
and U740 (N_740,N_701,N_665);
and U741 (N_741,N_712,N_681);
nor U742 (N_742,N_693,N_716);
and U743 (N_743,N_697,N_704);
nor U744 (N_744,N_691,N_675);
nand U745 (N_745,N_699,N_686);
nand U746 (N_746,N_711,N_667);
or U747 (N_747,N_664,N_676);
nand U748 (N_748,N_683,N_690);
and U749 (N_749,N_706,N_671);
or U750 (N_750,N_702,N_676);
nor U751 (N_751,N_675,N_718);
nand U752 (N_752,N_689,N_682);
or U753 (N_753,N_703,N_698);
and U754 (N_754,N_696,N_664);
or U755 (N_755,N_674,N_700);
nor U756 (N_756,N_662,N_690);
xnor U757 (N_757,N_686,N_689);
nand U758 (N_758,N_695,N_712);
and U759 (N_759,N_700,N_661);
nand U760 (N_760,N_699,N_666);
and U761 (N_761,N_719,N_672);
and U762 (N_762,N_661,N_710);
nor U763 (N_763,N_707,N_701);
or U764 (N_764,N_705,N_714);
and U765 (N_765,N_696,N_713);
and U766 (N_766,N_682,N_704);
nand U767 (N_767,N_700,N_718);
nand U768 (N_768,N_679,N_688);
or U769 (N_769,N_710,N_700);
and U770 (N_770,N_706,N_716);
and U771 (N_771,N_713,N_717);
and U772 (N_772,N_709,N_704);
nor U773 (N_773,N_673,N_705);
nor U774 (N_774,N_673,N_717);
nand U775 (N_775,N_710,N_718);
nor U776 (N_776,N_675,N_670);
or U777 (N_777,N_681,N_663);
or U778 (N_778,N_676,N_719);
nand U779 (N_779,N_677,N_689);
and U780 (N_780,N_729,N_770);
nand U781 (N_781,N_751,N_779);
and U782 (N_782,N_722,N_743);
nand U783 (N_783,N_745,N_734);
and U784 (N_784,N_721,N_767);
xnor U785 (N_785,N_761,N_758);
nand U786 (N_786,N_750,N_733);
or U787 (N_787,N_731,N_742);
nand U788 (N_788,N_772,N_764);
nand U789 (N_789,N_773,N_741);
nor U790 (N_790,N_724,N_725);
nor U791 (N_791,N_777,N_775);
and U792 (N_792,N_723,N_753);
or U793 (N_793,N_765,N_762);
or U794 (N_794,N_740,N_763);
or U795 (N_795,N_726,N_749);
or U796 (N_796,N_759,N_776);
nand U797 (N_797,N_768,N_747);
nand U798 (N_798,N_735,N_737);
nor U799 (N_799,N_736,N_755);
and U800 (N_800,N_730,N_752);
nor U801 (N_801,N_744,N_774);
nand U802 (N_802,N_771,N_728);
or U803 (N_803,N_760,N_748);
and U804 (N_804,N_757,N_732);
nor U805 (N_805,N_756,N_727);
nor U806 (N_806,N_754,N_769);
and U807 (N_807,N_766,N_720);
nand U808 (N_808,N_739,N_746);
or U809 (N_809,N_778,N_738);
nor U810 (N_810,N_739,N_775);
nor U811 (N_811,N_770,N_758);
and U812 (N_812,N_749,N_754);
and U813 (N_813,N_756,N_740);
nor U814 (N_814,N_776,N_779);
nand U815 (N_815,N_753,N_775);
and U816 (N_816,N_776,N_747);
or U817 (N_817,N_767,N_778);
nor U818 (N_818,N_725,N_779);
or U819 (N_819,N_763,N_760);
nand U820 (N_820,N_746,N_738);
nand U821 (N_821,N_721,N_745);
and U822 (N_822,N_758,N_741);
nor U823 (N_823,N_765,N_721);
or U824 (N_824,N_777,N_759);
or U825 (N_825,N_734,N_773);
nor U826 (N_826,N_754,N_728);
and U827 (N_827,N_733,N_721);
or U828 (N_828,N_756,N_772);
and U829 (N_829,N_750,N_745);
nand U830 (N_830,N_750,N_759);
nor U831 (N_831,N_768,N_760);
nand U832 (N_832,N_740,N_730);
or U833 (N_833,N_743,N_773);
nand U834 (N_834,N_744,N_778);
or U835 (N_835,N_756,N_732);
or U836 (N_836,N_774,N_739);
nor U837 (N_837,N_755,N_772);
nand U838 (N_838,N_760,N_772);
or U839 (N_839,N_751,N_764);
nor U840 (N_840,N_810,N_815);
and U841 (N_841,N_784,N_811);
and U842 (N_842,N_823,N_838);
or U843 (N_843,N_827,N_804);
nand U844 (N_844,N_817,N_835);
and U845 (N_845,N_783,N_795);
nand U846 (N_846,N_808,N_809);
nor U847 (N_847,N_813,N_794);
and U848 (N_848,N_806,N_820);
and U849 (N_849,N_802,N_785);
nor U850 (N_850,N_781,N_819);
or U851 (N_851,N_824,N_826);
and U852 (N_852,N_816,N_798);
nor U853 (N_853,N_796,N_807);
nand U854 (N_854,N_829,N_833);
or U855 (N_855,N_786,N_793);
nor U856 (N_856,N_831,N_799);
and U857 (N_857,N_787,N_832);
nor U858 (N_858,N_801,N_821);
and U859 (N_859,N_818,N_834);
nor U860 (N_860,N_822,N_814);
nand U861 (N_861,N_803,N_828);
nor U862 (N_862,N_800,N_780);
nand U863 (N_863,N_839,N_788);
nand U864 (N_864,N_836,N_791);
or U865 (N_865,N_797,N_782);
and U866 (N_866,N_789,N_825);
and U867 (N_867,N_837,N_830);
nand U868 (N_868,N_812,N_792);
or U869 (N_869,N_805,N_790);
and U870 (N_870,N_828,N_808);
nand U871 (N_871,N_783,N_791);
and U872 (N_872,N_831,N_823);
and U873 (N_873,N_819,N_806);
nand U874 (N_874,N_831,N_810);
nor U875 (N_875,N_799,N_823);
nor U876 (N_876,N_808,N_801);
and U877 (N_877,N_820,N_833);
nor U878 (N_878,N_814,N_815);
nand U879 (N_879,N_830,N_809);
nor U880 (N_880,N_830,N_832);
or U881 (N_881,N_819,N_833);
nand U882 (N_882,N_815,N_836);
nor U883 (N_883,N_809,N_837);
or U884 (N_884,N_833,N_788);
nand U885 (N_885,N_787,N_824);
and U886 (N_886,N_794,N_821);
xor U887 (N_887,N_790,N_808);
or U888 (N_888,N_791,N_805);
or U889 (N_889,N_827,N_829);
nand U890 (N_890,N_839,N_801);
or U891 (N_891,N_800,N_833);
nand U892 (N_892,N_834,N_788);
nand U893 (N_893,N_839,N_794);
and U894 (N_894,N_837,N_797);
or U895 (N_895,N_798,N_807);
or U896 (N_896,N_791,N_798);
or U897 (N_897,N_782,N_790);
nand U898 (N_898,N_788,N_810);
nor U899 (N_899,N_812,N_838);
and U900 (N_900,N_857,N_846);
or U901 (N_901,N_878,N_866);
and U902 (N_902,N_884,N_886);
or U903 (N_903,N_841,N_844);
nor U904 (N_904,N_862,N_871);
nor U905 (N_905,N_861,N_860);
and U906 (N_906,N_891,N_864);
and U907 (N_907,N_850,N_895);
and U908 (N_908,N_897,N_855);
and U909 (N_909,N_856,N_892);
or U910 (N_910,N_868,N_840);
or U911 (N_911,N_875,N_843);
or U912 (N_912,N_848,N_881);
or U913 (N_913,N_893,N_845);
nand U914 (N_914,N_869,N_852);
nor U915 (N_915,N_896,N_898);
nor U916 (N_916,N_858,N_876);
nor U917 (N_917,N_859,N_867);
nor U918 (N_918,N_899,N_894);
nand U919 (N_919,N_883,N_847);
nor U920 (N_920,N_854,N_872);
nand U921 (N_921,N_863,N_889);
nor U922 (N_922,N_849,N_870);
nand U923 (N_923,N_865,N_842);
and U924 (N_924,N_882,N_880);
and U925 (N_925,N_853,N_851);
nor U926 (N_926,N_887,N_874);
nor U927 (N_927,N_877,N_888);
nor U928 (N_928,N_885,N_873);
nor U929 (N_929,N_890,N_879);
or U930 (N_930,N_878,N_887);
or U931 (N_931,N_872,N_890);
nand U932 (N_932,N_849,N_895);
or U933 (N_933,N_879,N_877);
or U934 (N_934,N_866,N_853);
and U935 (N_935,N_852,N_848);
and U936 (N_936,N_853,N_842);
nand U937 (N_937,N_873,N_896);
and U938 (N_938,N_872,N_864);
nand U939 (N_939,N_899,N_845);
or U940 (N_940,N_853,N_860);
and U941 (N_941,N_881,N_854);
nor U942 (N_942,N_894,N_865);
or U943 (N_943,N_886,N_881);
or U944 (N_944,N_875,N_882);
nor U945 (N_945,N_887,N_897);
or U946 (N_946,N_893,N_848);
and U947 (N_947,N_860,N_889);
and U948 (N_948,N_843,N_853);
or U949 (N_949,N_897,N_881);
and U950 (N_950,N_855,N_876);
nand U951 (N_951,N_887,N_886);
or U952 (N_952,N_880,N_890);
or U953 (N_953,N_853,N_892);
and U954 (N_954,N_876,N_877);
or U955 (N_955,N_888,N_860);
nand U956 (N_956,N_898,N_845);
nand U957 (N_957,N_881,N_872);
nor U958 (N_958,N_895,N_899);
or U959 (N_959,N_872,N_878);
and U960 (N_960,N_946,N_948);
nor U961 (N_961,N_902,N_921);
or U962 (N_962,N_944,N_923);
nor U963 (N_963,N_952,N_915);
or U964 (N_964,N_925,N_926);
and U965 (N_965,N_910,N_909);
nand U966 (N_966,N_945,N_932);
nor U967 (N_967,N_922,N_907);
and U968 (N_968,N_955,N_937);
or U969 (N_969,N_953,N_934);
nor U970 (N_970,N_956,N_958);
nand U971 (N_971,N_905,N_942);
nor U972 (N_972,N_901,N_912);
and U973 (N_973,N_919,N_914);
or U974 (N_974,N_935,N_959);
and U975 (N_975,N_911,N_927);
nand U976 (N_976,N_936,N_951);
nand U977 (N_977,N_930,N_900);
or U978 (N_978,N_904,N_928);
or U979 (N_979,N_938,N_917);
or U980 (N_980,N_906,N_933);
nor U981 (N_981,N_940,N_916);
nand U982 (N_982,N_939,N_929);
nand U983 (N_983,N_924,N_950);
and U984 (N_984,N_913,N_943);
nand U985 (N_985,N_920,N_908);
and U986 (N_986,N_903,N_918);
or U987 (N_987,N_931,N_947);
nor U988 (N_988,N_954,N_957);
nand U989 (N_989,N_941,N_949);
nand U990 (N_990,N_945,N_941);
nand U991 (N_991,N_929,N_936);
and U992 (N_992,N_946,N_935);
nand U993 (N_993,N_943,N_904);
or U994 (N_994,N_905,N_915);
nand U995 (N_995,N_932,N_922);
xor U996 (N_996,N_949,N_954);
nand U997 (N_997,N_954,N_914);
or U998 (N_998,N_927,N_905);
and U999 (N_999,N_935,N_904);
and U1000 (N_1000,N_957,N_901);
nand U1001 (N_1001,N_957,N_900);
nor U1002 (N_1002,N_940,N_929);
nor U1003 (N_1003,N_912,N_957);
or U1004 (N_1004,N_952,N_905);
and U1005 (N_1005,N_945,N_950);
nand U1006 (N_1006,N_913,N_954);
nor U1007 (N_1007,N_908,N_938);
or U1008 (N_1008,N_919,N_933);
nor U1009 (N_1009,N_959,N_955);
and U1010 (N_1010,N_913,N_917);
and U1011 (N_1011,N_927,N_956);
and U1012 (N_1012,N_959,N_901);
nor U1013 (N_1013,N_935,N_934);
nor U1014 (N_1014,N_935,N_909);
nand U1015 (N_1015,N_959,N_917);
or U1016 (N_1016,N_950,N_921);
nand U1017 (N_1017,N_920,N_952);
nand U1018 (N_1018,N_947,N_949);
nor U1019 (N_1019,N_923,N_946);
nor U1020 (N_1020,N_1007,N_975);
nor U1021 (N_1021,N_969,N_978);
nand U1022 (N_1022,N_964,N_1001);
or U1023 (N_1023,N_992,N_1017);
nor U1024 (N_1024,N_1016,N_990);
nor U1025 (N_1025,N_982,N_966);
and U1026 (N_1026,N_985,N_1005);
or U1027 (N_1027,N_1006,N_1009);
and U1028 (N_1028,N_1011,N_1015);
and U1029 (N_1029,N_994,N_1010);
or U1030 (N_1030,N_971,N_965);
nand U1031 (N_1031,N_989,N_974);
and U1032 (N_1032,N_997,N_999);
nand U1033 (N_1033,N_977,N_991);
xnor U1034 (N_1034,N_968,N_972);
or U1035 (N_1035,N_979,N_973);
or U1036 (N_1036,N_976,N_963);
nand U1037 (N_1037,N_980,N_967);
and U1038 (N_1038,N_993,N_988);
and U1039 (N_1039,N_984,N_1004);
or U1040 (N_1040,N_1018,N_998);
or U1041 (N_1041,N_1003,N_987);
and U1042 (N_1042,N_970,N_1012);
or U1043 (N_1043,N_961,N_1013);
nand U1044 (N_1044,N_981,N_1019);
nand U1045 (N_1045,N_962,N_1014);
and U1046 (N_1046,N_960,N_1008);
or U1047 (N_1047,N_995,N_1000);
nand U1048 (N_1048,N_983,N_1002);
and U1049 (N_1049,N_996,N_986);
or U1050 (N_1050,N_979,N_1004);
or U1051 (N_1051,N_991,N_982);
nand U1052 (N_1052,N_967,N_979);
or U1053 (N_1053,N_993,N_963);
and U1054 (N_1054,N_981,N_962);
nand U1055 (N_1055,N_979,N_1016);
nand U1056 (N_1056,N_1015,N_991);
nor U1057 (N_1057,N_1003,N_981);
or U1058 (N_1058,N_978,N_1010);
or U1059 (N_1059,N_968,N_975);
nor U1060 (N_1060,N_1012,N_991);
or U1061 (N_1061,N_964,N_994);
nor U1062 (N_1062,N_986,N_969);
nor U1063 (N_1063,N_968,N_970);
nor U1064 (N_1064,N_1018,N_979);
nor U1065 (N_1065,N_1018,N_980);
nand U1066 (N_1066,N_1018,N_999);
nand U1067 (N_1067,N_975,N_974);
or U1068 (N_1068,N_961,N_1003);
and U1069 (N_1069,N_999,N_980);
nor U1070 (N_1070,N_1015,N_982);
nor U1071 (N_1071,N_976,N_968);
nand U1072 (N_1072,N_1009,N_965);
nand U1073 (N_1073,N_963,N_962);
and U1074 (N_1074,N_1019,N_987);
nand U1075 (N_1075,N_963,N_1000);
nor U1076 (N_1076,N_960,N_989);
or U1077 (N_1077,N_989,N_1010);
nand U1078 (N_1078,N_1017,N_986);
nand U1079 (N_1079,N_979,N_976);
nor U1080 (N_1080,N_1077,N_1062);
nand U1081 (N_1081,N_1058,N_1076);
nand U1082 (N_1082,N_1021,N_1065);
nor U1083 (N_1083,N_1064,N_1079);
or U1084 (N_1084,N_1059,N_1067);
and U1085 (N_1085,N_1048,N_1052);
nor U1086 (N_1086,N_1068,N_1045);
nand U1087 (N_1087,N_1050,N_1035);
nor U1088 (N_1088,N_1022,N_1039);
or U1089 (N_1089,N_1032,N_1031);
nor U1090 (N_1090,N_1028,N_1053);
and U1091 (N_1091,N_1033,N_1049);
nor U1092 (N_1092,N_1072,N_1051);
nor U1093 (N_1093,N_1061,N_1060);
and U1094 (N_1094,N_1026,N_1040);
and U1095 (N_1095,N_1038,N_1070);
and U1096 (N_1096,N_1057,N_1066);
nand U1097 (N_1097,N_1044,N_1075);
and U1098 (N_1098,N_1025,N_1063);
or U1099 (N_1099,N_1042,N_1029);
or U1100 (N_1100,N_1078,N_1041);
nand U1101 (N_1101,N_1037,N_1030);
nor U1102 (N_1102,N_1055,N_1056);
nor U1103 (N_1103,N_1069,N_1054);
xnor U1104 (N_1104,N_1034,N_1047);
and U1105 (N_1105,N_1020,N_1024);
or U1106 (N_1106,N_1071,N_1074);
or U1107 (N_1107,N_1043,N_1073);
or U1108 (N_1108,N_1023,N_1036);
nand U1109 (N_1109,N_1046,N_1027);
nand U1110 (N_1110,N_1059,N_1021);
or U1111 (N_1111,N_1049,N_1035);
nand U1112 (N_1112,N_1071,N_1056);
or U1113 (N_1113,N_1071,N_1079);
nor U1114 (N_1114,N_1030,N_1067);
nor U1115 (N_1115,N_1026,N_1063);
nand U1116 (N_1116,N_1046,N_1073);
nand U1117 (N_1117,N_1030,N_1061);
nor U1118 (N_1118,N_1047,N_1066);
nand U1119 (N_1119,N_1038,N_1043);
nor U1120 (N_1120,N_1023,N_1077);
or U1121 (N_1121,N_1059,N_1075);
or U1122 (N_1122,N_1049,N_1071);
nand U1123 (N_1123,N_1068,N_1048);
xnor U1124 (N_1124,N_1026,N_1029);
xor U1125 (N_1125,N_1058,N_1055);
and U1126 (N_1126,N_1024,N_1028);
nor U1127 (N_1127,N_1024,N_1030);
nor U1128 (N_1128,N_1024,N_1063);
nor U1129 (N_1129,N_1026,N_1043);
and U1130 (N_1130,N_1034,N_1046);
nor U1131 (N_1131,N_1077,N_1067);
or U1132 (N_1132,N_1065,N_1047);
or U1133 (N_1133,N_1053,N_1063);
or U1134 (N_1134,N_1063,N_1038);
nand U1135 (N_1135,N_1059,N_1024);
or U1136 (N_1136,N_1071,N_1059);
and U1137 (N_1137,N_1077,N_1051);
or U1138 (N_1138,N_1053,N_1030);
nor U1139 (N_1139,N_1078,N_1076);
and U1140 (N_1140,N_1083,N_1126);
nor U1141 (N_1141,N_1115,N_1117);
or U1142 (N_1142,N_1134,N_1121);
nand U1143 (N_1143,N_1128,N_1086);
nor U1144 (N_1144,N_1123,N_1087);
or U1145 (N_1145,N_1080,N_1082);
nor U1146 (N_1146,N_1139,N_1116);
nor U1147 (N_1147,N_1081,N_1133);
nor U1148 (N_1148,N_1138,N_1135);
nor U1149 (N_1149,N_1127,N_1098);
nand U1150 (N_1150,N_1103,N_1122);
and U1151 (N_1151,N_1119,N_1118);
nand U1152 (N_1152,N_1102,N_1093);
nand U1153 (N_1153,N_1091,N_1090);
or U1154 (N_1154,N_1110,N_1111);
nor U1155 (N_1155,N_1131,N_1094);
and U1156 (N_1156,N_1100,N_1114);
nor U1157 (N_1157,N_1088,N_1109);
and U1158 (N_1158,N_1101,N_1095);
or U1159 (N_1159,N_1108,N_1105);
or U1160 (N_1160,N_1136,N_1112);
nor U1161 (N_1161,N_1113,N_1089);
or U1162 (N_1162,N_1099,N_1124);
nor U1163 (N_1163,N_1084,N_1130);
nand U1164 (N_1164,N_1125,N_1120);
nand U1165 (N_1165,N_1092,N_1129);
xor U1166 (N_1166,N_1104,N_1137);
nand U1167 (N_1167,N_1132,N_1085);
nand U1168 (N_1168,N_1106,N_1097);
and U1169 (N_1169,N_1096,N_1107);
or U1170 (N_1170,N_1090,N_1101);
nand U1171 (N_1171,N_1133,N_1086);
nor U1172 (N_1172,N_1107,N_1115);
nand U1173 (N_1173,N_1129,N_1111);
nor U1174 (N_1174,N_1132,N_1082);
and U1175 (N_1175,N_1106,N_1096);
nor U1176 (N_1176,N_1092,N_1084);
nand U1177 (N_1177,N_1091,N_1139);
nor U1178 (N_1178,N_1129,N_1131);
or U1179 (N_1179,N_1080,N_1093);
or U1180 (N_1180,N_1084,N_1121);
nor U1181 (N_1181,N_1131,N_1097);
nor U1182 (N_1182,N_1120,N_1082);
nand U1183 (N_1183,N_1117,N_1101);
and U1184 (N_1184,N_1115,N_1113);
or U1185 (N_1185,N_1134,N_1098);
nor U1186 (N_1186,N_1114,N_1091);
or U1187 (N_1187,N_1084,N_1131);
nor U1188 (N_1188,N_1111,N_1122);
and U1189 (N_1189,N_1105,N_1121);
nor U1190 (N_1190,N_1114,N_1115);
nor U1191 (N_1191,N_1112,N_1101);
nor U1192 (N_1192,N_1124,N_1111);
or U1193 (N_1193,N_1105,N_1081);
nand U1194 (N_1194,N_1111,N_1114);
or U1195 (N_1195,N_1124,N_1133);
and U1196 (N_1196,N_1134,N_1116);
nand U1197 (N_1197,N_1125,N_1138);
or U1198 (N_1198,N_1085,N_1113);
nor U1199 (N_1199,N_1106,N_1098);
nor U1200 (N_1200,N_1155,N_1147);
nand U1201 (N_1201,N_1198,N_1188);
nor U1202 (N_1202,N_1191,N_1152);
nand U1203 (N_1203,N_1150,N_1180);
and U1204 (N_1204,N_1193,N_1199);
and U1205 (N_1205,N_1179,N_1169);
and U1206 (N_1206,N_1149,N_1183);
nand U1207 (N_1207,N_1192,N_1151);
nand U1208 (N_1208,N_1161,N_1178);
and U1209 (N_1209,N_1166,N_1141);
nand U1210 (N_1210,N_1148,N_1196);
nand U1211 (N_1211,N_1158,N_1164);
or U1212 (N_1212,N_1140,N_1189);
or U1213 (N_1213,N_1176,N_1153);
nor U1214 (N_1214,N_1143,N_1187);
nor U1215 (N_1215,N_1163,N_1195);
nor U1216 (N_1216,N_1165,N_1162);
and U1217 (N_1217,N_1156,N_1190);
nor U1218 (N_1218,N_1184,N_1174);
and U1219 (N_1219,N_1177,N_1144);
nor U1220 (N_1220,N_1159,N_1181);
or U1221 (N_1221,N_1142,N_1154);
or U1222 (N_1222,N_1168,N_1186);
nand U1223 (N_1223,N_1172,N_1175);
nand U1224 (N_1224,N_1145,N_1167);
and U1225 (N_1225,N_1170,N_1157);
nor U1226 (N_1226,N_1173,N_1171);
nor U1227 (N_1227,N_1194,N_1146);
and U1228 (N_1228,N_1185,N_1182);
nor U1229 (N_1229,N_1160,N_1197);
nor U1230 (N_1230,N_1153,N_1169);
nor U1231 (N_1231,N_1172,N_1191);
nor U1232 (N_1232,N_1145,N_1161);
nor U1233 (N_1233,N_1162,N_1175);
nor U1234 (N_1234,N_1171,N_1196);
nor U1235 (N_1235,N_1187,N_1198);
and U1236 (N_1236,N_1161,N_1191);
nor U1237 (N_1237,N_1166,N_1196);
and U1238 (N_1238,N_1152,N_1186);
nor U1239 (N_1239,N_1156,N_1183);
and U1240 (N_1240,N_1146,N_1196);
nor U1241 (N_1241,N_1170,N_1169);
nor U1242 (N_1242,N_1159,N_1199);
or U1243 (N_1243,N_1150,N_1194);
or U1244 (N_1244,N_1148,N_1187);
or U1245 (N_1245,N_1192,N_1187);
nand U1246 (N_1246,N_1145,N_1168);
nand U1247 (N_1247,N_1180,N_1154);
and U1248 (N_1248,N_1163,N_1188);
nand U1249 (N_1249,N_1159,N_1175);
nand U1250 (N_1250,N_1177,N_1196);
and U1251 (N_1251,N_1198,N_1163);
nand U1252 (N_1252,N_1168,N_1146);
nand U1253 (N_1253,N_1170,N_1184);
nor U1254 (N_1254,N_1181,N_1144);
or U1255 (N_1255,N_1168,N_1148);
nand U1256 (N_1256,N_1194,N_1141);
nand U1257 (N_1257,N_1196,N_1143);
nor U1258 (N_1258,N_1173,N_1166);
nand U1259 (N_1259,N_1184,N_1163);
nor U1260 (N_1260,N_1229,N_1230);
or U1261 (N_1261,N_1252,N_1245);
nand U1262 (N_1262,N_1207,N_1237);
and U1263 (N_1263,N_1223,N_1239);
and U1264 (N_1264,N_1201,N_1209);
nand U1265 (N_1265,N_1220,N_1203);
and U1266 (N_1266,N_1250,N_1249);
and U1267 (N_1267,N_1235,N_1225);
nor U1268 (N_1268,N_1242,N_1243);
nand U1269 (N_1269,N_1210,N_1231);
and U1270 (N_1270,N_1258,N_1246);
nor U1271 (N_1271,N_1253,N_1228);
nand U1272 (N_1272,N_1211,N_1219);
or U1273 (N_1273,N_1236,N_1257);
and U1274 (N_1274,N_1247,N_1254);
nand U1275 (N_1275,N_1200,N_1214);
nand U1276 (N_1276,N_1226,N_1208);
or U1277 (N_1277,N_1248,N_1202);
or U1278 (N_1278,N_1213,N_1204);
nor U1279 (N_1279,N_1234,N_1224);
and U1280 (N_1280,N_1218,N_1241);
nor U1281 (N_1281,N_1240,N_1215);
and U1282 (N_1282,N_1259,N_1212);
nor U1283 (N_1283,N_1206,N_1227);
and U1284 (N_1284,N_1251,N_1256);
nor U1285 (N_1285,N_1217,N_1205);
and U1286 (N_1286,N_1244,N_1238);
and U1287 (N_1287,N_1232,N_1216);
and U1288 (N_1288,N_1222,N_1255);
and U1289 (N_1289,N_1233,N_1221);
nand U1290 (N_1290,N_1230,N_1200);
or U1291 (N_1291,N_1253,N_1257);
nor U1292 (N_1292,N_1223,N_1247);
nand U1293 (N_1293,N_1211,N_1205);
and U1294 (N_1294,N_1231,N_1242);
and U1295 (N_1295,N_1253,N_1226);
nor U1296 (N_1296,N_1236,N_1224);
or U1297 (N_1297,N_1231,N_1253);
nor U1298 (N_1298,N_1205,N_1225);
nor U1299 (N_1299,N_1201,N_1236);
and U1300 (N_1300,N_1247,N_1233);
nor U1301 (N_1301,N_1250,N_1259);
or U1302 (N_1302,N_1246,N_1242);
and U1303 (N_1303,N_1223,N_1209);
or U1304 (N_1304,N_1231,N_1216);
and U1305 (N_1305,N_1248,N_1255);
or U1306 (N_1306,N_1245,N_1251);
nand U1307 (N_1307,N_1233,N_1206);
and U1308 (N_1308,N_1247,N_1207);
and U1309 (N_1309,N_1234,N_1205);
or U1310 (N_1310,N_1216,N_1246);
or U1311 (N_1311,N_1229,N_1259);
and U1312 (N_1312,N_1204,N_1207);
nor U1313 (N_1313,N_1231,N_1241);
or U1314 (N_1314,N_1232,N_1237);
and U1315 (N_1315,N_1207,N_1230);
nor U1316 (N_1316,N_1233,N_1220);
nand U1317 (N_1317,N_1257,N_1206);
or U1318 (N_1318,N_1232,N_1209);
or U1319 (N_1319,N_1200,N_1241);
or U1320 (N_1320,N_1310,N_1311);
nand U1321 (N_1321,N_1317,N_1290);
nand U1322 (N_1322,N_1295,N_1308);
and U1323 (N_1323,N_1287,N_1291);
and U1324 (N_1324,N_1284,N_1269);
nor U1325 (N_1325,N_1271,N_1283);
or U1326 (N_1326,N_1301,N_1260);
nor U1327 (N_1327,N_1270,N_1263);
nor U1328 (N_1328,N_1307,N_1305);
or U1329 (N_1329,N_1277,N_1304);
and U1330 (N_1330,N_1318,N_1265);
or U1331 (N_1331,N_1306,N_1285);
nor U1332 (N_1332,N_1275,N_1294);
nand U1333 (N_1333,N_1274,N_1273);
or U1334 (N_1334,N_1282,N_1268);
nand U1335 (N_1335,N_1312,N_1264);
and U1336 (N_1336,N_1276,N_1267);
or U1337 (N_1337,N_1313,N_1261);
xor U1338 (N_1338,N_1293,N_1302);
nor U1339 (N_1339,N_1309,N_1292);
and U1340 (N_1340,N_1288,N_1298);
or U1341 (N_1341,N_1319,N_1280);
and U1342 (N_1342,N_1303,N_1278);
nor U1343 (N_1343,N_1262,N_1316);
nand U1344 (N_1344,N_1266,N_1300);
nor U1345 (N_1345,N_1296,N_1279);
and U1346 (N_1346,N_1281,N_1297);
and U1347 (N_1347,N_1272,N_1299);
nand U1348 (N_1348,N_1286,N_1315);
nand U1349 (N_1349,N_1289,N_1314);
nand U1350 (N_1350,N_1309,N_1293);
and U1351 (N_1351,N_1270,N_1304);
and U1352 (N_1352,N_1270,N_1272);
nand U1353 (N_1353,N_1276,N_1277);
nand U1354 (N_1354,N_1260,N_1290);
nor U1355 (N_1355,N_1310,N_1269);
and U1356 (N_1356,N_1316,N_1269);
and U1357 (N_1357,N_1286,N_1287);
xor U1358 (N_1358,N_1268,N_1296);
nor U1359 (N_1359,N_1313,N_1288);
and U1360 (N_1360,N_1312,N_1271);
nand U1361 (N_1361,N_1316,N_1286);
and U1362 (N_1362,N_1319,N_1303);
nor U1363 (N_1363,N_1312,N_1262);
or U1364 (N_1364,N_1299,N_1303);
and U1365 (N_1365,N_1313,N_1287);
and U1366 (N_1366,N_1302,N_1313);
nand U1367 (N_1367,N_1297,N_1303);
nand U1368 (N_1368,N_1306,N_1265);
or U1369 (N_1369,N_1283,N_1287);
or U1370 (N_1370,N_1260,N_1319);
nand U1371 (N_1371,N_1310,N_1291);
nand U1372 (N_1372,N_1275,N_1268);
or U1373 (N_1373,N_1291,N_1297);
nor U1374 (N_1374,N_1278,N_1309);
and U1375 (N_1375,N_1278,N_1306);
and U1376 (N_1376,N_1304,N_1303);
or U1377 (N_1377,N_1262,N_1295);
nand U1378 (N_1378,N_1277,N_1297);
and U1379 (N_1379,N_1279,N_1262);
or U1380 (N_1380,N_1322,N_1363);
nand U1381 (N_1381,N_1324,N_1355);
and U1382 (N_1382,N_1369,N_1368);
nand U1383 (N_1383,N_1338,N_1336);
nor U1384 (N_1384,N_1323,N_1328);
nor U1385 (N_1385,N_1343,N_1345);
and U1386 (N_1386,N_1378,N_1358);
or U1387 (N_1387,N_1351,N_1367);
and U1388 (N_1388,N_1346,N_1337);
and U1389 (N_1389,N_1379,N_1362);
nor U1390 (N_1390,N_1370,N_1376);
nand U1391 (N_1391,N_1333,N_1347);
and U1392 (N_1392,N_1354,N_1342);
and U1393 (N_1393,N_1360,N_1357);
and U1394 (N_1394,N_1341,N_1352);
or U1395 (N_1395,N_1375,N_1332);
nand U1396 (N_1396,N_1356,N_1326);
nand U1397 (N_1397,N_1335,N_1373);
nand U1398 (N_1398,N_1359,N_1366);
nor U1399 (N_1399,N_1349,N_1321);
and U1400 (N_1400,N_1327,N_1320);
or U1401 (N_1401,N_1330,N_1325);
or U1402 (N_1402,N_1344,N_1329);
or U1403 (N_1403,N_1340,N_1348);
or U1404 (N_1404,N_1361,N_1350);
and U1405 (N_1405,N_1353,N_1339);
and U1406 (N_1406,N_1372,N_1331);
or U1407 (N_1407,N_1374,N_1371);
and U1408 (N_1408,N_1377,N_1365);
nand U1409 (N_1409,N_1364,N_1334);
nand U1410 (N_1410,N_1366,N_1320);
nand U1411 (N_1411,N_1321,N_1365);
and U1412 (N_1412,N_1323,N_1361);
nand U1413 (N_1413,N_1334,N_1321);
and U1414 (N_1414,N_1366,N_1333);
nor U1415 (N_1415,N_1337,N_1334);
and U1416 (N_1416,N_1379,N_1365);
nor U1417 (N_1417,N_1355,N_1339);
nand U1418 (N_1418,N_1350,N_1329);
nand U1419 (N_1419,N_1365,N_1331);
and U1420 (N_1420,N_1354,N_1327);
and U1421 (N_1421,N_1377,N_1321);
and U1422 (N_1422,N_1344,N_1320);
or U1423 (N_1423,N_1329,N_1356);
and U1424 (N_1424,N_1363,N_1379);
and U1425 (N_1425,N_1346,N_1351);
nand U1426 (N_1426,N_1330,N_1364);
or U1427 (N_1427,N_1339,N_1359);
or U1428 (N_1428,N_1377,N_1374);
nor U1429 (N_1429,N_1337,N_1378);
and U1430 (N_1430,N_1328,N_1354);
and U1431 (N_1431,N_1322,N_1335);
nor U1432 (N_1432,N_1325,N_1346);
nor U1433 (N_1433,N_1376,N_1366);
nand U1434 (N_1434,N_1325,N_1369);
or U1435 (N_1435,N_1350,N_1347);
or U1436 (N_1436,N_1347,N_1325);
and U1437 (N_1437,N_1323,N_1355);
or U1438 (N_1438,N_1372,N_1352);
and U1439 (N_1439,N_1359,N_1340);
nor U1440 (N_1440,N_1416,N_1435);
or U1441 (N_1441,N_1432,N_1422);
or U1442 (N_1442,N_1400,N_1402);
or U1443 (N_1443,N_1401,N_1388);
or U1444 (N_1444,N_1380,N_1409);
nand U1445 (N_1445,N_1398,N_1417);
nor U1446 (N_1446,N_1411,N_1433);
or U1447 (N_1447,N_1413,N_1412);
and U1448 (N_1448,N_1387,N_1389);
or U1449 (N_1449,N_1431,N_1426);
nand U1450 (N_1450,N_1390,N_1399);
nor U1451 (N_1451,N_1385,N_1428);
nand U1452 (N_1452,N_1434,N_1425);
nor U1453 (N_1453,N_1439,N_1421);
and U1454 (N_1454,N_1407,N_1386);
or U1455 (N_1455,N_1418,N_1414);
nor U1456 (N_1456,N_1429,N_1403);
nand U1457 (N_1457,N_1436,N_1423);
nand U1458 (N_1458,N_1381,N_1406);
nor U1459 (N_1459,N_1395,N_1438);
and U1460 (N_1460,N_1382,N_1393);
or U1461 (N_1461,N_1420,N_1427);
nor U1462 (N_1462,N_1408,N_1430);
and U1463 (N_1463,N_1391,N_1396);
and U1464 (N_1464,N_1397,N_1419);
nand U1465 (N_1465,N_1415,N_1392);
nor U1466 (N_1466,N_1410,N_1404);
nor U1467 (N_1467,N_1437,N_1383);
nand U1468 (N_1468,N_1424,N_1405);
and U1469 (N_1469,N_1394,N_1384);
nor U1470 (N_1470,N_1435,N_1438);
nand U1471 (N_1471,N_1396,N_1436);
and U1472 (N_1472,N_1405,N_1389);
and U1473 (N_1473,N_1381,N_1420);
and U1474 (N_1474,N_1408,N_1413);
nand U1475 (N_1475,N_1383,N_1411);
nand U1476 (N_1476,N_1401,N_1404);
and U1477 (N_1477,N_1406,N_1431);
or U1478 (N_1478,N_1430,N_1406);
nor U1479 (N_1479,N_1400,N_1394);
and U1480 (N_1480,N_1391,N_1425);
nor U1481 (N_1481,N_1428,N_1400);
nor U1482 (N_1482,N_1385,N_1422);
or U1483 (N_1483,N_1387,N_1422);
nor U1484 (N_1484,N_1386,N_1399);
nand U1485 (N_1485,N_1387,N_1432);
and U1486 (N_1486,N_1432,N_1389);
nor U1487 (N_1487,N_1396,N_1426);
nor U1488 (N_1488,N_1432,N_1420);
nor U1489 (N_1489,N_1382,N_1400);
and U1490 (N_1490,N_1401,N_1436);
nor U1491 (N_1491,N_1420,N_1423);
nor U1492 (N_1492,N_1430,N_1403);
nand U1493 (N_1493,N_1421,N_1404);
nand U1494 (N_1494,N_1418,N_1385);
nor U1495 (N_1495,N_1397,N_1387);
or U1496 (N_1496,N_1412,N_1438);
nor U1497 (N_1497,N_1437,N_1435);
and U1498 (N_1498,N_1437,N_1407);
nor U1499 (N_1499,N_1439,N_1400);
and U1500 (N_1500,N_1463,N_1475);
and U1501 (N_1501,N_1441,N_1481);
or U1502 (N_1502,N_1484,N_1461);
nor U1503 (N_1503,N_1486,N_1454);
or U1504 (N_1504,N_1449,N_1442);
or U1505 (N_1505,N_1452,N_1480);
or U1506 (N_1506,N_1467,N_1456);
xnor U1507 (N_1507,N_1466,N_1451);
and U1508 (N_1508,N_1457,N_1447);
or U1509 (N_1509,N_1478,N_1488);
and U1510 (N_1510,N_1464,N_1473);
or U1511 (N_1511,N_1477,N_1495);
nand U1512 (N_1512,N_1444,N_1446);
and U1513 (N_1513,N_1497,N_1453);
and U1514 (N_1514,N_1483,N_1470);
or U1515 (N_1515,N_1491,N_1455);
nand U1516 (N_1516,N_1487,N_1468);
nand U1517 (N_1517,N_1476,N_1458);
nand U1518 (N_1518,N_1440,N_1479);
or U1519 (N_1519,N_1498,N_1490);
and U1520 (N_1520,N_1462,N_1493);
and U1521 (N_1521,N_1448,N_1465);
and U1522 (N_1522,N_1485,N_1459);
nand U1523 (N_1523,N_1494,N_1445);
and U1524 (N_1524,N_1450,N_1496);
nand U1525 (N_1525,N_1443,N_1474);
or U1526 (N_1526,N_1469,N_1472);
or U1527 (N_1527,N_1489,N_1471);
nor U1528 (N_1528,N_1460,N_1482);
nand U1529 (N_1529,N_1492,N_1499);
and U1530 (N_1530,N_1481,N_1442);
and U1531 (N_1531,N_1497,N_1460);
nor U1532 (N_1532,N_1471,N_1461);
or U1533 (N_1533,N_1493,N_1494);
or U1534 (N_1534,N_1475,N_1464);
and U1535 (N_1535,N_1446,N_1477);
or U1536 (N_1536,N_1452,N_1496);
and U1537 (N_1537,N_1478,N_1461);
or U1538 (N_1538,N_1489,N_1449);
and U1539 (N_1539,N_1467,N_1462);
and U1540 (N_1540,N_1498,N_1479);
nor U1541 (N_1541,N_1484,N_1443);
nor U1542 (N_1542,N_1477,N_1454);
and U1543 (N_1543,N_1444,N_1469);
nor U1544 (N_1544,N_1493,N_1459);
nor U1545 (N_1545,N_1476,N_1487);
nand U1546 (N_1546,N_1485,N_1484);
nand U1547 (N_1547,N_1486,N_1452);
nor U1548 (N_1548,N_1448,N_1491);
and U1549 (N_1549,N_1482,N_1470);
or U1550 (N_1550,N_1456,N_1487);
and U1551 (N_1551,N_1487,N_1440);
and U1552 (N_1552,N_1446,N_1471);
and U1553 (N_1553,N_1440,N_1475);
and U1554 (N_1554,N_1453,N_1483);
and U1555 (N_1555,N_1482,N_1467);
nand U1556 (N_1556,N_1470,N_1475);
nor U1557 (N_1557,N_1491,N_1499);
and U1558 (N_1558,N_1468,N_1469);
nor U1559 (N_1559,N_1467,N_1458);
or U1560 (N_1560,N_1512,N_1546);
and U1561 (N_1561,N_1513,N_1532);
and U1562 (N_1562,N_1549,N_1539);
or U1563 (N_1563,N_1538,N_1509);
nand U1564 (N_1564,N_1518,N_1502);
and U1565 (N_1565,N_1519,N_1511);
and U1566 (N_1566,N_1529,N_1535);
or U1567 (N_1567,N_1533,N_1543);
and U1568 (N_1568,N_1517,N_1553);
or U1569 (N_1569,N_1527,N_1505);
nor U1570 (N_1570,N_1542,N_1540);
nand U1571 (N_1571,N_1537,N_1506);
or U1572 (N_1572,N_1516,N_1548);
or U1573 (N_1573,N_1515,N_1536);
nor U1574 (N_1574,N_1526,N_1558);
nor U1575 (N_1575,N_1555,N_1528);
nand U1576 (N_1576,N_1503,N_1547);
nor U1577 (N_1577,N_1504,N_1554);
and U1578 (N_1578,N_1508,N_1544);
or U1579 (N_1579,N_1510,N_1551);
nor U1580 (N_1580,N_1521,N_1514);
and U1581 (N_1581,N_1530,N_1522);
nand U1582 (N_1582,N_1556,N_1520);
nand U1583 (N_1583,N_1550,N_1500);
xnor U1584 (N_1584,N_1525,N_1507);
xnor U1585 (N_1585,N_1541,N_1545);
nand U1586 (N_1586,N_1534,N_1501);
and U1587 (N_1587,N_1531,N_1552);
nor U1588 (N_1588,N_1557,N_1559);
and U1589 (N_1589,N_1523,N_1524);
nor U1590 (N_1590,N_1530,N_1509);
or U1591 (N_1591,N_1535,N_1552);
or U1592 (N_1592,N_1507,N_1550);
nand U1593 (N_1593,N_1516,N_1538);
nand U1594 (N_1594,N_1538,N_1510);
nor U1595 (N_1595,N_1528,N_1530);
or U1596 (N_1596,N_1516,N_1532);
and U1597 (N_1597,N_1525,N_1500);
or U1598 (N_1598,N_1509,N_1537);
nor U1599 (N_1599,N_1553,N_1519);
and U1600 (N_1600,N_1515,N_1502);
nand U1601 (N_1601,N_1517,N_1500);
nand U1602 (N_1602,N_1543,N_1517);
and U1603 (N_1603,N_1527,N_1542);
and U1604 (N_1604,N_1558,N_1509);
nand U1605 (N_1605,N_1509,N_1541);
or U1606 (N_1606,N_1516,N_1528);
or U1607 (N_1607,N_1527,N_1526);
nand U1608 (N_1608,N_1540,N_1511);
and U1609 (N_1609,N_1556,N_1541);
and U1610 (N_1610,N_1558,N_1501);
nor U1611 (N_1611,N_1547,N_1538);
and U1612 (N_1612,N_1542,N_1537);
and U1613 (N_1613,N_1500,N_1549);
nor U1614 (N_1614,N_1557,N_1556);
nor U1615 (N_1615,N_1556,N_1538);
nand U1616 (N_1616,N_1503,N_1516);
and U1617 (N_1617,N_1507,N_1517);
nor U1618 (N_1618,N_1529,N_1519);
nand U1619 (N_1619,N_1501,N_1520);
or U1620 (N_1620,N_1609,N_1562);
and U1621 (N_1621,N_1587,N_1611);
and U1622 (N_1622,N_1576,N_1568);
nand U1623 (N_1623,N_1574,N_1612);
nor U1624 (N_1624,N_1580,N_1598);
nor U1625 (N_1625,N_1581,N_1599);
or U1626 (N_1626,N_1601,N_1583);
nand U1627 (N_1627,N_1584,N_1604);
and U1628 (N_1628,N_1573,N_1614);
nand U1629 (N_1629,N_1605,N_1610);
or U1630 (N_1630,N_1561,N_1592);
and U1631 (N_1631,N_1570,N_1607);
or U1632 (N_1632,N_1618,N_1596);
and U1633 (N_1633,N_1589,N_1560);
or U1634 (N_1634,N_1572,N_1571);
and U1635 (N_1635,N_1602,N_1575);
nand U1636 (N_1636,N_1585,N_1586);
nand U1637 (N_1637,N_1603,N_1564);
nand U1638 (N_1638,N_1577,N_1569);
or U1639 (N_1639,N_1619,N_1613);
nand U1640 (N_1640,N_1608,N_1600);
and U1641 (N_1641,N_1566,N_1595);
or U1642 (N_1642,N_1594,N_1615);
nand U1643 (N_1643,N_1593,N_1588);
or U1644 (N_1644,N_1590,N_1565);
and U1645 (N_1645,N_1567,N_1578);
nor U1646 (N_1646,N_1617,N_1597);
nand U1647 (N_1647,N_1563,N_1616);
or U1648 (N_1648,N_1579,N_1582);
and U1649 (N_1649,N_1591,N_1606);
nand U1650 (N_1650,N_1601,N_1567);
and U1651 (N_1651,N_1571,N_1598);
or U1652 (N_1652,N_1613,N_1615);
or U1653 (N_1653,N_1569,N_1618);
or U1654 (N_1654,N_1572,N_1619);
nand U1655 (N_1655,N_1575,N_1608);
nand U1656 (N_1656,N_1592,N_1596);
nor U1657 (N_1657,N_1595,N_1579);
nor U1658 (N_1658,N_1580,N_1575);
nor U1659 (N_1659,N_1583,N_1597);
or U1660 (N_1660,N_1587,N_1563);
and U1661 (N_1661,N_1565,N_1608);
or U1662 (N_1662,N_1613,N_1589);
or U1663 (N_1663,N_1575,N_1565);
nor U1664 (N_1664,N_1619,N_1602);
nand U1665 (N_1665,N_1571,N_1574);
nor U1666 (N_1666,N_1567,N_1599);
and U1667 (N_1667,N_1601,N_1590);
or U1668 (N_1668,N_1566,N_1564);
nand U1669 (N_1669,N_1578,N_1587);
or U1670 (N_1670,N_1582,N_1569);
or U1671 (N_1671,N_1582,N_1561);
or U1672 (N_1672,N_1603,N_1605);
or U1673 (N_1673,N_1582,N_1604);
nor U1674 (N_1674,N_1580,N_1612);
nor U1675 (N_1675,N_1613,N_1616);
nor U1676 (N_1676,N_1614,N_1615);
or U1677 (N_1677,N_1616,N_1581);
or U1678 (N_1678,N_1577,N_1595);
nor U1679 (N_1679,N_1575,N_1569);
or U1680 (N_1680,N_1671,N_1643);
or U1681 (N_1681,N_1629,N_1631);
nand U1682 (N_1682,N_1666,N_1673);
nand U1683 (N_1683,N_1641,N_1642);
or U1684 (N_1684,N_1645,N_1652);
nand U1685 (N_1685,N_1622,N_1636);
and U1686 (N_1686,N_1660,N_1635);
nand U1687 (N_1687,N_1656,N_1663);
nor U1688 (N_1688,N_1634,N_1640);
or U1689 (N_1689,N_1650,N_1632);
and U1690 (N_1690,N_1647,N_1651);
nor U1691 (N_1691,N_1628,N_1633);
or U1692 (N_1692,N_1675,N_1669);
nor U1693 (N_1693,N_1646,N_1658);
or U1694 (N_1694,N_1630,N_1626);
or U1695 (N_1695,N_1627,N_1657);
nor U1696 (N_1696,N_1649,N_1661);
nor U1697 (N_1697,N_1679,N_1672);
nand U1698 (N_1698,N_1620,N_1678);
or U1699 (N_1699,N_1667,N_1625);
and U1700 (N_1700,N_1639,N_1623);
or U1701 (N_1701,N_1624,N_1648);
nor U1702 (N_1702,N_1665,N_1662);
and U1703 (N_1703,N_1638,N_1659);
nor U1704 (N_1704,N_1670,N_1654);
nor U1705 (N_1705,N_1653,N_1668);
and U1706 (N_1706,N_1637,N_1644);
nand U1707 (N_1707,N_1674,N_1655);
or U1708 (N_1708,N_1664,N_1676);
and U1709 (N_1709,N_1621,N_1677);
and U1710 (N_1710,N_1666,N_1632);
or U1711 (N_1711,N_1647,N_1622);
nor U1712 (N_1712,N_1657,N_1639);
or U1713 (N_1713,N_1677,N_1627);
and U1714 (N_1714,N_1678,N_1645);
or U1715 (N_1715,N_1674,N_1630);
and U1716 (N_1716,N_1626,N_1622);
nand U1717 (N_1717,N_1628,N_1653);
nor U1718 (N_1718,N_1647,N_1648);
nor U1719 (N_1719,N_1672,N_1651);
nand U1720 (N_1720,N_1663,N_1631);
and U1721 (N_1721,N_1648,N_1667);
and U1722 (N_1722,N_1664,N_1644);
nor U1723 (N_1723,N_1669,N_1632);
and U1724 (N_1724,N_1630,N_1647);
or U1725 (N_1725,N_1631,N_1625);
nor U1726 (N_1726,N_1652,N_1664);
or U1727 (N_1727,N_1642,N_1639);
or U1728 (N_1728,N_1621,N_1667);
or U1729 (N_1729,N_1641,N_1631);
and U1730 (N_1730,N_1637,N_1620);
or U1731 (N_1731,N_1662,N_1638);
xor U1732 (N_1732,N_1667,N_1664);
nand U1733 (N_1733,N_1648,N_1662);
and U1734 (N_1734,N_1665,N_1655);
nand U1735 (N_1735,N_1653,N_1631);
or U1736 (N_1736,N_1641,N_1636);
nand U1737 (N_1737,N_1663,N_1632);
nor U1738 (N_1738,N_1620,N_1633);
nand U1739 (N_1739,N_1637,N_1658);
nor U1740 (N_1740,N_1726,N_1718);
and U1741 (N_1741,N_1722,N_1716);
nand U1742 (N_1742,N_1702,N_1706);
nor U1743 (N_1743,N_1703,N_1700);
nor U1744 (N_1744,N_1738,N_1701);
or U1745 (N_1745,N_1708,N_1737);
and U1746 (N_1746,N_1732,N_1705);
nand U1747 (N_1747,N_1683,N_1721);
or U1748 (N_1748,N_1724,N_1719);
and U1749 (N_1749,N_1727,N_1692);
nand U1750 (N_1750,N_1685,N_1689);
and U1751 (N_1751,N_1730,N_1707);
or U1752 (N_1752,N_1725,N_1690);
or U1753 (N_1753,N_1733,N_1687);
nand U1754 (N_1754,N_1688,N_1694);
or U1755 (N_1755,N_1680,N_1693);
nor U1756 (N_1756,N_1704,N_1739);
or U1757 (N_1757,N_1720,N_1717);
and U1758 (N_1758,N_1710,N_1736);
nand U1759 (N_1759,N_1686,N_1731);
or U1760 (N_1760,N_1691,N_1711);
or U1761 (N_1761,N_1735,N_1729);
and U1762 (N_1762,N_1698,N_1681);
nand U1763 (N_1763,N_1696,N_1712);
nor U1764 (N_1764,N_1682,N_1728);
and U1765 (N_1765,N_1697,N_1714);
nand U1766 (N_1766,N_1713,N_1699);
or U1767 (N_1767,N_1723,N_1734);
nand U1768 (N_1768,N_1684,N_1695);
nor U1769 (N_1769,N_1709,N_1715);
or U1770 (N_1770,N_1683,N_1706);
nand U1771 (N_1771,N_1715,N_1724);
or U1772 (N_1772,N_1737,N_1717);
and U1773 (N_1773,N_1686,N_1712);
and U1774 (N_1774,N_1733,N_1704);
or U1775 (N_1775,N_1717,N_1734);
or U1776 (N_1776,N_1682,N_1736);
nand U1777 (N_1777,N_1734,N_1711);
nand U1778 (N_1778,N_1727,N_1685);
nor U1779 (N_1779,N_1732,N_1712);
or U1780 (N_1780,N_1693,N_1690);
nor U1781 (N_1781,N_1688,N_1681);
or U1782 (N_1782,N_1712,N_1724);
and U1783 (N_1783,N_1736,N_1717);
and U1784 (N_1784,N_1734,N_1737);
or U1785 (N_1785,N_1684,N_1724);
nand U1786 (N_1786,N_1680,N_1710);
or U1787 (N_1787,N_1699,N_1711);
nand U1788 (N_1788,N_1688,N_1723);
nand U1789 (N_1789,N_1733,N_1693);
nand U1790 (N_1790,N_1735,N_1715);
nand U1791 (N_1791,N_1717,N_1722);
or U1792 (N_1792,N_1699,N_1728);
nand U1793 (N_1793,N_1704,N_1710);
and U1794 (N_1794,N_1712,N_1685);
or U1795 (N_1795,N_1683,N_1704);
nor U1796 (N_1796,N_1699,N_1708);
xor U1797 (N_1797,N_1713,N_1684);
nand U1798 (N_1798,N_1694,N_1724);
or U1799 (N_1799,N_1690,N_1726);
nor U1800 (N_1800,N_1746,N_1771);
or U1801 (N_1801,N_1792,N_1748);
xor U1802 (N_1802,N_1768,N_1752);
and U1803 (N_1803,N_1776,N_1744);
nor U1804 (N_1804,N_1755,N_1761);
nand U1805 (N_1805,N_1757,N_1789);
and U1806 (N_1806,N_1753,N_1749);
nor U1807 (N_1807,N_1786,N_1743);
nand U1808 (N_1808,N_1772,N_1742);
nand U1809 (N_1809,N_1783,N_1788);
nand U1810 (N_1810,N_1762,N_1796);
nand U1811 (N_1811,N_1740,N_1780);
nand U1812 (N_1812,N_1774,N_1764);
and U1813 (N_1813,N_1777,N_1765);
nand U1814 (N_1814,N_1790,N_1756);
or U1815 (N_1815,N_1763,N_1794);
xor U1816 (N_1816,N_1787,N_1745);
and U1817 (N_1817,N_1751,N_1747);
or U1818 (N_1818,N_1797,N_1795);
and U1819 (N_1819,N_1760,N_1769);
nor U1820 (N_1820,N_1785,N_1779);
nand U1821 (N_1821,N_1798,N_1793);
nor U1822 (N_1822,N_1781,N_1773);
nor U1823 (N_1823,N_1758,N_1770);
or U1824 (N_1824,N_1784,N_1754);
nand U1825 (N_1825,N_1778,N_1759);
or U1826 (N_1826,N_1750,N_1766);
nor U1827 (N_1827,N_1799,N_1791);
or U1828 (N_1828,N_1782,N_1775);
and U1829 (N_1829,N_1767,N_1741);
nor U1830 (N_1830,N_1762,N_1781);
or U1831 (N_1831,N_1762,N_1740);
nor U1832 (N_1832,N_1774,N_1770);
nor U1833 (N_1833,N_1795,N_1757);
and U1834 (N_1834,N_1785,N_1752);
and U1835 (N_1835,N_1766,N_1761);
nor U1836 (N_1836,N_1756,N_1747);
nor U1837 (N_1837,N_1773,N_1785);
nand U1838 (N_1838,N_1760,N_1779);
nand U1839 (N_1839,N_1762,N_1779);
nor U1840 (N_1840,N_1740,N_1752);
and U1841 (N_1841,N_1761,N_1773);
nor U1842 (N_1842,N_1794,N_1748);
and U1843 (N_1843,N_1791,N_1745);
and U1844 (N_1844,N_1743,N_1773);
nand U1845 (N_1845,N_1768,N_1788);
nor U1846 (N_1846,N_1776,N_1795);
nor U1847 (N_1847,N_1769,N_1798);
and U1848 (N_1848,N_1747,N_1769);
nand U1849 (N_1849,N_1780,N_1790);
or U1850 (N_1850,N_1773,N_1766);
or U1851 (N_1851,N_1774,N_1785);
or U1852 (N_1852,N_1755,N_1747);
or U1853 (N_1853,N_1756,N_1743);
nand U1854 (N_1854,N_1765,N_1791);
or U1855 (N_1855,N_1794,N_1755);
or U1856 (N_1856,N_1779,N_1787);
nand U1857 (N_1857,N_1756,N_1759);
and U1858 (N_1858,N_1752,N_1796);
nor U1859 (N_1859,N_1769,N_1752);
nand U1860 (N_1860,N_1844,N_1810);
or U1861 (N_1861,N_1829,N_1811);
or U1862 (N_1862,N_1822,N_1823);
nand U1863 (N_1863,N_1859,N_1819);
and U1864 (N_1864,N_1838,N_1849);
nor U1865 (N_1865,N_1853,N_1852);
nand U1866 (N_1866,N_1833,N_1814);
nor U1867 (N_1867,N_1827,N_1834);
nor U1868 (N_1868,N_1820,N_1825);
and U1869 (N_1869,N_1803,N_1857);
nor U1870 (N_1870,N_1809,N_1841);
nor U1871 (N_1871,N_1821,N_1808);
nor U1872 (N_1872,N_1824,N_1845);
nand U1873 (N_1873,N_1804,N_1842);
nand U1874 (N_1874,N_1826,N_1816);
nor U1875 (N_1875,N_1805,N_1830);
nand U1876 (N_1876,N_1847,N_1817);
nor U1877 (N_1877,N_1851,N_1854);
or U1878 (N_1878,N_1836,N_1858);
or U1879 (N_1879,N_1839,N_1807);
or U1880 (N_1880,N_1855,N_1806);
or U1881 (N_1881,N_1828,N_1815);
or U1882 (N_1882,N_1800,N_1813);
or U1883 (N_1883,N_1848,N_1831);
nor U1884 (N_1884,N_1801,N_1837);
nor U1885 (N_1885,N_1832,N_1840);
and U1886 (N_1886,N_1818,N_1843);
nand U1887 (N_1887,N_1835,N_1850);
nor U1888 (N_1888,N_1802,N_1846);
or U1889 (N_1889,N_1856,N_1812);
xor U1890 (N_1890,N_1841,N_1817);
nor U1891 (N_1891,N_1809,N_1807);
nor U1892 (N_1892,N_1825,N_1843);
nor U1893 (N_1893,N_1849,N_1810);
nand U1894 (N_1894,N_1834,N_1859);
nor U1895 (N_1895,N_1836,N_1847);
and U1896 (N_1896,N_1847,N_1806);
or U1897 (N_1897,N_1814,N_1821);
nand U1898 (N_1898,N_1812,N_1811);
nor U1899 (N_1899,N_1848,N_1833);
or U1900 (N_1900,N_1842,N_1857);
nand U1901 (N_1901,N_1832,N_1842);
nor U1902 (N_1902,N_1831,N_1836);
nand U1903 (N_1903,N_1856,N_1815);
nand U1904 (N_1904,N_1813,N_1801);
nor U1905 (N_1905,N_1801,N_1807);
nand U1906 (N_1906,N_1815,N_1849);
nand U1907 (N_1907,N_1807,N_1854);
and U1908 (N_1908,N_1824,N_1837);
nand U1909 (N_1909,N_1859,N_1849);
nor U1910 (N_1910,N_1812,N_1857);
and U1911 (N_1911,N_1851,N_1857);
or U1912 (N_1912,N_1806,N_1827);
or U1913 (N_1913,N_1811,N_1853);
or U1914 (N_1914,N_1806,N_1835);
nor U1915 (N_1915,N_1846,N_1822);
xnor U1916 (N_1916,N_1842,N_1835);
and U1917 (N_1917,N_1827,N_1836);
or U1918 (N_1918,N_1819,N_1840);
nand U1919 (N_1919,N_1813,N_1814);
nor U1920 (N_1920,N_1879,N_1873);
and U1921 (N_1921,N_1910,N_1866);
nor U1922 (N_1922,N_1894,N_1875);
or U1923 (N_1923,N_1895,N_1912);
and U1924 (N_1924,N_1898,N_1911);
nor U1925 (N_1925,N_1908,N_1913);
nand U1926 (N_1926,N_1904,N_1869);
and U1927 (N_1927,N_1881,N_1878);
nor U1928 (N_1928,N_1872,N_1882);
and U1929 (N_1929,N_1861,N_1897);
nor U1930 (N_1930,N_1893,N_1909);
and U1931 (N_1931,N_1884,N_1890);
or U1932 (N_1932,N_1919,N_1864);
nand U1933 (N_1933,N_1862,N_1886);
or U1934 (N_1934,N_1860,N_1870);
and U1935 (N_1935,N_1865,N_1896);
nand U1936 (N_1936,N_1868,N_1880);
or U1937 (N_1937,N_1916,N_1907);
xnor U1938 (N_1938,N_1891,N_1887);
and U1939 (N_1939,N_1863,N_1877);
or U1940 (N_1940,N_1889,N_1915);
xnor U1941 (N_1941,N_1903,N_1885);
and U1942 (N_1942,N_1899,N_1905);
or U1943 (N_1943,N_1917,N_1876);
or U1944 (N_1944,N_1871,N_1892);
or U1945 (N_1945,N_1900,N_1867);
or U1946 (N_1946,N_1883,N_1914);
nor U1947 (N_1947,N_1888,N_1906);
or U1948 (N_1948,N_1874,N_1918);
nor U1949 (N_1949,N_1901,N_1902);
nor U1950 (N_1950,N_1866,N_1861);
or U1951 (N_1951,N_1907,N_1901);
nand U1952 (N_1952,N_1917,N_1884);
nor U1953 (N_1953,N_1873,N_1894);
nor U1954 (N_1954,N_1917,N_1912);
and U1955 (N_1955,N_1913,N_1899);
or U1956 (N_1956,N_1864,N_1870);
nor U1957 (N_1957,N_1872,N_1866);
and U1958 (N_1958,N_1890,N_1894);
and U1959 (N_1959,N_1914,N_1919);
or U1960 (N_1960,N_1870,N_1895);
nand U1961 (N_1961,N_1861,N_1914);
nand U1962 (N_1962,N_1902,N_1866);
and U1963 (N_1963,N_1875,N_1878);
and U1964 (N_1964,N_1892,N_1901);
or U1965 (N_1965,N_1884,N_1899);
nor U1966 (N_1966,N_1887,N_1883);
and U1967 (N_1967,N_1903,N_1867);
or U1968 (N_1968,N_1888,N_1862);
nand U1969 (N_1969,N_1903,N_1878);
nor U1970 (N_1970,N_1898,N_1915);
and U1971 (N_1971,N_1870,N_1883);
and U1972 (N_1972,N_1896,N_1870);
nand U1973 (N_1973,N_1895,N_1880);
nor U1974 (N_1974,N_1881,N_1898);
nand U1975 (N_1975,N_1873,N_1868);
nand U1976 (N_1976,N_1897,N_1862);
nor U1977 (N_1977,N_1916,N_1891);
or U1978 (N_1978,N_1889,N_1891);
nor U1979 (N_1979,N_1913,N_1904);
nand U1980 (N_1980,N_1949,N_1936);
nor U1981 (N_1981,N_1927,N_1940);
and U1982 (N_1982,N_1941,N_1977);
nor U1983 (N_1983,N_1966,N_1968);
or U1984 (N_1984,N_1925,N_1931);
and U1985 (N_1985,N_1972,N_1920);
nor U1986 (N_1986,N_1923,N_1951);
and U1987 (N_1987,N_1950,N_1969);
and U1988 (N_1988,N_1971,N_1976);
or U1989 (N_1989,N_1922,N_1928);
nand U1990 (N_1990,N_1960,N_1939);
or U1991 (N_1991,N_1929,N_1934);
and U1992 (N_1992,N_1963,N_1942);
or U1993 (N_1993,N_1945,N_1978);
and U1994 (N_1994,N_1979,N_1938);
nand U1995 (N_1995,N_1921,N_1959);
and U1996 (N_1996,N_1955,N_1961);
nand U1997 (N_1997,N_1962,N_1935);
nor U1998 (N_1998,N_1943,N_1933);
nand U1999 (N_1999,N_1967,N_1953);
nor U2000 (N_2000,N_1944,N_1930);
or U2001 (N_2001,N_1954,N_1958);
nand U2002 (N_2002,N_1975,N_1947);
nor U2003 (N_2003,N_1957,N_1924);
nor U2004 (N_2004,N_1946,N_1970);
and U2005 (N_2005,N_1952,N_1932);
xor U2006 (N_2006,N_1937,N_1973);
and U2007 (N_2007,N_1964,N_1965);
or U2008 (N_2008,N_1974,N_1926);
or U2009 (N_2009,N_1956,N_1948);
nand U2010 (N_2010,N_1937,N_1941);
nand U2011 (N_2011,N_1940,N_1947);
nor U2012 (N_2012,N_1946,N_1962);
or U2013 (N_2013,N_1944,N_1966);
nor U2014 (N_2014,N_1929,N_1943);
nand U2015 (N_2015,N_1947,N_1923);
nor U2016 (N_2016,N_1925,N_1932);
nor U2017 (N_2017,N_1975,N_1965);
nand U2018 (N_2018,N_1954,N_1976);
nand U2019 (N_2019,N_1948,N_1978);
nor U2020 (N_2020,N_1970,N_1965);
or U2021 (N_2021,N_1922,N_1939);
nor U2022 (N_2022,N_1961,N_1965);
and U2023 (N_2023,N_1951,N_1932);
nand U2024 (N_2024,N_1928,N_1937);
nor U2025 (N_2025,N_1940,N_1952);
xor U2026 (N_2026,N_1964,N_1950);
nand U2027 (N_2027,N_1928,N_1975);
and U2028 (N_2028,N_1971,N_1921);
or U2029 (N_2029,N_1931,N_1948);
or U2030 (N_2030,N_1972,N_1977);
or U2031 (N_2031,N_1932,N_1924);
nand U2032 (N_2032,N_1962,N_1967);
and U2033 (N_2033,N_1925,N_1938);
or U2034 (N_2034,N_1960,N_1959);
nor U2035 (N_2035,N_1941,N_1942);
nor U2036 (N_2036,N_1921,N_1973);
nand U2037 (N_2037,N_1975,N_1929);
nor U2038 (N_2038,N_1927,N_1928);
nand U2039 (N_2039,N_1935,N_1925);
nor U2040 (N_2040,N_2011,N_1992);
and U2041 (N_2041,N_1994,N_1987);
nor U2042 (N_2042,N_2017,N_2034);
xor U2043 (N_2043,N_2036,N_2018);
nor U2044 (N_2044,N_1985,N_2027);
nor U2045 (N_2045,N_2037,N_1986);
nand U2046 (N_2046,N_1997,N_2029);
nand U2047 (N_2047,N_1983,N_2002);
or U2048 (N_2048,N_2028,N_2009);
xnor U2049 (N_2049,N_1993,N_2025);
nor U2050 (N_2050,N_1999,N_2016);
and U2051 (N_2051,N_2035,N_2022);
nor U2052 (N_2052,N_2010,N_2039);
nand U2053 (N_2053,N_2021,N_2031);
and U2054 (N_2054,N_2008,N_1990);
or U2055 (N_2055,N_2013,N_2001);
or U2056 (N_2056,N_2032,N_2000);
or U2057 (N_2057,N_2020,N_1989);
nor U2058 (N_2058,N_2026,N_2023);
nand U2059 (N_2059,N_1995,N_1980);
nor U2060 (N_2060,N_2007,N_2006);
nor U2061 (N_2061,N_1988,N_1996);
and U2062 (N_2062,N_2012,N_2014);
or U2063 (N_2063,N_2038,N_2015);
and U2064 (N_2064,N_2003,N_2030);
nor U2065 (N_2065,N_1998,N_2019);
and U2066 (N_2066,N_2005,N_2024);
and U2067 (N_2067,N_2004,N_1991);
and U2068 (N_2068,N_2033,N_1981);
and U2069 (N_2069,N_1984,N_1982);
nor U2070 (N_2070,N_2035,N_1998);
nor U2071 (N_2071,N_2002,N_2008);
nand U2072 (N_2072,N_2020,N_2033);
and U2073 (N_2073,N_2002,N_2004);
and U2074 (N_2074,N_2006,N_2038);
nor U2075 (N_2075,N_1981,N_2031);
and U2076 (N_2076,N_2005,N_1995);
nor U2077 (N_2077,N_1991,N_2008);
and U2078 (N_2078,N_2026,N_2027);
and U2079 (N_2079,N_2007,N_2000);
nor U2080 (N_2080,N_2013,N_2022);
nand U2081 (N_2081,N_2001,N_1999);
and U2082 (N_2082,N_2027,N_1991);
or U2083 (N_2083,N_2036,N_1999);
and U2084 (N_2084,N_1988,N_1987);
nor U2085 (N_2085,N_2007,N_2026);
and U2086 (N_2086,N_2007,N_2011);
and U2087 (N_2087,N_2001,N_2006);
and U2088 (N_2088,N_2028,N_1980);
nand U2089 (N_2089,N_1980,N_1981);
and U2090 (N_2090,N_2016,N_1980);
nand U2091 (N_2091,N_2006,N_2030);
nand U2092 (N_2092,N_1995,N_1984);
nand U2093 (N_2093,N_2002,N_2025);
and U2094 (N_2094,N_2017,N_1986);
or U2095 (N_2095,N_2019,N_1981);
and U2096 (N_2096,N_1996,N_2005);
nand U2097 (N_2097,N_2016,N_2023);
nand U2098 (N_2098,N_2023,N_2010);
nor U2099 (N_2099,N_2008,N_2016);
nand U2100 (N_2100,N_2090,N_2059);
or U2101 (N_2101,N_2089,N_2071);
nand U2102 (N_2102,N_2062,N_2096);
nand U2103 (N_2103,N_2078,N_2079);
and U2104 (N_2104,N_2040,N_2060);
and U2105 (N_2105,N_2048,N_2054);
nor U2106 (N_2106,N_2043,N_2064);
and U2107 (N_2107,N_2063,N_2068);
and U2108 (N_2108,N_2098,N_2076);
nand U2109 (N_2109,N_2044,N_2087);
nand U2110 (N_2110,N_2075,N_2050);
and U2111 (N_2111,N_2082,N_2070);
nor U2112 (N_2112,N_2073,N_2099);
nor U2113 (N_2113,N_2080,N_2066);
and U2114 (N_2114,N_2041,N_2086);
nand U2115 (N_2115,N_2052,N_2053);
nand U2116 (N_2116,N_2077,N_2045);
nor U2117 (N_2117,N_2092,N_2097);
nor U2118 (N_2118,N_2056,N_2042);
nand U2119 (N_2119,N_2083,N_2046);
or U2120 (N_2120,N_2095,N_2081);
nand U2121 (N_2121,N_2093,N_2055);
or U2122 (N_2122,N_2049,N_2084);
and U2123 (N_2123,N_2072,N_2047);
nand U2124 (N_2124,N_2067,N_2091);
nand U2125 (N_2125,N_2061,N_2065);
nand U2126 (N_2126,N_2074,N_2088);
nand U2127 (N_2127,N_2057,N_2094);
nor U2128 (N_2128,N_2085,N_2069);
or U2129 (N_2129,N_2051,N_2058);
and U2130 (N_2130,N_2043,N_2082);
and U2131 (N_2131,N_2096,N_2069);
nor U2132 (N_2132,N_2086,N_2079);
and U2133 (N_2133,N_2049,N_2096);
or U2134 (N_2134,N_2065,N_2085);
nand U2135 (N_2135,N_2085,N_2067);
and U2136 (N_2136,N_2047,N_2051);
or U2137 (N_2137,N_2090,N_2043);
or U2138 (N_2138,N_2078,N_2055);
and U2139 (N_2139,N_2048,N_2096);
nand U2140 (N_2140,N_2084,N_2063);
or U2141 (N_2141,N_2090,N_2056);
nand U2142 (N_2142,N_2073,N_2092);
nor U2143 (N_2143,N_2052,N_2040);
nor U2144 (N_2144,N_2048,N_2094);
and U2145 (N_2145,N_2084,N_2055);
nand U2146 (N_2146,N_2058,N_2070);
or U2147 (N_2147,N_2071,N_2088);
nor U2148 (N_2148,N_2054,N_2061);
nand U2149 (N_2149,N_2066,N_2078);
or U2150 (N_2150,N_2076,N_2084);
nand U2151 (N_2151,N_2042,N_2066);
or U2152 (N_2152,N_2044,N_2096);
and U2153 (N_2153,N_2048,N_2077);
nor U2154 (N_2154,N_2042,N_2043);
nand U2155 (N_2155,N_2040,N_2054);
nor U2156 (N_2156,N_2089,N_2068);
and U2157 (N_2157,N_2081,N_2048);
nand U2158 (N_2158,N_2056,N_2069);
and U2159 (N_2159,N_2050,N_2046);
and U2160 (N_2160,N_2146,N_2124);
nor U2161 (N_2161,N_2150,N_2102);
nor U2162 (N_2162,N_2105,N_2145);
or U2163 (N_2163,N_2122,N_2114);
or U2164 (N_2164,N_2117,N_2107);
or U2165 (N_2165,N_2101,N_2147);
or U2166 (N_2166,N_2138,N_2137);
nor U2167 (N_2167,N_2136,N_2115);
nor U2168 (N_2168,N_2152,N_2106);
or U2169 (N_2169,N_2156,N_2135);
or U2170 (N_2170,N_2143,N_2148);
nor U2171 (N_2171,N_2155,N_2144);
nor U2172 (N_2172,N_2140,N_2131);
nand U2173 (N_2173,N_2125,N_2153);
and U2174 (N_2174,N_2110,N_2134);
nand U2175 (N_2175,N_2128,N_2100);
and U2176 (N_2176,N_2113,N_2149);
nand U2177 (N_2177,N_2103,N_2139);
nand U2178 (N_2178,N_2151,N_2120);
and U2179 (N_2179,N_2112,N_2141);
nand U2180 (N_2180,N_2121,N_2158);
and U2181 (N_2181,N_2119,N_2132);
nor U2182 (N_2182,N_2104,N_2157);
nor U2183 (N_2183,N_2116,N_2127);
nor U2184 (N_2184,N_2109,N_2123);
nor U2185 (N_2185,N_2118,N_2130);
nand U2186 (N_2186,N_2108,N_2154);
or U2187 (N_2187,N_2129,N_2133);
nand U2188 (N_2188,N_2142,N_2126);
nand U2189 (N_2189,N_2159,N_2111);
nor U2190 (N_2190,N_2157,N_2135);
xor U2191 (N_2191,N_2113,N_2140);
nand U2192 (N_2192,N_2151,N_2111);
and U2193 (N_2193,N_2106,N_2145);
and U2194 (N_2194,N_2125,N_2100);
and U2195 (N_2195,N_2152,N_2145);
or U2196 (N_2196,N_2108,N_2104);
nand U2197 (N_2197,N_2144,N_2116);
or U2198 (N_2198,N_2150,N_2148);
nand U2199 (N_2199,N_2108,N_2135);
and U2200 (N_2200,N_2142,N_2155);
nand U2201 (N_2201,N_2107,N_2114);
nand U2202 (N_2202,N_2111,N_2116);
or U2203 (N_2203,N_2109,N_2114);
and U2204 (N_2204,N_2105,N_2112);
and U2205 (N_2205,N_2136,N_2156);
nand U2206 (N_2206,N_2128,N_2153);
and U2207 (N_2207,N_2130,N_2132);
nor U2208 (N_2208,N_2102,N_2151);
nor U2209 (N_2209,N_2149,N_2154);
nand U2210 (N_2210,N_2128,N_2151);
or U2211 (N_2211,N_2157,N_2131);
nand U2212 (N_2212,N_2147,N_2104);
and U2213 (N_2213,N_2159,N_2123);
nand U2214 (N_2214,N_2109,N_2103);
xor U2215 (N_2215,N_2137,N_2149);
nor U2216 (N_2216,N_2115,N_2150);
and U2217 (N_2217,N_2110,N_2113);
and U2218 (N_2218,N_2124,N_2140);
or U2219 (N_2219,N_2105,N_2123);
or U2220 (N_2220,N_2194,N_2195);
nor U2221 (N_2221,N_2204,N_2167);
or U2222 (N_2222,N_2180,N_2171);
nor U2223 (N_2223,N_2212,N_2187);
and U2224 (N_2224,N_2176,N_2218);
nand U2225 (N_2225,N_2188,N_2183);
nor U2226 (N_2226,N_2217,N_2196);
and U2227 (N_2227,N_2170,N_2213);
nand U2228 (N_2228,N_2162,N_2173);
and U2229 (N_2229,N_2179,N_2185);
nor U2230 (N_2230,N_2165,N_2160);
nor U2231 (N_2231,N_2178,N_2197);
and U2232 (N_2232,N_2192,N_2163);
nor U2233 (N_2233,N_2209,N_2168);
or U2234 (N_2234,N_2198,N_2199);
or U2235 (N_2235,N_2206,N_2174);
nand U2236 (N_2236,N_2175,N_2191);
nand U2237 (N_2237,N_2169,N_2166);
xor U2238 (N_2238,N_2203,N_2193);
nor U2239 (N_2239,N_2181,N_2207);
and U2240 (N_2240,N_2210,N_2216);
or U2241 (N_2241,N_2189,N_2172);
or U2242 (N_2242,N_2219,N_2200);
nor U2243 (N_2243,N_2211,N_2202);
or U2244 (N_2244,N_2214,N_2161);
and U2245 (N_2245,N_2182,N_2186);
nand U2246 (N_2246,N_2201,N_2177);
nor U2247 (N_2247,N_2208,N_2215);
or U2248 (N_2248,N_2184,N_2205);
nor U2249 (N_2249,N_2190,N_2164);
or U2250 (N_2250,N_2199,N_2170);
and U2251 (N_2251,N_2208,N_2193);
or U2252 (N_2252,N_2180,N_2213);
and U2253 (N_2253,N_2219,N_2197);
and U2254 (N_2254,N_2174,N_2171);
and U2255 (N_2255,N_2210,N_2200);
and U2256 (N_2256,N_2185,N_2166);
or U2257 (N_2257,N_2189,N_2175);
and U2258 (N_2258,N_2218,N_2212);
nand U2259 (N_2259,N_2163,N_2193);
nand U2260 (N_2260,N_2180,N_2218);
nor U2261 (N_2261,N_2161,N_2186);
and U2262 (N_2262,N_2178,N_2180);
and U2263 (N_2263,N_2197,N_2216);
or U2264 (N_2264,N_2163,N_2164);
or U2265 (N_2265,N_2170,N_2210);
nor U2266 (N_2266,N_2168,N_2199);
nor U2267 (N_2267,N_2170,N_2177);
or U2268 (N_2268,N_2214,N_2211);
nor U2269 (N_2269,N_2162,N_2214);
nor U2270 (N_2270,N_2213,N_2190);
or U2271 (N_2271,N_2173,N_2217);
nor U2272 (N_2272,N_2174,N_2166);
nor U2273 (N_2273,N_2201,N_2173);
nand U2274 (N_2274,N_2210,N_2162);
and U2275 (N_2275,N_2160,N_2205);
or U2276 (N_2276,N_2188,N_2206);
nand U2277 (N_2277,N_2209,N_2186);
nor U2278 (N_2278,N_2211,N_2198);
nor U2279 (N_2279,N_2215,N_2164);
and U2280 (N_2280,N_2267,N_2263);
nand U2281 (N_2281,N_2225,N_2253);
nor U2282 (N_2282,N_2241,N_2239);
or U2283 (N_2283,N_2255,N_2258);
nor U2284 (N_2284,N_2251,N_2270);
or U2285 (N_2285,N_2240,N_2268);
and U2286 (N_2286,N_2262,N_2274);
nand U2287 (N_2287,N_2221,N_2246);
and U2288 (N_2288,N_2232,N_2271);
nor U2289 (N_2289,N_2254,N_2250);
or U2290 (N_2290,N_2257,N_2234);
and U2291 (N_2291,N_2272,N_2222);
nor U2292 (N_2292,N_2275,N_2244);
or U2293 (N_2293,N_2278,N_2242);
and U2294 (N_2294,N_2220,N_2248);
nor U2295 (N_2295,N_2259,N_2233);
nand U2296 (N_2296,N_2264,N_2235);
nor U2297 (N_2297,N_2252,N_2269);
nand U2298 (N_2298,N_2277,N_2226);
or U2299 (N_2299,N_2231,N_2227);
and U2300 (N_2300,N_2228,N_2230);
nand U2301 (N_2301,N_2265,N_2276);
and U2302 (N_2302,N_2224,N_2279);
nor U2303 (N_2303,N_2243,N_2249);
and U2304 (N_2304,N_2236,N_2245);
or U2305 (N_2305,N_2260,N_2229);
nand U2306 (N_2306,N_2266,N_2273);
nand U2307 (N_2307,N_2238,N_2247);
and U2308 (N_2308,N_2256,N_2223);
and U2309 (N_2309,N_2261,N_2237);
nor U2310 (N_2310,N_2236,N_2242);
nand U2311 (N_2311,N_2260,N_2246);
or U2312 (N_2312,N_2255,N_2225);
or U2313 (N_2313,N_2222,N_2228);
and U2314 (N_2314,N_2262,N_2221);
and U2315 (N_2315,N_2267,N_2231);
and U2316 (N_2316,N_2223,N_2254);
nand U2317 (N_2317,N_2226,N_2262);
or U2318 (N_2318,N_2259,N_2272);
or U2319 (N_2319,N_2223,N_2271);
nand U2320 (N_2320,N_2241,N_2268);
nor U2321 (N_2321,N_2249,N_2262);
and U2322 (N_2322,N_2249,N_2270);
nor U2323 (N_2323,N_2263,N_2227);
or U2324 (N_2324,N_2247,N_2257);
or U2325 (N_2325,N_2241,N_2261);
or U2326 (N_2326,N_2230,N_2270);
and U2327 (N_2327,N_2278,N_2269);
and U2328 (N_2328,N_2232,N_2258);
nor U2329 (N_2329,N_2240,N_2226);
nor U2330 (N_2330,N_2230,N_2248);
or U2331 (N_2331,N_2235,N_2254);
nand U2332 (N_2332,N_2266,N_2228);
and U2333 (N_2333,N_2273,N_2261);
or U2334 (N_2334,N_2240,N_2251);
or U2335 (N_2335,N_2246,N_2264);
nor U2336 (N_2336,N_2277,N_2249);
or U2337 (N_2337,N_2244,N_2242);
or U2338 (N_2338,N_2246,N_2240);
xor U2339 (N_2339,N_2254,N_2229);
and U2340 (N_2340,N_2305,N_2334);
nand U2341 (N_2341,N_2288,N_2335);
or U2342 (N_2342,N_2325,N_2287);
and U2343 (N_2343,N_2326,N_2280);
and U2344 (N_2344,N_2285,N_2301);
or U2345 (N_2345,N_2327,N_2282);
nor U2346 (N_2346,N_2291,N_2286);
and U2347 (N_2347,N_2281,N_2317);
and U2348 (N_2348,N_2302,N_2309);
nor U2349 (N_2349,N_2292,N_2320);
or U2350 (N_2350,N_2328,N_2306);
nor U2351 (N_2351,N_2300,N_2310);
or U2352 (N_2352,N_2294,N_2338);
nand U2353 (N_2353,N_2313,N_2331);
nor U2354 (N_2354,N_2299,N_2339);
nor U2355 (N_2355,N_2304,N_2314);
nand U2356 (N_2356,N_2312,N_2315);
or U2357 (N_2357,N_2308,N_2295);
and U2358 (N_2358,N_2293,N_2307);
and U2359 (N_2359,N_2283,N_2322);
and U2360 (N_2360,N_2316,N_2298);
or U2361 (N_2361,N_2336,N_2337);
or U2362 (N_2362,N_2311,N_2289);
or U2363 (N_2363,N_2324,N_2303);
nand U2364 (N_2364,N_2318,N_2290);
and U2365 (N_2365,N_2330,N_2297);
nor U2366 (N_2366,N_2296,N_2329);
or U2367 (N_2367,N_2284,N_2323);
nand U2368 (N_2368,N_2332,N_2333);
xnor U2369 (N_2369,N_2319,N_2321);
or U2370 (N_2370,N_2333,N_2318);
nor U2371 (N_2371,N_2324,N_2287);
and U2372 (N_2372,N_2284,N_2295);
and U2373 (N_2373,N_2288,N_2302);
or U2374 (N_2374,N_2326,N_2337);
nor U2375 (N_2375,N_2312,N_2306);
nand U2376 (N_2376,N_2292,N_2323);
and U2377 (N_2377,N_2299,N_2338);
or U2378 (N_2378,N_2328,N_2331);
and U2379 (N_2379,N_2291,N_2282);
and U2380 (N_2380,N_2301,N_2312);
and U2381 (N_2381,N_2303,N_2327);
nor U2382 (N_2382,N_2327,N_2308);
nor U2383 (N_2383,N_2291,N_2329);
nor U2384 (N_2384,N_2324,N_2306);
nor U2385 (N_2385,N_2330,N_2313);
or U2386 (N_2386,N_2328,N_2307);
xnor U2387 (N_2387,N_2329,N_2305);
or U2388 (N_2388,N_2290,N_2304);
nand U2389 (N_2389,N_2323,N_2316);
and U2390 (N_2390,N_2330,N_2319);
or U2391 (N_2391,N_2335,N_2314);
nand U2392 (N_2392,N_2290,N_2314);
and U2393 (N_2393,N_2322,N_2306);
xor U2394 (N_2394,N_2286,N_2334);
and U2395 (N_2395,N_2316,N_2281);
nand U2396 (N_2396,N_2312,N_2324);
nor U2397 (N_2397,N_2281,N_2314);
or U2398 (N_2398,N_2339,N_2285);
or U2399 (N_2399,N_2334,N_2284);
or U2400 (N_2400,N_2379,N_2351);
nand U2401 (N_2401,N_2358,N_2382);
nor U2402 (N_2402,N_2396,N_2355);
and U2403 (N_2403,N_2366,N_2345);
or U2404 (N_2404,N_2344,N_2373);
and U2405 (N_2405,N_2368,N_2346);
or U2406 (N_2406,N_2349,N_2393);
or U2407 (N_2407,N_2354,N_2364);
nor U2408 (N_2408,N_2362,N_2360);
nand U2409 (N_2409,N_2386,N_2380);
nand U2410 (N_2410,N_2390,N_2377);
or U2411 (N_2411,N_2397,N_2392);
and U2412 (N_2412,N_2383,N_2391);
nand U2413 (N_2413,N_2361,N_2384);
nand U2414 (N_2414,N_2375,N_2381);
and U2415 (N_2415,N_2370,N_2342);
and U2416 (N_2416,N_2374,N_2347);
and U2417 (N_2417,N_2385,N_2363);
nand U2418 (N_2418,N_2387,N_2343);
and U2419 (N_2419,N_2388,N_2394);
nor U2420 (N_2420,N_2395,N_2372);
and U2421 (N_2421,N_2398,N_2353);
or U2422 (N_2422,N_2365,N_2356);
or U2423 (N_2423,N_2350,N_2357);
or U2424 (N_2424,N_2376,N_2352);
nand U2425 (N_2425,N_2369,N_2371);
and U2426 (N_2426,N_2389,N_2348);
nand U2427 (N_2427,N_2378,N_2399);
and U2428 (N_2428,N_2340,N_2359);
or U2429 (N_2429,N_2367,N_2341);
and U2430 (N_2430,N_2356,N_2364);
nor U2431 (N_2431,N_2382,N_2353);
nor U2432 (N_2432,N_2381,N_2371);
or U2433 (N_2433,N_2344,N_2397);
nor U2434 (N_2434,N_2392,N_2378);
and U2435 (N_2435,N_2353,N_2389);
and U2436 (N_2436,N_2352,N_2377);
nand U2437 (N_2437,N_2363,N_2377);
nand U2438 (N_2438,N_2359,N_2362);
or U2439 (N_2439,N_2367,N_2343);
and U2440 (N_2440,N_2399,N_2396);
nand U2441 (N_2441,N_2395,N_2353);
xor U2442 (N_2442,N_2385,N_2376);
or U2443 (N_2443,N_2376,N_2343);
nor U2444 (N_2444,N_2378,N_2398);
and U2445 (N_2445,N_2399,N_2364);
or U2446 (N_2446,N_2389,N_2386);
nor U2447 (N_2447,N_2352,N_2354);
nor U2448 (N_2448,N_2348,N_2356);
nor U2449 (N_2449,N_2381,N_2367);
nor U2450 (N_2450,N_2358,N_2356);
nor U2451 (N_2451,N_2350,N_2396);
or U2452 (N_2452,N_2378,N_2372);
nand U2453 (N_2453,N_2392,N_2379);
and U2454 (N_2454,N_2356,N_2396);
nand U2455 (N_2455,N_2371,N_2359);
and U2456 (N_2456,N_2343,N_2361);
nand U2457 (N_2457,N_2347,N_2394);
or U2458 (N_2458,N_2393,N_2390);
nor U2459 (N_2459,N_2386,N_2372);
nor U2460 (N_2460,N_2415,N_2401);
or U2461 (N_2461,N_2454,N_2409);
xor U2462 (N_2462,N_2453,N_2422);
or U2463 (N_2463,N_2416,N_2406);
nor U2464 (N_2464,N_2429,N_2418);
nand U2465 (N_2465,N_2433,N_2413);
and U2466 (N_2466,N_2427,N_2405);
and U2467 (N_2467,N_2414,N_2452);
and U2468 (N_2468,N_2444,N_2430);
or U2469 (N_2469,N_2423,N_2407);
or U2470 (N_2470,N_2408,N_2445);
or U2471 (N_2471,N_2419,N_2436);
nor U2472 (N_2472,N_2431,N_2439);
and U2473 (N_2473,N_2446,N_2447);
nor U2474 (N_2474,N_2425,N_2402);
nor U2475 (N_2475,N_2435,N_2412);
nor U2476 (N_2476,N_2449,N_2441);
nand U2477 (N_2477,N_2404,N_2417);
nand U2478 (N_2478,N_2437,N_2455);
nor U2479 (N_2479,N_2426,N_2428);
nand U2480 (N_2480,N_2456,N_2411);
and U2481 (N_2481,N_2424,N_2421);
nor U2482 (N_2482,N_2432,N_2442);
nand U2483 (N_2483,N_2400,N_2403);
and U2484 (N_2484,N_2443,N_2438);
nor U2485 (N_2485,N_2450,N_2434);
nand U2486 (N_2486,N_2420,N_2451);
and U2487 (N_2487,N_2457,N_2448);
nand U2488 (N_2488,N_2410,N_2459);
or U2489 (N_2489,N_2440,N_2458);
nor U2490 (N_2490,N_2405,N_2445);
or U2491 (N_2491,N_2419,N_2407);
or U2492 (N_2492,N_2443,N_2421);
nor U2493 (N_2493,N_2425,N_2454);
nor U2494 (N_2494,N_2402,N_2419);
nor U2495 (N_2495,N_2432,N_2425);
nor U2496 (N_2496,N_2451,N_2406);
nand U2497 (N_2497,N_2453,N_2420);
nand U2498 (N_2498,N_2454,N_2430);
nor U2499 (N_2499,N_2426,N_2408);
nand U2500 (N_2500,N_2426,N_2439);
nand U2501 (N_2501,N_2451,N_2401);
and U2502 (N_2502,N_2451,N_2437);
nor U2503 (N_2503,N_2441,N_2421);
or U2504 (N_2504,N_2406,N_2402);
or U2505 (N_2505,N_2414,N_2459);
nor U2506 (N_2506,N_2423,N_2424);
nor U2507 (N_2507,N_2434,N_2420);
and U2508 (N_2508,N_2444,N_2445);
nand U2509 (N_2509,N_2401,N_2421);
and U2510 (N_2510,N_2456,N_2422);
nor U2511 (N_2511,N_2413,N_2431);
or U2512 (N_2512,N_2458,N_2416);
or U2513 (N_2513,N_2435,N_2458);
nor U2514 (N_2514,N_2405,N_2407);
and U2515 (N_2515,N_2422,N_2439);
and U2516 (N_2516,N_2448,N_2405);
or U2517 (N_2517,N_2411,N_2405);
and U2518 (N_2518,N_2423,N_2428);
nand U2519 (N_2519,N_2414,N_2438);
or U2520 (N_2520,N_2512,N_2493);
nor U2521 (N_2521,N_2474,N_2506);
or U2522 (N_2522,N_2492,N_2499);
nand U2523 (N_2523,N_2489,N_2510);
nand U2524 (N_2524,N_2488,N_2496);
or U2525 (N_2525,N_2513,N_2511);
nand U2526 (N_2526,N_2465,N_2501);
nor U2527 (N_2527,N_2509,N_2469);
nor U2528 (N_2528,N_2482,N_2504);
xor U2529 (N_2529,N_2477,N_2497);
nor U2530 (N_2530,N_2468,N_2483);
nor U2531 (N_2531,N_2460,N_2507);
nand U2532 (N_2532,N_2505,N_2471);
nor U2533 (N_2533,N_2470,N_2486);
nand U2534 (N_2534,N_2480,N_2494);
xor U2535 (N_2535,N_2518,N_2475);
nand U2536 (N_2536,N_2461,N_2503);
nand U2537 (N_2537,N_2490,N_2467);
nor U2538 (N_2538,N_2508,N_2514);
nor U2539 (N_2539,N_2463,N_2515);
nor U2540 (N_2540,N_2502,N_2498);
nand U2541 (N_2541,N_2472,N_2500);
nand U2542 (N_2542,N_2487,N_2462);
and U2543 (N_2543,N_2481,N_2495);
and U2544 (N_2544,N_2484,N_2517);
nor U2545 (N_2545,N_2466,N_2473);
nand U2546 (N_2546,N_2491,N_2476);
nand U2547 (N_2547,N_2519,N_2464);
or U2548 (N_2548,N_2479,N_2516);
and U2549 (N_2549,N_2485,N_2478);
or U2550 (N_2550,N_2499,N_2461);
nor U2551 (N_2551,N_2508,N_2500);
or U2552 (N_2552,N_2466,N_2472);
or U2553 (N_2553,N_2472,N_2506);
or U2554 (N_2554,N_2487,N_2499);
nor U2555 (N_2555,N_2510,N_2470);
and U2556 (N_2556,N_2460,N_2492);
and U2557 (N_2557,N_2515,N_2491);
and U2558 (N_2558,N_2511,N_2467);
nor U2559 (N_2559,N_2519,N_2469);
or U2560 (N_2560,N_2488,N_2490);
or U2561 (N_2561,N_2501,N_2507);
nand U2562 (N_2562,N_2462,N_2465);
or U2563 (N_2563,N_2496,N_2491);
nor U2564 (N_2564,N_2503,N_2507);
nand U2565 (N_2565,N_2480,N_2473);
or U2566 (N_2566,N_2463,N_2461);
nor U2567 (N_2567,N_2487,N_2510);
xor U2568 (N_2568,N_2494,N_2483);
nand U2569 (N_2569,N_2506,N_2496);
nand U2570 (N_2570,N_2514,N_2499);
or U2571 (N_2571,N_2517,N_2479);
xor U2572 (N_2572,N_2492,N_2510);
nand U2573 (N_2573,N_2519,N_2493);
and U2574 (N_2574,N_2516,N_2509);
nor U2575 (N_2575,N_2465,N_2519);
or U2576 (N_2576,N_2501,N_2511);
nand U2577 (N_2577,N_2484,N_2481);
and U2578 (N_2578,N_2513,N_2493);
nand U2579 (N_2579,N_2496,N_2464);
nand U2580 (N_2580,N_2527,N_2569);
and U2581 (N_2581,N_2521,N_2570);
nand U2582 (N_2582,N_2577,N_2541);
nor U2583 (N_2583,N_2538,N_2544);
and U2584 (N_2584,N_2560,N_2550);
nor U2585 (N_2585,N_2540,N_2531);
or U2586 (N_2586,N_2548,N_2537);
or U2587 (N_2587,N_2525,N_2542);
xnor U2588 (N_2588,N_2524,N_2559);
nand U2589 (N_2589,N_2546,N_2551);
nand U2590 (N_2590,N_2558,N_2578);
nand U2591 (N_2591,N_2561,N_2530);
or U2592 (N_2592,N_2567,N_2563);
nand U2593 (N_2593,N_2576,N_2565);
nand U2594 (N_2594,N_2552,N_2528);
nand U2595 (N_2595,N_2564,N_2532);
or U2596 (N_2596,N_2568,N_2566);
nor U2597 (N_2597,N_2575,N_2555);
or U2598 (N_2598,N_2534,N_2520);
nor U2599 (N_2599,N_2572,N_2553);
or U2600 (N_2600,N_2562,N_2557);
nor U2601 (N_2601,N_2529,N_2536);
nand U2602 (N_2602,N_2535,N_2573);
nand U2603 (N_2603,N_2579,N_2549);
nor U2604 (N_2604,N_2543,N_2574);
nand U2605 (N_2605,N_2554,N_2533);
nor U2606 (N_2606,N_2523,N_2547);
nor U2607 (N_2607,N_2571,N_2539);
nor U2608 (N_2608,N_2556,N_2545);
nand U2609 (N_2609,N_2526,N_2522);
and U2610 (N_2610,N_2543,N_2569);
nor U2611 (N_2611,N_2577,N_2524);
or U2612 (N_2612,N_2552,N_2579);
or U2613 (N_2613,N_2527,N_2562);
nand U2614 (N_2614,N_2578,N_2552);
and U2615 (N_2615,N_2559,N_2565);
and U2616 (N_2616,N_2566,N_2562);
nand U2617 (N_2617,N_2526,N_2530);
or U2618 (N_2618,N_2569,N_2563);
nor U2619 (N_2619,N_2576,N_2539);
or U2620 (N_2620,N_2572,N_2549);
nor U2621 (N_2621,N_2554,N_2571);
nor U2622 (N_2622,N_2577,N_2526);
or U2623 (N_2623,N_2534,N_2543);
nand U2624 (N_2624,N_2530,N_2527);
or U2625 (N_2625,N_2577,N_2536);
nor U2626 (N_2626,N_2552,N_2550);
nand U2627 (N_2627,N_2563,N_2536);
and U2628 (N_2628,N_2571,N_2553);
nor U2629 (N_2629,N_2552,N_2538);
nand U2630 (N_2630,N_2566,N_2540);
nor U2631 (N_2631,N_2538,N_2567);
nand U2632 (N_2632,N_2569,N_2547);
nor U2633 (N_2633,N_2578,N_2531);
and U2634 (N_2634,N_2566,N_2567);
nor U2635 (N_2635,N_2547,N_2557);
nor U2636 (N_2636,N_2547,N_2539);
nor U2637 (N_2637,N_2551,N_2521);
nand U2638 (N_2638,N_2557,N_2541);
nand U2639 (N_2639,N_2542,N_2547);
or U2640 (N_2640,N_2600,N_2587);
nand U2641 (N_2641,N_2632,N_2624);
and U2642 (N_2642,N_2613,N_2623);
and U2643 (N_2643,N_2589,N_2622);
nor U2644 (N_2644,N_2602,N_2618);
nand U2645 (N_2645,N_2591,N_2626);
or U2646 (N_2646,N_2583,N_2585);
and U2647 (N_2647,N_2593,N_2633);
and U2648 (N_2648,N_2584,N_2616);
nor U2649 (N_2649,N_2610,N_2595);
nor U2650 (N_2650,N_2592,N_2629);
nor U2651 (N_2651,N_2617,N_2637);
and U2652 (N_2652,N_2581,N_2611);
nand U2653 (N_2653,N_2634,N_2638);
nor U2654 (N_2654,N_2607,N_2601);
nor U2655 (N_2655,N_2605,N_2619);
nand U2656 (N_2656,N_2586,N_2582);
nor U2657 (N_2657,N_2604,N_2621);
or U2658 (N_2658,N_2594,N_2590);
nor U2659 (N_2659,N_2606,N_2599);
and U2660 (N_2660,N_2631,N_2598);
nor U2661 (N_2661,N_2614,N_2580);
nand U2662 (N_2662,N_2628,N_2597);
or U2663 (N_2663,N_2635,N_2639);
nand U2664 (N_2664,N_2630,N_2603);
and U2665 (N_2665,N_2588,N_2612);
nand U2666 (N_2666,N_2596,N_2620);
or U2667 (N_2667,N_2627,N_2609);
nor U2668 (N_2668,N_2608,N_2625);
nor U2669 (N_2669,N_2636,N_2615);
or U2670 (N_2670,N_2638,N_2583);
or U2671 (N_2671,N_2603,N_2633);
nor U2672 (N_2672,N_2583,N_2627);
and U2673 (N_2673,N_2614,N_2592);
nand U2674 (N_2674,N_2612,N_2600);
nor U2675 (N_2675,N_2581,N_2636);
and U2676 (N_2676,N_2622,N_2608);
and U2677 (N_2677,N_2586,N_2612);
nor U2678 (N_2678,N_2595,N_2612);
nor U2679 (N_2679,N_2610,N_2588);
and U2680 (N_2680,N_2638,N_2584);
and U2681 (N_2681,N_2587,N_2613);
nor U2682 (N_2682,N_2611,N_2609);
and U2683 (N_2683,N_2580,N_2621);
and U2684 (N_2684,N_2607,N_2627);
nor U2685 (N_2685,N_2610,N_2616);
and U2686 (N_2686,N_2612,N_2632);
nor U2687 (N_2687,N_2607,N_2609);
nand U2688 (N_2688,N_2619,N_2603);
nor U2689 (N_2689,N_2631,N_2594);
and U2690 (N_2690,N_2596,N_2607);
nand U2691 (N_2691,N_2588,N_2603);
nor U2692 (N_2692,N_2586,N_2628);
or U2693 (N_2693,N_2609,N_2625);
nor U2694 (N_2694,N_2635,N_2584);
nor U2695 (N_2695,N_2591,N_2625);
or U2696 (N_2696,N_2583,N_2607);
and U2697 (N_2697,N_2636,N_2591);
nand U2698 (N_2698,N_2611,N_2619);
nand U2699 (N_2699,N_2630,N_2583);
and U2700 (N_2700,N_2670,N_2643);
nor U2701 (N_2701,N_2671,N_2676);
nor U2702 (N_2702,N_2656,N_2691);
nand U2703 (N_2703,N_2677,N_2659);
and U2704 (N_2704,N_2696,N_2655);
nor U2705 (N_2705,N_2685,N_2699);
nor U2706 (N_2706,N_2681,N_2690);
nor U2707 (N_2707,N_2665,N_2667);
nand U2708 (N_2708,N_2679,N_2650);
or U2709 (N_2709,N_2662,N_2647);
or U2710 (N_2710,N_2675,N_2646);
nand U2711 (N_2711,N_2672,N_2658);
nand U2712 (N_2712,N_2645,N_2693);
nand U2713 (N_2713,N_2689,N_2695);
or U2714 (N_2714,N_2684,N_2678);
or U2715 (N_2715,N_2660,N_2680);
or U2716 (N_2716,N_2657,N_2652);
nor U2717 (N_2717,N_2687,N_2654);
nand U2718 (N_2718,N_2661,N_2648);
nor U2719 (N_2719,N_2651,N_2674);
or U2720 (N_2720,N_2644,N_2686);
or U2721 (N_2721,N_2653,N_2697);
or U2722 (N_2722,N_2694,N_2668);
or U2723 (N_2723,N_2692,N_2640);
nor U2724 (N_2724,N_2663,N_2682);
and U2725 (N_2725,N_2664,N_2649);
or U2726 (N_2726,N_2669,N_2666);
nor U2727 (N_2727,N_2641,N_2642);
and U2728 (N_2728,N_2688,N_2673);
or U2729 (N_2729,N_2683,N_2698);
and U2730 (N_2730,N_2655,N_2699);
and U2731 (N_2731,N_2648,N_2645);
or U2732 (N_2732,N_2668,N_2699);
or U2733 (N_2733,N_2659,N_2678);
or U2734 (N_2734,N_2640,N_2689);
and U2735 (N_2735,N_2649,N_2677);
xnor U2736 (N_2736,N_2688,N_2662);
nand U2737 (N_2737,N_2681,N_2673);
nor U2738 (N_2738,N_2677,N_2678);
or U2739 (N_2739,N_2687,N_2643);
nor U2740 (N_2740,N_2662,N_2667);
or U2741 (N_2741,N_2688,N_2678);
or U2742 (N_2742,N_2673,N_2679);
or U2743 (N_2743,N_2692,N_2685);
or U2744 (N_2744,N_2646,N_2692);
nor U2745 (N_2745,N_2695,N_2658);
or U2746 (N_2746,N_2685,N_2663);
or U2747 (N_2747,N_2662,N_2691);
nor U2748 (N_2748,N_2661,N_2651);
and U2749 (N_2749,N_2640,N_2679);
nor U2750 (N_2750,N_2654,N_2649);
nand U2751 (N_2751,N_2690,N_2661);
and U2752 (N_2752,N_2640,N_2677);
or U2753 (N_2753,N_2670,N_2645);
or U2754 (N_2754,N_2698,N_2670);
nand U2755 (N_2755,N_2647,N_2641);
nor U2756 (N_2756,N_2651,N_2672);
nor U2757 (N_2757,N_2691,N_2641);
nor U2758 (N_2758,N_2689,N_2651);
nor U2759 (N_2759,N_2682,N_2684);
and U2760 (N_2760,N_2718,N_2730);
nand U2761 (N_2761,N_2719,N_2740);
and U2762 (N_2762,N_2748,N_2758);
or U2763 (N_2763,N_2729,N_2734);
and U2764 (N_2764,N_2726,N_2741);
nand U2765 (N_2765,N_2701,N_2739);
nand U2766 (N_2766,N_2753,N_2724);
nand U2767 (N_2767,N_2700,N_2744);
nand U2768 (N_2768,N_2712,N_2754);
nor U2769 (N_2769,N_2756,N_2703);
nor U2770 (N_2770,N_2738,N_2722);
nor U2771 (N_2771,N_2725,N_2727);
and U2772 (N_2772,N_2716,N_2704);
or U2773 (N_2773,N_2747,N_2723);
or U2774 (N_2774,N_2751,N_2752);
or U2775 (N_2775,N_2737,N_2746);
or U2776 (N_2776,N_2728,N_2720);
nand U2777 (N_2777,N_2732,N_2735);
or U2778 (N_2778,N_2715,N_2749);
or U2779 (N_2779,N_2710,N_2757);
nand U2780 (N_2780,N_2745,N_2750);
and U2781 (N_2781,N_2707,N_2713);
and U2782 (N_2782,N_2714,N_2705);
or U2783 (N_2783,N_2733,N_2706);
or U2784 (N_2784,N_2731,N_2736);
and U2785 (N_2785,N_2708,N_2743);
nand U2786 (N_2786,N_2759,N_2717);
or U2787 (N_2787,N_2742,N_2709);
nor U2788 (N_2788,N_2702,N_2721);
nor U2789 (N_2789,N_2755,N_2711);
nor U2790 (N_2790,N_2751,N_2732);
nor U2791 (N_2791,N_2706,N_2729);
and U2792 (N_2792,N_2757,N_2745);
or U2793 (N_2793,N_2744,N_2725);
or U2794 (N_2794,N_2730,N_2719);
and U2795 (N_2795,N_2757,N_2707);
and U2796 (N_2796,N_2756,N_2706);
nor U2797 (N_2797,N_2747,N_2757);
or U2798 (N_2798,N_2717,N_2720);
nor U2799 (N_2799,N_2712,N_2707);
and U2800 (N_2800,N_2716,N_2757);
nor U2801 (N_2801,N_2758,N_2723);
or U2802 (N_2802,N_2705,N_2708);
or U2803 (N_2803,N_2721,N_2729);
nand U2804 (N_2804,N_2709,N_2758);
nand U2805 (N_2805,N_2743,N_2752);
nand U2806 (N_2806,N_2709,N_2723);
nor U2807 (N_2807,N_2748,N_2708);
or U2808 (N_2808,N_2753,N_2736);
and U2809 (N_2809,N_2754,N_2758);
and U2810 (N_2810,N_2749,N_2707);
nand U2811 (N_2811,N_2705,N_2719);
nor U2812 (N_2812,N_2718,N_2746);
nor U2813 (N_2813,N_2706,N_2710);
nand U2814 (N_2814,N_2747,N_2753);
nor U2815 (N_2815,N_2738,N_2730);
or U2816 (N_2816,N_2700,N_2752);
nand U2817 (N_2817,N_2701,N_2741);
and U2818 (N_2818,N_2726,N_2713);
and U2819 (N_2819,N_2709,N_2718);
nand U2820 (N_2820,N_2786,N_2783);
nor U2821 (N_2821,N_2794,N_2769);
nor U2822 (N_2822,N_2780,N_2810);
or U2823 (N_2823,N_2766,N_2788);
nand U2824 (N_2824,N_2803,N_2791);
nand U2825 (N_2825,N_2774,N_2819);
nor U2826 (N_2826,N_2805,N_2802);
or U2827 (N_2827,N_2777,N_2773);
and U2828 (N_2828,N_2812,N_2784);
and U2829 (N_2829,N_2775,N_2813);
or U2830 (N_2830,N_2761,N_2806);
and U2831 (N_2831,N_2772,N_2817);
nor U2832 (N_2832,N_2787,N_2809);
nand U2833 (N_2833,N_2771,N_2779);
nand U2834 (N_2834,N_2795,N_2760);
or U2835 (N_2835,N_2816,N_2799);
nor U2836 (N_2836,N_2808,N_2776);
or U2837 (N_2837,N_2764,N_2797);
or U2838 (N_2838,N_2765,N_2807);
or U2839 (N_2839,N_2770,N_2815);
nor U2840 (N_2840,N_2767,N_2796);
xnor U2841 (N_2841,N_2785,N_2798);
nand U2842 (N_2842,N_2793,N_2800);
nor U2843 (N_2843,N_2801,N_2778);
nor U2844 (N_2844,N_2790,N_2818);
nor U2845 (N_2845,N_2804,N_2768);
nand U2846 (N_2846,N_2781,N_2782);
or U2847 (N_2847,N_2792,N_2811);
and U2848 (N_2848,N_2789,N_2762);
nor U2849 (N_2849,N_2763,N_2814);
or U2850 (N_2850,N_2761,N_2764);
or U2851 (N_2851,N_2808,N_2815);
or U2852 (N_2852,N_2772,N_2800);
or U2853 (N_2853,N_2797,N_2781);
nand U2854 (N_2854,N_2790,N_2767);
or U2855 (N_2855,N_2811,N_2787);
nor U2856 (N_2856,N_2818,N_2803);
nor U2857 (N_2857,N_2765,N_2782);
or U2858 (N_2858,N_2772,N_2779);
nor U2859 (N_2859,N_2768,N_2798);
and U2860 (N_2860,N_2783,N_2763);
nand U2861 (N_2861,N_2798,N_2793);
or U2862 (N_2862,N_2788,N_2791);
nor U2863 (N_2863,N_2797,N_2776);
nor U2864 (N_2864,N_2803,N_2799);
nand U2865 (N_2865,N_2816,N_2785);
or U2866 (N_2866,N_2800,N_2796);
and U2867 (N_2867,N_2771,N_2785);
nor U2868 (N_2868,N_2799,N_2813);
nand U2869 (N_2869,N_2796,N_2815);
or U2870 (N_2870,N_2778,N_2769);
nand U2871 (N_2871,N_2807,N_2787);
nor U2872 (N_2872,N_2815,N_2810);
or U2873 (N_2873,N_2769,N_2761);
and U2874 (N_2874,N_2811,N_2785);
or U2875 (N_2875,N_2816,N_2798);
nand U2876 (N_2876,N_2775,N_2787);
nor U2877 (N_2877,N_2787,N_2798);
nand U2878 (N_2878,N_2763,N_2774);
nor U2879 (N_2879,N_2767,N_2806);
and U2880 (N_2880,N_2840,N_2842);
nor U2881 (N_2881,N_2831,N_2834);
nand U2882 (N_2882,N_2829,N_2835);
nor U2883 (N_2883,N_2879,N_2836);
nor U2884 (N_2884,N_2853,N_2859);
and U2885 (N_2885,N_2844,N_2846);
or U2886 (N_2886,N_2873,N_2822);
nand U2887 (N_2887,N_2866,N_2856);
and U2888 (N_2888,N_2841,N_2830);
nor U2889 (N_2889,N_2843,N_2850);
or U2890 (N_2890,N_2825,N_2839);
or U2891 (N_2891,N_2868,N_2874);
nand U2892 (N_2892,N_2824,N_2863);
nor U2893 (N_2893,N_2877,N_2871);
and U2894 (N_2894,N_2855,N_2849);
nor U2895 (N_2895,N_2872,N_2848);
nand U2896 (N_2896,N_2860,N_2865);
and U2897 (N_2897,N_2878,N_2851);
xnor U2898 (N_2898,N_2869,N_2864);
and U2899 (N_2899,N_2821,N_2870);
or U2900 (N_2900,N_2858,N_2820);
and U2901 (N_2901,N_2867,N_2857);
nor U2902 (N_2902,N_2875,N_2838);
nand U2903 (N_2903,N_2827,N_2862);
and U2904 (N_2904,N_2861,N_2876);
and U2905 (N_2905,N_2837,N_2832);
or U2906 (N_2906,N_2826,N_2854);
nand U2907 (N_2907,N_2833,N_2823);
or U2908 (N_2908,N_2847,N_2852);
and U2909 (N_2909,N_2845,N_2828);
nor U2910 (N_2910,N_2835,N_2827);
or U2911 (N_2911,N_2840,N_2873);
nand U2912 (N_2912,N_2825,N_2873);
or U2913 (N_2913,N_2865,N_2862);
or U2914 (N_2914,N_2867,N_2850);
or U2915 (N_2915,N_2831,N_2879);
nor U2916 (N_2916,N_2834,N_2846);
or U2917 (N_2917,N_2874,N_2830);
or U2918 (N_2918,N_2867,N_2841);
nand U2919 (N_2919,N_2829,N_2827);
nor U2920 (N_2920,N_2872,N_2851);
nor U2921 (N_2921,N_2852,N_2866);
nor U2922 (N_2922,N_2849,N_2823);
nor U2923 (N_2923,N_2861,N_2821);
or U2924 (N_2924,N_2834,N_2822);
nor U2925 (N_2925,N_2873,N_2862);
and U2926 (N_2926,N_2870,N_2833);
or U2927 (N_2927,N_2840,N_2820);
nand U2928 (N_2928,N_2879,N_2820);
nand U2929 (N_2929,N_2857,N_2859);
nor U2930 (N_2930,N_2858,N_2844);
and U2931 (N_2931,N_2849,N_2844);
nand U2932 (N_2932,N_2826,N_2838);
and U2933 (N_2933,N_2861,N_2826);
and U2934 (N_2934,N_2826,N_2851);
or U2935 (N_2935,N_2850,N_2862);
nor U2936 (N_2936,N_2851,N_2825);
and U2937 (N_2937,N_2865,N_2835);
nor U2938 (N_2938,N_2851,N_2869);
or U2939 (N_2939,N_2875,N_2856);
and U2940 (N_2940,N_2917,N_2901);
or U2941 (N_2941,N_2895,N_2920);
nor U2942 (N_2942,N_2939,N_2918);
nand U2943 (N_2943,N_2913,N_2911);
nor U2944 (N_2944,N_2908,N_2910);
and U2945 (N_2945,N_2925,N_2930);
and U2946 (N_2946,N_2897,N_2888);
and U2947 (N_2947,N_2905,N_2890);
nand U2948 (N_2948,N_2926,N_2903);
nand U2949 (N_2949,N_2919,N_2886);
or U2950 (N_2950,N_2882,N_2899);
and U2951 (N_2951,N_2892,N_2938);
nand U2952 (N_2952,N_2880,N_2889);
nor U2953 (N_2953,N_2928,N_2898);
and U2954 (N_2954,N_2914,N_2909);
nor U2955 (N_2955,N_2912,N_2923);
xnor U2956 (N_2956,N_2916,N_2936);
and U2957 (N_2957,N_2933,N_2904);
and U2958 (N_2958,N_2937,N_2893);
or U2959 (N_2959,N_2915,N_2934);
and U2960 (N_2960,N_2906,N_2931);
or U2961 (N_2961,N_2883,N_2927);
and U2962 (N_2962,N_2887,N_2884);
or U2963 (N_2963,N_2924,N_2929);
and U2964 (N_2964,N_2932,N_2907);
nand U2965 (N_2965,N_2885,N_2881);
and U2966 (N_2966,N_2896,N_2894);
or U2967 (N_2967,N_2935,N_2922);
nand U2968 (N_2968,N_2900,N_2921);
or U2969 (N_2969,N_2902,N_2891);
nand U2970 (N_2970,N_2897,N_2907);
nand U2971 (N_2971,N_2894,N_2919);
nor U2972 (N_2972,N_2911,N_2887);
or U2973 (N_2973,N_2909,N_2883);
nand U2974 (N_2974,N_2927,N_2925);
or U2975 (N_2975,N_2927,N_2906);
and U2976 (N_2976,N_2932,N_2921);
or U2977 (N_2977,N_2920,N_2889);
or U2978 (N_2978,N_2918,N_2891);
or U2979 (N_2979,N_2886,N_2929);
nand U2980 (N_2980,N_2935,N_2938);
nor U2981 (N_2981,N_2881,N_2900);
nand U2982 (N_2982,N_2905,N_2884);
and U2983 (N_2983,N_2887,N_2890);
nor U2984 (N_2984,N_2937,N_2884);
nor U2985 (N_2985,N_2897,N_2926);
nor U2986 (N_2986,N_2900,N_2913);
nand U2987 (N_2987,N_2929,N_2908);
or U2988 (N_2988,N_2935,N_2932);
or U2989 (N_2989,N_2919,N_2904);
nand U2990 (N_2990,N_2923,N_2884);
and U2991 (N_2991,N_2892,N_2928);
nand U2992 (N_2992,N_2907,N_2912);
nor U2993 (N_2993,N_2899,N_2924);
nor U2994 (N_2994,N_2931,N_2937);
and U2995 (N_2995,N_2901,N_2886);
nor U2996 (N_2996,N_2919,N_2912);
nor U2997 (N_2997,N_2902,N_2886);
and U2998 (N_2998,N_2886,N_2933);
nor U2999 (N_2999,N_2901,N_2933);
nor UO_0 (O_0,N_2979,N_2947);
nor UO_1 (O_1,N_2971,N_2969);
nand UO_2 (O_2,N_2992,N_2964);
nor UO_3 (O_3,N_2951,N_2948);
nand UO_4 (O_4,N_2982,N_2959);
nor UO_5 (O_5,N_2954,N_2945);
nor UO_6 (O_6,N_2967,N_2950);
nor UO_7 (O_7,N_2963,N_2995);
nor UO_8 (O_8,N_2949,N_2975);
nand UO_9 (O_9,N_2955,N_2978);
and UO_10 (O_10,N_2942,N_2998);
and UO_11 (O_11,N_2983,N_2952);
and UO_12 (O_12,N_2987,N_2993);
nand UO_13 (O_13,N_2960,N_2944);
nand UO_14 (O_14,N_2966,N_2980);
nand UO_15 (O_15,N_2943,N_2990);
and UO_16 (O_16,N_2970,N_2940);
or UO_17 (O_17,N_2957,N_2984);
nand UO_18 (O_18,N_2991,N_2981);
xor UO_19 (O_19,N_2977,N_2976);
and UO_20 (O_20,N_2956,N_2985);
nand UO_21 (O_21,N_2999,N_2965);
nor UO_22 (O_22,N_2953,N_2958);
nor UO_23 (O_23,N_2988,N_2973);
or UO_24 (O_24,N_2986,N_2941);
and UO_25 (O_25,N_2997,N_2961);
or UO_26 (O_26,N_2962,N_2974);
and UO_27 (O_27,N_2968,N_2946);
nor UO_28 (O_28,N_2989,N_2972);
and UO_29 (O_29,N_2994,N_2996);
and UO_30 (O_30,N_2992,N_2974);
nand UO_31 (O_31,N_2972,N_2978);
nand UO_32 (O_32,N_2971,N_2968);
nor UO_33 (O_33,N_2969,N_2983);
or UO_34 (O_34,N_2998,N_2979);
and UO_35 (O_35,N_2946,N_2960);
and UO_36 (O_36,N_2990,N_2973);
xnor UO_37 (O_37,N_2971,N_2964);
and UO_38 (O_38,N_2940,N_2946);
and UO_39 (O_39,N_2994,N_2956);
and UO_40 (O_40,N_2974,N_2980);
or UO_41 (O_41,N_2969,N_2964);
or UO_42 (O_42,N_2967,N_2990);
or UO_43 (O_43,N_2974,N_2958);
or UO_44 (O_44,N_2974,N_2979);
or UO_45 (O_45,N_2998,N_2964);
nor UO_46 (O_46,N_2948,N_2972);
nand UO_47 (O_47,N_2971,N_2983);
nor UO_48 (O_48,N_2981,N_2989);
nand UO_49 (O_49,N_2999,N_2989);
nor UO_50 (O_50,N_2942,N_2996);
or UO_51 (O_51,N_2957,N_2980);
and UO_52 (O_52,N_2972,N_2988);
or UO_53 (O_53,N_2942,N_2976);
nor UO_54 (O_54,N_2970,N_2950);
nand UO_55 (O_55,N_2984,N_2996);
or UO_56 (O_56,N_2942,N_2991);
or UO_57 (O_57,N_2960,N_2954);
or UO_58 (O_58,N_2959,N_2978);
and UO_59 (O_59,N_2963,N_2979);
or UO_60 (O_60,N_2984,N_2977);
nor UO_61 (O_61,N_2976,N_2960);
and UO_62 (O_62,N_2945,N_2984);
nor UO_63 (O_63,N_2958,N_2963);
nand UO_64 (O_64,N_2989,N_2958);
nand UO_65 (O_65,N_2975,N_2999);
or UO_66 (O_66,N_2987,N_2944);
and UO_67 (O_67,N_2972,N_2996);
or UO_68 (O_68,N_2989,N_2986);
nor UO_69 (O_69,N_2992,N_2943);
and UO_70 (O_70,N_2959,N_2954);
nand UO_71 (O_71,N_2981,N_2973);
or UO_72 (O_72,N_2960,N_2950);
and UO_73 (O_73,N_2983,N_2978);
xnor UO_74 (O_74,N_2994,N_2968);
nand UO_75 (O_75,N_2969,N_2941);
or UO_76 (O_76,N_2992,N_2947);
and UO_77 (O_77,N_2944,N_2958);
nor UO_78 (O_78,N_2977,N_2973);
and UO_79 (O_79,N_2951,N_2949);
nor UO_80 (O_80,N_2969,N_2998);
nand UO_81 (O_81,N_2956,N_2963);
or UO_82 (O_82,N_2944,N_2977);
and UO_83 (O_83,N_2948,N_2996);
nor UO_84 (O_84,N_2969,N_2986);
nand UO_85 (O_85,N_2971,N_2981);
and UO_86 (O_86,N_2961,N_2969);
and UO_87 (O_87,N_2958,N_2972);
and UO_88 (O_88,N_2980,N_2942);
nand UO_89 (O_89,N_2997,N_2956);
nand UO_90 (O_90,N_2957,N_2987);
or UO_91 (O_91,N_2963,N_2961);
and UO_92 (O_92,N_2987,N_2960);
and UO_93 (O_93,N_2976,N_2973);
nand UO_94 (O_94,N_2940,N_2991);
nand UO_95 (O_95,N_2949,N_2987);
and UO_96 (O_96,N_2972,N_2979);
or UO_97 (O_97,N_2995,N_2943);
nor UO_98 (O_98,N_2980,N_2970);
or UO_99 (O_99,N_2965,N_2982);
nand UO_100 (O_100,N_2986,N_2992);
nand UO_101 (O_101,N_2980,N_2993);
nand UO_102 (O_102,N_2992,N_2940);
and UO_103 (O_103,N_2955,N_2962);
or UO_104 (O_104,N_2983,N_2949);
nand UO_105 (O_105,N_2974,N_2999);
nor UO_106 (O_106,N_2976,N_2999);
and UO_107 (O_107,N_2990,N_2959);
or UO_108 (O_108,N_2981,N_2982);
or UO_109 (O_109,N_2998,N_2999);
nand UO_110 (O_110,N_2959,N_2969);
or UO_111 (O_111,N_2965,N_2940);
nor UO_112 (O_112,N_2971,N_2949);
nor UO_113 (O_113,N_2996,N_2973);
nor UO_114 (O_114,N_2986,N_2972);
or UO_115 (O_115,N_2968,N_2952);
and UO_116 (O_116,N_2969,N_2973);
nand UO_117 (O_117,N_2981,N_2974);
nand UO_118 (O_118,N_2948,N_2973);
nand UO_119 (O_119,N_2951,N_2990);
nor UO_120 (O_120,N_2963,N_2972);
and UO_121 (O_121,N_2944,N_2997);
nor UO_122 (O_122,N_2946,N_2962);
nor UO_123 (O_123,N_2979,N_2984);
nor UO_124 (O_124,N_2973,N_2942);
or UO_125 (O_125,N_2995,N_2999);
nor UO_126 (O_126,N_2961,N_2941);
nand UO_127 (O_127,N_2958,N_2947);
nand UO_128 (O_128,N_2982,N_2941);
xnor UO_129 (O_129,N_2953,N_2944);
or UO_130 (O_130,N_2944,N_2983);
nor UO_131 (O_131,N_2986,N_2940);
nand UO_132 (O_132,N_2944,N_2995);
and UO_133 (O_133,N_2974,N_2985);
and UO_134 (O_134,N_2998,N_2961);
or UO_135 (O_135,N_2961,N_2989);
nand UO_136 (O_136,N_2992,N_2953);
nand UO_137 (O_137,N_2979,N_2995);
or UO_138 (O_138,N_2941,N_2978);
nand UO_139 (O_139,N_2955,N_2954);
or UO_140 (O_140,N_2961,N_2979);
and UO_141 (O_141,N_2993,N_2971);
or UO_142 (O_142,N_2999,N_2984);
and UO_143 (O_143,N_2992,N_2999);
or UO_144 (O_144,N_2991,N_2954);
and UO_145 (O_145,N_2962,N_2999);
or UO_146 (O_146,N_2985,N_2961);
or UO_147 (O_147,N_2941,N_2975);
or UO_148 (O_148,N_2981,N_2947);
nand UO_149 (O_149,N_2941,N_2943);
nand UO_150 (O_150,N_2945,N_2977);
and UO_151 (O_151,N_2945,N_2986);
or UO_152 (O_152,N_2955,N_2990);
and UO_153 (O_153,N_2984,N_2997);
or UO_154 (O_154,N_2966,N_2992);
nand UO_155 (O_155,N_2978,N_2946);
nand UO_156 (O_156,N_2943,N_2960);
nand UO_157 (O_157,N_2996,N_2990);
or UO_158 (O_158,N_2985,N_2948);
nand UO_159 (O_159,N_2996,N_2954);
nand UO_160 (O_160,N_2977,N_2993);
nand UO_161 (O_161,N_2987,N_2956);
and UO_162 (O_162,N_2958,N_2993);
and UO_163 (O_163,N_2994,N_2946);
nor UO_164 (O_164,N_2997,N_2946);
or UO_165 (O_165,N_2965,N_2967);
or UO_166 (O_166,N_2950,N_2981);
or UO_167 (O_167,N_2953,N_2968);
nor UO_168 (O_168,N_2953,N_2996);
or UO_169 (O_169,N_2993,N_2988);
nand UO_170 (O_170,N_2980,N_2953);
nor UO_171 (O_171,N_2951,N_2968);
and UO_172 (O_172,N_2969,N_2956);
and UO_173 (O_173,N_2996,N_2985);
nand UO_174 (O_174,N_2943,N_2962);
and UO_175 (O_175,N_2986,N_2961);
nor UO_176 (O_176,N_2972,N_2943);
and UO_177 (O_177,N_2991,N_2967);
or UO_178 (O_178,N_2958,N_2946);
and UO_179 (O_179,N_2947,N_2996);
nor UO_180 (O_180,N_2971,N_2994);
or UO_181 (O_181,N_2942,N_2970);
nand UO_182 (O_182,N_2984,N_2948);
or UO_183 (O_183,N_2977,N_2942);
or UO_184 (O_184,N_2971,N_2973);
nor UO_185 (O_185,N_2955,N_2964);
nand UO_186 (O_186,N_2957,N_2990);
or UO_187 (O_187,N_2981,N_2952);
nand UO_188 (O_188,N_2950,N_2990);
nor UO_189 (O_189,N_2970,N_2956);
nand UO_190 (O_190,N_2946,N_2982);
nand UO_191 (O_191,N_2955,N_2984);
nand UO_192 (O_192,N_2963,N_2967);
nand UO_193 (O_193,N_2990,N_2964);
nand UO_194 (O_194,N_2960,N_2991);
or UO_195 (O_195,N_2977,N_2968);
or UO_196 (O_196,N_2944,N_2974);
nand UO_197 (O_197,N_2965,N_2954);
nor UO_198 (O_198,N_2972,N_2964);
and UO_199 (O_199,N_2942,N_2962);
or UO_200 (O_200,N_2981,N_2953);
and UO_201 (O_201,N_2998,N_2959);
nor UO_202 (O_202,N_2998,N_2990);
nor UO_203 (O_203,N_2972,N_2983);
nor UO_204 (O_204,N_2941,N_2944);
nor UO_205 (O_205,N_2963,N_2997);
nand UO_206 (O_206,N_2963,N_2960);
nor UO_207 (O_207,N_2980,N_2975);
nand UO_208 (O_208,N_2962,N_2996);
or UO_209 (O_209,N_2949,N_2958);
nand UO_210 (O_210,N_2967,N_2992);
and UO_211 (O_211,N_2991,N_2978);
nand UO_212 (O_212,N_2982,N_2952);
or UO_213 (O_213,N_2998,N_2971);
or UO_214 (O_214,N_2947,N_2957);
nand UO_215 (O_215,N_2962,N_2940);
nand UO_216 (O_216,N_2967,N_2972);
nor UO_217 (O_217,N_2992,N_2984);
nand UO_218 (O_218,N_2996,N_2960);
nor UO_219 (O_219,N_2945,N_2990);
or UO_220 (O_220,N_2940,N_2954);
nor UO_221 (O_221,N_2970,N_2997);
nor UO_222 (O_222,N_2954,N_2946);
or UO_223 (O_223,N_2982,N_2987);
or UO_224 (O_224,N_2985,N_2964);
or UO_225 (O_225,N_2952,N_2955);
and UO_226 (O_226,N_2990,N_2987);
nand UO_227 (O_227,N_2994,N_2972);
nand UO_228 (O_228,N_2980,N_2976);
and UO_229 (O_229,N_2965,N_2983);
nor UO_230 (O_230,N_2984,N_2988);
nor UO_231 (O_231,N_2944,N_2978);
or UO_232 (O_232,N_2959,N_2956);
nor UO_233 (O_233,N_2976,N_2969);
and UO_234 (O_234,N_2983,N_2968);
or UO_235 (O_235,N_2958,N_2950);
or UO_236 (O_236,N_2946,N_2979);
nor UO_237 (O_237,N_2953,N_2949);
or UO_238 (O_238,N_2975,N_2955);
and UO_239 (O_239,N_2958,N_2999);
and UO_240 (O_240,N_2972,N_2957);
nand UO_241 (O_241,N_2961,N_2995);
or UO_242 (O_242,N_2948,N_2946);
nor UO_243 (O_243,N_2988,N_2956);
nor UO_244 (O_244,N_2945,N_2968);
nor UO_245 (O_245,N_2968,N_2990);
or UO_246 (O_246,N_2967,N_2947);
nor UO_247 (O_247,N_2980,N_2996);
nand UO_248 (O_248,N_2961,N_2994);
and UO_249 (O_249,N_2972,N_2981);
nor UO_250 (O_250,N_2988,N_2975);
nand UO_251 (O_251,N_2966,N_2993);
and UO_252 (O_252,N_2945,N_2983);
nand UO_253 (O_253,N_2999,N_2982);
nand UO_254 (O_254,N_2978,N_2981);
nor UO_255 (O_255,N_2996,N_2969);
nand UO_256 (O_256,N_2976,N_2968);
or UO_257 (O_257,N_2940,N_2949);
or UO_258 (O_258,N_2990,N_2940);
nand UO_259 (O_259,N_2968,N_2998);
and UO_260 (O_260,N_2947,N_2964);
and UO_261 (O_261,N_2982,N_2971);
nand UO_262 (O_262,N_2949,N_2946);
and UO_263 (O_263,N_2965,N_2984);
nor UO_264 (O_264,N_2983,N_2999);
and UO_265 (O_265,N_2956,N_2973);
nor UO_266 (O_266,N_2971,N_2958);
nand UO_267 (O_267,N_2954,N_2947);
or UO_268 (O_268,N_2995,N_2976);
and UO_269 (O_269,N_2990,N_2953);
and UO_270 (O_270,N_2981,N_2976);
and UO_271 (O_271,N_2986,N_2955);
nor UO_272 (O_272,N_2990,N_2942);
nand UO_273 (O_273,N_2951,N_2995);
xor UO_274 (O_274,N_2983,N_2957);
nor UO_275 (O_275,N_2967,N_2993);
or UO_276 (O_276,N_2964,N_2941);
or UO_277 (O_277,N_2951,N_2980);
or UO_278 (O_278,N_2942,N_2950);
and UO_279 (O_279,N_2984,N_2947);
nand UO_280 (O_280,N_2948,N_2975);
nand UO_281 (O_281,N_2999,N_2996);
or UO_282 (O_282,N_2991,N_2984);
or UO_283 (O_283,N_2964,N_2989);
nand UO_284 (O_284,N_2956,N_2955);
nand UO_285 (O_285,N_2965,N_2992);
nand UO_286 (O_286,N_2974,N_2967);
nand UO_287 (O_287,N_2972,N_2990);
or UO_288 (O_288,N_2969,N_2947);
nand UO_289 (O_289,N_2972,N_2965);
and UO_290 (O_290,N_2955,N_2971);
or UO_291 (O_291,N_2953,N_2957);
or UO_292 (O_292,N_2991,N_2958);
and UO_293 (O_293,N_2986,N_2981);
and UO_294 (O_294,N_2984,N_2960);
nand UO_295 (O_295,N_2998,N_2962);
or UO_296 (O_296,N_2974,N_2965);
nand UO_297 (O_297,N_2979,N_2943);
and UO_298 (O_298,N_2964,N_2942);
and UO_299 (O_299,N_2968,N_2959);
or UO_300 (O_300,N_2952,N_2993);
and UO_301 (O_301,N_2973,N_2943);
and UO_302 (O_302,N_2989,N_2968);
nor UO_303 (O_303,N_2961,N_2982);
nand UO_304 (O_304,N_2948,N_2969);
or UO_305 (O_305,N_2996,N_2982);
and UO_306 (O_306,N_2981,N_2990);
and UO_307 (O_307,N_2987,N_2945);
nor UO_308 (O_308,N_2962,N_2978);
nor UO_309 (O_309,N_2956,N_2982);
nand UO_310 (O_310,N_2970,N_2994);
nand UO_311 (O_311,N_2979,N_2966);
and UO_312 (O_312,N_2949,N_2961);
nor UO_313 (O_313,N_2988,N_2942);
nand UO_314 (O_314,N_2991,N_2977);
nor UO_315 (O_315,N_2995,N_2970);
and UO_316 (O_316,N_2946,N_2976);
and UO_317 (O_317,N_2973,N_2947);
and UO_318 (O_318,N_2951,N_2955);
and UO_319 (O_319,N_2943,N_2940);
nand UO_320 (O_320,N_2971,N_2948);
or UO_321 (O_321,N_2985,N_2976);
or UO_322 (O_322,N_2948,N_2956);
nor UO_323 (O_323,N_2975,N_2960);
nand UO_324 (O_324,N_2995,N_2991);
nand UO_325 (O_325,N_2977,N_2955);
or UO_326 (O_326,N_2965,N_2950);
nor UO_327 (O_327,N_2991,N_2961);
nand UO_328 (O_328,N_2983,N_2997);
or UO_329 (O_329,N_2978,N_2975);
and UO_330 (O_330,N_2950,N_2982);
and UO_331 (O_331,N_2988,N_2998);
and UO_332 (O_332,N_2954,N_2967);
or UO_333 (O_333,N_2994,N_2986);
nand UO_334 (O_334,N_2998,N_2972);
nor UO_335 (O_335,N_2962,N_2950);
nor UO_336 (O_336,N_2957,N_2966);
nand UO_337 (O_337,N_2996,N_2971);
nand UO_338 (O_338,N_2984,N_2946);
nand UO_339 (O_339,N_2958,N_2997);
nand UO_340 (O_340,N_2969,N_2987);
nand UO_341 (O_341,N_2952,N_2943);
and UO_342 (O_342,N_2956,N_2998);
or UO_343 (O_343,N_2946,N_2980);
nand UO_344 (O_344,N_2967,N_2986);
nor UO_345 (O_345,N_2955,N_2948);
nor UO_346 (O_346,N_2970,N_2945);
nor UO_347 (O_347,N_2941,N_2949);
nor UO_348 (O_348,N_2956,N_2972);
nand UO_349 (O_349,N_2962,N_2992);
or UO_350 (O_350,N_2966,N_2944);
nand UO_351 (O_351,N_2974,N_2993);
nand UO_352 (O_352,N_2958,N_2943);
nand UO_353 (O_353,N_2952,N_2985);
or UO_354 (O_354,N_2961,N_2954);
or UO_355 (O_355,N_2963,N_2976);
nand UO_356 (O_356,N_2986,N_2952);
or UO_357 (O_357,N_2983,N_2975);
nor UO_358 (O_358,N_2952,N_2999);
nor UO_359 (O_359,N_2958,N_2998);
nand UO_360 (O_360,N_2965,N_2955);
nand UO_361 (O_361,N_2960,N_2990);
or UO_362 (O_362,N_2968,N_2985);
nand UO_363 (O_363,N_2988,N_2980);
nand UO_364 (O_364,N_2992,N_2997);
nor UO_365 (O_365,N_2969,N_2991);
or UO_366 (O_366,N_2960,N_2958);
nand UO_367 (O_367,N_2982,N_2990);
nor UO_368 (O_368,N_2962,N_2945);
nand UO_369 (O_369,N_2988,N_2992);
nand UO_370 (O_370,N_2978,N_2967);
or UO_371 (O_371,N_2992,N_2995);
or UO_372 (O_372,N_2999,N_2978);
nand UO_373 (O_373,N_2990,N_2978);
nor UO_374 (O_374,N_2992,N_2954);
or UO_375 (O_375,N_2999,N_2946);
nand UO_376 (O_376,N_2992,N_2942);
or UO_377 (O_377,N_2941,N_2956);
or UO_378 (O_378,N_2965,N_2942);
nor UO_379 (O_379,N_2989,N_2996);
nor UO_380 (O_380,N_2975,N_2998);
nor UO_381 (O_381,N_2988,N_2954);
nor UO_382 (O_382,N_2991,N_2974);
and UO_383 (O_383,N_2991,N_2994);
nand UO_384 (O_384,N_2972,N_2960);
or UO_385 (O_385,N_2985,N_2981);
and UO_386 (O_386,N_2956,N_2993);
nand UO_387 (O_387,N_2959,N_2949);
nand UO_388 (O_388,N_2950,N_2978);
or UO_389 (O_389,N_2959,N_2995);
nor UO_390 (O_390,N_2958,N_2995);
nand UO_391 (O_391,N_2997,N_2972);
nand UO_392 (O_392,N_2966,N_2990);
nand UO_393 (O_393,N_2953,N_2961);
and UO_394 (O_394,N_2987,N_2967);
nand UO_395 (O_395,N_2947,N_2953);
nand UO_396 (O_396,N_2943,N_2966);
and UO_397 (O_397,N_2954,N_2987);
or UO_398 (O_398,N_2940,N_2956);
and UO_399 (O_399,N_2947,N_2948);
nor UO_400 (O_400,N_2985,N_2970);
or UO_401 (O_401,N_2970,N_2976);
and UO_402 (O_402,N_2995,N_2975);
or UO_403 (O_403,N_2969,N_2988);
nor UO_404 (O_404,N_2972,N_2950);
and UO_405 (O_405,N_2990,N_2946);
and UO_406 (O_406,N_2942,N_2956);
nand UO_407 (O_407,N_2997,N_2978);
nor UO_408 (O_408,N_2999,N_2941);
and UO_409 (O_409,N_2952,N_2959);
nand UO_410 (O_410,N_2965,N_2991);
nand UO_411 (O_411,N_2953,N_2977);
or UO_412 (O_412,N_2982,N_2948);
and UO_413 (O_413,N_2955,N_2973);
or UO_414 (O_414,N_2986,N_2975);
and UO_415 (O_415,N_2954,N_2949);
nor UO_416 (O_416,N_2958,N_2986);
nand UO_417 (O_417,N_2994,N_2955);
and UO_418 (O_418,N_2959,N_2962);
or UO_419 (O_419,N_2999,N_2988);
or UO_420 (O_420,N_2954,N_2983);
nor UO_421 (O_421,N_2959,N_2944);
or UO_422 (O_422,N_2949,N_2993);
nor UO_423 (O_423,N_2976,N_2993);
and UO_424 (O_424,N_2951,N_2975);
and UO_425 (O_425,N_2942,N_2958);
nor UO_426 (O_426,N_2944,N_2968);
nand UO_427 (O_427,N_2999,N_2986);
and UO_428 (O_428,N_2956,N_2968);
nand UO_429 (O_429,N_2959,N_2986);
nand UO_430 (O_430,N_2943,N_2999);
or UO_431 (O_431,N_2984,N_2987);
nor UO_432 (O_432,N_2969,N_2940);
or UO_433 (O_433,N_2955,N_2976);
or UO_434 (O_434,N_2947,N_2978);
nor UO_435 (O_435,N_2955,N_2966);
nor UO_436 (O_436,N_2978,N_2945);
or UO_437 (O_437,N_2967,N_2997);
nand UO_438 (O_438,N_2942,N_2952);
nor UO_439 (O_439,N_2996,N_2956);
or UO_440 (O_440,N_2988,N_2997);
or UO_441 (O_441,N_2971,N_2987);
or UO_442 (O_442,N_2969,N_2945);
or UO_443 (O_443,N_2981,N_2980);
or UO_444 (O_444,N_2975,N_2966);
and UO_445 (O_445,N_2941,N_2992);
and UO_446 (O_446,N_2976,N_2987);
nor UO_447 (O_447,N_2978,N_2958);
nor UO_448 (O_448,N_2965,N_2963);
and UO_449 (O_449,N_2960,N_2992);
and UO_450 (O_450,N_2966,N_2951);
nor UO_451 (O_451,N_2996,N_2992);
nor UO_452 (O_452,N_2981,N_2943);
nor UO_453 (O_453,N_2942,N_2982);
nand UO_454 (O_454,N_2967,N_2948);
nand UO_455 (O_455,N_2941,N_2954);
and UO_456 (O_456,N_2991,N_2957);
nand UO_457 (O_457,N_2962,N_2956);
or UO_458 (O_458,N_2949,N_2962);
nor UO_459 (O_459,N_2966,N_2978);
nor UO_460 (O_460,N_2969,N_2984);
xor UO_461 (O_461,N_2988,N_2951);
nor UO_462 (O_462,N_2993,N_2992);
nand UO_463 (O_463,N_2955,N_2989);
or UO_464 (O_464,N_2984,N_2958);
or UO_465 (O_465,N_2997,N_2998);
nand UO_466 (O_466,N_2979,N_2970);
xnor UO_467 (O_467,N_2977,N_2979);
or UO_468 (O_468,N_2983,N_2985);
or UO_469 (O_469,N_2952,N_2979);
and UO_470 (O_470,N_2980,N_2955);
xnor UO_471 (O_471,N_2955,N_2944);
and UO_472 (O_472,N_2970,N_2974);
nand UO_473 (O_473,N_2988,N_2952);
nor UO_474 (O_474,N_2967,N_2956);
nand UO_475 (O_475,N_2959,N_2960);
nand UO_476 (O_476,N_2953,N_2960);
nand UO_477 (O_477,N_2959,N_2957);
and UO_478 (O_478,N_2941,N_2994);
nor UO_479 (O_479,N_2969,N_2993);
or UO_480 (O_480,N_2952,N_2965);
and UO_481 (O_481,N_2969,N_2960);
and UO_482 (O_482,N_2945,N_2981);
nor UO_483 (O_483,N_2989,N_2944);
or UO_484 (O_484,N_2995,N_2962);
and UO_485 (O_485,N_2961,N_2946);
and UO_486 (O_486,N_2971,N_2942);
or UO_487 (O_487,N_2981,N_2983);
nand UO_488 (O_488,N_2997,N_2940);
nand UO_489 (O_489,N_2963,N_2982);
nand UO_490 (O_490,N_2986,N_2951);
or UO_491 (O_491,N_2959,N_2972);
nor UO_492 (O_492,N_2943,N_2998);
or UO_493 (O_493,N_2940,N_2963);
nor UO_494 (O_494,N_2951,N_2957);
nor UO_495 (O_495,N_2951,N_2977);
and UO_496 (O_496,N_2973,N_2997);
nor UO_497 (O_497,N_2955,N_2998);
and UO_498 (O_498,N_2964,N_2994);
or UO_499 (O_499,N_2997,N_2989);
endmodule