module basic_1500_15000_2000_30_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1257,In_1064);
or U1 (N_1,In_1162,In_347);
or U2 (N_2,In_877,In_1316);
nand U3 (N_3,In_372,In_702);
and U4 (N_4,In_1336,In_549);
nand U5 (N_5,In_1118,In_1068);
xnor U6 (N_6,In_669,In_1281);
nand U7 (N_7,In_74,In_1279);
nand U8 (N_8,In_1361,In_381);
xor U9 (N_9,In_1368,In_162);
nand U10 (N_10,In_970,In_466);
nand U11 (N_11,In_493,In_1180);
nor U12 (N_12,In_979,In_86);
xor U13 (N_13,In_704,In_713);
nand U14 (N_14,In_849,In_1052);
or U15 (N_15,In_257,In_241);
or U16 (N_16,In_1049,In_606);
and U17 (N_17,In_777,In_760);
xnor U18 (N_18,In_734,In_277);
nor U19 (N_19,In_1110,In_487);
or U20 (N_20,In_1353,In_117);
xor U21 (N_21,In_327,In_525);
nand U22 (N_22,In_844,In_450);
xor U23 (N_23,In_716,In_12);
and U24 (N_24,In_216,In_628);
and U25 (N_25,In_1311,In_260);
and U26 (N_26,In_884,In_1307);
nor U27 (N_27,In_715,In_1053);
or U28 (N_28,In_664,In_977);
and U29 (N_29,In_682,In_1133);
nor U30 (N_30,In_133,In_1456);
and U31 (N_31,In_126,In_146);
and U32 (N_32,In_395,In_1481);
nor U33 (N_33,In_382,In_1009);
nand U34 (N_34,In_1117,In_1426);
and U35 (N_35,In_1337,In_784);
xnor U36 (N_36,In_168,In_489);
xor U37 (N_37,In_523,In_570);
and U38 (N_38,In_6,In_615);
nor U39 (N_39,In_703,In_272);
xor U40 (N_40,In_1200,In_1343);
or U41 (N_41,In_255,In_107);
xnor U42 (N_42,In_1192,In_891);
nand U43 (N_43,In_513,In_843);
or U44 (N_44,In_1472,In_828);
and U45 (N_45,In_1010,In_1402);
or U46 (N_46,In_9,In_1264);
nand U47 (N_47,In_616,In_826);
nand U48 (N_48,In_353,In_839);
and U49 (N_49,In_1225,In_1002);
nor U50 (N_50,In_573,In_797);
nand U51 (N_51,In_756,In_1342);
or U52 (N_52,In_90,In_1000);
and U53 (N_53,In_875,In_343);
nand U54 (N_54,In_534,In_1289);
or U55 (N_55,In_31,In_217);
and U56 (N_56,In_780,In_148);
and U57 (N_57,In_961,In_793);
or U58 (N_58,In_1242,In_403);
and U59 (N_59,In_1255,In_1288);
or U60 (N_60,In_1109,In_794);
nand U61 (N_61,In_1467,In_1172);
or U62 (N_62,In_253,In_219);
or U63 (N_63,In_1313,In_1135);
xnor U64 (N_64,In_655,In_215);
nand U65 (N_65,In_899,In_1143);
or U66 (N_66,In_663,In_1403);
xnor U67 (N_67,In_437,In_890);
nor U68 (N_68,In_1410,In_984);
nand U69 (N_69,In_490,In_1006);
or U70 (N_70,In_1360,In_366);
nor U71 (N_71,In_939,In_1465);
and U72 (N_72,In_973,In_122);
xor U73 (N_73,In_1186,In_385);
or U74 (N_74,In_1461,In_825);
and U75 (N_75,In_1114,In_1479);
and U76 (N_76,In_1260,In_532);
nor U77 (N_77,In_634,In_696);
or U78 (N_78,In_1454,In_1246);
and U79 (N_79,In_1483,In_313);
nor U80 (N_80,In_1325,In_701);
nor U81 (N_81,In_595,In_566);
and U82 (N_82,In_1005,In_76);
or U83 (N_83,In_907,In_562);
xor U84 (N_84,In_30,In_81);
nor U85 (N_85,In_1477,In_1161);
xnor U86 (N_86,In_789,In_312);
xor U87 (N_87,In_441,In_103);
or U88 (N_88,In_752,In_354);
or U89 (N_89,In_174,In_0);
xnor U90 (N_90,In_131,In_1160);
nand U91 (N_91,In_291,In_447);
and U92 (N_92,In_193,In_645);
and U93 (N_93,In_228,In_321);
nand U94 (N_94,In_496,In_1004);
nand U95 (N_95,In_1338,In_888);
nor U96 (N_96,In_350,In_252);
nor U97 (N_97,In_1333,In_709);
or U98 (N_98,In_720,In_738);
and U99 (N_99,In_1026,In_1462);
nor U100 (N_100,In_779,In_1072);
or U101 (N_101,In_932,In_273);
and U102 (N_102,In_809,In_1438);
nor U103 (N_103,In_908,In_344);
nand U104 (N_104,In_421,In_205);
nor U105 (N_105,In_603,In_914);
nor U106 (N_106,In_1443,In_1098);
xor U107 (N_107,In_19,In_317);
nor U108 (N_108,In_1491,In_1440);
xor U109 (N_109,In_1136,In_310);
nor U110 (N_110,In_432,In_998);
xor U111 (N_111,In_1156,In_36);
nor U112 (N_112,In_1344,In_765);
xnor U113 (N_113,In_1083,In_590);
and U114 (N_114,In_944,In_21);
or U115 (N_115,In_1398,In_725);
and U116 (N_116,In_1131,In_906);
nor U117 (N_117,In_1191,In_680);
xor U118 (N_118,In_771,In_1453);
nand U119 (N_119,In_1207,In_1210);
and U120 (N_120,In_1354,In_783);
nor U121 (N_121,In_316,In_1038);
xnor U122 (N_122,In_587,In_859);
nor U123 (N_123,In_499,In_922);
nand U124 (N_124,In_613,In_957);
and U125 (N_125,In_1113,In_807);
nand U126 (N_126,In_855,In_1022);
nand U127 (N_127,In_1074,In_1101);
nand U128 (N_128,In_504,In_1039);
xnor U129 (N_129,In_770,In_1229);
xnor U130 (N_130,In_279,In_142);
nand U131 (N_131,In_911,In_172);
and U132 (N_132,In_325,In_1201);
nand U133 (N_133,In_226,In_451);
xor U134 (N_134,In_512,In_431);
and U135 (N_135,In_1226,In_87);
nand U136 (N_136,In_185,In_1216);
and U137 (N_137,In_736,In_555);
xor U138 (N_138,In_70,In_82);
nand U139 (N_139,In_1065,In_218);
nand U140 (N_140,In_1094,In_851);
nand U141 (N_141,In_1014,In_15);
xor U142 (N_142,In_22,In_544);
nand U143 (N_143,In_341,In_258);
nor U144 (N_144,In_231,In_230);
or U145 (N_145,In_1017,In_547);
and U146 (N_146,In_1170,In_1315);
or U147 (N_147,In_73,In_369);
nand U148 (N_148,In_101,In_788);
and U149 (N_149,In_671,In_1271);
nor U150 (N_150,In_761,In_905);
xor U151 (N_151,In_163,In_1031);
nand U152 (N_152,In_274,In_44);
xor U153 (N_153,In_1405,In_471);
or U154 (N_154,In_975,In_636);
xnor U155 (N_155,In_189,In_654);
xor U156 (N_156,In_746,In_872);
nor U157 (N_157,In_108,In_278);
or U158 (N_158,In_198,In_619);
xor U159 (N_159,In_427,In_407);
or U160 (N_160,In_1495,In_340);
xnor U161 (N_161,In_1469,In_1097);
nand U162 (N_162,In_91,In_601);
or U163 (N_163,In_94,In_1243);
nand U164 (N_164,In_1308,In_717);
xor U165 (N_165,In_640,In_1046);
nand U166 (N_166,In_1449,In_208);
and U167 (N_167,In_743,In_237);
or U168 (N_168,In_904,In_857);
and U169 (N_169,In_1211,In_405);
xor U170 (N_170,In_1486,In_1339);
nand U171 (N_171,In_1450,In_1208);
xnor U172 (N_172,In_781,In_1287);
or U173 (N_173,In_1286,In_1394);
nand U174 (N_174,In_842,In_598);
or U175 (N_175,In_847,In_878);
nand U176 (N_176,In_585,In_753);
and U177 (N_177,In_666,In_591);
xor U178 (N_178,In_604,In_988);
xor U179 (N_179,In_283,In_652);
nor U180 (N_180,In_507,In_1250);
or U181 (N_181,In_1376,In_722);
nor U182 (N_182,In_229,In_1239);
and U183 (N_183,In_438,In_800);
nand U184 (N_184,In_79,In_302);
xor U185 (N_185,In_799,In_1050);
xnor U186 (N_186,In_649,In_1388);
nand U187 (N_187,In_990,In_120);
xor U188 (N_188,In_1066,In_428);
or U189 (N_189,In_225,In_1427);
nor U190 (N_190,In_1340,In_196);
nand U191 (N_191,In_635,In_178);
nor U192 (N_192,In_1298,In_220);
xor U193 (N_193,In_516,In_536);
xnor U194 (N_194,In_326,In_1051);
nor U195 (N_195,In_24,In_829);
nand U196 (N_196,In_778,In_731);
nor U197 (N_197,In_1367,In_668);
nand U198 (N_198,In_1032,In_84);
nor U199 (N_199,In_305,In_212);
xnor U200 (N_200,In_486,In_398);
or U201 (N_201,In_894,In_314);
and U202 (N_202,In_1396,In_768);
nand U203 (N_203,In_330,In_1409);
nor U204 (N_204,In_687,In_850);
nor U205 (N_205,In_695,In_488);
or U206 (N_206,In_1452,In_334);
xor U207 (N_207,In_1227,In_77);
and U208 (N_208,In_1302,In_1366);
or U209 (N_209,In_1122,In_600);
nand U210 (N_210,In_48,In_361);
xnor U211 (N_211,In_1375,In_1231);
xor U212 (N_212,In_651,In_764);
nand U213 (N_213,In_1103,In_589);
and U214 (N_214,In_759,In_389);
xor U215 (N_215,In_125,In_32);
xnor U216 (N_216,In_578,In_404);
and U217 (N_217,In_102,In_331);
and U218 (N_218,In_71,In_565);
nor U219 (N_219,In_1164,In_1327);
and U220 (N_220,In_1492,In_45);
nand U221 (N_221,In_785,In_266);
and U222 (N_222,In_430,In_690);
nand U223 (N_223,In_989,In_724);
xor U224 (N_224,In_1218,In_1324);
nor U225 (N_225,In_1067,In_397);
nand U226 (N_226,In_1124,In_62);
and U227 (N_227,In_1480,In_1259);
nand U228 (N_228,In_559,In_1334);
nor U229 (N_229,In_1235,In_714);
and U230 (N_230,In_527,In_502);
nor U231 (N_231,In_991,In_356);
nor U232 (N_232,In_897,In_1087);
xnor U233 (N_233,In_1464,In_1309);
and U234 (N_234,In_538,In_363);
or U235 (N_235,In_319,In_819);
nand U236 (N_236,In_864,In_608);
or U237 (N_237,In_235,In_966);
and U238 (N_238,In_199,In_1140);
xor U239 (N_239,In_706,In_236);
nand U240 (N_240,In_923,In_965);
or U241 (N_241,In_251,In_1252);
xor U242 (N_242,In_836,In_424);
nand U243 (N_243,In_662,In_835);
nor U244 (N_244,In_848,In_41);
and U245 (N_245,In_201,In_104);
and U246 (N_246,In_194,In_678);
or U247 (N_247,In_1152,In_295);
and U248 (N_248,In_811,In_109);
nor U249 (N_249,In_766,In_1176);
nor U250 (N_250,In_1416,In_942);
xnor U251 (N_251,In_883,In_357);
and U252 (N_252,In_1362,In_192);
or U253 (N_253,In_328,In_515);
or U254 (N_254,In_296,In_75);
nand U255 (N_255,In_698,In_386);
nand U256 (N_256,In_881,In_1439);
nand U257 (N_257,In_453,In_263);
xnor U258 (N_258,In_337,In_1173);
nor U259 (N_259,In_834,In_898);
nand U260 (N_260,In_648,In_1267);
nand U261 (N_261,In_1137,In_1015);
and U262 (N_262,In_463,In_1434);
nand U263 (N_263,In_1433,In_1436);
nor U264 (N_264,In_1071,In_469);
nand U265 (N_265,In_54,In_1193);
xnor U266 (N_266,In_733,In_594);
nor U267 (N_267,In_983,In_978);
nor U268 (N_268,In_1330,In_621);
or U269 (N_269,In_1442,In_358);
xor U270 (N_270,In_1085,In_1059);
and U271 (N_271,In_896,In_1301);
xor U272 (N_272,In_599,In_1012);
xor U273 (N_273,In_996,In_744);
nor U274 (N_274,In_1323,In_741);
and U275 (N_275,In_1157,In_1035);
xor U276 (N_276,In_1299,In_400);
and U277 (N_277,In_392,In_29);
or U278 (N_278,In_452,In_845);
or U279 (N_279,In_412,In_670);
nor U280 (N_280,In_1418,In_1300);
or U281 (N_281,In_611,In_958);
and U282 (N_282,In_946,In_554);
nand U283 (N_283,In_98,In_203);
or U284 (N_284,In_63,In_658);
nor U285 (N_285,In_728,In_380);
nand U286 (N_286,In_1003,In_1168);
and U287 (N_287,In_1223,In_823);
nand U288 (N_288,In_415,In_1273);
or U289 (N_289,In_647,In_1189);
or U290 (N_290,In_239,In_976);
xnor U291 (N_291,In_1188,In_458);
and U292 (N_292,In_169,In_339);
xor U293 (N_293,In_1370,In_1319);
xnor U294 (N_294,In_1013,In_188);
xnor U295 (N_295,In_541,In_88);
nand U296 (N_296,In_1034,In_822);
nand U297 (N_297,In_200,In_900);
xor U298 (N_298,In_256,In_1149);
nand U299 (N_299,In_1322,In_533);
or U300 (N_300,In_726,In_987);
or U301 (N_301,In_1057,In_749);
nand U302 (N_302,In_446,In_917);
nor U303 (N_303,In_1373,In_521);
nor U304 (N_304,In_1146,In_1238);
or U305 (N_305,In_1384,In_1248);
and U306 (N_306,In_1202,In_299);
nor U307 (N_307,In_986,In_1455);
nand U308 (N_308,In_1318,In_1147);
xor U309 (N_309,In_1305,In_1033);
nor U310 (N_310,In_1167,In_627);
and U311 (N_311,In_941,In_755);
xnor U312 (N_312,In_1431,In_40);
xnor U313 (N_313,In_439,In_249);
nor U314 (N_314,In_892,In_754);
or U315 (N_315,In_1247,In_1044);
nand U316 (N_316,In_85,In_876);
and U317 (N_317,In_1116,In_1215);
nor U318 (N_318,In_355,In_1023);
nor U319 (N_319,In_113,In_1422);
nand U320 (N_320,In_1030,In_360);
nand U321 (N_321,In_186,In_478);
xnor U322 (N_322,In_110,In_1310);
xor U323 (N_323,In_425,In_121);
and U324 (N_324,In_423,In_1179);
nand U325 (N_325,In_213,In_336);
or U326 (N_326,In_592,In_831);
xnor U327 (N_327,In_1292,In_391);
xor U328 (N_328,In_92,In_481);
xnor U329 (N_329,In_1488,In_732);
nand U330 (N_330,In_535,In_602);
and U331 (N_331,In_1185,In_948);
or U332 (N_332,In_903,In_920);
nor U333 (N_333,In_653,In_177);
xor U334 (N_334,In_1141,In_265);
and U335 (N_335,In_4,In_1056);
and U336 (N_336,In_51,In_545);
and U337 (N_337,In_1007,In_477);
nor U338 (N_338,In_1236,In_820);
nand U339 (N_339,In_919,In_959);
nor U340 (N_340,In_322,In_1446);
and U341 (N_341,In_967,In_963);
nor U342 (N_342,In_596,In_1391);
or U343 (N_343,In_164,In_1417);
xor U344 (N_344,In_53,In_1233);
nand U345 (N_345,In_871,In_115);
nor U346 (N_346,In_1275,In_727);
nand U347 (N_347,In_1401,In_1159);
nor U348 (N_348,In_65,In_1352);
nand U349 (N_349,In_303,In_762);
and U350 (N_350,In_867,In_588);
nand U351 (N_351,In_1036,In_461);
or U352 (N_352,In_1198,In_1349);
and U353 (N_353,In_1256,In_1237);
or U354 (N_354,In_1195,In_183);
and U355 (N_355,In_558,In_1425);
nand U356 (N_356,In_491,In_1341);
nand U357 (N_357,In_748,In_971);
or U358 (N_358,In_83,In_1241);
nor U359 (N_359,In_982,In_569);
and U360 (N_360,In_1441,In_1285);
xor U361 (N_361,In_1411,In_124);
and U362 (N_362,In_750,In_1213);
nor U363 (N_363,In_1214,In_500);
or U364 (N_364,In_1385,In_479);
nand U365 (N_365,In_681,In_1395);
and U366 (N_366,In_1084,In_633);
nand U367 (N_367,In_1016,In_775);
xnor U368 (N_368,In_817,In_721);
xor U369 (N_369,In_1011,In_112);
xor U370 (N_370,In_384,In_557);
or U371 (N_371,In_1008,In_1364);
or U372 (N_372,In_1304,In_442);
xnor U373 (N_373,In_773,In_1382);
xor U374 (N_374,In_35,In_868);
nand U375 (N_375,In_1054,In_1263);
and U376 (N_376,In_563,In_1268);
and U377 (N_377,In_248,In_292);
and U378 (N_378,In_1144,In_1169);
or U379 (N_379,In_806,In_1478);
or U380 (N_380,In_786,In_259);
nand U381 (N_381,In_42,In_16);
nand U382 (N_382,In_1348,In_915);
and U383 (N_383,In_324,In_846);
and U384 (N_384,In_1108,In_333);
nor U385 (N_385,In_1206,In_969);
or U386 (N_386,In_134,In_832);
and U387 (N_387,In_1493,In_1069);
xnor U388 (N_388,In_1412,In_548);
nor U389 (N_389,In_980,In_556);
or U390 (N_390,In_1445,In_69);
and U391 (N_391,In_539,In_307);
nand U392 (N_392,In_1269,In_705);
nand U393 (N_393,In_282,In_329);
nand U394 (N_394,In_1086,In_393);
nor U395 (N_395,In_723,In_1166);
nor U396 (N_396,In_184,In_508);
nor U397 (N_397,In_390,In_297);
and U398 (N_398,In_546,In_351);
nand U399 (N_399,In_947,In_729);
nand U400 (N_400,In_830,In_1404);
nor U401 (N_401,In_805,In_742);
nor U402 (N_402,In_1457,In_1119);
and U403 (N_403,In_204,In_238);
xnor U404 (N_404,In_1386,In_206);
xnor U405 (N_405,In_926,In_901);
xor U406 (N_406,In_1048,In_190);
nor U407 (N_407,In_694,In_1475);
xor U408 (N_408,In_456,In_93);
and U409 (N_409,In_105,In_804);
and U410 (N_410,In_20,In_250);
xor U411 (N_411,In_129,In_943);
nand U412 (N_412,In_462,In_476);
nand U413 (N_413,In_882,In_1463);
or U414 (N_414,In_1165,In_243);
nand U415 (N_415,In_61,In_99);
xnor U416 (N_416,In_795,In_1484);
nand U417 (N_417,In_568,In_609);
nand U418 (N_418,In_197,In_306);
or U419 (N_419,In_156,In_885);
nor U420 (N_420,In_1027,In_1374);
and U421 (N_421,In_1400,In_684);
nand U422 (N_422,In_1096,In_473);
xnor U423 (N_423,In_365,In_1181);
nor U424 (N_424,In_1219,In_676);
nor U425 (N_425,In_614,In_787);
or U426 (N_426,In_52,In_1199);
nand U427 (N_427,In_264,In_457);
nor U428 (N_428,In_246,In_950);
nor U429 (N_429,In_1099,In_100);
and U430 (N_430,In_1024,In_1055);
xor U431 (N_431,In_509,In_1230);
nor U432 (N_432,In_1280,In_1204);
or U433 (N_433,In_497,In_1081);
and U434 (N_434,In_449,In_593);
and U435 (N_435,In_1134,In_95);
nor U436 (N_436,In_345,In_464);
nand U437 (N_437,In_537,In_1487);
or U438 (N_438,In_149,In_1496);
and U439 (N_439,In_1217,In_1);
nor U440 (N_440,In_1019,In_1102);
nand U441 (N_441,In_170,In_791);
or U442 (N_442,In_529,In_997);
nand U443 (N_443,In_673,In_1092);
xor U444 (N_444,In_840,In_949);
nand U445 (N_445,In_1490,In_78);
xor U446 (N_446,In_860,In_276);
or U447 (N_447,In_782,In_414);
and U448 (N_448,In_1419,In_1132);
xor U449 (N_449,In_503,In_550);
xnor U450 (N_450,In_342,In_1332);
nand U451 (N_451,In_1451,In_1088);
nor U452 (N_452,In_992,In_567);
nand U453 (N_453,In_1460,In_56);
xor U454 (N_454,In_518,In_17);
or U455 (N_455,In_1345,In_597);
nor U456 (N_456,In_774,In_271);
nor U457 (N_457,In_1320,In_422);
xnor U458 (N_458,In_13,In_1107);
or U459 (N_459,In_1407,In_612);
nand U460 (N_460,In_359,In_1177);
nand U461 (N_461,In_1129,In_68);
nor U462 (N_462,In_222,In_419);
nor U463 (N_463,In_543,In_1497);
nor U464 (N_464,In_1234,In_1029);
xnor U465 (N_465,In_1205,In_1078);
or U466 (N_466,In_165,In_798);
xnor U467 (N_467,In_610,In_175);
xnor U468 (N_468,In_1379,In_1314);
or U469 (N_469,In_388,In_889);
xor U470 (N_470,In_39,In_368);
and U471 (N_471,In_1155,In_893);
nor U472 (N_472,In_1125,In_3);
or U473 (N_473,In_952,In_1355);
nor U474 (N_474,In_644,In_37);
nand U475 (N_475,In_571,In_1100);
and U476 (N_476,In_155,In_994);
nor U477 (N_477,In_176,In_38);
xor U478 (N_478,In_1414,In_288);
nor U479 (N_479,In_145,In_1282);
and U480 (N_480,In_929,In_261);
and U481 (N_481,In_650,In_909);
or U482 (N_482,In_298,In_679);
and U483 (N_483,In_924,In_114);
nand U484 (N_484,In_553,In_583);
nor U485 (N_485,In_1190,In_376);
and U486 (N_486,In_300,In_123);
nand U487 (N_487,In_1251,In_524);
nand U488 (N_488,In_711,In_551);
xor U489 (N_489,In_617,In_993);
nor U490 (N_490,In_910,In_116);
xor U491 (N_491,In_667,In_335);
xnor U492 (N_492,In_181,In_945);
nor U493 (N_493,In_699,In_852);
xnor U494 (N_494,In_60,In_1221);
and U495 (N_495,In_1197,In_1042);
nand U496 (N_496,In_1021,In_304);
nand U497 (N_497,In_769,In_710);
and U498 (N_498,In_352,In_269);
xor U499 (N_499,In_1145,In_375);
or U500 (N_500,In_492,In_519);
xnor U501 (N_501,In_1277,In_232);
xor U502 (N_502,N_116,N_32);
nand U503 (N_503,N_80,N_74);
nand U504 (N_504,N_371,In_933);
or U505 (N_505,N_81,In_1430);
nor U506 (N_506,In_1060,N_369);
or U507 (N_507,N_491,In_1112);
nor U508 (N_508,In_254,N_338);
nand U509 (N_509,In_171,In_758);
or U510 (N_510,In_227,N_394);
or U511 (N_511,In_962,In_281);
or U512 (N_512,N_378,In_526);
nor U513 (N_513,In_1111,In_1474);
and U514 (N_514,N_155,N_275);
xnor U515 (N_515,N_319,N_277);
xnor U516 (N_516,In_607,N_263);
nand U517 (N_517,N_99,In_373);
and U518 (N_518,In_130,In_402);
nand U519 (N_519,In_1130,N_17);
nand U520 (N_520,In_26,N_484);
nor U521 (N_521,In_1494,N_247);
nor U522 (N_522,N_434,N_210);
or U523 (N_523,N_309,N_38);
nor U524 (N_524,N_442,N_269);
nor U525 (N_525,In_1075,N_224);
nor U526 (N_526,In_801,N_153);
nor U527 (N_527,In_494,In_584);
nand U528 (N_528,N_383,In_154);
and U529 (N_529,In_72,N_53);
nor U530 (N_530,In_1389,In_1466);
or U531 (N_531,In_426,N_284);
and U532 (N_532,In_879,N_102);
or U533 (N_533,In_28,In_498);
nand U534 (N_534,N_315,In_688);
and U535 (N_535,N_202,In_311);
nor U536 (N_536,In_139,N_447);
xnor U537 (N_537,N_310,In_144);
and U538 (N_538,N_429,In_1183);
or U539 (N_539,In_1148,N_470);
nand U540 (N_540,N_301,In_1306);
nor U541 (N_541,In_790,In_665);
or U542 (N_542,N_415,In_1377);
xor U543 (N_543,N_352,In_240);
or U544 (N_544,N_449,In_718);
nand U545 (N_545,N_300,N_316);
xnor U546 (N_546,In_913,In_863);
and U547 (N_547,N_425,In_895);
nor U548 (N_548,N_493,In_140);
or U549 (N_549,N_193,In_854);
xor U550 (N_550,N_10,In_861);
and U551 (N_551,N_201,N_250);
xor U552 (N_552,N_313,In_1171);
nor U553 (N_553,N_173,N_452);
xor U554 (N_554,In_912,In_1061);
xnor U555 (N_555,N_483,N_402);
nor U556 (N_556,In_33,N_114);
nand U557 (N_557,In_173,In_1358);
xor U558 (N_558,N_298,In_67);
nand U559 (N_559,N_437,In_46);
nor U560 (N_560,N_262,In_159);
or U561 (N_561,In_520,In_865);
nand U562 (N_562,In_1458,N_289);
nor U563 (N_563,In_294,In_1079);
or U564 (N_564,In_686,N_137);
and U565 (N_565,N_264,N_171);
xor U566 (N_566,N_374,In_1328);
or U567 (N_567,N_189,N_51);
or U568 (N_568,In_182,In_887);
nand U569 (N_569,In_1104,N_459);
and U570 (N_570,N_65,In_564);
nor U571 (N_571,N_227,In_833);
or U572 (N_572,N_121,N_13);
nor U573 (N_573,In_1115,In_951);
xnor U574 (N_574,In_406,N_100);
or U575 (N_575,In_309,In_1187);
or U576 (N_576,N_200,N_311);
nor U577 (N_577,N_477,N_400);
and U578 (N_578,N_329,In_692);
and U579 (N_579,In_938,In_370);
xor U580 (N_580,N_8,In_136);
nor U581 (N_581,In_873,N_205);
xor U582 (N_582,N_290,In_377);
xnor U583 (N_583,N_337,In_118);
or U584 (N_584,N_265,N_236);
nor U585 (N_585,N_478,In_1232);
nand U586 (N_586,In_286,In_1356);
and U587 (N_587,N_27,N_197);
nor U588 (N_588,In_1106,In_626);
or U589 (N_589,N_3,N_398);
xor U590 (N_590,N_128,In_880);
or U591 (N_591,N_7,In_632);
nor U592 (N_592,In_866,N_186);
nor U593 (N_593,N_397,In_1142);
nor U594 (N_594,N_14,In_960);
nor U595 (N_595,N_431,N_382);
nand U596 (N_596,In_210,In_956);
nand U597 (N_597,N_444,In_1154);
xor U598 (N_598,In_1347,N_416);
nor U599 (N_599,In_55,In_964);
nand U600 (N_600,N_448,In_436);
xor U601 (N_601,N_423,N_462);
xnor U602 (N_602,N_390,N_59);
or U603 (N_603,N_246,In_1076);
xnor U604 (N_604,In_1138,In_763);
and U605 (N_605,In_981,In_1399);
or U606 (N_606,In_1043,N_77);
and U607 (N_607,In_1392,N_208);
and U608 (N_608,In_1018,In_1435);
and U609 (N_609,N_76,In_572);
and U610 (N_610,N_258,N_238);
and U611 (N_611,In_25,N_362);
nand U612 (N_612,In_517,In_89);
nor U613 (N_613,N_465,In_936);
and U614 (N_614,In_501,N_36);
nand U615 (N_615,N_97,N_133);
nor U616 (N_616,In_49,N_92);
and U617 (N_617,N_156,In_815);
xnor U618 (N_618,In_1120,N_367);
or U619 (N_619,In_1224,N_123);
nor U620 (N_620,N_174,N_216);
and U621 (N_621,N_21,In_708);
and U622 (N_622,N_451,N_405);
or U623 (N_623,N_379,N_359);
xnor U624 (N_624,N_120,N_242);
nand U625 (N_625,N_450,In_674);
and U626 (N_626,In_582,In_772);
nor U627 (N_627,N_281,N_468);
nor U628 (N_628,In_1139,N_222);
xnor U629 (N_629,In_379,N_190);
xor U630 (N_630,In_459,In_1413);
and U631 (N_631,N_487,In_1397);
and U632 (N_632,N_165,N_341);
or U633 (N_633,N_419,In_158);
xor U634 (N_634,In_1473,N_119);
xor U635 (N_635,In_1274,N_333);
and U636 (N_636,In_1262,In_1093);
nand U637 (N_637,In_638,In_480);
and U638 (N_638,In_646,In_1062);
nand U639 (N_639,In_374,In_207);
or U640 (N_640,N_296,In_167);
nand U641 (N_641,N_6,In_510);
nor U642 (N_642,N_260,In_1447);
nor U643 (N_643,N_293,N_71);
and U644 (N_644,N_261,N_385);
nand U645 (N_645,N_220,N_166);
nor U646 (N_646,In_1359,In_1203);
or U647 (N_647,In_1499,In_1128);
and U648 (N_648,In_267,N_228);
and U649 (N_649,In_869,In_625);
xor U650 (N_650,N_170,N_182);
xnor U651 (N_651,In_972,In_1365);
nor U652 (N_652,In_474,N_375);
nor U653 (N_653,N_469,In_1432);
nor U654 (N_654,N_117,N_373);
nor U655 (N_655,In_1346,N_443);
nor U656 (N_656,N_203,In_1258);
nand U657 (N_657,In_530,In_1182);
or U658 (N_658,In_467,N_388);
nand U659 (N_659,N_157,N_178);
nand U660 (N_660,In_856,N_164);
xnor U661 (N_661,N_302,In_221);
and U662 (N_662,In_34,In_1089);
nor U663 (N_663,In_802,In_577);
nor U664 (N_664,In_410,N_215);
nor U665 (N_665,In_2,N_94);
nand U666 (N_666,In_433,In_349);
and U667 (N_667,In_808,In_47);
nand U668 (N_668,In_135,In_270);
and U669 (N_669,In_576,N_172);
nand U670 (N_670,In_338,N_50);
nor U671 (N_671,N_295,N_66);
or U672 (N_672,N_145,In_1228);
and U673 (N_673,In_151,In_66);
nor U674 (N_674,In_858,In_862);
nor U675 (N_675,In_1240,In_1001);
nand U676 (N_676,In_242,In_1123);
and U677 (N_677,In_1082,N_62);
nand U678 (N_678,N_494,In_11);
xnor U679 (N_679,In_472,In_1184);
nor U680 (N_680,In_816,In_1293);
or U681 (N_681,In_886,N_254);
and U682 (N_682,N_492,N_144);
nor U683 (N_683,In_629,In_106);
xor U684 (N_684,N_141,In_739);
xnor U685 (N_685,N_357,N_18);
and U686 (N_686,In_1424,In_730);
nand U687 (N_687,In_138,In_401);
xor U688 (N_688,In_58,N_499);
nor U689 (N_689,In_1270,In_659);
or U690 (N_690,N_115,N_372);
xor U691 (N_691,N_251,In_641);
xnor U692 (N_692,In_792,In_751);
nand U693 (N_693,In_1423,In_1459);
or U694 (N_694,In_693,N_328);
xnor U695 (N_695,N_433,In_1266);
and U696 (N_696,In_1150,In_928);
xnor U697 (N_697,In_1178,N_486);
or U698 (N_698,N_24,In_1470);
nand U699 (N_699,In_202,N_321);
xnor U700 (N_700,N_111,N_95);
xor U701 (N_701,N_196,N_435);
nand U702 (N_702,In_1291,N_47);
nor U703 (N_703,In_293,N_54);
and U704 (N_704,N_5,N_386);
or U705 (N_705,N_317,N_88);
and U706 (N_706,N_461,In_657);
nor U707 (N_707,In_1244,N_48);
nand U708 (N_708,In_935,N_140);
nor U709 (N_709,In_179,In_841);
or U710 (N_710,N_9,N_85);
nor U711 (N_711,N_93,N_473);
xnor U712 (N_712,N_314,In_1153);
and U713 (N_713,In_191,In_639);
nand U714 (N_714,N_253,N_346);
nand U715 (N_715,N_343,N_0);
xnor U716 (N_716,N_413,N_240);
and U717 (N_717,In_418,N_113);
xor U718 (N_718,N_199,N_482);
nand U719 (N_719,N_411,N_29);
xor U720 (N_720,N_475,In_137);
nor U721 (N_721,In_5,N_219);
and U722 (N_722,In_127,N_446);
or U723 (N_723,N_306,In_707);
and U724 (N_724,In_417,N_55);
and U725 (N_725,In_1489,N_244);
nor U726 (N_726,N_4,N_72);
nand U727 (N_727,N_154,N_368);
and U728 (N_728,N_312,N_334);
nor U729 (N_729,In_18,In_1429);
nand U730 (N_730,N_125,N_331);
and U731 (N_731,N_282,N_332);
and U732 (N_732,In_396,In_735);
nor U733 (N_733,N_351,In_399);
or U734 (N_734,In_1028,N_287);
or U735 (N_735,N_424,N_392);
nor U736 (N_736,In_1276,In_289);
and U737 (N_737,In_579,N_252);
nand U738 (N_738,N_107,N_151);
xor U739 (N_739,In_111,N_37);
nand U740 (N_740,In_371,N_396);
xnor U741 (N_741,In_870,In_1312);
or U742 (N_742,In_747,In_1321);
and U743 (N_743,N_432,N_83);
nor U744 (N_744,In_50,N_11);
nor U745 (N_745,In_280,In_318);
nand U746 (N_746,N_68,N_230);
nand U747 (N_747,In_482,N_105);
or U748 (N_748,In_362,N_335);
or U749 (N_749,In_642,In_1294);
or U750 (N_750,In_1468,N_195);
xnor U751 (N_751,N_270,In_506);
or U752 (N_752,In_812,In_367);
nand U753 (N_753,N_35,In_180);
nand U754 (N_754,In_287,In_244);
nor U755 (N_755,In_1378,N_112);
nand U756 (N_756,N_403,N_428);
nand U757 (N_757,In_814,N_498);
nand U758 (N_758,In_1220,In_245);
nand U759 (N_759,In_153,In_1393);
nor U760 (N_760,In_64,N_322);
or U761 (N_761,In_59,N_198);
or U762 (N_762,In_630,N_146);
xnor U763 (N_763,N_61,N_279);
and U764 (N_764,N_129,In_689);
nand U765 (N_765,In_620,In_618);
nand U766 (N_766,N_417,In_1070);
xnor U767 (N_767,N_214,In_1045);
xor U768 (N_768,In_285,N_348);
nor U769 (N_769,In_1380,In_460);
nand U770 (N_770,In_685,N_28);
xor U771 (N_771,N_30,N_56);
nand U772 (N_772,In_1063,N_350);
nor U773 (N_773,In_902,N_234);
nand U774 (N_774,N_466,In_187);
nand U775 (N_775,In_416,N_122);
and U776 (N_776,In_455,In_1387);
or U777 (N_777,In_315,N_180);
and U778 (N_778,N_90,In_1209);
nand U779 (N_779,N_285,In_1091);
and U780 (N_780,N_118,In_1303);
or U781 (N_781,In_995,In_838);
and U782 (N_782,In_465,In_1278);
and U783 (N_783,N_267,In_1290);
nand U784 (N_784,N_496,N_381);
and U785 (N_785,N_176,N_278);
and U786 (N_786,N_58,In_767);
nor U787 (N_787,N_57,In_672);
xor U788 (N_788,In_1297,In_697);
and U789 (N_789,In_408,In_435);
and U790 (N_790,In_1383,N_366);
xor U791 (N_791,N_126,N_330);
nor U792 (N_792,N_420,In_1381);
xor U793 (N_793,In_346,N_22);
and U794 (N_794,N_365,In_209);
or U795 (N_795,N_349,N_231);
nor U796 (N_796,In_1476,In_1420);
nand U797 (N_797,N_187,N_454);
and U798 (N_798,N_307,In_737);
nor U799 (N_799,In_1127,N_464);
or U800 (N_800,In_1025,N_471);
nand U801 (N_801,In_757,N_438);
nor U802 (N_802,In_968,N_393);
or U803 (N_803,N_163,N_336);
xor U804 (N_804,In_937,N_2);
nor U805 (N_805,N_142,N_147);
nor U806 (N_806,N_63,N_25);
or U807 (N_807,In_444,In_387);
and U808 (N_808,N_256,N_213);
xnor U809 (N_809,In_128,In_1194);
and U810 (N_810,N_401,N_280);
or U811 (N_811,N_266,N_64);
or U812 (N_812,N_138,N_422);
nand U813 (N_813,N_456,N_354);
nand U814 (N_814,In_1212,N_179);
nor U815 (N_815,In_586,In_119);
or U816 (N_816,N_271,In_195);
or U817 (N_817,In_552,N_42);
nor U818 (N_818,In_1317,N_273);
nand U819 (N_819,In_1174,N_152);
and U820 (N_820,N_481,In_745);
and U821 (N_821,N_23,N_288);
xor U822 (N_822,In_1126,N_325);
xnor U823 (N_823,N_212,In_1261);
nor U824 (N_824,In_930,N_237);
nand U825 (N_825,N_223,N_421);
and U826 (N_826,In_1371,In_23);
nor U827 (N_827,N_497,In_1329);
nand U828 (N_828,In_383,In_1080);
or U829 (N_829,N_84,N_218);
and U830 (N_830,N_124,N_460);
xnor U831 (N_831,In_623,N_407);
and U832 (N_832,N_356,In_1406);
or U833 (N_833,N_41,N_160);
xnor U834 (N_834,N_327,In_1357);
and U835 (N_835,N_360,In_409);
nand U836 (N_836,N_130,In_953);
and U837 (N_837,In_96,In_1408);
nor U838 (N_838,In_443,N_490);
and U839 (N_839,In_813,In_824);
and U840 (N_840,In_7,In_147);
or U841 (N_841,N_131,N_347);
or U842 (N_842,In_214,N_31);
nor U843 (N_843,In_580,N_225);
nor U844 (N_844,In_853,N_355);
nand U845 (N_845,N_318,In_1498);
nor U846 (N_846,N_206,N_184);
nand U847 (N_847,In_348,N_323);
and U848 (N_848,N_132,N_409);
nand U849 (N_849,N_60,N_221);
nand U850 (N_850,In_80,N_15);
nand U851 (N_851,N_134,N_363);
and U852 (N_852,In_157,N_489);
and U853 (N_853,In_448,In_332);
and U854 (N_854,In_1296,N_217);
and U855 (N_855,N_19,In_284);
or U856 (N_856,N_274,In_660);
or U857 (N_857,In_1095,N_418);
nand U858 (N_858,N_387,In_624);
nor U859 (N_859,N_159,In_301);
and U860 (N_860,In_1326,In_740);
or U861 (N_861,N_297,In_542);
and U862 (N_862,In_776,In_1272);
and U863 (N_863,N_391,N_79);
nor U864 (N_864,N_430,N_283);
and U865 (N_865,N_457,N_412);
or U866 (N_866,In_954,In_560);
nor U867 (N_867,In_925,N_168);
nand U868 (N_868,N_175,N_226);
nor U869 (N_869,N_148,N_135);
nand U870 (N_870,In_622,In_656);
xnor U871 (N_871,N_479,N_384);
or U872 (N_872,N_320,N_404);
xnor U873 (N_873,N_272,In_511);
xor U874 (N_874,In_1363,N_162);
or U875 (N_875,In_675,In_161);
or U876 (N_876,In_1421,In_1283);
nand U877 (N_877,In_308,N_103);
nor U878 (N_878,In_561,In_268);
xor U879 (N_879,In_43,In_57);
xor U880 (N_880,In_927,N_345);
nand U881 (N_881,N_139,N_476);
nand U882 (N_882,N_257,N_149);
nand U883 (N_883,N_67,In_837);
nand U884 (N_884,In_97,N_45);
and U885 (N_885,N_427,In_1369);
nor U886 (N_886,N_467,In_683);
xnor U887 (N_887,N_33,N_229);
or U888 (N_888,N_110,N_395);
nand U889 (N_889,N_1,In_150);
and U890 (N_890,In_1037,In_700);
and U891 (N_891,N_440,N_75);
nor U892 (N_892,In_152,In_827);
nor U893 (N_893,N_191,N_408);
nor U894 (N_894,In_1265,In_874);
xor U895 (N_895,N_188,In_323);
xor U896 (N_896,In_429,N_304);
nand U897 (N_897,In_275,N_445);
xor U898 (N_898,In_1428,In_141);
and U899 (N_899,In_378,N_495);
or U900 (N_900,N_364,In_434);
nand U901 (N_901,N_453,N_108);
xnor U902 (N_902,N_339,In_411);
and U903 (N_903,In_528,N_361);
xnor U904 (N_904,In_712,N_291);
and U905 (N_905,N_44,In_661);
nand U906 (N_906,In_796,N_43);
and U907 (N_907,In_918,In_505);
or U908 (N_908,In_1058,In_1351);
or U909 (N_909,N_485,N_52);
nand U910 (N_910,N_104,N_249);
nor U911 (N_911,N_358,N_16);
nor U912 (N_912,N_89,In_1390);
nor U913 (N_913,N_324,N_399);
xor U914 (N_914,N_211,N_239);
xnor U915 (N_915,N_167,N_294);
and U916 (N_916,N_241,In_440);
xnor U917 (N_917,N_39,In_27);
and U918 (N_918,In_1151,N_370);
nand U919 (N_919,In_1196,N_474);
nand U920 (N_920,In_233,In_921);
nand U921 (N_921,In_1437,N_169);
and U922 (N_922,N_87,In_290);
nand U923 (N_923,In_10,In_637);
nand U924 (N_924,In_211,N_158);
or U925 (N_925,In_320,N_410);
and U926 (N_926,N_380,In_1372);
nand U927 (N_927,In_420,In_1284);
or U928 (N_928,N_305,In_8);
nor U929 (N_929,N_276,In_810);
or U930 (N_930,N_73,In_522);
and U931 (N_931,N_480,In_575);
nand U932 (N_932,N_20,N_342);
nand U933 (N_933,In_166,N_243);
xnor U934 (N_934,N_150,N_248);
nor U935 (N_935,In_14,In_475);
nand U936 (N_936,In_1253,N_69);
xor U937 (N_937,In_234,N_82);
or U938 (N_938,In_1163,In_1415);
nor U939 (N_939,In_1158,In_468);
xor U940 (N_940,In_364,In_1482);
nand U941 (N_941,N_49,In_1020);
nand U942 (N_942,In_143,N_183);
nand U943 (N_943,N_299,In_224);
nand U944 (N_944,N_488,N_255);
xor U945 (N_945,N_232,N_441);
or U946 (N_946,N_233,N_101);
nand U947 (N_947,N_376,N_34);
xnor U948 (N_948,N_177,N_245);
or U949 (N_949,N_472,In_1444);
nor U950 (N_950,In_719,In_931);
nor U951 (N_951,In_514,In_934);
xor U952 (N_952,N_12,N_344);
or U953 (N_953,N_127,In_540);
or U954 (N_954,N_463,N_70);
nand U955 (N_955,N_109,In_631);
nor U956 (N_956,In_484,In_916);
xor U957 (N_957,In_413,In_1350);
or U958 (N_958,N_209,In_1073);
xor U959 (N_959,N_91,N_181);
and U960 (N_960,In_483,N_194);
and U961 (N_961,In_1040,In_495);
and U962 (N_962,N_259,N_143);
nand U963 (N_963,N_426,N_377);
or U964 (N_964,In_677,N_303);
or U965 (N_965,In_531,In_247);
xor U966 (N_966,In_394,N_98);
and U967 (N_967,In_1105,N_458);
xnor U968 (N_968,N_106,N_235);
xor U969 (N_969,N_292,In_1047);
or U970 (N_970,In_574,N_455);
nand U971 (N_971,In_1471,In_470);
nor U972 (N_972,N_326,In_454);
xor U973 (N_973,In_1041,In_1295);
xor U974 (N_974,In_1331,In_445);
nand U975 (N_975,N_286,In_1077);
nor U976 (N_976,N_340,In_1090);
or U977 (N_977,In_1485,N_96);
or U978 (N_978,N_353,In_160);
xnor U979 (N_979,In_132,In_985);
xor U980 (N_980,In_974,In_643);
xor U981 (N_981,In_1335,N_439);
nand U982 (N_982,In_223,N_26);
and U983 (N_983,N_204,N_406);
nand U984 (N_984,N_436,N_414);
xor U985 (N_985,In_1245,In_1175);
nand U986 (N_986,In_955,In_1121);
xor U987 (N_987,In_1254,N_46);
nor U988 (N_988,N_136,In_485);
nor U989 (N_989,N_40,In_1222);
or U990 (N_990,In_1249,In_818);
xor U991 (N_991,N_78,In_605);
or U992 (N_992,In_691,N_207);
xor U993 (N_993,N_389,N_161);
nand U994 (N_994,N_185,In_581);
nand U995 (N_995,In_1448,In_821);
nand U996 (N_996,N_268,In_262);
nand U997 (N_997,In_940,N_86);
nand U998 (N_998,In_999,In_803);
nor U999 (N_999,N_308,N_192);
nor U1000 (N_1000,N_955,N_983);
and U1001 (N_1001,N_913,N_799);
xnor U1002 (N_1002,N_851,N_641);
nor U1003 (N_1003,N_823,N_790);
nor U1004 (N_1004,N_747,N_727);
or U1005 (N_1005,N_758,N_996);
xor U1006 (N_1006,N_662,N_699);
nand U1007 (N_1007,N_909,N_872);
nor U1008 (N_1008,N_785,N_515);
and U1009 (N_1009,N_791,N_868);
nor U1010 (N_1010,N_682,N_952);
nand U1011 (N_1011,N_653,N_689);
or U1012 (N_1012,N_992,N_899);
or U1013 (N_1013,N_576,N_776);
or U1014 (N_1014,N_646,N_563);
and U1015 (N_1015,N_878,N_757);
nor U1016 (N_1016,N_549,N_882);
nor U1017 (N_1017,N_663,N_597);
xnor U1018 (N_1018,N_853,N_753);
and U1019 (N_1019,N_650,N_966);
xnor U1020 (N_1020,N_583,N_715);
nor U1021 (N_1021,N_947,N_845);
nor U1022 (N_1022,N_574,N_770);
nor U1023 (N_1023,N_973,N_844);
nand U1024 (N_1024,N_739,N_986);
and U1025 (N_1025,N_554,N_755);
and U1026 (N_1026,N_516,N_590);
nor U1027 (N_1027,N_988,N_731);
xor U1028 (N_1028,N_936,N_562);
or U1029 (N_1029,N_568,N_933);
nor U1030 (N_1030,N_814,N_671);
and U1031 (N_1031,N_617,N_709);
nand U1032 (N_1032,N_927,N_692);
and U1033 (N_1033,N_541,N_948);
xnor U1034 (N_1034,N_884,N_807);
nand U1035 (N_1035,N_539,N_921);
or U1036 (N_1036,N_874,N_904);
or U1037 (N_1037,N_522,N_934);
or U1038 (N_1038,N_660,N_839);
or U1039 (N_1039,N_866,N_600);
and U1040 (N_1040,N_767,N_775);
xnor U1041 (N_1041,N_707,N_683);
xor U1042 (N_1042,N_889,N_726);
nand U1043 (N_1043,N_593,N_582);
nand U1044 (N_1044,N_993,N_959);
and U1045 (N_1045,N_728,N_990);
or U1046 (N_1046,N_512,N_931);
or U1047 (N_1047,N_840,N_538);
and U1048 (N_1048,N_756,N_781);
and U1049 (N_1049,N_524,N_902);
nand U1050 (N_1050,N_951,N_849);
nand U1051 (N_1051,N_942,N_752);
xor U1052 (N_1052,N_928,N_615);
or U1053 (N_1053,N_564,N_620);
or U1054 (N_1054,N_648,N_673);
or U1055 (N_1055,N_519,N_822);
nor U1056 (N_1056,N_975,N_510);
nand U1057 (N_1057,N_808,N_824);
xnor U1058 (N_1058,N_675,N_880);
nor U1059 (N_1059,N_837,N_635);
nand U1060 (N_1060,N_654,N_954);
nor U1061 (N_1061,N_801,N_651);
or U1062 (N_1062,N_890,N_528);
and U1063 (N_1063,N_613,N_879);
and U1064 (N_1064,N_883,N_508);
nand U1065 (N_1065,N_924,N_587);
nand U1066 (N_1066,N_970,N_609);
nand U1067 (N_1067,N_905,N_687);
xnor U1068 (N_1068,N_532,N_714);
or U1069 (N_1069,N_831,N_566);
and U1070 (N_1070,N_690,N_596);
or U1071 (N_1071,N_926,N_720);
nand U1072 (N_1072,N_636,N_804);
xnor U1073 (N_1073,N_779,N_847);
or U1074 (N_1074,N_751,N_718);
or U1075 (N_1075,N_830,N_693);
or U1076 (N_1076,N_547,N_502);
or U1077 (N_1077,N_594,N_531);
or U1078 (N_1078,N_588,N_944);
nand U1079 (N_1079,N_935,N_796);
and U1080 (N_1080,N_901,N_891);
nand U1081 (N_1081,N_833,N_865);
nor U1082 (N_1082,N_634,N_614);
or U1083 (N_1083,N_703,N_961);
nor U1084 (N_1084,N_545,N_567);
nand U1085 (N_1085,N_786,N_920);
nand U1086 (N_1086,N_592,N_619);
or U1087 (N_1087,N_559,N_772);
or U1088 (N_1088,N_644,N_643);
nor U1089 (N_1089,N_965,N_577);
nand U1090 (N_1090,N_806,N_979);
nor U1091 (N_1091,N_639,N_676);
and U1092 (N_1092,N_730,N_842);
or U1093 (N_1093,N_680,N_907);
nand U1094 (N_1094,N_584,N_700);
nor U1095 (N_1095,N_881,N_998);
or U1096 (N_1096,N_809,N_957);
or U1097 (N_1097,N_789,N_744);
and U1098 (N_1098,N_886,N_710);
or U1099 (N_1099,N_871,N_638);
or U1100 (N_1100,N_774,N_761);
and U1101 (N_1101,N_740,N_828);
xor U1102 (N_1102,N_919,N_616);
or U1103 (N_1103,N_794,N_598);
or U1104 (N_1104,N_949,N_537);
or U1105 (N_1105,N_713,N_533);
xor U1106 (N_1106,N_685,N_606);
xnor U1107 (N_1107,N_869,N_610);
or U1108 (N_1108,N_511,N_820);
nor U1109 (N_1109,N_963,N_657);
or U1110 (N_1110,N_500,N_585);
nor U1111 (N_1111,N_678,N_893);
xnor U1112 (N_1112,N_586,N_503);
nand U1113 (N_1113,N_642,N_631);
xor U1114 (N_1114,N_704,N_906);
nand U1115 (N_1115,N_708,N_754);
xor U1116 (N_1116,N_798,N_721);
nand U1117 (N_1117,N_723,N_725);
nor U1118 (N_1118,N_958,N_735);
xor U1119 (N_1119,N_867,N_797);
nand U1120 (N_1120,N_552,N_581);
or U1121 (N_1121,N_625,N_938);
xnor U1122 (N_1122,N_764,N_826);
nor U1123 (N_1123,N_923,N_981);
xnor U1124 (N_1124,N_705,N_911);
xor U1125 (N_1125,N_940,N_939);
xor U1126 (N_1126,N_895,N_759);
or U1127 (N_1127,N_737,N_802);
or U1128 (N_1128,N_733,N_624);
nor U1129 (N_1129,N_558,N_819);
or U1130 (N_1130,N_969,N_914);
xnor U1131 (N_1131,N_748,N_556);
and U1132 (N_1132,N_507,N_857);
or U1133 (N_1133,N_551,N_862);
nor U1134 (N_1134,N_745,N_898);
nand U1135 (N_1135,N_670,N_557);
and U1136 (N_1136,N_722,N_570);
nand U1137 (N_1137,N_605,N_523);
xor U1138 (N_1138,N_813,N_976);
nand U1139 (N_1139,N_829,N_529);
or U1140 (N_1140,N_945,N_621);
or U1141 (N_1141,N_688,N_892);
xor U1142 (N_1142,N_572,N_719);
nand U1143 (N_1143,N_623,N_825);
nand U1144 (N_1144,N_603,N_627);
nor U1145 (N_1145,N_553,N_929);
nand U1146 (N_1146,N_749,N_543);
xor U1147 (N_1147,N_738,N_604);
xor U1148 (N_1148,N_548,N_659);
or U1149 (N_1149,N_504,N_991);
xor U1150 (N_1150,N_972,N_542);
nand U1151 (N_1151,N_578,N_922);
and U1152 (N_1152,N_870,N_812);
nand U1153 (N_1153,N_937,N_915);
or U1154 (N_1154,N_854,N_527);
or U1155 (N_1155,N_746,N_985);
nand U1156 (N_1156,N_956,N_974);
and U1157 (N_1157,N_815,N_697);
and U1158 (N_1158,N_787,N_967);
or U1159 (N_1159,N_652,N_711);
nor U1160 (N_1160,N_505,N_987);
or U1161 (N_1161,N_864,N_701);
nand U1162 (N_1162,N_736,N_821);
or U1163 (N_1163,N_618,N_964);
and U1164 (N_1164,N_912,N_877);
nor U1165 (N_1165,N_827,N_784);
and U1166 (N_1166,N_832,N_875);
nand U1167 (N_1167,N_803,N_950);
xnor U1168 (N_1168,N_978,N_580);
nand U1169 (N_1169,N_897,N_766);
or U1170 (N_1170,N_916,N_816);
xor U1171 (N_1171,N_571,N_655);
or U1172 (N_1172,N_521,N_530);
nand U1173 (N_1173,N_702,N_540);
or U1174 (N_1174,N_595,N_888);
or U1175 (N_1175,N_918,N_626);
xnor U1176 (N_1176,N_599,N_971);
nand U1177 (N_1177,N_835,N_661);
or U1178 (N_1178,N_903,N_691);
and U1179 (N_1179,N_795,N_834);
nand U1180 (N_1180,N_649,N_666);
or U1181 (N_1181,N_729,N_656);
xor U1182 (N_1182,N_763,N_658);
and U1183 (N_1183,N_995,N_777);
nand U1184 (N_1184,N_743,N_546);
xnor U1185 (N_1185,N_518,N_667);
and U1186 (N_1186,N_999,N_535);
xnor U1187 (N_1187,N_716,N_607);
and U1188 (N_1188,N_765,N_896);
and U1189 (N_1189,N_885,N_984);
and U1190 (N_1190,N_941,N_672);
or U1191 (N_1191,N_750,N_873);
nand U1192 (N_1192,N_953,N_677);
nor U1193 (N_1193,N_555,N_622);
or U1194 (N_1194,N_810,N_805);
xor U1195 (N_1195,N_525,N_561);
nand U1196 (N_1196,N_946,N_741);
and U1197 (N_1197,N_856,N_669);
and U1198 (N_1198,N_501,N_811);
xnor U1199 (N_1199,N_836,N_506);
and U1200 (N_1200,N_611,N_608);
or U1201 (N_1201,N_647,N_968);
nor U1202 (N_1202,N_633,N_681);
xnor U1203 (N_1203,N_855,N_717);
nand U1204 (N_1204,N_569,N_989);
xor U1205 (N_1205,N_742,N_860);
nor U1206 (N_1206,N_637,N_818);
and U1207 (N_1207,N_997,N_630);
nor U1208 (N_1208,N_910,N_579);
or U1209 (N_1209,N_917,N_843);
nor U1210 (N_1210,N_930,N_788);
and U1211 (N_1211,N_664,N_712);
nor U1212 (N_1212,N_526,N_778);
and U1213 (N_1213,N_632,N_800);
nor U1214 (N_1214,N_565,N_544);
nand U1215 (N_1215,N_696,N_852);
and U1216 (N_1216,N_679,N_550);
and U1217 (N_1217,N_846,N_977);
and U1218 (N_1218,N_876,N_674);
nor U1219 (N_1219,N_925,N_520);
or U1220 (N_1220,N_793,N_602);
and U1221 (N_1221,N_665,N_980);
nor U1222 (N_1222,N_994,N_724);
xor U1223 (N_1223,N_762,N_573);
and U1224 (N_1224,N_645,N_960);
nand U1225 (N_1225,N_612,N_782);
or U1226 (N_1226,N_560,N_841);
or U1227 (N_1227,N_792,N_848);
nand U1228 (N_1228,N_859,N_694);
xnor U1229 (N_1229,N_536,N_838);
nor U1230 (N_1230,N_684,N_509);
and U1231 (N_1231,N_900,N_514);
nor U1232 (N_1232,N_734,N_698);
nand U1233 (N_1233,N_589,N_601);
xnor U1234 (N_1234,N_771,N_686);
or U1235 (N_1235,N_962,N_850);
nand U1236 (N_1236,N_943,N_783);
and U1237 (N_1237,N_517,N_732);
xor U1238 (N_1238,N_760,N_861);
nand U1239 (N_1239,N_668,N_858);
nor U1240 (N_1240,N_768,N_894);
and U1241 (N_1241,N_863,N_706);
or U1242 (N_1242,N_575,N_817);
nor U1243 (N_1243,N_640,N_513);
or U1244 (N_1244,N_773,N_628);
nand U1245 (N_1245,N_780,N_932);
xor U1246 (N_1246,N_908,N_982);
or U1247 (N_1247,N_591,N_769);
or U1248 (N_1248,N_695,N_887);
xnor U1249 (N_1249,N_629,N_534);
and U1250 (N_1250,N_857,N_923);
or U1251 (N_1251,N_715,N_856);
and U1252 (N_1252,N_845,N_607);
xnor U1253 (N_1253,N_674,N_695);
nand U1254 (N_1254,N_646,N_583);
or U1255 (N_1255,N_744,N_547);
and U1256 (N_1256,N_539,N_725);
nor U1257 (N_1257,N_899,N_707);
and U1258 (N_1258,N_737,N_770);
nor U1259 (N_1259,N_702,N_850);
and U1260 (N_1260,N_895,N_877);
nand U1261 (N_1261,N_658,N_727);
nand U1262 (N_1262,N_640,N_699);
and U1263 (N_1263,N_633,N_838);
and U1264 (N_1264,N_542,N_952);
nand U1265 (N_1265,N_632,N_945);
nor U1266 (N_1266,N_876,N_694);
and U1267 (N_1267,N_899,N_948);
nor U1268 (N_1268,N_522,N_996);
nor U1269 (N_1269,N_666,N_870);
nor U1270 (N_1270,N_901,N_798);
xor U1271 (N_1271,N_584,N_777);
nand U1272 (N_1272,N_557,N_816);
xnor U1273 (N_1273,N_640,N_778);
xnor U1274 (N_1274,N_940,N_620);
nand U1275 (N_1275,N_754,N_702);
nand U1276 (N_1276,N_682,N_894);
and U1277 (N_1277,N_618,N_603);
nand U1278 (N_1278,N_508,N_711);
nand U1279 (N_1279,N_680,N_575);
and U1280 (N_1280,N_613,N_527);
xnor U1281 (N_1281,N_677,N_729);
or U1282 (N_1282,N_573,N_564);
and U1283 (N_1283,N_617,N_874);
nand U1284 (N_1284,N_854,N_765);
xor U1285 (N_1285,N_912,N_758);
nand U1286 (N_1286,N_601,N_545);
and U1287 (N_1287,N_636,N_893);
xor U1288 (N_1288,N_521,N_799);
nor U1289 (N_1289,N_642,N_527);
nand U1290 (N_1290,N_977,N_614);
nor U1291 (N_1291,N_827,N_781);
nor U1292 (N_1292,N_634,N_635);
and U1293 (N_1293,N_871,N_790);
nor U1294 (N_1294,N_635,N_642);
and U1295 (N_1295,N_783,N_987);
xor U1296 (N_1296,N_693,N_972);
nand U1297 (N_1297,N_621,N_640);
nand U1298 (N_1298,N_987,N_578);
xnor U1299 (N_1299,N_873,N_981);
or U1300 (N_1300,N_905,N_950);
or U1301 (N_1301,N_505,N_609);
xnor U1302 (N_1302,N_808,N_667);
nor U1303 (N_1303,N_921,N_582);
and U1304 (N_1304,N_857,N_789);
xor U1305 (N_1305,N_657,N_634);
xor U1306 (N_1306,N_573,N_994);
and U1307 (N_1307,N_762,N_555);
or U1308 (N_1308,N_637,N_963);
nor U1309 (N_1309,N_643,N_920);
and U1310 (N_1310,N_993,N_886);
nand U1311 (N_1311,N_838,N_620);
nor U1312 (N_1312,N_944,N_930);
and U1313 (N_1313,N_940,N_805);
nand U1314 (N_1314,N_911,N_676);
or U1315 (N_1315,N_968,N_937);
nand U1316 (N_1316,N_659,N_741);
xor U1317 (N_1317,N_600,N_669);
xnor U1318 (N_1318,N_688,N_605);
and U1319 (N_1319,N_938,N_775);
or U1320 (N_1320,N_581,N_621);
xor U1321 (N_1321,N_937,N_946);
or U1322 (N_1322,N_872,N_781);
nand U1323 (N_1323,N_613,N_530);
and U1324 (N_1324,N_509,N_864);
nor U1325 (N_1325,N_541,N_831);
nand U1326 (N_1326,N_727,N_611);
xnor U1327 (N_1327,N_914,N_786);
or U1328 (N_1328,N_751,N_607);
nand U1329 (N_1329,N_568,N_601);
nor U1330 (N_1330,N_604,N_906);
nor U1331 (N_1331,N_570,N_756);
and U1332 (N_1332,N_527,N_961);
nand U1333 (N_1333,N_789,N_796);
nand U1334 (N_1334,N_945,N_593);
or U1335 (N_1335,N_822,N_940);
nor U1336 (N_1336,N_775,N_530);
nand U1337 (N_1337,N_720,N_997);
xnor U1338 (N_1338,N_969,N_844);
xor U1339 (N_1339,N_796,N_779);
xnor U1340 (N_1340,N_683,N_983);
xnor U1341 (N_1341,N_916,N_658);
or U1342 (N_1342,N_594,N_574);
xor U1343 (N_1343,N_784,N_988);
nor U1344 (N_1344,N_898,N_805);
or U1345 (N_1345,N_652,N_803);
or U1346 (N_1346,N_544,N_921);
and U1347 (N_1347,N_638,N_884);
and U1348 (N_1348,N_914,N_541);
or U1349 (N_1349,N_751,N_733);
nor U1350 (N_1350,N_511,N_697);
xor U1351 (N_1351,N_778,N_906);
nor U1352 (N_1352,N_684,N_834);
or U1353 (N_1353,N_957,N_736);
and U1354 (N_1354,N_835,N_868);
xnor U1355 (N_1355,N_695,N_537);
nand U1356 (N_1356,N_640,N_620);
nor U1357 (N_1357,N_642,N_717);
xor U1358 (N_1358,N_933,N_682);
or U1359 (N_1359,N_734,N_724);
xor U1360 (N_1360,N_851,N_663);
or U1361 (N_1361,N_714,N_900);
nand U1362 (N_1362,N_889,N_839);
nor U1363 (N_1363,N_630,N_798);
nor U1364 (N_1364,N_612,N_836);
xnor U1365 (N_1365,N_809,N_586);
and U1366 (N_1366,N_869,N_588);
nor U1367 (N_1367,N_906,N_616);
or U1368 (N_1368,N_930,N_650);
and U1369 (N_1369,N_728,N_754);
xor U1370 (N_1370,N_796,N_877);
xnor U1371 (N_1371,N_938,N_662);
or U1372 (N_1372,N_780,N_622);
nor U1373 (N_1373,N_652,N_540);
nor U1374 (N_1374,N_964,N_814);
and U1375 (N_1375,N_922,N_772);
and U1376 (N_1376,N_565,N_504);
nor U1377 (N_1377,N_589,N_795);
nor U1378 (N_1378,N_691,N_519);
nor U1379 (N_1379,N_700,N_790);
nand U1380 (N_1380,N_503,N_703);
xnor U1381 (N_1381,N_771,N_960);
nand U1382 (N_1382,N_821,N_623);
or U1383 (N_1383,N_604,N_581);
nor U1384 (N_1384,N_539,N_963);
xor U1385 (N_1385,N_883,N_820);
nand U1386 (N_1386,N_694,N_599);
and U1387 (N_1387,N_565,N_863);
xnor U1388 (N_1388,N_825,N_992);
nor U1389 (N_1389,N_716,N_720);
or U1390 (N_1390,N_986,N_554);
xor U1391 (N_1391,N_590,N_909);
xnor U1392 (N_1392,N_920,N_728);
or U1393 (N_1393,N_563,N_824);
xnor U1394 (N_1394,N_941,N_803);
nor U1395 (N_1395,N_585,N_545);
and U1396 (N_1396,N_520,N_587);
nor U1397 (N_1397,N_677,N_705);
nand U1398 (N_1398,N_848,N_984);
or U1399 (N_1399,N_598,N_999);
or U1400 (N_1400,N_779,N_540);
xor U1401 (N_1401,N_804,N_776);
nand U1402 (N_1402,N_956,N_714);
xnor U1403 (N_1403,N_680,N_655);
xnor U1404 (N_1404,N_846,N_611);
or U1405 (N_1405,N_966,N_571);
xnor U1406 (N_1406,N_765,N_773);
nor U1407 (N_1407,N_854,N_509);
nor U1408 (N_1408,N_592,N_909);
nor U1409 (N_1409,N_508,N_836);
and U1410 (N_1410,N_948,N_965);
and U1411 (N_1411,N_887,N_606);
xor U1412 (N_1412,N_943,N_849);
and U1413 (N_1413,N_794,N_835);
and U1414 (N_1414,N_622,N_626);
nand U1415 (N_1415,N_594,N_695);
xor U1416 (N_1416,N_864,N_644);
xnor U1417 (N_1417,N_825,N_948);
nor U1418 (N_1418,N_895,N_818);
nor U1419 (N_1419,N_680,N_560);
nor U1420 (N_1420,N_608,N_973);
and U1421 (N_1421,N_821,N_680);
nand U1422 (N_1422,N_936,N_789);
and U1423 (N_1423,N_799,N_528);
xor U1424 (N_1424,N_674,N_500);
nand U1425 (N_1425,N_748,N_527);
nor U1426 (N_1426,N_973,N_525);
xnor U1427 (N_1427,N_893,N_823);
xor U1428 (N_1428,N_753,N_628);
xnor U1429 (N_1429,N_946,N_687);
xor U1430 (N_1430,N_913,N_680);
or U1431 (N_1431,N_925,N_604);
nor U1432 (N_1432,N_692,N_552);
or U1433 (N_1433,N_989,N_865);
and U1434 (N_1434,N_880,N_849);
and U1435 (N_1435,N_631,N_915);
xor U1436 (N_1436,N_680,N_662);
nand U1437 (N_1437,N_736,N_609);
nand U1438 (N_1438,N_999,N_577);
and U1439 (N_1439,N_956,N_624);
and U1440 (N_1440,N_958,N_505);
and U1441 (N_1441,N_859,N_741);
nor U1442 (N_1442,N_777,N_677);
nand U1443 (N_1443,N_558,N_582);
nor U1444 (N_1444,N_588,N_699);
nor U1445 (N_1445,N_912,N_871);
nor U1446 (N_1446,N_605,N_942);
nor U1447 (N_1447,N_801,N_664);
or U1448 (N_1448,N_950,N_847);
nor U1449 (N_1449,N_770,N_907);
xor U1450 (N_1450,N_574,N_867);
and U1451 (N_1451,N_699,N_644);
and U1452 (N_1452,N_857,N_834);
or U1453 (N_1453,N_780,N_640);
xor U1454 (N_1454,N_548,N_590);
nor U1455 (N_1455,N_871,N_727);
xor U1456 (N_1456,N_614,N_566);
nand U1457 (N_1457,N_865,N_628);
nor U1458 (N_1458,N_715,N_828);
or U1459 (N_1459,N_644,N_913);
xnor U1460 (N_1460,N_825,N_973);
or U1461 (N_1461,N_513,N_608);
and U1462 (N_1462,N_629,N_701);
or U1463 (N_1463,N_972,N_597);
nand U1464 (N_1464,N_627,N_664);
or U1465 (N_1465,N_776,N_785);
xor U1466 (N_1466,N_587,N_832);
and U1467 (N_1467,N_772,N_564);
xor U1468 (N_1468,N_636,N_591);
nor U1469 (N_1469,N_774,N_684);
xor U1470 (N_1470,N_782,N_726);
or U1471 (N_1471,N_866,N_929);
and U1472 (N_1472,N_789,N_934);
and U1473 (N_1473,N_744,N_705);
nand U1474 (N_1474,N_960,N_775);
nand U1475 (N_1475,N_600,N_900);
xnor U1476 (N_1476,N_902,N_985);
and U1477 (N_1477,N_778,N_531);
nand U1478 (N_1478,N_805,N_913);
or U1479 (N_1479,N_739,N_551);
xor U1480 (N_1480,N_939,N_835);
nor U1481 (N_1481,N_643,N_680);
nor U1482 (N_1482,N_747,N_852);
xnor U1483 (N_1483,N_528,N_538);
and U1484 (N_1484,N_926,N_999);
or U1485 (N_1485,N_558,N_533);
or U1486 (N_1486,N_812,N_959);
xor U1487 (N_1487,N_732,N_725);
nand U1488 (N_1488,N_807,N_651);
nor U1489 (N_1489,N_500,N_995);
xor U1490 (N_1490,N_773,N_724);
or U1491 (N_1491,N_621,N_635);
xor U1492 (N_1492,N_506,N_863);
or U1493 (N_1493,N_928,N_526);
nor U1494 (N_1494,N_730,N_645);
nor U1495 (N_1495,N_530,N_500);
or U1496 (N_1496,N_569,N_667);
nor U1497 (N_1497,N_585,N_818);
xnor U1498 (N_1498,N_556,N_836);
or U1499 (N_1499,N_817,N_954);
xnor U1500 (N_1500,N_1355,N_1122);
nor U1501 (N_1501,N_1104,N_1013);
nor U1502 (N_1502,N_1123,N_1117);
nand U1503 (N_1503,N_1134,N_1114);
and U1504 (N_1504,N_1020,N_1177);
xor U1505 (N_1505,N_1178,N_1248);
or U1506 (N_1506,N_1046,N_1499);
or U1507 (N_1507,N_1314,N_1026);
and U1508 (N_1508,N_1307,N_1469);
or U1509 (N_1509,N_1411,N_1197);
and U1510 (N_1510,N_1113,N_1128);
or U1511 (N_1511,N_1472,N_1310);
and U1512 (N_1512,N_1403,N_1031);
or U1513 (N_1513,N_1230,N_1231);
or U1514 (N_1514,N_1004,N_1022);
nand U1515 (N_1515,N_1101,N_1321);
and U1516 (N_1516,N_1485,N_1090);
nand U1517 (N_1517,N_1143,N_1312);
or U1518 (N_1518,N_1270,N_1408);
and U1519 (N_1519,N_1381,N_1445);
or U1520 (N_1520,N_1169,N_1131);
or U1521 (N_1521,N_1171,N_1133);
nand U1522 (N_1522,N_1191,N_1125);
and U1523 (N_1523,N_1423,N_1359);
or U1524 (N_1524,N_1144,N_1220);
and U1525 (N_1525,N_1348,N_1461);
and U1526 (N_1526,N_1433,N_1049);
nor U1527 (N_1527,N_1202,N_1268);
and U1528 (N_1528,N_1300,N_1458);
nor U1529 (N_1529,N_1465,N_1391);
and U1530 (N_1530,N_1079,N_1162);
nor U1531 (N_1531,N_1100,N_1301);
nand U1532 (N_1532,N_1373,N_1141);
or U1533 (N_1533,N_1152,N_1137);
and U1534 (N_1534,N_1368,N_1416);
xnor U1535 (N_1535,N_1328,N_1192);
xnor U1536 (N_1536,N_1102,N_1120);
or U1537 (N_1537,N_1014,N_1116);
or U1538 (N_1538,N_1454,N_1198);
or U1539 (N_1539,N_1062,N_1462);
and U1540 (N_1540,N_1306,N_1057);
and U1541 (N_1541,N_1167,N_1394);
and U1542 (N_1542,N_1303,N_1362);
nand U1543 (N_1543,N_1324,N_1074);
and U1544 (N_1544,N_1332,N_1228);
and U1545 (N_1545,N_1369,N_1160);
or U1546 (N_1546,N_1339,N_1241);
xor U1547 (N_1547,N_1080,N_1235);
xor U1548 (N_1548,N_1098,N_1239);
or U1549 (N_1549,N_1407,N_1092);
and U1550 (N_1550,N_1190,N_1233);
nor U1551 (N_1551,N_1290,N_1262);
nor U1552 (N_1552,N_1259,N_1015);
xor U1553 (N_1553,N_1376,N_1099);
nand U1554 (N_1554,N_1088,N_1367);
nand U1555 (N_1555,N_1110,N_1495);
or U1556 (N_1556,N_1449,N_1371);
or U1557 (N_1557,N_1294,N_1149);
nor U1558 (N_1558,N_1135,N_1164);
and U1559 (N_1559,N_1345,N_1442);
xor U1560 (N_1560,N_1217,N_1209);
or U1561 (N_1561,N_1253,N_1444);
xnor U1562 (N_1562,N_1374,N_1398);
nor U1563 (N_1563,N_1382,N_1288);
and U1564 (N_1564,N_1023,N_1224);
or U1565 (N_1565,N_1330,N_1068);
nand U1566 (N_1566,N_1446,N_1419);
and U1567 (N_1567,N_1103,N_1346);
and U1568 (N_1568,N_1042,N_1184);
nor U1569 (N_1569,N_1308,N_1161);
xnor U1570 (N_1570,N_1280,N_1482);
nand U1571 (N_1571,N_1352,N_1410);
nand U1572 (N_1572,N_1199,N_1414);
and U1573 (N_1573,N_1127,N_1347);
and U1574 (N_1574,N_1287,N_1093);
or U1575 (N_1575,N_1138,N_1201);
nor U1576 (N_1576,N_1395,N_1058);
or U1577 (N_1577,N_1354,N_1071);
nor U1578 (N_1578,N_1147,N_1072);
nor U1579 (N_1579,N_1305,N_1335);
or U1580 (N_1580,N_1492,N_1342);
nand U1581 (N_1581,N_1226,N_1258);
nor U1582 (N_1582,N_1256,N_1351);
xor U1583 (N_1583,N_1174,N_1084);
nand U1584 (N_1584,N_1487,N_1337);
nor U1585 (N_1585,N_1195,N_1457);
nand U1586 (N_1586,N_1311,N_1349);
and U1587 (N_1587,N_1431,N_1210);
nor U1588 (N_1588,N_1263,N_1309);
xor U1589 (N_1589,N_1393,N_1139);
and U1590 (N_1590,N_1343,N_1254);
or U1591 (N_1591,N_1331,N_1471);
xor U1592 (N_1592,N_1405,N_1075);
and U1593 (N_1593,N_1420,N_1064);
and U1594 (N_1594,N_1432,N_1397);
or U1595 (N_1595,N_1142,N_1063);
and U1596 (N_1596,N_1183,N_1082);
nand U1597 (N_1597,N_1059,N_1281);
and U1598 (N_1598,N_1245,N_1404);
nand U1599 (N_1599,N_1479,N_1238);
and U1600 (N_1600,N_1484,N_1317);
and U1601 (N_1601,N_1086,N_1412);
nand U1602 (N_1602,N_1402,N_1054);
nand U1603 (N_1603,N_1112,N_1474);
or U1604 (N_1604,N_1051,N_1315);
nand U1605 (N_1605,N_1165,N_1400);
xnor U1606 (N_1606,N_1021,N_1399);
and U1607 (N_1607,N_1157,N_1111);
and U1608 (N_1608,N_1477,N_1409);
and U1609 (N_1609,N_1194,N_1237);
or U1610 (N_1610,N_1247,N_1480);
nor U1611 (N_1611,N_1200,N_1163);
nand U1612 (N_1612,N_1413,N_1003);
and U1613 (N_1613,N_1221,N_1406);
and U1614 (N_1614,N_1272,N_1207);
nand U1615 (N_1615,N_1363,N_1214);
or U1616 (N_1616,N_1069,N_1212);
nand U1617 (N_1617,N_1279,N_1087);
and U1618 (N_1618,N_1481,N_1322);
and U1619 (N_1619,N_1118,N_1229);
nor U1620 (N_1620,N_1091,N_1129);
xnor U1621 (N_1621,N_1286,N_1034);
nor U1622 (N_1622,N_1425,N_1105);
and U1623 (N_1623,N_1298,N_1089);
nand U1624 (N_1624,N_1044,N_1204);
or U1625 (N_1625,N_1260,N_1379);
nor U1626 (N_1626,N_1437,N_1292);
nand U1627 (N_1627,N_1269,N_1353);
nand U1628 (N_1628,N_1033,N_1327);
nor U1629 (N_1629,N_1271,N_1356);
and U1630 (N_1630,N_1140,N_1490);
xor U1631 (N_1631,N_1418,N_1340);
or U1632 (N_1632,N_1032,N_1187);
xnor U1633 (N_1633,N_1040,N_1218);
and U1634 (N_1634,N_1106,N_1296);
nand U1635 (N_1635,N_1056,N_1430);
nor U1636 (N_1636,N_1483,N_1284);
nor U1637 (N_1637,N_1266,N_1037);
nand U1638 (N_1638,N_1424,N_1278);
and U1639 (N_1639,N_1028,N_1486);
nand U1640 (N_1640,N_1428,N_1264);
xor U1641 (N_1641,N_1323,N_1146);
nor U1642 (N_1642,N_1196,N_1460);
or U1643 (N_1643,N_1030,N_1320);
xor U1644 (N_1644,N_1243,N_1316);
or U1645 (N_1645,N_1273,N_1094);
or U1646 (N_1646,N_1350,N_1211);
xnor U1647 (N_1647,N_1473,N_1488);
nand U1648 (N_1648,N_1427,N_1456);
or U1649 (N_1649,N_1277,N_1150);
or U1650 (N_1650,N_1297,N_1438);
nor U1651 (N_1651,N_1396,N_1024);
nand U1652 (N_1652,N_1010,N_1050);
nand U1653 (N_1653,N_1401,N_1159);
xor U1654 (N_1654,N_1372,N_1038);
and U1655 (N_1655,N_1006,N_1045);
xor U1656 (N_1656,N_1452,N_1180);
nand U1657 (N_1657,N_1291,N_1225);
nand U1658 (N_1658,N_1203,N_1078);
nor U1659 (N_1659,N_1083,N_1333);
or U1660 (N_1660,N_1453,N_1007);
nor U1661 (N_1661,N_1166,N_1012);
nand U1662 (N_1662,N_1389,N_1336);
nor U1663 (N_1663,N_1383,N_1421);
or U1664 (N_1664,N_1464,N_1377);
or U1665 (N_1665,N_1170,N_1041);
xor U1666 (N_1666,N_1326,N_1455);
nor U1667 (N_1667,N_1478,N_1148);
or U1668 (N_1668,N_1334,N_1039);
nor U1669 (N_1669,N_1188,N_1017);
xor U1670 (N_1670,N_1009,N_1047);
nor U1671 (N_1671,N_1358,N_1151);
nand U1672 (N_1672,N_1341,N_1344);
nand U1673 (N_1673,N_1095,N_1491);
xor U1674 (N_1674,N_1215,N_1249);
xor U1675 (N_1675,N_1441,N_1386);
or U1676 (N_1676,N_1126,N_1498);
or U1677 (N_1677,N_1206,N_1276);
or U1678 (N_1678,N_1066,N_1476);
xor U1679 (N_1679,N_1076,N_1463);
and U1680 (N_1680,N_1029,N_1459);
nor U1681 (N_1681,N_1246,N_1440);
nand U1682 (N_1682,N_1222,N_1065);
and U1683 (N_1683,N_1053,N_1475);
xor U1684 (N_1684,N_1018,N_1319);
or U1685 (N_1685,N_1275,N_1274);
nor U1686 (N_1686,N_1067,N_1357);
or U1687 (N_1687,N_1005,N_1216);
nand U1688 (N_1688,N_1257,N_1283);
and U1689 (N_1689,N_1497,N_1002);
and U1690 (N_1690,N_1434,N_1107);
xor U1691 (N_1691,N_1435,N_1097);
xor U1692 (N_1692,N_1213,N_1136);
and U1693 (N_1693,N_1267,N_1392);
and U1694 (N_1694,N_1360,N_1450);
nor U1695 (N_1695,N_1158,N_1130);
nor U1696 (N_1696,N_1390,N_1329);
or U1697 (N_1697,N_1132,N_1155);
xor U1698 (N_1698,N_1467,N_1109);
and U1699 (N_1699,N_1077,N_1115);
xor U1700 (N_1700,N_1001,N_1365);
nand U1701 (N_1701,N_1185,N_1154);
xor U1702 (N_1702,N_1375,N_1289);
nand U1703 (N_1703,N_1186,N_1055);
nor U1704 (N_1704,N_1299,N_1035);
or U1705 (N_1705,N_1470,N_1124);
nand U1706 (N_1706,N_1008,N_1081);
or U1707 (N_1707,N_1227,N_1388);
xor U1708 (N_1708,N_1179,N_1338);
xnor U1709 (N_1709,N_1366,N_1240);
xor U1710 (N_1710,N_1378,N_1466);
nand U1711 (N_1711,N_1043,N_1182);
nor U1712 (N_1712,N_1380,N_1153);
nor U1713 (N_1713,N_1108,N_1489);
xnor U1714 (N_1714,N_1293,N_1181);
or U1715 (N_1715,N_1244,N_1302);
and U1716 (N_1716,N_1384,N_1493);
nor U1717 (N_1717,N_1000,N_1168);
or U1718 (N_1718,N_1261,N_1027);
nor U1719 (N_1719,N_1193,N_1208);
or U1720 (N_1720,N_1325,N_1304);
nand U1721 (N_1721,N_1385,N_1025);
or U1722 (N_1722,N_1119,N_1250);
or U1723 (N_1723,N_1447,N_1219);
xnor U1724 (N_1724,N_1295,N_1036);
and U1725 (N_1725,N_1451,N_1156);
or U1726 (N_1726,N_1448,N_1172);
nand U1727 (N_1727,N_1234,N_1016);
xor U1728 (N_1728,N_1236,N_1052);
nand U1729 (N_1729,N_1189,N_1426);
nor U1730 (N_1730,N_1242,N_1422);
and U1731 (N_1731,N_1255,N_1443);
nor U1732 (N_1732,N_1173,N_1494);
nor U1733 (N_1733,N_1313,N_1468);
and U1734 (N_1734,N_1251,N_1232);
and U1735 (N_1735,N_1085,N_1387);
xnor U1736 (N_1736,N_1048,N_1252);
or U1737 (N_1737,N_1096,N_1361);
or U1738 (N_1738,N_1223,N_1176);
or U1739 (N_1739,N_1282,N_1205);
nor U1740 (N_1740,N_1364,N_1265);
xnor U1741 (N_1741,N_1011,N_1285);
xor U1742 (N_1742,N_1370,N_1439);
nand U1743 (N_1743,N_1436,N_1429);
or U1744 (N_1744,N_1175,N_1070);
nand U1745 (N_1745,N_1417,N_1145);
nand U1746 (N_1746,N_1073,N_1061);
nand U1747 (N_1747,N_1415,N_1060);
or U1748 (N_1748,N_1318,N_1019);
xnor U1749 (N_1749,N_1496,N_1121);
or U1750 (N_1750,N_1108,N_1462);
xnor U1751 (N_1751,N_1163,N_1133);
nand U1752 (N_1752,N_1087,N_1320);
and U1753 (N_1753,N_1081,N_1171);
xnor U1754 (N_1754,N_1139,N_1259);
nand U1755 (N_1755,N_1224,N_1016);
or U1756 (N_1756,N_1059,N_1048);
xor U1757 (N_1757,N_1088,N_1317);
and U1758 (N_1758,N_1189,N_1455);
nor U1759 (N_1759,N_1005,N_1349);
nand U1760 (N_1760,N_1292,N_1391);
nor U1761 (N_1761,N_1489,N_1141);
xor U1762 (N_1762,N_1056,N_1180);
nand U1763 (N_1763,N_1377,N_1010);
nor U1764 (N_1764,N_1431,N_1070);
nand U1765 (N_1765,N_1476,N_1104);
nor U1766 (N_1766,N_1429,N_1485);
nor U1767 (N_1767,N_1495,N_1134);
or U1768 (N_1768,N_1306,N_1163);
nand U1769 (N_1769,N_1203,N_1100);
nand U1770 (N_1770,N_1264,N_1028);
xnor U1771 (N_1771,N_1432,N_1357);
nor U1772 (N_1772,N_1334,N_1445);
xor U1773 (N_1773,N_1091,N_1304);
nand U1774 (N_1774,N_1224,N_1279);
nor U1775 (N_1775,N_1243,N_1228);
and U1776 (N_1776,N_1165,N_1255);
or U1777 (N_1777,N_1400,N_1451);
xor U1778 (N_1778,N_1479,N_1241);
xor U1779 (N_1779,N_1471,N_1025);
nor U1780 (N_1780,N_1256,N_1437);
nand U1781 (N_1781,N_1416,N_1354);
xnor U1782 (N_1782,N_1299,N_1294);
nand U1783 (N_1783,N_1473,N_1187);
xnor U1784 (N_1784,N_1451,N_1142);
and U1785 (N_1785,N_1373,N_1057);
nor U1786 (N_1786,N_1328,N_1199);
and U1787 (N_1787,N_1391,N_1097);
nor U1788 (N_1788,N_1053,N_1287);
and U1789 (N_1789,N_1351,N_1172);
nor U1790 (N_1790,N_1091,N_1319);
or U1791 (N_1791,N_1472,N_1196);
xnor U1792 (N_1792,N_1499,N_1228);
nor U1793 (N_1793,N_1244,N_1493);
nor U1794 (N_1794,N_1214,N_1316);
xor U1795 (N_1795,N_1400,N_1111);
nor U1796 (N_1796,N_1236,N_1301);
and U1797 (N_1797,N_1276,N_1416);
and U1798 (N_1798,N_1056,N_1117);
nand U1799 (N_1799,N_1316,N_1231);
and U1800 (N_1800,N_1192,N_1039);
nand U1801 (N_1801,N_1386,N_1323);
nor U1802 (N_1802,N_1299,N_1103);
nor U1803 (N_1803,N_1227,N_1107);
xnor U1804 (N_1804,N_1484,N_1496);
or U1805 (N_1805,N_1247,N_1402);
xnor U1806 (N_1806,N_1078,N_1394);
nor U1807 (N_1807,N_1367,N_1427);
or U1808 (N_1808,N_1068,N_1413);
nand U1809 (N_1809,N_1098,N_1000);
or U1810 (N_1810,N_1076,N_1108);
nand U1811 (N_1811,N_1258,N_1056);
nor U1812 (N_1812,N_1121,N_1082);
nand U1813 (N_1813,N_1381,N_1452);
or U1814 (N_1814,N_1424,N_1233);
nor U1815 (N_1815,N_1111,N_1418);
nor U1816 (N_1816,N_1291,N_1401);
and U1817 (N_1817,N_1211,N_1466);
nor U1818 (N_1818,N_1491,N_1221);
nand U1819 (N_1819,N_1194,N_1138);
nor U1820 (N_1820,N_1373,N_1451);
xor U1821 (N_1821,N_1384,N_1150);
xor U1822 (N_1822,N_1323,N_1413);
nand U1823 (N_1823,N_1430,N_1027);
xor U1824 (N_1824,N_1234,N_1396);
or U1825 (N_1825,N_1347,N_1475);
or U1826 (N_1826,N_1011,N_1317);
and U1827 (N_1827,N_1323,N_1145);
xnor U1828 (N_1828,N_1041,N_1229);
nor U1829 (N_1829,N_1277,N_1372);
nor U1830 (N_1830,N_1281,N_1056);
or U1831 (N_1831,N_1199,N_1332);
nand U1832 (N_1832,N_1404,N_1355);
xor U1833 (N_1833,N_1252,N_1406);
and U1834 (N_1834,N_1487,N_1458);
and U1835 (N_1835,N_1414,N_1278);
nor U1836 (N_1836,N_1466,N_1289);
xnor U1837 (N_1837,N_1011,N_1124);
nor U1838 (N_1838,N_1211,N_1475);
nand U1839 (N_1839,N_1051,N_1232);
xnor U1840 (N_1840,N_1017,N_1312);
or U1841 (N_1841,N_1279,N_1339);
or U1842 (N_1842,N_1046,N_1429);
nand U1843 (N_1843,N_1261,N_1427);
nand U1844 (N_1844,N_1130,N_1105);
nand U1845 (N_1845,N_1003,N_1159);
nor U1846 (N_1846,N_1325,N_1192);
nand U1847 (N_1847,N_1116,N_1498);
nand U1848 (N_1848,N_1088,N_1328);
nand U1849 (N_1849,N_1001,N_1451);
or U1850 (N_1850,N_1159,N_1219);
or U1851 (N_1851,N_1390,N_1037);
xor U1852 (N_1852,N_1259,N_1375);
xnor U1853 (N_1853,N_1292,N_1011);
nand U1854 (N_1854,N_1153,N_1300);
nand U1855 (N_1855,N_1008,N_1139);
nor U1856 (N_1856,N_1490,N_1443);
or U1857 (N_1857,N_1001,N_1136);
nand U1858 (N_1858,N_1496,N_1124);
and U1859 (N_1859,N_1345,N_1148);
nand U1860 (N_1860,N_1294,N_1235);
or U1861 (N_1861,N_1004,N_1098);
nor U1862 (N_1862,N_1472,N_1049);
or U1863 (N_1863,N_1343,N_1172);
nand U1864 (N_1864,N_1163,N_1469);
and U1865 (N_1865,N_1091,N_1323);
xor U1866 (N_1866,N_1256,N_1056);
nor U1867 (N_1867,N_1135,N_1179);
and U1868 (N_1868,N_1349,N_1019);
and U1869 (N_1869,N_1129,N_1202);
nor U1870 (N_1870,N_1326,N_1361);
nand U1871 (N_1871,N_1375,N_1185);
xor U1872 (N_1872,N_1089,N_1224);
or U1873 (N_1873,N_1407,N_1153);
xor U1874 (N_1874,N_1410,N_1309);
xor U1875 (N_1875,N_1240,N_1373);
xnor U1876 (N_1876,N_1456,N_1412);
or U1877 (N_1877,N_1066,N_1252);
nor U1878 (N_1878,N_1325,N_1329);
xor U1879 (N_1879,N_1260,N_1276);
nor U1880 (N_1880,N_1170,N_1198);
nand U1881 (N_1881,N_1382,N_1006);
and U1882 (N_1882,N_1296,N_1202);
or U1883 (N_1883,N_1494,N_1277);
nand U1884 (N_1884,N_1452,N_1147);
xor U1885 (N_1885,N_1284,N_1216);
nor U1886 (N_1886,N_1266,N_1095);
or U1887 (N_1887,N_1306,N_1176);
and U1888 (N_1888,N_1193,N_1406);
xnor U1889 (N_1889,N_1418,N_1016);
or U1890 (N_1890,N_1354,N_1310);
or U1891 (N_1891,N_1019,N_1270);
nand U1892 (N_1892,N_1458,N_1041);
xnor U1893 (N_1893,N_1120,N_1476);
or U1894 (N_1894,N_1429,N_1360);
xor U1895 (N_1895,N_1325,N_1054);
and U1896 (N_1896,N_1435,N_1331);
and U1897 (N_1897,N_1447,N_1448);
xnor U1898 (N_1898,N_1413,N_1498);
nand U1899 (N_1899,N_1072,N_1429);
and U1900 (N_1900,N_1234,N_1189);
and U1901 (N_1901,N_1362,N_1144);
or U1902 (N_1902,N_1327,N_1059);
and U1903 (N_1903,N_1016,N_1451);
nand U1904 (N_1904,N_1394,N_1462);
and U1905 (N_1905,N_1122,N_1276);
and U1906 (N_1906,N_1040,N_1162);
xor U1907 (N_1907,N_1499,N_1035);
or U1908 (N_1908,N_1446,N_1425);
and U1909 (N_1909,N_1163,N_1498);
xor U1910 (N_1910,N_1127,N_1213);
xor U1911 (N_1911,N_1395,N_1324);
xor U1912 (N_1912,N_1282,N_1437);
xor U1913 (N_1913,N_1484,N_1230);
or U1914 (N_1914,N_1353,N_1059);
nor U1915 (N_1915,N_1275,N_1111);
xnor U1916 (N_1916,N_1283,N_1342);
nor U1917 (N_1917,N_1478,N_1018);
nand U1918 (N_1918,N_1055,N_1099);
or U1919 (N_1919,N_1174,N_1196);
xnor U1920 (N_1920,N_1381,N_1151);
xor U1921 (N_1921,N_1485,N_1282);
or U1922 (N_1922,N_1197,N_1187);
nor U1923 (N_1923,N_1379,N_1157);
nor U1924 (N_1924,N_1331,N_1179);
and U1925 (N_1925,N_1499,N_1446);
nor U1926 (N_1926,N_1229,N_1421);
nor U1927 (N_1927,N_1495,N_1316);
nor U1928 (N_1928,N_1155,N_1497);
or U1929 (N_1929,N_1352,N_1295);
nor U1930 (N_1930,N_1032,N_1241);
xnor U1931 (N_1931,N_1267,N_1349);
and U1932 (N_1932,N_1337,N_1268);
and U1933 (N_1933,N_1214,N_1074);
nor U1934 (N_1934,N_1211,N_1385);
xor U1935 (N_1935,N_1310,N_1346);
nand U1936 (N_1936,N_1101,N_1332);
and U1937 (N_1937,N_1219,N_1141);
xnor U1938 (N_1938,N_1028,N_1016);
or U1939 (N_1939,N_1366,N_1167);
nand U1940 (N_1940,N_1146,N_1221);
xor U1941 (N_1941,N_1012,N_1146);
nor U1942 (N_1942,N_1318,N_1471);
nand U1943 (N_1943,N_1221,N_1196);
xor U1944 (N_1944,N_1189,N_1383);
nor U1945 (N_1945,N_1036,N_1345);
xor U1946 (N_1946,N_1445,N_1472);
and U1947 (N_1947,N_1471,N_1121);
and U1948 (N_1948,N_1328,N_1062);
nor U1949 (N_1949,N_1146,N_1105);
nor U1950 (N_1950,N_1115,N_1446);
nor U1951 (N_1951,N_1353,N_1168);
and U1952 (N_1952,N_1105,N_1366);
or U1953 (N_1953,N_1133,N_1060);
xor U1954 (N_1954,N_1442,N_1395);
nor U1955 (N_1955,N_1343,N_1127);
nor U1956 (N_1956,N_1375,N_1346);
nor U1957 (N_1957,N_1025,N_1284);
xor U1958 (N_1958,N_1265,N_1213);
nand U1959 (N_1959,N_1144,N_1394);
nand U1960 (N_1960,N_1097,N_1083);
and U1961 (N_1961,N_1331,N_1119);
and U1962 (N_1962,N_1256,N_1010);
xnor U1963 (N_1963,N_1064,N_1117);
and U1964 (N_1964,N_1244,N_1292);
or U1965 (N_1965,N_1051,N_1034);
xnor U1966 (N_1966,N_1334,N_1394);
and U1967 (N_1967,N_1467,N_1205);
and U1968 (N_1968,N_1241,N_1005);
nand U1969 (N_1969,N_1283,N_1206);
or U1970 (N_1970,N_1119,N_1053);
xor U1971 (N_1971,N_1263,N_1005);
xnor U1972 (N_1972,N_1032,N_1139);
nor U1973 (N_1973,N_1032,N_1054);
nor U1974 (N_1974,N_1111,N_1255);
nor U1975 (N_1975,N_1276,N_1350);
nand U1976 (N_1976,N_1257,N_1175);
xnor U1977 (N_1977,N_1391,N_1018);
nor U1978 (N_1978,N_1448,N_1496);
or U1979 (N_1979,N_1056,N_1475);
or U1980 (N_1980,N_1052,N_1375);
or U1981 (N_1981,N_1333,N_1378);
nor U1982 (N_1982,N_1120,N_1317);
and U1983 (N_1983,N_1468,N_1017);
xor U1984 (N_1984,N_1196,N_1290);
and U1985 (N_1985,N_1494,N_1118);
nor U1986 (N_1986,N_1455,N_1098);
or U1987 (N_1987,N_1473,N_1109);
nor U1988 (N_1988,N_1159,N_1324);
xor U1989 (N_1989,N_1250,N_1363);
nand U1990 (N_1990,N_1311,N_1312);
and U1991 (N_1991,N_1164,N_1450);
nor U1992 (N_1992,N_1367,N_1468);
or U1993 (N_1993,N_1486,N_1313);
nor U1994 (N_1994,N_1237,N_1079);
nand U1995 (N_1995,N_1185,N_1491);
nor U1996 (N_1996,N_1408,N_1313);
nor U1997 (N_1997,N_1152,N_1328);
xnor U1998 (N_1998,N_1411,N_1366);
and U1999 (N_1999,N_1440,N_1331);
xor U2000 (N_2000,N_1680,N_1975);
nor U2001 (N_2001,N_1718,N_1646);
nor U2002 (N_2002,N_1681,N_1561);
and U2003 (N_2003,N_1583,N_1668);
nand U2004 (N_2004,N_1632,N_1542);
and U2005 (N_2005,N_1886,N_1928);
xor U2006 (N_2006,N_1837,N_1774);
xnor U2007 (N_2007,N_1764,N_1920);
or U2008 (N_2008,N_1981,N_1741);
and U2009 (N_2009,N_1734,N_1631);
xor U2010 (N_2010,N_1840,N_1563);
and U2011 (N_2011,N_1897,N_1969);
nand U2012 (N_2012,N_1825,N_1566);
or U2013 (N_2013,N_1937,N_1623);
nor U2014 (N_2014,N_1884,N_1751);
or U2015 (N_2015,N_1709,N_1992);
or U2016 (N_2016,N_1649,N_1761);
nand U2017 (N_2017,N_1826,N_1870);
nor U2018 (N_2018,N_1727,N_1807);
nand U2019 (N_2019,N_1833,N_1985);
and U2020 (N_2020,N_1890,N_1629);
nand U2021 (N_2021,N_1590,N_1683);
nor U2022 (N_2022,N_1919,N_1706);
xnor U2023 (N_2023,N_1508,N_1754);
xor U2024 (N_2024,N_1777,N_1996);
nand U2025 (N_2025,N_1801,N_1509);
or U2026 (N_2026,N_1970,N_1627);
xor U2027 (N_2027,N_1516,N_1607);
and U2028 (N_2028,N_1726,N_1567);
xor U2029 (N_2029,N_1959,N_1584);
and U2030 (N_2030,N_1560,N_1795);
or U2031 (N_2031,N_1735,N_1908);
nor U2032 (N_2032,N_1995,N_1591);
nand U2033 (N_2033,N_1809,N_1847);
or U2034 (N_2034,N_1934,N_1711);
and U2035 (N_2035,N_1982,N_1792);
or U2036 (N_2036,N_1917,N_1511);
nand U2037 (N_2037,N_1518,N_1834);
xor U2038 (N_2038,N_1503,N_1608);
nor U2039 (N_2039,N_1666,N_1948);
xor U2040 (N_2040,N_1913,N_1881);
or U2041 (N_2041,N_1505,N_1987);
or U2042 (N_2042,N_1656,N_1543);
nand U2043 (N_2043,N_1941,N_1615);
or U2044 (N_2044,N_1783,N_1785);
nor U2045 (N_2045,N_1760,N_1635);
and U2046 (N_2046,N_1979,N_1555);
xor U2047 (N_2047,N_1918,N_1603);
and U2048 (N_2048,N_1697,N_1710);
and U2049 (N_2049,N_1796,N_1605);
nand U2050 (N_2050,N_1977,N_1626);
xor U2051 (N_2051,N_1658,N_1874);
xor U2052 (N_2052,N_1880,N_1685);
and U2053 (N_2053,N_1581,N_1883);
or U2054 (N_2054,N_1578,N_1758);
or U2055 (N_2055,N_1851,N_1643);
xor U2056 (N_2056,N_1703,N_1850);
and U2057 (N_2057,N_1867,N_1830);
or U2058 (N_2058,N_1855,N_1765);
nand U2059 (N_2059,N_1818,N_1604);
and U2060 (N_2060,N_1642,N_1541);
and U2061 (N_2061,N_1790,N_1600);
or U2062 (N_2062,N_1576,N_1788);
xor U2063 (N_2063,N_1953,N_1708);
xor U2064 (N_2064,N_1964,N_1553);
and U2065 (N_2065,N_1749,N_1906);
or U2066 (N_2066,N_1817,N_1621);
xor U2067 (N_2067,N_1699,N_1854);
nor U2068 (N_2068,N_1848,N_1610);
and U2069 (N_2069,N_1927,N_1701);
or U2070 (N_2070,N_1771,N_1939);
and U2071 (N_2071,N_1596,N_1958);
nand U2072 (N_2072,N_1779,N_1533);
nand U2073 (N_2073,N_1672,N_1641);
nand U2074 (N_2074,N_1993,N_1510);
and U2075 (N_2075,N_1989,N_1821);
and U2076 (N_2076,N_1942,N_1716);
and U2077 (N_2077,N_1574,N_1690);
or U2078 (N_2078,N_1824,N_1732);
and U2079 (N_2079,N_1620,N_1704);
or U2080 (N_2080,N_1962,N_1684);
or U2081 (N_2081,N_1956,N_1525);
or U2082 (N_2082,N_1748,N_1705);
and U2083 (N_2083,N_1857,N_1951);
nor U2084 (N_2084,N_1844,N_1924);
and U2085 (N_2085,N_1994,N_1647);
or U2086 (N_2086,N_1831,N_1967);
or U2087 (N_2087,N_1501,N_1973);
and U2088 (N_2088,N_1843,N_1873);
nor U2089 (N_2089,N_1770,N_1823);
or U2090 (N_2090,N_1529,N_1902);
nor U2091 (N_2091,N_1827,N_1618);
or U2092 (N_2092,N_1715,N_1677);
nand U2093 (N_2093,N_1839,N_1721);
and U2094 (N_2094,N_1500,N_1720);
xor U2095 (N_2095,N_1805,N_1628);
xor U2096 (N_2096,N_1592,N_1546);
nand U2097 (N_2097,N_1651,N_1587);
or U2098 (N_2098,N_1955,N_1523);
nand U2099 (N_2099,N_1856,N_1661);
xor U2100 (N_2100,N_1864,N_1986);
nor U2101 (N_2101,N_1582,N_1815);
nand U2102 (N_2102,N_1935,N_1655);
or U2103 (N_2103,N_1717,N_1691);
and U2104 (N_2104,N_1804,N_1686);
nor U2105 (N_2105,N_1997,N_1526);
or U2106 (N_2106,N_1909,N_1719);
nand U2107 (N_2107,N_1916,N_1838);
xor U2108 (N_2108,N_1766,N_1812);
xor U2109 (N_2109,N_1822,N_1921);
or U2110 (N_2110,N_1550,N_1876);
nor U2111 (N_2111,N_1502,N_1957);
nand U2112 (N_2112,N_1961,N_1965);
or U2113 (N_2113,N_1789,N_1580);
nand U2114 (N_2114,N_1863,N_1910);
nor U2115 (N_2115,N_1534,N_1858);
xor U2116 (N_2116,N_1861,N_1619);
nor U2117 (N_2117,N_1769,N_1527);
or U2118 (N_2118,N_1729,N_1852);
nor U2119 (N_2119,N_1682,N_1936);
xnor U2120 (N_2120,N_1901,N_1507);
nor U2121 (N_2121,N_1520,N_1938);
xor U2122 (N_2122,N_1894,N_1696);
and U2123 (N_2123,N_1506,N_1586);
xnor U2124 (N_2124,N_1798,N_1800);
xor U2125 (N_2125,N_1637,N_1725);
nand U2126 (N_2126,N_1663,N_1613);
nand U2127 (N_2127,N_1521,N_1875);
xor U2128 (N_2128,N_1673,N_1778);
or U2129 (N_2129,N_1519,N_1745);
xnor U2130 (N_2130,N_1791,N_1888);
nor U2131 (N_2131,N_1943,N_1814);
xnor U2132 (N_2132,N_1776,N_1653);
nor U2133 (N_2133,N_1923,N_1907);
or U2134 (N_2134,N_1899,N_1537);
nand U2135 (N_2135,N_1531,N_1517);
nor U2136 (N_2136,N_1669,N_1885);
or U2137 (N_2137,N_1564,N_1872);
nor U2138 (N_2138,N_1750,N_1693);
xnor U2139 (N_2139,N_1535,N_1638);
and U2140 (N_2140,N_1976,N_1657);
and U2141 (N_2141,N_1540,N_1879);
nor U2142 (N_2142,N_1835,N_1536);
xnor U2143 (N_2143,N_1860,N_1636);
nand U2144 (N_2144,N_1676,N_1538);
nor U2145 (N_2145,N_1594,N_1554);
nor U2146 (N_2146,N_1579,N_1904);
nor U2147 (N_2147,N_1674,N_1900);
or U2148 (N_2148,N_1782,N_1869);
and U2149 (N_2149,N_1645,N_1816);
xor U2150 (N_2150,N_1640,N_1772);
nand U2151 (N_2151,N_1794,N_1755);
or U2152 (N_2152,N_1650,N_1742);
nor U2153 (N_2153,N_1671,N_1648);
nor U2154 (N_2154,N_1700,N_1926);
or U2155 (N_2155,N_1723,N_1713);
nand U2156 (N_2156,N_1552,N_1692);
and U2157 (N_2157,N_1606,N_1895);
and U2158 (N_2158,N_1998,N_1945);
and U2159 (N_2159,N_1722,N_1966);
xnor U2160 (N_2160,N_1634,N_1802);
nor U2161 (N_2161,N_1547,N_1625);
and U2162 (N_2162,N_1797,N_1744);
xnor U2163 (N_2163,N_1545,N_1665);
nand U2164 (N_2164,N_1695,N_1687);
and U2165 (N_2165,N_1978,N_1763);
xor U2166 (N_2166,N_1549,N_1787);
nand U2167 (N_2167,N_1712,N_1746);
xor U2168 (N_2168,N_1905,N_1612);
nor U2169 (N_2169,N_1846,N_1731);
or U2170 (N_2170,N_1999,N_1922);
and U2171 (N_2171,N_1565,N_1522);
nor U2172 (N_2172,N_1639,N_1753);
nand U2173 (N_2173,N_1609,N_1557);
or U2174 (N_2174,N_1601,N_1532);
xor U2175 (N_2175,N_1762,N_1781);
and U2176 (N_2176,N_1950,N_1736);
or U2177 (N_2177,N_1597,N_1929);
or U2178 (N_2178,N_1733,N_1990);
and U2179 (N_2179,N_1914,N_1862);
nand U2180 (N_2180,N_1984,N_1868);
nor U2181 (N_2181,N_1893,N_1896);
and U2182 (N_2182,N_1739,N_1940);
nand U2183 (N_2183,N_1614,N_1630);
and U2184 (N_2184,N_1903,N_1842);
or U2185 (N_2185,N_1622,N_1963);
or U2186 (N_2186,N_1968,N_1756);
and U2187 (N_2187,N_1911,N_1515);
nand U2188 (N_2188,N_1980,N_1780);
nand U2189 (N_2189,N_1946,N_1757);
or U2190 (N_2190,N_1678,N_1949);
xnor U2191 (N_2191,N_1664,N_1784);
nor U2192 (N_2192,N_1747,N_1539);
and U2193 (N_2193,N_1829,N_1889);
and U2194 (N_2194,N_1877,N_1932);
nand U2195 (N_2195,N_1933,N_1925);
and U2196 (N_2196,N_1786,N_1944);
or U2197 (N_2197,N_1595,N_1882);
nand U2198 (N_2198,N_1806,N_1811);
and U2199 (N_2199,N_1912,N_1570);
or U2200 (N_2200,N_1859,N_1819);
nor U2201 (N_2201,N_1808,N_1577);
xor U2202 (N_2202,N_1514,N_1849);
nand U2203 (N_2203,N_1575,N_1589);
nand U2204 (N_2204,N_1743,N_1667);
or U2205 (N_2205,N_1954,N_1698);
xnor U2206 (N_2206,N_1974,N_1513);
xor U2207 (N_2207,N_1752,N_1707);
nand U2208 (N_2208,N_1983,N_1845);
xnor U2209 (N_2209,N_1799,N_1599);
nand U2210 (N_2210,N_1654,N_1689);
and U2211 (N_2211,N_1887,N_1573);
and U2212 (N_2212,N_1688,N_1730);
or U2213 (N_2213,N_1593,N_1878);
or U2214 (N_2214,N_1644,N_1544);
nand U2215 (N_2215,N_1714,N_1866);
or U2216 (N_2216,N_1915,N_1865);
or U2217 (N_2217,N_1931,N_1832);
nand U2218 (N_2218,N_1558,N_1670);
xnor U2219 (N_2219,N_1853,N_1836);
or U2220 (N_2220,N_1598,N_1810);
nand U2221 (N_2221,N_1569,N_1793);
and U2222 (N_2222,N_1611,N_1891);
xor U2223 (N_2223,N_1988,N_1633);
or U2224 (N_2224,N_1971,N_1803);
nand U2225 (N_2225,N_1504,N_1679);
nor U2226 (N_2226,N_1616,N_1724);
or U2227 (N_2227,N_1588,N_1585);
and U2228 (N_2228,N_1524,N_1559);
or U2229 (N_2229,N_1571,N_1659);
or U2230 (N_2230,N_1528,N_1767);
nand U2231 (N_2231,N_1841,N_1728);
nand U2232 (N_2232,N_1820,N_1898);
nor U2233 (N_2233,N_1991,N_1568);
nand U2234 (N_2234,N_1773,N_1960);
xnor U2235 (N_2235,N_1562,N_1759);
nor U2236 (N_2236,N_1775,N_1737);
or U2237 (N_2237,N_1972,N_1512);
and U2238 (N_2238,N_1660,N_1952);
nor U2239 (N_2239,N_1662,N_1828);
xnor U2240 (N_2240,N_1947,N_1871);
xnor U2241 (N_2241,N_1930,N_1551);
or U2242 (N_2242,N_1740,N_1548);
nor U2243 (N_2243,N_1702,N_1572);
nor U2244 (N_2244,N_1694,N_1813);
and U2245 (N_2245,N_1892,N_1617);
nor U2246 (N_2246,N_1530,N_1556);
xor U2247 (N_2247,N_1675,N_1624);
xor U2248 (N_2248,N_1652,N_1768);
nor U2249 (N_2249,N_1738,N_1602);
or U2250 (N_2250,N_1786,N_1559);
nand U2251 (N_2251,N_1978,N_1958);
nand U2252 (N_2252,N_1847,N_1542);
nor U2253 (N_2253,N_1574,N_1614);
xnor U2254 (N_2254,N_1620,N_1559);
xnor U2255 (N_2255,N_1963,N_1691);
nand U2256 (N_2256,N_1945,N_1770);
nand U2257 (N_2257,N_1856,N_1877);
or U2258 (N_2258,N_1919,N_1953);
nor U2259 (N_2259,N_1697,N_1867);
and U2260 (N_2260,N_1564,N_1509);
nand U2261 (N_2261,N_1551,N_1640);
nand U2262 (N_2262,N_1883,N_1629);
and U2263 (N_2263,N_1906,N_1977);
and U2264 (N_2264,N_1903,N_1661);
xnor U2265 (N_2265,N_1542,N_1731);
nand U2266 (N_2266,N_1740,N_1697);
xor U2267 (N_2267,N_1599,N_1832);
nor U2268 (N_2268,N_1697,N_1983);
xnor U2269 (N_2269,N_1781,N_1828);
and U2270 (N_2270,N_1735,N_1692);
and U2271 (N_2271,N_1690,N_1525);
xnor U2272 (N_2272,N_1876,N_1996);
and U2273 (N_2273,N_1706,N_1650);
and U2274 (N_2274,N_1815,N_1535);
nand U2275 (N_2275,N_1980,N_1954);
and U2276 (N_2276,N_1890,N_1547);
nand U2277 (N_2277,N_1850,N_1773);
nor U2278 (N_2278,N_1858,N_1631);
nor U2279 (N_2279,N_1974,N_1900);
or U2280 (N_2280,N_1810,N_1597);
xnor U2281 (N_2281,N_1780,N_1964);
xor U2282 (N_2282,N_1889,N_1725);
or U2283 (N_2283,N_1517,N_1509);
and U2284 (N_2284,N_1737,N_1788);
or U2285 (N_2285,N_1965,N_1935);
nor U2286 (N_2286,N_1894,N_1741);
nand U2287 (N_2287,N_1787,N_1580);
nand U2288 (N_2288,N_1564,N_1723);
nor U2289 (N_2289,N_1661,N_1916);
xnor U2290 (N_2290,N_1787,N_1509);
xor U2291 (N_2291,N_1533,N_1973);
nor U2292 (N_2292,N_1840,N_1807);
or U2293 (N_2293,N_1560,N_1596);
nand U2294 (N_2294,N_1783,N_1723);
and U2295 (N_2295,N_1580,N_1664);
xor U2296 (N_2296,N_1530,N_1633);
xor U2297 (N_2297,N_1952,N_1587);
or U2298 (N_2298,N_1617,N_1914);
or U2299 (N_2299,N_1845,N_1754);
or U2300 (N_2300,N_1656,N_1752);
nand U2301 (N_2301,N_1765,N_1806);
or U2302 (N_2302,N_1971,N_1635);
xnor U2303 (N_2303,N_1803,N_1657);
nand U2304 (N_2304,N_1822,N_1775);
and U2305 (N_2305,N_1712,N_1519);
xor U2306 (N_2306,N_1604,N_1787);
or U2307 (N_2307,N_1678,N_1523);
xnor U2308 (N_2308,N_1717,N_1945);
xnor U2309 (N_2309,N_1700,N_1568);
or U2310 (N_2310,N_1992,N_1916);
nand U2311 (N_2311,N_1859,N_1515);
nor U2312 (N_2312,N_1580,N_1701);
nor U2313 (N_2313,N_1504,N_1874);
or U2314 (N_2314,N_1841,N_1869);
xor U2315 (N_2315,N_1614,N_1632);
or U2316 (N_2316,N_1911,N_1809);
or U2317 (N_2317,N_1793,N_1588);
xnor U2318 (N_2318,N_1951,N_1800);
or U2319 (N_2319,N_1634,N_1964);
xor U2320 (N_2320,N_1652,N_1756);
or U2321 (N_2321,N_1716,N_1811);
or U2322 (N_2322,N_1967,N_1544);
xnor U2323 (N_2323,N_1971,N_1591);
and U2324 (N_2324,N_1536,N_1710);
xnor U2325 (N_2325,N_1582,N_1546);
nor U2326 (N_2326,N_1927,N_1634);
and U2327 (N_2327,N_1827,N_1697);
nor U2328 (N_2328,N_1625,N_1991);
and U2329 (N_2329,N_1612,N_1708);
nor U2330 (N_2330,N_1955,N_1942);
or U2331 (N_2331,N_1683,N_1524);
nor U2332 (N_2332,N_1693,N_1780);
nor U2333 (N_2333,N_1859,N_1586);
and U2334 (N_2334,N_1741,N_1508);
nand U2335 (N_2335,N_1924,N_1709);
xor U2336 (N_2336,N_1985,N_1559);
xor U2337 (N_2337,N_1922,N_1767);
nand U2338 (N_2338,N_1661,N_1658);
xor U2339 (N_2339,N_1939,N_1602);
nor U2340 (N_2340,N_1777,N_1876);
nor U2341 (N_2341,N_1659,N_1972);
nand U2342 (N_2342,N_1843,N_1928);
nor U2343 (N_2343,N_1935,N_1842);
nand U2344 (N_2344,N_1587,N_1609);
and U2345 (N_2345,N_1768,N_1712);
or U2346 (N_2346,N_1768,N_1597);
xor U2347 (N_2347,N_1968,N_1843);
and U2348 (N_2348,N_1875,N_1868);
or U2349 (N_2349,N_1982,N_1900);
xnor U2350 (N_2350,N_1896,N_1662);
nand U2351 (N_2351,N_1761,N_1989);
nand U2352 (N_2352,N_1965,N_1511);
or U2353 (N_2353,N_1938,N_1837);
nor U2354 (N_2354,N_1829,N_1520);
and U2355 (N_2355,N_1530,N_1542);
nor U2356 (N_2356,N_1612,N_1908);
or U2357 (N_2357,N_1693,N_1762);
and U2358 (N_2358,N_1765,N_1676);
and U2359 (N_2359,N_1916,N_1515);
or U2360 (N_2360,N_1620,N_1880);
and U2361 (N_2361,N_1728,N_1545);
nand U2362 (N_2362,N_1749,N_1860);
nand U2363 (N_2363,N_1697,N_1892);
nor U2364 (N_2364,N_1572,N_1845);
or U2365 (N_2365,N_1560,N_1659);
xnor U2366 (N_2366,N_1808,N_1532);
nor U2367 (N_2367,N_1549,N_1506);
xnor U2368 (N_2368,N_1780,N_1760);
and U2369 (N_2369,N_1954,N_1890);
nor U2370 (N_2370,N_1991,N_1689);
and U2371 (N_2371,N_1970,N_1927);
nor U2372 (N_2372,N_1786,N_1600);
nor U2373 (N_2373,N_1665,N_1959);
and U2374 (N_2374,N_1605,N_1746);
xor U2375 (N_2375,N_1773,N_1711);
nand U2376 (N_2376,N_1572,N_1794);
or U2377 (N_2377,N_1902,N_1680);
and U2378 (N_2378,N_1758,N_1968);
xor U2379 (N_2379,N_1942,N_1702);
nor U2380 (N_2380,N_1730,N_1853);
nor U2381 (N_2381,N_1504,N_1970);
and U2382 (N_2382,N_1697,N_1797);
and U2383 (N_2383,N_1987,N_1629);
or U2384 (N_2384,N_1674,N_1845);
nand U2385 (N_2385,N_1842,N_1675);
nor U2386 (N_2386,N_1520,N_1543);
and U2387 (N_2387,N_1617,N_1962);
xnor U2388 (N_2388,N_1893,N_1761);
nor U2389 (N_2389,N_1826,N_1567);
or U2390 (N_2390,N_1644,N_1859);
or U2391 (N_2391,N_1699,N_1537);
or U2392 (N_2392,N_1987,N_1795);
xor U2393 (N_2393,N_1865,N_1666);
and U2394 (N_2394,N_1874,N_1665);
and U2395 (N_2395,N_1525,N_1806);
and U2396 (N_2396,N_1594,N_1908);
and U2397 (N_2397,N_1574,N_1711);
or U2398 (N_2398,N_1573,N_1562);
nand U2399 (N_2399,N_1989,N_1548);
or U2400 (N_2400,N_1592,N_1698);
nor U2401 (N_2401,N_1903,N_1836);
or U2402 (N_2402,N_1914,N_1596);
and U2403 (N_2403,N_1752,N_1574);
and U2404 (N_2404,N_1598,N_1868);
and U2405 (N_2405,N_1593,N_1504);
nand U2406 (N_2406,N_1741,N_1583);
nand U2407 (N_2407,N_1573,N_1953);
or U2408 (N_2408,N_1879,N_1971);
nand U2409 (N_2409,N_1664,N_1850);
nor U2410 (N_2410,N_1652,N_1649);
or U2411 (N_2411,N_1558,N_1876);
nand U2412 (N_2412,N_1904,N_1920);
or U2413 (N_2413,N_1517,N_1784);
or U2414 (N_2414,N_1966,N_1536);
or U2415 (N_2415,N_1965,N_1714);
xnor U2416 (N_2416,N_1746,N_1771);
or U2417 (N_2417,N_1615,N_1737);
and U2418 (N_2418,N_1904,N_1761);
nand U2419 (N_2419,N_1563,N_1612);
nand U2420 (N_2420,N_1621,N_1526);
nand U2421 (N_2421,N_1587,N_1510);
or U2422 (N_2422,N_1970,N_1509);
xor U2423 (N_2423,N_1619,N_1791);
and U2424 (N_2424,N_1527,N_1681);
and U2425 (N_2425,N_1553,N_1640);
or U2426 (N_2426,N_1972,N_1996);
nor U2427 (N_2427,N_1845,N_1631);
nor U2428 (N_2428,N_1743,N_1885);
or U2429 (N_2429,N_1546,N_1527);
and U2430 (N_2430,N_1561,N_1850);
nand U2431 (N_2431,N_1920,N_1653);
xnor U2432 (N_2432,N_1724,N_1572);
xnor U2433 (N_2433,N_1937,N_1949);
or U2434 (N_2434,N_1707,N_1655);
and U2435 (N_2435,N_1944,N_1867);
or U2436 (N_2436,N_1908,N_1681);
or U2437 (N_2437,N_1577,N_1705);
xnor U2438 (N_2438,N_1917,N_1550);
or U2439 (N_2439,N_1786,N_1529);
nand U2440 (N_2440,N_1602,N_1622);
or U2441 (N_2441,N_1970,N_1632);
or U2442 (N_2442,N_1807,N_1920);
xnor U2443 (N_2443,N_1559,N_1596);
xor U2444 (N_2444,N_1569,N_1600);
nand U2445 (N_2445,N_1546,N_1839);
or U2446 (N_2446,N_1579,N_1897);
and U2447 (N_2447,N_1567,N_1519);
xor U2448 (N_2448,N_1964,N_1528);
nor U2449 (N_2449,N_1947,N_1646);
and U2450 (N_2450,N_1580,N_1925);
nor U2451 (N_2451,N_1867,N_1677);
nand U2452 (N_2452,N_1720,N_1782);
xnor U2453 (N_2453,N_1656,N_1896);
nor U2454 (N_2454,N_1938,N_1956);
and U2455 (N_2455,N_1754,N_1678);
xnor U2456 (N_2456,N_1691,N_1650);
nor U2457 (N_2457,N_1728,N_1667);
nor U2458 (N_2458,N_1764,N_1511);
nor U2459 (N_2459,N_1883,N_1708);
or U2460 (N_2460,N_1690,N_1609);
nand U2461 (N_2461,N_1647,N_1574);
or U2462 (N_2462,N_1572,N_1554);
and U2463 (N_2463,N_1787,N_1903);
xnor U2464 (N_2464,N_1669,N_1943);
nand U2465 (N_2465,N_1830,N_1754);
or U2466 (N_2466,N_1802,N_1738);
nor U2467 (N_2467,N_1838,N_1614);
nand U2468 (N_2468,N_1613,N_1825);
and U2469 (N_2469,N_1513,N_1747);
or U2470 (N_2470,N_1509,N_1875);
nor U2471 (N_2471,N_1779,N_1693);
xor U2472 (N_2472,N_1805,N_1973);
nand U2473 (N_2473,N_1573,N_1663);
and U2474 (N_2474,N_1787,N_1657);
nor U2475 (N_2475,N_1822,N_1909);
nor U2476 (N_2476,N_1691,N_1855);
or U2477 (N_2477,N_1977,N_1662);
nor U2478 (N_2478,N_1889,N_1546);
or U2479 (N_2479,N_1956,N_1824);
or U2480 (N_2480,N_1585,N_1633);
nor U2481 (N_2481,N_1786,N_1590);
nand U2482 (N_2482,N_1792,N_1757);
or U2483 (N_2483,N_1937,N_1555);
xor U2484 (N_2484,N_1816,N_1669);
nand U2485 (N_2485,N_1507,N_1759);
nand U2486 (N_2486,N_1732,N_1522);
xor U2487 (N_2487,N_1578,N_1946);
or U2488 (N_2488,N_1977,N_1958);
xor U2489 (N_2489,N_1748,N_1861);
xor U2490 (N_2490,N_1804,N_1920);
xor U2491 (N_2491,N_1554,N_1652);
or U2492 (N_2492,N_1780,N_1664);
xor U2493 (N_2493,N_1700,N_1860);
nor U2494 (N_2494,N_1859,N_1676);
nor U2495 (N_2495,N_1584,N_1800);
xnor U2496 (N_2496,N_1568,N_1556);
or U2497 (N_2497,N_1786,N_1524);
or U2498 (N_2498,N_1550,N_1793);
and U2499 (N_2499,N_1660,N_1901);
nor U2500 (N_2500,N_2203,N_2097);
or U2501 (N_2501,N_2155,N_2244);
nor U2502 (N_2502,N_2405,N_2284);
or U2503 (N_2503,N_2006,N_2471);
nor U2504 (N_2504,N_2032,N_2236);
xor U2505 (N_2505,N_2337,N_2490);
nand U2506 (N_2506,N_2468,N_2260);
nor U2507 (N_2507,N_2355,N_2197);
and U2508 (N_2508,N_2073,N_2251);
or U2509 (N_2509,N_2220,N_2011);
nor U2510 (N_2510,N_2333,N_2198);
and U2511 (N_2511,N_2283,N_2301);
or U2512 (N_2512,N_2314,N_2353);
nor U2513 (N_2513,N_2361,N_2122);
nor U2514 (N_2514,N_2018,N_2201);
nand U2515 (N_2515,N_2208,N_2446);
nand U2516 (N_2516,N_2484,N_2033);
nor U2517 (N_2517,N_2436,N_2210);
nand U2518 (N_2518,N_2108,N_2420);
xnor U2519 (N_2519,N_2266,N_2163);
nor U2520 (N_2520,N_2076,N_2124);
nor U2521 (N_2521,N_2125,N_2000);
xnor U2522 (N_2522,N_2069,N_2085);
nand U2523 (N_2523,N_2037,N_2106);
and U2524 (N_2524,N_2185,N_2116);
xnor U2525 (N_2525,N_2055,N_2336);
nand U2526 (N_2526,N_2335,N_2448);
or U2527 (N_2527,N_2499,N_2056);
nor U2528 (N_2528,N_2217,N_2365);
or U2529 (N_2529,N_2144,N_2092);
nand U2530 (N_2530,N_2035,N_2271);
nor U2531 (N_2531,N_2231,N_2014);
nor U2532 (N_2532,N_2247,N_2312);
xnor U2533 (N_2533,N_2078,N_2239);
xor U2534 (N_2534,N_2046,N_2051);
nor U2535 (N_2535,N_2215,N_2151);
nand U2536 (N_2536,N_2091,N_2386);
or U2537 (N_2537,N_2118,N_2315);
or U2538 (N_2538,N_2299,N_2346);
or U2539 (N_2539,N_2443,N_2395);
nor U2540 (N_2540,N_2376,N_2235);
xnor U2541 (N_2541,N_2470,N_2173);
and U2542 (N_2542,N_2067,N_2227);
nor U2543 (N_2543,N_2149,N_2019);
xnor U2544 (N_2544,N_2045,N_2318);
and U2545 (N_2545,N_2322,N_2321);
and U2546 (N_2546,N_2021,N_2358);
nor U2547 (N_2547,N_2370,N_2418);
xor U2548 (N_2548,N_2205,N_2063);
nand U2549 (N_2549,N_2096,N_2160);
or U2550 (N_2550,N_2427,N_2042);
nor U2551 (N_2551,N_2012,N_2473);
nand U2552 (N_2552,N_2372,N_2306);
nand U2553 (N_2553,N_2466,N_2123);
xnor U2554 (N_2554,N_2478,N_2364);
nor U2555 (N_2555,N_2302,N_2411);
and U2556 (N_2556,N_2022,N_2360);
nand U2557 (N_2557,N_2325,N_2457);
nor U2558 (N_2558,N_2451,N_2406);
and U2559 (N_2559,N_2342,N_2391);
and U2560 (N_2560,N_2297,N_2437);
nand U2561 (N_2561,N_2435,N_2417);
xnor U2562 (N_2562,N_2463,N_2054);
nand U2563 (N_2563,N_2485,N_2319);
nand U2564 (N_2564,N_2390,N_2275);
and U2565 (N_2565,N_2426,N_2273);
nand U2566 (N_2566,N_2348,N_2261);
xnor U2567 (N_2567,N_2379,N_2290);
xnor U2568 (N_2568,N_2059,N_2289);
nand U2569 (N_2569,N_2385,N_2262);
xor U2570 (N_2570,N_2147,N_2060);
and U2571 (N_2571,N_2267,N_2025);
nor U2572 (N_2572,N_2193,N_2121);
nor U2573 (N_2573,N_2387,N_2071);
xnor U2574 (N_2574,N_2214,N_2162);
and U2575 (N_2575,N_2438,N_2334);
or U2576 (N_2576,N_2199,N_2008);
xnor U2577 (N_2577,N_2324,N_2007);
xnor U2578 (N_2578,N_2410,N_2287);
xor U2579 (N_2579,N_2292,N_2344);
nor U2580 (N_2580,N_2282,N_2293);
nand U2581 (N_2581,N_2294,N_2304);
nand U2582 (N_2582,N_2475,N_2039);
xnor U2583 (N_2583,N_2206,N_2066);
and U2584 (N_2584,N_2137,N_2087);
xnor U2585 (N_2585,N_2493,N_2279);
xnor U2586 (N_2586,N_2223,N_2209);
and U2587 (N_2587,N_2101,N_2442);
nand U2588 (N_2588,N_2157,N_2452);
or U2589 (N_2589,N_2238,N_2113);
or U2590 (N_2590,N_2168,N_2093);
and U2591 (N_2591,N_2053,N_2183);
nor U2592 (N_2592,N_2119,N_2187);
and U2593 (N_2593,N_2002,N_2152);
nand U2594 (N_2594,N_2171,N_2276);
and U2595 (N_2595,N_2347,N_2425);
xnor U2596 (N_2596,N_2256,N_2178);
and U2597 (N_2597,N_2422,N_2009);
and U2598 (N_2598,N_2479,N_2459);
and U2599 (N_2599,N_2225,N_2083);
nor U2600 (N_2600,N_2296,N_2146);
nor U2601 (N_2601,N_2270,N_2281);
nor U2602 (N_2602,N_2481,N_2246);
or U2603 (N_2603,N_2132,N_2382);
nand U2604 (N_2604,N_2100,N_2028);
nand U2605 (N_2605,N_2213,N_2449);
and U2606 (N_2606,N_2263,N_2234);
nor U2607 (N_2607,N_2090,N_2222);
nand U2608 (N_2608,N_2305,N_2327);
nor U2609 (N_2609,N_2064,N_2415);
nand U2610 (N_2610,N_2068,N_2228);
and U2611 (N_2611,N_2313,N_2316);
and U2612 (N_2612,N_2062,N_2182);
nor U2613 (N_2613,N_2001,N_2403);
nand U2614 (N_2614,N_2111,N_2052);
nor U2615 (N_2615,N_2419,N_2476);
and U2616 (N_2616,N_2170,N_2202);
nor U2617 (N_2617,N_2191,N_2458);
or U2618 (N_2618,N_2491,N_2127);
and U2619 (N_2619,N_2095,N_2080);
nand U2620 (N_2620,N_2268,N_2207);
xor U2621 (N_2621,N_2138,N_2444);
xor U2622 (N_2622,N_2079,N_2194);
or U2623 (N_2623,N_2140,N_2243);
and U2624 (N_2624,N_2176,N_2329);
nand U2625 (N_2625,N_2134,N_2130);
nand U2626 (N_2626,N_2392,N_2255);
or U2627 (N_2627,N_2323,N_2226);
xor U2628 (N_2628,N_2303,N_2274);
nor U2629 (N_2629,N_2402,N_2328);
xnor U2630 (N_2630,N_2082,N_2003);
or U2631 (N_2631,N_2399,N_2024);
xor U2632 (N_2632,N_2421,N_2423);
or U2633 (N_2633,N_2343,N_2005);
and U2634 (N_2634,N_2020,N_2248);
nand U2635 (N_2635,N_2483,N_2110);
or U2636 (N_2636,N_2269,N_2249);
xnor U2637 (N_2637,N_2326,N_2285);
xor U2638 (N_2638,N_2219,N_2258);
nand U2639 (N_2639,N_2161,N_2181);
or U2640 (N_2640,N_2142,N_2397);
and U2641 (N_2641,N_2345,N_2363);
nor U2642 (N_2642,N_2156,N_2034);
xnor U2643 (N_2643,N_2331,N_2041);
nor U2644 (N_2644,N_2272,N_2004);
or U2645 (N_2645,N_2357,N_2145);
xor U2646 (N_2646,N_2309,N_2413);
nor U2647 (N_2647,N_2043,N_2280);
nor U2648 (N_2648,N_2186,N_2240);
xnor U2649 (N_2649,N_2494,N_2307);
xnor U2650 (N_2650,N_2467,N_2434);
and U2651 (N_2651,N_2167,N_2254);
and U2652 (N_2652,N_2013,N_2378);
nand U2653 (N_2653,N_2453,N_2031);
nand U2654 (N_2654,N_2218,N_2356);
and U2655 (N_2655,N_2172,N_2371);
or U2656 (N_2656,N_2424,N_2384);
xor U2657 (N_2657,N_2373,N_2441);
and U2658 (N_2658,N_2115,N_2350);
and U2659 (N_2659,N_2396,N_2158);
nor U2660 (N_2660,N_2368,N_2094);
or U2661 (N_2661,N_2196,N_2221);
and U2662 (N_2662,N_2088,N_2401);
xor U2663 (N_2663,N_2474,N_2128);
xnor U2664 (N_2664,N_2291,N_2232);
or U2665 (N_2665,N_2259,N_2278);
or U2666 (N_2666,N_2489,N_2166);
nand U2667 (N_2667,N_2252,N_2131);
or U2668 (N_2668,N_2389,N_2109);
or U2669 (N_2669,N_2461,N_2180);
nor U2670 (N_2670,N_2135,N_2086);
nand U2671 (N_2671,N_2129,N_2414);
nand U2672 (N_2672,N_2233,N_2027);
nand U2673 (N_2673,N_2098,N_2174);
or U2674 (N_2674,N_2044,N_2114);
nor U2675 (N_2675,N_2099,N_2430);
nor U2676 (N_2676,N_2036,N_2143);
or U2677 (N_2677,N_2105,N_2250);
and U2678 (N_2678,N_2230,N_2469);
nor U2679 (N_2679,N_2184,N_2341);
xnor U2680 (N_2680,N_2159,N_2126);
xor U2681 (N_2681,N_2015,N_2447);
xor U2682 (N_2682,N_2089,N_2030);
nor U2683 (N_2683,N_2487,N_2047);
or U2684 (N_2684,N_2317,N_2103);
or U2685 (N_2685,N_2454,N_2477);
and U2686 (N_2686,N_2058,N_2374);
and U2687 (N_2687,N_2048,N_2486);
and U2688 (N_2688,N_2456,N_2311);
xor U2689 (N_2689,N_2351,N_2288);
xor U2690 (N_2690,N_2308,N_2264);
xor U2691 (N_2691,N_2084,N_2366);
or U2692 (N_2692,N_2412,N_2102);
nor U2693 (N_2693,N_2165,N_2429);
or U2694 (N_2694,N_2211,N_2029);
xnor U2695 (N_2695,N_2455,N_2359);
or U2696 (N_2696,N_2295,N_2237);
and U2697 (N_2697,N_2192,N_2398);
nand U2698 (N_2698,N_2440,N_2388);
nor U2699 (N_2699,N_2367,N_2408);
and U2700 (N_2700,N_2061,N_2383);
nand U2701 (N_2701,N_2409,N_2349);
and U2702 (N_2702,N_2375,N_2298);
nand U2703 (N_2703,N_2286,N_2016);
xor U2704 (N_2704,N_2179,N_2362);
or U2705 (N_2705,N_2050,N_2393);
or U2706 (N_2706,N_2017,N_2104);
nand U2707 (N_2707,N_2169,N_2204);
or U2708 (N_2708,N_2465,N_2265);
and U2709 (N_2709,N_2190,N_2075);
or U2710 (N_2710,N_2300,N_2010);
nor U2711 (N_2711,N_2112,N_2332);
or U2712 (N_2712,N_2216,N_2462);
xor U2713 (N_2713,N_2340,N_2150);
xor U2714 (N_2714,N_2394,N_2139);
nand U2715 (N_2715,N_2141,N_2177);
nor U2716 (N_2716,N_2472,N_2040);
xor U2717 (N_2717,N_2339,N_2492);
or U2718 (N_2718,N_2154,N_2038);
or U2719 (N_2719,N_2338,N_2354);
xnor U2720 (N_2720,N_2212,N_2107);
nor U2721 (N_2721,N_2369,N_2133);
xnor U2722 (N_2722,N_2070,N_2242);
nor U2723 (N_2723,N_2428,N_2377);
nor U2724 (N_2724,N_2195,N_2495);
and U2725 (N_2725,N_2431,N_2120);
and U2726 (N_2726,N_2416,N_2320);
or U2727 (N_2727,N_2241,N_2049);
and U2728 (N_2728,N_2445,N_2257);
or U2729 (N_2729,N_2432,N_2074);
or U2730 (N_2730,N_2072,N_2057);
nand U2731 (N_2731,N_2407,N_2188);
or U2732 (N_2732,N_2433,N_2330);
or U2733 (N_2733,N_2117,N_2148);
nor U2734 (N_2734,N_2023,N_2497);
nor U2735 (N_2735,N_2189,N_2439);
or U2736 (N_2736,N_2381,N_2065);
and U2737 (N_2737,N_2480,N_2498);
nor U2738 (N_2738,N_2464,N_2460);
xor U2739 (N_2739,N_2136,N_2450);
nand U2740 (N_2740,N_2229,N_2164);
nand U2741 (N_2741,N_2400,N_2077);
or U2742 (N_2742,N_2277,N_2224);
nand U2743 (N_2743,N_2081,N_2496);
nor U2744 (N_2744,N_2245,N_2352);
nor U2745 (N_2745,N_2153,N_2253);
and U2746 (N_2746,N_2310,N_2482);
or U2747 (N_2747,N_2404,N_2200);
xor U2748 (N_2748,N_2380,N_2175);
and U2749 (N_2749,N_2488,N_2026);
nor U2750 (N_2750,N_2087,N_2398);
and U2751 (N_2751,N_2233,N_2341);
nand U2752 (N_2752,N_2432,N_2137);
or U2753 (N_2753,N_2162,N_2132);
nand U2754 (N_2754,N_2012,N_2300);
and U2755 (N_2755,N_2029,N_2043);
or U2756 (N_2756,N_2097,N_2357);
nor U2757 (N_2757,N_2467,N_2449);
nor U2758 (N_2758,N_2216,N_2379);
or U2759 (N_2759,N_2362,N_2185);
and U2760 (N_2760,N_2405,N_2346);
nor U2761 (N_2761,N_2080,N_2050);
nand U2762 (N_2762,N_2020,N_2494);
and U2763 (N_2763,N_2444,N_2203);
and U2764 (N_2764,N_2017,N_2257);
nand U2765 (N_2765,N_2021,N_2298);
nand U2766 (N_2766,N_2219,N_2106);
nand U2767 (N_2767,N_2169,N_2348);
nand U2768 (N_2768,N_2196,N_2380);
xor U2769 (N_2769,N_2307,N_2160);
xor U2770 (N_2770,N_2439,N_2319);
nor U2771 (N_2771,N_2107,N_2115);
or U2772 (N_2772,N_2029,N_2274);
nor U2773 (N_2773,N_2313,N_2217);
and U2774 (N_2774,N_2001,N_2186);
xnor U2775 (N_2775,N_2449,N_2283);
nor U2776 (N_2776,N_2314,N_2364);
nor U2777 (N_2777,N_2233,N_2310);
or U2778 (N_2778,N_2475,N_2371);
xor U2779 (N_2779,N_2347,N_2082);
nand U2780 (N_2780,N_2399,N_2270);
nor U2781 (N_2781,N_2436,N_2155);
xor U2782 (N_2782,N_2143,N_2482);
xor U2783 (N_2783,N_2278,N_2391);
nand U2784 (N_2784,N_2306,N_2238);
xor U2785 (N_2785,N_2343,N_2174);
nand U2786 (N_2786,N_2200,N_2108);
xnor U2787 (N_2787,N_2182,N_2165);
xnor U2788 (N_2788,N_2106,N_2430);
xor U2789 (N_2789,N_2343,N_2243);
nor U2790 (N_2790,N_2166,N_2458);
or U2791 (N_2791,N_2151,N_2238);
nor U2792 (N_2792,N_2005,N_2205);
and U2793 (N_2793,N_2342,N_2252);
nand U2794 (N_2794,N_2296,N_2401);
xnor U2795 (N_2795,N_2135,N_2109);
or U2796 (N_2796,N_2221,N_2322);
or U2797 (N_2797,N_2078,N_2464);
and U2798 (N_2798,N_2139,N_2207);
nor U2799 (N_2799,N_2007,N_2299);
nor U2800 (N_2800,N_2020,N_2206);
nand U2801 (N_2801,N_2114,N_2095);
or U2802 (N_2802,N_2367,N_2362);
nand U2803 (N_2803,N_2457,N_2203);
xnor U2804 (N_2804,N_2018,N_2314);
or U2805 (N_2805,N_2273,N_2396);
nor U2806 (N_2806,N_2286,N_2056);
xor U2807 (N_2807,N_2093,N_2001);
or U2808 (N_2808,N_2287,N_2494);
or U2809 (N_2809,N_2352,N_2425);
or U2810 (N_2810,N_2241,N_2384);
nand U2811 (N_2811,N_2234,N_2351);
xnor U2812 (N_2812,N_2306,N_2178);
nor U2813 (N_2813,N_2444,N_2078);
nor U2814 (N_2814,N_2347,N_2433);
and U2815 (N_2815,N_2389,N_2072);
or U2816 (N_2816,N_2340,N_2279);
or U2817 (N_2817,N_2367,N_2201);
or U2818 (N_2818,N_2287,N_2130);
xor U2819 (N_2819,N_2223,N_2457);
nor U2820 (N_2820,N_2321,N_2476);
xor U2821 (N_2821,N_2485,N_2009);
or U2822 (N_2822,N_2053,N_2363);
and U2823 (N_2823,N_2408,N_2240);
nor U2824 (N_2824,N_2198,N_2143);
xnor U2825 (N_2825,N_2213,N_2188);
and U2826 (N_2826,N_2107,N_2457);
and U2827 (N_2827,N_2073,N_2169);
nor U2828 (N_2828,N_2007,N_2244);
xor U2829 (N_2829,N_2102,N_2326);
nor U2830 (N_2830,N_2018,N_2260);
or U2831 (N_2831,N_2215,N_2251);
nand U2832 (N_2832,N_2143,N_2159);
or U2833 (N_2833,N_2320,N_2361);
nand U2834 (N_2834,N_2407,N_2009);
nor U2835 (N_2835,N_2029,N_2214);
nand U2836 (N_2836,N_2495,N_2192);
nand U2837 (N_2837,N_2278,N_2199);
or U2838 (N_2838,N_2111,N_2061);
or U2839 (N_2839,N_2443,N_2091);
xor U2840 (N_2840,N_2288,N_2199);
xnor U2841 (N_2841,N_2047,N_2271);
or U2842 (N_2842,N_2348,N_2136);
and U2843 (N_2843,N_2372,N_2284);
or U2844 (N_2844,N_2303,N_2325);
nor U2845 (N_2845,N_2325,N_2460);
and U2846 (N_2846,N_2098,N_2222);
nand U2847 (N_2847,N_2405,N_2408);
xnor U2848 (N_2848,N_2484,N_2160);
nor U2849 (N_2849,N_2461,N_2362);
nor U2850 (N_2850,N_2303,N_2308);
xnor U2851 (N_2851,N_2419,N_2455);
xnor U2852 (N_2852,N_2024,N_2068);
xnor U2853 (N_2853,N_2003,N_2473);
and U2854 (N_2854,N_2405,N_2171);
or U2855 (N_2855,N_2053,N_2331);
nor U2856 (N_2856,N_2234,N_2125);
nor U2857 (N_2857,N_2490,N_2300);
nor U2858 (N_2858,N_2380,N_2303);
nor U2859 (N_2859,N_2283,N_2398);
nor U2860 (N_2860,N_2113,N_2297);
nand U2861 (N_2861,N_2232,N_2105);
and U2862 (N_2862,N_2089,N_2263);
xnor U2863 (N_2863,N_2443,N_2268);
and U2864 (N_2864,N_2222,N_2023);
or U2865 (N_2865,N_2391,N_2141);
nand U2866 (N_2866,N_2241,N_2410);
nand U2867 (N_2867,N_2474,N_2076);
or U2868 (N_2868,N_2471,N_2344);
nor U2869 (N_2869,N_2480,N_2038);
nor U2870 (N_2870,N_2182,N_2250);
nand U2871 (N_2871,N_2044,N_2281);
nor U2872 (N_2872,N_2443,N_2345);
nor U2873 (N_2873,N_2278,N_2462);
xor U2874 (N_2874,N_2318,N_2213);
xor U2875 (N_2875,N_2443,N_2128);
nand U2876 (N_2876,N_2108,N_2170);
and U2877 (N_2877,N_2029,N_2066);
xor U2878 (N_2878,N_2303,N_2247);
and U2879 (N_2879,N_2478,N_2391);
nand U2880 (N_2880,N_2319,N_2282);
and U2881 (N_2881,N_2045,N_2080);
or U2882 (N_2882,N_2356,N_2178);
nor U2883 (N_2883,N_2382,N_2104);
and U2884 (N_2884,N_2401,N_2001);
or U2885 (N_2885,N_2482,N_2309);
nor U2886 (N_2886,N_2414,N_2209);
and U2887 (N_2887,N_2459,N_2080);
nand U2888 (N_2888,N_2491,N_2200);
or U2889 (N_2889,N_2175,N_2493);
xor U2890 (N_2890,N_2391,N_2305);
xnor U2891 (N_2891,N_2270,N_2484);
and U2892 (N_2892,N_2424,N_2237);
xor U2893 (N_2893,N_2283,N_2161);
and U2894 (N_2894,N_2166,N_2448);
nand U2895 (N_2895,N_2188,N_2324);
or U2896 (N_2896,N_2171,N_2333);
and U2897 (N_2897,N_2082,N_2171);
xor U2898 (N_2898,N_2072,N_2419);
or U2899 (N_2899,N_2257,N_2356);
and U2900 (N_2900,N_2481,N_2027);
and U2901 (N_2901,N_2140,N_2260);
xor U2902 (N_2902,N_2467,N_2231);
or U2903 (N_2903,N_2057,N_2191);
xnor U2904 (N_2904,N_2485,N_2041);
xnor U2905 (N_2905,N_2236,N_2265);
or U2906 (N_2906,N_2352,N_2269);
and U2907 (N_2907,N_2141,N_2467);
and U2908 (N_2908,N_2266,N_2242);
or U2909 (N_2909,N_2138,N_2192);
or U2910 (N_2910,N_2476,N_2110);
and U2911 (N_2911,N_2277,N_2040);
nor U2912 (N_2912,N_2244,N_2466);
nor U2913 (N_2913,N_2396,N_2274);
and U2914 (N_2914,N_2160,N_2049);
and U2915 (N_2915,N_2471,N_2152);
and U2916 (N_2916,N_2295,N_2278);
nand U2917 (N_2917,N_2357,N_2402);
nand U2918 (N_2918,N_2148,N_2401);
and U2919 (N_2919,N_2186,N_2345);
or U2920 (N_2920,N_2044,N_2299);
and U2921 (N_2921,N_2221,N_2346);
or U2922 (N_2922,N_2173,N_2493);
nor U2923 (N_2923,N_2493,N_2396);
nor U2924 (N_2924,N_2339,N_2254);
nor U2925 (N_2925,N_2099,N_2437);
nor U2926 (N_2926,N_2062,N_2274);
or U2927 (N_2927,N_2372,N_2276);
and U2928 (N_2928,N_2168,N_2328);
nor U2929 (N_2929,N_2130,N_2072);
nand U2930 (N_2930,N_2262,N_2100);
nand U2931 (N_2931,N_2440,N_2152);
nand U2932 (N_2932,N_2073,N_2120);
and U2933 (N_2933,N_2186,N_2437);
nand U2934 (N_2934,N_2098,N_2062);
or U2935 (N_2935,N_2468,N_2168);
nand U2936 (N_2936,N_2339,N_2007);
nor U2937 (N_2937,N_2275,N_2414);
and U2938 (N_2938,N_2072,N_2280);
nand U2939 (N_2939,N_2487,N_2127);
and U2940 (N_2940,N_2192,N_2006);
xor U2941 (N_2941,N_2150,N_2408);
or U2942 (N_2942,N_2402,N_2407);
nor U2943 (N_2943,N_2366,N_2325);
nor U2944 (N_2944,N_2461,N_2181);
nand U2945 (N_2945,N_2223,N_2285);
or U2946 (N_2946,N_2206,N_2204);
nand U2947 (N_2947,N_2150,N_2024);
and U2948 (N_2948,N_2455,N_2283);
or U2949 (N_2949,N_2367,N_2223);
nor U2950 (N_2950,N_2037,N_2056);
or U2951 (N_2951,N_2191,N_2394);
or U2952 (N_2952,N_2240,N_2135);
nand U2953 (N_2953,N_2210,N_2040);
or U2954 (N_2954,N_2439,N_2481);
or U2955 (N_2955,N_2185,N_2339);
xor U2956 (N_2956,N_2365,N_2490);
nand U2957 (N_2957,N_2133,N_2223);
xnor U2958 (N_2958,N_2065,N_2022);
or U2959 (N_2959,N_2326,N_2332);
and U2960 (N_2960,N_2498,N_2347);
nand U2961 (N_2961,N_2343,N_2412);
nor U2962 (N_2962,N_2301,N_2063);
nand U2963 (N_2963,N_2467,N_2002);
xor U2964 (N_2964,N_2063,N_2056);
and U2965 (N_2965,N_2173,N_2336);
nor U2966 (N_2966,N_2400,N_2453);
and U2967 (N_2967,N_2440,N_2255);
and U2968 (N_2968,N_2045,N_2356);
xor U2969 (N_2969,N_2008,N_2021);
nor U2970 (N_2970,N_2140,N_2413);
nor U2971 (N_2971,N_2379,N_2276);
or U2972 (N_2972,N_2041,N_2249);
nand U2973 (N_2973,N_2199,N_2160);
and U2974 (N_2974,N_2413,N_2093);
nor U2975 (N_2975,N_2469,N_2027);
nor U2976 (N_2976,N_2038,N_2419);
or U2977 (N_2977,N_2408,N_2041);
xor U2978 (N_2978,N_2401,N_2498);
or U2979 (N_2979,N_2112,N_2062);
nand U2980 (N_2980,N_2200,N_2349);
xor U2981 (N_2981,N_2087,N_2462);
nand U2982 (N_2982,N_2018,N_2014);
or U2983 (N_2983,N_2372,N_2130);
nor U2984 (N_2984,N_2309,N_2097);
or U2985 (N_2985,N_2488,N_2065);
xnor U2986 (N_2986,N_2164,N_2386);
nor U2987 (N_2987,N_2279,N_2242);
or U2988 (N_2988,N_2000,N_2453);
nor U2989 (N_2989,N_2397,N_2492);
nand U2990 (N_2990,N_2226,N_2078);
xor U2991 (N_2991,N_2221,N_2334);
xnor U2992 (N_2992,N_2059,N_2262);
nand U2993 (N_2993,N_2218,N_2340);
nor U2994 (N_2994,N_2213,N_2301);
or U2995 (N_2995,N_2405,N_2162);
nand U2996 (N_2996,N_2022,N_2146);
xnor U2997 (N_2997,N_2083,N_2357);
and U2998 (N_2998,N_2474,N_2379);
and U2999 (N_2999,N_2009,N_2438);
or U3000 (N_3000,N_2835,N_2903);
or U3001 (N_3001,N_2536,N_2776);
xnor U3002 (N_3002,N_2565,N_2628);
nor U3003 (N_3003,N_2516,N_2504);
or U3004 (N_3004,N_2796,N_2638);
nor U3005 (N_3005,N_2674,N_2688);
nand U3006 (N_3006,N_2522,N_2625);
or U3007 (N_3007,N_2897,N_2898);
nor U3008 (N_3008,N_2510,N_2500);
nor U3009 (N_3009,N_2734,N_2823);
or U3010 (N_3010,N_2738,N_2816);
nand U3011 (N_3011,N_2704,N_2800);
nand U3012 (N_3012,N_2735,N_2590);
nor U3013 (N_3013,N_2801,N_2846);
or U3014 (N_3014,N_2677,N_2950);
nand U3015 (N_3015,N_2719,N_2843);
or U3016 (N_3016,N_2660,N_2792);
nor U3017 (N_3017,N_2953,N_2617);
xnor U3018 (N_3018,N_2965,N_2567);
xnor U3019 (N_3019,N_2794,N_2747);
xnor U3020 (N_3020,N_2515,N_2751);
or U3021 (N_3021,N_2624,N_2913);
xor U3022 (N_3022,N_2845,N_2940);
nor U3023 (N_3023,N_2725,N_2805);
nor U3024 (N_3024,N_2616,N_2929);
xnor U3025 (N_3025,N_2851,N_2618);
xnor U3026 (N_3026,N_2682,N_2525);
or U3027 (N_3027,N_2795,N_2773);
or U3028 (N_3028,N_2727,N_2692);
nor U3029 (N_3029,N_2887,N_2707);
nand U3030 (N_3030,N_2778,N_2882);
nor U3031 (N_3031,N_2596,N_2764);
or U3032 (N_3032,N_2875,N_2543);
nor U3033 (N_3033,N_2765,N_2948);
nand U3034 (N_3034,N_2675,N_2741);
nor U3035 (N_3035,N_2626,N_2972);
nand U3036 (N_3036,N_2827,N_2676);
nand U3037 (N_3037,N_2505,N_2553);
xnor U3038 (N_3038,N_2895,N_2663);
or U3039 (N_3039,N_2886,N_2756);
nand U3040 (N_3040,N_2894,N_2771);
and U3041 (N_3041,N_2755,N_2931);
and U3042 (N_3042,N_2668,N_2540);
xnor U3043 (N_3043,N_2981,N_2770);
or U3044 (N_3044,N_2813,N_2694);
nor U3045 (N_3045,N_2957,N_2870);
or U3046 (N_3046,N_2680,N_2621);
and U3047 (N_3047,N_2508,N_2554);
and U3048 (N_3048,N_2938,N_2612);
xor U3049 (N_3049,N_2592,N_2943);
nand U3050 (N_3050,N_2721,N_2996);
xnor U3051 (N_3051,N_2526,N_2927);
or U3052 (N_3052,N_2980,N_2605);
nor U3053 (N_3053,N_2817,N_2635);
or U3054 (N_3054,N_2549,N_2574);
or U3055 (N_3055,N_2569,N_2824);
and U3056 (N_3056,N_2865,N_2836);
nor U3057 (N_3057,N_2872,N_2761);
or U3058 (N_3058,N_2854,N_2924);
nand U3059 (N_3059,N_2608,N_2664);
nor U3060 (N_3060,N_2720,N_2842);
or U3061 (N_3061,N_2715,N_2766);
nand U3062 (N_3062,N_2534,N_2945);
nand U3063 (N_3063,N_2859,N_2669);
xor U3064 (N_3064,N_2809,N_2670);
xor U3065 (N_3065,N_2891,N_2806);
nand U3066 (N_3066,N_2511,N_2550);
nand U3067 (N_3067,N_2685,N_2821);
nand U3068 (N_3068,N_2702,N_2812);
nand U3069 (N_3069,N_2678,N_2822);
nand U3070 (N_3070,N_2873,N_2956);
nor U3071 (N_3071,N_2568,N_2671);
and U3072 (N_3072,N_2593,N_2701);
xnor U3073 (N_3073,N_2633,N_2620);
or U3074 (N_3074,N_2705,N_2629);
nand U3075 (N_3075,N_2687,N_2990);
or U3076 (N_3076,N_2867,N_2728);
xor U3077 (N_3077,N_2968,N_2757);
or U3078 (N_3078,N_2597,N_2934);
nor U3079 (N_3079,N_2700,N_2856);
xnor U3080 (N_3080,N_2802,N_2775);
nor U3081 (N_3081,N_2768,N_2863);
xor U3082 (N_3082,N_2529,N_2716);
nand U3083 (N_3083,N_2906,N_2706);
and U3084 (N_3084,N_2955,N_2695);
and U3085 (N_3085,N_2847,N_2651);
nand U3086 (N_3086,N_2967,N_2623);
nand U3087 (N_3087,N_2979,N_2935);
xnor U3088 (N_3088,N_2852,N_2922);
or U3089 (N_3089,N_2658,N_2912);
nor U3090 (N_3090,N_2781,N_2519);
and U3091 (N_3091,N_2864,N_2958);
xor U3092 (N_3092,N_2787,N_2793);
or U3093 (N_3093,N_2636,N_2960);
or U3094 (N_3094,N_2837,N_2502);
nand U3095 (N_3095,N_2532,N_2820);
nor U3096 (N_3096,N_2791,N_2901);
nor U3097 (N_3097,N_2542,N_2853);
nand U3098 (N_3098,N_2850,N_2782);
nor U3099 (N_3099,N_2807,N_2883);
or U3100 (N_3100,N_2578,N_2577);
or U3101 (N_3101,N_2932,N_2575);
and U3102 (N_3102,N_2690,N_2900);
nor U3103 (N_3103,N_2841,N_2866);
nand U3104 (N_3104,N_2926,N_2507);
or U3105 (N_3105,N_2609,N_2643);
or U3106 (N_3106,N_2644,N_2523);
xnor U3107 (N_3107,N_2966,N_2645);
and U3108 (N_3108,N_2995,N_2840);
nand U3109 (N_3109,N_2797,N_2533);
xor U3110 (N_3110,N_2518,N_2648);
or U3111 (N_3111,N_2888,N_2989);
xor U3112 (N_3112,N_2649,N_2632);
nand U3113 (N_3113,N_2910,N_2646);
and U3114 (N_3114,N_2889,N_2546);
and U3115 (N_3115,N_2760,N_2641);
or U3116 (N_3116,N_2524,N_2833);
nor U3117 (N_3117,N_2961,N_2581);
xnor U3118 (N_3118,N_2743,N_2509);
nor U3119 (N_3119,N_2538,N_2947);
nand U3120 (N_3120,N_2528,N_2637);
or U3121 (N_3121,N_2919,N_2893);
nand U3122 (N_3122,N_2928,N_2858);
nor U3123 (N_3123,N_2703,N_2642);
or U3124 (N_3124,N_2890,N_2537);
xor U3125 (N_3125,N_2871,N_2607);
or U3126 (N_3126,N_2750,N_2659);
and U3127 (N_3127,N_2964,N_2684);
xnor U3128 (N_3128,N_2804,N_2602);
nor U3129 (N_3129,N_2610,N_2829);
and U3130 (N_3130,N_2718,N_2923);
xor U3131 (N_3131,N_2552,N_2652);
nor U3132 (N_3132,N_2530,N_2949);
and U3133 (N_3133,N_2603,N_2733);
nand U3134 (N_3134,N_2595,N_2868);
nand U3135 (N_3135,N_2613,N_2724);
nand U3136 (N_3136,N_2885,N_2994);
nand U3137 (N_3137,N_2861,N_2634);
and U3138 (N_3138,N_2786,N_2539);
and U3139 (N_3139,N_2978,N_2899);
or U3140 (N_3140,N_2977,N_2656);
nor U3141 (N_3141,N_2828,N_2666);
or U3142 (N_3142,N_2580,N_2942);
or U3143 (N_3143,N_2679,N_2606);
xnor U3144 (N_3144,N_2937,N_2586);
or U3145 (N_3145,N_2521,N_2892);
nor U3146 (N_3146,N_2591,N_2561);
xor U3147 (N_3147,N_2564,N_2814);
xor U3148 (N_3148,N_2650,N_2832);
or U3149 (N_3149,N_2573,N_2544);
xnor U3150 (N_3150,N_2681,N_2905);
xnor U3151 (N_3151,N_2551,N_2514);
and U3152 (N_3152,N_2627,N_2789);
and U3153 (N_3153,N_2512,N_2848);
nor U3154 (N_3154,N_2811,N_2788);
xor U3155 (N_3155,N_2693,N_2944);
or U3156 (N_3156,N_2691,N_2984);
and U3157 (N_3157,N_2963,N_2876);
xnor U3158 (N_3158,N_2982,N_2556);
nor U3159 (N_3159,N_2983,N_2619);
or U3160 (N_3160,N_2601,N_2976);
xnor U3161 (N_3161,N_2520,N_2737);
nand U3162 (N_3162,N_2558,N_2709);
xnor U3163 (N_3163,N_2729,N_2630);
xnor U3164 (N_3164,N_2672,N_2600);
and U3165 (N_3165,N_2908,N_2742);
nand U3166 (N_3166,N_2710,N_2951);
and U3167 (N_3167,N_2917,N_2884);
nand U3168 (N_3168,N_2952,N_2655);
nor U3169 (N_3169,N_2783,N_2946);
or U3170 (N_3170,N_2686,N_2611);
and U3171 (N_3171,N_2974,N_2914);
or U3172 (N_3172,N_2583,N_2902);
or U3173 (N_3173,N_2639,N_2810);
xor U3174 (N_3174,N_2711,N_2826);
and U3175 (N_3175,N_2769,N_2631);
or U3176 (N_3176,N_2745,N_2818);
nand U3177 (N_3177,N_2665,N_2844);
and U3178 (N_3178,N_2896,N_2973);
nor U3179 (N_3179,N_2535,N_2683);
xor U3180 (N_3180,N_2599,N_2654);
or U3181 (N_3181,N_2723,N_2936);
nor U3182 (N_3182,N_2501,N_2772);
nor U3183 (N_3183,N_2999,N_2998);
nor U3184 (N_3184,N_2991,N_2547);
and U3185 (N_3185,N_2941,N_2753);
nor U3186 (N_3186,N_2736,N_2920);
nor U3187 (N_3187,N_2988,N_2767);
and U3188 (N_3188,N_2808,N_2878);
xor U3189 (N_3189,N_2752,N_2732);
xnor U3190 (N_3190,N_2740,N_2986);
xnor U3191 (N_3191,N_2784,N_2830);
nand U3192 (N_3192,N_2662,N_2722);
or U3193 (N_3193,N_2915,N_2777);
xnor U3194 (N_3194,N_2557,N_2726);
or U3195 (N_3195,N_2527,N_2708);
nand U3196 (N_3196,N_2874,N_2667);
nand U3197 (N_3197,N_2962,N_2657);
and U3198 (N_3198,N_2993,N_2661);
and U3199 (N_3199,N_2798,N_2614);
nand U3200 (N_3200,N_2831,N_2975);
or U3201 (N_3201,N_2696,N_2780);
and U3202 (N_3202,N_2647,N_2563);
xor U3203 (N_3203,N_2779,N_2925);
or U3204 (N_3204,N_2731,N_2748);
and U3205 (N_3205,N_2572,N_2839);
xor U3206 (N_3206,N_2604,N_2589);
nor U3207 (N_3207,N_2598,N_2918);
and U3208 (N_3208,N_2689,N_2517);
nor U3209 (N_3209,N_2699,N_2548);
and U3210 (N_3210,N_2559,N_2673);
nand U3211 (N_3211,N_2959,N_2774);
and U3212 (N_3212,N_2754,N_2555);
nand U3213 (N_3213,N_2579,N_2911);
nand U3214 (N_3214,N_2571,N_2758);
xnor U3215 (N_3215,N_2566,N_2933);
xnor U3216 (N_3216,N_2615,N_2746);
xnor U3217 (N_3217,N_2877,N_2594);
and U3218 (N_3218,N_2562,N_2970);
nor U3219 (N_3219,N_2907,N_2869);
or U3220 (N_3220,N_2803,N_2541);
or U3221 (N_3221,N_2576,N_2939);
nand U3222 (N_3222,N_2785,N_2640);
and U3223 (N_3223,N_2744,N_2712);
nand U3224 (N_3224,N_2992,N_2584);
and U3225 (N_3225,N_2531,N_2730);
nor U3226 (N_3226,N_2713,N_2997);
xor U3227 (N_3227,N_2799,N_2763);
or U3228 (N_3228,N_2857,N_2985);
and U3229 (N_3229,N_2653,N_2971);
nand U3230 (N_3230,N_2585,N_2909);
or U3231 (N_3231,N_2739,N_2860);
nand U3232 (N_3232,N_2503,N_2513);
nand U3233 (N_3233,N_2880,N_2825);
nor U3234 (N_3234,N_2717,N_2790);
nor U3235 (N_3235,N_2904,N_2987);
and U3236 (N_3236,N_2749,N_2815);
or U3237 (N_3237,N_2714,N_2879);
nand U3238 (N_3238,N_2570,N_2698);
xor U3239 (N_3239,N_2969,N_2881);
xnor U3240 (N_3240,N_2697,N_2849);
nand U3241 (N_3241,N_2862,N_2930);
nor U3242 (N_3242,N_2759,N_2545);
nor U3243 (N_3243,N_2622,N_2916);
xnor U3244 (N_3244,N_2954,N_2582);
nor U3245 (N_3245,N_2588,N_2560);
and U3246 (N_3246,N_2762,N_2819);
or U3247 (N_3247,N_2506,N_2587);
or U3248 (N_3248,N_2921,N_2855);
or U3249 (N_3249,N_2838,N_2834);
nor U3250 (N_3250,N_2516,N_2827);
nor U3251 (N_3251,N_2930,N_2814);
and U3252 (N_3252,N_2858,N_2519);
and U3253 (N_3253,N_2676,N_2843);
xnor U3254 (N_3254,N_2573,N_2769);
or U3255 (N_3255,N_2751,N_2872);
and U3256 (N_3256,N_2926,N_2975);
nor U3257 (N_3257,N_2879,N_2905);
nor U3258 (N_3258,N_2810,N_2856);
nand U3259 (N_3259,N_2537,N_2996);
and U3260 (N_3260,N_2626,N_2606);
nor U3261 (N_3261,N_2882,N_2506);
and U3262 (N_3262,N_2744,N_2573);
nand U3263 (N_3263,N_2650,N_2777);
nor U3264 (N_3264,N_2886,N_2520);
xor U3265 (N_3265,N_2683,N_2694);
or U3266 (N_3266,N_2994,N_2586);
xor U3267 (N_3267,N_2760,N_2532);
or U3268 (N_3268,N_2810,N_2748);
nand U3269 (N_3269,N_2587,N_2709);
nor U3270 (N_3270,N_2986,N_2659);
nand U3271 (N_3271,N_2993,N_2503);
and U3272 (N_3272,N_2780,N_2883);
nor U3273 (N_3273,N_2564,N_2950);
or U3274 (N_3274,N_2626,N_2962);
and U3275 (N_3275,N_2563,N_2806);
nand U3276 (N_3276,N_2595,N_2729);
nand U3277 (N_3277,N_2539,N_2626);
nand U3278 (N_3278,N_2717,N_2512);
xor U3279 (N_3279,N_2599,N_2724);
and U3280 (N_3280,N_2960,N_2821);
or U3281 (N_3281,N_2941,N_2599);
xnor U3282 (N_3282,N_2845,N_2584);
nor U3283 (N_3283,N_2539,N_2817);
and U3284 (N_3284,N_2719,N_2753);
or U3285 (N_3285,N_2739,N_2746);
nand U3286 (N_3286,N_2560,N_2661);
and U3287 (N_3287,N_2892,N_2962);
nor U3288 (N_3288,N_2641,N_2813);
xor U3289 (N_3289,N_2834,N_2540);
and U3290 (N_3290,N_2951,N_2738);
nor U3291 (N_3291,N_2671,N_2505);
nand U3292 (N_3292,N_2524,N_2766);
nand U3293 (N_3293,N_2658,N_2793);
nor U3294 (N_3294,N_2602,N_2862);
xor U3295 (N_3295,N_2650,N_2748);
nand U3296 (N_3296,N_2528,N_2511);
nor U3297 (N_3297,N_2647,N_2622);
xnor U3298 (N_3298,N_2874,N_2643);
nand U3299 (N_3299,N_2982,N_2686);
or U3300 (N_3300,N_2928,N_2503);
xor U3301 (N_3301,N_2734,N_2672);
nor U3302 (N_3302,N_2600,N_2793);
nand U3303 (N_3303,N_2899,N_2773);
nor U3304 (N_3304,N_2621,N_2713);
nor U3305 (N_3305,N_2610,N_2521);
and U3306 (N_3306,N_2892,N_2690);
or U3307 (N_3307,N_2761,N_2504);
or U3308 (N_3308,N_2998,N_2552);
nand U3309 (N_3309,N_2839,N_2774);
nor U3310 (N_3310,N_2806,N_2716);
nor U3311 (N_3311,N_2970,N_2688);
and U3312 (N_3312,N_2824,N_2768);
or U3313 (N_3313,N_2721,N_2745);
or U3314 (N_3314,N_2603,N_2588);
or U3315 (N_3315,N_2847,N_2953);
xnor U3316 (N_3316,N_2693,N_2534);
nand U3317 (N_3317,N_2906,N_2646);
xnor U3318 (N_3318,N_2685,N_2765);
and U3319 (N_3319,N_2553,N_2541);
and U3320 (N_3320,N_2543,N_2855);
nor U3321 (N_3321,N_2791,N_2699);
or U3322 (N_3322,N_2623,N_2591);
nor U3323 (N_3323,N_2933,N_2661);
nor U3324 (N_3324,N_2732,N_2600);
or U3325 (N_3325,N_2578,N_2524);
xnor U3326 (N_3326,N_2750,N_2787);
nand U3327 (N_3327,N_2820,N_2645);
nand U3328 (N_3328,N_2857,N_2987);
nand U3329 (N_3329,N_2681,N_2944);
nor U3330 (N_3330,N_2633,N_2594);
xor U3331 (N_3331,N_2563,N_2777);
and U3332 (N_3332,N_2625,N_2568);
xnor U3333 (N_3333,N_2671,N_2976);
xnor U3334 (N_3334,N_2865,N_2950);
xnor U3335 (N_3335,N_2907,N_2826);
xor U3336 (N_3336,N_2794,N_2714);
nor U3337 (N_3337,N_2764,N_2658);
xor U3338 (N_3338,N_2553,N_2539);
nand U3339 (N_3339,N_2895,N_2744);
nand U3340 (N_3340,N_2641,N_2979);
xor U3341 (N_3341,N_2861,N_2857);
nor U3342 (N_3342,N_2667,N_2839);
or U3343 (N_3343,N_2578,N_2571);
nand U3344 (N_3344,N_2863,N_2874);
nand U3345 (N_3345,N_2753,N_2939);
nor U3346 (N_3346,N_2988,N_2968);
and U3347 (N_3347,N_2918,N_2927);
and U3348 (N_3348,N_2511,N_2527);
and U3349 (N_3349,N_2610,N_2868);
and U3350 (N_3350,N_2589,N_2913);
nor U3351 (N_3351,N_2803,N_2577);
and U3352 (N_3352,N_2831,N_2702);
or U3353 (N_3353,N_2662,N_2838);
xor U3354 (N_3354,N_2614,N_2605);
xnor U3355 (N_3355,N_2940,N_2680);
xnor U3356 (N_3356,N_2756,N_2738);
xnor U3357 (N_3357,N_2959,N_2692);
or U3358 (N_3358,N_2954,N_2766);
and U3359 (N_3359,N_2832,N_2889);
nand U3360 (N_3360,N_2523,N_2692);
xor U3361 (N_3361,N_2728,N_2611);
nand U3362 (N_3362,N_2522,N_2955);
and U3363 (N_3363,N_2861,N_2557);
and U3364 (N_3364,N_2642,N_2958);
or U3365 (N_3365,N_2608,N_2707);
nand U3366 (N_3366,N_2554,N_2818);
and U3367 (N_3367,N_2736,N_2899);
nand U3368 (N_3368,N_2571,N_2825);
or U3369 (N_3369,N_2630,N_2880);
xnor U3370 (N_3370,N_2855,N_2523);
and U3371 (N_3371,N_2504,N_2548);
nand U3372 (N_3372,N_2801,N_2872);
and U3373 (N_3373,N_2845,N_2999);
or U3374 (N_3374,N_2979,N_2656);
and U3375 (N_3375,N_2879,N_2881);
nor U3376 (N_3376,N_2794,N_2912);
nor U3377 (N_3377,N_2758,N_2556);
or U3378 (N_3378,N_2907,N_2573);
and U3379 (N_3379,N_2862,N_2754);
nor U3380 (N_3380,N_2941,N_2701);
and U3381 (N_3381,N_2796,N_2591);
and U3382 (N_3382,N_2945,N_2503);
nand U3383 (N_3383,N_2932,N_2691);
and U3384 (N_3384,N_2842,N_2816);
nor U3385 (N_3385,N_2752,N_2959);
and U3386 (N_3386,N_2732,N_2581);
and U3387 (N_3387,N_2733,N_2562);
nor U3388 (N_3388,N_2897,N_2730);
or U3389 (N_3389,N_2552,N_2550);
nand U3390 (N_3390,N_2751,N_2693);
and U3391 (N_3391,N_2555,N_2891);
and U3392 (N_3392,N_2616,N_2773);
or U3393 (N_3393,N_2816,N_2967);
or U3394 (N_3394,N_2634,N_2588);
and U3395 (N_3395,N_2899,N_2961);
nor U3396 (N_3396,N_2895,N_2816);
or U3397 (N_3397,N_2838,N_2591);
nor U3398 (N_3398,N_2896,N_2854);
and U3399 (N_3399,N_2593,N_2549);
nor U3400 (N_3400,N_2612,N_2773);
nor U3401 (N_3401,N_2930,N_2538);
nand U3402 (N_3402,N_2880,N_2990);
or U3403 (N_3403,N_2803,N_2944);
and U3404 (N_3404,N_2639,N_2985);
and U3405 (N_3405,N_2599,N_2986);
or U3406 (N_3406,N_2729,N_2817);
and U3407 (N_3407,N_2518,N_2537);
nand U3408 (N_3408,N_2929,N_2505);
and U3409 (N_3409,N_2964,N_2976);
nor U3410 (N_3410,N_2701,N_2778);
or U3411 (N_3411,N_2517,N_2626);
nand U3412 (N_3412,N_2763,N_2830);
nand U3413 (N_3413,N_2981,N_2844);
or U3414 (N_3414,N_2710,N_2818);
xor U3415 (N_3415,N_2720,N_2654);
and U3416 (N_3416,N_2666,N_2673);
or U3417 (N_3417,N_2985,N_2589);
xnor U3418 (N_3418,N_2745,N_2664);
nor U3419 (N_3419,N_2549,N_2960);
or U3420 (N_3420,N_2750,N_2732);
and U3421 (N_3421,N_2885,N_2814);
xor U3422 (N_3422,N_2864,N_2603);
and U3423 (N_3423,N_2601,N_2967);
and U3424 (N_3424,N_2823,N_2513);
or U3425 (N_3425,N_2794,N_2973);
or U3426 (N_3426,N_2547,N_2981);
nand U3427 (N_3427,N_2820,N_2979);
and U3428 (N_3428,N_2615,N_2856);
and U3429 (N_3429,N_2694,N_2888);
nor U3430 (N_3430,N_2732,N_2998);
nand U3431 (N_3431,N_2887,N_2556);
nand U3432 (N_3432,N_2651,N_2805);
and U3433 (N_3433,N_2881,N_2532);
nor U3434 (N_3434,N_2804,N_2803);
xor U3435 (N_3435,N_2853,N_2558);
nor U3436 (N_3436,N_2699,N_2769);
and U3437 (N_3437,N_2579,N_2750);
and U3438 (N_3438,N_2580,N_2683);
xor U3439 (N_3439,N_2900,N_2813);
nand U3440 (N_3440,N_2778,N_2876);
nor U3441 (N_3441,N_2956,N_2538);
nor U3442 (N_3442,N_2923,N_2688);
nand U3443 (N_3443,N_2620,N_2565);
nor U3444 (N_3444,N_2823,N_2860);
nand U3445 (N_3445,N_2974,N_2584);
xnor U3446 (N_3446,N_2890,N_2952);
xor U3447 (N_3447,N_2830,N_2658);
or U3448 (N_3448,N_2765,N_2989);
nand U3449 (N_3449,N_2846,N_2835);
xor U3450 (N_3450,N_2880,N_2923);
or U3451 (N_3451,N_2649,N_2761);
or U3452 (N_3452,N_2858,N_2923);
and U3453 (N_3453,N_2633,N_2593);
xnor U3454 (N_3454,N_2782,N_2858);
xnor U3455 (N_3455,N_2796,N_2585);
nand U3456 (N_3456,N_2989,N_2728);
nor U3457 (N_3457,N_2800,N_2506);
nor U3458 (N_3458,N_2993,N_2855);
xor U3459 (N_3459,N_2694,N_2746);
or U3460 (N_3460,N_2731,N_2746);
xor U3461 (N_3461,N_2534,N_2674);
xor U3462 (N_3462,N_2775,N_2785);
or U3463 (N_3463,N_2998,N_2723);
nor U3464 (N_3464,N_2740,N_2829);
and U3465 (N_3465,N_2711,N_2872);
nand U3466 (N_3466,N_2984,N_2976);
and U3467 (N_3467,N_2960,N_2760);
and U3468 (N_3468,N_2747,N_2873);
and U3469 (N_3469,N_2774,N_2513);
xnor U3470 (N_3470,N_2907,N_2821);
and U3471 (N_3471,N_2900,N_2720);
or U3472 (N_3472,N_2884,N_2531);
nor U3473 (N_3473,N_2507,N_2646);
and U3474 (N_3474,N_2829,N_2581);
nor U3475 (N_3475,N_2661,N_2746);
xor U3476 (N_3476,N_2928,N_2622);
or U3477 (N_3477,N_2759,N_2707);
or U3478 (N_3478,N_2500,N_2942);
xnor U3479 (N_3479,N_2813,N_2658);
nor U3480 (N_3480,N_2811,N_2727);
or U3481 (N_3481,N_2704,N_2531);
or U3482 (N_3482,N_2737,N_2718);
and U3483 (N_3483,N_2994,N_2546);
or U3484 (N_3484,N_2924,N_2719);
and U3485 (N_3485,N_2694,N_2744);
xor U3486 (N_3486,N_2810,N_2894);
xnor U3487 (N_3487,N_2830,N_2554);
or U3488 (N_3488,N_2761,N_2601);
or U3489 (N_3489,N_2619,N_2572);
nand U3490 (N_3490,N_2685,N_2620);
nor U3491 (N_3491,N_2632,N_2972);
nand U3492 (N_3492,N_2886,N_2730);
and U3493 (N_3493,N_2977,N_2703);
nand U3494 (N_3494,N_2561,N_2553);
or U3495 (N_3495,N_2577,N_2500);
nor U3496 (N_3496,N_2970,N_2547);
and U3497 (N_3497,N_2819,N_2590);
or U3498 (N_3498,N_2523,N_2731);
xnor U3499 (N_3499,N_2890,N_2981);
nand U3500 (N_3500,N_3044,N_3252);
and U3501 (N_3501,N_3060,N_3399);
nor U3502 (N_3502,N_3131,N_3178);
and U3503 (N_3503,N_3404,N_3299);
or U3504 (N_3504,N_3211,N_3014);
or U3505 (N_3505,N_3141,N_3076);
nand U3506 (N_3506,N_3132,N_3296);
or U3507 (N_3507,N_3104,N_3357);
or U3508 (N_3508,N_3054,N_3109);
nand U3509 (N_3509,N_3158,N_3200);
nand U3510 (N_3510,N_3469,N_3359);
nand U3511 (N_3511,N_3069,N_3019);
or U3512 (N_3512,N_3315,N_3038);
or U3513 (N_3513,N_3456,N_3274);
and U3514 (N_3514,N_3080,N_3460);
xnor U3515 (N_3515,N_3089,N_3325);
and U3516 (N_3516,N_3249,N_3198);
xor U3517 (N_3517,N_3427,N_3475);
or U3518 (N_3518,N_3018,N_3229);
nor U3519 (N_3519,N_3270,N_3128);
nor U3520 (N_3520,N_3424,N_3217);
and U3521 (N_3521,N_3147,N_3232);
xor U3522 (N_3522,N_3119,N_3191);
xor U3523 (N_3523,N_3115,N_3334);
or U3524 (N_3524,N_3219,N_3015);
xor U3525 (N_3525,N_3367,N_3140);
or U3526 (N_3526,N_3477,N_3250);
and U3527 (N_3527,N_3073,N_3055);
nand U3528 (N_3528,N_3068,N_3067);
nand U3529 (N_3529,N_3478,N_3387);
nand U3530 (N_3530,N_3336,N_3177);
and U3531 (N_3531,N_3319,N_3451);
nand U3532 (N_3532,N_3352,N_3483);
or U3533 (N_3533,N_3335,N_3444);
xnor U3534 (N_3534,N_3281,N_3340);
or U3535 (N_3535,N_3300,N_3123);
and U3536 (N_3536,N_3492,N_3025);
nand U3537 (N_3537,N_3101,N_3129);
xor U3538 (N_3538,N_3280,N_3084);
xnor U3539 (N_3539,N_3182,N_3405);
and U3540 (N_3540,N_3351,N_3180);
or U3541 (N_3541,N_3066,N_3439);
and U3542 (N_3542,N_3017,N_3188);
nor U3543 (N_3543,N_3380,N_3390);
xor U3544 (N_3544,N_3048,N_3433);
and U3545 (N_3545,N_3116,N_3401);
xor U3546 (N_3546,N_3309,N_3453);
xor U3547 (N_3547,N_3423,N_3096);
xnor U3548 (N_3548,N_3005,N_3108);
nand U3549 (N_3549,N_3485,N_3279);
and U3550 (N_3550,N_3022,N_3432);
nor U3551 (N_3551,N_3410,N_3434);
or U3552 (N_3552,N_3041,N_3481);
nand U3553 (N_3553,N_3001,N_3402);
and U3554 (N_3554,N_3320,N_3409);
or U3555 (N_3555,N_3127,N_3455);
nand U3556 (N_3556,N_3465,N_3070);
xor U3557 (N_3557,N_3006,N_3457);
nor U3558 (N_3558,N_3375,N_3161);
xor U3559 (N_3559,N_3329,N_3298);
and U3560 (N_3560,N_3491,N_3083);
xnor U3561 (N_3561,N_3011,N_3356);
nor U3562 (N_3562,N_3471,N_3310);
nand U3563 (N_3563,N_3165,N_3151);
xor U3564 (N_3564,N_3149,N_3239);
nor U3565 (N_3565,N_3228,N_3024);
nor U3566 (N_3566,N_3266,N_3092);
nor U3567 (N_3567,N_3134,N_3138);
and U3568 (N_3568,N_3071,N_3064);
xor U3569 (N_3569,N_3350,N_3111);
and U3570 (N_3570,N_3220,N_3153);
or U3571 (N_3571,N_3400,N_3181);
nand U3572 (N_3572,N_3487,N_3323);
nand U3573 (N_3573,N_3259,N_3088);
or U3574 (N_3574,N_3332,N_3347);
and U3575 (N_3575,N_3371,N_3376);
nand U3576 (N_3576,N_3470,N_3099);
or U3577 (N_3577,N_3366,N_3360);
nor U3578 (N_3578,N_3205,N_3124);
or U3579 (N_3579,N_3030,N_3263);
and U3580 (N_3580,N_3321,N_3476);
and U3581 (N_3581,N_3372,N_3035);
nor U3582 (N_3582,N_3341,N_3303);
xor U3583 (N_3583,N_3098,N_3474);
xor U3584 (N_3584,N_3349,N_3408);
or U3585 (N_3585,N_3373,N_3110);
nor U3586 (N_3586,N_3130,N_3114);
nand U3587 (N_3587,N_3365,N_3020);
xnor U3588 (N_3588,N_3311,N_3327);
nor U3589 (N_3589,N_3265,N_3497);
nand U3590 (N_3590,N_3216,N_3369);
nor U3591 (N_3591,N_3186,N_3425);
or U3592 (N_3592,N_3192,N_3053);
nand U3593 (N_3593,N_3324,N_3489);
nor U3594 (N_3594,N_3395,N_3148);
and U3595 (N_3595,N_3461,N_3183);
nand U3596 (N_3596,N_3193,N_3154);
nand U3597 (N_3597,N_3046,N_3251);
nand U3598 (N_3598,N_3295,N_3312);
and U3599 (N_3599,N_3185,N_3137);
xnor U3600 (N_3600,N_3440,N_3330);
nor U3601 (N_3601,N_3314,N_3464);
nor U3602 (N_3602,N_3164,N_3264);
xnor U3603 (N_3603,N_3415,N_3466);
nor U3604 (N_3604,N_3026,N_3291);
or U3605 (N_3605,N_3246,N_3145);
nor U3606 (N_3606,N_3081,N_3037);
nor U3607 (N_3607,N_3087,N_3482);
or U3608 (N_3608,N_3036,N_3418);
nand U3609 (N_3609,N_3438,N_3258);
nor U3610 (N_3610,N_3117,N_3097);
or U3611 (N_3611,N_3480,N_3225);
xor U3612 (N_3612,N_3388,N_3441);
or U3613 (N_3613,N_3284,N_3195);
nor U3614 (N_3614,N_3428,N_3121);
and U3615 (N_3615,N_3029,N_3215);
or U3616 (N_3616,N_3223,N_3093);
nor U3617 (N_3617,N_3361,N_3374);
nor U3618 (N_3618,N_3275,N_3496);
and U3619 (N_3619,N_3162,N_3050);
xor U3620 (N_3620,N_3452,N_3257);
nand U3621 (N_3621,N_3398,N_3004);
nand U3622 (N_3622,N_3412,N_3448);
nand U3623 (N_3623,N_3176,N_3458);
nand U3624 (N_3624,N_3394,N_3459);
and U3625 (N_3625,N_3112,N_3430);
xor U3626 (N_3626,N_3422,N_3316);
or U3627 (N_3627,N_3245,N_3077);
and U3628 (N_3628,N_3328,N_3339);
and U3629 (N_3629,N_3146,N_3007);
xor U3630 (N_3630,N_3021,N_3343);
nor U3631 (N_3631,N_3243,N_3344);
nand U3632 (N_3632,N_3079,N_3454);
xnor U3633 (N_3633,N_3345,N_3212);
or U3634 (N_3634,N_3013,N_3468);
xor U3635 (N_3635,N_3317,N_3268);
and U3636 (N_3636,N_3382,N_3133);
xor U3637 (N_3637,N_3113,N_3307);
nor U3638 (N_3638,N_3260,N_3143);
nand U3639 (N_3639,N_3306,N_3012);
and U3640 (N_3640,N_3269,N_3169);
nor U3641 (N_3641,N_3144,N_3156);
and U3642 (N_3642,N_3033,N_3179);
nor U3643 (N_3643,N_3290,N_3059);
and U3644 (N_3644,N_3392,N_3479);
and U3645 (N_3645,N_3166,N_3125);
or U3646 (N_3646,N_3287,N_3009);
nor U3647 (N_3647,N_3197,N_3493);
or U3648 (N_3648,N_3381,N_3342);
or U3649 (N_3649,N_3234,N_3027);
xnor U3650 (N_3650,N_3206,N_3285);
nor U3651 (N_3651,N_3233,N_3413);
nor U3652 (N_3652,N_3237,N_3032);
and U3653 (N_3653,N_3331,N_3364);
and U3654 (N_3654,N_3196,N_3039);
nand U3655 (N_3655,N_3391,N_3043);
nand U3656 (N_3656,N_3254,N_3122);
nor U3657 (N_3657,N_3277,N_3201);
and U3658 (N_3658,N_3222,N_3155);
xnor U3659 (N_3659,N_3486,N_3389);
nand U3660 (N_3660,N_3411,N_3484);
nand U3661 (N_3661,N_3106,N_3184);
and U3662 (N_3662,N_3318,N_3028);
and U3663 (N_3663,N_3003,N_3214);
or U3664 (N_3664,N_3213,N_3247);
and U3665 (N_3665,N_3354,N_3337);
xor U3666 (N_3666,N_3058,N_3086);
nand U3667 (N_3667,N_3355,N_3172);
nand U3668 (N_3668,N_3305,N_3000);
or U3669 (N_3669,N_3126,N_3010);
nor U3670 (N_3670,N_3174,N_3283);
nand U3671 (N_3671,N_3338,N_3209);
nor U3672 (N_3672,N_3218,N_3304);
xor U3673 (N_3673,N_3091,N_3383);
or U3674 (N_3674,N_3210,N_3498);
nand U3675 (N_3675,N_3288,N_3107);
or U3676 (N_3676,N_3173,N_3346);
nor U3677 (N_3677,N_3231,N_3139);
nand U3678 (N_3678,N_3135,N_3202);
xnor U3679 (N_3679,N_3008,N_3170);
xor U3680 (N_3680,N_3204,N_3241);
and U3681 (N_3681,N_3421,N_3253);
nand U3682 (N_3682,N_3462,N_3157);
and U3683 (N_3683,N_3378,N_3272);
nor U3684 (N_3684,N_3194,N_3152);
or U3685 (N_3685,N_3235,N_3322);
nand U3686 (N_3686,N_3159,N_3207);
and U3687 (N_3687,N_3100,N_3403);
or U3688 (N_3688,N_3150,N_3463);
nor U3689 (N_3689,N_3102,N_3442);
and U3690 (N_3690,N_3445,N_3057);
or U3691 (N_3691,N_3160,N_3436);
xnor U3692 (N_3692,N_3446,N_3226);
or U3693 (N_3693,N_3377,N_3203);
or U3694 (N_3694,N_3042,N_3082);
nand U3695 (N_3695,N_3384,N_3419);
nor U3696 (N_3696,N_3063,N_3045);
and U3697 (N_3697,N_3199,N_3326);
xnor U3698 (N_3698,N_3467,N_3016);
nor U3699 (N_3699,N_3171,N_3267);
nor U3700 (N_3700,N_3308,N_3348);
nand U3701 (N_3701,N_3406,N_3051);
or U3702 (N_3702,N_3292,N_3034);
or U3703 (N_3703,N_3435,N_3065);
xor U3704 (N_3704,N_3286,N_3368);
nor U3705 (N_3705,N_3227,N_3293);
nor U3706 (N_3706,N_3447,N_3420);
xor U3707 (N_3707,N_3333,N_3449);
and U3708 (N_3708,N_3118,N_3120);
nor U3709 (N_3709,N_3370,N_3056);
nand U3710 (N_3710,N_3386,N_3393);
or U3711 (N_3711,N_3238,N_3499);
xnor U3712 (N_3712,N_3495,N_3078);
xnor U3713 (N_3713,N_3002,N_3095);
nor U3714 (N_3714,N_3472,N_3136);
or U3715 (N_3715,N_3090,N_3248);
and U3716 (N_3716,N_3049,N_3074);
and U3717 (N_3717,N_3443,N_3494);
nand U3718 (N_3718,N_3208,N_3450);
and U3719 (N_3719,N_3061,N_3175);
nor U3720 (N_3720,N_3103,N_3397);
or U3721 (N_3721,N_3072,N_3302);
or U3722 (N_3722,N_3221,N_3473);
nor U3723 (N_3723,N_3353,N_3282);
xor U3724 (N_3724,N_3261,N_3262);
or U3725 (N_3725,N_3236,N_3429);
and U3726 (N_3726,N_3240,N_3244);
nand U3727 (N_3727,N_3488,N_3490);
or U3728 (N_3728,N_3075,N_3407);
xnor U3729 (N_3729,N_3437,N_3385);
xor U3730 (N_3730,N_3190,N_3230);
xnor U3731 (N_3731,N_3363,N_3416);
nand U3732 (N_3732,N_3168,N_3167);
and U3733 (N_3733,N_3294,N_3426);
or U3734 (N_3734,N_3062,N_3040);
or U3735 (N_3735,N_3414,N_3031);
nor U3736 (N_3736,N_3278,N_3189);
or U3737 (N_3737,N_3273,N_3224);
nor U3738 (N_3738,N_3094,N_3142);
nor U3739 (N_3739,N_3396,N_3271);
nand U3740 (N_3740,N_3085,N_3297);
and U3741 (N_3741,N_3431,N_3187);
or U3742 (N_3742,N_3289,N_3023);
or U3743 (N_3743,N_3163,N_3417);
or U3744 (N_3744,N_3256,N_3362);
nor U3745 (N_3745,N_3276,N_3105);
nand U3746 (N_3746,N_3047,N_3313);
xor U3747 (N_3747,N_3242,N_3052);
or U3748 (N_3748,N_3358,N_3379);
nor U3749 (N_3749,N_3255,N_3301);
nand U3750 (N_3750,N_3278,N_3323);
xnor U3751 (N_3751,N_3233,N_3146);
nor U3752 (N_3752,N_3211,N_3261);
nand U3753 (N_3753,N_3112,N_3156);
nor U3754 (N_3754,N_3365,N_3239);
nor U3755 (N_3755,N_3421,N_3149);
xnor U3756 (N_3756,N_3449,N_3385);
nand U3757 (N_3757,N_3405,N_3122);
or U3758 (N_3758,N_3278,N_3328);
or U3759 (N_3759,N_3036,N_3365);
nand U3760 (N_3760,N_3077,N_3494);
nor U3761 (N_3761,N_3355,N_3100);
nand U3762 (N_3762,N_3213,N_3122);
xnor U3763 (N_3763,N_3479,N_3072);
or U3764 (N_3764,N_3187,N_3299);
and U3765 (N_3765,N_3160,N_3291);
or U3766 (N_3766,N_3033,N_3230);
nand U3767 (N_3767,N_3152,N_3150);
nand U3768 (N_3768,N_3420,N_3272);
xnor U3769 (N_3769,N_3030,N_3335);
and U3770 (N_3770,N_3205,N_3384);
nor U3771 (N_3771,N_3031,N_3497);
nand U3772 (N_3772,N_3441,N_3213);
and U3773 (N_3773,N_3452,N_3198);
and U3774 (N_3774,N_3134,N_3072);
nor U3775 (N_3775,N_3210,N_3127);
nand U3776 (N_3776,N_3311,N_3430);
nor U3777 (N_3777,N_3326,N_3047);
or U3778 (N_3778,N_3040,N_3164);
xor U3779 (N_3779,N_3340,N_3187);
or U3780 (N_3780,N_3210,N_3041);
and U3781 (N_3781,N_3281,N_3006);
nor U3782 (N_3782,N_3070,N_3230);
nor U3783 (N_3783,N_3327,N_3472);
and U3784 (N_3784,N_3156,N_3423);
or U3785 (N_3785,N_3492,N_3411);
and U3786 (N_3786,N_3069,N_3195);
nand U3787 (N_3787,N_3443,N_3187);
nor U3788 (N_3788,N_3340,N_3133);
and U3789 (N_3789,N_3375,N_3483);
xnor U3790 (N_3790,N_3284,N_3136);
and U3791 (N_3791,N_3215,N_3448);
nand U3792 (N_3792,N_3374,N_3084);
and U3793 (N_3793,N_3048,N_3348);
nand U3794 (N_3794,N_3044,N_3063);
or U3795 (N_3795,N_3457,N_3078);
nand U3796 (N_3796,N_3140,N_3189);
and U3797 (N_3797,N_3424,N_3195);
nand U3798 (N_3798,N_3295,N_3376);
and U3799 (N_3799,N_3414,N_3183);
and U3800 (N_3800,N_3099,N_3111);
nor U3801 (N_3801,N_3094,N_3202);
xnor U3802 (N_3802,N_3310,N_3332);
nand U3803 (N_3803,N_3251,N_3497);
nor U3804 (N_3804,N_3003,N_3151);
and U3805 (N_3805,N_3065,N_3177);
nor U3806 (N_3806,N_3480,N_3164);
xor U3807 (N_3807,N_3240,N_3140);
and U3808 (N_3808,N_3328,N_3077);
and U3809 (N_3809,N_3383,N_3271);
nand U3810 (N_3810,N_3210,N_3155);
nand U3811 (N_3811,N_3008,N_3102);
xnor U3812 (N_3812,N_3437,N_3472);
xnor U3813 (N_3813,N_3096,N_3115);
or U3814 (N_3814,N_3383,N_3159);
and U3815 (N_3815,N_3134,N_3095);
xnor U3816 (N_3816,N_3397,N_3291);
and U3817 (N_3817,N_3033,N_3030);
nand U3818 (N_3818,N_3097,N_3356);
and U3819 (N_3819,N_3458,N_3175);
xor U3820 (N_3820,N_3314,N_3122);
nor U3821 (N_3821,N_3102,N_3175);
nor U3822 (N_3822,N_3056,N_3225);
and U3823 (N_3823,N_3421,N_3029);
or U3824 (N_3824,N_3271,N_3170);
nand U3825 (N_3825,N_3205,N_3189);
or U3826 (N_3826,N_3333,N_3337);
or U3827 (N_3827,N_3014,N_3087);
xnor U3828 (N_3828,N_3460,N_3193);
or U3829 (N_3829,N_3167,N_3471);
or U3830 (N_3830,N_3053,N_3034);
or U3831 (N_3831,N_3457,N_3481);
xor U3832 (N_3832,N_3175,N_3132);
xor U3833 (N_3833,N_3213,N_3120);
and U3834 (N_3834,N_3340,N_3193);
nor U3835 (N_3835,N_3012,N_3462);
or U3836 (N_3836,N_3264,N_3097);
and U3837 (N_3837,N_3159,N_3201);
nor U3838 (N_3838,N_3075,N_3406);
and U3839 (N_3839,N_3065,N_3012);
nand U3840 (N_3840,N_3499,N_3318);
nand U3841 (N_3841,N_3224,N_3303);
or U3842 (N_3842,N_3101,N_3206);
and U3843 (N_3843,N_3074,N_3250);
or U3844 (N_3844,N_3438,N_3270);
nor U3845 (N_3845,N_3161,N_3109);
xnor U3846 (N_3846,N_3424,N_3028);
nor U3847 (N_3847,N_3002,N_3295);
nand U3848 (N_3848,N_3136,N_3091);
xor U3849 (N_3849,N_3361,N_3429);
or U3850 (N_3850,N_3353,N_3267);
nor U3851 (N_3851,N_3066,N_3164);
or U3852 (N_3852,N_3319,N_3322);
xor U3853 (N_3853,N_3062,N_3460);
nand U3854 (N_3854,N_3468,N_3070);
xor U3855 (N_3855,N_3290,N_3126);
and U3856 (N_3856,N_3243,N_3222);
or U3857 (N_3857,N_3286,N_3298);
or U3858 (N_3858,N_3103,N_3437);
nor U3859 (N_3859,N_3386,N_3058);
and U3860 (N_3860,N_3014,N_3203);
nand U3861 (N_3861,N_3180,N_3419);
xnor U3862 (N_3862,N_3254,N_3230);
nand U3863 (N_3863,N_3399,N_3008);
nor U3864 (N_3864,N_3033,N_3049);
xnor U3865 (N_3865,N_3084,N_3472);
nand U3866 (N_3866,N_3167,N_3151);
and U3867 (N_3867,N_3469,N_3422);
nand U3868 (N_3868,N_3394,N_3398);
xnor U3869 (N_3869,N_3031,N_3264);
and U3870 (N_3870,N_3284,N_3472);
xnor U3871 (N_3871,N_3066,N_3494);
nor U3872 (N_3872,N_3475,N_3042);
nor U3873 (N_3873,N_3050,N_3371);
xor U3874 (N_3874,N_3202,N_3155);
nand U3875 (N_3875,N_3232,N_3077);
and U3876 (N_3876,N_3372,N_3497);
and U3877 (N_3877,N_3279,N_3251);
nand U3878 (N_3878,N_3190,N_3284);
nor U3879 (N_3879,N_3346,N_3499);
nand U3880 (N_3880,N_3488,N_3419);
nand U3881 (N_3881,N_3026,N_3337);
nor U3882 (N_3882,N_3025,N_3337);
xor U3883 (N_3883,N_3295,N_3130);
nor U3884 (N_3884,N_3038,N_3264);
nor U3885 (N_3885,N_3121,N_3151);
nand U3886 (N_3886,N_3208,N_3279);
xor U3887 (N_3887,N_3156,N_3380);
nor U3888 (N_3888,N_3083,N_3377);
xor U3889 (N_3889,N_3062,N_3347);
nor U3890 (N_3890,N_3497,N_3269);
or U3891 (N_3891,N_3398,N_3039);
nand U3892 (N_3892,N_3310,N_3258);
nand U3893 (N_3893,N_3396,N_3309);
xor U3894 (N_3894,N_3256,N_3309);
nand U3895 (N_3895,N_3406,N_3464);
xnor U3896 (N_3896,N_3205,N_3425);
and U3897 (N_3897,N_3484,N_3204);
nor U3898 (N_3898,N_3010,N_3209);
or U3899 (N_3899,N_3273,N_3432);
nand U3900 (N_3900,N_3143,N_3115);
and U3901 (N_3901,N_3045,N_3190);
or U3902 (N_3902,N_3112,N_3325);
and U3903 (N_3903,N_3051,N_3042);
and U3904 (N_3904,N_3098,N_3263);
nand U3905 (N_3905,N_3271,N_3319);
nand U3906 (N_3906,N_3295,N_3265);
or U3907 (N_3907,N_3127,N_3449);
xnor U3908 (N_3908,N_3276,N_3138);
nand U3909 (N_3909,N_3136,N_3495);
nand U3910 (N_3910,N_3297,N_3125);
xor U3911 (N_3911,N_3436,N_3163);
or U3912 (N_3912,N_3304,N_3222);
xor U3913 (N_3913,N_3017,N_3260);
nand U3914 (N_3914,N_3073,N_3380);
and U3915 (N_3915,N_3117,N_3478);
and U3916 (N_3916,N_3334,N_3093);
or U3917 (N_3917,N_3431,N_3374);
nand U3918 (N_3918,N_3264,N_3057);
xor U3919 (N_3919,N_3372,N_3264);
xor U3920 (N_3920,N_3020,N_3437);
or U3921 (N_3921,N_3014,N_3484);
or U3922 (N_3922,N_3466,N_3327);
or U3923 (N_3923,N_3085,N_3320);
or U3924 (N_3924,N_3148,N_3132);
and U3925 (N_3925,N_3319,N_3065);
or U3926 (N_3926,N_3273,N_3111);
xnor U3927 (N_3927,N_3485,N_3053);
nor U3928 (N_3928,N_3095,N_3208);
xnor U3929 (N_3929,N_3174,N_3195);
and U3930 (N_3930,N_3021,N_3184);
nand U3931 (N_3931,N_3352,N_3194);
nand U3932 (N_3932,N_3141,N_3448);
and U3933 (N_3933,N_3499,N_3070);
xor U3934 (N_3934,N_3008,N_3035);
nand U3935 (N_3935,N_3013,N_3194);
and U3936 (N_3936,N_3242,N_3450);
nor U3937 (N_3937,N_3331,N_3385);
or U3938 (N_3938,N_3031,N_3145);
xnor U3939 (N_3939,N_3430,N_3228);
and U3940 (N_3940,N_3431,N_3250);
or U3941 (N_3941,N_3020,N_3360);
and U3942 (N_3942,N_3129,N_3369);
xnor U3943 (N_3943,N_3284,N_3199);
or U3944 (N_3944,N_3366,N_3374);
and U3945 (N_3945,N_3129,N_3358);
or U3946 (N_3946,N_3438,N_3378);
and U3947 (N_3947,N_3135,N_3223);
nor U3948 (N_3948,N_3383,N_3205);
and U3949 (N_3949,N_3353,N_3058);
nor U3950 (N_3950,N_3204,N_3454);
xnor U3951 (N_3951,N_3128,N_3213);
xor U3952 (N_3952,N_3053,N_3039);
nand U3953 (N_3953,N_3126,N_3461);
xor U3954 (N_3954,N_3221,N_3028);
nor U3955 (N_3955,N_3035,N_3232);
nand U3956 (N_3956,N_3056,N_3395);
or U3957 (N_3957,N_3161,N_3290);
nor U3958 (N_3958,N_3354,N_3038);
and U3959 (N_3959,N_3135,N_3487);
nand U3960 (N_3960,N_3428,N_3172);
nor U3961 (N_3961,N_3261,N_3044);
or U3962 (N_3962,N_3249,N_3239);
nor U3963 (N_3963,N_3085,N_3310);
nor U3964 (N_3964,N_3035,N_3007);
nand U3965 (N_3965,N_3050,N_3399);
xor U3966 (N_3966,N_3062,N_3456);
or U3967 (N_3967,N_3196,N_3471);
and U3968 (N_3968,N_3047,N_3220);
or U3969 (N_3969,N_3289,N_3384);
or U3970 (N_3970,N_3440,N_3342);
and U3971 (N_3971,N_3384,N_3328);
nor U3972 (N_3972,N_3301,N_3049);
nand U3973 (N_3973,N_3234,N_3182);
and U3974 (N_3974,N_3173,N_3408);
nor U3975 (N_3975,N_3210,N_3142);
nor U3976 (N_3976,N_3273,N_3340);
nand U3977 (N_3977,N_3488,N_3384);
or U3978 (N_3978,N_3458,N_3422);
or U3979 (N_3979,N_3083,N_3414);
xnor U3980 (N_3980,N_3201,N_3397);
and U3981 (N_3981,N_3373,N_3320);
nor U3982 (N_3982,N_3337,N_3382);
and U3983 (N_3983,N_3422,N_3244);
xnor U3984 (N_3984,N_3023,N_3376);
and U3985 (N_3985,N_3456,N_3491);
nand U3986 (N_3986,N_3077,N_3051);
xor U3987 (N_3987,N_3287,N_3075);
xor U3988 (N_3988,N_3386,N_3160);
xnor U3989 (N_3989,N_3172,N_3378);
or U3990 (N_3990,N_3228,N_3083);
nor U3991 (N_3991,N_3402,N_3031);
and U3992 (N_3992,N_3277,N_3028);
nand U3993 (N_3993,N_3454,N_3391);
and U3994 (N_3994,N_3237,N_3310);
nor U3995 (N_3995,N_3180,N_3080);
and U3996 (N_3996,N_3315,N_3338);
and U3997 (N_3997,N_3201,N_3320);
or U3998 (N_3998,N_3247,N_3060);
xnor U3999 (N_3999,N_3032,N_3373);
and U4000 (N_4000,N_3904,N_3558);
xnor U4001 (N_4001,N_3929,N_3534);
xnor U4002 (N_4002,N_3999,N_3885);
or U4003 (N_4003,N_3935,N_3646);
nor U4004 (N_4004,N_3568,N_3987);
nand U4005 (N_4005,N_3712,N_3598);
xnor U4006 (N_4006,N_3862,N_3849);
and U4007 (N_4007,N_3516,N_3892);
or U4008 (N_4008,N_3551,N_3599);
nand U4009 (N_4009,N_3776,N_3941);
nand U4010 (N_4010,N_3930,N_3691);
or U4011 (N_4011,N_3847,N_3798);
nand U4012 (N_4012,N_3890,N_3926);
or U4013 (N_4013,N_3730,N_3963);
nand U4014 (N_4014,N_3992,N_3834);
xor U4015 (N_4015,N_3986,N_3556);
nand U4016 (N_4016,N_3734,N_3920);
xor U4017 (N_4017,N_3616,N_3886);
xnor U4018 (N_4018,N_3677,N_3718);
xnor U4019 (N_4019,N_3803,N_3825);
xor U4020 (N_4020,N_3510,N_3619);
nor U4021 (N_4021,N_3660,N_3531);
or U4022 (N_4022,N_3940,N_3919);
nand U4023 (N_4023,N_3550,N_3770);
nand U4024 (N_4024,N_3968,N_3786);
xor U4025 (N_4025,N_3831,N_3756);
and U4026 (N_4026,N_3662,N_3910);
nand U4027 (N_4027,N_3896,N_3741);
and U4028 (N_4028,N_3864,N_3707);
and U4029 (N_4029,N_3539,N_3656);
or U4030 (N_4030,N_3973,N_3828);
nor U4031 (N_4031,N_3563,N_3580);
nand U4032 (N_4032,N_3965,N_3578);
and U4033 (N_4033,N_3693,N_3977);
or U4034 (N_4034,N_3735,N_3898);
or U4035 (N_4035,N_3912,N_3883);
nor U4036 (N_4036,N_3840,N_3713);
or U4037 (N_4037,N_3857,N_3674);
xor U4038 (N_4038,N_3595,N_3690);
xnor U4039 (N_4039,N_3855,N_3611);
nor U4040 (N_4040,N_3954,N_3975);
or U4041 (N_4041,N_3624,N_3789);
nand U4042 (N_4042,N_3925,N_3994);
nor U4043 (N_4043,N_3628,N_3879);
xor U4044 (N_4044,N_3924,N_3723);
nor U4045 (N_4045,N_3799,N_3811);
or U4046 (N_4046,N_3714,N_3873);
and U4047 (N_4047,N_3746,N_3576);
xnor U4048 (N_4048,N_3738,N_3805);
and U4049 (N_4049,N_3922,N_3774);
nand U4050 (N_4050,N_3566,N_3729);
nand U4051 (N_4051,N_3969,N_3715);
nand U4052 (N_4052,N_3848,N_3705);
and U4053 (N_4053,N_3983,N_3932);
nand U4054 (N_4054,N_3949,N_3654);
or U4055 (N_4055,N_3943,N_3856);
xor U4056 (N_4056,N_3765,N_3687);
nand U4057 (N_4057,N_3661,N_3575);
and U4058 (N_4058,N_3717,N_3570);
or U4059 (N_4059,N_3976,N_3638);
or U4060 (N_4060,N_3763,N_3518);
nor U4061 (N_4061,N_3870,N_3978);
and U4062 (N_4062,N_3988,N_3793);
or U4063 (N_4063,N_3683,N_3720);
or U4064 (N_4064,N_3569,N_3980);
xor U4065 (N_4065,N_3945,N_3821);
and U4066 (N_4066,N_3812,N_3685);
xnor U4067 (N_4067,N_3990,N_3801);
and U4068 (N_4068,N_3901,N_3752);
nor U4069 (N_4069,N_3525,N_3944);
nor U4070 (N_4070,N_3701,N_3547);
xnor U4071 (N_4071,N_3500,N_3727);
nor U4072 (N_4072,N_3546,N_3952);
and U4073 (N_4073,N_3582,N_3911);
nand U4074 (N_4074,N_3989,N_3744);
nor U4075 (N_4075,N_3652,N_3958);
or U4076 (N_4076,N_3647,N_3781);
and U4077 (N_4077,N_3863,N_3917);
nor U4078 (N_4078,N_3553,N_3900);
nand U4079 (N_4079,N_3617,N_3884);
nand U4080 (N_4080,N_3692,N_3615);
and U4081 (N_4081,N_3841,N_3521);
xnor U4082 (N_4082,N_3505,N_3782);
xor U4083 (N_4083,N_3875,N_3796);
or U4084 (N_4084,N_3626,N_3893);
xor U4085 (N_4085,N_3645,N_3508);
or U4086 (N_4086,N_3565,N_3621);
and U4087 (N_4087,N_3915,N_3750);
and U4088 (N_4088,N_3544,N_3775);
xor U4089 (N_4089,N_3788,N_3827);
nor U4090 (N_4090,N_3514,N_3633);
or U4091 (N_4091,N_3991,N_3676);
or U4092 (N_4092,N_3607,N_3635);
xnor U4093 (N_4093,N_3623,N_3842);
or U4094 (N_4094,N_3532,N_3529);
or U4095 (N_4095,N_3522,N_3536);
xor U4096 (N_4096,N_3506,N_3794);
nand U4097 (N_4097,N_3942,N_3609);
and U4098 (N_4098,N_3610,N_3533);
or U4099 (N_4099,N_3631,N_3970);
nand U4100 (N_4100,N_3806,N_3823);
and U4101 (N_4101,N_3923,N_3948);
or U4102 (N_4102,N_3585,N_3928);
nor U4103 (N_4103,N_3588,N_3903);
xnor U4104 (N_4104,N_3689,N_3972);
or U4105 (N_4105,N_3780,N_3622);
nand U4106 (N_4106,N_3916,N_3829);
nand U4107 (N_4107,N_3837,N_3725);
nor U4108 (N_4108,N_3555,N_3597);
nor U4109 (N_4109,N_3709,N_3760);
nor U4110 (N_4110,N_3982,N_3981);
nor U4111 (N_4111,N_3680,N_3759);
nand U4112 (N_4112,N_3613,N_3955);
nor U4113 (N_4113,N_3951,N_3519);
nor U4114 (N_4114,N_3655,N_3854);
nor U4115 (N_4115,N_3634,N_3636);
nor U4116 (N_4116,N_3542,N_3913);
and U4117 (N_4117,N_3785,N_3927);
and U4118 (N_4118,N_3814,N_3858);
nand U4119 (N_4119,N_3504,N_3523);
nor U4120 (N_4120,N_3888,N_3846);
nand U4121 (N_4121,N_3771,N_3819);
xnor U4122 (N_4122,N_3953,N_3562);
nand U4123 (N_4123,N_3853,N_3810);
nand U4124 (N_4124,N_3758,N_3743);
xor U4125 (N_4125,N_3754,N_3665);
or U4126 (N_4126,N_3807,N_3719);
nand U4127 (N_4127,N_3722,N_3669);
nand U4128 (N_4128,N_3843,N_3509);
nor U4129 (N_4129,N_3632,N_3543);
or U4130 (N_4130,N_3748,N_3561);
nand U4131 (N_4131,N_3699,N_3820);
xor U4132 (N_4132,N_3902,N_3637);
and U4133 (N_4133,N_3600,N_3502);
nand U4134 (N_4134,N_3675,N_3962);
nand U4135 (N_4135,N_3557,N_3947);
and U4136 (N_4136,N_3753,N_3737);
and U4137 (N_4137,N_3618,N_3700);
or U4138 (N_4138,N_3587,N_3844);
xor U4139 (N_4139,N_3629,N_3710);
nor U4140 (N_4140,N_3967,N_3736);
or U4141 (N_4141,N_3959,N_3804);
nor U4142 (N_4142,N_3696,N_3815);
xnor U4143 (N_4143,N_3984,N_3653);
nand U4144 (N_4144,N_3868,N_3559);
and U4145 (N_4145,N_3914,N_3836);
xnor U4146 (N_4146,N_3605,N_3596);
nand U4147 (N_4147,N_3797,N_3956);
or U4148 (N_4148,N_3809,N_3768);
nor U4149 (N_4149,N_3839,N_3971);
nor U4150 (N_4150,N_3520,N_3957);
nand U4151 (N_4151,N_3998,N_3874);
or U4152 (N_4152,N_3581,N_3603);
nor U4153 (N_4153,N_3790,N_3591);
xnor U4154 (N_4154,N_3711,N_3740);
nor U4155 (N_4155,N_3688,N_3933);
and U4156 (N_4156,N_3813,N_3643);
and U4157 (N_4157,N_3777,N_3937);
nand U4158 (N_4158,N_3800,N_3871);
nor U4159 (N_4159,N_3921,N_3572);
and U4160 (N_4160,N_3650,N_3757);
and U4161 (N_4161,N_3515,N_3501);
xor U4162 (N_4162,N_3835,N_3918);
nor U4163 (N_4163,N_3627,N_3540);
nor U4164 (N_4164,N_3589,N_3802);
nand U4165 (N_4165,N_3773,N_3644);
xnor U4166 (N_4166,N_3877,N_3878);
xnor U4167 (N_4167,N_3684,N_3818);
nand U4168 (N_4168,N_3851,N_3946);
or U4169 (N_4169,N_3649,N_3733);
nand U4170 (N_4170,N_3865,N_3961);
xor U4171 (N_4171,N_3985,N_3538);
and U4172 (N_4172,N_3511,N_3872);
nor U4173 (N_4173,N_3996,N_3779);
nand U4174 (N_4174,N_3584,N_3887);
and U4175 (N_4175,N_3824,N_3755);
xnor U4176 (N_4176,N_3974,N_3826);
and U4177 (N_4177,N_3641,N_3663);
xor U4178 (N_4178,N_3784,N_3880);
nand U4179 (N_4179,N_3860,N_3772);
nor U4180 (N_4180,N_3528,N_3651);
nor U4181 (N_4181,N_3751,N_3664);
and U4182 (N_4182,N_3537,N_3778);
xor U4183 (N_4183,N_3728,N_3545);
and U4184 (N_4184,N_3732,N_3833);
nand U4185 (N_4185,N_3672,N_3995);
and U4186 (N_4186,N_3716,N_3808);
xor U4187 (N_4187,N_3724,N_3592);
xor U4188 (N_4188,N_3869,N_3993);
nand U4189 (N_4189,N_3642,N_3666);
nand U4190 (N_4190,N_3747,N_3601);
nand U4191 (N_4191,N_3731,N_3608);
nor U4192 (N_4192,N_3934,N_3979);
xnor U4193 (N_4193,N_3960,N_3697);
nand U4194 (N_4194,N_3703,N_3671);
xor U4195 (N_4195,N_3614,N_3548);
and U4196 (N_4196,N_3891,N_3657);
nand U4197 (N_4197,N_3907,N_3630);
and U4198 (N_4198,N_3567,N_3742);
or U4199 (N_4199,N_3560,N_3861);
or U4200 (N_4200,N_3706,N_3530);
or U4201 (N_4201,N_3524,N_3552);
and U4202 (N_4202,N_3507,N_3964);
and U4203 (N_4203,N_3698,N_3606);
nand U4204 (N_4204,N_3909,N_3830);
nor U4205 (N_4205,N_3586,N_3850);
or U4206 (N_4206,N_3702,N_3997);
and U4207 (N_4207,N_3517,N_3554);
and U4208 (N_4208,N_3764,N_3593);
xnor U4209 (N_4209,N_3549,N_3721);
nor U4210 (N_4210,N_3658,N_3604);
and U4211 (N_4211,N_3881,N_3761);
nor U4212 (N_4212,N_3571,N_3620);
xnor U4213 (N_4213,N_3648,N_3749);
nand U4214 (N_4214,N_3708,N_3897);
nor U4215 (N_4215,N_3899,N_3704);
nor U4216 (N_4216,N_3667,N_3859);
or U4217 (N_4217,N_3938,N_3577);
xnor U4218 (N_4218,N_3791,N_3678);
nand U4219 (N_4219,N_3822,N_3762);
nor U4220 (N_4220,N_3889,N_3590);
or U4221 (N_4221,N_3838,N_3659);
and U4222 (N_4222,N_3866,N_3845);
xnor U4223 (N_4223,N_3908,N_3745);
or U4224 (N_4224,N_3939,N_3679);
xnor U4225 (N_4225,N_3906,N_3931);
nand U4226 (N_4226,N_3695,N_3640);
xor U4227 (N_4227,N_3950,N_3513);
and U4228 (N_4228,N_3668,N_3816);
xor U4229 (N_4229,N_3579,N_3726);
and U4230 (N_4230,N_3876,N_3795);
nor U4231 (N_4231,N_3612,N_3512);
nor U4232 (N_4232,N_3882,N_3527);
and U4233 (N_4233,N_3766,N_3686);
xnor U4234 (N_4234,N_3594,N_3852);
xnor U4235 (N_4235,N_3625,N_3867);
nor U4236 (N_4236,N_3574,N_3966);
and U4237 (N_4237,N_3767,N_3895);
and U4238 (N_4238,N_3670,N_3503);
xnor U4239 (N_4239,N_3832,N_3681);
nor U4240 (N_4240,N_3535,N_3526);
xnor U4241 (N_4241,N_3682,N_3787);
and U4242 (N_4242,N_3783,N_3792);
nor U4243 (N_4243,N_3769,N_3564);
or U4244 (N_4244,N_3673,N_3694);
nand U4245 (N_4245,N_3936,N_3573);
nand U4246 (N_4246,N_3639,N_3817);
or U4247 (N_4247,N_3583,N_3602);
nand U4248 (N_4248,N_3541,N_3739);
nor U4249 (N_4249,N_3905,N_3894);
xor U4250 (N_4250,N_3554,N_3769);
xor U4251 (N_4251,N_3843,N_3850);
nand U4252 (N_4252,N_3660,N_3933);
and U4253 (N_4253,N_3669,N_3698);
and U4254 (N_4254,N_3534,N_3839);
xnor U4255 (N_4255,N_3829,N_3651);
nor U4256 (N_4256,N_3843,N_3608);
nor U4257 (N_4257,N_3864,N_3603);
nor U4258 (N_4258,N_3692,N_3728);
or U4259 (N_4259,N_3629,N_3860);
xnor U4260 (N_4260,N_3801,N_3675);
and U4261 (N_4261,N_3847,N_3581);
nand U4262 (N_4262,N_3690,N_3985);
and U4263 (N_4263,N_3836,N_3530);
nand U4264 (N_4264,N_3584,N_3793);
and U4265 (N_4265,N_3789,N_3766);
nor U4266 (N_4266,N_3594,N_3887);
nor U4267 (N_4267,N_3519,N_3752);
nor U4268 (N_4268,N_3832,N_3811);
nand U4269 (N_4269,N_3704,N_3867);
or U4270 (N_4270,N_3587,N_3664);
xnor U4271 (N_4271,N_3739,N_3917);
xnor U4272 (N_4272,N_3605,N_3837);
xor U4273 (N_4273,N_3999,N_3972);
and U4274 (N_4274,N_3921,N_3530);
xor U4275 (N_4275,N_3684,N_3946);
and U4276 (N_4276,N_3970,N_3750);
xnor U4277 (N_4277,N_3579,N_3905);
or U4278 (N_4278,N_3890,N_3641);
and U4279 (N_4279,N_3827,N_3815);
nor U4280 (N_4280,N_3753,N_3760);
nor U4281 (N_4281,N_3732,N_3663);
and U4282 (N_4282,N_3969,N_3920);
nand U4283 (N_4283,N_3760,N_3663);
nand U4284 (N_4284,N_3930,N_3945);
nand U4285 (N_4285,N_3928,N_3627);
nor U4286 (N_4286,N_3693,N_3667);
xor U4287 (N_4287,N_3981,N_3878);
nor U4288 (N_4288,N_3572,N_3504);
nand U4289 (N_4289,N_3725,N_3621);
and U4290 (N_4290,N_3971,N_3786);
xor U4291 (N_4291,N_3529,N_3628);
nand U4292 (N_4292,N_3999,N_3547);
and U4293 (N_4293,N_3614,N_3722);
nor U4294 (N_4294,N_3986,N_3745);
or U4295 (N_4295,N_3922,N_3991);
or U4296 (N_4296,N_3713,N_3962);
xor U4297 (N_4297,N_3551,N_3670);
and U4298 (N_4298,N_3986,N_3981);
nand U4299 (N_4299,N_3598,N_3833);
or U4300 (N_4300,N_3513,N_3566);
xnor U4301 (N_4301,N_3910,N_3863);
xnor U4302 (N_4302,N_3747,N_3502);
nand U4303 (N_4303,N_3641,N_3510);
nand U4304 (N_4304,N_3525,N_3740);
xor U4305 (N_4305,N_3876,N_3532);
nor U4306 (N_4306,N_3887,N_3555);
and U4307 (N_4307,N_3514,N_3962);
and U4308 (N_4308,N_3509,N_3629);
nor U4309 (N_4309,N_3690,N_3960);
nor U4310 (N_4310,N_3803,N_3968);
or U4311 (N_4311,N_3712,N_3908);
nand U4312 (N_4312,N_3818,N_3756);
nor U4313 (N_4313,N_3924,N_3783);
nand U4314 (N_4314,N_3516,N_3614);
nor U4315 (N_4315,N_3685,N_3507);
xor U4316 (N_4316,N_3668,N_3932);
nor U4317 (N_4317,N_3935,N_3752);
nand U4318 (N_4318,N_3758,N_3842);
xor U4319 (N_4319,N_3905,N_3790);
and U4320 (N_4320,N_3909,N_3975);
or U4321 (N_4321,N_3684,N_3829);
nand U4322 (N_4322,N_3670,N_3847);
nand U4323 (N_4323,N_3954,N_3918);
and U4324 (N_4324,N_3782,N_3619);
and U4325 (N_4325,N_3638,N_3820);
and U4326 (N_4326,N_3532,N_3973);
or U4327 (N_4327,N_3688,N_3574);
and U4328 (N_4328,N_3521,N_3924);
xor U4329 (N_4329,N_3977,N_3757);
xnor U4330 (N_4330,N_3532,N_3796);
nand U4331 (N_4331,N_3621,N_3936);
and U4332 (N_4332,N_3782,N_3617);
and U4333 (N_4333,N_3919,N_3733);
or U4334 (N_4334,N_3817,N_3913);
or U4335 (N_4335,N_3682,N_3708);
and U4336 (N_4336,N_3880,N_3664);
nand U4337 (N_4337,N_3900,N_3870);
nand U4338 (N_4338,N_3631,N_3913);
nand U4339 (N_4339,N_3977,N_3792);
or U4340 (N_4340,N_3715,N_3917);
xnor U4341 (N_4341,N_3685,N_3970);
or U4342 (N_4342,N_3845,N_3943);
or U4343 (N_4343,N_3559,N_3583);
and U4344 (N_4344,N_3854,N_3573);
nor U4345 (N_4345,N_3827,N_3727);
nor U4346 (N_4346,N_3515,N_3566);
or U4347 (N_4347,N_3831,N_3615);
or U4348 (N_4348,N_3536,N_3792);
nand U4349 (N_4349,N_3942,N_3528);
nand U4350 (N_4350,N_3796,N_3540);
or U4351 (N_4351,N_3554,N_3861);
nor U4352 (N_4352,N_3569,N_3620);
nor U4353 (N_4353,N_3942,N_3627);
or U4354 (N_4354,N_3909,N_3856);
or U4355 (N_4355,N_3903,N_3513);
and U4356 (N_4356,N_3889,N_3943);
and U4357 (N_4357,N_3533,N_3548);
xor U4358 (N_4358,N_3816,N_3961);
nand U4359 (N_4359,N_3862,N_3541);
nand U4360 (N_4360,N_3662,N_3892);
nor U4361 (N_4361,N_3827,N_3865);
or U4362 (N_4362,N_3610,N_3906);
nor U4363 (N_4363,N_3809,N_3720);
nand U4364 (N_4364,N_3534,N_3758);
nor U4365 (N_4365,N_3620,N_3528);
nand U4366 (N_4366,N_3900,N_3824);
nor U4367 (N_4367,N_3696,N_3855);
xnor U4368 (N_4368,N_3703,N_3717);
and U4369 (N_4369,N_3906,N_3972);
nor U4370 (N_4370,N_3610,N_3621);
nand U4371 (N_4371,N_3589,N_3645);
and U4372 (N_4372,N_3531,N_3617);
xor U4373 (N_4373,N_3896,N_3703);
xor U4374 (N_4374,N_3936,N_3575);
xnor U4375 (N_4375,N_3856,N_3872);
nor U4376 (N_4376,N_3594,N_3763);
or U4377 (N_4377,N_3612,N_3609);
or U4378 (N_4378,N_3674,N_3855);
nand U4379 (N_4379,N_3665,N_3880);
and U4380 (N_4380,N_3717,N_3810);
and U4381 (N_4381,N_3616,N_3769);
xor U4382 (N_4382,N_3911,N_3528);
nand U4383 (N_4383,N_3548,N_3877);
nor U4384 (N_4384,N_3680,N_3843);
nor U4385 (N_4385,N_3806,N_3659);
nand U4386 (N_4386,N_3660,N_3976);
nand U4387 (N_4387,N_3503,N_3613);
and U4388 (N_4388,N_3833,N_3713);
and U4389 (N_4389,N_3850,N_3858);
and U4390 (N_4390,N_3546,N_3698);
nand U4391 (N_4391,N_3742,N_3919);
nand U4392 (N_4392,N_3924,N_3713);
nand U4393 (N_4393,N_3733,N_3760);
and U4394 (N_4394,N_3934,N_3917);
xnor U4395 (N_4395,N_3527,N_3757);
nand U4396 (N_4396,N_3739,N_3660);
nand U4397 (N_4397,N_3751,N_3669);
or U4398 (N_4398,N_3866,N_3615);
xnor U4399 (N_4399,N_3519,N_3719);
xor U4400 (N_4400,N_3909,N_3820);
and U4401 (N_4401,N_3998,N_3875);
nor U4402 (N_4402,N_3574,N_3683);
xor U4403 (N_4403,N_3502,N_3858);
nor U4404 (N_4404,N_3941,N_3896);
and U4405 (N_4405,N_3759,N_3728);
nand U4406 (N_4406,N_3555,N_3552);
xor U4407 (N_4407,N_3609,N_3761);
xnor U4408 (N_4408,N_3689,N_3887);
or U4409 (N_4409,N_3846,N_3690);
nand U4410 (N_4410,N_3938,N_3766);
nor U4411 (N_4411,N_3560,N_3602);
nor U4412 (N_4412,N_3874,N_3628);
nor U4413 (N_4413,N_3565,N_3806);
and U4414 (N_4414,N_3814,N_3589);
nand U4415 (N_4415,N_3943,N_3728);
or U4416 (N_4416,N_3729,N_3839);
nand U4417 (N_4417,N_3595,N_3713);
and U4418 (N_4418,N_3691,N_3803);
nor U4419 (N_4419,N_3828,N_3700);
xor U4420 (N_4420,N_3935,N_3728);
or U4421 (N_4421,N_3805,N_3876);
and U4422 (N_4422,N_3617,N_3844);
and U4423 (N_4423,N_3635,N_3544);
xor U4424 (N_4424,N_3708,N_3909);
or U4425 (N_4425,N_3704,N_3709);
nand U4426 (N_4426,N_3590,N_3979);
nand U4427 (N_4427,N_3505,N_3699);
or U4428 (N_4428,N_3656,N_3954);
and U4429 (N_4429,N_3790,N_3963);
xnor U4430 (N_4430,N_3906,N_3934);
and U4431 (N_4431,N_3556,N_3799);
xor U4432 (N_4432,N_3545,N_3618);
or U4433 (N_4433,N_3588,N_3634);
nand U4434 (N_4434,N_3551,N_3829);
or U4435 (N_4435,N_3743,N_3576);
nor U4436 (N_4436,N_3672,N_3736);
nor U4437 (N_4437,N_3713,N_3887);
nor U4438 (N_4438,N_3651,N_3580);
and U4439 (N_4439,N_3799,N_3797);
and U4440 (N_4440,N_3534,N_3658);
nor U4441 (N_4441,N_3720,N_3830);
and U4442 (N_4442,N_3556,N_3977);
nand U4443 (N_4443,N_3669,N_3640);
nand U4444 (N_4444,N_3969,N_3859);
xnor U4445 (N_4445,N_3517,N_3557);
or U4446 (N_4446,N_3923,N_3798);
nor U4447 (N_4447,N_3857,N_3507);
nand U4448 (N_4448,N_3672,N_3692);
xor U4449 (N_4449,N_3959,N_3668);
or U4450 (N_4450,N_3682,N_3978);
xnor U4451 (N_4451,N_3818,N_3585);
xor U4452 (N_4452,N_3594,N_3901);
and U4453 (N_4453,N_3573,N_3630);
nand U4454 (N_4454,N_3910,N_3739);
or U4455 (N_4455,N_3507,N_3687);
or U4456 (N_4456,N_3676,N_3926);
nor U4457 (N_4457,N_3949,N_3988);
nor U4458 (N_4458,N_3641,N_3976);
xnor U4459 (N_4459,N_3837,N_3796);
or U4460 (N_4460,N_3746,N_3769);
or U4461 (N_4461,N_3664,N_3780);
and U4462 (N_4462,N_3852,N_3581);
xnor U4463 (N_4463,N_3817,N_3648);
or U4464 (N_4464,N_3615,N_3686);
nand U4465 (N_4465,N_3654,N_3572);
nor U4466 (N_4466,N_3695,N_3791);
nand U4467 (N_4467,N_3648,N_3885);
and U4468 (N_4468,N_3724,N_3807);
nand U4469 (N_4469,N_3877,N_3945);
or U4470 (N_4470,N_3935,N_3809);
or U4471 (N_4471,N_3504,N_3998);
and U4472 (N_4472,N_3563,N_3585);
or U4473 (N_4473,N_3890,N_3980);
and U4474 (N_4474,N_3877,N_3671);
and U4475 (N_4475,N_3662,N_3549);
nor U4476 (N_4476,N_3913,N_3816);
or U4477 (N_4477,N_3962,N_3669);
nor U4478 (N_4478,N_3951,N_3768);
xnor U4479 (N_4479,N_3550,N_3949);
or U4480 (N_4480,N_3824,N_3666);
and U4481 (N_4481,N_3775,N_3761);
xor U4482 (N_4482,N_3718,N_3748);
and U4483 (N_4483,N_3699,N_3731);
nor U4484 (N_4484,N_3608,N_3974);
or U4485 (N_4485,N_3574,N_3840);
or U4486 (N_4486,N_3745,N_3771);
xnor U4487 (N_4487,N_3678,N_3507);
xnor U4488 (N_4488,N_3942,N_3553);
nand U4489 (N_4489,N_3869,N_3888);
nor U4490 (N_4490,N_3919,N_3955);
or U4491 (N_4491,N_3904,N_3658);
or U4492 (N_4492,N_3992,N_3720);
or U4493 (N_4493,N_3604,N_3646);
nand U4494 (N_4494,N_3841,N_3538);
nand U4495 (N_4495,N_3830,N_3520);
or U4496 (N_4496,N_3970,N_3834);
nor U4497 (N_4497,N_3592,N_3524);
and U4498 (N_4498,N_3530,N_3930);
nor U4499 (N_4499,N_3731,N_3625);
nor U4500 (N_4500,N_4205,N_4360);
xnor U4501 (N_4501,N_4022,N_4366);
xor U4502 (N_4502,N_4142,N_4035);
nor U4503 (N_4503,N_4485,N_4181);
nor U4504 (N_4504,N_4212,N_4400);
nand U4505 (N_4505,N_4418,N_4389);
or U4506 (N_4506,N_4325,N_4337);
nand U4507 (N_4507,N_4346,N_4017);
nand U4508 (N_4508,N_4206,N_4277);
or U4509 (N_4509,N_4042,N_4156);
xor U4510 (N_4510,N_4113,N_4241);
or U4511 (N_4511,N_4476,N_4008);
nor U4512 (N_4512,N_4315,N_4031);
nor U4513 (N_4513,N_4417,N_4421);
nor U4514 (N_4514,N_4268,N_4061);
and U4515 (N_4515,N_4353,N_4459);
or U4516 (N_4516,N_4495,N_4221);
xor U4517 (N_4517,N_4146,N_4333);
nand U4518 (N_4518,N_4180,N_4135);
nand U4519 (N_4519,N_4129,N_4009);
nand U4520 (N_4520,N_4455,N_4356);
xnor U4521 (N_4521,N_4000,N_4154);
nor U4522 (N_4522,N_4380,N_4460);
and U4523 (N_4523,N_4060,N_4342);
xor U4524 (N_4524,N_4273,N_4287);
xnor U4525 (N_4525,N_4139,N_4238);
xor U4526 (N_4526,N_4313,N_4046);
nand U4527 (N_4527,N_4102,N_4321);
or U4528 (N_4528,N_4453,N_4219);
xnor U4529 (N_4529,N_4288,N_4168);
nor U4530 (N_4530,N_4249,N_4236);
nor U4531 (N_4531,N_4263,N_4220);
nand U4532 (N_4532,N_4014,N_4422);
and U4533 (N_4533,N_4358,N_4178);
nor U4534 (N_4534,N_4209,N_4449);
xnor U4535 (N_4535,N_4292,N_4493);
and U4536 (N_4536,N_4222,N_4271);
nand U4537 (N_4537,N_4118,N_4062);
xnor U4538 (N_4538,N_4368,N_4450);
or U4539 (N_4539,N_4112,N_4085);
and U4540 (N_4540,N_4413,N_4006);
or U4541 (N_4541,N_4210,N_4057);
xnor U4542 (N_4542,N_4053,N_4433);
nand U4543 (N_4543,N_4120,N_4477);
and U4544 (N_4544,N_4410,N_4279);
nor U4545 (N_4545,N_4496,N_4303);
xnor U4546 (N_4546,N_4441,N_4378);
nand U4547 (N_4547,N_4174,N_4081);
and U4548 (N_4548,N_4444,N_4474);
xor U4549 (N_4549,N_4141,N_4247);
xnor U4550 (N_4550,N_4003,N_4098);
or U4551 (N_4551,N_4392,N_4470);
nand U4552 (N_4552,N_4038,N_4276);
nor U4553 (N_4553,N_4225,N_4330);
and U4554 (N_4554,N_4369,N_4281);
nor U4555 (N_4555,N_4432,N_4108);
nor U4556 (N_4556,N_4160,N_4448);
or U4557 (N_4557,N_4072,N_4213);
nor U4558 (N_4558,N_4004,N_4089);
nand U4559 (N_4559,N_4403,N_4078);
and U4560 (N_4560,N_4295,N_4111);
or U4561 (N_4561,N_4254,N_4335);
nand U4562 (N_4562,N_4483,N_4384);
and U4563 (N_4563,N_4040,N_4037);
or U4564 (N_4564,N_4179,N_4253);
xnor U4565 (N_4565,N_4059,N_4331);
nor U4566 (N_4566,N_4188,N_4486);
nor U4567 (N_4567,N_4226,N_4364);
or U4568 (N_4568,N_4322,N_4068);
nor U4569 (N_4569,N_4116,N_4355);
nand U4570 (N_4570,N_4257,N_4001);
xor U4571 (N_4571,N_4186,N_4265);
or U4572 (N_4572,N_4039,N_4250);
and U4573 (N_4573,N_4045,N_4148);
nor U4574 (N_4574,N_4434,N_4379);
or U4575 (N_4575,N_4291,N_4164);
xor U4576 (N_4576,N_4370,N_4352);
and U4577 (N_4577,N_4310,N_4475);
and U4578 (N_4578,N_4324,N_4391);
nand U4579 (N_4579,N_4165,N_4282);
nor U4580 (N_4580,N_4275,N_4077);
and U4581 (N_4581,N_4079,N_4056);
nand U4582 (N_4582,N_4018,N_4147);
or U4583 (N_4583,N_4308,N_4130);
xnor U4584 (N_4584,N_4013,N_4076);
and U4585 (N_4585,N_4479,N_4248);
and U4586 (N_4586,N_4350,N_4131);
or U4587 (N_4587,N_4065,N_4176);
nor U4588 (N_4588,N_4399,N_4159);
and U4589 (N_4589,N_4161,N_4363);
xnor U4590 (N_4590,N_4240,N_4233);
and U4591 (N_4591,N_4052,N_4266);
nor U4592 (N_4592,N_4471,N_4465);
nor U4593 (N_4593,N_4468,N_4122);
and U4594 (N_4594,N_4357,N_4151);
or U4595 (N_4595,N_4223,N_4019);
nor U4596 (N_4596,N_4296,N_4317);
nor U4597 (N_4597,N_4411,N_4182);
xnor U4598 (N_4598,N_4497,N_4283);
nand U4599 (N_4599,N_4442,N_4184);
xor U4600 (N_4600,N_4105,N_4446);
nor U4601 (N_4601,N_4099,N_4383);
and U4602 (N_4602,N_4048,N_4203);
and U4603 (N_4603,N_4096,N_4478);
and U4604 (N_4604,N_4304,N_4242);
nor U4605 (N_4605,N_4097,N_4447);
and U4606 (N_4606,N_4101,N_4239);
nand U4607 (N_4607,N_4351,N_4034);
nor U4608 (N_4608,N_4149,N_4030);
or U4609 (N_4609,N_4067,N_4252);
nand U4610 (N_4610,N_4426,N_4316);
and U4611 (N_4611,N_4211,N_4466);
or U4612 (N_4612,N_4187,N_4332);
and U4613 (N_4613,N_4454,N_4290);
nor U4614 (N_4614,N_4153,N_4336);
or U4615 (N_4615,N_4145,N_4472);
xnor U4616 (N_4616,N_4199,N_4372);
or U4617 (N_4617,N_4484,N_4436);
nand U4618 (N_4618,N_4083,N_4082);
or U4619 (N_4619,N_4069,N_4329);
nand U4620 (N_4620,N_4104,N_4347);
or U4621 (N_4621,N_4150,N_4367);
xor U4622 (N_4622,N_4393,N_4469);
xnor U4623 (N_4623,N_4404,N_4086);
nor U4624 (N_4624,N_4084,N_4032);
or U4625 (N_4625,N_4138,N_4216);
and U4626 (N_4626,N_4488,N_4390);
or U4627 (N_4627,N_4259,N_4464);
and U4628 (N_4628,N_4396,N_4088);
or U4629 (N_4629,N_4294,N_4318);
or U4630 (N_4630,N_4415,N_4299);
and U4631 (N_4631,N_4215,N_4015);
xnor U4632 (N_4632,N_4090,N_4409);
nand U4633 (N_4633,N_4091,N_4002);
and U4634 (N_4634,N_4467,N_4234);
xnor U4635 (N_4635,N_4232,N_4406);
xor U4636 (N_4636,N_4043,N_4218);
nor U4637 (N_4637,N_4094,N_4445);
nor U4638 (N_4638,N_4058,N_4201);
xor U4639 (N_4639,N_4024,N_4298);
nor U4640 (N_4640,N_4049,N_4498);
xor U4641 (N_4641,N_4345,N_4386);
nor U4642 (N_4642,N_4115,N_4319);
xnor U4643 (N_4643,N_4231,N_4439);
or U4644 (N_4644,N_4388,N_4229);
or U4645 (N_4645,N_4327,N_4286);
or U4646 (N_4646,N_4284,N_4246);
or U4647 (N_4647,N_4051,N_4354);
nor U4648 (N_4648,N_4121,N_4026);
nand U4649 (N_4649,N_4152,N_4087);
nor U4650 (N_4650,N_4126,N_4425);
nand U4651 (N_4651,N_4012,N_4258);
nor U4652 (N_4652,N_4103,N_4424);
xnor U4653 (N_4653,N_4193,N_4237);
xor U4654 (N_4654,N_4341,N_4143);
and U4655 (N_4655,N_4194,N_4419);
nand U4656 (N_4656,N_4323,N_4050);
or U4657 (N_4657,N_4029,N_4124);
and U4658 (N_4658,N_4344,N_4371);
nor U4659 (N_4659,N_4423,N_4414);
nor U4660 (N_4660,N_4270,N_4499);
and U4661 (N_4661,N_4402,N_4398);
nand U4662 (N_4662,N_4093,N_4462);
and U4663 (N_4663,N_4373,N_4440);
nor U4664 (N_4664,N_4492,N_4195);
xnor U4665 (N_4665,N_4463,N_4071);
nand U4666 (N_4666,N_4243,N_4457);
nand U4667 (N_4667,N_4262,N_4267);
nand U4668 (N_4668,N_4311,N_4016);
and U4669 (N_4669,N_4044,N_4197);
nand U4670 (N_4670,N_4169,N_4435);
and U4671 (N_4671,N_4166,N_4438);
nand U4672 (N_4672,N_4487,N_4306);
nand U4673 (N_4673,N_4280,N_4170);
nor U4674 (N_4674,N_4244,N_4010);
or U4675 (N_4675,N_4027,N_4070);
nand U4676 (N_4676,N_4293,N_4494);
nor U4677 (N_4677,N_4063,N_4173);
nand U4678 (N_4678,N_4359,N_4005);
nor U4679 (N_4679,N_4309,N_4451);
and U4680 (N_4680,N_4461,N_4066);
nor U4681 (N_4681,N_4054,N_4362);
and U4682 (N_4682,N_4140,N_4007);
or U4683 (N_4683,N_4274,N_4167);
and U4684 (N_4684,N_4123,N_4340);
and U4685 (N_4685,N_4036,N_4075);
or U4686 (N_4686,N_4204,N_4264);
nand U4687 (N_4687,N_4109,N_4202);
or U4688 (N_4688,N_4261,N_4397);
and U4689 (N_4689,N_4020,N_4339);
nor U4690 (N_4690,N_4155,N_4128);
nor U4691 (N_4691,N_4385,N_4073);
nor U4692 (N_4692,N_4443,N_4033);
or U4693 (N_4693,N_4177,N_4133);
xor U4694 (N_4694,N_4348,N_4100);
and U4695 (N_4695,N_4055,N_4480);
xor U4696 (N_4696,N_4437,N_4134);
or U4697 (N_4697,N_4365,N_4387);
nand U4698 (N_4698,N_4300,N_4207);
nand U4699 (N_4699,N_4278,N_4183);
nor U4700 (N_4700,N_4107,N_4456);
xnor U4701 (N_4701,N_4080,N_4431);
xor U4702 (N_4702,N_4190,N_4458);
and U4703 (N_4703,N_4428,N_4407);
or U4704 (N_4704,N_4191,N_4256);
and U4705 (N_4705,N_4157,N_4320);
nand U4706 (N_4706,N_4158,N_4095);
nor U4707 (N_4707,N_4289,N_4361);
nor U4708 (N_4708,N_4416,N_4137);
or U4709 (N_4709,N_4338,N_4343);
and U4710 (N_4710,N_4011,N_4175);
and U4711 (N_4711,N_4047,N_4021);
and U4712 (N_4712,N_4114,N_4376);
nor U4713 (N_4713,N_4189,N_4028);
nor U4714 (N_4714,N_4196,N_4490);
xor U4715 (N_4715,N_4375,N_4132);
xor U4716 (N_4716,N_4214,N_4395);
nor U4717 (N_4717,N_4307,N_4489);
or U4718 (N_4718,N_4305,N_4382);
xnor U4719 (N_4719,N_4227,N_4230);
or U4720 (N_4720,N_4023,N_4117);
xnor U4721 (N_4721,N_4427,N_4074);
or U4722 (N_4722,N_4334,N_4326);
xor U4723 (N_4723,N_4285,N_4041);
nor U4724 (N_4724,N_4217,N_4125);
xor U4725 (N_4725,N_4255,N_4198);
or U4726 (N_4726,N_4110,N_4144);
xnor U4727 (N_4727,N_4163,N_4235);
nand U4728 (N_4728,N_4208,N_4245);
nor U4729 (N_4729,N_4312,N_4482);
nor U4730 (N_4730,N_4473,N_4430);
or U4731 (N_4731,N_4136,N_4251);
nand U4732 (N_4732,N_4412,N_4260);
nor U4733 (N_4733,N_4272,N_4200);
xor U4734 (N_4734,N_4374,N_4394);
nand U4735 (N_4735,N_4092,N_4224);
nand U4736 (N_4736,N_4401,N_4405);
nor U4737 (N_4737,N_4185,N_4162);
and U4738 (N_4738,N_4127,N_4314);
and U4739 (N_4739,N_4106,N_4297);
nor U4740 (N_4740,N_4269,N_4420);
or U4741 (N_4741,N_4119,N_4408);
xor U4742 (N_4742,N_4025,N_4328);
nor U4743 (N_4743,N_4429,N_4302);
nand U4744 (N_4744,N_4301,N_4377);
xnor U4745 (N_4745,N_4064,N_4481);
or U4746 (N_4746,N_4228,N_4349);
nor U4747 (N_4747,N_4452,N_4381);
xnor U4748 (N_4748,N_4491,N_4171);
nand U4749 (N_4749,N_4172,N_4192);
nor U4750 (N_4750,N_4020,N_4183);
xor U4751 (N_4751,N_4066,N_4264);
xnor U4752 (N_4752,N_4261,N_4111);
or U4753 (N_4753,N_4483,N_4242);
nor U4754 (N_4754,N_4447,N_4067);
nand U4755 (N_4755,N_4070,N_4359);
nand U4756 (N_4756,N_4244,N_4121);
nand U4757 (N_4757,N_4068,N_4014);
nor U4758 (N_4758,N_4280,N_4480);
nand U4759 (N_4759,N_4472,N_4085);
xnor U4760 (N_4760,N_4318,N_4075);
xor U4761 (N_4761,N_4090,N_4375);
nand U4762 (N_4762,N_4080,N_4344);
nor U4763 (N_4763,N_4275,N_4306);
or U4764 (N_4764,N_4184,N_4086);
and U4765 (N_4765,N_4071,N_4141);
or U4766 (N_4766,N_4203,N_4293);
or U4767 (N_4767,N_4421,N_4020);
and U4768 (N_4768,N_4396,N_4420);
nand U4769 (N_4769,N_4231,N_4054);
xor U4770 (N_4770,N_4445,N_4311);
or U4771 (N_4771,N_4381,N_4016);
xnor U4772 (N_4772,N_4193,N_4037);
xnor U4773 (N_4773,N_4458,N_4162);
and U4774 (N_4774,N_4349,N_4321);
nand U4775 (N_4775,N_4443,N_4316);
or U4776 (N_4776,N_4301,N_4207);
and U4777 (N_4777,N_4099,N_4177);
or U4778 (N_4778,N_4117,N_4331);
xnor U4779 (N_4779,N_4342,N_4117);
nor U4780 (N_4780,N_4454,N_4173);
and U4781 (N_4781,N_4062,N_4037);
nor U4782 (N_4782,N_4197,N_4066);
or U4783 (N_4783,N_4479,N_4045);
or U4784 (N_4784,N_4484,N_4476);
xor U4785 (N_4785,N_4241,N_4447);
xnor U4786 (N_4786,N_4073,N_4387);
nand U4787 (N_4787,N_4448,N_4073);
nor U4788 (N_4788,N_4322,N_4053);
and U4789 (N_4789,N_4152,N_4490);
or U4790 (N_4790,N_4207,N_4410);
and U4791 (N_4791,N_4090,N_4454);
nor U4792 (N_4792,N_4190,N_4424);
or U4793 (N_4793,N_4109,N_4212);
xor U4794 (N_4794,N_4440,N_4406);
xnor U4795 (N_4795,N_4098,N_4282);
nand U4796 (N_4796,N_4131,N_4344);
nor U4797 (N_4797,N_4422,N_4235);
or U4798 (N_4798,N_4380,N_4119);
nor U4799 (N_4799,N_4477,N_4118);
xor U4800 (N_4800,N_4491,N_4295);
and U4801 (N_4801,N_4051,N_4154);
xnor U4802 (N_4802,N_4370,N_4240);
nor U4803 (N_4803,N_4370,N_4083);
or U4804 (N_4804,N_4213,N_4469);
or U4805 (N_4805,N_4134,N_4112);
nor U4806 (N_4806,N_4146,N_4263);
nand U4807 (N_4807,N_4121,N_4100);
nand U4808 (N_4808,N_4278,N_4174);
nand U4809 (N_4809,N_4399,N_4400);
or U4810 (N_4810,N_4421,N_4374);
and U4811 (N_4811,N_4441,N_4035);
or U4812 (N_4812,N_4015,N_4485);
or U4813 (N_4813,N_4481,N_4390);
and U4814 (N_4814,N_4107,N_4230);
xnor U4815 (N_4815,N_4481,N_4420);
and U4816 (N_4816,N_4239,N_4479);
xnor U4817 (N_4817,N_4010,N_4298);
nor U4818 (N_4818,N_4306,N_4029);
nor U4819 (N_4819,N_4468,N_4258);
xor U4820 (N_4820,N_4032,N_4265);
or U4821 (N_4821,N_4193,N_4312);
or U4822 (N_4822,N_4360,N_4093);
or U4823 (N_4823,N_4393,N_4499);
nor U4824 (N_4824,N_4098,N_4493);
xor U4825 (N_4825,N_4483,N_4354);
nand U4826 (N_4826,N_4225,N_4233);
nor U4827 (N_4827,N_4491,N_4381);
nor U4828 (N_4828,N_4485,N_4410);
xnor U4829 (N_4829,N_4141,N_4273);
nor U4830 (N_4830,N_4320,N_4387);
xnor U4831 (N_4831,N_4069,N_4193);
nor U4832 (N_4832,N_4454,N_4424);
nor U4833 (N_4833,N_4418,N_4157);
nand U4834 (N_4834,N_4195,N_4183);
xor U4835 (N_4835,N_4326,N_4376);
nand U4836 (N_4836,N_4021,N_4432);
nand U4837 (N_4837,N_4064,N_4421);
and U4838 (N_4838,N_4263,N_4362);
nor U4839 (N_4839,N_4117,N_4120);
nor U4840 (N_4840,N_4330,N_4340);
or U4841 (N_4841,N_4362,N_4377);
nor U4842 (N_4842,N_4012,N_4084);
and U4843 (N_4843,N_4337,N_4219);
nand U4844 (N_4844,N_4315,N_4454);
xnor U4845 (N_4845,N_4147,N_4141);
or U4846 (N_4846,N_4459,N_4014);
or U4847 (N_4847,N_4494,N_4388);
nand U4848 (N_4848,N_4252,N_4384);
nand U4849 (N_4849,N_4478,N_4397);
and U4850 (N_4850,N_4129,N_4139);
or U4851 (N_4851,N_4193,N_4097);
xnor U4852 (N_4852,N_4015,N_4442);
xnor U4853 (N_4853,N_4402,N_4285);
nor U4854 (N_4854,N_4005,N_4307);
or U4855 (N_4855,N_4444,N_4083);
nor U4856 (N_4856,N_4119,N_4090);
xor U4857 (N_4857,N_4151,N_4279);
and U4858 (N_4858,N_4071,N_4041);
nand U4859 (N_4859,N_4304,N_4315);
or U4860 (N_4860,N_4470,N_4403);
nand U4861 (N_4861,N_4410,N_4221);
xor U4862 (N_4862,N_4108,N_4150);
and U4863 (N_4863,N_4283,N_4019);
or U4864 (N_4864,N_4281,N_4366);
nor U4865 (N_4865,N_4342,N_4355);
nor U4866 (N_4866,N_4315,N_4215);
and U4867 (N_4867,N_4417,N_4447);
and U4868 (N_4868,N_4288,N_4365);
or U4869 (N_4869,N_4317,N_4130);
xnor U4870 (N_4870,N_4287,N_4283);
or U4871 (N_4871,N_4069,N_4466);
nor U4872 (N_4872,N_4101,N_4430);
xor U4873 (N_4873,N_4053,N_4499);
nor U4874 (N_4874,N_4106,N_4007);
xor U4875 (N_4875,N_4271,N_4424);
or U4876 (N_4876,N_4242,N_4138);
xnor U4877 (N_4877,N_4116,N_4035);
xor U4878 (N_4878,N_4444,N_4107);
and U4879 (N_4879,N_4404,N_4464);
or U4880 (N_4880,N_4335,N_4033);
and U4881 (N_4881,N_4245,N_4465);
xor U4882 (N_4882,N_4402,N_4416);
or U4883 (N_4883,N_4309,N_4377);
and U4884 (N_4884,N_4183,N_4346);
and U4885 (N_4885,N_4283,N_4127);
nand U4886 (N_4886,N_4443,N_4026);
nand U4887 (N_4887,N_4451,N_4035);
nor U4888 (N_4888,N_4420,N_4046);
xnor U4889 (N_4889,N_4475,N_4315);
nand U4890 (N_4890,N_4253,N_4426);
nand U4891 (N_4891,N_4388,N_4192);
or U4892 (N_4892,N_4005,N_4275);
or U4893 (N_4893,N_4205,N_4219);
nand U4894 (N_4894,N_4406,N_4126);
nor U4895 (N_4895,N_4160,N_4050);
nor U4896 (N_4896,N_4168,N_4320);
or U4897 (N_4897,N_4001,N_4312);
and U4898 (N_4898,N_4112,N_4121);
or U4899 (N_4899,N_4345,N_4268);
xor U4900 (N_4900,N_4363,N_4254);
xor U4901 (N_4901,N_4232,N_4125);
nand U4902 (N_4902,N_4072,N_4250);
or U4903 (N_4903,N_4038,N_4464);
nand U4904 (N_4904,N_4263,N_4441);
or U4905 (N_4905,N_4460,N_4490);
nor U4906 (N_4906,N_4495,N_4039);
and U4907 (N_4907,N_4120,N_4001);
and U4908 (N_4908,N_4408,N_4155);
and U4909 (N_4909,N_4171,N_4359);
and U4910 (N_4910,N_4461,N_4340);
nand U4911 (N_4911,N_4418,N_4212);
xnor U4912 (N_4912,N_4374,N_4165);
nand U4913 (N_4913,N_4182,N_4214);
or U4914 (N_4914,N_4380,N_4084);
xnor U4915 (N_4915,N_4359,N_4024);
or U4916 (N_4916,N_4051,N_4102);
or U4917 (N_4917,N_4278,N_4214);
xor U4918 (N_4918,N_4148,N_4170);
or U4919 (N_4919,N_4032,N_4169);
or U4920 (N_4920,N_4448,N_4437);
and U4921 (N_4921,N_4200,N_4415);
and U4922 (N_4922,N_4330,N_4199);
or U4923 (N_4923,N_4372,N_4080);
xor U4924 (N_4924,N_4088,N_4388);
xnor U4925 (N_4925,N_4052,N_4147);
or U4926 (N_4926,N_4207,N_4051);
or U4927 (N_4927,N_4023,N_4267);
and U4928 (N_4928,N_4254,N_4324);
nand U4929 (N_4929,N_4013,N_4304);
and U4930 (N_4930,N_4088,N_4231);
and U4931 (N_4931,N_4355,N_4000);
or U4932 (N_4932,N_4397,N_4153);
or U4933 (N_4933,N_4451,N_4169);
or U4934 (N_4934,N_4140,N_4151);
nand U4935 (N_4935,N_4470,N_4063);
nand U4936 (N_4936,N_4359,N_4097);
nand U4937 (N_4937,N_4340,N_4166);
xnor U4938 (N_4938,N_4016,N_4047);
xor U4939 (N_4939,N_4064,N_4343);
xnor U4940 (N_4940,N_4050,N_4266);
and U4941 (N_4941,N_4175,N_4295);
xor U4942 (N_4942,N_4184,N_4357);
or U4943 (N_4943,N_4095,N_4257);
nor U4944 (N_4944,N_4459,N_4412);
and U4945 (N_4945,N_4240,N_4419);
nor U4946 (N_4946,N_4265,N_4447);
or U4947 (N_4947,N_4423,N_4022);
xor U4948 (N_4948,N_4355,N_4036);
nand U4949 (N_4949,N_4361,N_4499);
nand U4950 (N_4950,N_4285,N_4491);
xor U4951 (N_4951,N_4362,N_4095);
or U4952 (N_4952,N_4135,N_4130);
nor U4953 (N_4953,N_4412,N_4455);
nor U4954 (N_4954,N_4345,N_4176);
nor U4955 (N_4955,N_4055,N_4312);
xor U4956 (N_4956,N_4129,N_4084);
nand U4957 (N_4957,N_4433,N_4089);
nor U4958 (N_4958,N_4212,N_4181);
and U4959 (N_4959,N_4147,N_4109);
xor U4960 (N_4960,N_4279,N_4306);
nand U4961 (N_4961,N_4125,N_4285);
and U4962 (N_4962,N_4335,N_4059);
nand U4963 (N_4963,N_4465,N_4053);
and U4964 (N_4964,N_4048,N_4015);
or U4965 (N_4965,N_4418,N_4189);
and U4966 (N_4966,N_4442,N_4296);
and U4967 (N_4967,N_4355,N_4090);
and U4968 (N_4968,N_4137,N_4104);
nand U4969 (N_4969,N_4341,N_4069);
and U4970 (N_4970,N_4365,N_4151);
or U4971 (N_4971,N_4112,N_4118);
xnor U4972 (N_4972,N_4417,N_4435);
nor U4973 (N_4973,N_4262,N_4401);
nand U4974 (N_4974,N_4260,N_4282);
nor U4975 (N_4975,N_4485,N_4391);
nor U4976 (N_4976,N_4138,N_4352);
or U4977 (N_4977,N_4025,N_4271);
nor U4978 (N_4978,N_4016,N_4253);
nor U4979 (N_4979,N_4339,N_4119);
and U4980 (N_4980,N_4426,N_4415);
or U4981 (N_4981,N_4455,N_4272);
or U4982 (N_4982,N_4464,N_4388);
nand U4983 (N_4983,N_4330,N_4089);
nor U4984 (N_4984,N_4203,N_4056);
xnor U4985 (N_4985,N_4032,N_4354);
xnor U4986 (N_4986,N_4442,N_4160);
nor U4987 (N_4987,N_4199,N_4038);
nand U4988 (N_4988,N_4058,N_4399);
or U4989 (N_4989,N_4289,N_4034);
or U4990 (N_4990,N_4070,N_4378);
and U4991 (N_4991,N_4093,N_4481);
and U4992 (N_4992,N_4382,N_4192);
or U4993 (N_4993,N_4177,N_4296);
or U4994 (N_4994,N_4321,N_4108);
xor U4995 (N_4995,N_4124,N_4164);
nand U4996 (N_4996,N_4092,N_4054);
xor U4997 (N_4997,N_4121,N_4270);
or U4998 (N_4998,N_4228,N_4135);
xnor U4999 (N_4999,N_4115,N_4157);
or U5000 (N_5000,N_4725,N_4604);
nand U5001 (N_5001,N_4614,N_4846);
nor U5002 (N_5002,N_4525,N_4896);
nand U5003 (N_5003,N_4920,N_4961);
xor U5004 (N_5004,N_4880,N_4892);
nor U5005 (N_5005,N_4541,N_4546);
or U5006 (N_5006,N_4972,N_4763);
or U5007 (N_5007,N_4963,N_4694);
nand U5008 (N_5008,N_4615,N_4752);
xnor U5009 (N_5009,N_4741,N_4794);
nand U5010 (N_5010,N_4597,N_4878);
nor U5011 (N_5011,N_4974,N_4513);
nand U5012 (N_5012,N_4904,N_4610);
or U5013 (N_5013,N_4970,N_4567);
or U5014 (N_5014,N_4825,N_4927);
nor U5015 (N_5015,N_4891,N_4737);
nand U5016 (N_5016,N_4671,N_4831);
nand U5017 (N_5017,N_4953,N_4800);
nor U5018 (N_5018,N_4555,N_4523);
nor U5019 (N_5019,N_4876,N_4673);
nand U5020 (N_5020,N_4652,N_4720);
or U5021 (N_5021,N_4564,N_4528);
or U5022 (N_5022,N_4804,N_4793);
and U5023 (N_5023,N_4550,N_4886);
or U5024 (N_5024,N_4576,N_4750);
nor U5025 (N_5025,N_4786,N_4502);
xor U5026 (N_5026,N_4785,N_4556);
nor U5027 (N_5027,N_4844,N_4653);
and U5028 (N_5028,N_4612,N_4657);
nor U5029 (N_5029,N_4894,N_4557);
nor U5030 (N_5030,N_4888,N_4634);
and U5031 (N_5031,N_4887,N_4924);
nand U5032 (N_5032,N_4828,N_4582);
and U5033 (N_5033,N_4636,N_4706);
or U5034 (N_5034,N_4635,N_4631);
xnor U5035 (N_5035,N_4868,N_4715);
and U5036 (N_5036,N_4861,N_4940);
or U5037 (N_5037,N_4664,N_4575);
nor U5038 (N_5038,N_4792,N_4625);
or U5039 (N_5039,N_4922,N_4701);
xor U5040 (N_5040,N_4526,N_4545);
nand U5041 (N_5041,N_4791,N_4761);
nand U5042 (N_5042,N_4860,N_4722);
and U5043 (N_5043,N_4820,N_4787);
nor U5044 (N_5044,N_4933,N_4911);
or U5045 (N_5045,N_4570,N_4799);
and U5046 (N_5046,N_4928,N_4930);
or U5047 (N_5047,N_4921,N_4856);
nand U5048 (N_5048,N_4757,N_4690);
nand U5049 (N_5049,N_4516,N_4695);
xnor U5050 (N_5050,N_4932,N_4938);
nor U5051 (N_5051,N_4500,N_4683);
or U5052 (N_5052,N_4986,N_4668);
xnor U5053 (N_5053,N_4889,N_4739);
and U5054 (N_5054,N_4912,N_4633);
xor U5055 (N_5055,N_4733,N_4865);
or U5056 (N_5056,N_4707,N_4562);
xor U5057 (N_5057,N_4897,N_4943);
nand U5058 (N_5058,N_4819,N_4632);
and U5059 (N_5059,N_4540,N_4817);
nand U5060 (N_5060,N_4874,N_4951);
nand U5061 (N_5061,N_4734,N_4603);
nand U5062 (N_5062,N_4906,N_4646);
and U5063 (N_5063,N_4531,N_4539);
nor U5064 (N_5064,N_4881,N_4775);
nor U5065 (N_5065,N_4867,N_4973);
xnor U5066 (N_5066,N_4997,N_4659);
or U5067 (N_5067,N_4693,N_4835);
and U5068 (N_5068,N_4747,N_4915);
and U5069 (N_5069,N_4527,N_4669);
xnor U5070 (N_5070,N_4608,N_4518);
nor U5071 (N_5071,N_4611,N_4600);
or U5072 (N_5072,N_4682,N_4858);
xnor U5073 (N_5073,N_4660,N_4758);
or U5074 (N_5074,N_4998,N_4956);
nand U5075 (N_5075,N_4935,N_4736);
and U5076 (N_5076,N_4766,N_4939);
nor U5077 (N_5077,N_4981,N_4782);
nor U5078 (N_5078,N_4853,N_4849);
and U5079 (N_5079,N_4821,N_4537);
and U5080 (N_5080,N_4764,N_4520);
nand U5081 (N_5081,N_4988,N_4812);
and U5082 (N_5082,N_4581,N_4969);
xnor U5083 (N_5083,N_4883,N_4511);
nor U5084 (N_5084,N_4929,N_4590);
nand U5085 (N_5085,N_4805,N_4514);
nor U5086 (N_5086,N_4721,N_4679);
nand U5087 (N_5087,N_4572,N_4808);
and U5088 (N_5088,N_4521,N_4620);
nand U5089 (N_5089,N_4962,N_4565);
nor U5090 (N_5090,N_4798,N_4696);
xnor U5091 (N_5091,N_4670,N_4830);
nand U5092 (N_5092,N_4640,N_4697);
and U5093 (N_5093,N_4999,N_4702);
nand U5094 (N_5094,N_4649,N_4918);
xor U5095 (N_5095,N_4993,N_4847);
xor U5096 (N_5096,N_4743,N_4688);
nand U5097 (N_5097,N_4959,N_4806);
and U5098 (N_5098,N_4810,N_4723);
nor U5099 (N_5099,N_4755,N_4579);
nand U5100 (N_5100,N_4762,N_4773);
nor U5101 (N_5101,N_4801,N_4599);
xor U5102 (N_5102,N_4913,N_4709);
or U5103 (N_5103,N_4698,N_4925);
or U5104 (N_5104,N_4729,N_4585);
nor U5105 (N_5105,N_4584,N_4829);
nor U5106 (N_5106,N_4967,N_4742);
or U5107 (N_5107,N_4765,N_4719);
nand U5108 (N_5108,N_4834,N_4983);
and U5109 (N_5109,N_4987,N_4756);
nand U5110 (N_5110,N_4833,N_4872);
xor U5111 (N_5111,N_4602,N_4795);
nand U5112 (N_5112,N_4826,N_4548);
or U5113 (N_5113,N_4838,N_4841);
or U5114 (N_5114,N_4989,N_4958);
or U5115 (N_5115,N_4917,N_4642);
and U5116 (N_5116,N_4971,N_4573);
nand U5117 (N_5117,N_4621,N_4965);
or U5118 (N_5118,N_4837,N_4661);
xnor U5119 (N_5119,N_4866,N_4945);
or U5120 (N_5120,N_4811,N_4789);
and U5121 (N_5121,N_4544,N_4542);
and U5122 (N_5122,N_4623,N_4524);
nor U5123 (N_5123,N_4593,N_4979);
or U5124 (N_5124,N_4992,N_4647);
xor U5125 (N_5125,N_4784,N_4991);
nor U5126 (N_5126,N_4882,N_4984);
nand U5127 (N_5127,N_4596,N_4666);
xnor U5128 (N_5128,N_4727,N_4717);
and U5129 (N_5129,N_4960,N_4827);
and U5130 (N_5130,N_4583,N_4704);
xnor U5131 (N_5131,N_4873,N_4580);
xnor U5132 (N_5132,N_4862,N_4508);
or U5133 (N_5133,N_4687,N_4899);
nor U5134 (N_5134,N_4517,N_4779);
nand U5135 (N_5135,N_4818,N_4654);
and U5136 (N_5136,N_4607,N_4754);
nor U5137 (N_5137,N_4947,N_4941);
xor U5138 (N_5138,N_4676,N_4898);
nor U5139 (N_5139,N_4595,N_4522);
and U5140 (N_5140,N_4885,N_4895);
and U5141 (N_5141,N_4824,N_4815);
nor U5142 (N_5142,N_4748,N_4901);
xnor U5143 (N_5143,N_4780,N_4594);
xnor U5144 (N_5144,N_4994,N_4839);
nor U5145 (N_5145,N_4678,N_4716);
nand U5146 (N_5146,N_4705,N_4535);
nor U5147 (N_5147,N_4622,N_4760);
and U5148 (N_5148,N_4955,N_4560);
or U5149 (N_5149,N_4626,N_4515);
nor U5150 (N_5150,N_4767,N_4845);
nand U5151 (N_5151,N_4547,N_4589);
nor U5152 (N_5152,N_4832,N_4504);
nand U5153 (N_5153,N_4728,N_4996);
nor U5154 (N_5154,N_4977,N_4900);
nand U5155 (N_5155,N_4549,N_4753);
and U5156 (N_5156,N_4744,N_4797);
and U5157 (N_5157,N_4648,N_4512);
or U5158 (N_5158,N_4875,N_4995);
nand U5159 (N_5159,N_4708,N_4908);
xnor U5160 (N_5160,N_4534,N_4803);
xor U5161 (N_5161,N_4561,N_4909);
and U5162 (N_5162,N_4712,N_4854);
nor U5163 (N_5163,N_4536,N_4871);
nor U5164 (N_5164,N_4617,N_4724);
xnor U5165 (N_5165,N_4822,N_4776);
nor U5166 (N_5166,N_4658,N_4667);
xnor U5167 (N_5167,N_4577,N_4650);
xnor U5168 (N_5168,N_4533,N_4843);
nand U5169 (N_5169,N_4950,N_4543);
or U5170 (N_5170,N_4796,N_4601);
xnor U5171 (N_5171,N_4745,N_4551);
and U5172 (N_5172,N_4691,N_4644);
nor U5173 (N_5173,N_4902,N_4732);
nor U5174 (N_5174,N_4884,N_4759);
and U5175 (N_5175,N_4957,N_4507);
and U5176 (N_5176,N_4916,N_4919);
and U5177 (N_5177,N_4978,N_4689);
nor U5178 (N_5178,N_4783,N_4863);
nor U5179 (N_5179,N_4770,N_4619);
or U5180 (N_5180,N_4613,N_4869);
nor U5181 (N_5181,N_4768,N_4735);
xnor U5182 (N_5182,N_4718,N_4942);
and U5183 (N_5183,N_4836,N_4692);
nand U5184 (N_5184,N_4774,N_4864);
xor U5185 (N_5185,N_4809,N_4624);
xor U5186 (N_5186,N_4529,N_4510);
nor U5187 (N_5187,N_4628,N_4591);
xor U5188 (N_5188,N_4982,N_4966);
nand U5189 (N_5189,N_4656,N_4559);
nor U5190 (N_5190,N_4588,N_4877);
nor U5191 (N_5191,N_4772,N_4711);
xor U5192 (N_5192,N_4554,N_4855);
nand U5193 (N_5193,N_4751,N_4879);
or U5194 (N_5194,N_4553,N_4907);
nand U5195 (N_5195,N_4641,N_4677);
or U5196 (N_5196,N_4569,N_4914);
and U5197 (N_5197,N_4509,N_4629);
and U5198 (N_5198,N_4639,N_4842);
and U5199 (N_5199,N_4566,N_4954);
and U5200 (N_5200,N_4616,N_4713);
nand U5201 (N_5201,N_4807,N_4730);
and U5202 (N_5202,N_4870,N_4980);
xnor U5203 (N_5203,N_4505,N_4618);
nor U5204 (N_5204,N_4592,N_4605);
xnor U5205 (N_5205,N_4681,N_4609);
xor U5206 (N_5206,N_4675,N_4655);
and U5207 (N_5207,N_4674,N_4519);
nand U5208 (N_5208,N_4574,N_4685);
nor U5209 (N_5209,N_4823,N_4643);
nand U5210 (N_5210,N_4501,N_4651);
and U5211 (N_5211,N_4964,N_4771);
xnor U5212 (N_5212,N_4663,N_4630);
nor U5213 (N_5213,N_4749,N_4563);
xnor U5214 (N_5214,N_4851,N_4703);
xnor U5215 (N_5215,N_4990,N_4627);
and U5216 (N_5216,N_4568,N_4777);
xnor U5217 (N_5217,N_4738,N_4944);
or U5218 (N_5218,N_4506,N_4975);
nand U5219 (N_5219,N_4532,N_4788);
and U5220 (N_5220,N_4680,N_4816);
xnor U5221 (N_5221,N_4700,N_4852);
xnor U5222 (N_5222,N_4905,N_4662);
xor U5223 (N_5223,N_4731,N_4586);
nor U5224 (N_5224,N_4949,N_4790);
nor U5225 (N_5225,N_4746,N_4538);
or U5226 (N_5226,N_4598,N_4769);
nand U5227 (N_5227,N_4814,N_4571);
nor U5228 (N_5228,N_4802,N_4699);
nand U5229 (N_5229,N_4859,N_4558);
xor U5230 (N_5230,N_4850,N_4684);
and U5231 (N_5231,N_4638,N_4778);
and U5232 (N_5232,N_4985,N_4931);
nor U5233 (N_5233,N_4530,N_4781);
or U5234 (N_5234,N_4893,N_4934);
nand U5235 (N_5235,N_4903,N_4968);
or U5236 (N_5236,N_4686,N_4910);
nand U5237 (N_5237,N_4740,N_4813);
or U5238 (N_5238,N_4578,N_4890);
xor U5239 (N_5239,N_4710,N_4840);
xor U5240 (N_5240,N_4606,N_4926);
nor U5241 (N_5241,N_4726,N_4857);
xnor U5242 (N_5242,N_4848,N_4503);
nand U5243 (N_5243,N_4665,N_4645);
nor U5244 (N_5244,N_4937,N_4714);
nor U5245 (N_5245,N_4948,N_4672);
xnor U5246 (N_5246,N_4587,N_4946);
xnor U5247 (N_5247,N_4552,N_4923);
xnor U5248 (N_5248,N_4952,N_4637);
nand U5249 (N_5249,N_4976,N_4936);
xor U5250 (N_5250,N_4670,N_4697);
nand U5251 (N_5251,N_4654,N_4870);
xor U5252 (N_5252,N_4913,N_4750);
nor U5253 (N_5253,N_4507,N_4879);
nor U5254 (N_5254,N_4945,N_4639);
nand U5255 (N_5255,N_4797,N_4698);
and U5256 (N_5256,N_4550,N_4568);
nand U5257 (N_5257,N_4580,N_4955);
and U5258 (N_5258,N_4533,N_4783);
and U5259 (N_5259,N_4520,N_4644);
and U5260 (N_5260,N_4761,N_4657);
or U5261 (N_5261,N_4993,N_4933);
nor U5262 (N_5262,N_4637,N_4980);
and U5263 (N_5263,N_4811,N_4986);
or U5264 (N_5264,N_4944,N_4542);
and U5265 (N_5265,N_4744,N_4743);
xnor U5266 (N_5266,N_4959,N_4874);
or U5267 (N_5267,N_4907,N_4762);
nor U5268 (N_5268,N_4885,N_4928);
or U5269 (N_5269,N_4714,N_4653);
or U5270 (N_5270,N_4906,N_4589);
nor U5271 (N_5271,N_4968,N_4856);
nand U5272 (N_5272,N_4644,N_4647);
nand U5273 (N_5273,N_4941,N_4887);
and U5274 (N_5274,N_4883,N_4502);
and U5275 (N_5275,N_4828,N_4778);
nand U5276 (N_5276,N_4506,N_4673);
nand U5277 (N_5277,N_4613,N_4514);
xor U5278 (N_5278,N_4669,N_4879);
nand U5279 (N_5279,N_4763,N_4502);
or U5280 (N_5280,N_4639,N_4660);
nor U5281 (N_5281,N_4788,N_4700);
or U5282 (N_5282,N_4562,N_4615);
nand U5283 (N_5283,N_4598,N_4588);
xnor U5284 (N_5284,N_4593,N_4846);
nand U5285 (N_5285,N_4574,N_4511);
or U5286 (N_5286,N_4883,N_4946);
nand U5287 (N_5287,N_4855,N_4851);
xnor U5288 (N_5288,N_4906,N_4574);
or U5289 (N_5289,N_4750,N_4792);
and U5290 (N_5290,N_4998,N_4958);
or U5291 (N_5291,N_4590,N_4874);
and U5292 (N_5292,N_4980,N_4687);
xnor U5293 (N_5293,N_4609,N_4827);
xnor U5294 (N_5294,N_4929,N_4918);
and U5295 (N_5295,N_4912,N_4964);
and U5296 (N_5296,N_4565,N_4682);
nand U5297 (N_5297,N_4593,N_4592);
and U5298 (N_5298,N_4525,N_4650);
xor U5299 (N_5299,N_4831,N_4700);
and U5300 (N_5300,N_4673,N_4664);
and U5301 (N_5301,N_4901,N_4554);
xnor U5302 (N_5302,N_4902,N_4556);
nand U5303 (N_5303,N_4555,N_4964);
or U5304 (N_5304,N_4684,N_4910);
nor U5305 (N_5305,N_4852,N_4998);
nor U5306 (N_5306,N_4726,N_4734);
or U5307 (N_5307,N_4878,N_4688);
or U5308 (N_5308,N_4730,N_4826);
and U5309 (N_5309,N_4655,N_4834);
nand U5310 (N_5310,N_4523,N_4924);
and U5311 (N_5311,N_4999,N_4903);
nand U5312 (N_5312,N_4540,N_4717);
or U5313 (N_5313,N_4571,N_4603);
nand U5314 (N_5314,N_4604,N_4693);
and U5315 (N_5315,N_4751,N_4679);
nand U5316 (N_5316,N_4560,N_4742);
xor U5317 (N_5317,N_4521,N_4947);
nand U5318 (N_5318,N_4619,N_4994);
nand U5319 (N_5319,N_4870,N_4962);
xnor U5320 (N_5320,N_4645,N_4973);
or U5321 (N_5321,N_4846,N_4979);
nor U5322 (N_5322,N_4713,N_4538);
nor U5323 (N_5323,N_4913,N_4760);
nor U5324 (N_5324,N_4640,N_4557);
or U5325 (N_5325,N_4950,N_4544);
nor U5326 (N_5326,N_4805,N_4923);
nand U5327 (N_5327,N_4596,N_4850);
nand U5328 (N_5328,N_4630,N_4588);
and U5329 (N_5329,N_4780,N_4936);
nor U5330 (N_5330,N_4615,N_4677);
and U5331 (N_5331,N_4947,N_4937);
xnor U5332 (N_5332,N_4820,N_4622);
xnor U5333 (N_5333,N_4848,N_4909);
or U5334 (N_5334,N_4679,N_4558);
nand U5335 (N_5335,N_4803,N_4643);
nor U5336 (N_5336,N_4678,N_4842);
nor U5337 (N_5337,N_4692,N_4764);
or U5338 (N_5338,N_4827,N_4687);
nor U5339 (N_5339,N_4965,N_4665);
nand U5340 (N_5340,N_4801,N_4586);
xor U5341 (N_5341,N_4678,N_4654);
and U5342 (N_5342,N_4971,N_4643);
and U5343 (N_5343,N_4744,N_4595);
and U5344 (N_5344,N_4688,N_4548);
and U5345 (N_5345,N_4966,N_4789);
or U5346 (N_5346,N_4578,N_4833);
and U5347 (N_5347,N_4553,N_4557);
nand U5348 (N_5348,N_4581,N_4946);
or U5349 (N_5349,N_4876,N_4943);
xnor U5350 (N_5350,N_4520,N_4816);
or U5351 (N_5351,N_4654,N_4519);
nor U5352 (N_5352,N_4757,N_4514);
or U5353 (N_5353,N_4778,N_4639);
nor U5354 (N_5354,N_4940,N_4613);
and U5355 (N_5355,N_4897,N_4693);
xnor U5356 (N_5356,N_4996,N_4739);
and U5357 (N_5357,N_4890,N_4551);
nand U5358 (N_5358,N_4621,N_4838);
or U5359 (N_5359,N_4828,N_4790);
and U5360 (N_5360,N_4762,N_4633);
or U5361 (N_5361,N_4646,N_4645);
and U5362 (N_5362,N_4768,N_4769);
and U5363 (N_5363,N_4734,N_4848);
nor U5364 (N_5364,N_4657,N_4811);
nand U5365 (N_5365,N_4824,N_4877);
or U5366 (N_5366,N_4798,N_4838);
nor U5367 (N_5367,N_4986,N_4756);
and U5368 (N_5368,N_4900,N_4633);
xnor U5369 (N_5369,N_4604,N_4510);
nand U5370 (N_5370,N_4917,N_4551);
and U5371 (N_5371,N_4581,N_4801);
xor U5372 (N_5372,N_4717,N_4925);
xnor U5373 (N_5373,N_4927,N_4871);
nor U5374 (N_5374,N_4681,N_4733);
xnor U5375 (N_5375,N_4821,N_4919);
xnor U5376 (N_5376,N_4779,N_4858);
xnor U5377 (N_5377,N_4604,N_4814);
nor U5378 (N_5378,N_4566,N_4515);
xor U5379 (N_5379,N_4544,N_4924);
nand U5380 (N_5380,N_4921,N_4598);
and U5381 (N_5381,N_4579,N_4597);
nand U5382 (N_5382,N_4626,N_4996);
nor U5383 (N_5383,N_4932,N_4554);
nand U5384 (N_5384,N_4625,N_4668);
and U5385 (N_5385,N_4656,N_4636);
xnor U5386 (N_5386,N_4532,N_4844);
xor U5387 (N_5387,N_4586,N_4912);
nand U5388 (N_5388,N_4646,N_4980);
nor U5389 (N_5389,N_4977,N_4577);
xnor U5390 (N_5390,N_4706,N_4708);
nand U5391 (N_5391,N_4584,N_4788);
xnor U5392 (N_5392,N_4949,N_4636);
xnor U5393 (N_5393,N_4916,N_4938);
xor U5394 (N_5394,N_4720,N_4867);
nor U5395 (N_5395,N_4927,N_4620);
nor U5396 (N_5396,N_4886,N_4979);
nand U5397 (N_5397,N_4612,N_4686);
nor U5398 (N_5398,N_4501,N_4505);
nand U5399 (N_5399,N_4570,N_4820);
nand U5400 (N_5400,N_4882,N_4586);
xor U5401 (N_5401,N_4634,N_4667);
nor U5402 (N_5402,N_4714,N_4581);
nand U5403 (N_5403,N_4548,N_4584);
nand U5404 (N_5404,N_4597,N_4886);
nor U5405 (N_5405,N_4648,N_4689);
xor U5406 (N_5406,N_4761,N_4803);
nor U5407 (N_5407,N_4993,N_4845);
nor U5408 (N_5408,N_4766,N_4537);
nor U5409 (N_5409,N_4632,N_4728);
nor U5410 (N_5410,N_4519,N_4880);
nand U5411 (N_5411,N_4689,N_4922);
nor U5412 (N_5412,N_4725,N_4945);
nand U5413 (N_5413,N_4606,N_4956);
nor U5414 (N_5414,N_4890,N_4641);
xnor U5415 (N_5415,N_4614,N_4991);
and U5416 (N_5416,N_4572,N_4563);
xor U5417 (N_5417,N_4780,N_4718);
nand U5418 (N_5418,N_4649,N_4809);
xnor U5419 (N_5419,N_4561,N_4791);
xor U5420 (N_5420,N_4746,N_4894);
nand U5421 (N_5421,N_4903,N_4516);
and U5422 (N_5422,N_4881,N_4611);
or U5423 (N_5423,N_4808,N_4667);
nor U5424 (N_5424,N_4884,N_4987);
and U5425 (N_5425,N_4885,N_4947);
or U5426 (N_5426,N_4565,N_4729);
xor U5427 (N_5427,N_4867,N_4634);
or U5428 (N_5428,N_4875,N_4894);
nor U5429 (N_5429,N_4566,N_4682);
nand U5430 (N_5430,N_4709,N_4722);
nor U5431 (N_5431,N_4534,N_4956);
or U5432 (N_5432,N_4610,N_4504);
xnor U5433 (N_5433,N_4814,N_4948);
or U5434 (N_5434,N_4553,N_4584);
or U5435 (N_5435,N_4782,N_4941);
nand U5436 (N_5436,N_4914,N_4506);
nor U5437 (N_5437,N_4874,N_4570);
or U5438 (N_5438,N_4815,N_4700);
and U5439 (N_5439,N_4738,N_4586);
and U5440 (N_5440,N_4982,N_4615);
xor U5441 (N_5441,N_4832,N_4627);
xnor U5442 (N_5442,N_4522,N_4833);
nor U5443 (N_5443,N_4863,N_4994);
and U5444 (N_5444,N_4580,N_4939);
nor U5445 (N_5445,N_4758,N_4954);
or U5446 (N_5446,N_4571,N_4682);
or U5447 (N_5447,N_4928,N_4549);
nor U5448 (N_5448,N_4607,N_4968);
nor U5449 (N_5449,N_4519,N_4951);
nand U5450 (N_5450,N_4949,N_4967);
xor U5451 (N_5451,N_4701,N_4852);
nor U5452 (N_5452,N_4590,N_4954);
nand U5453 (N_5453,N_4732,N_4678);
nand U5454 (N_5454,N_4796,N_4831);
nand U5455 (N_5455,N_4757,N_4915);
and U5456 (N_5456,N_4695,N_4709);
xor U5457 (N_5457,N_4661,N_4986);
nor U5458 (N_5458,N_4996,N_4740);
nand U5459 (N_5459,N_4878,N_4643);
and U5460 (N_5460,N_4970,N_4894);
nand U5461 (N_5461,N_4998,N_4899);
nor U5462 (N_5462,N_4995,N_4727);
and U5463 (N_5463,N_4715,N_4536);
or U5464 (N_5464,N_4708,N_4964);
or U5465 (N_5465,N_4938,N_4689);
and U5466 (N_5466,N_4602,N_4869);
nand U5467 (N_5467,N_4838,N_4998);
or U5468 (N_5468,N_4731,N_4621);
or U5469 (N_5469,N_4755,N_4563);
nand U5470 (N_5470,N_4900,N_4903);
xnor U5471 (N_5471,N_4502,N_4940);
or U5472 (N_5472,N_4972,N_4533);
nand U5473 (N_5473,N_4910,N_4536);
nor U5474 (N_5474,N_4660,N_4931);
nor U5475 (N_5475,N_4825,N_4633);
and U5476 (N_5476,N_4782,N_4809);
nor U5477 (N_5477,N_4852,N_4552);
or U5478 (N_5478,N_4908,N_4882);
or U5479 (N_5479,N_4649,N_4801);
and U5480 (N_5480,N_4623,N_4870);
xor U5481 (N_5481,N_4875,N_4738);
nand U5482 (N_5482,N_4626,N_4951);
xor U5483 (N_5483,N_4879,N_4941);
and U5484 (N_5484,N_4590,N_4936);
nand U5485 (N_5485,N_4586,N_4780);
xor U5486 (N_5486,N_4783,N_4853);
nor U5487 (N_5487,N_4754,N_4609);
xor U5488 (N_5488,N_4668,N_4857);
or U5489 (N_5489,N_4864,N_4879);
or U5490 (N_5490,N_4651,N_4692);
and U5491 (N_5491,N_4649,N_4745);
nand U5492 (N_5492,N_4903,N_4895);
or U5493 (N_5493,N_4564,N_4718);
and U5494 (N_5494,N_4816,N_4566);
or U5495 (N_5495,N_4516,N_4559);
and U5496 (N_5496,N_4694,N_4921);
nand U5497 (N_5497,N_4961,N_4647);
xnor U5498 (N_5498,N_4942,N_4970);
and U5499 (N_5499,N_4824,N_4902);
xnor U5500 (N_5500,N_5189,N_5246);
nand U5501 (N_5501,N_5163,N_5295);
nor U5502 (N_5502,N_5289,N_5329);
nand U5503 (N_5503,N_5167,N_5300);
or U5504 (N_5504,N_5335,N_5127);
or U5505 (N_5505,N_5409,N_5022);
and U5506 (N_5506,N_5312,N_5252);
nand U5507 (N_5507,N_5370,N_5260);
xor U5508 (N_5508,N_5058,N_5109);
nor U5509 (N_5509,N_5294,N_5489);
and U5510 (N_5510,N_5180,N_5073);
or U5511 (N_5511,N_5057,N_5244);
and U5512 (N_5512,N_5385,N_5288);
xnor U5513 (N_5513,N_5028,N_5471);
nand U5514 (N_5514,N_5496,N_5110);
or U5515 (N_5515,N_5266,N_5334);
nor U5516 (N_5516,N_5021,N_5147);
xor U5517 (N_5517,N_5078,N_5197);
nor U5518 (N_5518,N_5133,N_5041);
nor U5519 (N_5519,N_5187,N_5221);
and U5520 (N_5520,N_5213,N_5402);
nand U5521 (N_5521,N_5411,N_5045);
nand U5522 (N_5522,N_5201,N_5414);
or U5523 (N_5523,N_5333,N_5004);
and U5524 (N_5524,N_5378,N_5023);
or U5525 (N_5525,N_5410,N_5362);
or U5526 (N_5526,N_5337,N_5426);
and U5527 (N_5527,N_5444,N_5292);
nand U5528 (N_5528,N_5322,N_5148);
and U5529 (N_5529,N_5231,N_5276);
xnor U5530 (N_5530,N_5157,N_5065);
or U5531 (N_5531,N_5238,N_5119);
xor U5532 (N_5532,N_5382,N_5264);
nand U5533 (N_5533,N_5481,N_5139);
xor U5534 (N_5534,N_5018,N_5176);
nor U5535 (N_5535,N_5227,N_5394);
nor U5536 (N_5536,N_5474,N_5466);
or U5537 (N_5537,N_5226,N_5166);
and U5538 (N_5538,N_5283,N_5388);
nor U5539 (N_5539,N_5425,N_5241);
xor U5540 (N_5540,N_5458,N_5026);
nor U5541 (N_5541,N_5239,N_5164);
xnor U5542 (N_5542,N_5342,N_5060);
and U5543 (N_5543,N_5107,N_5014);
nor U5544 (N_5544,N_5150,N_5493);
and U5545 (N_5545,N_5171,N_5095);
and U5546 (N_5546,N_5429,N_5498);
nand U5547 (N_5547,N_5223,N_5096);
xor U5548 (N_5548,N_5233,N_5416);
and U5549 (N_5549,N_5042,N_5428);
and U5550 (N_5550,N_5430,N_5450);
nor U5551 (N_5551,N_5325,N_5181);
and U5552 (N_5552,N_5105,N_5358);
nor U5553 (N_5553,N_5206,N_5256);
or U5554 (N_5554,N_5359,N_5070);
nor U5555 (N_5555,N_5321,N_5236);
xor U5556 (N_5556,N_5437,N_5002);
xnor U5557 (N_5557,N_5054,N_5379);
nor U5558 (N_5558,N_5056,N_5237);
nor U5559 (N_5559,N_5027,N_5199);
nand U5560 (N_5560,N_5268,N_5030);
nor U5561 (N_5561,N_5116,N_5093);
or U5562 (N_5562,N_5316,N_5285);
nor U5563 (N_5563,N_5254,N_5081);
or U5564 (N_5564,N_5098,N_5467);
or U5565 (N_5565,N_5305,N_5432);
nor U5566 (N_5566,N_5203,N_5219);
nand U5567 (N_5567,N_5470,N_5019);
nor U5568 (N_5568,N_5386,N_5101);
nor U5569 (N_5569,N_5029,N_5357);
or U5570 (N_5570,N_5247,N_5468);
nand U5571 (N_5571,N_5330,N_5209);
xnor U5572 (N_5572,N_5345,N_5068);
xor U5573 (N_5573,N_5207,N_5082);
nor U5574 (N_5574,N_5061,N_5265);
xor U5575 (N_5575,N_5353,N_5297);
and U5576 (N_5576,N_5348,N_5145);
nor U5577 (N_5577,N_5000,N_5490);
nand U5578 (N_5578,N_5215,N_5461);
nor U5579 (N_5579,N_5383,N_5132);
nand U5580 (N_5580,N_5311,N_5212);
nand U5581 (N_5581,N_5195,N_5158);
nand U5582 (N_5582,N_5140,N_5261);
nor U5583 (N_5583,N_5415,N_5459);
nand U5584 (N_5584,N_5007,N_5462);
and U5585 (N_5585,N_5012,N_5317);
nand U5586 (N_5586,N_5135,N_5438);
nand U5587 (N_5587,N_5210,N_5074);
or U5588 (N_5588,N_5401,N_5480);
nand U5589 (N_5589,N_5040,N_5131);
nand U5590 (N_5590,N_5282,N_5198);
or U5591 (N_5591,N_5126,N_5473);
nand U5592 (N_5592,N_5419,N_5306);
nand U5593 (N_5593,N_5124,N_5435);
nor U5594 (N_5594,N_5138,N_5063);
xnor U5595 (N_5595,N_5043,N_5072);
nor U5596 (N_5596,N_5304,N_5249);
nand U5597 (N_5597,N_5303,N_5454);
nor U5598 (N_5598,N_5491,N_5130);
nand U5599 (N_5599,N_5477,N_5153);
nand U5600 (N_5600,N_5134,N_5332);
nand U5601 (N_5601,N_5024,N_5296);
or U5602 (N_5602,N_5299,N_5038);
nand U5603 (N_5603,N_5235,N_5214);
and U5604 (N_5604,N_5344,N_5286);
or U5605 (N_5605,N_5472,N_5412);
nor U5606 (N_5606,N_5165,N_5381);
and U5607 (N_5607,N_5400,N_5397);
or U5608 (N_5608,N_5418,N_5059);
nor U5609 (N_5609,N_5087,N_5088);
xnor U5610 (N_5610,N_5447,N_5141);
nor U5611 (N_5611,N_5032,N_5262);
xnor U5612 (N_5612,N_5486,N_5441);
or U5613 (N_5613,N_5273,N_5280);
xnor U5614 (N_5614,N_5281,N_5044);
and U5615 (N_5615,N_5159,N_5177);
nand U5616 (N_5616,N_5067,N_5174);
or U5617 (N_5617,N_5373,N_5062);
nand U5618 (N_5618,N_5035,N_5320);
nor U5619 (N_5619,N_5403,N_5192);
xnor U5620 (N_5620,N_5017,N_5079);
xor U5621 (N_5621,N_5125,N_5089);
xor U5622 (N_5622,N_5046,N_5049);
nand U5623 (N_5623,N_5390,N_5271);
xor U5624 (N_5624,N_5031,N_5050);
or U5625 (N_5625,N_5250,N_5008);
or U5626 (N_5626,N_5376,N_5055);
nor U5627 (N_5627,N_5279,N_5443);
nor U5628 (N_5628,N_5298,N_5278);
or U5629 (N_5629,N_5104,N_5393);
nand U5630 (N_5630,N_5431,N_5439);
and U5631 (N_5631,N_5338,N_5003);
nand U5632 (N_5632,N_5451,N_5277);
or U5633 (N_5633,N_5367,N_5423);
and U5634 (N_5634,N_5188,N_5071);
nor U5635 (N_5635,N_5408,N_5118);
and U5636 (N_5636,N_5113,N_5488);
or U5637 (N_5637,N_5083,N_5160);
or U5638 (N_5638,N_5396,N_5398);
nor U5639 (N_5639,N_5085,N_5413);
nand U5640 (N_5640,N_5048,N_5037);
or U5641 (N_5641,N_5284,N_5346);
nand U5642 (N_5642,N_5064,N_5010);
and U5643 (N_5643,N_5094,N_5034);
nand U5644 (N_5644,N_5336,N_5436);
nand U5645 (N_5645,N_5205,N_5009);
and U5646 (N_5646,N_5449,N_5421);
or U5647 (N_5647,N_5374,N_5090);
nand U5648 (N_5648,N_5066,N_5162);
nand U5649 (N_5649,N_5255,N_5169);
xnor U5650 (N_5650,N_5194,N_5361);
nand U5651 (N_5651,N_5420,N_5293);
and U5652 (N_5652,N_5076,N_5220);
and U5653 (N_5653,N_5106,N_5445);
and U5654 (N_5654,N_5455,N_5091);
xor U5655 (N_5655,N_5355,N_5483);
and U5656 (N_5656,N_5154,N_5456);
or U5657 (N_5657,N_5216,N_5387);
nor U5658 (N_5658,N_5146,N_5230);
nand U5659 (N_5659,N_5417,N_5123);
xor U5660 (N_5660,N_5463,N_5331);
and U5661 (N_5661,N_5446,N_5352);
nand U5662 (N_5662,N_5240,N_5097);
or U5663 (N_5663,N_5077,N_5270);
nand U5664 (N_5664,N_5075,N_5399);
and U5665 (N_5665,N_5313,N_5407);
xor U5666 (N_5666,N_5120,N_5122);
nand U5667 (N_5667,N_5005,N_5433);
xor U5668 (N_5668,N_5354,N_5340);
nor U5669 (N_5669,N_5084,N_5051);
or U5670 (N_5670,N_5404,N_5469);
or U5671 (N_5671,N_5185,N_5368);
or U5672 (N_5672,N_5341,N_5365);
nand U5673 (N_5673,N_5327,N_5324);
and U5674 (N_5674,N_5484,N_5190);
or U5675 (N_5675,N_5291,N_5172);
or U5676 (N_5676,N_5155,N_5248);
nand U5677 (N_5677,N_5015,N_5170);
or U5678 (N_5678,N_5224,N_5251);
or U5679 (N_5679,N_5100,N_5350);
nand U5680 (N_5680,N_5482,N_5080);
nor U5681 (N_5681,N_5323,N_5395);
nand U5682 (N_5682,N_5319,N_5360);
xnor U5683 (N_5683,N_5476,N_5364);
xor U5684 (N_5684,N_5103,N_5011);
xnor U5685 (N_5685,N_5151,N_5302);
and U5686 (N_5686,N_5274,N_5121);
nor U5687 (N_5687,N_5128,N_5479);
xnor U5688 (N_5688,N_5161,N_5242);
xor U5689 (N_5689,N_5405,N_5202);
or U5690 (N_5690,N_5228,N_5328);
xnor U5691 (N_5691,N_5112,N_5092);
xor U5692 (N_5692,N_5307,N_5310);
or U5693 (N_5693,N_5314,N_5392);
nand U5694 (N_5694,N_5052,N_5384);
or U5695 (N_5695,N_5391,N_5108);
xnor U5696 (N_5696,N_5152,N_5309);
xor U5697 (N_5697,N_5406,N_5200);
and U5698 (N_5698,N_5225,N_5001);
nand U5699 (N_5699,N_5326,N_5442);
xor U5700 (N_5700,N_5253,N_5184);
and U5701 (N_5701,N_5142,N_5427);
nor U5702 (N_5702,N_5053,N_5229);
nor U5703 (N_5703,N_5372,N_5149);
and U5704 (N_5704,N_5269,N_5315);
or U5705 (N_5705,N_5478,N_5245);
nor U5706 (N_5706,N_5186,N_5308);
or U5707 (N_5707,N_5485,N_5290);
and U5708 (N_5708,N_5424,N_5086);
nor U5709 (N_5709,N_5033,N_5179);
xor U5710 (N_5710,N_5452,N_5193);
nand U5711 (N_5711,N_5117,N_5006);
and U5712 (N_5712,N_5339,N_5196);
and U5713 (N_5713,N_5222,N_5183);
and U5714 (N_5714,N_5143,N_5137);
nor U5715 (N_5715,N_5475,N_5272);
or U5716 (N_5716,N_5375,N_5448);
nand U5717 (N_5717,N_5243,N_5102);
nor U5718 (N_5718,N_5173,N_5208);
nand U5719 (N_5719,N_5275,N_5389);
or U5720 (N_5720,N_5232,N_5366);
xnor U5721 (N_5721,N_5234,N_5175);
nand U5722 (N_5722,N_5460,N_5039);
nand U5723 (N_5723,N_5434,N_5347);
nand U5724 (N_5724,N_5144,N_5259);
nand U5725 (N_5725,N_5016,N_5069);
xor U5726 (N_5726,N_5495,N_5218);
nor U5727 (N_5727,N_5440,N_5047);
xor U5728 (N_5728,N_5422,N_5351);
and U5729 (N_5729,N_5464,N_5494);
nor U5730 (N_5730,N_5497,N_5114);
nand U5731 (N_5731,N_5267,N_5465);
nand U5732 (N_5732,N_5115,N_5287);
and U5733 (N_5733,N_5380,N_5263);
nor U5734 (N_5734,N_5371,N_5168);
xnor U5735 (N_5735,N_5217,N_5111);
nand U5736 (N_5736,N_5025,N_5363);
nor U5737 (N_5737,N_5258,N_5036);
or U5738 (N_5738,N_5369,N_5457);
and U5739 (N_5739,N_5156,N_5487);
nand U5740 (N_5740,N_5013,N_5178);
or U5741 (N_5741,N_5211,N_5257);
or U5742 (N_5742,N_5129,N_5301);
nand U5743 (N_5743,N_5343,N_5453);
nor U5744 (N_5744,N_5191,N_5182);
nor U5745 (N_5745,N_5499,N_5318);
nand U5746 (N_5746,N_5020,N_5356);
nand U5747 (N_5747,N_5136,N_5204);
xor U5748 (N_5748,N_5349,N_5377);
nor U5749 (N_5749,N_5099,N_5492);
nor U5750 (N_5750,N_5290,N_5051);
nor U5751 (N_5751,N_5205,N_5057);
nor U5752 (N_5752,N_5119,N_5421);
xor U5753 (N_5753,N_5493,N_5251);
nand U5754 (N_5754,N_5207,N_5193);
or U5755 (N_5755,N_5020,N_5249);
and U5756 (N_5756,N_5091,N_5247);
and U5757 (N_5757,N_5462,N_5435);
and U5758 (N_5758,N_5079,N_5250);
or U5759 (N_5759,N_5354,N_5465);
or U5760 (N_5760,N_5382,N_5116);
or U5761 (N_5761,N_5165,N_5322);
nand U5762 (N_5762,N_5055,N_5113);
nor U5763 (N_5763,N_5375,N_5398);
or U5764 (N_5764,N_5302,N_5345);
or U5765 (N_5765,N_5373,N_5351);
and U5766 (N_5766,N_5235,N_5464);
nand U5767 (N_5767,N_5094,N_5262);
nor U5768 (N_5768,N_5352,N_5304);
nor U5769 (N_5769,N_5290,N_5120);
xnor U5770 (N_5770,N_5378,N_5485);
nand U5771 (N_5771,N_5200,N_5124);
nand U5772 (N_5772,N_5276,N_5474);
nor U5773 (N_5773,N_5321,N_5078);
or U5774 (N_5774,N_5457,N_5437);
or U5775 (N_5775,N_5278,N_5414);
and U5776 (N_5776,N_5060,N_5120);
and U5777 (N_5777,N_5205,N_5338);
nor U5778 (N_5778,N_5079,N_5464);
nand U5779 (N_5779,N_5423,N_5128);
nor U5780 (N_5780,N_5097,N_5269);
and U5781 (N_5781,N_5195,N_5388);
and U5782 (N_5782,N_5235,N_5189);
nand U5783 (N_5783,N_5050,N_5450);
and U5784 (N_5784,N_5022,N_5356);
nor U5785 (N_5785,N_5354,N_5422);
xnor U5786 (N_5786,N_5369,N_5140);
and U5787 (N_5787,N_5478,N_5049);
or U5788 (N_5788,N_5307,N_5007);
nor U5789 (N_5789,N_5276,N_5385);
or U5790 (N_5790,N_5063,N_5432);
nor U5791 (N_5791,N_5436,N_5104);
nor U5792 (N_5792,N_5311,N_5494);
and U5793 (N_5793,N_5353,N_5361);
xor U5794 (N_5794,N_5419,N_5128);
nand U5795 (N_5795,N_5452,N_5484);
xor U5796 (N_5796,N_5067,N_5150);
xnor U5797 (N_5797,N_5216,N_5183);
or U5798 (N_5798,N_5315,N_5010);
xor U5799 (N_5799,N_5342,N_5326);
nand U5800 (N_5800,N_5137,N_5356);
and U5801 (N_5801,N_5077,N_5415);
nand U5802 (N_5802,N_5212,N_5047);
or U5803 (N_5803,N_5283,N_5362);
or U5804 (N_5804,N_5484,N_5380);
nor U5805 (N_5805,N_5116,N_5385);
nand U5806 (N_5806,N_5179,N_5326);
and U5807 (N_5807,N_5200,N_5381);
nor U5808 (N_5808,N_5282,N_5363);
xnor U5809 (N_5809,N_5458,N_5378);
nor U5810 (N_5810,N_5382,N_5006);
or U5811 (N_5811,N_5375,N_5407);
and U5812 (N_5812,N_5220,N_5245);
or U5813 (N_5813,N_5357,N_5208);
or U5814 (N_5814,N_5177,N_5380);
nand U5815 (N_5815,N_5166,N_5239);
xnor U5816 (N_5816,N_5023,N_5213);
xnor U5817 (N_5817,N_5356,N_5443);
and U5818 (N_5818,N_5185,N_5147);
nor U5819 (N_5819,N_5436,N_5406);
nor U5820 (N_5820,N_5391,N_5065);
nor U5821 (N_5821,N_5377,N_5374);
xnor U5822 (N_5822,N_5217,N_5069);
xnor U5823 (N_5823,N_5290,N_5270);
xor U5824 (N_5824,N_5196,N_5298);
xnor U5825 (N_5825,N_5378,N_5207);
nor U5826 (N_5826,N_5129,N_5299);
nor U5827 (N_5827,N_5434,N_5460);
or U5828 (N_5828,N_5356,N_5415);
and U5829 (N_5829,N_5214,N_5367);
xnor U5830 (N_5830,N_5208,N_5175);
or U5831 (N_5831,N_5493,N_5453);
and U5832 (N_5832,N_5489,N_5462);
or U5833 (N_5833,N_5465,N_5066);
and U5834 (N_5834,N_5313,N_5491);
and U5835 (N_5835,N_5125,N_5301);
xnor U5836 (N_5836,N_5209,N_5364);
nand U5837 (N_5837,N_5281,N_5413);
nand U5838 (N_5838,N_5091,N_5274);
xnor U5839 (N_5839,N_5463,N_5468);
xnor U5840 (N_5840,N_5137,N_5470);
and U5841 (N_5841,N_5265,N_5302);
nand U5842 (N_5842,N_5092,N_5447);
nor U5843 (N_5843,N_5267,N_5446);
nand U5844 (N_5844,N_5322,N_5013);
or U5845 (N_5845,N_5364,N_5235);
and U5846 (N_5846,N_5404,N_5044);
nand U5847 (N_5847,N_5474,N_5236);
nand U5848 (N_5848,N_5161,N_5476);
xor U5849 (N_5849,N_5439,N_5321);
nor U5850 (N_5850,N_5351,N_5017);
xor U5851 (N_5851,N_5488,N_5485);
xnor U5852 (N_5852,N_5189,N_5360);
or U5853 (N_5853,N_5223,N_5286);
nand U5854 (N_5854,N_5185,N_5217);
nor U5855 (N_5855,N_5363,N_5449);
nor U5856 (N_5856,N_5305,N_5060);
nand U5857 (N_5857,N_5302,N_5395);
or U5858 (N_5858,N_5248,N_5436);
nand U5859 (N_5859,N_5165,N_5255);
or U5860 (N_5860,N_5155,N_5302);
or U5861 (N_5861,N_5388,N_5037);
nand U5862 (N_5862,N_5328,N_5416);
xor U5863 (N_5863,N_5186,N_5409);
nand U5864 (N_5864,N_5490,N_5454);
or U5865 (N_5865,N_5158,N_5474);
or U5866 (N_5866,N_5347,N_5295);
xnor U5867 (N_5867,N_5030,N_5214);
nor U5868 (N_5868,N_5210,N_5241);
and U5869 (N_5869,N_5088,N_5182);
xor U5870 (N_5870,N_5048,N_5312);
xor U5871 (N_5871,N_5499,N_5398);
or U5872 (N_5872,N_5203,N_5200);
or U5873 (N_5873,N_5196,N_5167);
nor U5874 (N_5874,N_5118,N_5204);
nor U5875 (N_5875,N_5416,N_5107);
nand U5876 (N_5876,N_5413,N_5317);
nor U5877 (N_5877,N_5015,N_5346);
nand U5878 (N_5878,N_5315,N_5374);
and U5879 (N_5879,N_5286,N_5205);
and U5880 (N_5880,N_5130,N_5076);
and U5881 (N_5881,N_5411,N_5249);
nor U5882 (N_5882,N_5023,N_5148);
or U5883 (N_5883,N_5072,N_5279);
xor U5884 (N_5884,N_5101,N_5131);
or U5885 (N_5885,N_5330,N_5438);
nor U5886 (N_5886,N_5007,N_5492);
xnor U5887 (N_5887,N_5116,N_5468);
and U5888 (N_5888,N_5398,N_5343);
or U5889 (N_5889,N_5171,N_5266);
or U5890 (N_5890,N_5065,N_5244);
nor U5891 (N_5891,N_5207,N_5418);
nor U5892 (N_5892,N_5268,N_5356);
nor U5893 (N_5893,N_5368,N_5465);
or U5894 (N_5894,N_5140,N_5367);
or U5895 (N_5895,N_5195,N_5367);
nand U5896 (N_5896,N_5478,N_5212);
xor U5897 (N_5897,N_5161,N_5001);
xor U5898 (N_5898,N_5235,N_5023);
or U5899 (N_5899,N_5250,N_5253);
nor U5900 (N_5900,N_5043,N_5000);
nand U5901 (N_5901,N_5278,N_5188);
or U5902 (N_5902,N_5318,N_5012);
nor U5903 (N_5903,N_5188,N_5394);
or U5904 (N_5904,N_5311,N_5114);
nand U5905 (N_5905,N_5071,N_5326);
or U5906 (N_5906,N_5495,N_5030);
or U5907 (N_5907,N_5375,N_5489);
or U5908 (N_5908,N_5498,N_5479);
nor U5909 (N_5909,N_5453,N_5274);
or U5910 (N_5910,N_5315,N_5038);
nor U5911 (N_5911,N_5297,N_5338);
or U5912 (N_5912,N_5211,N_5127);
nor U5913 (N_5913,N_5070,N_5272);
nor U5914 (N_5914,N_5084,N_5239);
nor U5915 (N_5915,N_5435,N_5148);
and U5916 (N_5916,N_5247,N_5275);
xor U5917 (N_5917,N_5450,N_5211);
nand U5918 (N_5918,N_5045,N_5375);
or U5919 (N_5919,N_5248,N_5071);
and U5920 (N_5920,N_5245,N_5271);
xor U5921 (N_5921,N_5095,N_5253);
nor U5922 (N_5922,N_5269,N_5107);
nand U5923 (N_5923,N_5219,N_5227);
xnor U5924 (N_5924,N_5312,N_5245);
and U5925 (N_5925,N_5342,N_5166);
and U5926 (N_5926,N_5109,N_5369);
xor U5927 (N_5927,N_5073,N_5484);
xor U5928 (N_5928,N_5098,N_5195);
nor U5929 (N_5929,N_5168,N_5217);
nor U5930 (N_5930,N_5196,N_5192);
and U5931 (N_5931,N_5248,N_5305);
nand U5932 (N_5932,N_5255,N_5454);
nand U5933 (N_5933,N_5151,N_5089);
and U5934 (N_5934,N_5046,N_5312);
and U5935 (N_5935,N_5014,N_5332);
or U5936 (N_5936,N_5162,N_5253);
xor U5937 (N_5937,N_5007,N_5430);
or U5938 (N_5938,N_5117,N_5421);
or U5939 (N_5939,N_5232,N_5476);
and U5940 (N_5940,N_5169,N_5340);
nand U5941 (N_5941,N_5088,N_5211);
and U5942 (N_5942,N_5302,N_5217);
and U5943 (N_5943,N_5487,N_5352);
xnor U5944 (N_5944,N_5298,N_5233);
nor U5945 (N_5945,N_5063,N_5319);
xor U5946 (N_5946,N_5374,N_5061);
nor U5947 (N_5947,N_5038,N_5185);
or U5948 (N_5948,N_5060,N_5076);
and U5949 (N_5949,N_5391,N_5409);
and U5950 (N_5950,N_5286,N_5494);
xnor U5951 (N_5951,N_5229,N_5351);
xor U5952 (N_5952,N_5497,N_5043);
xor U5953 (N_5953,N_5410,N_5088);
nand U5954 (N_5954,N_5082,N_5117);
nor U5955 (N_5955,N_5351,N_5468);
and U5956 (N_5956,N_5209,N_5387);
or U5957 (N_5957,N_5446,N_5102);
nand U5958 (N_5958,N_5128,N_5202);
nor U5959 (N_5959,N_5287,N_5110);
xor U5960 (N_5960,N_5001,N_5048);
and U5961 (N_5961,N_5073,N_5026);
and U5962 (N_5962,N_5021,N_5023);
nor U5963 (N_5963,N_5381,N_5128);
and U5964 (N_5964,N_5412,N_5306);
or U5965 (N_5965,N_5039,N_5287);
or U5966 (N_5966,N_5494,N_5017);
nand U5967 (N_5967,N_5436,N_5021);
or U5968 (N_5968,N_5210,N_5300);
xor U5969 (N_5969,N_5232,N_5496);
nand U5970 (N_5970,N_5276,N_5255);
or U5971 (N_5971,N_5247,N_5225);
or U5972 (N_5972,N_5408,N_5095);
and U5973 (N_5973,N_5295,N_5142);
nor U5974 (N_5974,N_5251,N_5278);
nand U5975 (N_5975,N_5097,N_5162);
and U5976 (N_5976,N_5470,N_5261);
nor U5977 (N_5977,N_5487,N_5016);
nand U5978 (N_5978,N_5017,N_5244);
and U5979 (N_5979,N_5421,N_5050);
and U5980 (N_5980,N_5381,N_5153);
nor U5981 (N_5981,N_5440,N_5108);
nand U5982 (N_5982,N_5368,N_5019);
xor U5983 (N_5983,N_5365,N_5145);
or U5984 (N_5984,N_5047,N_5330);
xnor U5985 (N_5985,N_5051,N_5082);
nor U5986 (N_5986,N_5052,N_5477);
and U5987 (N_5987,N_5352,N_5193);
nand U5988 (N_5988,N_5173,N_5234);
and U5989 (N_5989,N_5372,N_5035);
nand U5990 (N_5990,N_5223,N_5161);
or U5991 (N_5991,N_5102,N_5348);
nand U5992 (N_5992,N_5426,N_5057);
nand U5993 (N_5993,N_5004,N_5146);
or U5994 (N_5994,N_5461,N_5171);
and U5995 (N_5995,N_5207,N_5329);
and U5996 (N_5996,N_5303,N_5294);
nand U5997 (N_5997,N_5498,N_5108);
xnor U5998 (N_5998,N_5294,N_5477);
nand U5999 (N_5999,N_5041,N_5179);
xor U6000 (N_6000,N_5874,N_5506);
xor U6001 (N_6001,N_5784,N_5601);
or U6002 (N_6002,N_5642,N_5779);
xor U6003 (N_6003,N_5804,N_5820);
xor U6004 (N_6004,N_5731,N_5600);
nor U6005 (N_6005,N_5537,N_5615);
nand U6006 (N_6006,N_5596,N_5764);
or U6007 (N_6007,N_5751,N_5792);
nor U6008 (N_6008,N_5554,N_5602);
xnor U6009 (N_6009,N_5721,N_5909);
or U6010 (N_6010,N_5933,N_5884);
xor U6011 (N_6011,N_5746,N_5844);
or U6012 (N_6012,N_5572,N_5611);
nand U6013 (N_6013,N_5523,N_5743);
nor U6014 (N_6014,N_5950,N_5802);
and U6015 (N_6015,N_5949,N_5952);
nor U6016 (N_6016,N_5684,N_5795);
xor U6017 (N_6017,N_5593,N_5984);
xor U6018 (N_6018,N_5906,N_5893);
or U6019 (N_6019,N_5843,N_5740);
nor U6020 (N_6020,N_5834,N_5819);
or U6021 (N_6021,N_5534,N_5903);
nand U6022 (N_6022,N_5667,N_5693);
nor U6023 (N_6023,N_5570,N_5846);
nand U6024 (N_6024,N_5956,N_5787);
xor U6025 (N_6025,N_5977,N_5877);
xor U6026 (N_6026,N_5864,N_5586);
nor U6027 (N_6027,N_5962,N_5747);
nand U6028 (N_6028,N_5744,N_5953);
or U6029 (N_6029,N_5649,N_5697);
and U6030 (N_6030,N_5641,N_5979);
xnor U6031 (N_6031,N_5808,N_5917);
or U6032 (N_6032,N_5587,N_5821);
nor U6033 (N_6033,N_5723,N_5910);
nand U6034 (N_6034,N_5876,N_5741);
xnor U6035 (N_6035,N_5826,N_5734);
or U6036 (N_6036,N_5509,N_5553);
nand U6037 (N_6037,N_5813,N_5840);
and U6038 (N_6038,N_5612,N_5915);
nand U6039 (N_6039,N_5580,N_5563);
or U6040 (N_6040,N_5644,N_5632);
and U6041 (N_6041,N_5951,N_5797);
or U6042 (N_6042,N_5637,N_5980);
nand U6043 (N_6043,N_5898,N_5573);
nand U6044 (N_6044,N_5860,N_5548);
or U6045 (N_6045,N_5786,N_5881);
xor U6046 (N_6046,N_5681,N_5560);
nor U6047 (N_6047,N_5664,N_5790);
or U6048 (N_6048,N_5619,N_5945);
and U6049 (N_6049,N_5545,N_5831);
and U6050 (N_6050,N_5916,N_5712);
nand U6051 (N_6051,N_5861,N_5995);
nor U6052 (N_6052,N_5647,N_5827);
or U6053 (N_6053,N_5970,N_5608);
and U6054 (N_6054,N_5630,N_5558);
or U6055 (N_6055,N_5807,N_5661);
nand U6056 (N_6056,N_5568,N_5845);
nand U6057 (N_6057,N_5891,N_5908);
nor U6058 (N_6058,N_5607,N_5948);
or U6059 (N_6059,N_5894,N_5668);
or U6060 (N_6060,N_5559,N_5606);
nor U6061 (N_6061,N_5530,N_5782);
nor U6062 (N_6062,N_5849,N_5789);
and U6063 (N_6063,N_5886,N_5870);
or U6064 (N_6064,N_5645,N_5550);
and U6065 (N_6065,N_5708,N_5718);
or U6066 (N_6066,N_5830,N_5946);
or U6067 (N_6067,N_5540,N_5928);
nand U6068 (N_6068,N_5699,N_5932);
nand U6069 (N_6069,N_5502,N_5942);
and U6070 (N_6070,N_5594,N_5522);
xnor U6071 (N_6071,N_5643,N_5590);
nor U6072 (N_6072,N_5837,N_5521);
or U6073 (N_6073,N_5672,N_5887);
xnor U6074 (N_6074,N_5758,N_5666);
xor U6075 (N_6075,N_5639,N_5713);
nand U6076 (N_6076,N_5981,N_5996);
or U6077 (N_6077,N_5679,N_5759);
and U6078 (N_6078,N_5926,N_5774);
and U6079 (N_6079,N_5687,N_5833);
and U6080 (N_6080,N_5745,N_5581);
or U6081 (N_6081,N_5508,N_5655);
or U6082 (N_6082,N_5756,N_5503);
nor U6083 (N_6083,N_5957,N_5685);
or U6084 (N_6084,N_5654,N_5993);
nand U6085 (N_6085,N_5754,N_5850);
nor U6086 (N_6086,N_5562,N_5960);
and U6087 (N_6087,N_5737,N_5766);
or U6088 (N_6088,N_5662,N_5597);
nand U6089 (N_6089,N_5866,N_5825);
and U6090 (N_6090,N_5565,N_5800);
or U6091 (N_6091,N_5769,N_5620);
nand U6092 (N_6092,N_5511,N_5646);
nand U6093 (N_6093,N_5694,N_5609);
xnor U6094 (N_6094,N_5552,N_5736);
and U6095 (N_6095,N_5629,N_5829);
nor U6096 (N_6096,N_5780,N_5618);
or U6097 (N_6097,N_5576,N_5954);
nor U6098 (N_6098,N_5939,N_5986);
and U6099 (N_6099,N_5990,N_5923);
nor U6100 (N_6100,N_5934,N_5636);
nor U6101 (N_6101,N_5651,N_5564);
xor U6102 (N_6102,N_5892,N_5504);
and U6103 (N_6103,N_5624,N_5716);
nand U6104 (N_6104,N_5710,N_5542);
and U6105 (N_6105,N_5582,N_5991);
nand U6106 (N_6106,N_5879,N_5770);
or U6107 (N_6107,N_5863,N_5663);
or U6108 (N_6108,N_5640,N_5763);
nand U6109 (N_6109,N_5854,N_5930);
nand U6110 (N_6110,N_5714,N_5905);
and U6111 (N_6111,N_5706,N_5535);
xnor U6112 (N_6112,N_5623,N_5806);
or U6113 (N_6113,N_5505,N_5816);
nand U6114 (N_6114,N_5638,N_5883);
and U6115 (N_6115,N_5931,N_5677);
nand U6116 (N_6116,N_5867,N_5569);
xor U6117 (N_6117,N_5768,N_5822);
or U6118 (N_6118,N_5767,N_5895);
xnor U6119 (N_6119,N_5762,N_5616);
or U6120 (N_6120,N_5711,N_5755);
and U6121 (N_6121,N_5533,N_5815);
nand U6122 (N_6122,N_5901,N_5828);
nor U6123 (N_6123,N_5584,N_5812);
xnor U6124 (N_6124,N_5625,N_5914);
nand U6125 (N_6125,N_5622,N_5902);
nor U6126 (N_6126,N_5720,N_5670);
and U6127 (N_6127,N_5835,N_5518);
xnor U6128 (N_6128,N_5682,N_5858);
or U6129 (N_6129,N_5941,N_5727);
xor U6130 (N_6130,N_5785,N_5888);
nand U6131 (N_6131,N_5617,N_5865);
nand U6132 (N_6132,N_5555,N_5935);
nand U6133 (N_6133,N_5961,N_5730);
or U6134 (N_6134,N_5913,N_5673);
nand U6135 (N_6135,N_5652,N_5753);
or U6136 (N_6136,N_5695,N_5702);
and U6137 (N_6137,N_5947,N_5544);
nand U6138 (N_6138,N_5675,N_5976);
nor U6139 (N_6139,N_5583,N_5538);
xor U6140 (N_6140,N_5703,N_5817);
xor U6141 (N_6141,N_5631,N_5704);
nor U6142 (N_6142,N_5627,N_5818);
xnor U6143 (N_6143,N_5717,N_5796);
nand U6144 (N_6144,N_5724,N_5574);
and U6145 (N_6145,N_5680,N_5614);
nand U6146 (N_6146,N_5696,N_5547);
or U6147 (N_6147,N_5987,N_5579);
and U6148 (N_6148,N_5880,N_5899);
xor U6149 (N_6149,N_5603,N_5925);
nor U6150 (N_6150,N_5669,N_5878);
and U6151 (N_6151,N_5633,N_5551);
or U6152 (N_6152,N_5659,N_5674);
and U6153 (N_6153,N_5676,N_5805);
nor U6154 (N_6154,N_5875,N_5726);
nand U6155 (N_6155,N_5958,N_5873);
or U6156 (N_6156,N_5777,N_5648);
nand U6157 (N_6157,N_5885,N_5626);
or U6158 (N_6158,N_5823,N_5968);
nand U6159 (N_6159,N_5515,N_5973);
or U6160 (N_6160,N_5918,N_5911);
or U6161 (N_6161,N_5859,N_5965);
xnor U6162 (N_6162,N_5571,N_5512);
nor U6163 (N_6163,N_5869,N_5520);
nand U6164 (N_6164,N_5985,N_5824);
nor U6165 (N_6165,N_5683,N_5715);
and U6166 (N_6166,N_5656,N_5539);
nor U6167 (N_6167,N_5994,N_5733);
nand U6168 (N_6168,N_5709,N_5549);
xnor U6169 (N_6169,N_5577,N_5526);
xor U6170 (N_6170,N_5671,N_5929);
and U6171 (N_6171,N_5955,N_5966);
nor U6172 (N_6172,N_5514,N_5997);
xnor U6173 (N_6173,N_5937,N_5660);
nor U6174 (N_6174,N_5513,N_5904);
nand U6175 (N_6175,N_5771,N_5978);
nand U6176 (N_6176,N_5591,N_5847);
and U6177 (N_6177,N_5944,N_5621);
or U6178 (N_6178,N_5814,N_5842);
nand U6179 (N_6179,N_5788,N_5974);
and U6180 (N_6180,N_5851,N_5566);
nand U6181 (N_6181,N_5732,N_5868);
xnor U6182 (N_6182,N_5938,N_5510);
or U6183 (N_6183,N_5856,N_5811);
nand U6184 (N_6184,N_5783,N_5665);
or U6185 (N_6185,N_5781,N_5516);
nor U6186 (N_6186,N_5738,N_5742);
or U6187 (N_6187,N_5527,N_5752);
xor U6188 (N_6188,N_5739,N_5776);
xnor U6189 (N_6189,N_5536,N_5912);
xnor U6190 (N_6190,N_5848,N_5871);
and U6191 (N_6191,N_5963,N_5969);
nand U6192 (N_6192,N_5841,N_5532);
nor U6193 (N_6193,N_5561,N_5613);
and U6194 (N_6194,N_5598,N_5921);
nand U6195 (N_6195,N_5857,N_5940);
or U6196 (N_6196,N_5772,N_5943);
and U6197 (N_6197,N_5757,N_5728);
xor U6198 (N_6198,N_5798,N_5595);
nor U6199 (N_6199,N_5778,N_5525);
or U6200 (N_6200,N_5999,N_5793);
nor U6201 (N_6201,N_5517,N_5964);
xnor U6202 (N_6202,N_5889,N_5907);
nand U6203 (N_6203,N_5604,N_5689);
and U6204 (N_6204,N_5688,N_5700);
and U6205 (N_6205,N_5852,N_5546);
or U6206 (N_6206,N_5634,N_5982);
xnor U6207 (N_6207,N_5575,N_5543);
xor U6208 (N_6208,N_5722,N_5524);
nor U6209 (N_6209,N_5983,N_5589);
and U6210 (N_6210,N_5988,N_5920);
or U6211 (N_6211,N_5810,N_5705);
or U6212 (N_6212,N_5872,N_5975);
nor U6213 (N_6213,N_5760,N_5919);
nand U6214 (N_6214,N_5605,N_5698);
or U6215 (N_6215,N_5799,N_5972);
and U6216 (N_6216,N_5959,N_5836);
and U6217 (N_6217,N_5610,N_5500);
or U6218 (N_6218,N_5599,N_5927);
nor U6219 (N_6219,N_5761,N_5557);
nand U6220 (N_6220,N_5882,N_5989);
nor U6221 (N_6221,N_5794,N_5690);
nor U6222 (N_6222,N_5748,N_5890);
nor U6223 (N_6223,N_5686,N_5853);
and U6224 (N_6224,N_5588,N_5650);
xor U6225 (N_6225,N_5529,N_5936);
and U6226 (N_6226,N_5775,N_5692);
nor U6227 (N_6227,N_5922,N_5635);
nand U6228 (N_6228,N_5541,N_5992);
xor U6229 (N_6229,N_5971,N_5585);
or U6230 (N_6230,N_5567,N_5658);
and U6231 (N_6231,N_5801,N_5657);
nand U6232 (N_6232,N_5765,N_5719);
and U6233 (N_6233,N_5924,N_5653);
and U6234 (N_6234,N_5729,N_5897);
nor U6235 (N_6235,N_5528,N_5838);
or U6236 (N_6236,N_5707,N_5735);
or U6237 (N_6237,N_5809,N_5998);
or U6238 (N_6238,N_5678,N_5592);
nand U6239 (N_6239,N_5896,N_5791);
nor U6240 (N_6240,N_5862,N_5531);
nor U6241 (N_6241,N_5501,N_5691);
nor U6242 (N_6242,N_5773,N_5832);
or U6243 (N_6243,N_5803,N_5556);
nand U6244 (N_6244,N_5750,N_5839);
and U6245 (N_6245,N_5578,N_5519);
xnor U6246 (N_6246,N_5507,N_5725);
nand U6247 (N_6247,N_5701,N_5967);
xnor U6248 (N_6248,N_5900,N_5855);
xor U6249 (N_6249,N_5628,N_5749);
or U6250 (N_6250,N_5751,N_5552);
nand U6251 (N_6251,N_5700,N_5963);
and U6252 (N_6252,N_5788,N_5663);
or U6253 (N_6253,N_5904,N_5631);
nor U6254 (N_6254,N_5933,N_5883);
nand U6255 (N_6255,N_5760,N_5758);
nor U6256 (N_6256,N_5976,N_5908);
or U6257 (N_6257,N_5639,N_5652);
nor U6258 (N_6258,N_5807,N_5715);
and U6259 (N_6259,N_5902,N_5603);
nand U6260 (N_6260,N_5908,N_5918);
xor U6261 (N_6261,N_5899,N_5948);
or U6262 (N_6262,N_5529,N_5512);
nor U6263 (N_6263,N_5753,N_5826);
nor U6264 (N_6264,N_5859,N_5714);
and U6265 (N_6265,N_5619,N_5957);
and U6266 (N_6266,N_5753,N_5977);
xor U6267 (N_6267,N_5789,N_5863);
nor U6268 (N_6268,N_5638,N_5523);
or U6269 (N_6269,N_5832,N_5958);
and U6270 (N_6270,N_5680,N_5809);
nand U6271 (N_6271,N_5807,N_5625);
or U6272 (N_6272,N_5799,N_5681);
and U6273 (N_6273,N_5633,N_5976);
nand U6274 (N_6274,N_5883,N_5653);
and U6275 (N_6275,N_5643,N_5627);
or U6276 (N_6276,N_5508,N_5748);
nand U6277 (N_6277,N_5873,N_5617);
nand U6278 (N_6278,N_5718,N_5821);
or U6279 (N_6279,N_5542,N_5667);
or U6280 (N_6280,N_5501,N_5826);
nor U6281 (N_6281,N_5645,N_5977);
nand U6282 (N_6282,N_5625,N_5811);
nand U6283 (N_6283,N_5601,N_5942);
xor U6284 (N_6284,N_5673,N_5600);
nand U6285 (N_6285,N_5876,N_5758);
and U6286 (N_6286,N_5533,N_5515);
and U6287 (N_6287,N_5886,N_5636);
xor U6288 (N_6288,N_5869,N_5682);
xor U6289 (N_6289,N_5940,N_5699);
or U6290 (N_6290,N_5840,N_5942);
and U6291 (N_6291,N_5508,N_5773);
and U6292 (N_6292,N_5944,N_5879);
nand U6293 (N_6293,N_5964,N_5910);
nor U6294 (N_6294,N_5763,N_5973);
xor U6295 (N_6295,N_5616,N_5621);
nor U6296 (N_6296,N_5786,N_5870);
xnor U6297 (N_6297,N_5993,N_5615);
nor U6298 (N_6298,N_5630,N_5798);
and U6299 (N_6299,N_5873,N_5649);
nand U6300 (N_6300,N_5806,N_5573);
and U6301 (N_6301,N_5766,N_5816);
nor U6302 (N_6302,N_5763,N_5591);
nor U6303 (N_6303,N_5659,N_5826);
xnor U6304 (N_6304,N_5522,N_5754);
nor U6305 (N_6305,N_5638,N_5864);
xnor U6306 (N_6306,N_5518,N_5655);
nand U6307 (N_6307,N_5807,N_5671);
xor U6308 (N_6308,N_5593,N_5860);
nor U6309 (N_6309,N_5503,N_5813);
xnor U6310 (N_6310,N_5800,N_5803);
nand U6311 (N_6311,N_5500,N_5702);
or U6312 (N_6312,N_5906,N_5508);
or U6313 (N_6313,N_5508,N_5676);
nor U6314 (N_6314,N_5560,N_5622);
and U6315 (N_6315,N_5753,N_5909);
nor U6316 (N_6316,N_5981,N_5602);
nor U6317 (N_6317,N_5574,N_5514);
nor U6318 (N_6318,N_5919,N_5548);
or U6319 (N_6319,N_5579,N_5774);
and U6320 (N_6320,N_5749,N_5983);
nor U6321 (N_6321,N_5908,N_5706);
nand U6322 (N_6322,N_5715,N_5684);
or U6323 (N_6323,N_5582,N_5879);
nand U6324 (N_6324,N_5599,N_5860);
or U6325 (N_6325,N_5610,N_5855);
nor U6326 (N_6326,N_5762,N_5941);
nor U6327 (N_6327,N_5536,N_5510);
and U6328 (N_6328,N_5835,N_5836);
xnor U6329 (N_6329,N_5721,N_5534);
nand U6330 (N_6330,N_5856,N_5592);
and U6331 (N_6331,N_5941,N_5992);
xor U6332 (N_6332,N_5814,N_5696);
nor U6333 (N_6333,N_5571,N_5777);
and U6334 (N_6334,N_5795,N_5998);
xnor U6335 (N_6335,N_5962,N_5817);
nand U6336 (N_6336,N_5955,N_5840);
xnor U6337 (N_6337,N_5890,N_5517);
nand U6338 (N_6338,N_5768,N_5504);
xnor U6339 (N_6339,N_5729,N_5982);
nand U6340 (N_6340,N_5572,N_5669);
nor U6341 (N_6341,N_5678,N_5696);
nand U6342 (N_6342,N_5796,N_5662);
and U6343 (N_6343,N_5688,N_5991);
nand U6344 (N_6344,N_5951,N_5647);
xnor U6345 (N_6345,N_5831,N_5754);
or U6346 (N_6346,N_5999,N_5570);
xor U6347 (N_6347,N_5740,N_5786);
and U6348 (N_6348,N_5976,N_5863);
or U6349 (N_6349,N_5824,N_5631);
and U6350 (N_6350,N_5981,N_5541);
xnor U6351 (N_6351,N_5553,N_5960);
and U6352 (N_6352,N_5687,N_5792);
nand U6353 (N_6353,N_5903,N_5576);
nand U6354 (N_6354,N_5814,N_5960);
xor U6355 (N_6355,N_5741,N_5660);
and U6356 (N_6356,N_5892,N_5822);
xnor U6357 (N_6357,N_5870,N_5788);
nand U6358 (N_6358,N_5599,N_5830);
xnor U6359 (N_6359,N_5852,N_5770);
and U6360 (N_6360,N_5767,N_5785);
or U6361 (N_6361,N_5745,N_5518);
and U6362 (N_6362,N_5685,N_5673);
xnor U6363 (N_6363,N_5744,N_5982);
nor U6364 (N_6364,N_5625,N_5570);
or U6365 (N_6365,N_5857,N_5992);
or U6366 (N_6366,N_5937,N_5958);
and U6367 (N_6367,N_5808,N_5532);
or U6368 (N_6368,N_5796,N_5782);
nor U6369 (N_6369,N_5965,N_5870);
nor U6370 (N_6370,N_5833,N_5594);
or U6371 (N_6371,N_5812,N_5587);
or U6372 (N_6372,N_5660,N_5851);
and U6373 (N_6373,N_5537,N_5624);
or U6374 (N_6374,N_5740,N_5652);
and U6375 (N_6375,N_5713,N_5765);
nand U6376 (N_6376,N_5840,N_5875);
or U6377 (N_6377,N_5783,N_5605);
and U6378 (N_6378,N_5947,N_5991);
xnor U6379 (N_6379,N_5713,N_5903);
and U6380 (N_6380,N_5862,N_5743);
nor U6381 (N_6381,N_5696,N_5873);
and U6382 (N_6382,N_5585,N_5912);
or U6383 (N_6383,N_5837,N_5693);
nand U6384 (N_6384,N_5752,N_5755);
nand U6385 (N_6385,N_5573,N_5544);
and U6386 (N_6386,N_5777,N_5787);
xnor U6387 (N_6387,N_5906,N_5614);
nand U6388 (N_6388,N_5967,N_5528);
nand U6389 (N_6389,N_5554,N_5687);
and U6390 (N_6390,N_5683,N_5642);
and U6391 (N_6391,N_5858,N_5646);
nor U6392 (N_6392,N_5705,N_5527);
nand U6393 (N_6393,N_5963,N_5633);
nand U6394 (N_6394,N_5805,N_5950);
nor U6395 (N_6395,N_5790,N_5775);
xnor U6396 (N_6396,N_5692,N_5764);
and U6397 (N_6397,N_5848,N_5846);
and U6398 (N_6398,N_5979,N_5729);
and U6399 (N_6399,N_5748,N_5531);
nand U6400 (N_6400,N_5864,N_5664);
nand U6401 (N_6401,N_5766,N_5762);
and U6402 (N_6402,N_5657,N_5722);
nand U6403 (N_6403,N_5834,N_5879);
xnor U6404 (N_6404,N_5511,N_5849);
or U6405 (N_6405,N_5956,N_5503);
xnor U6406 (N_6406,N_5763,N_5728);
nor U6407 (N_6407,N_5949,N_5893);
and U6408 (N_6408,N_5627,N_5960);
nor U6409 (N_6409,N_5596,N_5501);
nand U6410 (N_6410,N_5577,N_5795);
xor U6411 (N_6411,N_5678,N_5955);
or U6412 (N_6412,N_5590,N_5923);
nand U6413 (N_6413,N_5834,N_5530);
nand U6414 (N_6414,N_5846,N_5646);
nor U6415 (N_6415,N_5924,N_5545);
nand U6416 (N_6416,N_5612,N_5791);
nand U6417 (N_6417,N_5617,N_5944);
nor U6418 (N_6418,N_5571,N_5563);
or U6419 (N_6419,N_5762,N_5788);
xnor U6420 (N_6420,N_5900,N_5901);
or U6421 (N_6421,N_5693,N_5639);
xnor U6422 (N_6422,N_5523,N_5649);
nor U6423 (N_6423,N_5676,N_5534);
or U6424 (N_6424,N_5962,N_5838);
xnor U6425 (N_6425,N_5730,N_5752);
xor U6426 (N_6426,N_5707,N_5872);
xnor U6427 (N_6427,N_5566,N_5521);
nand U6428 (N_6428,N_5861,N_5640);
or U6429 (N_6429,N_5739,N_5867);
and U6430 (N_6430,N_5755,N_5666);
and U6431 (N_6431,N_5505,N_5654);
nand U6432 (N_6432,N_5511,N_5508);
nor U6433 (N_6433,N_5616,N_5588);
and U6434 (N_6434,N_5734,N_5555);
nand U6435 (N_6435,N_5920,N_5772);
nand U6436 (N_6436,N_5606,N_5604);
or U6437 (N_6437,N_5583,N_5986);
nand U6438 (N_6438,N_5756,N_5743);
and U6439 (N_6439,N_5759,N_5819);
nand U6440 (N_6440,N_5968,N_5960);
nor U6441 (N_6441,N_5615,N_5765);
or U6442 (N_6442,N_5950,N_5750);
xnor U6443 (N_6443,N_5864,N_5866);
xor U6444 (N_6444,N_5802,N_5537);
or U6445 (N_6445,N_5683,N_5808);
xor U6446 (N_6446,N_5820,N_5843);
xor U6447 (N_6447,N_5573,N_5607);
and U6448 (N_6448,N_5860,N_5945);
nor U6449 (N_6449,N_5837,N_5565);
xnor U6450 (N_6450,N_5698,N_5937);
xnor U6451 (N_6451,N_5942,N_5990);
nand U6452 (N_6452,N_5797,N_5661);
xnor U6453 (N_6453,N_5775,N_5752);
xnor U6454 (N_6454,N_5823,N_5664);
nor U6455 (N_6455,N_5761,N_5658);
or U6456 (N_6456,N_5962,N_5832);
xnor U6457 (N_6457,N_5905,N_5658);
nor U6458 (N_6458,N_5933,N_5639);
and U6459 (N_6459,N_5545,N_5606);
xor U6460 (N_6460,N_5840,N_5781);
nor U6461 (N_6461,N_5560,N_5929);
xnor U6462 (N_6462,N_5995,N_5764);
nand U6463 (N_6463,N_5503,N_5736);
xor U6464 (N_6464,N_5688,N_5862);
nand U6465 (N_6465,N_5667,N_5632);
nor U6466 (N_6466,N_5685,N_5844);
or U6467 (N_6467,N_5660,N_5798);
nand U6468 (N_6468,N_5725,N_5712);
xor U6469 (N_6469,N_5505,N_5959);
and U6470 (N_6470,N_5912,N_5844);
or U6471 (N_6471,N_5898,N_5650);
or U6472 (N_6472,N_5923,N_5684);
nor U6473 (N_6473,N_5562,N_5882);
or U6474 (N_6474,N_5557,N_5593);
xor U6475 (N_6475,N_5929,N_5825);
xnor U6476 (N_6476,N_5696,N_5911);
nand U6477 (N_6477,N_5595,N_5650);
xor U6478 (N_6478,N_5860,N_5927);
xor U6479 (N_6479,N_5927,N_5982);
nand U6480 (N_6480,N_5667,N_5626);
or U6481 (N_6481,N_5833,N_5523);
xnor U6482 (N_6482,N_5978,N_5973);
xor U6483 (N_6483,N_5841,N_5898);
nor U6484 (N_6484,N_5680,N_5972);
nor U6485 (N_6485,N_5536,N_5578);
or U6486 (N_6486,N_5603,N_5753);
xnor U6487 (N_6487,N_5731,N_5956);
or U6488 (N_6488,N_5766,N_5858);
and U6489 (N_6489,N_5534,N_5932);
and U6490 (N_6490,N_5957,N_5951);
or U6491 (N_6491,N_5937,N_5642);
and U6492 (N_6492,N_5624,N_5546);
xnor U6493 (N_6493,N_5917,N_5920);
nor U6494 (N_6494,N_5652,N_5536);
or U6495 (N_6495,N_5705,N_5995);
nor U6496 (N_6496,N_5657,N_5636);
xnor U6497 (N_6497,N_5596,N_5955);
and U6498 (N_6498,N_5975,N_5927);
xnor U6499 (N_6499,N_5844,N_5795);
nand U6500 (N_6500,N_6385,N_6274);
xnor U6501 (N_6501,N_6227,N_6279);
nor U6502 (N_6502,N_6293,N_6225);
nor U6503 (N_6503,N_6264,N_6401);
or U6504 (N_6504,N_6381,N_6424);
or U6505 (N_6505,N_6246,N_6085);
nor U6506 (N_6506,N_6162,N_6257);
and U6507 (N_6507,N_6319,N_6355);
nor U6508 (N_6508,N_6129,N_6062);
and U6509 (N_6509,N_6393,N_6300);
nor U6510 (N_6510,N_6347,N_6171);
and U6511 (N_6511,N_6294,N_6242);
xor U6512 (N_6512,N_6166,N_6406);
nand U6513 (N_6513,N_6275,N_6057);
xor U6514 (N_6514,N_6405,N_6445);
nand U6515 (N_6515,N_6025,N_6286);
xnor U6516 (N_6516,N_6343,N_6188);
nor U6517 (N_6517,N_6098,N_6441);
and U6518 (N_6518,N_6459,N_6449);
xnor U6519 (N_6519,N_6408,N_6303);
and U6520 (N_6520,N_6462,N_6452);
xor U6521 (N_6521,N_6439,N_6335);
or U6522 (N_6522,N_6460,N_6316);
xor U6523 (N_6523,N_6486,N_6193);
nand U6524 (N_6524,N_6321,N_6147);
nand U6525 (N_6525,N_6172,N_6397);
nand U6526 (N_6526,N_6291,N_6498);
nor U6527 (N_6527,N_6083,N_6099);
nor U6528 (N_6528,N_6182,N_6320);
nand U6529 (N_6529,N_6280,N_6387);
nor U6530 (N_6530,N_6283,N_6238);
nor U6531 (N_6531,N_6032,N_6113);
nor U6532 (N_6532,N_6499,N_6281);
xnor U6533 (N_6533,N_6164,N_6497);
or U6534 (N_6534,N_6383,N_6042);
nor U6535 (N_6535,N_6268,N_6101);
or U6536 (N_6536,N_6369,N_6103);
or U6537 (N_6537,N_6107,N_6327);
and U6538 (N_6538,N_6465,N_6448);
and U6539 (N_6539,N_6367,N_6248);
and U6540 (N_6540,N_6375,N_6218);
xnor U6541 (N_6541,N_6191,N_6346);
and U6542 (N_6542,N_6488,N_6469);
and U6543 (N_6543,N_6458,N_6413);
nand U6544 (N_6544,N_6019,N_6230);
xor U6545 (N_6545,N_6338,N_6040);
and U6546 (N_6546,N_6376,N_6250);
or U6547 (N_6547,N_6144,N_6084);
nor U6548 (N_6548,N_6466,N_6145);
or U6549 (N_6549,N_6453,N_6152);
nand U6550 (N_6550,N_6051,N_6208);
nor U6551 (N_6551,N_6111,N_6484);
nand U6552 (N_6552,N_6239,N_6259);
xor U6553 (N_6553,N_6349,N_6070);
nor U6554 (N_6554,N_6154,N_6296);
and U6555 (N_6555,N_6136,N_6480);
and U6556 (N_6556,N_6059,N_6391);
and U6557 (N_6557,N_6295,N_6022);
and U6558 (N_6558,N_6194,N_6024);
or U6559 (N_6559,N_6241,N_6287);
xnor U6560 (N_6560,N_6026,N_6243);
nand U6561 (N_6561,N_6033,N_6472);
or U6562 (N_6562,N_6461,N_6456);
or U6563 (N_6563,N_6000,N_6282);
nor U6564 (N_6564,N_6245,N_6065);
and U6565 (N_6565,N_6487,N_6148);
and U6566 (N_6566,N_6322,N_6077);
xor U6567 (N_6567,N_6262,N_6035);
nor U6568 (N_6568,N_6211,N_6201);
and U6569 (N_6569,N_6039,N_6117);
nor U6570 (N_6570,N_6273,N_6203);
nand U6571 (N_6571,N_6324,N_6180);
nand U6572 (N_6572,N_6217,N_6097);
nor U6573 (N_6573,N_6265,N_6421);
and U6574 (N_6574,N_6003,N_6046);
xor U6575 (N_6575,N_6011,N_6207);
and U6576 (N_6576,N_6244,N_6030);
nand U6577 (N_6577,N_6185,N_6336);
or U6578 (N_6578,N_6231,N_6373);
nor U6579 (N_6579,N_6197,N_6204);
nor U6580 (N_6580,N_6072,N_6108);
and U6581 (N_6581,N_6475,N_6457);
and U6582 (N_6582,N_6429,N_6183);
nor U6583 (N_6583,N_6087,N_6356);
nand U6584 (N_6584,N_6184,N_6482);
or U6585 (N_6585,N_6410,N_6261);
xnor U6586 (N_6586,N_6292,N_6044);
nand U6587 (N_6587,N_6403,N_6399);
and U6588 (N_6588,N_6012,N_6020);
and U6589 (N_6589,N_6006,N_6306);
xor U6590 (N_6590,N_6431,N_6390);
xnor U6591 (N_6591,N_6029,N_6134);
xnor U6592 (N_6592,N_6080,N_6340);
xor U6593 (N_6593,N_6221,N_6168);
and U6594 (N_6594,N_6314,N_6366);
and U6595 (N_6595,N_6068,N_6483);
or U6596 (N_6596,N_6198,N_6414);
xor U6597 (N_6597,N_6229,N_6008);
nand U6598 (N_6598,N_6380,N_6119);
nor U6599 (N_6599,N_6137,N_6474);
nand U6600 (N_6600,N_6021,N_6337);
nor U6601 (N_6601,N_6061,N_6023);
nand U6602 (N_6602,N_6444,N_6330);
or U6603 (N_6603,N_6386,N_6479);
or U6604 (N_6604,N_6496,N_6492);
xor U6605 (N_6605,N_6156,N_6052);
xnor U6606 (N_6606,N_6140,N_6210);
xnor U6607 (N_6607,N_6446,N_6277);
xor U6608 (N_6608,N_6240,N_6106);
xnor U6609 (N_6609,N_6220,N_6278);
nor U6610 (N_6610,N_6071,N_6426);
xor U6611 (N_6611,N_6195,N_6471);
and U6612 (N_6612,N_6269,N_6133);
xnor U6613 (N_6613,N_6089,N_6345);
nor U6614 (N_6614,N_6150,N_6377);
nand U6615 (N_6615,N_6223,N_6001);
and U6616 (N_6616,N_6402,N_6212);
xnor U6617 (N_6617,N_6213,N_6132);
and U6618 (N_6618,N_6031,N_6219);
xnor U6619 (N_6619,N_6468,N_6120);
and U6620 (N_6620,N_6232,N_6114);
xor U6621 (N_6621,N_6477,N_6216);
nor U6622 (N_6622,N_6224,N_6396);
nor U6623 (N_6623,N_6272,N_6297);
xnor U6624 (N_6624,N_6334,N_6090);
or U6625 (N_6625,N_6249,N_6360);
or U6626 (N_6626,N_6374,N_6010);
xnor U6627 (N_6627,N_6434,N_6435);
nand U6628 (N_6628,N_6313,N_6094);
xor U6629 (N_6629,N_6004,N_6473);
xor U6630 (N_6630,N_6491,N_6058);
or U6631 (N_6631,N_6371,N_6438);
and U6632 (N_6632,N_6308,N_6440);
xnor U6633 (N_6633,N_6161,N_6494);
nor U6634 (N_6634,N_6315,N_6476);
or U6635 (N_6635,N_6155,N_6237);
and U6636 (N_6636,N_6088,N_6454);
nor U6637 (N_6637,N_6384,N_6290);
and U6638 (N_6638,N_6153,N_6309);
or U6639 (N_6639,N_6190,N_6192);
nand U6640 (N_6640,N_6187,N_6395);
or U6641 (N_6641,N_6093,N_6017);
or U6642 (N_6642,N_6339,N_6102);
nand U6643 (N_6643,N_6159,N_6368);
nand U6644 (N_6644,N_6415,N_6307);
xnor U6645 (N_6645,N_6422,N_6049);
nand U6646 (N_6646,N_6143,N_6370);
nand U6647 (N_6647,N_6382,N_6412);
and U6648 (N_6648,N_6121,N_6357);
nor U6649 (N_6649,N_6247,N_6178);
nand U6650 (N_6650,N_6091,N_6214);
nor U6651 (N_6651,N_6354,N_6236);
xor U6652 (N_6652,N_6416,N_6151);
nand U6653 (N_6653,N_6331,N_6251);
nor U6654 (N_6654,N_6116,N_6455);
nand U6655 (N_6655,N_6299,N_6350);
or U6656 (N_6656,N_6173,N_6222);
nand U6657 (N_6657,N_6018,N_6199);
nand U6658 (N_6658,N_6418,N_6060);
nand U6659 (N_6659,N_6430,N_6392);
xnor U6660 (N_6660,N_6139,N_6054);
and U6661 (N_6661,N_6045,N_6149);
xor U6662 (N_6662,N_6353,N_6053);
nor U6663 (N_6663,N_6342,N_6228);
xnor U6664 (N_6664,N_6082,N_6398);
xnor U6665 (N_6665,N_6043,N_6409);
nor U6666 (N_6666,N_6163,N_6433);
xnor U6667 (N_6667,N_6005,N_6263);
and U6668 (N_6668,N_6419,N_6305);
nor U6669 (N_6669,N_6495,N_6425);
and U6670 (N_6670,N_6362,N_6411);
nand U6671 (N_6671,N_6186,N_6447);
xor U6672 (N_6672,N_6179,N_6170);
or U6673 (N_6673,N_6302,N_6311);
nor U6674 (N_6674,N_6141,N_6036);
xor U6675 (N_6675,N_6007,N_6235);
nor U6676 (N_6676,N_6378,N_6437);
or U6677 (N_6677,N_6365,N_6325);
nor U6678 (N_6678,N_6196,N_6048);
or U6679 (N_6679,N_6205,N_6358);
and U6680 (N_6680,N_6432,N_6389);
and U6681 (N_6681,N_6009,N_6451);
and U6682 (N_6682,N_6128,N_6013);
xor U6683 (N_6683,N_6326,N_6436);
and U6684 (N_6684,N_6127,N_6014);
or U6685 (N_6685,N_6165,N_6189);
nand U6686 (N_6686,N_6252,N_6075);
or U6687 (N_6687,N_6328,N_6233);
nand U6688 (N_6688,N_6086,N_6174);
xnor U6689 (N_6689,N_6142,N_6038);
or U6690 (N_6690,N_6267,N_6135);
nand U6691 (N_6691,N_6323,N_6427);
xor U6692 (N_6692,N_6276,N_6400);
and U6693 (N_6693,N_6420,N_6177);
and U6694 (N_6694,N_6055,N_6226);
and U6695 (N_6695,N_6175,N_6125);
nand U6696 (N_6696,N_6074,N_6359);
xnor U6697 (N_6697,N_6379,N_6363);
and U6698 (N_6698,N_6417,N_6002);
nor U6699 (N_6699,N_6206,N_6202);
or U6700 (N_6700,N_6123,N_6064);
xnor U6701 (N_6701,N_6289,N_6388);
nand U6702 (N_6702,N_6200,N_6463);
nor U6703 (N_6703,N_6255,N_6442);
or U6704 (N_6704,N_6100,N_6104);
and U6705 (N_6705,N_6122,N_6169);
nor U6706 (N_6706,N_6467,N_6318);
and U6707 (N_6707,N_6176,N_6041);
or U6708 (N_6708,N_6364,N_6481);
nand U6709 (N_6709,N_6266,N_6493);
xor U6710 (N_6710,N_6450,N_6352);
and U6711 (N_6711,N_6181,N_6095);
xnor U6712 (N_6712,N_6490,N_6160);
xnor U6713 (N_6713,N_6284,N_6271);
xor U6714 (N_6714,N_6050,N_6146);
nor U6715 (N_6715,N_6047,N_6258);
xor U6716 (N_6716,N_6407,N_6478);
and U6717 (N_6717,N_6270,N_6254);
or U6718 (N_6718,N_6076,N_6037);
nand U6719 (N_6719,N_6361,N_6063);
nand U6720 (N_6720,N_6130,N_6118);
or U6721 (N_6721,N_6167,N_6348);
nand U6722 (N_6722,N_6404,N_6288);
or U6723 (N_6723,N_6256,N_6301);
xor U6724 (N_6724,N_6110,N_6351);
or U6725 (N_6725,N_6310,N_6423);
or U6726 (N_6726,N_6027,N_6285);
nand U6727 (N_6727,N_6138,N_6443);
or U6728 (N_6728,N_6109,N_6372);
nor U6729 (N_6729,N_6332,N_6464);
xnor U6730 (N_6730,N_6105,N_6428);
nand U6731 (N_6731,N_6344,N_6333);
and U6732 (N_6732,N_6394,N_6158);
or U6733 (N_6733,N_6253,N_6073);
or U6734 (N_6734,N_6312,N_6470);
xor U6735 (N_6735,N_6034,N_6131);
nor U6736 (N_6736,N_6078,N_6304);
and U6737 (N_6737,N_6489,N_6298);
xor U6738 (N_6738,N_6079,N_6260);
xnor U6739 (N_6739,N_6081,N_6096);
or U6740 (N_6740,N_6069,N_6067);
or U6741 (N_6741,N_6092,N_6028);
and U6742 (N_6742,N_6234,N_6341);
nand U6743 (N_6743,N_6329,N_6485);
nand U6744 (N_6744,N_6015,N_6209);
or U6745 (N_6745,N_6112,N_6126);
or U6746 (N_6746,N_6317,N_6157);
or U6747 (N_6747,N_6124,N_6016);
xnor U6748 (N_6748,N_6056,N_6215);
xnor U6749 (N_6749,N_6115,N_6066);
and U6750 (N_6750,N_6337,N_6072);
or U6751 (N_6751,N_6190,N_6264);
nor U6752 (N_6752,N_6235,N_6171);
xnor U6753 (N_6753,N_6200,N_6017);
nand U6754 (N_6754,N_6360,N_6405);
xor U6755 (N_6755,N_6362,N_6225);
nor U6756 (N_6756,N_6382,N_6462);
xor U6757 (N_6757,N_6384,N_6292);
or U6758 (N_6758,N_6003,N_6273);
and U6759 (N_6759,N_6015,N_6310);
and U6760 (N_6760,N_6064,N_6051);
or U6761 (N_6761,N_6072,N_6412);
or U6762 (N_6762,N_6252,N_6416);
xnor U6763 (N_6763,N_6158,N_6353);
nor U6764 (N_6764,N_6286,N_6166);
or U6765 (N_6765,N_6490,N_6134);
xnor U6766 (N_6766,N_6103,N_6290);
nor U6767 (N_6767,N_6138,N_6257);
nor U6768 (N_6768,N_6454,N_6143);
xnor U6769 (N_6769,N_6413,N_6201);
nand U6770 (N_6770,N_6133,N_6475);
and U6771 (N_6771,N_6370,N_6081);
xnor U6772 (N_6772,N_6498,N_6299);
nand U6773 (N_6773,N_6295,N_6390);
and U6774 (N_6774,N_6202,N_6008);
xnor U6775 (N_6775,N_6330,N_6434);
and U6776 (N_6776,N_6033,N_6111);
and U6777 (N_6777,N_6177,N_6257);
nand U6778 (N_6778,N_6061,N_6361);
or U6779 (N_6779,N_6181,N_6469);
and U6780 (N_6780,N_6116,N_6472);
nand U6781 (N_6781,N_6290,N_6458);
nor U6782 (N_6782,N_6211,N_6188);
and U6783 (N_6783,N_6187,N_6231);
nand U6784 (N_6784,N_6496,N_6159);
and U6785 (N_6785,N_6294,N_6487);
xor U6786 (N_6786,N_6191,N_6207);
xnor U6787 (N_6787,N_6401,N_6320);
nor U6788 (N_6788,N_6202,N_6268);
nor U6789 (N_6789,N_6215,N_6311);
or U6790 (N_6790,N_6258,N_6434);
nand U6791 (N_6791,N_6410,N_6047);
or U6792 (N_6792,N_6398,N_6437);
nand U6793 (N_6793,N_6263,N_6470);
nand U6794 (N_6794,N_6090,N_6158);
and U6795 (N_6795,N_6175,N_6285);
nor U6796 (N_6796,N_6270,N_6155);
and U6797 (N_6797,N_6179,N_6400);
and U6798 (N_6798,N_6073,N_6144);
xnor U6799 (N_6799,N_6019,N_6155);
and U6800 (N_6800,N_6444,N_6431);
nand U6801 (N_6801,N_6300,N_6321);
nor U6802 (N_6802,N_6314,N_6469);
nand U6803 (N_6803,N_6326,N_6467);
nand U6804 (N_6804,N_6142,N_6185);
nor U6805 (N_6805,N_6280,N_6270);
nand U6806 (N_6806,N_6079,N_6176);
and U6807 (N_6807,N_6062,N_6340);
nor U6808 (N_6808,N_6341,N_6101);
and U6809 (N_6809,N_6161,N_6414);
nor U6810 (N_6810,N_6471,N_6039);
nor U6811 (N_6811,N_6231,N_6378);
nand U6812 (N_6812,N_6057,N_6334);
xnor U6813 (N_6813,N_6188,N_6139);
or U6814 (N_6814,N_6477,N_6393);
xor U6815 (N_6815,N_6161,N_6151);
or U6816 (N_6816,N_6131,N_6221);
and U6817 (N_6817,N_6087,N_6186);
xnor U6818 (N_6818,N_6431,N_6367);
nand U6819 (N_6819,N_6151,N_6195);
and U6820 (N_6820,N_6194,N_6493);
nand U6821 (N_6821,N_6058,N_6275);
nor U6822 (N_6822,N_6156,N_6408);
xor U6823 (N_6823,N_6276,N_6478);
and U6824 (N_6824,N_6333,N_6225);
and U6825 (N_6825,N_6470,N_6059);
or U6826 (N_6826,N_6224,N_6214);
xor U6827 (N_6827,N_6466,N_6215);
and U6828 (N_6828,N_6387,N_6086);
xor U6829 (N_6829,N_6367,N_6470);
xnor U6830 (N_6830,N_6492,N_6081);
nand U6831 (N_6831,N_6195,N_6103);
or U6832 (N_6832,N_6147,N_6172);
nand U6833 (N_6833,N_6323,N_6017);
nor U6834 (N_6834,N_6031,N_6340);
or U6835 (N_6835,N_6445,N_6492);
xnor U6836 (N_6836,N_6397,N_6132);
and U6837 (N_6837,N_6063,N_6067);
xnor U6838 (N_6838,N_6199,N_6176);
nor U6839 (N_6839,N_6286,N_6311);
nor U6840 (N_6840,N_6402,N_6032);
and U6841 (N_6841,N_6200,N_6399);
and U6842 (N_6842,N_6312,N_6259);
and U6843 (N_6843,N_6384,N_6314);
xor U6844 (N_6844,N_6307,N_6341);
xor U6845 (N_6845,N_6412,N_6313);
or U6846 (N_6846,N_6161,N_6123);
nand U6847 (N_6847,N_6352,N_6078);
nor U6848 (N_6848,N_6283,N_6035);
nand U6849 (N_6849,N_6491,N_6104);
and U6850 (N_6850,N_6314,N_6232);
xor U6851 (N_6851,N_6129,N_6329);
nor U6852 (N_6852,N_6073,N_6098);
or U6853 (N_6853,N_6419,N_6224);
xnor U6854 (N_6854,N_6110,N_6184);
nand U6855 (N_6855,N_6411,N_6367);
or U6856 (N_6856,N_6228,N_6000);
xnor U6857 (N_6857,N_6147,N_6063);
nand U6858 (N_6858,N_6191,N_6445);
nor U6859 (N_6859,N_6045,N_6168);
nand U6860 (N_6860,N_6489,N_6006);
nor U6861 (N_6861,N_6012,N_6173);
nor U6862 (N_6862,N_6409,N_6491);
nor U6863 (N_6863,N_6348,N_6353);
xnor U6864 (N_6864,N_6102,N_6109);
nor U6865 (N_6865,N_6008,N_6010);
nor U6866 (N_6866,N_6220,N_6066);
nand U6867 (N_6867,N_6391,N_6394);
and U6868 (N_6868,N_6270,N_6069);
and U6869 (N_6869,N_6076,N_6326);
xor U6870 (N_6870,N_6040,N_6134);
nand U6871 (N_6871,N_6472,N_6299);
and U6872 (N_6872,N_6406,N_6304);
nand U6873 (N_6873,N_6302,N_6424);
and U6874 (N_6874,N_6399,N_6152);
nand U6875 (N_6875,N_6378,N_6072);
nor U6876 (N_6876,N_6318,N_6255);
xor U6877 (N_6877,N_6012,N_6134);
and U6878 (N_6878,N_6015,N_6041);
nand U6879 (N_6879,N_6036,N_6207);
nand U6880 (N_6880,N_6347,N_6080);
or U6881 (N_6881,N_6110,N_6290);
nor U6882 (N_6882,N_6457,N_6344);
xnor U6883 (N_6883,N_6280,N_6061);
nand U6884 (N_6884,N_6168,N_6366);
nand U6885 (N_6885,N_6126,N_6398);
or U6886 (N_6886,N_6355,N_6249);
or U6887 (N_6887,N_6183,N_6143);
or U6888 (N_6888,N_6305,N_6131);
and U6889 (N_6889,N_6353,N_6088);
or U6890 (N_6890,N_6034,N_6417);
nand U6891 (N_6891,N_6169,N_6045);
xnor U6892 (N_6892,N_6345,N_6249);
nand U6893 (N_6893,N_6476,N_6087);
or U6894 (N_6894,N_6270,N_6175);
and U6895 (N_6895,N_6222,N_6144);
xnor U6896 (N_6896,N_6264,N_6140);
or U6897 (N_6897,N_6302,N_6108);
xnor U6898 (N_6898,N_6403,N_6255);
nand U6899 (N_6899,N_6364,N_6330);
nand U6900 (N_6900,N_6360,N_6369);
nor U6901 (N_6901,N_6466,N_6237);
nor U6902 (N_6902,N_6145,N_6270);
nor U6903 (N_6903,N_6138,N_6193);
and U6904 (N_6904,N_6412,N_6374);
nor U6905 (N_6905,N_6187,N_6382);
and U6906 (N_6906,N_6040,N_6250);
nand U6907 (N_6907,N_6366,N_6109);
xor U6908 (N_6908,N_6324,N_6356);
nand U6909 (N_6909,N_6456,N_6179);
nor U6910 (N_6910,N_6406,N_6498);
and U6911 (N_6911,N_6211,N_6294);
and U6912 (N_6912,N_6131,N_6317);
xnor U6913 (N_6913,N_6021,N_6484);
or U6914 (N_6914,N_6332,N_6289);
and U6915 (N_6915,N_6088,N_6293);
and U6916 (N_6916,N_6172,N_6141);
nor U6917 (N_6917,N_6377,N_6122);
and U6918 (N_6918,N_6320,N_6125);
nand U6919 (N_6919,N_6150,N_6284);
or U6920 (N_6920,N_6095,N_6308);
nand U6921 (N_6921,N_6261,N_6308);
nor U6922 (N_6922,N_6133,N_6300);
nand U6923 (N_6923,N_6112,N_6039);
and U6924 (N_6924,N_6010,N_6377);
xor U6925 (N_6925,N_6186,N_6219);
or U6926 (N_6926,N_6462,N_6000);
nor U6927 (N_6927,N_6006,N_6354);
or U6928 (N_6928,N_6158,N_6043);
or U6929 (N_6929,N_6266,N_6321);
and U6930 (N_6930,N_6383,N_6385);
xnor U6931 (N_6931,N_6275,N_6262);
nor U6932 (N_6932,N_6397,N_6273);
and U6933 (N_6933,N_6091,N_6065);
or U6934 (N_6934,N_6150,N_6425);
xnor U6935 (N_6935,N_6497,N_6249);
xor U6936 (N_6936,N_6223,N_6082);
nor U6937 (N_6937,N_6132,N_6467);
xor U6938 (N_6938,N_6437,N_6403);
nand U6939 (N_6939,N_6117,N_6372);
xor U6940 (N_6940,N_6048,N_6430);
xor U6941 (N_6941,N_6381,N_6014);
nor U6942 (N_6942,N_6200,N_6182);
and U6943 (N_6943,N_6245,N_6460);
xnor U6944 (N_6944,N_6088,N_6377);
and U6945 (N_6945,N_6298,N_6137);
or U6946 (N_6946,N_6087,N_6267);
xnor U6947 (N_6947,N_6130,N_6170);
nor U6948 (N_6948,N_6201,N_6161);
nor U6949 (N_6949,N_6309,N_6191);
and U6950 (N_6950,N_6480,N_6424);
xor U6951 (N_6951,N_6167,N_6074);
xor U6952 (N_6952,N_6461,N_6401);
or U6953 (N_6953,N_6130,N_6288);
or U6954 (N_6954,N_6376,N_6490);
nor U6955 (N_6955,N_6327,N_6191);
nand U6956 (N_6956,N_6091,N_6137);
nand U6957 (N_6957,N_6092,N_6227);
or U6958 (N_6958,N_6404,N_6196);
nand U6959 (N_6959,N_6417,N_6237);
and U6960 (N_6960,N_6334,N_6336);
or U6961 (N_6961,N_6202,N_6167);
nand U6962 (N_6962,N_6393,N_6298);
and U6963 (N_6963,N_6106,N_6493);
nor U6964 (N_6964,N_6041,N_6461);
nand U6965 (N_6965,N_6490,N_6440);
and U6966 (N_6966,N_6416,N_6322);
nor U6967 (N_6967,N_6460,N_6377);
xnor U6968 (N_6968,N_6023,N_6359);
or U6969 (N_6969,N_6061,N_6019);
xor U6970 (N_6970,N_6127,N_6142);
nor U6971 (N_6971,N_6227,N_6274);
nor U6972 (N_6972,N_6010,N_6174);
nand U6973 (N_6973,N_6282,N_6343);
nor U6974 (N_6974,N_6438,N_6065);
nor U6975 (N_6975,N_6482,N_6293);
nand U6976 (N_6976,N_6473,N_6393);
nand U6977 (N_6977,N_6145,N_6396);
or U6978 (N_6978,N_6307,N_6030);
nand U6979 (N_6979,N_6069,N_6040);
and U6980 (N_6980,N_6330,N_6036);
and U6981 (N_6981,N_6330,N_6161);
nor U6982 (N_6982,N_6443,N_6294);
nand U6983 (N_6983,N_6127,N_6085);
nand U6984 (N_6984,N_6289,N_6081);
and U6985 (N_6985,N_6321,N_6024);
xor U6986 (N_6986,N_6375,N_6272);
nand U6987 (N_6987,N_6264,N_6344);
xor U6988 (N_6988,N_6323,N_6169);
nand U6989 (N_6989,N_6248,N_6359);
nand U6990 (N_6990,N_6339,N_6409);
xnor U6991 (N_6991,N_6324,N_6106);
xor U6992 (N_6992,N_6397,N_6201);
and U6993 (N_6993,N_6130,N_6439);
and U6994 (N_6994,N_6323,N_6194);
and U6995 (N_6995,N_6069,N_6339);
nor U6996 (N_6996,N_6322,N_6013);
nand U6997 (N_6997,N_6329,N_6202);
nand U6998 (N_6998,N_6394,N_6012);
xor U6999 (N_6999,N_6250,N_6345);
or U7000 (N_7000,N_6622,N_6577);
and U7001 (N_7001,N_6960,N_6867);
nor U7002 (N_7002,N_6701,N_6978);
or U7003 (N_7003,N_6989,N_6783);
xnor U7004 (N_7004,N_6579,N_6687);
nor U7005 (N_7005,N_6980,N_6886);
and U7006 (N_7006,N_6694,N_6606);
or U7007 (N_7007,N_6559,N_6778);
nor U7008 (N_7008,N_6809,N_6772);
nor U7009 (N_7009,N_6658,N_6927);
or U7010 (N_7010,N_6561,N_6776);
and U7011 (N_7011,N_6923,N_6562);
or U7012 (N_7012,N_6620,N_6727);
and U7013 (N_7013,N_6864,N_6839);
nand U7014 (N_7014,N_6901,N_6899);
xor U7015 (N_7015,N_6844,N_6972);
nand U7016 (N_7016,N_6734,N_6878);
or U7017 (N_7017,N_6615,N_6906);
xor U7018 (N_7018,N_6806,N_6730);
or U7019 (N_7019,N_6888,N_6711);
nand U7020 (N_7020,N_6702,N_6507);
nor U7021 (N_7021,N_6852,N_6969);
or U7022 (N_7022,N_6721,N_6657);
or U7023 (N_7023,N_6576,N_6633);
and U7024 (N_7024,N_6858,N_6638);
xnor U7025 (N_7025,N_6760,N_6926);
and U7026 (N_7026,N_6509,N_6933);
xnor U7027 (N_7027,N_6823,N_6765);
or U7028 (N_7028,N_6982,N_6555);
or U7029 (N_7029,N_6900,N_6924);
nor U7030 (N_7030,N_6985,N_6803);
nor U7031 (N_7031,N_6649,N_6580);
or U7032 (N_7032,N_6748,N_6767);
and U7033 (N_7033,N_6594,N_6801);
nor U7034 (N_7034,N_6522,N_6849);
nand U7035 (N_7035,N_6533,N_6909);
and U7036 (N_7036,N_6531,N_6920);
xor U7037 (N_7037,N_6644,N_6530);
or U7038 (N_7038,N_6796,N_6655);
xor U7039 (N_7039,N_6674,N_6830);
and U7040 (N_7040,N_6520,N_6557);
nor U7041 (N_7041,N_6877,N_6722);
and U7042 (N_7042,N_6570,N_6661);
and U7043 (N_7043,N_6546,N_6527);
nand U7044 (N_7044,N_6681,N_6846);
and U7045 (N_7045,N_6784,N_6810);
or U7046 (N_7046,N_6829,N_6571);
and U7047 (N_7047,N_6952,N_6769);
xnor U7048 (N_7048,N_6607,N_6564);
or U7049 (N_7049,N_6912,N_6551);
xnor U7050 (N_7050,N_6516,N_6632);
nor U7051 (N_7051,N_6587,N_6928);
nand U7052 (N_7052,N_6792,N_6671);
nor U7053 (N_7053,N_6874,N_6515);
xor U7054 (N_7054,N_6932,N_6735);
or U7055 (N_7055,N_6905,N_6707);
nor U7056 (N_7056,N_6501,N_6938);
or U7057 (N_7057,N_6870,N_6930);
or U7058 (N_7058,N_6731,N_6944);
nand U7059 (N_7059,N_6981,N_6517);
xor U7060 (N_7060,N_6907,N_6887);
nand U7061 (N_7061,N_6959,N_6768);
and U7062 (N_7062,N_6510,N_6773);
xor U7063 (N_7063,N_6684,N_6962);
or U7064 (N_7064,N_6758,N_6903);
nand U7065 (N_7065,N_6793,N_6934);
nand U7066 (N_7066,N_6610,N_6569);
or U7067 (N_7067,N_6508,N_6774);
or U7068 (N_7068,N_6789,N_6815);
nand U7069 (N_7069,N_6602,N_6936);
xor U7070 (N_7070,N_6619,N_6635);
and U7071 (N_7071,N_6800,N_6832);
and U7072 (N_7072,N_6756,N_6554);
or U7073 (N_7073,N_6827,N_6566);
xor U7074 (N_7074,N_6572,N_6629);
or U7075 (N_7075,N_6560,N_6593);
and U7076 (N_7076,N_6745,N_6750);
or U7077 (N_7077,N_6940,N_6715);
xnor U7078 (N_7078,N_6718,N_6617);
and U7079 (N_7079,N_6670,N_6910);
or U7080 (N_7080,N_6514,N_6763);
or U7081 (N_7081,N_6616,N_6775);
or U7082 (N_7082,N_6642,N_6683);
nand U7083 (N_7083,N_6770,N_6637);
or U7084 (N_7084,N_6675,N_6820);
xnor U7085 (N_7085,N_6976,N_6866);
nand U7086 (N_7086,N_6558,N_6521);
nor U7087 (N_7087,N_6737,N_6691);
nor U7088 (N_7088,N_6951,N_6581);
or U7089 (N_7089,N_6709,N_6967);
or U7090 (N_7090,N_6697,N_6714);
nand U7091 (N_7091,N_6712,N_6964);
or U7092 (N_7092,N_6808,N_6998);
nand U7093 (N_7093,N_6672,N_6623);
or U7094 (N_7094,N_6854,N_6540);
and U7095 (N_7095,N_6818,N_6502);
nand U7096 (N_7096,N_6652,N_6720);
nor U7097 (N_7097,N_6685,N_6786);
nand U7098 (N_7098,N_6876,N_6692);
xor U7099 (N_7099,N_6535,N_6994);
xnor U7100 (N_7100,N_6591,N_6857);
and U7101 (N_7101,N_6791,N_6821);
and U7102 (N_7102,N_6575,N_6641);
and U7103 (N_7103,N_6603,N_6524);
and U7104 (N_7104,N_6855,N_6590);
nor U7105 (N_7105,N_6992,N_6825);
nand U7106 (N_7106,N_6659,N_6814);
xnor U7107 (N_7107,N_6879,N_6973);
and U7108 (N_7108,N_6863,N_6664);
and U7109 (N_7109,N_6654,N_6706);
xnor U7110 (N_7110,N_6598,N_6541);
or U7111 (N_7111,N_6653,N_6717);
and U7112 (N_7112,N_6826,N_6596);
nor U7113 (N_7113,N_6668,N_6724);
and U7114 (N_7114,N_6988,N_6816);
nor U7115 (N_7115,N_6677,N_6889);
nand U7116 (N_7116,N_6828,N_6640);
nor U7117 (N_7117,N_6713,N_6842);
xor U7118 (N_7118,N_6682,N_6780);
nand U7119 (N_7119,N_6662,N_6904);
or U7120 (N_7120,N_6553,N_6996);
and U7121 (N_7121,N_6979,N_6568);
and U7122 (N_7122,N_6666,N_6759);
and U7123 (N_7123,N_6704,N_6939);
xnor U7124 (N_7124,N_6545,N_6543);
nor U7125 (N_7125,N_6946,N_6585);
xor U7126 (N_7126,N_6751,N_6977);
and U7127 (N_7127,N_6529,N_6512);
nand U7128 (N_7128,N_6987,N_6891);
nand U7129 (N_7129,N_6650,N_6710);
or U7130 (N_7130,N_6833,N_6817);
nor U7131 (N_7131,N_6911,N_6537);
and U7132 (N_7132,N_6958,N_6798);
nand U7133 (N_7133,N_6646,N_6782);
nor U7134 (N_7134,N_6813,N_6504);
nor U7135 (N_7135,N_6563,N_6628);
nand U7136 (N_7136,N_6890,N_6582);
and U7137 (N_7137,N_6639,N_6941);
nor U7138 (N_7138,N_6539,N_6990);
or U7139 (N_7139,N_6971,N_6908);
nor U7140 (N_7140,N_6732,N_6937);
nand U7141 (N_7141,N_6736,N_6609);
and U7142 (N_7142,N_6614,N_6895);
nand U7143 (N_7143,N_6893,N_6807);
xnor U7144 (N_7144,N_6738,N_6506);
and U7145 (N_7145,N_6779,N_6700);
and U7146 (N_7146,N_6573,N_6550);
or U7147 (N_7147,N_6667,N_6708);
and U7148 (N_7148,N_6785,N_6942);
or U7149 (N_7149,N_6761,N_6588);
nor U7150 (N_7150,N_6755,N_6943);
or U7151 (N_7151,N_6999,N_6880);
and U7152 (N_7152,N_6766,N_6678);
xnor U7153 (N_7153,N_6845,N_6754);
nor U7154 (N_7154,N_6892,N_6565);
xnor U7155 (N_7155,N_6651,N_6841);
and U7156 (N_7156,N_6975,N_6824);
or U7157 (N_7157,N_6984,N_6723);
nand U7158 (N_7158,N_6947,N_6729);
or U7159 (N_7159,N_6838,N_6624);
and U7160 (N_7160,N_6913,N_6993);
nand U7161 (N_7161,N_6753,N_6995);
and U7162 (N_7162,N_6955,N_6850);
nand U7163 (N_7163,N_6592,N_6871);
nor U7164 (N_7164,N_6621,N_6812);
or U7165 (N_7165,N_6918,N_6836);
nand U7166 (N_7166,N_6847,N_6705);
xnor U7167 (N_7167,N_6665,N_6549);
nor U7168 (N_7168,N_6511,N_6599);
or U7169 (N_7169,N_6719,N_6746);
xnor U7170 (N_7170,N_6586,N_6949);
xnor U7171 (N_7171,N_6698,N_6505);
nor U7172 (N_7172,N_6991,N_6532);
and U7173 (N_7173,N_6542,N_6526);
xnor U7174 (N_7174,N_6853,N_6795);
and U7175 (N_7175,N_6881,N_6648);
nor U7176 (N_7176,N_6945,N_6997);
xnor U7177 (N_7177,N_6950,N_6686);
or U7178 (N_7178,N_6690,N_6618);
nor U7179 (N_7179,N_6764,N_6601);
nand U7180 (N_7180,N_6851,N_6548);
or U7181 (N_7181,N_6525,N_6916);
nor U7182 (N_7182,N_6986,N_6983);
nand U7183 (N_7183,N_6669,N_6538);
xnor U7184 (N_7184,N_6869,N_6631);
nor U7185 (N_7185,N_6797,N_6584);
or U7186 (N_7186,N_6600,N_6931);
xor U7187 (N_7187,N_6552,N_6567);
or U7188 (N_7188,N_6663,N_6703);
nor U7189 (N_7189,N_6897,N_6819);
and U7190 (N_7190,N_6699,N_6733);
and U7191 (N_7191,N_6885,N_6896);
or U7192 (N_7192,N_6788,N_6805);
and U7193 (N_7193,N_6741,N_6605);
and U7194 (N_7194,N_6519,N_6523);
nor U7195 (N_7195,N_6676,N_6608);
or U7196 (N_7196,N_6856,N_6749);
and U7197 (N_7197,N_6884,N_6957);
or U7198 (N_7198,N_6966,N_6929);
nand U7199 (N_7199,N_6898,N_6625);
nand U7200 (N_7200,N_6693,N_6862);
or U7201 (N_7201,N_6953,N_6811);
or U7202 (N_7202,N_6919,N_6583);
nand U7203 (N_7203,N_6915,N_6500);
and U7204 (N_7204,N_6762,N_6518);
nor U7205 (N_7205,N_6794,N_6882);
or U7206 (N_7206,N_6503,N_6673);
xor U7207 (N_7207,N_6611,N_6747);
and U7208 (N_7208,N_6834,N_6589);
xnor U7209 (N_7209,N_6831,N_6771);
nand U7210 (N_7210,N_6725,N_6739);
nor U7211 (N_7211,N_6660,N_6536);
nor U7212 (N_7212,N_6875,N_6643);
xor U7213 (N_7213,N_6740,N_6921);
nand U7214 (N_7214,N_6802,N_6917);
nand U7215 (N_7215,N_6883,N_6688);
xor U7216 (N_7216,N_6528,N_6689);
and U7217 (N_7217,N_6513,N_6695);
xor U7218 (N_7218,N_6835,N_6728);
nor U7219 (N_7219,N_6925,N_6840);
xnor U7220 (N_7220,N_6578,N_6868);
nor U7221 (N_7221,N_6612,N_6604);
and U7222 (N_7222,N_6822,N_6627);
nand U7223 (N_7223,N_6894,N_6799);
nand U7224 (N_7224,N_6656,N_6787);
and U7225 (N_7225,N_6743,N_6961);
nor U7226 (N_7226,N_6804,N_6922);
or U7227 (N_7227,N_6970,N_6860);
nor U7228 (N_7228,N_6861,N_6843);
or U7229 (N_7229,N_6556,N_6595);
and U7230 (N_7230,N_6757,N_6630);
xnor U7231 (N_7231,N_6948,N_6790);
and U7232 (N_7232,N_6752,N_6574);
nor U7233 (N_7233,N_6848,N_6865);
nand U7234 (N_7234,N_6696,N_6837);
nor U7235 (N_7235,N_6954,N_6726);
nor U7236 (N_7236,N_6613,N_6645);
nand U7237 (N_7237,N_6647,N_6716);
nand U7238 (N_7238,N_6914,N_6968);
and U7239 (N_7239,N_6873,N_6974);
nand U7240 (N_7240,N_6636,N_6902);
nand U7241 (N_7241,N_6680,N_6547);
and U7242 (N_7242,N_6544,N_6781);
and U7243 (N_7243,N_6965,N_6859);
or U7244 (N_7244,N_6534,N_6634);
and U7245 (N_7245,N_6956,N_6626);
or U7246 (N_7246,N_6742,N_6597);
and U7247 (N_7247,N_6679,N_6744);
or U7248 (N_7248,N_6872,N_6777);
nand U7249 (N_7249,N_6963,N_6935);
or U7250 (N_7250,N_6847,N_6630);
nand U7251 (N_7251,N_6734,N_6912);
nor U7252 (N_7252,N_6622,N_6632);
xnor U7253 (N_7253,N_6693,N_6562);
and U7254 (N_7254,N_6976,N_6863);
nor U7255 (N_7255,N_6907,N_6903);
nand U7256 (N_7256,N_6857,N_6649);
or U7257 (N_7257,N_6909,N_6782);
or U7258 (N_7258,N_6654,N_6894);
or U7259 (N_7259,N_6959,N_6549);
xor U7260 (N_7260,N_6879,N_6759);
or U7261 (N_7261,N_6896,N_6519);
and U7262 (N_7262,N_6873,N_6965);
and U7263 (N_7263,N_6777,N_6916);
and U7264 (N_7264,N_6701,N_6668);
nor U7265 (N_7265,N_6636,N_6663);
xor U7266 (N_7266,N_6937,N_6500);
nand U7267 (N_7267,N_6610,N_6681);
nor U7268 (N_7268,N_6896,N_6602);
and U7269 (N_7269,N_6861,N_6605);
nand U7270 (N_7270,N_6669,N_6923);
or U7271 (N_7271,N_6716,N_6825);
and U7272 (N_7272,N_6808,N_6791);
and U7273 (N_7273,N_6836,N_6971);
nor U7274 (N_7274,N_6909,N_6881);
nand U7275 (N_7275,N_6547,N_6642);
and U7276 (N_7276,N_6958,N_6775);
nand U7277 (N_7277,N_6749,N_6710);
nor U7278 (N_7278,N_6967,N_6835);
and U7279 (N_7279,N_6900,N_6520);
xor U7280 (N_7280,N_6616,N_6643);
nand U7281 (N_7281,N_6894,N_6725);
or U7282 (N_7282,N_6776,N_6598);
nand U7283 (N_7283,N_6940,N_6705);
and U7284 (N_7284,N_6854,N_6534);
nand U7285 (N_7285,N_6541,N_6791);
nor U7286 (N_7286,N_6652,N_6666);
and U7287 (N_7287,N_6567,N_6512);
and U7288 (N_7288,N_6598,N_6536);
xor U7289 (N_7289,N_6955,N_6708);
or U7290 (N_7290,N_6749,N_6610);
or U7291 (N_7291,N_6636,N_6882);
or U7292 (N_7292,N_6923,N_6551);
nand U7293 (N_7293,N_6668,N_6795);
or U7294 (N_7294,N_6601,N_6660);
or U7295 (N_7295,N_6529,N_6504);
nor U7296 (N_7296,N_6743,N_6522);
or U7297 (N_7297,N_6901,N_6603);
nand U7298 (N_7298,N_6865,N_6585);
nor U7299 (N_7299,N_6667,N_6566);
and U7300 (N_7300,N_6574,N_6508);
xor U7301 (N_7301,N_6558,N_6643);
or U7302 (N_7302,N_6706,N_6549);
xnor U7303 (N_7303,N_6804,N_6807);
xor U7304 (N_7304,N_6653,N_6548);
and U7305 (N_7305,N_6552,N_6848);
or U7306 (N_7306,N_6968,N_6944);
nor U7307 (N_7307,N_6539,N_6511);
nand U7308 (N_7308,N_6968,N_6792);
and U7309 (N_7309,N_6549,N_6625);
nor U7310 (N_7310,N_6530,N_6748);
or U7311 (N_7311,N_6682,N_6633);
xnor U7312 (N_7312,N_6578,N_6635);
nor U7313 (N_7313,N_6565,N_6863);
xor U7314 (N_7314,N_6564,N_6594);
nand U7315 (N_7315,N_6844,N_6989);
or U7316 (N_7316,N_6564,N_6934);
nor U7317 (N_7317,N_6569,N_6597);
xnor U7318 (N_7318,N_6842,N_6554);
and U7319 (N_7319,N_6766,N_6890);
and U7320 (N_7320,N_6717,N_6767);
nor U7321 (N_7321,N_6764,N_6998);
xor U7322 (N_7322,N_6870,N_6750);
xor U7323 (N_7323,N_6909,N_6527);
nand U7324 (N_7324,N_6746,N_6745);
nor U7325 (N_7325,N_6932,N_6827);
xor U7326 (N_7326,N_6770,N_6644);
nor U7327 (N_7327,N_6508,N_6780);
nor U7328 (N_7328,N_6980,N_6836);
and U7329 (N_7329,N_6641,N_6584);
nor U7330 (N_7330,N_6508,N_6789);
nor U7331 (N_7331,N_6897,N_6636);
nor U7332 (N_7332,N_6759,N_6825);
nor U7333 (N_7333,N_6892,N_6528);
or U7334 (N_7334,N_6591,N_6578);
nand U7335 (N_7335,N_6618,N_6793);
xnor U7336 (N_7336,N_6757,N_6883);
and U7337 (N_7337,N_6978,N_6702);
xnor U7338 (N_7338,N_6565,N_6726);
nand U7339 (N_7339,N_6774,N_6666);
nand U7340 (N_7340,N_6995,N_6792);
nand U7341 (N_7341,N_6685,N_6824);
xor U7342 (N_7342,N_6920,N_6965);
nor U7343 (N_7343,N_6568,N_6667);
nand U7344 (N_7344,N_6720,N_6951);
or U7345 (N_7345,N_6705,N_6570);
or U7346 (N_7346,N_6871,N_6887);
or U7347 (N_7347,N_6558,N_6800);
and U7348 (N_7348,N_6792,N_6593);
nand U7349 (N_7349,N_6773,N_6693);
xor U7350 (N_7350,N_6720,N_6859);
xnor U7351 (N_7351,N_6899,N_6863);
or U7352 (N_7352,N_6646,N_6568);
or U7353 (N_7353,N_6671,N_6974);
or U7354 (N_7354,N_6540,N_6822);
xor U7355 (N_7355,N_6771,N_6539);
nand U7356 (N_7356,N_6753,N_6559);
and U7357 (N_7357,N_6586,N_6791);
nand U7358 (N_7358,N_6819,N_6658);
and U7359 (N_7359,N_6620,N_6672);
or U7360 (N_7360,N_6662,N_6816);
xor U7361 (N_7361,N_6967,N_6983);
nor U7362 (N_7362,N_6769,N_6532);
xnor U7363 (N_7363,N_6683,N_6685);
and U7364 (N_7364,N_6745,N_6935);
nor U7365 (N_7365,N_6823,N_6701);
nor U7366 (N_7366,N_6920,N_6839);
nand U7367 (N_7367,N_6567,N_6533);
xnor U7368 (N_7368,N_6713,N_6738);
nand U7369 (N_7369,N_6707,N_6585);
nand U7370 (N_7370,N_6696,N_6634);
and U7371 (N_7371,N_6621,N_6560);
nor U7372 (N_7372,N_6903,N_6884);
or U7373 (N_7373,N_6938,N_6910);
and U7374 (N_7374,N_6771,N_6577);
xnor U7375 (N_7375,N_6626,N_6649);
nand U7376 (N_7376,N_6959,N_6973);
nor U7377 (N_7377,N_6739,N_6709);
nand U7378 (N_7378,N_6949,N_6547);
nor U7379 (N_7379,N_6798,N_6594);
xor U7380 (N_7380,N_6789,N_6818);
and U7381 (N_7381,N_6992,N_6878);
xor U7382 (N_7382,N_6773,N_6623);
xnor U7383 (N_7383,N_6595,N_6955);
or U7384 (N_7384,N_6994,N_6610);
or U7385 (N_7385,N_6516,N_6593);
nor U7386 (N_7386,N_6802,N_6923);
or U7387 (N_7387,N_6923,N_6874);
nor U7388 (N_7388,N_6667,N_6510);
and U7389 (N_7389,N_6901,N_6575);
and U7390 (N_7390,N_6799,N_6535);
nor U7391 (N_7391,N_6969,N_6581);
xnor U7392 (N_7392,N_6888,N_6872);
nand U7393 (N_7393,N_6673,N_6812);
and U7394 (N_7394,N_6885,N_6630);
nand U7395 (N_7395,N_6847,N_6720);
or U7396 (N_7396,N_6756,N_6694);
xor U7397 (N_7397,N_6734,N_6989);
or U7398 (N_7398,N_6840,N_6799);
nor U7399 (N_7399,N_6806,N_6925);
nor U7400 (N_7400,N_6723,N_6941);
or U7401 (N_7401,N_6657,N_6800);
xnor U7402 (N_7402,N_6567,N_6853);
xnor U7403 (N_7403,N_6919,N_6701);
nand U7404 (N_7404,N_6515,N_6924);
and U7405 (N_7405,N_6845,N_6521);
xor U7406 (N_7406,N_6645,N_6558);
nor U7407 (N_7407,N_6757,N_6528);
or U7408 (N_7408,N_6976,N_6832);
xnor U7409 (N_7409,N_6865,N_6958);
nand U7410 (N_7410,N_6836,N_6983);
nand U7411 (N_7411,N_6590,N_6877);
nand U7412 (N_7412,N_6650,N_6619);
and U7413 (N_7413,N_6895,N_6854);
nor U7414 (N_7414,N_6587,N_6752);
and U7415 (N_7415,N_6921,N_6871);
nand U7416 (N_7416,N_6709,N_6916);
xor U7417 (N_7417,N_6649,N_6847);
or U7418 (N_7418,N_6897,N_6921);
nand U7419 (N_7419,N_6649,N_6740);
nand U7420 (N_7420,N_6653,N_6823);
xnor U7421 (N_7421,N_6866,N_6514);
xnor U7422 (N_7422,N_6813,N_6689);
nand U7423 (N_7423,N_6711,N_6692);
and U7424 (N_7424,N_6885,N_6768);
or U7425 (N_7425,N_6561,N_6723);
or U7426 (N_7426,N_6885,N_6939);
nor U7427 (N_7427,N_6540,N_6508);
or U7428 (N_7428,N_6676,N_6877);
and U7429 (N_7429,N_6549,N_6814);
nor U7430 (N_7430,N_6917,N_6729);
nand U7431 (N_7431,N_6696,N_6597);
nor U7432 (N_7432,N_6608,N_6785);
xor U7433 (N_7433,N_6829,N_6783);
nand U7434 (N_7434,N_6920,N_6690);
nand U7435 (N_7435,N_6587,N_6571);
xnor U7436 (N_7436,N_6521,N_6543);
nor U7437 (N_7437,N_6682,N_6852);
nor U7438 (N_7438,N_6892,N_6864);
nor U7439 (N_7439,N_6597,N_6854);
xnor U7440 (N_7440,N_6656,N_6582);
xor U7441 (N_7441,N_6696,N_6567);
and U7442 (N_7442,N_6802,N_6575);
nand U7443 (N_7443,N_6931,N_6745);
and U7444 (N_7444,N_6887,N_6501);
nor U7445 (N_7445,N_6905,N_6659);
or U7446 (N_7446,N_6680,N_6506);
and U7447 (N_7447,N_6733,N_6778);
nor U7448 (N_7448,N_6770,N_6831);
nor U7449 (N_7449,N_6679,N_6966);
and U7450 (N_7450,N_6914,N_6591);
and U7451 (N_7451,N_6688,N_6671);
nor U7452 (N_7452,N_6702,N_6865);
and U7453 (N_7453,N_6945,N_6733);
xnor U7454 (N_7454,N_6962,N_6733);
nand U7455 (N_7455,N_6591,N_6663);
xor U7456 (N_7456,N_6645,N_6718);
nand U7457 (N_7457,N_6845,N_6555);
and U7458 (N_7458,N_6662,N_6874);
nor U7459 (N_7459,N_6581,N_6981);
and U7460 (N_7460,N_6772,N_6780);
or U7461 (N_7461,N_6759,N_6634);
nor U7462 (N_7462,N_6591,N_6878);
nand U7463 (N_7463,N_6671,N_6944);
or U7464 (N_7464,N_6631,N_6828);
nand U7465 (N_7465,N_6833,N_6513);
nor U7466 (N_7466,N_6674,N_6737);
nor U7467 (N_7467,N_6810,N_6614);
xor U7468 (N_7468,N_6726,N_6697);
nand U7469 (N_7469,N_6628,N_6739);
nand U7470 (N_7470,N_6750,N_6909);
nand U7471 (N_7471,N_6914,N_6558);
nor U7472 (N_7472,N_6613,N_6823);
nand U7473 (N_7473,N_6958,N_6860);
or U7474 (N_7474,N_6936,N_6855);
and U7475 (N_7475,N_6651,N_6614);
nand U7476 (N_7476,N_6678,N_6936);
nor U7477 (N_7477,N_6690,N_6663);
or U7478 (N_7478,N_6734,N_6709);
xor U7479 (N_7479,N_6837,N_6830);
nor U7480 (N_7480,N_6578,N_6953);
nand U7481 (N_7481,N_6500,N_6967);
nor U7482 (N_7482,N_6708,N_6803);
or U7483 (N_7483,N_6507,N_6605);
nand U7484 (N_7484,N_6555,N_6736);
or U7485 (N_7485,N_6694,N_6948);
nor U7486 (N_7486,N_6652,N_6555);
xnor U7487 (N_7487,N_6987,N_6913);
xor U7488 (N_7488,N_6597,N_6500);
and U7489 (N_7489,N_6565,N_6629);
xnor U7490 (N_7490,N_6844,N_6589);
xnor U7491 (N_7491,N_6715,N_6787);
nor U7492 (N_7492,N_6624,N_6560);
xnor U7493 (N_7493,N_6582,N_6848);
nor U7494 (N_7494,N_6508,N_6916);
nand U7495 (N_7495,N_6743,N_6832);
and U7496 (N_7496,N_6552,N_6991);
nand U7497 (N_7497,N_6975,N_6717);
and U7498 (N_7498,N_6590,N_6979);
and U7499 (N_7499,N_6825,N_6941);
and U7500 (N_7500,N_7139,N_7138);
xor U7501 (N_7501,N_7128,N_7033);
nand U7502 (N_7502,N_7355,N_7254);
xnor U7503 (N_7503,N_7277,N_7311);
and U7504 (N_7504,N_7097,N_7253);
xnor U7505 (N_7505,N_7262,N_7270);
nand U7506 (N_7506,N_7247,N_7259);
nand U7507 (N_7507,N_7154,N_7145);
or U7508 (N_7508,N_7170,N_7172);
nand U7509 (N_7509,N_7209,N_7055);
xnor U7510 (N_7510,N_7294,N_7443);
xor U7511 (N_7511,N_7332,N_7263);
nor U7512 (N_7512,N_7059,N_7021);
nand U7513 (N_7513,N_7053,N_7383);
nor U7514 (N_7514,N_7297,N_7474);
nor U7515 (N_7515,N_7268,N_7372);
nand U7516 (N_7516,N_7119,N_7228);
nor U7517 (N_7517,N_7337,N_7168);
and U7518 (N_7518,N_7285,N_7278);
xnor U7519 (N_7519,N_7157,N_7110);
or U7520 (N_7520,N_7237,N_7213);
xor U7521 (N_7521,N_7130,N_7425);
nor U7522 (N_7522,N_7420,N_7488);
or U7523 (N_7523,N_7075,N_7256);
or U7524 (N_7524,N_7123,N_7473);
nor U7525 (N_7525,N_7409,N_7344);
nand U7526 (N_7526,N_7363,N_7476);
xor U7527 (N_7527,N_7320,N_7088);
and U7528 (N_7528,N_7431,N_7408);
xnor U7529 (N_7529,N_7229,N_7137);
or U7530 (N_7530,N_7466,N_7378);
or U7531 (N_7531,N_7177,N_7068);
or U7532 (N_7532,N_7260,N_7220);
nor U7533 (N_7533,N_7370,N_7341);
and U7534 (N_7534,N_7102,N_7005);
nor U7535 (N_7535,N_7445,N_7246);
xor U7536 (N_7536,N_7233,N_7191);
and U7537 (N_7537,N_7339,N_7205);
xnor U7538 (N_7538,N_7389,N_7090);
nor U7539 (N_7539,N_7415,N_7452);
xnor U7540 (N_7540,N_7018,N_7424);
and U7541 (N_7541,N_7351,N_7221);
nor U7542 (N_7542,N_7036,N_7173);
nor U7543 (N_7543,N_7313,N_7083);
nand U7544 (N_7544,N_7106,N_7045);
and U7545 (N_7545,N_7103,N_7180);
and U7546 (N_7546,N_7164,N_7171);
and U7547 (N_7547,N_7096,N_7052);
and U7548 (N_7548,N_7034,N_7468);
xnor U7549 (N_7549,N_7000,N_7039);
nor U7550 (N_7550,N_7235,N_7010);
xor U7551 (N_7551,N_7366,N_7276);
xor U7552 (N_7552,N_7250,N_7151);
or U7553 (N_7553,N_7141,N_7491);
nand U7554 (N_7554,N_7025,N_7219);
nand U7555 (N_7555,N_7477,N_7426);
xor U7556 (N_7556,N_7436,N_7248);
or U7557 (N_7557,N_7046,N_7117);
xnor U7558 (N_7558,N_7307,N_7062);
xor U7559 (N_7559,N_7072,N_7416);
xor U7560 (N_7560,N_7079,N_7331);
or U7561 (N_7561,N_7175,N_7043);
xor U7562 (N_7562,N_7155,N_7027);
and U7563 (N_7563,N_7441,N_7356);
nor U7564 (N_7564,N_7190,N_7298);
xor U7565 (N_7565,N_7413,N_7342);
nor U7566 (N_7566,N_7126,N_7293);
nand U7567 (N_7567,N_7115,N_7368);
or U7568 (N_7568,N_7401,N_7350);
nand U7569 (N_7569,N_7377,N_7004);
xnor U7570 (N_7570,N_7086,N_7183);
xor U7571 (N_7571,N_7391,N_7269);
nand U7572 (N_7572,N_7241,N_7029);
xnor U7573 (N_7573,N_7357,N_7159);
nand U7574 (N_7574,N_7349,N_7174);
nor U7575 (N_7575,N_7487,N_7129);
and U7576 (N_7576,N_7133,N_7214);
or U7577 (N_7577,N_7390,N_7201);
nor U7578 (N_7578,N_7020,N_7371);
xor U7579 (N_7579,N_7442,N_7003);
nand U7580 (N_7580,N_7189,N_7230);
nor U7581 (N_7581,N_7279,N_7380);
and U7582 (N_7582,N_7317,N_7135);
xor U7583 (N_7583,N_7042,N_7116);
nor U7584 (N_7584,N_7404,N_7185);
or U7585 (N_7585,N_7153,N_7472);
nor U7586 (N_7586,N_7440,N_7244);
and U7587 (N_7587,N_7218,N_7446);
nor U7588 (N_7588,N_7496,N_7319);
xnor U7589 (N_7589,N_7362,N_7121);
or U7590 (N_7590,N_7300,N_7343);
or U7591 (N_7591,N_7322,N_7194);
nand U7592 (N_7592,N_7315,N_7176);
and U7593 (N_7593,N_7384,N_7124);
nor U7594 (N_7594,N_7225,N_7435);
xor U7595 (N_7595,N_7376,N_7217);
and U7596 (N_7596,N_7463,N_7108);
nand U7597 (N_7597,N_7202,N_7193);
nand U7598 (N_7598,N_7026,N_7295);
nor U7599 (N_7599,N_7136,N_7063);
and U7600 (N_7600,N_7287,N_7469);
or U7601 (N_7601,N_7458,N_7333);
xor U7602 (N_7602,N_7481,N_7492);
xor U7603 (N_7603,N_7249,N_7456);
xor U7604 (N_7604,N_7134,N_7016);
or U7605 (N_7605,N_7299,N_7432);
nand U7606 (N_7606,N_7467,N_7184);
xnor U7607 (N_7607,N_7284,N_7210);
nand U7608 (N_7608,N_7077,N_7140);
nor U7609 (N_7609,N_7447,N_7231);
or U7610 (N_7610,N_7082,N_7281);
nand U7611 (N_7611,N_7316,N_7251);
nand U7612 (N_7612,N_7358,N_7289);
and U7613 (N_7613,N_7165,N_7092);
nor U7614 (N_7614,N_7014,N_7282);
and U7615 (N_7615,N_7204,N_7245);
and U7616 (N_7616,N_7464,N_7132);
nor U7617 (N_7617,N_7179,N_7147);
nand U7618 (N_7618,N_7169,N_7008);
nor U7619 (N_7619,N_7149,N_7273);
nand U7620 (N_7620,N_7433,N_7489);
nor U7621 (N_7621,N_7483,N_7069);
nand U7622 (N_7622,N_7450,N_7242);
nand U7623 (N_7623,N_7255,N_7122);
nor U7624 (N_7624,N_7001,N_7470);
nor U7625 (N_7625,N_7482,N_7111);
nand U7626 (N_7626,N_7475,N_7291);
or U7627 (N_7627,N_7310,N_7051);
nand U7628 (N_7628,N_7375,N_7054);
xnor U7629 (N_7629,N_7038,N_7002);
nor U7630 (N_7630,N_7288,N_7381);
xnor U7631 (N_7631,N_7261,N_7037);
nand U7632 (N_7632,N_7178,N_7076);
nand U7633 (N_7633,N_7089,N_7335);
nor U7634 (N_7634,N_7336,N_7462);
or U7635 (N_7635,N_7144,N_7486);
and U7636 (N_7636,N_7098,N_7421);
nand U7637 (N_7637,N_7419,N_7120);
and U7638 (N_7638,N_7305,N_7150);
or U7639 (N_7639,N_7146,N_7417);
or U7640 (N_7640,N_7405,N_7498);
nor U7641 (N_7641,N_7353,N_7074);
nand U7642 (N_7642,N_7394,N_7334);
and U7643 (N_7643,N_7427,N_7023);
nor U7644 (N_7644,N_7304,N_7329);
or U7645 (N_7645,N_7104,N_7465);
nor U7646 (N_7646,N_7444,N_7430);
xnor U7647 (N_7647,N_7346,N_7402);
or U7648 (N_7648,N_7114,N_7407);
and U7649 (N_7649,N_7067,N_7275);
xnor U7650 (N_7650,N_7418,N_7318);
and U7651 (N_7651,N_7412,N_7187);
and U7652 (N_7652,N_7095,N_7049);
nand U7653 (N_7653,N_7406,N_7495);
or U7654 (N_7654,N_7028,N_7196);
xor U7655 (N_7655,N_7094,N_7107);
and U7656 (N_7656,N_7397,N_7118);
xnor U7657 (N_7657,N_7499,N_7301);
nor U7658 (N_7658,N_7267,N_7238);
and U7659 (N_7659,N_7453,N_7112);
or U7660 (N_7660,N_7080,N_7490);
xor U7661 (N_7661,N_7099,N_7274);
xor U7662 (N_7662,N_7485,N_7188);
nor U7663 (N_7663,N_7057,N_7031);
and U7664 (N_7664,N_7239,N_7439);
nor U7665 (N_7665,N_7266,N_7222);
nor U7666 (N_7666,N_7379,N_7399);
or U7667 (N_7667,N_7302,N_7422);
or U7668 (N_7668,N_7367,N_7073);
and U7669 (N_7669,N_7484,N_7497);
and U7670 (N_7670,N_7360,N_7236);
and U7671 (N_7671,N_7131,N_7041);
nor U7672 (N_7672,N_7388,N_7087);
nor U7673 (N_7673,N_7065,N_7460);
xnor U7674 (N_7674,N_7398,N_7015);
and U7675 (N_7675,N_7182,N_7395);
and U7676 (N_7676,N_7286,N_7454);
and U7677 (N_7677,N_7451,N_7265);
nor U7678 (N_7678,N_7032,N_7226);
or U7679 (N_7679,N_7100,N_7438);
xor U7680 (N_7680,N_7414,N_7227);
and U7681 (N_7681,N_7243,N_7060);
and U7682 (N_7682,N_7428,N_7324);
nor U7683 (N_7683,N_7396,N_7400);
and U7684 (N_7684,N_7006,N_7264);
nor U7685 (N_7685,N_7163,N_7423);
nor U7686 (N_7686,N_7312,N_7361);
xor U7687 (N_7687,N_7314,N_7048);
nor U7688 (N_7688,N_7017,N_7078);
nand U7689 (N_7689,N_7479,N_7009);
and U7690 (N_7690,N_7461,N_7125);
xor U7691 (N_7691,N_7035,N_7208);
and U7692 (N_7692,N_7061,N_7434);
nand U7693 (N_7693,N_7056,N_7162);
nor U7694 (N_7694,N_7365,N_7385);
nand U7695 (N_7695,N_7448,N_7411);
and U7696 (N_7696,N_7364,N_7203);
xnor U7697 (N_7697,N_7321,N_7013);
xnor U7698 (N_7698,N_7166,N_7308);
xnor U7699 (N_7699,N_7197,N_7303);
nor U7700 (N_7700,N_7403,N_7296);
nor U7701 (N_7701,N_7340,N_7181);
nor U7702 (N_7702,N_7494,N_7240);
and U7703 (N_7703,N_7345,N_7216);
xnor U7704 (N_7704,N_7410,N_7148);
or U7705 (N_7705,N_7352,N_7471);
or U7706 (N_7706,N_7030,N_7212);
xor U7707 (N_7707,N_7093,N_7323);
nand U7708 (N_7708,N_7186,N_7058);
nor U7709 (N_7709,N_7455,N_7457);
or U7710 (N_7710,N_7022,N_7347);
nor U7711 (N_7711,N_7195,N_7393);
and U7712 (N_7712,N_7234,N_7387);
nand U7713 (N_7713,N_7429,N_7480);
nor U7714 (N_7714,N_7354,N_7338);
nand U7715 (N_7715,N_7306,N_7200);
and U7716 (N_7716,N_7105,N_7493);
and U7717 (N_7717,N_7252,N_7206);
or U7718 (N_7718,N_7101,N_7192);
nand U7719 (N_7719,N_7066,N_7437);
and U7720 (N_7720,N_7326,N_7271);
nor U7721 (N_7721,N_7084,N_7327);
or U7722 (N_7722,N_7330,N_7386);
nor U7723 (N_7723,N_7071,N_7007);
nor U7724 (N_7724,N_7109,N_7143);
or U7725 (N_7725,N_7127,N_7374);
and U7726 (N_7726,N_7283,N_7478);
nand U7727 (N_7727,N_7359,N_7224);
or U7728 (N_7728,N_7091,N_7160);
xnor U7729 (N_7729,N_7309,N_7348);
xnor U7730 (N_7730,N_7198,N_7019);
nand U7731 (N_7731,N_7369,N_7272);
nor U7732 (N_7732,N_7156,N_7373);
nor U7733 (N_7733,N_7158,N_7012);
and U7734 (N_7734,N_7449,N_7211);
nand U7735 (N_7735,N_7290,N_7392);
nand U7736 (N_7736,N_7257,N_7113);
xor U7737 (N_7737,N_7070,N_7085);
or U7738 (N_7738,N_7024,N_7050);
or U7739 (N_7739,N_7199,N_7292);
nor U7740 (N_7740,N_7325,N_7215);
xnor U7741 (N_7741,N_7081,N_7223);
and U7742 (N_7742,N_7232,N_7040);
and U7743 (N_7743,N_7152,N_7011);
or U7744 (N_7744,N_7258,N_7167);
nor U7745 (N_7745,N_7064,N_7161);
or U7746 (N_7746,N_7328,N_7459);
and U7747 (N_7747,N_7044,N_7382);
and U7748 (N_7748,N_7207,N_7047);
nand U7749 (N_7749,N_7280,N_7142);
and U7750 (N_7750,N_7257,N_7040);
nand U7751 (N_7751,N_7365,N_7404);
xor U7752 (N_7752,N_7062,N_7140);
or U7753 (N_7753,N_7336,N_7377);
and U7754 (N_7754,N_7363,N_7079);
nor U7755 (N_7755,N_7088,N_7008);
nor U7756 (N_7756,N_7187,N_7011);
xor U7757 (N_7757,N_7020,N_7394);
xnor U7758 (N_7758,N_7231,N_7043);
xor U7759 (N_7759,N_7490,N_7295);
or U7760 (N_7760,N_7237,N_7107);
nand U7761 (N_7761,N_7347,N_7494);
nand U7762 (N_7762,N_7288,N_7184);
nand U7763 (N_7763,N_7000,N_7108);
xor U7764 (N_7764,N_7174,N_7340);
nor U7765 (N_7765,N_7267,N_7070);
and U7766 (N_7766,N_7022,N_7248);
or U7767 (N_7767,N_7056,N_7028);
or U7768 (N_7768,N_7215,N_7076);
and U7769 (N_7769,N_7098,N_7226);
and U7770 (N_7770,N_7439,N_7175);
nand U7771 (N_7771,N_7062,N_7163);
xor U7772 (N_7772,N_7180,N_7241);
xnor U7773 (N_7773,N_7193,N_7359);
xnor U7774 (N_7774,N_7333,N_7129);
nor U7775 (N_7775,N_7309,N_7105);
nand U7776 (N_7776,N_7454,N_7089);
nor U7777 (N_7777,N_7034,N_7473);
nand U7778 (N_7778,N_7114,N_7212);
or U7779 (N_7779,N_7080,N_7123);
or U7780 (N_7780,N_7153,N_7029);
xnor U7781 (N_7781,N_7393,N_7153);
and U7782 (N_7782,N_7493,N_7019);
xor U7783 (N_7783,N_7257,N_7122);
nor U7784 (N_7784,N_7202,N_7497);
and U7785 (N_7785,N_7279,N_7169);
or U7786 (N_7786,N_7212,N_7021);
xor U7787 (N_7787,N_7162,N_7498);
and U7788 (N_7788,N_7210,N_7215);
and U7789 (N_7789,N_7261,N_7258);
xor U7790 (N_7790,N_7175,N_7325);
xnor U7791 (N_7791,N_7414,N_7119);
or U7792 (N_7792,N_7329,N_7346);
nor U7793 (N_7793,N_7449,N_7217);
nor U7794 (N_7794,N_7004,N_7347);
and U7795 (N_7795,N_7479,N_7127);
xor U7796 (N_7796,N_7363,N_7029);
xor U7797 (N_7797,N_7480,N_7062);
xor U7798 (N_7798,N_7203,N_7282);
nor U7799 (N_7799,N_7177,N_7499);
nor U7800 (N_7800,N_7440,N_7114);
or U7801 (N_7801,N_7054,N_7361);
xnor U7802 (N_7802,N_7316,N_7147);
xnor U7803 (N_7803,N_7430,N_7208);
nand U7804 (N_7804,N_7121,N_7080);
xor U7805 (N_7805,N_7260,N_7464);
nor U7806 (N_7806,N_7475,N_7051);
or U7807 (N_7807,N_7309,N_7421);
xor U7808 (N_7808,N_7341,N_7192);
or U7809 (N_7809,N_7259,N_7229);
or U7810 (N_7810,N_7443,N_7001);
nand U7811 (N_7811,N_7318,N_7261);
nand U7812 (N_7812,N_7143,N_7401);
xnor U7813 (N_7813,N_7282,N_7180);
and U7814 (N_7814,N_7051,N_7219);
nor U7815 (N_7815,N_7002,N_7125);
xnor U7816 (N_7816,N_7276,N_7347);
nor U7817 (N_7817,N_7061,N_7110);
nor U7818 (N_7818,N_7415,N_7091);
or U7819 (N_7819,N_7067,N_7446);
nor U7820 (N_7820,N_7386,N_7283);
xor U7821 (N_7821,N_7082,N_7062);
nand U7822 (N_7822,N_7331,N_7464);
nor U7823 (N_7823,N_7181,N_7423);
nand U7824 (N_7824,N_7095,N_7275);
or U7825 (N_7825,N_7214,N_7048);
xor U7826 (N_7826,N_7255,N_7383);
nand U7827 (N_7827,N_7468,N_7469);
and U7828 (N_7828,N_7443,N_7243);
or U7829 (N_7829,N_7140,N_7357);
xnor U7830 (N_7830,N_7154,N_7099);
nor U7831 (N_7831,N_7326,N_7107);
nand U7832 (N_7832,N_7196,N_7103);
xor U7833 (N_7833,N_7269,N_7355);
nand U7834 (N_7834,N_7178,N_7086);
or U7835 (N_7835,N_7375,N_7168);
xnor U7836 (N_7836,N_7459,N_7449);
nor U7837 (N_7837,N_7064,N_7130);
xnor U7838 (N_7838,N_7421,N_7444);
or U7839 (N_7839,N_7309,N_7416);
and U7840 (N_7840,N_7069,N_7428);
xnor U7841 (N_7841,N_7436,N_7019);
or U7842 (N_7842,N_7413,N_7136);
and U7843 (N_7843,N_7258,N_7462);
nor U7844 (N_7844,N_7065,N_7112);
or U7845 (N_7845,N_7257,N_7477);
nor U7846 (N_7846,N_7158,N_7372);
or U7847 (N_7847,N_7079,N_7237);
xor U7848 (N_7848,N_7421,N_7402);
nand U7849 (N_7849,N_7001,N_7477);
nand U7850 (N_7850,N_7183,N_7162);
nor U7851 (N_7851,N_7414,N_7100);
nor U7852 (N_7852,N_7019,N_7483);
or U7853 (N_7853,N_7202,N_7209);
xor U7854 (N_7854,N_7228,N_7444);
and U7855 (N_7855,N_7307,N_7475);
and U7856 (N_7856,N_7242,N_7141);
xor U7857 (N_7857,N_7177,N_7141);
nor U7858 (N_7858,N_7439,N_7406);
nand U7859 (N_7859,N_7382,N_7067);
and U7860 (N_7860,N_7048,N_7177);
or U7861 (N_7861,N_7069,N_7082);
nor U7862 (N_7862,N_7081,N_7228);
xnor U7863 (N_7863,N_7015,N_7050);
xnor U7864 (N_7864,N_7049,N_7136);
xor U7865 (N_7865,N_7198,N_7238);
and U7866 (N_7866,N_7329,N_7085);
nor U7867 (N_7867,N_7141,N_7309);
nor U7868 (N_7868,N_7125,N_7147);
nand U7869 (N_7869,N_7335,N_7124);
nor U7870 (N_7870,N_7358,N_7194);
xor U7871 (N_7871,N_7439,N_7456);
nand U7872 (N_7872,N_7231,N_7429);
nor U7873 (N_7873,N_7424,N_7254);
and U7874 (N_7874,N_7072,N_7167);
and U7875 (N_7875,N_7083,N_7037);
xnor U7876 (N_7876,N_7002,N_7301);
and U7877 (N_7877,N_7456,N_7343);
and U7878 (N_7878,N_7201,N_7009);
nor U7879 (N_7879,N_7177,N_7123);
and U7880 (N_7880,N_7041,N_7388);
or U7881 (N_7881,N_7404,N_7226);
or U7882 (N_7882,N_7188,N_7415);
xor U7883 (N_7883,N_7090,N_7070);
and U7884 (N_7884,N_7118,N_7028);
or U7885 (N_7885,N_7254,N_7467);
xnor U7886 (N_7886,N_7180,N_7427);
nor U7887 (N_7887,N_7018,N_7285);
and U7888 (N_7888,N_7494,N_7056);
or U7889 (N_7889,N_7030,N_7438);
or U7890 (N_7890,N_7079,N_7376);
or U7891 (N_7891,N_7107,N_7488);
nor U7892 (N_7892,N_7407,N_7466);
and U7893 (N_7893,N_7366,N_7004);
or U7894 (N_7894,N_7307,N_7236);
and U7895 (N_7895,N_7147,N_7122);
and U7896 (N_7896,N_7114,N_7342);
xnor U7897 (N_7897,N_7123,N_7478);
nand U7898 (N_7898,N_7214,N_7456);
xor U7899 (N_7899,N_7458,N_7085);
nor U7900 (N_7900,N_7125,N_7381);
nor U7901 (N_7901,N_7415,N_7454);
xnor U7902 (N_7902,N_7349,N_7289);
and U7903 (N_7903,N_7406,N_7160);
or U7904 (N_7904,N_7306,N_7251);
and U7905 (N_7905,N_7141,N_7173);
nor U7906 (N_7906,N_7199,N_7396);
xor U7907 (N_7907,N_7494,N_7341);
nor U7908 (N_7908,N_7239,N_7419);
nand U7909 (N_7909,N_7262,N_7367);
or U7910 (N_7910,N_7134,N_7203);
nor U7911 (N_7911,N_7384,N_7235);
xnor U7912 (N_7912,N_7189,N_7181);
and U7913 (N_7913,N_7361,N_7487);
and U7914 (N_7914,N_7249,N_7303);
xnor U7915 (N_7915,N_7278,N_7166);
nand U7916 (N_7916,N_7048,N_7494);
or U7917 (N_7917,N_7434,N_7069);
xor U7918 (N_7918,N_7474,N_7276);
xor U7919 (N_7919,N_7494,N_7344);
and U7920 (N_7920,N_7245,N_7128);
nand U7921 (N_7921,N_7453,N_7270);
nor U7922 (N_7922,N_7185,N_7435);
or U7923 (N_7923,N_7268,N_7477);
xor U7924 (N_7924,N_7432,N_7104);
or U7925 (N_7925,N_7242,N_7203);
or U7926 (N_7926,N_7481,N_7266);
xnor U7927 (N_7927,N_7134,N_7244);
nor U7928 (N_7928,N_7015,N_7273);
nand U7929 (N_7929,N_7081,N_7070);
nor U7930 (N_7930,N_7303,N_7230);
or U7931 (N_7931,N_7410,N_7154);
xor U7932 (N_7932,N_7336,N_7350);
nor U7933 (N_7933,N_7094,N_7312);
xor U7934 (N_7934,N_7190,N_7426);
xor U7935 (N_7935,N_7220,N_7197);
nor U7936 (N_7936,N_7371,N_7011);
nor U7937 (N_7937,N_7216,N_7486);
nor U7938 (N_7938,N_7378,N_7341);
nor U7939 (N_7939,N_7020,N_7274);
xor U7940 (N_7940,N_7003,N_7268);
and U7941 (N_7941,N_7089,N_7279);
xnor U7942 (N_7942,N_7235,N_7128);
nor U7943 (N_7943,N_7424,N_7161);
nor U7944 (N_7944,N_7410,N_7164);
xor U7945 (N_7945,N_7281,N_7117);
nor U7946 (N_7946,N_7220,N_7173);
xnor U7947 (N_7947,N_7173,N_7385);
or U7948 (N_7948,N_7285,N_7404);
nand U7949 (N_7949,N_7312,N_7201);
xor U7950 (N_7950,N_7315,N_7299);
and U7951 (N_7951,N_7072,N_7363);
and U7952 (N_7952,N_7421,N_7063);
xnor U7953 (N_7953,N_7475,N_7241);
nor U7954 (N_7954,N_7035,N_7447);
nand U7955 (N_7955,N_7472,N_7233);
nand U7956 (N_7956,N_7031,N_7379);
and U7957 (N_7957,N_7477,N_7267);
xor U7958 (N_7958,N_7440,N_7319);
nand U7959 (N_7959,N_7182,N_7419);
xor U7960 (N_7960,N_7483,N_7096);
or U7961 (N_7961,N_7255,N_7264);
or U7962 (N_7962,N_7119,N_7256);
or U7963 (N_7963,N_7161,N_7322);
and U7964 (N_7964,N_7344,N_7152);
xnor U7965 (N_7965,N_7018,N_7482);
xor U7966 (N_7966,N_7151,N_7336);
and U7967 (N_7967,N_7374,N_7038);
or U7968 (N_7968,N_7130,N_7034);
or U7969 (N_7969,N_7230,N_7177);
or U7970 (N_7970,N_7415,N_7059);
and U7971 (N_7971,N_7065,N_7122);
or U7972 (N_7972,N_7367,N_7056);
nand U7973 (N_7973,N_7413,N_7071);
xnor U7974 (N_7974,N_7065,N_7049);
and U7975 (N_7975,N_7027,N_7140);
nor U7976 (N_7976,N_7436,N_7398);
nor U7977 (N_7977,N_7452,N_7188);
nor U7978 (N_7978,N_7059,N_7417);
or U7979 (N_7979,N_7182,N_7192);
xor U7980 (N_7980,N_7147,N_7117);
nand U7981 (N_7981,N_7151,N_7020);
and U7982 (N_7982,N_7300,N_7244);
or U7983 (N_7983,N_7257,N_7210);
and U7984 (N_7984,N_7295,N_7355);
or U7985 (N_7985,N_7278,N_7234);
and U7986 (N_7986,N_7110,N_7194);
xor U7987 (N_7987,N_7216,N_7256);
and U7988 (N_7988,N_7001,N_7485);
and U7989 (N_7989,N_7296,N_7157);
nand U7990 (N_7990,N_7301,N_7323);
xor U7991 (N_7991,N_7377,N_7158);
nor U7992 (N_7992,N_7416,N_7080);
nor U7993 (N_7993,N_7093,N_7337);
xnor U7994 (N_7994,N_7066,N_7363);
and U7995 (N_7995,N_7486,N_7045);
nand U7996 (N_7996,N_7164,N_7169);
and U7997 (N_7997,N_7116,N_7337);
nor U7998 (N_7998,N_7153,N_7422);
xnor U7999 (N_7999,N_7254,N_7239);
or U8000 (N_8000,N_7728,N_7850);
nor U8001 (N_8001,N_7524,N_7731);
or U8002 (N_8002,N_7681,N_7973);
nor U8003 (N_8003,N_7686,N_7650);
nor U8004 (N_8004,N_7675,N_7913);
xnor U8005 (N_8005,N_7941,N_7876);
xor U8006 (N_8006,N_7967,N_7857);
nor U8007 (N_8007,N_7722,N_7611);
nor U8008 (N_8008,N_7636,N_7660);
or U8009 (N_8009,N_7511,N_7923);
or U8010 (N_8010,N_7961,N_7696);
xnor U8011 (N_8011,N_7791,N_7886);
nand U8012 (N_8012,N_7826,N_7666);
or U8013 (N_8013,N_7986,N_7786);
and U8014 (N_8014,N_7796,N_7725);
or U8015 (N_8015,N_7584,N_7859);
nor U8016 (N_8016,N_7995,N_7807);
and U8017 (N_8017,N_7860,N_7614);
xnor U8018 (N_8018,N_7702,N_7901);
and U8019 (N_8019,N_7750,N_7537);
and U8020 (N_8020,N_7918,N_7867);
xnor U8021 (N_8021,N_7974,N_7762);
or U8022 (N_8022,N_7792,N_7668);
nor U8023 (N_8023,N_7872,N_7645);
nor U8024 (N_8024,N_7892,N_7620);
or U8025 (N_8025,N_7904,N_7869);
nor U8026 (N_8026,N_7753,N_7720);
nand U8027 (N_8027,N_7649,N_7861);
or U8028 (N_8028,N_7761,N_7774);
and U8029 (N_8029,N_7884,N_7990);
nand U8030 (N_8030,N_7591,N_7562);
nor U8031 (N_8031,N_7657,N_7508);
nor U8032 (N_8032,N_7570,N_7794);
nand U8033 (N_8033,N_7780,N_7933);
and U8034 (N_8034,N_7832,N_7646);
xnor U8035 (N_8035,N_7515,N_7661);
nand U8036 (N_8036,N_7671,N_7532);
nand U8037 (N_8037,N_7775,N_7669);
or U8038 (N_8038,N_7573,N_7633);
or U8039 (N_8039,N_7572,N_7838);
and U8040 (N_8040,N_7991,N_7963);
xor U8041 (N_8041,N_7896,N_7905);
xnor U8042 (N_8042,N_7536,N_7970);
or U8043 (N_8043,N_7779,N_7946);
nand U8044 (N_8044,N_7739,N_7790);
or U8045 (N_8045,N_7639,N_7531);
nand U8046 (N_8046,N_7683,N_7804);
xor U8047 (N_8047,N_7592,N_7831);
xor U8048 (N_8048,N_7556,N_7625);
and U8049 (N_8049,N_7578,N_7898);
nor U8050 (N_8050,N_7707,N_7658);
xor U8051 (N_8051,N_7679,N_7777);
xor U8052 (N_8052,N_7677,N_7959);
and U8053 (N_8053,N_7878,N_7752);
nand U8054 (N_8054,N_7512,N_7772);
nor U8055 (N_8055,N_7656,N_7648);
nand U8056 (N_8056,N_7938,N_7875);
or U8057 (N_8057,N_7841,N_7984);
nand U8058 (N_8058,N_7528,N_7929);
or U8059 (N_8059,N_7843,N_7809);
nand U8060 (N_8060,N_7533,N_7757);
nor U8061 (N_8061,N_7542,N_7758);
nor U8062 (N_8062,N_7802,N_7603);
nand U8063 (N_8063,N_7763,N_7943);
or U8064 (N_8064,N_7713,N_7516);
and U8065 (N_8065,N_7577,N_7821);
nor U8066 (N_8066,N_7834,N_7927);
or U8067 (N_8067,N_7883,N_7977);
nand U8068 (N_8068,N_7643,N_7806);
or U8069 (N_8069,N_7824,N_7672);
or U8070 (N_8070,N_7799,N_7721);
nand U8071 (N_8071,N_7699,N_7983);
xor U8072 (N_8072,N_7817,N_7694);
nor U8073 (N_8073,N_7766,N_7553);
xor U8074 (N_8074,N_7814,N_7560);
nor U8075 (N_8075,N_7971,N_7855);
nand U8076 (N_8076,N_7972,N_7659);
xor U8077 (N_8077,N_7730,N_7877);
nor U8078 (N_8078,N_7698,N_7985);
nor U8079 (N_8079,N_7632,N_7980);
xnor U8080 (N_8080,N_7685,N_7979);
nor U8081 (N_8081,N_7705,N_7820);
or U8082 (N_8082,N_7998,N_7767);
nand U8083 (N_8083,N_7823,N_7551);
or U8084 (N_8084,N_7899,N_7715);
or U8085 (N_8085,N_7842,N_7789);
nor U8086 (N_8086,N_7853,N_7552);
xnor U8087 (N_8087,N_7798,N_7764);
and U8088 (N_8088,N_7595,N_7628);
nand U8089 (N_8089,N_7561,N_7978);
nand U8090 (N_8090,N_7719,N_7637);
and U8091 (N_8091,N_7783,N_7565);
nand U8092 (N_8092,N_7816,N_7909);
xor U8093 (N_8093,N_7893,N_7960);
nand U8094 (N_8094,N_7771,N_7793);
or U8095 (N_8095,N_7541,N_7514);
nor U8096 (N_8096,N_7781,N_7534);
xor U8097 (N_8097,N_7925,N_7631);
xor U8098 (N_8098,N_7574,N_7805);
nand U8099 (N_8099,N_7760,N_7629);
nor U8100 (N_8100,N_7526,N_7689);
and U8101 (N_8101,N_7955,N_7506);
and U8102 (N_8102,N_7529,N_7638);
nand U8103 (N_8103,N_7741,N_7505);
xor U8104 (N_8104,N_7844,N_7787);
or U8105 (N_8105,N_7989,N_7969);
nand U8106 (N_8106,N_7503,N_7922);
xor U8107 (N_8107,N_7527,N_7734);
nor U8108 (N_8108,N_7510,N_7932);
xnor U8109 (N_8109,N_7885,N_7801);
nor U8110 (N_8110,N_7564,N_7743);
or U8111 (N_8111,N_7848,N_7803);
and U8112 (N_8112,N_7852,N_7641);
and U8113 (N_8113,N_7900,N_7710);
xnor U8114 (N_8114,N_7504,N_7509);
nand U8115 (N_8115,N_7653,N_7964);
xnor U8116 (N_8116,N_7676,N_7755);
and U8117 (N_8117,N_7530,N_7812);
xnor U8118 (N_8118,N_7644,N_7711);
xnor U8119 (N_8119,N_7597,N_7576);
or U8120 (N_8120,N_7695,N_7742);
or U8121 (N_8121,N_7907,N_7535);
nor U8122 (N_8122,N_7851,N_7800);
xnor U8123 (N_8123,N_7776,N_7910);
nor U8124 (N_8124,N_7630,N_7606);
or U8125 (N_8125,N_7920,N_7651);
and U8126 (N_8126,N_7879,N_7994);
nor U8127 (N_8127,N_7714,N_7616);
nand U8128 (N_8128,N_7870,N_7594);
nor U8129 (N_8129,N_7951,N_7554);
and U8130 (N_8130,N_7996,N_7997);
or U8131 (N_8131,N_7655,N_7712);
nand U8132 (N_8132,N_7667,N_7624);
or U8133 (N_8133,N_7934,N_7839);
or U8134 (N_8134,N_7881,N_7880);
or U8135 (N_8135,N_7549,N_7912);
or U8136 (N_8136,N_7559,N_7992);
xnor U8137 (N_8137,N_7873,N_7599);
and U8138 (N_8138,N_7916,N_7948);
or U8139 (N_8139,N_7682,N_7500);
xnor U8140 (N_8140,N_7962,N_7785);
and U8141 (N_8141,N_7610,N_7521);
and U8142 (N_8142,N_7735,N_7864);
and U8143 (N_8143,N_7501,N_7558);
or U8144 (N_8144,N_7618,N_7836);
and U8145 (N_8145,N_7687,N_7586);
and U8146 (N_8146,N_7949,N_7993);
or U8147 (N_8147,N_7937,N_7768);
xnor U8148 (N_8148,N_7502,N_7888);
nand U8149 (N_8149,N_7982,N_7837);
nand U8150 (N_8150,N_7727,N_7684);
or U8151 (N_8151,N_7840,N_7627);
xor U8152 (N_8152,N_7897,N_7813);
and U8153 (N_8153,N_7733,N_7664);
nand U8154 (N_8154,N_7670,N_7581);
xnor U8155 (N_8155,N_7523,N_7548);
and U8156 (N_8156,N_7706,N_7903);
nor U8157 (N_8157,N_7874,N_7751);
nor U8158 (N_8158,N_7947,N_7847);
xor U8159 (N_8159,N_7652,N_7680);
and U8160 (N_8160,N_7845,N_7691);
xor U8161 (N_8161,N_7593,N_7737);
xor U8162 (N_8162,N_7708,N_7808);
nor U8163 (N_8163,N_7538,N_7862);
nor U8164 (N_8164,N_7835,N_7745);
nand U8165 (N_8165,N_7635,N_7911);
and U8166 (N_8166,N_7674,N_7609);
nor U8167 (N_8167,N_7858,N_7583);
or U8168 (N_8168,N_7965,N_7662);
and U8169 (N_8169,N_7950,N_7988);
nor U8170 (N_8170,N_7987,N_7818);
xnor U8171 (N_8171,N_7931,N_7585);
or U8172 (N_8172,N_7975,N_7784);
nand U8173 (N_8173,N_7953,N_7582);
nand U8174 (N_8174,N_7822,N_7957);
xor U8175 (N_8175,N_7863,N_7954);
nor U8176 (N_8176,N_7895,N_7520);
nand U8177 (N_8177,N_7747,N_7738);
xnor U8178 (N_8178,N_7703,N_7543);
xnor U8179 (N_8179,N_7981,N_7507);
and U8180 (N_8180,N_7539,N_7716);
and U8181 (N_8181,N_7902,N_7830);
nand U8182 (N_8182,N_7958,N_7619);
nor U8183 (N_8183,N_7587,N_7940);
xor U8184 (N_8184,N_7939,N_7871);
nand U8185 (N_8185,N_7555,N_7588);
and U8186 (N_8186,N_7746,N_7693);
and U8187 (N_8187,N_7605,N_7640);
nand U8188 (N_8188,N_7819,N_7944);
xor U8189 (N_8189,N_7810,N_7778);
or U8190 (N_8190,N_7849,N_7976);
nor U8191 (N_8191,N_7617,N_7795);
xnor U8192 (N_8192,N_7935,N_7914);
and U8193 (N_8193,N_7765,N_7665);
and U8194 (N_8194,N_7525,N_7522);
nor U8195 (N_8195,N_7917,N_7797);
xor U8196 (N_8196,N_7908,N_7856);
nand U8197 (N_8197,N_7782,N_7740);
and U8198 (N_8198,N_7906,N_7690);
xnor U8199 (N_8199,N_7654,N_7590);
xor U8200 (N_8200,N_7546,N_7854);
xnor U8201 (N_8201,N_7865,N_7829);
nand U8202 (N_8202,N_7887,N_7846);
or U8203 (N_8203,N_7568,N_7678);
or U8204 (N_8204,N_7890,N_7601);
xnor U8205 (N_8205,N_7749,N_7602);
and U8206 (N_8206,N_7513,N_7724);
and U8207 (N_8207,N_7748,N_7868);
xnor U8208 (N_8208,N_7517,N_7701);
nand U8209 (N_8209,N_7773,N_7930);
xnor U8210 (N_8210,N_7613,N_7942);
nand U8211 (N_8211,N_7709,N_7547);
nand U8212 (N_8212,N_7770,N_7615);
xor U8213 (N_8213,N_7894,N_7999);
nor U8214 (N_8214,N_7921,N_7754);
nand U8215 (N_8215,N_7598,N_7882);
nand U8216 (N_8216,N_7544,N_7612);
nor U8217 (N_8217,N_7756,N_7634);
nand U8218 (N_8218,N_7567,N_7642);
or U8219 (N_8219,N_7688,N_7569);
and U8220 (N_8220,N_7928,N_7540);
xnor U8221 (N_8221,N_7519,N_7744);
nand U8222 (N_8222,N_7557,N_7945);
xor U8223 (N_8223,N_7604,N_7622);
and U8224 (N_8224,N_7563,N_7828);
nor U8225 (N_8225,N_7600,N_7811);
nand U8226 (N_8226,N_7956,N_7579);
or U8227 (N_8227,N_7607,N_7924);
xnor U8228 (N_8228,N_7833,N_7926);
nor U8229 (N_8229,N_7717,N_7545);
nand U8230 (N_8230,N_7673,N_7729);
or U8231 (N_8231,N_7788,N_7919);
nor U8232 (N_8232,N_7825,N_7518);
and U8233 (N_8233,N_7936,N_7732);
nand U8234 (N_8234,N_7663,N_7623);
and U8235 (N_8235,N_7815,N_7889);
xor U8236 (N_8236,N_7759,N_7608);
and U8237 (N_8237,N_7647,N_7580);
and U8238 (N_8238,N_7915,N_7697);
xor U8239 (N_8239,N_7866,N_7566);
nand U8240 (N_8240,N_7891,N_7692);
or U8241 (N_8241,N_7968,N_7626);
nor U8242 (N_8242,N_7723,N_7575);
xor U8243 (N_8243,N_7736,N_7966);
and U8244 (N_8244,N_7700,N_7596);
nand U8245 (N_8245,N_7726,N_7571);
xor U8246 (N_8246,N_7704,N_7589);
nand U8247 (N_8247,N_7952,N_7550);
nand U8248 (N_8248,N_7718,N_7769);
or U8249 (N_8249,N_7621,N_7827);
xor U8250 (N_8250,N_7756,N_7518);
and U8251 (N_8251,N_7563,N_7838);
xnor U8252 (N_8252,N_7622,N_7514);
and U8253 (N_8253,N_7671,N_7610);
nor U8254 (N_8254,N_7782,N_7918);
xor U8255 (N_8255,N_7903,N_7988);
xnor U8256 (N_8256,N_7533,N_7954);
or U8257 (N_8257,N_7578,N_7719);
and U8258 (N_8258,N_7914,N_7633);
and U8259 (N_8259,N_7966,N_7910);
or U8260 (N_8260,N_7778,N_7677);
nor U8261 (N_8261,N_7564,N_7664);
or U8262 (N_8262,N_7507,N_7994);
nor U8263 (N_8263,N_7705,N_7728);
or U8264 (N_8264,N_7645,N_7526);
nor U8265 (N_8265,N_7655,N_7762);
or U8266 (N_8266,N_7898,N_7715);
xnor U8267 (N_8267,N_7734,N_7714);
nor U8268 (N_8268,N_7628,N_7710);
xnor U8269 (N_8269,N_7857,N_7888);
xor U8270 (N_8270,N_7895,N_7757);
or U8271 (N_8271,N_7666,N_7681);
xnor U8272 (N_8272,N_7792,N_7802);
or U8273 (N_8273,N_7841,N_7588);
nand U8274 (N_8274,N_7521,N_7553);
xor U8275 (N_8275,N_7968,N_7897);
and U8276 (N_8276,N_7963,N_7874);
nand U8277 (N_8277,N_7895,N_7567);
xor U8278 (N_8278,N_7931,N_7662);
and U8279 (N_8279,N_7585,N_7818);
nor U8280 (N_8280,N_7844,N_7858);
xor U8281 (N_8281,N_7519,N_7961);
nor U8282 (N_8282,N_7575,N_7909);
or U8283 (N_8283,N_7955,N_7909);
nor U8284 (N_8284,N_7982,N_7923);
and U8285 (N_8285,N_7799,N_7976);
or U8286 (N_8286,N_7593,N_7850);
nand U8287 (N_8287,N_7896,N_7815);
nor U8288 (N_8288,N_7727,N_7861);
nand U8289 (N_8289,N_7827,N_7682);
nor U8290 (N_8290,N_7632,N_7994);
and U8291 (N_8291,N_7559,N_7607);
and U8292 (N_8292,N_7720,N_7952);
xor U8293 (N_8293,N_7806,N_7614);
nand U8294 (N_8294,N_7840,N_7749);
nand U8295 (N_8295,N_7907,N_7947);
or U8296 (N_8296,N_7962,N_7701);
nand U8297 (N_8297,N_7992,N_7803);
and U8298 (N_8298,N_7861,N_7590);
xnor U8299 (N_8299,N_7677,N_7572);
nor U8300 (N_8300,N_7679,N_7543);
nand U8301 (N_8301,N_7524,N_7606);
or U8302 (N_8302,N_7613,N_7850);
nand U8303 (N_8303,N_7656,N_7855);
or U8304 (N_8304,N_7704,N_7980);
and U8305 (N_8305,N_7630,N_7809);
nand U8306 (N_8306,N_7700,N_7693);
or U8307 (N_8307,N_7907,N_7860);
nor U8308 (N_8308,N_7848,N_7818);
and U8309 (N_8309,N_7610,N_7736);
xor U8310 (N_8310,N_7634,N_7999);
nand U8311 (N_8311,N_7752,N_7619);
nor U8312 (N_8312,N_7708,N_7549);
nand U8313 (N_8313,N_7653,N_7881);
or U8314 (N_8314,N_7662,N_7616);
nor U8315 (N_8315,N_7802,N_7806);
and U8316 (N_8316,N_7690,N_7642);
nor U8317 (N_8317,N_7829,N_7742);
or U8318 (N_8318,N_7900,N_7506);
xor U8319 (N_8319,N_7762,N_7821);
nor U8320 (N_8320,N_7950,N_7923);
and U8321 (N_8321,N_7744,N_7571);
or U8322 (N_8322,N_7855,N_7910);
or U8323 (N_8323,N_7700,N_7925);
xnor U8324 (N_8324,N_7956,N_7895);
and U8325 (N_8325,N_7678,N_7913);
or U8326 (N_8326,N_7953,N_7870);
nand U8327 (N_8327,N_7810,N_7645);
nor U8328 (N_8328,N_7701,N_7547);
and U8329 (N_8329,N_7693,N_7727);
or U8330 (N_8330,N_7930,N_7628);
or U8331 (N_8331,N_7997,N_7548);
nand U8332 (N_8332,N_7735,N_7701);
nand U8333 (N_8333,N_7604,N_7552);
nand U8334 (N_8334,N_7717,N_7797);
and U8335 (N_8335,N_7932,N_7809);
nor U8336 (N_8336,N_7609,N_7995);
and U8337 (N_8337,N_7988,N_7852);
nand U8338 (N_8338,N_7864,N_7725);
nand U8339 (N_8339,N_7595,N_7802);
or U8340 (N_8340,N_7527,N_7942);
or U8341 (N_8341,N_7743,N_7804);
xnor U8342 (N_8342,N_7770,N_7824);
nand U8343 (N_8343,N_7655,N_7553);
nor U8344 (N_8344,N_7566,N_7651);
nand U8345 (N_8345,N_7908,N_7729);
nand U8346 (N_8346,N_7989,N_7581);
nand U8347 (N_8347,N_7875,N_7850);
and U8348 (N_8348,N_7611,N_7505);
nor U8349 (N_8349,N_7875,N_7589);
and U8350 (N_8350,N_7811,N_7708);
xnor U8351 (N_8351,N_7957,N_7737);
or U8352 (N_8352,N_7757,N_7750);
nor U8353 (N_8353,N_7545,N_7692);
xnor U8354 (N_8354,N_7553,N_7729);
nor U8355 (N_8355,N_7575,N_7963);
or U8356 (N_8356,N_7610,N_7667);
or U8357 (N_8357,N_7699,N_7974);
or U8358 (N_8358,N_7713,N_7961);
nor U8359 (N_8359,N_7938,N_7978);
and U8360 (N_8360,N_7599,N_7678);
or U8361 (N_8361,N_7645,N_7793);
nand U8362 (N_8362,N_7527,N_7790);
or U8363 (N_8363,N_7606,N_7771);
nand U8364 (N_8364,N_7849,N_7615);
nor U8365 (N_8365,N_7998,N_7808);
xor U8366 (N_8366,N_7828,N_7676);
nand U8367 (N_8367,N_7576,N_7569);
nand U8368 (N_8368,N_7964,N_7905);
and U8369 (N_8369,N_7856,N_7888);
xnor U8370 (N_8370,N_7689,N_7646);
nor U8371 (N_8371,N_7658,N_7642);
xnor U8372 (N_8372,N_7623,N_7845);
and U8373 (N_8373,N_7949,N_7685);
nor U8374 (N_8374,N_7793,N_7529);
nor U8375 (N_8375,N_7821,N_7845);
or U8376 (N_8376,N_7557,N_7724);
xnor U8377 (N_8377,N_7788,N_7671);
xnor U8378 (N_8378,N_7558,N_7605);
nand U8379 (N_8379,N_7570,N_7733);
nand U8380 (N_8380,N_7999,N_7744);
nor U8381 (N_8381,N_7943,N_7818);
and U8382 (N_8382,N_7679,N_7758);
or U8383 (N_8383,N_7620,N_7555);
xnor U8384 (N_8384,N_7885,N_7908);
nand U8385 (N_8385,N_7592,N_7838);
nor U8386 (N_8386,N_7874,N_7695);
and U8387 (N_8387,N_7566,N_7613);
or U8388 (N_8388,N_7748,N_7959);
or U8389 (N_8389,N_7829,N_7918);
or U8390 (N_8390,N_7518,N_7885);
nand U8391 (N_8391,N_7871,N_7878);
nor U8392 (N_8392,N_7558,N_7640);
or U8393 (N_8393,N_7936,N_7780);
nand U8394 (N_8394,N_7574,N_7629);
nor U8395 (N_8395,N_7519,N_7705);
or U8396 (N_8396,N_7712,N_7611);
nand U8397 (N_8397,N_7939,N_7563);
nor U8398 (N_8398,N_7509,N_7840);
xor U8399 (N_8399,N_7717,N_7895);
or U8400 (N_8400,N_7978,N_7808);
nand U8401 (N_8401,N_7522,N_7698);
and U8402 (N_8402,N_7789,N_7705);
nand U8403 (N_8403,N_7716,N_7964);
xnor U8404 (N_8404,N_7706,N_7518);
or U8405 (N_8405,N_7934,N_7559);
nor U8406 (N_8406,N_7756,N_7747);
xnor U8407 (N_8407,N_7652,N_7887);
xnor U8408 (N_8408,N_7505,N_7736);
nand U8409 (N_8409,N_7742,N_7853);
nand U8410 (N_8410,N_7913,N_7942);
or U8411 (N_8411,N_7657,N_7933);
xor U8412 (N_8412,N_7569,N_7783);
nand U8413 (N_8413,N_7608,N_7829);
and U8414 (N_8414,N_7500,N_7821);
nand U8415 (N_8415,N_7554,N_7625);
xor U8416 (N_8416,N_7756,N_7615);
xor U8417 (N_8417,N_7809,N_7705);
nor U8418 (N_8418,N_7692,N_7634);
or U8419 (N_8419,N_7503,N_7550);
and U8420 (N_8420,N_7845,N_7897);
or U8421 (N_8421,N_7939,N_7868);
and U8422 (N_8422,N_7594,N_7587);
or U8423 (N_8423,N_7839,N_7917);
and U8424 (N_8424,N_7632,N_7959);
and U8425 (N_8425,N_7616,N_7533);
nand U8426 (N_8426,N_7746,N_7776);
nor U8427 (N_8427,N_7697,N_7983);
nor U8428 (N_8428,N_7565,N_7811);
or U8429 (N_8429,N_7916,N_7865);
nor U8430 (N_8430,N_7720,N_7680);
xnor U8431 (N_8431,N_7540,N_7813);
nand U8432 (N_8432,N_7556,N_7846);
or U8433 (N_8433,N_7821,N_7501);
nand U8434 (N_8434,N_7852,N_7507);
and U8435 (N_8435,N_7759,N_7964);
nand U8436 (N_8436,N_7587,N_7961);
and U8437 (N_8437,N_7977,N_7831);
nand U8438 (N_8438,N_7728,N_7646);
xnor U8439 (N_8439,N_7762,N_7532);
nand U8440 (N_8440,N_7711,N_7918);
or U8441 (N_8441,N_7987,N_7682);
or U8442 (N_8442,N_7526,N_7866);
nand U8443 (N_8443,N_7595,N_7571);
or U8444 (N_8444,N_7502,N_7742);
nand U8445 (N_8445,N_7844,N_7603);
or U8446 (N_8446,N_7957,N_7754);
and U8447 (N_8447,N_7938,N_7593);
xor U8448 (N_8448,N_7666,N_7602);
or U8449 (N_8449,N_7841,N_7983);
or U8450 (N_8450,N_7758,N_7911);
xnor U8451 (N_8451,N_7685,N_7782);
and U8452 (N_8452,N_7683,N_7668);
nor U8453 (N_8453,N_7890,N_7558);
xnor U8454 (N_8454,N_7832,N_7864);
nand U8455 (N_8455,N_7990,N_7720);
xor U8456 (N_8456,N_7932,N_7863);
nand U8457 (N_8457,N_7875,N_7984);
and U8458 (N_8458,N_7655,N_7754);
and U8459 (N_8459,N_7553,N_7625);
nor U8460 (N_8460,N_7578,N_7664);
nor U8461 (N_8461,N_7538,N_7767);
nor U8462 (N_8462,N_7779,N_7959);
nor U8463 (N_8463,N_7541,N_7691);
and U8464 (N_8464,N_7907,N_7810);
or U8465 (N_8465,N_7608,N_7748);
nand U8466 (N_8466,N_7703,N_7943);
nand U8467 (N_8467,N_7955,N_7714);
nor U8468 (N_8468,N_7539,N_7909);
xor U8469 (N_8469,N_7907,N_7511);
and U8470 (N_8470,N_7953,N_7924);
and U8471 (N_8471,N_7764,N_7929);
xor U8472 (N_8472,N_7543,N_7992);
nor U8473 (N_8473,N_7843,N_7770);
nand U8474 (N_8474,N_7957,N_7949);
and U8475 (N_8475,N_7515,N_7898);
xor U8476 (N_8476,N_7580,N_7872);
nand U8477 (N_8477,N_7688,N_7942);
nand U8478 (N_8478,N_7538,N_7895);
nand U8479 (N_8479,N_7928,N_7611);
xnor U8480 (N_8480,N_7922,N_7662);
xor U8481 (N_8481,N_7758,N_7768);
or U8482 (N_8482,N_7539,N_7886);
nor U8483 (N_8483,N_7647,N_7584);
and U8484 (N_8484,N_7959,N_7769);
or U8485 (N_8485,N_7956,N_7767);
nand U8486 (N_8486,N_7615,N_7739);
and U8487 (N_8487,N_7610,N_7987);
and U8488 (N_8488,N_7834,N_7887);
xor U8489 (N_8489,N_7753,N_7739);
nand U8490 (N_8490,N_7857,N_7625);
and U8491 (N_8491,N_7826,N_7600);
nand U8492 (N_8492,N_7633,N_7930);
xor U8493 (N_8493,N_7685,N_7845);
xnor U8494 (N_8494,N_7599,N_7577);
or U8495 (N_8495,N_7712,N_7797);
xor U8496 (N_8496,N_7824,N_7613);
or U8497 (N_8497,N_7958,N_7779);
and U8498 (N_8498,N_7567,N_7600);
nand U8499 (N_8499,N_7824,N_7793);
nand U8500 (N_8500,N_8456,N_8286);
nor U8501 (N_8501,N_8100,N_8126);
nand U8502 (N_8502,N_8311,N_8047);
xor U8503 (N_8503,N_8184,N_8307);
xnor U8504 (N_8504,N_8165,N_8380);
or U8505 (N_8505,N_8221,N_8331);
and U8506 (N_8506,N_8214,N_8472);
or U8507 (N_8507,N_8190,N_8270);
nor U8508 (N_8508,N_8245,N_8243);
nand U8509 (N_8509,N_8082,N_8309);
nor U8510 (N_8510,N_8316,N_8239);
xor U8511 (N_8511,N_8088,N_8241);
nor U8512 (N_8512,N_8223,N_8193);
xor U8513 (N_8513,N_8199,N_8091);
nand U8514 (N_8514,N_8228,N_8012);
or U8515 (N_8515,N_8202,N_8115);
nor U8516 (N_8516,N_8086,N_8098);
xor U8517 (N_8517,N_8068,N_8256);
and U8518 (N_8518,N_8060,N_8341);
or U8519 (N_8519,N_8368,N_8417);
nand U8520 (N_8520,N_8322,N_8011);
xnor U8521 (N_8521,N_8033,N_8325);
nor U8522 (N_8522,N_8035,N_8030);
or U8523 (N_8523,N_8053,N_8477);
nand U8524 (N_8524,N_8216,N_8394);
xor U8525 (N_8525,N_8399,N_8273);
nand U8526 (N_8526,N_8112,N_8017);
nand U8527 (N_8527,N_8269,N_8428);
xor U8528 (N_8528,N_8015,N_8031);
and U8529 (N_8529,N_8084,N_8484);
or U8530 (N_8530,N_8146,N_8281);
and U8531 (N_8531,N_8094,N_8087);
nand U8532 (N_8532,N_8234,N_8345);
or U8533 (N_8533,N_8054,N_8395);
or U8534 (N_8534,N_8426,N_8267);
xor U8535 (N_8535,N_8268,N_8419);
nand U8536 (N_8536,N_8160,N_8324);
nand U8537 (N_8537,N_8032,N_8164);
or U8538 (N_8538,N_8219,N_8113);
nand U8539 (N_8539,N_8212,N_8018);
xor U8540 (N_8540,N_8173,N_8045);
nand U8541 (N_8541,N_8458,N_8282);
or U8542 (N_8542,N_8218,N_8029);
nor U8543 (N_8543,N_8253,N_8103);
nor U8544 (N_8544,N_8043,N_8416);
nand U8545 (N_8545,N_8377,N_8067);
nor U8546 (N_8546,N_8106,N_8476);
and U8547 (N_8547,N_8138,N_8162);
or U8548 (N_8548,N_8161,N_8152);
nor U8549 (N_8549,N_8287,N_8013);
or U8550 (N_8550,N_8050,N_8404);
nor U8551 (N_8551,N_8110,N_8066);
xnor U8552 (N_8552,N_8411,N_8305);
xor U8553 (N_8553,N_8246,N_8078);
nand U8554 (N_8554,N_8383,N_8024);
nand U8555 (N_8555,N_8376,N_8124);
nor U8556 (N_8556,N_8175,N_8023);
nand U8557 (N_8557,N_8107,N_8352);
or U8558 (N_8558,N_8276,N_8046);
and U8559 (N_8559,N_8284,N_8207);
or U8560 (N_8560,N_8460,N_8356);
or U8561 (N_8561,N_8180,N_8432);
xnor U8562 (N_8562,N_8034,N_8498);
xnor U8563 (N_8563,N_8137,N_8388);
nand U8564 (N_8564,N_8170,N_8257);
nor U8565 (N_8565,N_8187,N_8196);
and U8566 (N_8566,N_8453,N_8251);
nor U8567 (N_8567,N_8158,N_8020);
nor U8568 (N_8568,N_8142,N_8330);
xor U8569 (N_8569,N_8166,N_8332);
xnor U8570 (N_8570,N_8168,N_8497);
xnor U8571 (N_8571,N_8122,N_8262);
and U8572 (N_8572,N_8130,N_8457);
nor U8573 (N_8573,N_8454,N_8000);
xnor U8574 (N_8574,N_8490,N_8304);
nand U8575 (N_8575,N_8467,N_8292);
nand U8576 (N_8576,N_8249,N_8444);
xor U8577 (N_8577,N_8421,N_8492);
and U8578 (N_8578,N_8441,N_8489);
xor U8579 (N_8579,N_8038,N_8150);
and U8580 (N_8580,N_8374,N_8496);
xor U8581 (N_8581,N_8157,N_8001);
nand U8582 (N_8582,N_8295,N_8036);
xor U8583 (N_8583,N_8102,N_8208);
and U8584 (N_8584,N_8014,N_8144);
and U8585 (N_8585,N_8204,N_8039);
and U8586 (N_8586,N_8026,N_8155);
or U8587 (N_8587,N_8242,N_8255);
and U8588 (N_8588,N_8384,N_8041);
xnor U8589 (N_8589,N_8483,N_8367);
and U8590 (N_8590,N_8481,N_8231);
nor U8591 (N_8591,N_8378,N_8464);
and U8592 (N_8592,N_8342,N_8402);
nand U8593 (N_8593,N_8436,N_8308);
nand U8594 (N_8594,N_8401,N_8447);
nand U8595 (N_8595,N_8433,N_8149);
and U8596 (N_8596,N_8048,N_8429);
nand U8597 (N_8597,N_8412,N_8133);
nand U8598 (N_8598,N_8471,N_8079);
or U8599 (N_8599,N_8437,N_8357);
and U8600 (N_8600,N_8109,N_8037);
nor U8601 (N_8601,N_8451,N_8071);
xor U8602 (N_8602,N_8475,N_8346);
and U8603 (N_8603,N_8409,N_8366);
nor U8604 (N_8604,N_8336,N_8302);
nand U8605 (N_8605,N_8080,N_8056);
xnor U8606 (N_8606,N_8283,N_8201);
xnor U8607 (N_8607,N_8326,N_8226);
and U8608 (N_8608,N_8105,N_8480);
nor U8609 (N_8609,N_8435,N_8136);
nand U8610 (N_8610,N_8265,N_8317);
and U8611 (N_8611,N_8151,N_8468);
nor U8612 (N_8612,N_8025,N_8008);
or U8613 (N_8613,N_8057,N_8337);
and U8614 (N_8614,N_8355,N_8131);
or U8615 (N_8615,N_8272,N_8229);
xor U8616 (N_8616,N_8306,N_8237);
or U8617 (N_8617,N_8319,N_8063);
and U8618 (N_8618,N_8186,N_8009);
nand U8619 (N_8619,N_8363,N_8260);
xor U8620 (N_8620,N_8120,N_8089);
nand U8621 (N_8621,N_8117,N_8351);
nor U8622 (N_8622,N_8181,N_8121);
nor U8623 (N_8623,N_8123,N_8288);
and U8624 (N_8624,N_8129,N_8300);
nand U8625 (N_8625,N_8169,N_8189);
nand U8626 (N_8626,N_8271,N_8095);
xor U8627 (N_8627,N_8141,N_8299);
xnor U8628 (N_8628,N_8076,N_8312);
or U8629 (N_8629,N_8176,N_8019);
xor U8630 (N_8630,N_8358,N_8097);
xor U8631 (N_8631,N_8178,N_8420);
or U8632 (N_8632,N_8183,N_8390);
xnor U8633 (N_8633,N_8004,N_8266);
nand U8634 (N_8634,N_8128,N_8323);
xor U8635 (N_8635,N_8143,N_8371);
xor U8636 (N_8636,N_8290,N_8375);
nand U8637 (N_8637,N_8167,N_8213);
xnor U8638 (N_8638,N_8233,N_8474);
xnor U8639 (N_8639,N_8338,N_8148);
or U8640 (N_8640,N_8440,N_8301);
or U8641 (N_8641,N_8334,N_8227);
nor U8642 (N_8642,N_8360,N_8058);
nor U8643 (N_8643,N_8238,N_8232);
xor U8644 (N_8644,N_8459,N_8118);
or U8645 (N_8645,N_8425,N_8052);
nor U8646 (N_8646,N_8040,N_8473);
and U8647 (N_8647,N_8177,N_8081);
and U8648 (N_8648,N_8225,N_8006);
nand U8649 (N_8649,N_8406,N_8320);
nor U8650 (N_8650,N_8042,N_8397);
xor U8651 (N_8651,N_8359,N_8488);
nor U8652 (N_8652,N_8339,N_8247);
xnor U8653 (N_8653,N_8462,N_8494);
and U8654 (N_8654,N_8396,N_8373);
and U8655 (N_8655,N_8362,N_8348);
xor U8656 (N_8656,N_8210,N_8493);
nor U8657 (N_8657,N_8147,N_8179);
and U8658 (N_8658,N_8298,N_8470);
nand U8659 (N_8659,N_8463,N_8450);
nor U8660 (N_8660,N_8198,N_8073);
or U8661 (N_8661,N_8114,N_8314);
nor U8662 (N_8662,N_8051,N_8065);
or U8663 (N_8663,N_8111,N_8016);
xor U8664 (N_8664,N_8104,N_8403);
or U8665 (N_8665,N_8259,N_8072);
xor U8666 (N_8666,N_8279,N_8252);
nor U8667 (N_8667,N_8211,N_8487);
or U8668 (N_8668,N_8333,N_8478);
xor U8669 (N_8669,N_8389,N_8372);
nor U8670 (N_8670,N_8070,N_8209);
xor U8671 (N_8671,N_8485,N_8382);
nor U8672 (N_8672,N_8393,N_8439);
or U8673 (N_8673,N_8340,N_8264);
nand U8674 (N_8674,N_8294,N_8171);
and U8675 (N_8675,N_8250,N_8413);
and U8676 (N_8676,N_8127,N_8191);
or U8677 (N_8677,N_8491,N_8075);
nand U8678 (N_8678,N_8244,N_8116);
nor U8679 (N_8679,N_8407,N_8415);
nor U8680 (N_8680,N_8408,N_8379);
nor U8681 (N_8681,N_8313,N_8059);
nand U8682 (N_8682,N_8003,N_8230);
nor U8683 (N_8683,N_8466,N_8414);
or U8684 (N_8684,N_8172,N_8443);
xor U8685 (N_8685,N_8327,N_8200);
xnor U8686 (N_8686,N_8349,N_8495);
and U8687 (N_8687,N_8055,N_8442);
nand U8688 (N_8688,N_8044,N_8427);
or U8689 (N_8689,N_8278,N_8418);
or U8690 (N_8690,N_8027,N_8188);
xnor U8691 (N_8691,N_8064,N_8145);
or U8692 (N_8692,N_8153,N_8203);
xor U8693 (N_8693,N_8263,N_8185);
xnor U8694 (N_8694,N_8215,N_8434);
nor U8695 (N_8695,N_8364,N_8206);
or U8696 (N_8696,N_8438,N_8445);
or U8697 (N_8697,N_8315,N_8077);
nor U8698 (N_8698,N_8248,N_8085);
nor U8699 (N_8699,N_8021,N_8074);
or U8700 (N_8700,N_8062,N_8217);
nand U8701 (N_8701,N_8446,N_8277);
nor U8702 (N_8702,N_8261,N_8069);
and U8703 (N_8703,N_8499,N_8090);
xor U8704 (N_8704,N_8400,N_8318);
nor U8705 (N_8705,N_8205,N_8195);
or U8706 (N_8706,N_8174,N_8424);
xor U8707 (N_8707,N_8119,N_8154);
nand U8708 (N_8708,N_8386,N_8391);
xnor U8709 (N_8709,N_8344,N_8083);
or U8710 (N_8710,N_8354,N_8303);
xnor U8711 (N_8711,N_8285,N_8431);
nor U8712 (N_8712,N_8449,N_8274);
xor U8713 (N_8713,N_8254,N_8461);
xnor U8714 (N_8714,N_8159,N_8482);
or U8715 (N_8715,N_8101,N_8452);
or U8716 (N_8716,N_8108,N_8224);
nor U8717 (N_8717,N_8335,N_8297);
and U8718 (N_8718,N_8005,N_8465);
and U8719 (N_8719,N_8163,N_8156);
or U8720 (N_8720,N_8291,N_8448);
nand U8721 (N_8721,N_8002,N_8365);
xor U8722 (N_8722,N_8410,N_8347);
or U8723 (N_8723,N_8235,N_8469);
xnor U8724 (N_8724,N_8329,N_8385);
and U8725 (N_8725,N_8222,N_8125);
xor U8726 (N_8726,N_8010,N_8022);
or U8727 (N_8727,N_8328,N_8455);
and U8728 (N_8728,N_8139,N_8310);
or U8729 (N_8729,N_8422,N_8479);
xor U8730 (N_8730,N_8192,N_8343);
or U8731 (N_8731,N_8258,N_8392);
and U8732 (N_8732,N_8194,N_8369);
xnor U8733 (N_8733,N_8381,N_8132);
nor U8734 (N_8734,N_8061,N_8293);
xnor U8735 (N_8735,N_8220,N_8296);
nand U8736 (N_8736,N_8398,N_8430);
nor U8737 (N_8737,N_8140,N_8280);
nor U8738 (N_8738,N_8423,N_8361);
and U8739 (N_8739,N_8405,N_8486);
nand U8740 (N_8740,N_8353,N_8370);
or U8741 (N_8741,N_8197,N_8049);
nand U8742 (N_8742,N_8007,N_8350);
nand U8743 (N_8743,N_8236,N_8092);
and U8744 (N_8744,N_8240,N_8289);
xnor U8745 (N_8745,N_8093,N_8275);
nor U8746 (N_8746,N_8182,N_8387);
nand U8747 (N_8747,N_8135,N_8134);
nor U8748 (N_8748,N_8321,N_8028);
nand U8749 (N_8749,N_8099,N_8096);
nand U8750 (N_8750,N_8001,N_8015);
or U8751 (N_8751,N_8299,N_8249);
or U8752 (N_8752,N_8264,N_8434);
nor U8753 (N_8753,N_8454,N_8313);
nor U8754 (N_8754,N_8305,N_8309);
xor U8755 (N_8755,N_8028,N_8270);
xnor U8756 (N_8756,N_8485,N_8132);
nand U8757 (N_8757,N_8297,N_8129);
xnor U8758 (N_8758,N_8410,N_8291);
or U8759 (N_8759,N_8466,N_8214);
xnor U8760 (N_8760,N_8440,N_8432);
or U8761 (N_8761,N_8247,N_8088);
nor U8762 (N_8762,N_8069,N_8239);
and U8763 (N_8763,N_8384,N_8010);
nand U8764 (N_8764,N_8076,N_8416);
nor U8765 (N_8765,N_8375,N_8347);
nand U8766 (N_8766,N_8411,N_8239);
nor U8767 (N_8767,N_8482,N_8304);
and U8768 (N_8768,N_8119,N_8359);
xor U8769 (N_8769,N_8065,N_8373);
xnor U8770 (N_8770,N_8022,N_8167);
or U8771 (N_8771,N_8089,N_8091);
nor U8772 (N_8772,N_8463,N_8448);
or U8773 (N_8773,N_8112,N_8197);
and U8774 (N_8774,N_8068,N_8183);
or U8775 (N_8775,N_8091,N_8028);
and U8776 (N_8776,N_8351,N_8165);
xnor U8777 (N_8777,N_8065,N_8338);
or U8778 (N_8778,N_8265,N_8490);
nor U8779 (N_8779,N_8291,N_8425);
nor U8780 (N_8780,N_8230,N_8064);
nand U8781 (N_8781,N_8094,N_8269);
nor U8782 (N_8782,N_8106,N_8137);
and U8783 (N_8783,N_8455,N_8409);
or U8784 (N_8784,N_8070,N_8179);
and U8785 (N_8785,N_8043,N_8127);
and U8786 (N_8786,N_8387,N_8496);
and U8787 (N_8787,N_8332,N_8130);
nand U8788 (N_8788,N_8318,N_8055);
xor U8789 (N_8789,N_8238,N_8033);
nor U8790 (N_8790,N_8357,N_8351);
xor U8791 (N_8791,N_8127,N_8091);
xnor U8792 (N_8792,N_8469,N_8141);
or U8793 (N_8793,N_8219,N_8205);
and U8794 (N_8794,N_8387,N_8287);
nor U8795 (N_8795,N_8318,N_8404);
nand U8796 (N_8796,N_8373,N_8233);
or U8797 (N_8797,N_8493,N_8166);
nand U8798 (N_8798,N_8477,N_8398);
xor U8799 (N_8799,N_8480,N_8459);
and U8800 (N_8800,N_8150,N_8354);
xor U8801 (N_8801,N_8474,N_8338);
xnor U8802 (N_8802,N_8340,N_8206);
nor U8803 (N_8803,N_8013,N_8155);
or U8804 (N_8804,N_8180,N_8210);
or U8805 (N_8805,N_8487,N_8156);
nor U8806 (N_8806,N_8456,N_8293);
or U8807 (N_8807,N_8398,N_8338);
nor U8808 (N_8808,N_8144,N_8337);
nor U8809 (N_8809,N_8011,N_8023);
or U8810 (N_8810,N_8108,N_8475);
and U8811 (N_8811,N_8356,N_8132);
or U8812 (N_8812,N_8493,N_8015);
xor U8813 (N_8813,N_8063,N_8458);
xor U8814 (N_8814,N_8348,N_8292);
and U8815 (N_8815,N_8444,N_8406);
nand U8816 (N_8816,N_8055,N_8021);
nor U8817 (N_8817,N_8281,N_8156);
xor U8818 (N_8818,N_8488,N_8016);
and U8819 (N_8819,N_8204,N_8208);
nor U8820 (N_8820,N_8442,N_8329);
or U8821 (N_8821,N_8051,N_8056);
nor U8822 (N_8822,N_8047,N_8007);
or U8823 (N_8823,N_8192,N_8141);
xor U8824 (N_8824,N_8059,N_8492);
nor U8825 (N_8825,N_8265,N_8469);
nor U8826 (N_8826,N_8403,N_8173);
nand U8827 (N_8827,N_8361,N_8222);
nand U8828 (N_8828,N_8063,N_8233);
nor U8829 (N_8829,N_8098,N_8148);
nand U8830 (N_8830,N_8412,N_8216);
nor U8831 (N_8831,N_8077,N_8147);
nor U8832 (N_8832,N_8327,N_8170);
or U8833 (N_8833,N_8041,N_8032);
xor U8834 (N_8834,N_8199,N_8152);
and U8835 (N_8835,N_8430,N_8371);
nor U8836 (N_8836,N_8443,N_8466);
or U8837 (N_8837,N_8176,N_8491);
and U8838 (N_8838,N_8055,N_8079);
xor U8839 (N_8839,N_8425,N_8209);
nand U8840 (N_8840,N_8451,N_8282);
nor U8841 (N_8841,N_8195,N_8091);
nand U8842 (N_8842,N_8286,N_8288);
xor U8843 (N_8843,N_8457,N_8083);
or U8844 (N_8844,N_8160,N_8382);
nor U8845 (N_8845,N_8295,N_8222);
nand U8846 (N_8846,N_8079,N_8263);
xor U8847 (N_8847,N_8426,N_8301);
nor U8848 (N_8848,N_8031,N_8045);
nand U8849 (N_8849,N_8084,N_8347);
nand U8850 (N_8850,N_8282,N_8013);
or U8851 (N_8851,N_8448,N_8318);
and U8852 (N_8852,N_8180,N_8292);
and U8853 (N_8853,N_8148,N_8250);
nor U8854 (N_8854,N_8185,N_8150);
and U8855 (N_8855,N_8235,N_8060);
nand U8856 (N_8856,N_8025,N_8466);
xor U8857 (N_8857,N_8230,N_8418);
nor U8858 (N_8858,N_8174,N_8010);
or U8859 (N_8859,N_8444,N_8455);
and U8860 (N_8860,N_8489,N_8198);
nor U8861 (N_8861,N_8198,N_8211);
and U8862 (N_8862,N_8387,N_8153);
nand U8863 (N_8863,N_8307,N_8234);
or U8864 (N_8864,N_8191,N_8481);
nor U8865 (N_8865,N_8265,N_8436);
xor U8866 (N_8866,N_8468,N_8273);
nor U8867 (N_8867,N_8103,N_8424);
and U8868 (N_8868,N_8425,N_8100);
and U8869 (N_8869,N_8179,N_8286);
and U8870 (N_8870,N_8328,N_8187);
and U8871 (N_8871,N_8120,N_8174);
xnor U8872 (N_8872,N_8175,N_8101);
or U8873 (N_8873,N_8179,N_8441);
and U8874 (N_8874,N_8489,N_8288);
xor U8875 (N_8875,N_8294,N_8276);
nor U8876 (N_8876,N_8419,N_8493);
nor U8877 (N_8877,N_8025,N_8215);
xor U8878 (N_8878,N_8346,N_8343);
and U8879 (N_8879,N_8067,N_8223);
nand U8880 (N_8880,N_8233,N_8002);
xnor U8881 (N_8881,N_8141,N_8241);
nand U8882 (N_8882,N_8227,N_8299);
nor U8883 (N_8883,N_8119,N_8192);
nor U8884 (N_8884,N_8395,N_8191);
or U8885 (N_8885,N_8224,N_8384);
nor U8886 (N_8886,N_8410,N_8188);
and U8887 (N_8887,N_8275,N_8432);
nor U8888 (N_8888,N_8426,N_8094);
xor U8889 (N_8889,N_8415,N_8361);
or U8890 (N_8890,N_8240,N_8157);
xnor U8891 (N_8891,N_8170,N_8306);
or U8892 (N_8892,N_8021,N_8273);
nor U8893 (N_8893,N_8278,N_8338);
and U8894 (N_8894,N_8140,N_8485);
and U8895 (N_8895,N_8357,N_8391);
or U8896 (N_8896,N_8233,N_8105);
or U8897 (N_8897,N_8436,N_8300);
and U8898 (N_8898,N_8282,N_8425);
and U8899 (N_8899,N_8310,N_8404);
or U8900 (N_8900,N_8144,N_8331);
xor U8901 (N_8901,N_8247,N_8142);
and U8902 (N_8902,N_8059,N_8465);
nor U8903 (N_8903,N_8385,N_8193);
nor U8904 (N_8904,N_8171,N_8149);
nor U8905 (N_8905,N_8096,N_8163);
nor U8906 (N_8906,N_8438,N_8393);
nor U8907 (N_8907,N_8076,N_8332);
or U8908 (N_8908,N_8327,N_8078);
or U8909 (N_8909,N_8236,N_8295);
nor U8910 (N_8910,N_8112,N_8497);
and U8911 (N_8911,N_8126,N_8182);
or U8912 (N_8912,N_8440,N_8337);
nand U8913 (N_8913,N_8323,N_8173);
and U8914 (N_8914,N_8109,N_8452);
or U8915 (N_8915,N_8103,N_8286);
or U8916 (N_8916,N_8169,N_8079);
nand U8917 (N_8917,N_8454,N_8453);
nor U8918 (N_8918,N_8027,N_8229);
nand U8919 (N_8919,N_8231,N_8109);
and U8920 (N_8920,N_8365,N_8378);
or U8921 (N_8921,N_8005,N_8391);
xor U8922 (N_8922,N_8330,N_8094);
xnor U8923 (N_8923,N_8455,N_8104);
xor U8924 (N_8924,N_8402,N_8243);
nor U8925 (N_8925,N_8289,N_8439);
nand U8926 (N_8926,N_8228,N_8460);
and U8927 (N_8927,N_8020,N_8197);
nand U8928 (N_8928,N_8482,N_8487);
and U8929 (N_8929,N_8473,N_8233);
nor U8930 (N_8930,N_8241,N_8194);
xor U8931 (N_8931,N_8074,N_8298);
xor U8932 (N_8932,N_8125,N_8005);
xnor U8933 (N_8933,N_8340,N_8077);
and U8934 (N_8934,N_8096,N_8354);
and U8935 (N_8935,N_8036,N_8395);
nor U8936 (N_8936,N_8497,N_8334);
nand U8937 (N_8937,N_8370,N_8252);
nand U8938 (N_8938,N_8392,N_8216);
nand U8939 (N_8939,N_8306,N_8224);
or U8940 (N_8940,N_8097,N_8418);
nand U8941 (N_8941,N_8427,N_8397);
or U8942 (N_8942,N_8164,N_8428);
xnor U8943 (N_8943,N_8389,N_8351);
nor U8944 (N_8944,N_8354,N_8235);
nand U8945 (N_8945,N_8191,N_8309);
xnor U8946 (N_8946,N_8145,N_8202);
nand U8947 (N_8947,N_8401,N_8201);
nor U8948 (N_8948,N_8148,N_8245);
and U8949 (N_8949,N_8272,N_8186);
and U8950 (N_8950,N_8011,N_8253);
or U8951 (N_8951,N_8112,N_8194);
xnor U8952 (N_8952,N_8396,N_8310);
and U8953 (N_8953,N_8032,N_8251);
or U8954 (N_8954,N_8158,N_8423);
xnor U8955 (N_8955,N_8446,N_8314);
nand U8956 (N_8956,N_8040,N_8192);
xor U8957 (N_8957,N_8410,N_8127);
nand U8958 (N_8958,N_8119,N_8391);
nor U8959 (N_8959,N_8403,N_8359);
nor U8960 (N_8960,N_8330,N_8229);
nand U8961 (N_8961,N_8065,N_8339);
xor U8962 (N_8962,N_8350,N_8024);
or U8963 (N_8963,N_8275,N_8331);
nor U8964 (N_8964,N_8000,N_8165);
and U8965 (N_8965,N_8171,N_8218);
or U8966 (N_8966,N_8008,N_8235);
xor U8967 (N_8967,N_8276,N_8466);
nor U8968 (N_8968,N_8328,N_8296);
and U8969 (N_8969,N_8065,N_8096);
or U8970 (N_8970,N_8149,N_8292);
nand U8971 (N_8971,N_8167,N_8311);
nor U8972 (N_8972,N_8315,N_8374);
nand U8973 (N_8973,N_8289,N_8328);
nand U8974 (N_8974,N_8205,N_8163);
xnor U8975 (N_8975,N_8340,N_8186);
and U8976 (N_8976,N_8380,N_8072);
or U8977 (N_8977,N_8000,N_8172);
and U8978 (N_8978,N_8191,N_8067);
and U8979 (N_8979,N_8413,N_8339);
or U8980 (N_8980,N_8118,N_8181);
and U8981 (N_8981,N_8267,N_8359);
and U8982 (N_8982,N_8255,N_8405);
and U8983 (N_8983,N_8172,N_8310);
and U8984 (N_8984,N_8168,N_8121);
or U8985 (N_8985,N_8027,N_8367);
nand U8986 (N_8986,N_8290,N_8342);
nor U8987 (N_8987,N_8478,N_8033);
or U8988 (N_8988,N_8447,N_8230);
nor U8989 (N_8989,N_8291,N_8355);
and U8990 (N_8990,N_8147,N_8013);
nor U8991 (N_8991,N_8206,N_8199);
nand U8992 (N_8992,N_8025,N_8242);
nor U8993 (N_8993,N_8034,N_8200);
or U8994 (N_8994,N_8392,N_8205);
xnor U8995 (N_8995,N_8413,N_8208);
or U8996 (N_8996,N_8187,N_8366);
nand U8997 (N_8997,N_8039,N_8495);
and U8998 (N_8998,N_8098,N_8051);
nand U8999 (N_8999,N_8254,N_8477);
nand U9000 (N_9000,N_8803,N_8509);
xnor U9001 (N_9001,N_8665,N_8772);
xor U9002 (N_9002,N_8735,N_8513);
and U9003 (N_9003,N_8629,N_8973);
xnor U9004 (N_9004,N_8943,N_8972);
and U9005 (N_9005,N_8981,N_8628);
nand U9006 (N_9006,N_8500,N_8843);
nand U9007 (N_9007,N_8714,N_8773);
and U9008 (N_9008,N_8534,N_8904);
and U9009 (N_9009,N_8747,N_8991);
and U9010 (N_9010,N_8692,N_8979);
or U9011 (N_9011,N_8758,N_8977);
or U9012 (N_9012,N_8903,N_8530);
nand U9013 (N_9013,N_8937,N_8944);
and U9014 (N_9014,N_8797,N_8784);
nand U9015 (N_9015,N_8835,N_8709);
nand U9016 (N_9016,N_8865,N_8566);
xor U9017 (N_9017,N_8621,N_8616);
and U9018 (N_9018,N_8706,N_8587);
nand U9019 (N_9019,N_8820,N_8744);
xnor U9020 (N_9020,N_8674,N_8508);
and U9021 (N_9021,N_8823,N_8532);
nand U9022 (N_9022,N_8524,N_8716);
nor U9023 (N_9023,N_8883,N_8642);
or U9024 (N_9024,N_8808,N_8875);
xnor U9025 (N_9025,N_8559,N_8946);
nand U9026 (N_9026,N_8762,N_8544);
nor U9027 (N_9027,N_8565,N_8682);
xnor U9028 (N_9028,N_8792,N_8833);
xor U9029 (N_9029,N_8676,N_8531);
or U9030 (N_9030,N_8574,N_8677);
nand U9031 (N_9031,N_8660,N_8867);
xnor U9032 (N_9032,N_8745,N_8655);
xnor U9033 (N_9033,N_8759,N_8834);
and U9034 (N_9034,N_8811,N_8764);
and U9035 (N_9035,N_8970,N_8506);
and U9036 (N_9036,N_8750,N_8926);
and U9037 (N_9037,N_8888,N_8868);
xor U9038 (N_9038,N_8966,N_8552);
nor U9039 (N_9039,N_8778,N_8561);
and U9040 (N_9040,N_8684,N_8731);
or U9041 (N_9041,N_8732,N_8514);
xor U9042 (N_9042,N_8942,N_8869);
xor U9043 (N_9043,N_8839,N_8899);
nor U9044 (N_9044,N_8641,N_8549);
or U9045 (N_9045,N_8995,N_8688);
and U9046 (N_9046,N_8595,N_8892);
xnor U9047 (N_9047,N_8578,N_8623);
and U9048 (N_9048,N_8860,N_8902);
nand U9049 (N_9049,N_8504,N_8854);
nand U9050 (N_9050,N_8601,N_8829);
nor U9051 (N_9051,N_8915,N_8941);
nand U9052 (N_9052,N_8733,N_8765);
nor U9053 (N_9053,N_8841,N_8555);
nand U9054 (N_9054,N_8852,N_8567);
nor U9055 (N_9055,N_8525,N_8985);
and U9056 (N_9056,N_8689,N_8771);
and U9057 (N_9057,N_8901,N_8591);
nand U9058 (N_9058,N_8556,N_8592);
nor U9059 (N_9059,N_8712,N_8931);
and U9060 (N_9060,N_8611,N_8846);
or U9061 (N_9061,N_8840,N_8720);
and U9062 (N_9062,N_8551,N_8900);
nor U9063 (N_9063,N_8763,N_8550);
or U9064 (N_9064,N_8626,N_8945);
and U9065 (N_9065,N_8810,N_8956);
nand U9066 (N_9066,N_8769,N_8668);
nand U9067 (N_9067,N_8729,N_8636);
or U9068 (N_9068,N_8802,N_8622);
xor U9069 (N_9069,N_8739,N_8817);
and U9070 (N_9070,N_8805,N_8992);
xnor U9071 (N_9071,N_8889,N_8520);
and U9072 (N_9072,N_8515,N_8648);
nand U9073 (N_9073,N_8516,N_8569);
or U9074 (N_9074,N_8738,N_8603);
xor U9075 (N_9075,N_8962,N_8940);
xor U9076 (N_9076,N_8662,N_8861);
or U9077 (N_9077,N_8503,N_8678);
or U9078 (N_9078,N_8768,N_8886);
xnor U9079 (N_9079,N_8533,N_8830);
or U9080 (N_9080,N_8547,N_8734);
nand U9081 (N_9081,N_8652,N_8948);
nor U9082 (N_9082,N_8670,N_8816);
xnor U9083 (N_9083,N_8708,N_8653);
xnor U9084 (N_9084,N_8838,N_8698);
xor U9085 (N_9085,N_8675,N_8701);
xnor U9086 (N_9086,N_8850,N_8697);
or U9087 (N_9087,N_8934,N_8596);
xor U9088 (N_9088,N_8749,N_8971);
or U9089 (N_9089,N_8990,N_8667);
xor U9090 (N_9090,N_8983,N_8987);
nand U9091 (N_9091,N_8913,N_8960);
nor U9092 (N_9092,N_8519,N_8522);
nand U9093 (N_9093,N_8613,N_8502);
nand U9094 (N_9094,N_8725,N_8752);
nand U9095 (N_9095,N_8743,N_8878);
and U9096 (N_9096,N_8679,N_8954);
and U9097 (N_9097,N_8620,N_8666);
xnor U9098 (N_9098,N_8891,N_8862);
nand U9099 (N_9099,N_8627,N_8920);
and U9100 (N_9100,N_8543,N_8760);
nor U9101 (N_9101,N_8558,N_8952);
and U9102 (N_9102,N_8681,N_8707);
or U9103 (N_9103,N_8832,N_8510);
and U9104 (N_9104,N_8614,N_8896);
nand U9105 (N_9105,N_8780,N_8571);
and U9106 (N_9106,N_8807,N_8964);
nand U9107 (N_9107,N_8786,N_8562);
nor U9108 (N_9108,N_8767,N_8997);
nand U9109 (N_9109,N_8602,N_8849);
or U9110 (N_9110,N_8965,N_8967);
nand U9111 (N_9111,N_8593,N_8798);
xor U9112 (N_9112,N_8507,N_8882);
and U9113 (N_9113,N_8959,N_8597);
xor U9114 (N_9114,N_8686,N_8505);
or U9115 (N_9115,N_8586,N_8542);
nand U9116 (N_9116,N_8728,N_8950);
or U9117 (N_9117,N_8610,N_8528);
nor U9118 (N_9118,N_8872,N_8982);
or U9119 (N_9119,N_8564,N_8608);
nand U9120 (N_9120,N_8837,N_8615);
xor U9121 (N_9121,N_8723,N_8844);
or U9122 (N_9122,N_8700,N_8585);
nor U9123 (N_9123,N_8907,N_8927);
nor U9124 (N_9124,N_8770,N_8800);
xnor U9125 (N_9125,N_8821,N_8935);
and U9126 (N_9126,N_8909,N_8737);
nor U9127 (N_9127,N_8687,N_8703);
and U9128 (N_9128,N_8649,N_8819);
nand U9129 (N_9129,N_8887,N_8672);
nand U9130 (N_9130,N_8921,N_8788);
or U9131 (N_9131,N_8781,N_8584);
and U9132 (N_9132,N_8986,N_8580);
nor U9133 (N_9133,N_8570,N_8624);
xor U9134 (N_9134,N_8957,N_8836);
nor U9135 (N_9135,N_8646,N_8925);
xnor U9136 (N_9136,N_8951,N_8933);
xnor U9137 (N_9137,N_8748,N_8695);
xnor U9138 (N_9138,N_8908,N_8806);
nor U9139 (N_9139,N_8905,N_8809);
xor U9140 (N_9140,N_8710,N_8645);
nand U9141 (N_9141,N_8822,N_8815);
nand U9142 (N_9142,N_8791,N_8922);
nand U9143 (N_9143,N_8606,N_8897);
and U9144 (N_9144,N_8799,N_8717);
xor U9145 (N_9145,N_8523,N_8975);
and U9146 (N_9146,N_8742,N_8993);
nand U9147 (N_9147,N_8976,N_8978);
and U9148 (N_9148,N_8501,N_8855);
and U9149 (N_9149,N_8775,N_8919);
xnor U9150 (N_9150,N_8537,N_8604);
nor U9151 (N_9151,N_8661,N_8605);
xor U9152 (N_9152,N_8656,N_8658);
or U9153 (N_9153,N_8754,N_8782);
and U9154 (N_9154,N_8715,N_8912);
nand U9155 (N_9155,N_8635,N_8884);
and U9156 (N_9156,N_8851,N_8609);
and U9157 (N_9157,N_8877,N_8654);
xnor U9158 (N_9158,N_8890,N_8568);
or U9159 (N_9159,N_8774,N_8518);
and U9160 (N_9160,N_8651,N_8546);
or U9161 (N_9161,N_8989,N_8916);
nand U9162 (N_9162,N_8521,N_8705);
nand U9163 (N_9163,N_8751,N_8690);
and U9164 (N_9164,N_8563,N_8895);
xor U9165 (N_9165,N_8804,N_8826);
nor U9166 (N_9166,N_8711,N_8893);
nor U9167 (N_9167,N_8718,N_8577);
nand U9168 (N_9168,N_8526,N_8726);
or U9169 (N_9169,N_8793,N_8557);
nor U9170 (N_9170,N_8879,N_8873);
and U9171 (N_9171,N_8924,N_8573);
and U9172 (N_9172,N_8801,N_8633);
and U9173 (N_9173,N_8637,N_8980);
nor U9174 (N_9174,N_8831,N_8818);
nor U9175 (N_9175,N_8517,N_8864);
nand U9176 (N_9176,N_8812,N_8650);
and U9177 (N_9177,N_8612,N_8572);
nor U9178 (N_9178,N_8724,N_8827);
or U9179 (N_9179,N_8657,N_8755);
xnor U9180 (N_9180,N_8968,N_8664);
or U9181 (N_9181,N_8858,N_8647);
or U9182 (N_9182,N_8906,N_8848);
and U9183 (N_9183,N_8947,N_8625);
or U9184 (N_9184,N_8842,N_8880);
or U9185 (N_9185,N_8813,N_8691);
and U9186 (N_9186,N_8560,N_8581);
nor U9187 (N_9187,N_8790,N_8814);
nand U9188 (N_9188,N_8783,N_8730);
and U9189 (N_9189,N_8529,N_8669);
nor U9190 (N_9190,N_8631,N_8949);
and U9191 (N_9191,N_8512,N_8548);
xnor U9192 (N_9192,N_8961,N_8936);
and U9193 (N_9193,N_8999,N_8847);
and U9194 (N_9194,N_8885,N_8576);
xnor U9195 (N_9195,N_8988,N_8589);
and U9196 (N_9196,N_8994,N_8824);
xnor U9197 (N_9197,N_8955,N_8579);
and U9198 (N_9198,N_8618,N_8598);
or U9199 (N_9199,N_8756,N_8953);
nand U9200 (N_9200,N_8871,N_8859);
nor U9201 (N_9201,N_8535,N_8683);
or U9202 (N_9202,N_8619,N_8794);
nand U9203 (N_9203,N_8785,N_8766);
nand U9204 (N_9204,N_8538,N_8600);
xor U9205 (N_9205,N_8828,N_8643);
and U9206 (N_9206,N_8874,N_8939);
xor U9207 (N_9207,N_8876,N_8640);
or U9208 (N_9208,N_8638,N_8998);
or U9209 (N_9209,N_8554,N_8594);
and U9210 (N_9210,N_8588,N_8736);
and U9211 (N_9211,N_8540,N_8599);
xor U9212 (N_9212,N_8796,N_8541);
nand U9213 (N_9213,N_8795,N_8918);
or U9214 (N_9214,N_8787,N_8673);
xor U9215 (N_9215,N_8753,N_8761);
nor U9216 (N_9216,N_8853,N_8963);
nand U9217 (N_9217,N_8984,N_8974);
nor U9218 (N_9218,N_8938,N_8727);
nand U9219 (N_9219,N_8856,N_8923);
or U9220 (N_9220,N_8969,N_8644);
xnor U9221 (N_9221,N_8632,N_8536);
nor U9222 (N_9222,N_8545,N_8671);
nor U9223 (N_9223,N_8696,N_8575);
and U9224 (N_9224,N_8870,N_8917);
or U9225 (N_9225,N_8607,N_8929);
nor U9226 (N_9226,N_8617,N_8699);
nand U9227 (N_9227,N_8722,N_8958);
xor U9228 (N_9228,N_8898,N_8634);
nand U9229 (N_9229,N_8866,N_8863);
xnor U9230 (N_9230,N_8590,N_8910);
nand U9231 (N_9231,N_8857,N_8639);
nand U9232 (N_9232,N_8511,N_8741);
nand U9233 (N_9233,N_8713,N_8583);
nand U9234 (N_9234,N_8845,N_8996);
nor U9235 (N_9235,N_8685,N_8928);
nor U9236 (N_9236,N_8932,N_8881);
xnor U9237 (N_9237,N_8659,N_8582);
nor U9238 (N_9238,N_8779,N_8825);
and U9239 (N_9239,N_8630,N_8777);
or U9240 (N_9240,N_8776,N_8663);
and U9241 (N_9241,N_8740,N_8914);
and U9242 (N_9242,N_8894,N_8702);
or U9243 (N_9243,N_8911,N_8693);
or U9244 (N_9244,N_8704,N_8719);
xor U9245 (N_9245,N_8789,N_8553);
nor U9246 (N_9246,N_8930,N_8694);
nor U9247 (N_9247,N_8527,N_8746);
nand U9248 (N_9248,N_8680,N_8721);
and U9249 (N_9249,N_8757,N_8539);
xnor U9250 (N_9250,N_8760,N_8629);
or U9251 (N_9251,N_8502,N_8700);
xor U9252 (N_9252,N_8681,N_8806);
xor U9253 (N_9253,N_8548,N_8592);
nand U9254 (N_9254,N_8958,N_8696);
nand U9255 (N_9255,N_8735,N_8779);
xor U9256 (N_9256,N_8892,N_8620);
nor U9257 (N_9257,N_8897,N_8680);
nand U9258 (N_9258,N_8992,N_8630);
nand U9259 (N_9259,N_8618,N_8694);
and U9260 (N_9260,N_8574,N_8869);
and U9261 (N_9261,N_8803,N_8618);
nor U9262 (N_9262,N_8549,N_8610);
or U9263 (N_9263,N_8995,N_8591);
xor U9264 (N_9264,N_8978,N_8723);
and U9265 (N_9265,N_8743,N_8581);
nor U9266 (N_9266,N_8994,N_8546);
xnor U9267 (N_9267,N_8796,N_8860);
or U9268 (N_9268,N_8823,N_8659);
or U9269 (N_9269,N_8504,N_8892);
xor U9270 (N_9270,N_8833,N_8550);
and U9271 (N_9271,N_8935,N_8720);
xnor U9272 (N_9272,N_8676,N_8602);
nor U9273 (N_9273,N_8962,N_8765);
nor U9274 (N_9274,N_8911,N_8898);
xor U9275 (N_9275,N_8758,N_8940);
nand U9276 (N_9276,N_8934,N_8731);
nand U9277 (N_9277,N_8958,N_8948);
nor U9278 (N_9278,N_8918,N_8595);
or U9279 (N_9279,N_8634,N_8984);
or U9280 (N_9280,N_8752,N_8600);
and U9281 (N_9281,N_8650,N_8871);
or U9282 (N_9282,N_8535,N_8601);
and U9283 (N_9283,N_8718,N_8983);
nand U9284 (N_9284,N_8871,N_8680);
xor U9285 (N_9285,N_8815,N_8764);
nor U9286 (N_9286,N_8696,N_8780);
nand U9287 (N_9287,N_8828,N_8653);
and U9288 (N_9288,N_8948,N_8639);
nor U9289 (N_9289,N_8725,N_8959);
or U9290 (N_9290,N_8546,N_8841);
nand U9291 (N_9291,N_8705,N_8728);
nand U9292 (N_9292,N_8698,N_8738);
or U9293 (N_9293,N_8509,N_8513);
xor U9294 (N_9294,N_8557,N_8887);
and U9295 (N_9295,N_8971,N_8928);
and U9296 (N_9296,N_8853,N_8715);
xor U9297 (N_9297,N_8558,N_8803);
nand U9298 (N_9298,N_8506,N_8956);
nand U9299 (N_9299,N_8965,N_8891);
xnor U9300 (N_9300,N_8882,N_8609);
nor U9301 (N_9301,N_8999,N_8635);
or U9302 (N_9302,N_8586,N_8742);
xor U9303 (N_9303,N_8694,N_8610);
and U9304 (N_9304,N_8759,N_8821);
or U9305 (N_9305,N_8598,N_8890);
nand U9306 (N_9306,N_8990,N_8526);
and U9307 (N_9307,N_8733,N_8648);
nor U9308 (N_9308,N_8702,N_8606);
xor U9309 (N_9309,N_8689,N_8869);
nand U9310 (N_9310,N_8841,N_8889);
nand U9311 (N_9311,N_8980,N_8879);
or U9312 (N_9312,N_8526,N_8842);
and U9313 (N_9313,N_8651,N_8966);
nand U9314 (N_9314,N_8890,N_8608);
and U9315 (N_9315,N_8570,N_8597);
nor U9316 (N_9316,N_8503,N_8772);
or U9317 (N_9317,N_8671,N_8995);
and U9318 (N_9318,N_8750,N_8563);
nor U9319 (N_9319,N_8787,N_8829);
and U9320 (N_9320,N_8504,N_8975);
nor U9321 (N_9321,N_8923,N_8962);
nand U9322 (N_9322,N_8566,N_8810);
or U9323 (N_9323,N_8598,N_8933);
or U9324 (N_9324,N_8550,N_8777);
xor U9325 (N_9325,N_8713,N_8678);
nand U9326 (N_9326,N_8988,N_8719);
nor U9327 (N_9327,N_8975,N_8553);
or U9328 (N_9328,N_8587,N_8593);
nor U9329 (N_9329,N_8919,N_8717);
xor U9330 (N_9330,N_8682,N_8832);
or U9331 (N_9331,N_8819,N_8526);
nor U9332 (N_9332,N_8672,N_8860);
nor U9333 (N_9333,N_8848,N_8522);
xor U9334 (N_9334,N_8842,N_8556);
nand U9335 (N_9335,N_8745,N_8995);
or U9336 (N_9336,N_8613,N_8940);
xor U9337 (N_9337,N_8975,N_8725);
nand U9338 (N_9338,N_8658,N_8529);
nand U9339 (N_9339,N_8760,N_8998);
or U9340 (N_9340,N_8752,N_8874);
or U9341 (N_9341,N_8741,N_8795);
nand U9342 (N_9342,N_8941,N_8835);
and U9343 (N_9343,N_8544,N_8872);
or U9344 (N_9344,N_8690,N_8682);
nor U9345 (N_9345,N_8774,N_8993);
nor U9346 (N_9346,N_8735,N_8623);
and U9347 (N_9347,N_8600,N_8552);
nand U9348 (N_9348,N_8894,N_8989);
nand U9349 (N_9349,N_8579,N_8587);
xnor U9350 (N_9350,N_8962,N_8679);
or U9351 (N_9351,N_8907,N_8500);
and U9352 (N_9352,N_8661,N_8517);
nor U9353 (N_9353,N_8951,N_8628);
or U9354 (N_9354,N_8815,N_8787);
nand U9355 (N_9355,N_8931,N_8895);
and U9356 (N_9356,N_8629,N_8614);
nand U9357 (N_9357,N_8607,N_8518);
nor U9358 (N_9358,N_8908,N_8854);
or U9359 (N_9359,N_8619,N_8556);
and U9360 (N_9360,N_8894,N_8959);
nand U9361 (N_9361,N_8843,N_8588);
or U9362 (N_9362,N_8643,N_8789);
nand U9363 (N_9363,N_8508,N_8769);
nand U9364 (N_9364,N_8934,N_8534);
or U9365 (N_9365,N_8701,N_8762);
or U9366 (N_9366,N_8546,N_8783);
or U9367 (N_9367,N_8726,N_8594);
xor U9368 (N_9368,N_8623,N_8901);
nand U9369 (N_9369,N_8861,N_8774);
or U9370 (N_9370,N_8514,N_8813);
nor U9371 (N_9371,N_8884,N_8683);
nor U9372 (N_9372,N_8739,N_8856);
xnor U9373 (N_9373,N_8889,N_8749);
nor U9374 (N_9374,N_8804,N_8784);
and U9375 (N_9375,N_8836,N_8547);
nor U9376 (N_9376,N_8878,N_8777);
xnor U9377 (N_9377,N_8647,N_8821);
and U9378 (N_9378,N_8656,N_8665);
xnor U9379 (N_9379,N_8888,N_8909);
nor U9380 (N_9380,N_8672,N_8849);
and U9381 (N_9381,N_8922,N_8761);
nor U9382 (N_9382,N_8500,N_8933);
nand U9383 (N_9383,N_8844,N_8999);
nor U9384 (N_9384,N_8874,N_8709);
and U9385 (N_9385,N_8928,N_8796);
nand U9386 (N_9386,N_8884,N_8827);
nor U9387 (N_9387,N_8633,N_8660);
nor U9388 (N_9388,N_8640,N_8553);
nand U9389 (N_9389,N_8964,N_8589);
or U9390 (N_9390,N_8602,N_8777);
nand U9391 (N_9391,N_8740,N_8633);
xor U9392 (N_9392,N_8569,N_8834);
nand U9393 (N_9393,N_8571,N_8747);
nand U9394 (N_9394,N_8982,N_8579);
xor U9395 (N_9395,N_8811,N_8541);
and U9396 (N_9396,N_8694,N_8743);
nor U9397 (N_9397,N_8558,N_8900);
or U9398 (N_9398,N_8745,N_8817);
xnor U9399 (N_9399,N_8786,N_8761);
nand U9400 (N_9400,N_8708,N_8599);
nand U9401 (N_9401,N_8515,N_8714);
nand U9402 (N_9402,N_8628,N_8874);
or U9403 (N_9403,N_8880,N_8871);
and U9404 (N_9404,N_8714,N_8729);
and U9405 (N_9405,N_8608,N_8790);
or U9406 (N_9406,N_8609,N_8623);
nand U9407 (N_9407,N_8798,N_8885);
xor U9408 (N_9408,N_8910,N_8641);
nor U9409 (N_9409,N_8974,N_8543);
nand U9410 (N_9410,N_8579,N_8654);
and U9411 (N_9411,N_8616,N_8828);
and U9412 (N_9412,N_8613,N_8570);
nand U9413 (N_9413,N_8865,N_8574);
and U9414 (N_9414,N_8505,N_8715);
nor U9415 (N_9415,N_8827,N_8787);
and U9416 (N_9416,N_8516,N_8630);
nor U9417 (N_9417,N_8997,N_8883);
or U9418 (N_9418,N_8995,N_8848);
and U9419 (N_9419,N_8550,N_8836);
and U9420 (N_9420,N_8990,N_8818);
or U9421 (N_9421,N_8792,N_8838);
and U9422 (N_9422,N_8705,N_8576);
or U9423 (N_9423,N_8630,N_8824);
and U9424 (N_9424,N_8606,N_8544);
and U9425 (N_9425,N_8582,N_8640);
nand U9426 (N_9426,N_8976,N_8768);
or U9427 (N_9427,N_8507,N_8858);
nor U9428 (N_9428,N_8801,N_8907);
or U9429 (N_9429,N_8739,N_8570);
nor U9430 (N_9430,N_8549,N_8861);
nor U9431 (N_9431,N_8842,N_8912);
and U9432 (N_9432,N_8628,N_8728);
or U9433 (N_9433,N_8812,N_8852);
nand U9434 (N_9434,N_8562,N_8604);
or U9435 (N_9435,N_8756,N_8802);
nand U9436 (N_9436,N_8677,N_8800);
and U9437 (N_9437,N_8932,N_8805);
or U9438 (N_9438,N_8797,N_8653);
and U9439 (N_9439,N_8685,N_8747);
xnor U9440 (N_9440,N_8564,N_8777);
nor U9441 (N_9441,N_8822,N_8677);
xor U9442 (N_9442,N_8780,N_8645);
xnor U9443 (N_9443,N_8559,N_8729);
xnor U9444 (N_9444,N_8784,N_8819);
or U9445 (N_9445,N_8917,N_8841);
xnor U9446 (N_9446,N_8585,N_8888);
xor U9447 (N_9447,N_8966,N_8814);
and U9448 (N_9448,N_8664,N_8744);
or U9449 (N_9449,N_8728,N_8986);
and U9450 (N_9450,N_8917,N_8719);
nor U9451 (N_9451,N_8862,N_8501);
xnor U9452 (N_9452,N_8704,N_8578);
and U9453 (N_9453,N_8991,N_8707);
xnor U9454 (N_9454,N_8642,N_8938);
nand U9455 (N_9455,N_8775,N_8904);
and U9456 (N_9456,N_8717,N_8682);
nand U9457 (N_9457,N_8567,N_8608);
xnor U9458 (N_9458,N_8926,N_8773);
and U9459 (N_9459,N_8901,N_8643);
xor U9460 (N_9460,N_8515,N_8684);
nand U9461 (N_9461,N_8664,N_8643);
nor U9462 (N_9462,N_8936,N_8669);
and U9463 (N_9463,N_8517,N_8507);
or U9464 (N_9464,N_8757,N_8721);
nand U9465 (N_9465,N_8936,N_8712);
xor U9466 (N_9466,N_8975,N_8902);
and U9467 (N_9467,N_8709,N_8802);
and U9468 (N_9468,N_8834,N_8865);
nand U9469 (N_9469,N_8641,N_8739);
nand U9470 (N_9470,N_8804,N_8509);
xnor U9471 (N_9471,N_8535,N_8565);
or U9472 (N_9472,N_8631,N_8666);
nor U9473 (N_9473,N_8667,N_8993);
nand U9474 (N_9474,N_8833,N_8893);
xor U9475 (N_9475,N_8984,N_8669);
nor U9476 (N_9476,N_8708,N_8760);
and U9477 (N_9477,N_8668,N_8628);
or U9478 (N_9478,N_8959,N_8720);
nand U9479 (N_9479,N_8663,N_8846);
and U9480 (N_9480,N_8705,N_8899);
nand U9481 (N_9481,N_8997,N_8773);
or U9482 (N_9482,N_8678,N_8651);
or U9483 (N_9483,N_8909,N_8837);
or U9484 (N_9484,N_8511,N_8971);
and U9485 (N_9485,N_8584,N_8818);
xnor U9486 (N_9486,N_8598,N_8550);
and U9487 (N_9487,N_8568,N_8912);
xor U9488 (N_9488,N_8831,N_8510);
nor U9489 (N_9489,N_8826,N_8646);
nor U9490 (N_9490,N_8769,N_8573);
or U9491 (N_9491,N_8993,N_8791);
or U9492 (N_9492,N_8946,N_8943);
nor U9493 (N_9493,N_8511,N_8654);
nor U9494 (N_9494,N_8835,N_8655);
nor U9495 (N_9495,N_8878,N_8771);
nor U9496 (N_9496,N_8701,N_8582);
xnor U9497 (N_9497,N_8766,N_8836);
nand U9498 (N_9498,N_8585,N_8705);
nor U9499 (N_9499,N_8873,N_8831);
and U9500 (N_9500,N_9148,N_9125);
or U9501 (N_9501,N_9177,N_9365);
and U9502 (N_9502,N_9460,N_9438);
nand U9503 (N_9503,N_9263,N_9088);
nand U9504 (N_9504,N_9035,N_9222);
xnor U9505 (N_9505,N_9433,N_9131);
or U9506 (N_9506,N_9332,N_9347);
or U9507 (N_9507,N_9108,N_9363);
or U9508 (N_9508,N_9297,N_9368);
nand U9509 (N_9509,N_9086,N_9259);
or U9510 (N_9510,N_9164,N_9271);
and U9511 (N_9511,N_9009,N_9060);
and U9512 (N_9512,N_9380,N_9243);
or U9513 (N_9513,N_9483,N_9132);
and U9514 (N_9514,N_9495,N_9450);
or U9515 (N_9515,N_9190,N_9016);
nand U9516 (N_9516,N_9296,N_9264);
nand U9517 (N_9517,N_9270,N_9019);
xor U9518 (N_9518,N_9150,N_9452);
or U9519 (N_9519,N_9074,N_9487);
or U9520 (N_9520,N_9492,N_9135);
or U9521 (N_9521,N_9283,N_9308);
or U9522 (N_9522,N_9012,N_9289);
xnor U9523 (N_9523,N_9493,N_9003);
and U9524 (N_9524,N_9099,N_9298);
or U9525 (N_9525,N_9344,N_9302);
nor U9526 (N_9526,N_9025,N_9423);
xnor U9527 (N_9527,N_9334,N_9322);
xor U9528 (N_9528,N_9171,N_9402);
and U9529 (N_9529,N_9077,N_9038);
nand U9530 (N_9530,N_9370,N_9191);
and U9531 (N_9531,N_9040,N_9045);
and U9532 (N_9532,N_9189,N_9217);
nand U9533 (N_9533,N_9142,N_9482);
or U9534 (N_9534,N_9138,N_9096);
nand U9535 (N_9535,N_9439,N_9230);
and U9536 (N_9536,N_9239,N_9497);
or U9537 (N_9537,N_9319,N_9382);
and U9538 (N_9538,N_9377,N_9247);
nand U9539 (N_9539,N_9024,N_9202);
or U9540 (N_9540,N_9371,N_9224);
and U9541 (N_9541,N_9237,N_9461);
xnor U9542 (N_9542,N_9268,N_9213);
nor U9543 (N_9543,N_9220,N_9246);
nand U9544 (N_9544,N_9267,N_9105);
nand U9545 (N_9545,N_9093,N_9122);
xnor U9546 (N_9546,N_9185,N_9391);
and U9547 (N_9547,N_9133,N_9345);
or U9548 (N_9548,N_9199,N_9203);
or U9549 (N_9549,N_9274,N_9144);
xnor U9550 (N_9550,N_9485,N_9329);
nor U9551 (N_9551,N_9219,N_9136);
nand U9552 (N_9552,N_9376,N_9429);
xnor U9553 (N_9553,N_9078,N_9094);
or U9554 (N_9554,N_9355,N_9435);
and U9555 (N_9555,N_9163,N_9292);
or U9556 (N_9556,N_9303,N_9468);
nand U9557 (N_9557,N_9392,N_9054);
and U9558 (N_9558,N_9321,N_9113);
nor U9559 (N_9559,N_9462,N_9470);
xor U9560 (N_9560,N_9436,N_9286);
nand U9561 (N_9561,N_9425,N_9408);
xnor U9562 (N_9562,N_9258,N_9260);
or U9563 (N_9563,N_9159,N_9021);
and U9564 (N_9564,N_9106,N_9097);
xor U9565 (N_9565,N_9427,N_9070);
or U9566 (N_9566,N_9162,N_9204);
or U9567 (N_9567,N_9188,N_9001);
xnor U9568 (N_9568,N_9489,N_9445);
nand U9569 (N_9569,N_9410,N_9112);
or U9570 (N_9570,N_9442,N_9103);
nor U9571 (N_9571,N_9479,N_9053);
or U9572 (N_9572,N_9422,N_9209);
nor U9573 (N_9573,N_9323,N_9228);
or U9574 (N_9574,N_9212,N_9290);
or U9575 (N_9575,N_9172,N_9140);
and U9576 (N_9576,N_9169,N_9250);
nor U9577 (N_9577,N_9201,N_9284);
or U9578 (N_9578,N_9179,N_9387);
xnor U9579 (N_9579,N_9065,N_9279);
xor U9580 (N_9580,N_9475,N_9057);
xnor U9581 (N_9581,N_9134,N_9362);
or U9582 (N_9582,N_9155,N_9328);
xor U9583 (N_9583,N_9165,N_9443);
or U9584 (N_9584,N_9313,N_9197);
nand U9585 (N_9585,N_9018,N_9282);
and U9586 (N_9586,N_9413,N_9490);
xor U9587 (N_9587,N_9359,N_9110);
nand U9588 (N_9588,N_9488,N_9406);
nor U9589 (N_9589,N_9013,N_9364);
xor U9590 (N_9590,N_9494,N_9366);
or U9591 (N_9591,N_9389,N_9076);
nand U9592 (N_9592,N_9272,N_9111);
nand U9593 (N_9593,N_9154,N_9457);
or U9594 (N_9594,N_9466,N_9360);
or U9595 (N_9595,N_9027,N_9152);
or U9596 (N_9596,N_9474,N_9415);
and U9597 (N_9597,N_9449,N_9463);
and U9598 (N_9598,N_9428,N_9225);
xor U9599 (N_9599,N_9249,N_9081);
nand U9600 (N_9600,N_9126,N_9255);
nor U9601 (N_9601,N_9396,N_9398);
nand U9602 (N_9602,N_9030,N_9304);
xor U9603 (N_9603,N_9052,N_9102);
and U9604 (N_9604,N_9000,N_9129);
nand U9605 (N_9605,N_9346,N_9399);
nor U9606 (N_9606,N_9198,N_9299);
or U9607 (N_9607,N_9278,N_9082);
and U9608 (N_9608,N_9193,N_9014);
xnor U9609 (N_9609,N_9033,N_9234);
xnor U9610 (N_9610,N_9405,N_9119);
xnor U9611 (N_9611,N_9208,N_9448);
nor U9612 (N_9612,N_9083,N_9343);
nand U9613 (N_9613,N_9395,N_9161);
nand U9614 (N_9614,N_9117,N_9262);
nand U9615 (N_9615,N_9248,N_9307);
nand U9616 (N_9616,N_9068,N_9352);
nor U9617 (N_9617,N_9301,N_9409);
and U9618 (N_9618,N_9273,N_9420);
nor U9619 (N_9619,N_9090,N_9192);
or U9620 (N_9620,N_9098,N_9058);
nor U9621 (N_9621,N_9095,N_9059);
and U9622 (N_9622,N_9369,N_9484);
nand U9623 (N_9623,N_9141,N_9238);
or U9624 (N_9624,N_9156,N_9374);
xnor U9625 (N_9625,N_9062,N_9087);
and U9626 (N_9626,N_9143,N_9472);
nor U9627 (N_9627,N_9338,N_9080);
nand U9628 (N_9628,N_9048,N_9491);
and U9629 (N_9629,N_9256,N_9128);
or U9630 (N_9630,N_9123,N_9269);
nor U9631 (N_9631,N_9206,N_9385);
nand U9632 (N_9632,N_9381,N_9455);
nand U9633 (N_9633,N_9039,N_9372);
and U9634 (N_9634,N_9180,N_9157);
nand U9635 (N_9635,N_9186,N_9431);
nand U9636 (N_9636,N_9316,N_9240);
xor U9637 (N_9637,N_9022,N_9046);
nand U9638 (N_9638,N_9049,N_9418);
or U9639 (N_9639,N_9404,N_9215);
and U9640 (N_9640,N_9235,N_9383);
xor U9641 (N_9641,N_9459,N_9465);
and U9642 (N_9642,N_9414,N_9416);
xnor U9643 (N_9643,N_9244,N_9451);
nand U9644 (N_9644,N_9378,N_9348);
nor U9645 (N_9645,N_9139,N_9432);
nand U9646 (N_9646,N_9178,N_9417);
and U9647 (N_9647,N_9454,N_9285);
and U9648 (N_9648,N_9388,N_9453);
and U9649 (N_9649,N_9107,N_9333);
xnor U9650 (N_9650,N_9486,N_9480);
nor U9651 (N_9651,N_9120,N_9124);
nand U9652 (N_9652,N_9075,N_9275);
nand U9653 (N_9653,N_9358,N_9341);
and U9654 (N_9654,N_9481,N_9421);
or U9655 (N_9655,N_9373,N_9187);
nand U9656 (N_9656,N_9444,N_9434);
nor U9657 (N_9657,N_9261,N_9073);
or U9658 (N_9658,N_9056,N_9147);
xnor U9659 (N_9659,N_9233,N_9069);
or U9660 (N_9660,N_9393,N_9335);
and U9661 (N_9661,N_9175,N_9194);
or U9662 (N_9662,N_9477,N_9200);
xor U9663 (N_9663,N_9280,N_9288);
nand U9664 (N_9664,N_9079,N_9310);
xor U9665 (N_9665,N_9166,N_9085);
nor U9666 (N_9666,N_9253,N_9170);
nor U9667 (N_9667,N_9214,N_9337);
xor U9668 (N_9668,N_9036,N_9023);
or U9669 (N_9669,N_9211,N_9205);
or U9670 (N_9670,N_9309,N_9361);
or U9671 (N_9671,N_9037,N_9181);
nor U9672 (N_9672,N_9456,N_9340);
and U9673 (N_9673,N_9447,N_9017);
or U9674 (N_9674,N_9121,N_9051);
or U9675 (N_9675,N_9311,N_9407);
nor U9676 (N_9676,N_9061,N_9050);
nand U9677 (N_9677,N_9160,N_9379);
nand U9678 (N_9678,N_9458,N_9227);
or U9679 (N_9679,N_9331,N_9092);
and U9680 (N_9680,N_9118,N_9357);
nor U9681 (N_9681,N_9218,N_9067);
or U9682 (N_9682,N_9294,N_9401);
nor U9683 (N_9683,N_9412,N_9020);
nor U9684 (N_9684,N_9008,N_9446);
or U9685 (N_9685,N_9029,N_9173);
or U9686 (N_9686,N_9104,N_9295);
nor U9687 (N_9687,N_9047,N_9471);
or U9688 (N_9688,N_9252,N_9114);
xnor U9689 (N_9689,N_9183,N_9390);
xor U9690 (N_9690,N_9089,N_9276);
and U9691 (N_9691,N_9216,N_9440);
xnor U9692 (N_9692,N_9031,N_9137);
xor U9693 (N_9693,N_9010,N_9498);
nor U9694 (N_9694,N_9293,N_9127);
and U9695 (N_9695,N_9257,N_9320);
xor U9696 (N_9696,N_9091,N_9207);
nor U9697 (N_9697,N_9317,N_9291);
nor U9698 (N_9698,N_9349,N_9026);
nand U9699 (N_9699,N_9375,N_9149);
nor U9700 (N_9700,N_9354,N_9426);
and U9701 (N_9701,N_9318,N_9007);
nand U9702 (N_9702,N_9315,N_9330);
xor U9703 (N_9703,N_9100,N_9245);
nand U9704 (N_9704,N_9351,N_9015);
nand U9705 (N_9705,N_9336,N_9353);
nand U9706 (N_9706,N_9281,N_9116);
and U9707 (N_9707,N_9242,N_9419);
nor U9708 (N_9708,N_9305,N_9437);
and U9709 (N_9709,N_9394,N_9071);
or U9710 (N_9710,N_9044,N_9063);
and U9711 (N_9711,N_9006,N_9226);
and U9712 (N_9712,N_9195,N_9174);
or U9713 (N_9713,N_9032,N_9241);
nand U9714 (N_9714,N_9084,N_9251);
nor U9715 (N_9715,N_9145,N_9397);
nor U9716 (N_9716,N_9055,N_9478);
nand U9717 (N_9717,N_9011,N_9034);
nand U9718 (N_9718,N_9499,N_9064);
and U9719 (N_9719,N_9042,N_9411);
nor U9720 (N_9720,N_9004,N_9384);
and U9721 (N_9721,N_9167,N_9356);
or U9722 (N_9722,N_9158,N_9314);
nand U9723 (N_9723,N_9130,N_9496);
nor U9724 (N_9724,N_9287,N_9367);
or U9725 (N_9725,N_9231,N_9469);
and U9726 (N_9726,N_9182,N_9430);
or U9727 (N_9727,N_9400,N_9342);
nor U9728 (N_9728,N_9386,N_9254);
xnor U9729 (N_9729,N_9043,N_9151);
and U9730 (N_9730,N_9176,N_9300);
xor U9731 (N_9731,N_9476,N_9168);
or U9732 (N_9732,N_9115,N_9306);
and U9733 (N_9733,N_9326,N_9350);
and U9734 (N_9734,N_9232,N_9153);
xor U9735 (N_9735,N_9184,N_9146);
and U9736 (N_9736,N_9002,N_9464);
xor U9737 (N_9737,N_9441,N_9265);
and U9738 (N_9738,N_9066,N_9109);
xor U9739 (N_9739,N_9312,N_9072);
xnor U9740 (N_9740,N_9424,N_9339);
or U9741 (N_9741,N_9028,N_9221);
or U9742 (N_9742,N_9324,N_9101);
nor U9743 (N_9743,N_9266,N_9325);
nand U9744 (N_9744,N_9236,N_9473);
nand U9745 (N_9745,N_9277,N_9005);
nand U9746 (N_9746,N_9327,N_9229);
xnor U9747 (N_9747,N_9196,N_9041);
or U9748 (N_9748,N_9467,N_9403);
nor U9749 (N_9749,N_9210,N_9223);
or U9750 (N_9750,N_9144,N_9196);
xnor U9751 (N_9751,N_9176,N_9431);
or U9752 (N_9752,N_9426,N_9310);
nor U9753 (N_9753,N_9295,N_9083);
and U9754 (N_9754,N_9236,N_9182);
or U9755 (N_9755,N_9301,N_9396);
nand U9756 (N_9756,N_9130,N_9442);
nor U9757 (N_9757,N_9147,N_9251);
xnor U9758 (N_9758,N_9039,N_9310);
and U9759 (N_9759,N_9130,N_9415);
nor U9760 (N_9760,N_9372,N_9134);
and U9761 (N_9761,N_9338,N_9208);
and U9762 (N_9762,N_9372,N_9207);
or U9763 (N_9763,N_9421,N_9422);
nand U9764 (N_9764,N_9450,N_9447);
nor U9765 (N_9765,N_9050,N_9241);
xnor U9766 (N_9766,N_9161,N_9102);
nor U9767 (N_9767,N_9217,N_9148);
nand U9768 (N_9768,N_9252,N_9020);
nor U9769 (N_9769,N_9136,N_9383);
xnor U9770 (N_9770,N_9034,N_9073);
nor U9771 (N_9771,N_9083,N_9086);
nand U9772 (N_9772,N_9219,N_9267);
and U9773 (N_9773,N_9356,N_9347);
or U9774 (N_9774,N_9337,N_9180);
nor U9775 (N_9775,N_9001,N_9322);
or U9776 (N_9776,N_9096,N_9183);
xnor U9777 (N_9777,N_9247,N_9033);
or U9778 (N_9778,N_9271,N_9396);
or U9779 (N_9779,N_9478,N_9336);
and U9780 (N_9780,N_9092,N_9482);
nand U9781 (N_9781,N_9433,N_9362);
xor U9782 (N_9782,N_9266,N_9082);
and U9783 (N_9783,N_9138,N_9129);
nor U9784 (N_9784,N_9012,N_9232);
xor U9785 (N_9785,N_9094,N_9432);
nor U9786 (N_9786,N_9044,N_9417);
nand U9787 (N_9787,N_9415,N_9056);
nand U9788 (N_9788,N_9202,N_9042);
or U9789 (N_9789,N_9100,N_9121);
and U9790 (N_9790,N_9395,N_9401);
or U9791 (N_9791,N_9259,N_9429);
and U9792 (N_9792,N_9473,N_9445);
xor U9793 (N_9793,N_9226,N_9172);
xor U9794 (N_9794,N_9445,N_9300);
and U9795 (N_9795,N_9289,N_9128);
xnor U9796 (N_9796,N_9285,N_9098);
and U9797 (N_9797,N_9381,N_9433);
or U9798 (N_9798,N_9496,N_9452);
xnor U9799 (N_9799,N_9446,N_9289);
or U9800 (N_9800,N_9149,N_9204);
nand U9801 (N_9801,N_9397,N_9135);
xor U9802 (N_9802,N_9428,N_9101);
or U9803 (N_9803,N_9001,N_9150);
xor U9804 (N_9804,N_9054,N_9442);
xnor U9805 (N_9805,N_9489,N_9340);
nor U9806 (N_9806,N_9409,N_9112);
nand U9807 (N_9807,N_9313,N_9329);
xor U9808 (N_9808,N_9222,N_9166);
or U9809 (N_9809,N_9281,N_9494);
nand U9810 (N_9810,N_9460,N_9379);
nor U9811 (N_9811,N_9210,N_9379);
nand U9812 (N_9812,N_9377,N_9065);
or U9813 (N_9813,N_9443,N_9037);
and U9814 (N_9814,N_9292,N_9380);
nor U9815 (N_9815,N_9185,N_9470);
nand U9816 (N_9816,N_9206,N_9187);
nor U9817 (N_9817,N_9350,N_9134);
xnor U9818 (N_9818,N_9185,N_9407);
or U9819 (N_9819,N_9284,N_9493);
xor U9820 (N_9820,N_9126,N_9343);
xnor U9821 (N_9821,N_9275,N_9189);
xor U9822 (N_9822,N_9255,N_9235);
nor U9823 (N_9823,N_9327,N_9010);
and U9824 (N_9824,N_9375,N_9210);
xor U9825 (N_9825,N_9135,N_9132);
xor U9826 (N_9826,N_9405,N_9253);
xor U9827 (N_9827,N_9429,N_9476);
nor U9828 (N_9828,N_9243,N_9484);
and U9829 (N_9829,N_9099,N_9211);
xor U9830 (N_9830,N_9320,N_9393);
and U9831 (N_9831,N_9126,N_9415);
or U9832 (N_9832,N_9081,N_9281);
and U9833 (N_9833,N_9290,N_9045);
or U9834 (N_9834,N_9299,N_9339);
and U9835 (N_9835,N_9017,N_9450);
nand U9836 (N_9836,N_9063,N_9474);
xnor U9837 (N_9837,N_9270,N_9188);
nor U9838 (N_9838,N_9068,N_9107);
and U9839 (N_9839,N_9378,N_9187);
nor U9840 (N_9840,N_9499,N_9172);
nor U9841 (N_9841,N_9096,N_9025);
and U9842 (N_9842,N_9361,N_9214);
nor U9843 (N_9843,N_9015,N_9064);
and U9844 (N_9844,N_9042,N_9492);
xor U9845 (N_9845,N_9039,N_9158);
nor U9846 (N_9846,N_9264,N_9386);
nor U9847 (N_9847,N_9263,N_9245);
nor U9848 (N_9848,N_9344,N_9154);
nand U9849 (N_9849,N_9173,N_9347);
xor U9850 (N_9850,N_9330,N_9020);
xor U9851 (N_9851,N_9190,N_9012);
or U9852 (N_9852,N_9475,N_9272);
or U9853 (N_9853,N_9038,N_9020);
or U9854 (N_9854,N_9286,N_9332);
nand U9855 (N_9855,N_9359,N_9130);
or U9856 (N_9856,N_9249,N_9263);
nand U9857 (N_9857,N_9081,N_9049);
nand U9858 (N_9858,N_9039,N_9252);
nand U9859 (N_9859,N_9093,N_9435);
or U9860 (N_9860,N_9265,N_9289);
nor U9861 (N_9861,N_9247,N_9050);
or U9862 (N_9862,N_9456,N_9279);
nor U9863 (N_9863,N_9380,N_9297);
nor U9864 (N_9864,N_9388,N_9076);
and U9865 (N_9865,N_9051,N_9391);
and U9866 (N_9866,N_9014,N_9205);
and U9867 (N_9867,N_9422,N_9302);
and U9868 (N_9868,N_9039,N_9453);
xnor U9869 (N_9869,N_9230,N_9367);
nor U9870 (N_9870,N_9072,N_9426);
nand U9871 (N_9871,N_9332,N_9436);
xor U9872 (N_9872,N_9018,N_9496);
xor U9873 (N_9873,N_9401,N_9363);
or U9874 (N_9874,N_9279,N_9039);
or U9875 (N_9875,N_9142,N_9386);
and U9876 (N_9876,N_9419,N_9483);
and U9877 (N_9877,N_9082,N_9239);
and U9878 (N_9878,N_9192,N_9275);
and U9879 (N_9879,N_9106,N_9439);
nor U9880 (N_9880,N_9140,N_9193);
xor U9881 (N_9881,N_9134,N_9387);
nand U9882 (N_9882,N_9120,N_9235);
xor U9883 (N_9883,N_9088,N_9440);
nand U9884 (N_9884,N_9352,N_9018);
or U9885 (N_9885,N_9020,N_9146);
nand U9886 (N_9886,N_9371,N_9262);
nand U9887 (N_9887,N_9354,N_9218);
xnor U9888 (N_9888,N_9218,N_9321);
nor U9889 (N_9889,N_9466,N_9379);
nand U9890 (N_9890,N_9033,N_9212);
xor U9891 (N_9891,N_9037,N_9310);
or U9892 (N_9892,N_9151,N_9345);
and U9893 (N_9893,N_9495,N_9435);
nor U9894 (N_9894,N_9001,N_9100);
or U9895 (N_9895,N_9441,N_9454);
and U9896 (N_9896,N_9069,N_9280);
or U9897 (N_9897,N_9409,N_9277);
nor U9898 (N_9898,N_9324,N_9373);
nor U9899 (N_9899,N_9202,N_9320);
or U9900 (N_9900,N_9336,N_9150);
and U9901 (N_9901,N_9412,N_9228);
nand U9902 (N_9902,N_9332,N_9416);
nor U9903 (N_9903,N_9182,N_9209);
and U9904 (N_9904,N_9322,N_9373);
nor U9905 (N_9905,N_9092,N_9143);
xnor U9906 (N_9906,N_9360,N_9022);
and U9907 (N_9907,N_9397,N_9073);
and U9908 (N_9908,N_9407,N_9494);
xnor U9909 (N_9909,N_9453,N_9394);
and U9910 (N_9910,N_9034,N_9435);
nor U9911 (N_9911,N_9321,N_9016);
xnor U9912 (N_9912,N_9468,N_9472);
and U9913 (N_9913,N_9137,N_9184);
or U9914 (N_9914,N_9124,N_9406);
xnor U9915 (N_9915,N_9207,N_9065);
nand U9916 (N_9916,N_9385,N_9182);
xnor U9917 (N_9917,N_9474,N_9235);
nor U9918 (N_9918,N_9246,N_9337);
or U9919 (N_9919,N_9224,N_9123);
and U9920 (N_9920,N_9469,N_9228);
and U9921 (N_9921,N_9003,N_9025);
nor U9922 (N_9922,N_9330,N_9304);
and U9923 (N_9923,N_9059,N_9319);
or U9924 (N_9924,N_9230,N_9380);
nor U9925 (N_9925,N_9013,N_9258);
nor U9926 (N_9926,N_9058,N_9486);
or U9927 (N_9927,N_9166,N_9405);
nand U9928 (N_9928,N_9017,N_9283);
or U9929 (N_9929,N_9334,N_9422);
nor U9930 (N_9930,N_9363,N_9031);
or U9931 (N_9931,N_9493,N_9108);
nand U9932 (N_9932,N_9364,N_9285);
xnor U9933 (N_9933,N_9200,N_9391);
and U9934 (N_9934,N_9095,N_9028);
or U9935 (N_9935,N_9193,N_9327);
nand U9936 (N_9936,N_9025,N_9435);
nor U9937 (N_9937,N_9250,N_9102);
or U9938 (N_9938,N_9416,N_9273);
nand U9939 (N_9939,N_9477,N_9085);
and U9940 (N_9940,N_9424,N_9215);
xor U9941 (N_9941,N_9084,N_9466);
xor U9942 (N_9942,N_9052,N_9353);
nor U9943 (N_9943,N_9164,N_9435);
xor U9944 (N_9944,N_9185,N_9010);
xnor U9945 (N_9945,N_9317,N_9067);
nor U9946 (N_9946,N_9447,N_9372);
nor U9947 (N_9947,N_9349,N_9377);
or U9948 (N_9948,N_9089,N_9188);
nand U9949 (N_9949,N_9141,N_9483);
or U9950 (N_9950,N_9496,N_9294);
xnor U9951 (N_9951,N_9103,N_9135);
nand U9952 (N_9952,N_9108,N_9076);
or U9953 (N_9953,N_9393,N_9087);
and U9954 (N_9954,N_9356,N_9360);
xnor U9955 (N_9955,N_9355,N_9139);
nor U9956 (N_9956,N_9243,N_9060);
nand U9957 (N_9957,N_9079,N_9440);
nand U9958 (N_9958,N_9190,N_9207);
nor U9959 (N_9959,N_9194,N_9063);
xnor U9960 (N_9960,N_9227,N_9457);
and U9961 (N_9961,N_9382,N_9291);
and U9962 (N_9962,N_9489,N_9300);
nor U9963 (N_9963,N_9329,N_9434);
and U9964 (N_9964,N_9349,N_9483);
xor U9965 (N_9965,N_9369,N_9062);
nor U9966 (N_9966,N_9218,N_9134);
xor U9967 (N_9967,N_9483,N_9398);
xor U9968 (N_9968,N_9223,N_9418);
nor U9969 (N_9969,N_9147,N_9185);
or U9970 (N_9970,N_9254,N_9186);
or U9971 (N_9971,N_9019,N_9428);
nand U9972 (N_9972,N_9037,N_9314);
or U9973 (N_9973,N_9069,N_9299);
nand U9974 (N_9974,N_9316,N_9457);
or U9975 (N_9975,N_9141,N_9269);
or U9976 (N_9976,N_9413,N_9021);
and U9977 (N_9977,N_9143,N_9410);
and U9978 (N_9978,N_9198,N_9359);
and U9979 (N_9979,N_9470,N_9214);
nand U9980 (N_9980,N_9476,N_9138);
nand U9981 (N_9981,N_9024,N_9476);
nand U9982 (N_9982,N_9011,N_9097);
nor U9983 (N_9983,N_9263,N_9462);
xnor U9984 (N_9984,N_9141,N_9267);
and U9985 (N_9985,N_9249,N_9356);
and U9986 (N_9986,N_9141,N_9201);
and U9987 (N_9987,N_9017,N_9212);
and U9988 (N_9988,N_9214,N_9183);
or U9989 (N_9989,N_9319,N_9318);
and U9990 (N_9990,N_9119,N_9028);
nand U9991 (N_9991,N_9200,N_9345);
nand U9992 (N_9992,N_9249,N_9272);
and U9993 (N_9993,N_9350,N_9157);
or U9994 (N_9994,N_9244,N_9398);
nor U9995 (N_9995,N_9364,N_9205);
and U9996 (N_9996,N_9180,N_9447);
xnor U9997 (N_9997,N_9390,N_9004);
xnor U9998 (N_9998,N_9159,N_9066);
or U9999 (N_9999,N_9401,N_9406);
and U10000 (N_10000,N_9636,N_9564);
nand U10001 (N_10001,N_9551,N_9709);
nor U10002 (N_10002,N_9622,N_9864);
and U10003 (N_10003,N_9582,N_9578);
nand U10004 (N_10004,N_9653,N_9510);
and U10005 (N_10005,N_9832,N_9612);
and U10006 (N_10006,N_9581,N_9735);
xor U10007 (N_10007,N_9856,N_9773);
or U10008 (N_10008,N_9512,N_9802);
nand U10009 (N_10009,N_9809,N_9794);
and U10010 (N_10010,N_9952,N_9939);
or U10011 (N_10011,N_9865,N_9876);
xnor U10012 (N_10012,N_9772,N_9786);
nor U10013 (N_10013,N_9693,N_9732);
or U10014 (N_10014,N_9689,N_9758);
xor U10015 (N_10015,N_9966,N_9765);
xor U10016 (N_10016,N_9590,N_9515);
nand U10017 (N_10017,N_9897,N_9924);
nand U10018 (N_10018,N_9671,N_9766);
nand U10019 (N_10019,N_9894,N_9635);
xor U10020 (N_10020,N_9533,N_9759);
nand U10021 (N_10021,N_9921,N_9988);
and U10022 (N_10022,N_9630,N_9841);
nor U10023 (N_10023,N_9613,N_9669);
nor U10024 (N_10024,N_9995,N_9906);
and U10025 (N_10025,N_9568,N_9545);
xor U10026 (N_10026,N_9723,N_9609);
nand U10027 (N_10027,N_9827,N_9690);
nand U10028 (N_10028,N_9826,N_9900);
and U10029 (N_10029,N_9695,N_9987);
nor U10030 (N_10030,N_9985,N_9867);
and U10031 (N_10031,N_9840,N_9945);
and U10032 (N_10032,N_9925,N_9784);
xor U10033 (N_10033,N_9508,N_9909);
xor U10034 (N_10034,N_9598,N_9678);
nand U10035 (N_10035,N_9757,N_9775);
nand U10036 (N_10036,N_9806,N_9659);
nor U10037 (N_10037,N_9778,N_9654);
or U10038 (N_10038,N_9641,N_9628);
nor U10039 (N_10039,N_9926,N_9594);
nor U10040 (N_10040,N_9792,N_9623);
xnor U10041 (N_10041,N_9937,N_9569);
and U10042 (N_10042,N_9661,N_9575);
and U10043 (N_10043,N_9696,N_9991);
and U10044 (N_10044,N_9566,N_9767);
or U10045 (N_10045,N_9965,N_9514);
and U10046 (N_10046,N_9591,N_9912);
xnor U10047 (N_10047,N_9842,N_9592);
nand U10048 (N_10048,N_9729,N_9934);
nor U10049 (N_10049,N_9700,N_9951);
nand U10050 (N_10050,N_9740,N_9670);
and U10051 (N_10051,N_9871,N_9500);
xnor U10052 (N_10052,N_9764,N_9969);
and U10053 (N_10053,N_9967,N_9577);
and U10054 (N_10054,N_9873,N_9632);
and U10055 (N_10055,N_9953,N_9916);
nand U10056 (N_10056,N_9721,N_9529);
nand U10057 (N_10057,N_9583,N_9717);
nand U10058 (N_10058,N_9790,N_9895);
or U10059 (N_10059,N_9535,N_9823);
and U10060 (N_10060,N_9703,N_9844);
nor U10061 (N_10061,N_9797,N_9960);
or U10062 (N_10062,N_9676,N_9686);
nand U10063 (N_10063,N_9893,N_9885);
xor U10064 (N_10064,N_9640,N_9989);
or U10065 (N_10065,N_9933,N_9907);
or U10066 (N_10066,N_9993,N_9940);
xor U10067 (N_10067,N_9996,N_9610);
nand U10068 (N_10068,N_9601,N_9860);
xor U10069 (N_10069,N_9663,N_9714);
and U10070 (N_10070,N_9847,N_9702);
nand U10071 (N_10071,N_9611,N_9616);
nor U10072 (N_10072,N_9553,N_9785);
and U10073 (N_10073,N_9980,N_9911);
nor U10074 (N_10074,N_9532,N_9502);
xor U10075 (N_10075,N_9872,N_9731);
nor U10076 (N_10076,N_9838,N_9970);
nor U10077 (N_10077,N_9959,N_9505);
xnor U10078 (N_10078,N_9923,N_9927);
xor U10079 (N_10079,N_9855,N_9835);
nor U10080 (N_10080,N_9862,N_9585);
nand U10081 (N_10081,N_9803,N_9781);
nor U10082 (N_10082,N_9554,N_9843);
or U10083 (N_10083,N_9990,N_9600);
nor U10084 (N_10084,N_9534,N_9718);
or U10085 (N_10085,N_9683,N_9710);
nor U10086 (N_10086,N_9739,N_9753);
or U10087 (N_10087,N_9536,N_9810);
or U10088 (N_10088,N_9964,N_9537);
and U10089 (N_10089,N_9523,N_9946);
and U10090 (N_10090,N_9639,N_9821);
xnor U10091 (N_10091,N_9874,N_9942);
nand U10092 (N_10092,N_9816,N_9931);
nand U10093 (N_10093,N_9808,N_9620);
nand U10094 (N_10094,N_9530,N_9837);
nor U10095 (N_10095,N_9602,N_9807);
xnor U10096 (N_10096,N_9851,N_9615);
nor U10097 (N_10097,N_9722,N_9800);
nor U10098 (N_10098,N_9643,N_9685);
nand U10099 (N_10099,N_9576,N_9956);
xor U10100 (N_10100,N_9558,N_9813);
or U10101 (N_10101,N_9652,N_9677);
nand U10102 (N_10102,N_9692,N_9517);
xnor U10103 (N_10103,N_9656,N_9928);
or U10104 (N_10104,N_9644,N_9999);
xor U10105 (N_10105,N_9698,N_9579);
and U10106 (N_10106,N_9795,N_9749);
xor U10107 (N_10107,N_9506,N_9662);
and U10108 (N_10108,N_9556,N_9561);
or U10109 (N_10109,N_9978,N_9829);
xnor U10110 (N_10110,N_9540,N_9666);
and U10111 (N_10111,N_9599,N_9550);
nor U10112 (N_10112,N_9948,N_9713);
and U10113 (N_10113,N_9730,N_9848);
nor U10114 (N_10114,N_9762,N_9680);
and U10115 (N_10115,N_9760,N_9646);
nand U10116 (N_10116,N_9629,N_9606);
nand U10117 (N_10117,N_9888,N_9982);
nor U10118 (N_10118,N_9751,N_9504);
and U10119 (N_10119,N_9984,N_9815);
nand U10120 (N_10120,N_9589,N_9527);
or U10121 (N_10121,N_9950,N_9793);
xnor U10122 (N_10122,N_9697,N_9524);
nand U10123 (N_10123,N_9649,N_9746);
or U10124 (N_10124,N_9920,N_9828);
and U10125 (N_10125,N_9801,N_9768);
and U10126 (N_10126,N_9743,N_9830);
nand U10127 (N_10127,N_9846,N_9614);
nand U10128 (N_10128,N_9563,N_9539);
nor U10129 (N_10129,N_9691,N_9892);
xor U10130 (N_10130,N_9910,N_9922);
xor U10131 (N_10131,N_9902,N_9845);
xnor U10132 (N_10132,N_9783,N_9503);
nor U10133 (N_10133,N_9752,N_9675);
xor U10134 (N_10134,N_9889,N_9774);
and U10135 (N_10135,N_9682,N_9555);
nand U10136 (N_10136,N_9549,N_9694);
or U10137 (N_10137,N_9861,N_9998);
xnor U10138 (N_10138,N_9944,N_9918);
xor U10139 (N_10139,N_9771,N_9852);
nor U10140 (N_10140,N_9705,N_9637);
nand U10141 (N_10141,N_9825,N_9604);
and U10142 (N_10142,N_9780,N_9886);
and U10143 (N_10143,N_9595,N_9870);
or U10144 (N_10144,N_9736,N_9777);
xnor U10145 (N_10145,N_9501,N_9586);
and U10146 (N_10146,N_9699,N_9908);
nor U10147 (N_10147,N_9704,N_9706);
or U10148 (N_10148,N_9650,N_9850);
or U10149 (N_10149,N_9858,N_9811);
nor U10150 (N_10150,N_9520,N_9547);
xor U10151 (N_10151,N_9930,N_9932);
nor U10152 (N_10152,N_9727,N_9761);
or U10153 (N_10153,N_9621,N_9805);
or U10154 (N_10154,N_9672,N_9779);
or U10155 (N_10155,N_9839,N_9798);
nand U10156 (N_10156,N_9608,N_9903);
or U10157 (N_10157,N_9943,N_9657);
xor U10158 (N_10158,N_9546,N_9708);
or U10159 (N_10159,N_9726,N_9881);
nor U10160 (N_10160,N_9868,N_9814);
nand U10161 (N_10161,N_9742,N_9603);
nor U10162 (N_10162,N_9804,N_9812);
and U10163 (N_10163,N_9645,N_9716);
nand U10164 (N_10164,N_9770,N_9679);
or U10165 (N_10165,N_9525,N_9979);
and U10166 (N_10166,N_9642,N_9507);
nand U10167 (N_10167,N_9593,N_9914);
and U10168 (N_10168,N_9935,N_9719);
and U10169 (N_10169,N_9552,N_9658);
nand U10170 (N_10170,N_9973,N_9833);
and U10171 (N_10171,N_9791,N_9562);
and U10172 (N_10172,N_9516,N_9559);
nand U10173 (N_10173,N_9531,N_9627);
or U10174 (N_10174,N_9567,N_9882);
or U10175 (N_10175,N_9971,N_9992);
or U10176 (N_10176,N_9941,N_9887);
nor U10177 (N_10177,N_9511,N_9949);
nand U10178 (N_10178,N_9544,N_9631);
nor U10179 (N_10179,N_9607,N_9728);
xnor U10180 (N_10180,N_9880,N_9619);
nor U10181 (N_10181,N_9879,N_9747);
and U10182 (N_10182,N_9681,N_9905);
xor U10183 (N_10183,N_9560,N_9521);
nor U10184 (N_10184,N_9573,N_9854);
or U10185 (N_10185,N_9513,N_9624);
and U10186 (N_10186,N_9597,N_9981);
or U10187 (N_10187,N_9877,N_9557);
nand U10188 (N_10188,N_9660,N_9986);
nand U10189 (N_10189,N_9684,N_9955);
or U10190 (N_10190,N_9711,N_9754);
xor U10191 (N_10191,N_9799,N_9976);
xnor U10192 (N_10192,N_9565,N_9617);
and U10193 (N_10193,N_9542,N_9673);
or U10194 (N_10194,N_9541,N_9822);
nor U10195 (N_10195,N_9929,N_9899);
or U10196 (N_10196,N_9664,N_9518);
or U10197 (N_10197,N_9633,N_9744);
nor U10198 (N_10198,N_9974,N_9947);
and U10199 (N_10199,N_9571,N_9853);
nand U10200 (N_10200,N_9674,N_9519);
and U10201 (N_10201,N_9526,N_9528);
and U10202 (N_10202,N_9548,N_9915);
xor U10203 (N_10203,N_9509,N_9878);
nor U10204 (N_10204,N_9733,N_9574);
xnor U10205 (N_10205,N_9588,N_9638);
nor U10206 (N_10206,N_9712,N_9725);
nand U10207 (N_10207,N_9884,N_9648);
nand U10208 (N_10208,N_9738,N_9667);
nor U10209 (N_10209,N_9818,N_9596);
nor U10210 (N_10210,N_9957,N_9715);
and U10211 (N_10211,N_9625,N_9634);
nand U10212 (N_10212,N_9817,N_9750);
and U10213 (N_10213,N_9572,N_9782);
and U10214 (N_10214,N_9668,N_9788);
or U10215 (N_10215,N_9891,N_9745);
nand U10216 (N_10216,N_9954,N_9580);
nand U10217 (N_10217,N_9836,N_9688);
or U10218 (N_10218,N_9890,N_9824);
and U10219 (N_10219,N_9958,N_9748);
or U10220 (N_10220,N_9522,N_9883);
nor U10221 (N_10221,N_9936,N_9896);
xor U10222 (N_10222,N_9776,N_9570);
nand U10223 (N_10223,N_9831,N_9819);
xor U10224 (N_10224,N_9869,N_9741);
nor U10225 (N_10225,N_9605,N_9737);
xnor U10226 (N_10226,N_9962,N_9834);
and U10227 (N_10227,N_9724,N_9863);
or U10228 (N_10228,N_9787,N_9963);
nor U10229 (N_10229,N_9898,N_9587);
and U10230 (N_10230,N_9618,N_9994);
and U10231 (N_10231,N_9647,N_9720);
and U10232 (N_10232,N_9651,N_9849);
xnor U10233 (N_10233,N_9796,N_9997);
nand U10234 (N_10234,N_9756,N_9901);
nor U10235 (N_10235,N_9734,N_9917);
nor U10236 (N_10236,N_9875,N_9983);
and U10237 (N_10237,N_9859,N_9701);
or U10238 (N_10238,N_9655,N_9913);
or U10239 (N_10239,N_9763,N_9789);
and U10240 (N_10240,N_9626,N_9857);
xor U10241 (N_10241,N_9904,N_9543);
and U10242 (N_10242,N_9972,N_9820);
xnor U10243 (N_10243,N_9968,N_9687);
nand U10244 (N_10244,N_9961,N_9707);
xnor U10245 (N_10245,N_9538,N_9769);
nor U10246 (N_10246,N_9665,N_9755);
and U10247 (N_10247,N_9584,N_9938);
nand U10248 (N_10248,N_9975,N_9919);
or U10249 (N_10249,N_9977,N_9866);
nor U10250 (N_10250,N_9697,N_9712);
nand U10251 (N_10251,N_9502,N_9865);
nand U10252 (N_10252,N_9903,N_9761);
and U10253 (N_10253,N_9504,N_9965);
xor U10254 (N_10254,N_9762,N_9799);
nor U10255 (N_10255,N_9753,N_9922);
or U10256 (N_10256,N_9812,N_9996);
xnor U10257 (N_10257,N_9548,N_9572);
xnor U10258 (N_10258,N_9678,N_9981);
nand U10259 (N_10259,N_9633,N_9616);
nand U10260 (N_10260,N_9899,N_9775);
nand U10261 (N_10261,N_9868,N_9856);
xnor U10262 (N_10262,N_9533,N_9698);
nand U10263 (N_10263,N_9762,N_9963);
xnor U10264 (N_10264,N_9993,N_9938);
nand U10265 (N_10265,N_9859,N_9892);
or U10266 (N_10266,N_9618,N_9696);
or U10267 (N_10267,N_9594,N_9911);
nor U10268 (N_10268,N_9876,N_9613);
and U10269 (N_10269,N_9839,N_9545);
nand U10270 (N_10270,N_9728,N_9714);
nor U10271 (N_10271,N_9615,N_9773);
or U10272 (N_10272,N_9863,N_9809);
nand U10273 (N_10273,N_9947,N_9832);
nand U10274 (N_10274,N_9629,N_9639);
xor U10275 (N_10275,N_9746,N_9629);
or U10276 (N_10276,N_9706,N_9920);
and U10277 (N_10277,N_9875,N_9613);
and U10278 (N_10278,N_9960,N_9786);
xor U10279 (N_10279,N_9556,N_9780);
nand U10280 (N_10280,N_9697,N_9652);
nand U10281 (N_10281,N_9951,N_9806);
xor U10282 (N_10282,N_9657,N_9696);
nand U10283 (N_10283,N_9597,N_9932);
nand U10284 (N_10284,N_9958,N_9869);
nand U10285 (N_10285,N_9561,N_9594);
nor U10286 (N_10286,N_9904,N_9945);
nand U10287 (N_10287,N_9940,N_9782);
nand U10288 (N_10288,N_9813,N_9852);
nand U10289 (N_10289,N_9896,N_9649);
nand U10290 (N_10290,N_9657,N_9641);
nand U10291 (N_10291,N_9804,N_9868);
xor U10292 (N_10292,N_9644,N_9705);
xor U10293 (N_10293,N_9926,N_9834);
nand U10294 (N_10294,N_9951,N_9618);
and U10295 (N_10295,N_9566,N_9542);
xnor U10296 (N_10296,N_9910,N_9851);
or U10297 (N_10297,N_9742,N_9624);
or U10298 (N_10298,N_9617,N_9689);
nor U10299 (N_10299,N_9768,N_9910);
and U10300 (N_10300,N_9766,N_9823);
nand U10301 (N_10301,N_9844,N_9766);
nor U10302 (N_10302,N_9781,N_9925);
or U10303 (N_10303,N_9794,N_9702);
and U10304 (N_10304,N_9695,N_9544);
xnor U10305 (N_10305,N_9708,N_9539);
and U10306 (N_10306,N_9581,N_9564);
or U10307 (N_10307,N_9585,N_9607);
and U10308 (N_10308,N_9713,N_9635);
or U10309 (N_10309,N_9748,N_9661);
and U10310 (N_10310,N_9760,N_9758);
xor U10311 (N_10311,N_9918,N_9726);
xnor U10312 (N_10312,N_9710,N_9995);
nor U10313 (N_10313,N_9667,N_9784);
or U10314 (N_10314,N_9542,N_9635);
and U10315 (N_10315,N_9624,N_9608);
xnor U10316 (N_10316,N_9704,N_9659);
or U10317 (N_10317,N_9927,N_9727);
or U10318 (N_10318,N_9554,N_9708);
and U10319 (N_10319,N_9514,N_9927);
or U10320 (N_10320,N_9978,N_9725);
or U10321 (N_10321,N_9897,N_9727);
nor U10322 (N_10322,N_9565,N_9777);
or U10323 (N_10323,N_9773,N_9656);
nor U10324 (N_10324,N_9995,N_9527);
xor U10325 (N_10325,N_9996,N_9754);
nand U10326 (N_10326,N_9547,N_9521);
nor U10327 (N_10327,N_9723,N_9725);
xor U10328 (N_10328,N_9500,N_9589);
nor U10329 (N_10329,N_9772,N_9586);
xnor U10330 (N_10330,N_9823,N_9985);
xor U10331 (N_10331,N_9938,N_9902);
nor U10332 (N_10332,N_9518,N_9671);
xor U10333 (N_10333,N_9834,N_9928);
xor U10334 (N_10334,N_9552,N_9960);
nand U10335 (N_10335,N_9866,N_9952);
nand U10336 (N_10336,N_9811,N_9689);
xnor U10337 (N_10337,N_9568,N_9778);
xnor U10338 (N_10338,N_9802,N_9854);
xnor U10339 (N_10339,N_9592,N_9520);
xor U10340 (N_10340,N_9886,N_9803);
nand U10341 (N_10341,N_9802,N_9532);
xor U10342 (N_10342,N_9843,N_9988);
and U10343 (N_10343,N_9514,N_9610);
xor U10344 (N_10344,N_9805,N_9846);
nor U10345 (N_10345,N_9588,N_9550);
or U10346 (N_10346,N_9787,N_9849);
and U10347 (N_10347,N_9793,N_9897);
nor U10348 (N_10348,N_9839,N_9807);
nor U10349 (N_10349,N_9557,N_9906);
nor U10350 (N_10350,N_9637,N_9697);
nand U10351 (N_10351,N_9789,N_9569);
xnor U10352 (N_10352,N_9601,N_9615);
nand U10353 (N_10353,N_9819,N_9662);
xnor U10354 (N_10354,N_9704,N_9835);
xor U10355 (N_10355,N_9974,N_9854);
and U10356 (N_10356,N_9893,N_9993);
or U10357 (N_10357,N_9729,N_9940);
xor U10358 (N_10358,N_9768,N_9751);
xnor U10359 (N_10359,N_9928,N_9683);
nor U10360 (N_10360,N_9988,N_9907);
or U10361 (N_10361,N_9515,N_9763);
or U10362 (N_10362,N_9856,N_9721);
xnor U10363 (N_10363,N_9793,N_9876);
and U10364 (N_10364,N_9880,N_9971);
xnor U10365 (N_10365,N_9810,N_9537);
or U10366 (N_10366,N_9851,N_9557);
or U10367 (N_10367,N_9861,N_9692);
xor U10368 (N_10368,N_9563,N_9707);
or U10369 (N_10369,N_9987,N_9819);
nor U10370 (N_10370,N_9838,N_9818);
or U10371 (N_10371,N_9615,N_9930);
and U10372 (N_10372,N_9603,N_9730);
and U10373 (N_10373,N_9758,N_9583);
and U10374 (N_10374,N_9842,N_9909);
nand U10375 (N_10375,N_9625,N_9631);
and U10376 (N_10376,N_9519,N_9735);
or U10377 (N_10377,N_9724,N_9950);
or U10378 (N_10378,N_9552,N_9676);
xnor U10379 (N_10379,N_9533,N_9660);
or U10380 (N_10380,N_9801,N_9819);
xor U10381 (N_10381,N_9950,N_9761);
and U10382 (N_10382,N_9982,N_9867);
xor U10383 (N_10383,N_9615,N_9763);
nand U10384 (N_10384,N_9954,N_9716);
xnor U10385 (N_10385,N_9687,N_9523);
xor U10386 (N_10386,N_9561,N_9946);
xor U10387 (N_10387,N_9503,N_9711);
xnor U10388 (N_10388,N_9590,N_9777);
and U10389 (N_10389,N_9794,N_9887);
or U10390 (N_10390,N_9997,N_9859);
or U10391 (N_10391,N_9580,N_9618);
or U10392 (N_10392,N_9745,N_9709);
or U10393 (N_10393,N_9575,N_9535);
or U10394 (N_10394,N_9641,N_9929);
and U10395 (N_10395,N_9846,N_9648);
xnor U10396 (N_10396,N_9563,N_9880);
or U10397 (N_10397,N_9730,N_9695);
nand U10398 (N_10398,N_9947,N_9936);
nand U10399 (N_10399,N_9711,N_9846);
nand U10400 (N_10400,N_9866,N_9574);
xor U10401 (N_10401,N_9810,N_9574);
or U10402 (N_10402,N_9847,N_9731);
and U10403 (N_10403,N_9714,N_9811);
or U10404 (N_10404,N_9894,N_9567);
or U10405 (N_10405,N_9799,N_9992);
and U10406 (N_10406,N_9849,N_9563);
nor U10407 (N_10407,N_9551,N_9777);
nor U10408 (N_10408,N_9962,N_9510);
and U10409 (N_10409,N_9927,N_9731);
or U10410 (N_10410,N_9597,N_9765);
nand U10411 (N_10411,N_9595,N_9796);
nor U10412 (N_10412,N_9788,N_9802);
xor U10413 (N_10413,N_9770,N_9874);
nor U10414 (N_10414,N_9770,N_9991);
xor U10415 (N_10415,N_9851,N_9679);
and U10416 (N_10416,N_9882,N_9517);
nand U10417 (N_10417,N_9946,N_9953);
or U10418 (N_10418,N_9722,N_9895);
xor U10419 (N_10419,N_9940,N_9641);
nand U10420 (N_10420,N_9749,N_9958);
nor U10421 (N_10421,N_9754,N_9786);
nor U10422 (N_10422,N_9501,N_9904);
nand U10423 (N_10423,N_9752,N_9680);
or U10424 (N_10424,N_9845,N_9856);
nand U10425 (N_10425,N_9831,N_9725);
and U10426 (N_10426,N_9992,N_9786);
or U10427 (N_10427,N_9969,N_9946);
nand U10428 (N_10428,N_9972,N_9515);
or U10429 (N_10429,N_9883,N_9889);
or U10430 (N_10430,N_9675,N_9725);
xnor U10431 (N_10431,N_9745,N_9513);
nor U10432 (N_10432,N_9908,N_9539);
and U10433 (N_10433,N_9772,N_9743);
nand U10434 (N_10434,N_9978,N_9870);
or U10435 (N_10435,N_9750,N_9586);
or U10436 (N_10436,N_9865,N_9776);
nand U10437 (N_10437,N_9901,N_9894);
nor U10438 (N_10438,N_9858,N_9714);
xnor U10439 (N_10439,N_9570,N_9871);
nor U10440 (N_10440,N_9981,N_9580);
nand U10441 (N_10441,N_9948,N_9743);
or U10442 (N_10442,N_9571,N_9670);
or U10443 (N_10443,N_9932,N_9807);
nor U10444 (N_10444,N_9823,N_9660);
and U10445 (N_10445,N_9947,N_9921);
or U10446 (N_10446,N_9614,N_9656);
or U10447 (N_10447,N_9987,N_9754);
nor U10448 (N_10448,N_9703,N_9930);
nand U10449 (N_10449,N_9827,N_9566);
nor U10450 (N_10450,N_9934,N_9935);
and U10451 (N_10451,N_9867,N_9544);
xor U10452 (N_10452,N_9884,N_9661);
nand U10453 (N_10453,N_9788,N_9943);
and U10454 (N_10454,N_9601,N_9685);
or U10455 (N_10455,N_9573,N_9542);
and U10456 (N_10456,N_9551,N_9639);
nor U10457 (N_10457,N_9717,N_9600);
nand U10458 (N_10458,N_9607,N_9862);
or U10459 (N_10459,N_9912,N_9672);
and U10460 (N_10460,N_9600,N_9803);
xnor U10461 (N_10461,N_9579,N_9933);
nor U10462 (N_10462,N_9934,N_9858);
nand U10463 (N_10463,N_9856,N_9545);
xor U10464 (N_10464,N_9628,N_9781);
and U10465 (N_10465,N_9831,N_9761);
nand U10466 (N_10466,N_9788,N_9882);
xor U10467 (N_10467,N_9656,N_9913);
nor U10468 (N_10468,N_9991,N_9951);
xnor U10469 (N_10469,N_9717,N_9783);
nor U10470 (N_10470,N_9563,N_9548);
xor U10471 (N_10471,N_9670,N_9950);
nand U10472 (N_10472,N_9632,N_9591);
xnor U10473 (N_10473,N_9763,N_9750);
or U10474 (N_10474,N_9635,N_9724);
xnor U10475 (N_10475,N_9595,N_9634);
xor U10476 (N_10476,N_9927,N_9643);
or U10477 (N_10477,N_9754,N_9635);
nand U10478 (N_10478,N_9652,N_9796);
and U10479 (N_10479,N_9619,N_9939);
and U10480 (N_10480,N_9535,N_9914);
nand U10481 (N_10481,N_9700,N_9587);
nand U10482 (N_10482,N_9749,N_9659);
nand U10483 (N_10483,N_9716,N_9934);
and U10484 (N_10484,N_9811,N_9542);
or U10485 (N_10485,N_9630,N_9656);
nand U10486 (N_10486,N_9619,N_9713);
xor U10487 (N_10487,N_9584,N_9795);
xnor U10488 (N_10488,N_9637,N_9532);
nor U10489 (N_10489,N_9934,N_9823);
nor U10490 (N_10490,N_9692,N_9563);
and U10491 (N_10491,N_9883,N_9590);
or U10492 (N_10492,N_9578,N_9834);
xor U10493 (N_10493,N_9793,N_9948);
xnor U10494 (N_10494,N_9756,N_9793);
or U10495 (N_10495,N_9762,N_9776);
nor U10496 (N_10496,N_9972,N_9800);
nor U10497 (N_10497,N_9620,N_9926);
xor U10498 (N_10498,N_9593,N_9509);
nand U10499 (N_10499,N_9939,N_9504);
or U10500 (N_10500,N_10458,N_10017);
xor U10501 (N_10501,N_10446,N_10154);
and U10502 (N_10502,N_10205,N_10224);
nor U10503 (N_10503,N_10064,N_10113);
nand U10504 (N_10504,N_10341,N_10157);
or U10505 (N_10505,N_10015,N_10161);
or U10506 (N_10506,N_10125,N_10063);
xor U10507 (N_10507,N_10068,N_10404);
nor U10508 (N_10508,N_10010,N_10432);
xor U10509 (N_10509,N_10261,N_10189);
nor U10510 (N_10510,N_10320,N_10426);
or U10511 (N_10511,N_10184,N_10008);
and U10512 (N_10512,N_10175,N_10133);
nand U10513 (N_10513,N_10303,N_10114);
nor U10514 (N_10514,N_10111,N_10347);
or U10515 (N_10515,N_10307,N_10499);
nand U10516 (N_10516,N_10109,N_10260);
or U10517 (N_10517,N_10074,N_10086);
or U10518 (N_10518,N_10098,N_10209);
nor U10519 (N_10519,N_10288,N_10372);
nor U10520 (N_10520,N_10156,N_10211);
and U10521 (N_10521,N_10193,N_10252);
nand U10522 (N_10522,N_10453,N_10406);
xor U10523 (N_10523,N_10278,N_10019);
nor U10524 (N_10524,N_10444,N_10066);
xnor U10525 (N_10525,N_10199,N_10387);
nor U10526 (N_10526,N_10435,N_10409);
and U10527 (N_10527,N_10459,N_10182);
nand U10528 (N_10528,N_10322,N_10047);
nand U10529 (N_10529,N_10243,N_10408);
or U10530 (N_10530,N_10096,N_10423);
or U10531 (N_10531,N_10007,N_10198);
and U10532 (N_10532,N_10119,N_10302);
nand U10533 (N_10533,N_10427,N_10152);
nand U10534 (N_10534,N_10353,N_10037);
nor U10535 (N_10535,N_10229,N_10263);
or U10536 (N_10536,N_10178,N_10070);
nand U10537 (N_10537,N_10494,N_10497);
nor U10538 (N_10538,N_10144,N_10221);
xnor U10539 (N_10539,N_10318,N_10496);
nand U10540 (N_10540,N_10428,N_10438);
nor U10541 (N_10541,N_10140,N_10054);
and U10542 (N_10542,N_10386,N_10150);
or U10543 (N_10543,N_10448,N_10466);
or U10544 (N_10544,N_10331,N_10329);
nor U10545 (N_10545,N_10327,N_10418);
nand U10546 (N_10546,N_10227,N_10089);
xor U10547 (N_10547,N_10285,N_10004);
nand U10548 (N_10548,N_10402,N_10490);
nor U10549 (N_10549,N_10169,N_10363);
nor U10550 (N_10550,N_10286,N_10391);
and U10551 (N_10551,N_10042,N_10348);
xor U10552 (N_10552,N_10056,N_10094);
nand U10553 (N_10553,N_10388,N_10158);
or U10554 (N_10554,N_10162,N_10251);
or U10555 (N_10555,N_10276,N_10396);
nor U10556 (N_10556,N_10220,N_10166);
and U10557 (N_10557,N_10240,N_10367);
nand U10558 (N_10558,N_10151,N_10005);
nor U10559 (N_10559,N_10413,N_10139);
or U10560 (N_10560,N_10312,N_10003);
nor U10561 (N_10561,N_10434,N_10325);
or U10562 (N_10562,N_10065,N_10044);
xor U10563 (N_10563,N_10346,N_10023);
nor U10564 (N_10564,N_10180,N_10040);
or U10565 (N_10565,N_10101,N_10362);
or U10566 (N_10566,N_10217,N_10360);
nor U10567 (N_10567,N_10465,N_10234);
xnor U10568 (N_10568,N_10480,N_10002);
or U10569 (N_10569,N_10077,N_10293);
and U10570 (N_10570,N_10081,N_10097);
or U10571 (N_10571,N_10401,N_10447);
nand U10572 (N_10572,N_10128,N_10377);
and U10573 (N_10573,N_10174,N_10210);
nor U10574 (N_10574,N_10394,N_10087);
nand U10575 (N_10575,N_10366,N_10476);
or U10576 (N_10576,N_10439,N_10279);
nor U10577 (N_10577,N_10395,N_10107);
nor U10578 (N_10578,N_10046,N_10200);
and U10579 (N_10579,N_10488,N_10265);
nand U10580 (N_10580,N_10084,N_10300);
nor U10581 (N_10581,N_10324,N_10283);
nand U10582 (N_10582,N_10163,N_10254);
and U10583 (N_10583,N_10354,N_10148);
nor U10584 (N_10584,N_10121,N_10131);
xor U10585 (N_10585,N_10208,N_10333);
xor U10586 (N_10586,N_10268,N_10299);
and U10587 (N_10587,N_10412,N_10138);
nor U10588 (N_10588,N_10455,N_10379);
and U10589 (N_10589,N_10027,N_10323);
xnor U10590 (N_10590,N_10335,N_10328);
nor U10591 (N_10591,N_10464,N_10429);
nand U10592 (N_10592,N_10264,N_10168);
nor U10593 (N_10593,N_10030,N_10203);
and U10594 (N_10594,N_10470,N_10126);
or U10595 (N_10595,N_10011,N_10226);
nand U10596 (N_10596,N_10306,N_10117);
and U10597 (N_10597,N_10053,N_10454);
nor U10598 (N_10598,N_10246,N_10146);
or U10599 (N_10599,N_10034,N_10228);
xor U10600 (N_10600,N_10233,N_10076);
nor U10601 (N_10601,N_10475,N_10356);
or U10602 (N_10602,N_10093,N_10219);
nand U10603 (N_10603,N_10308,N_10222);
or U10604 (N_10604,N_10104,N_10242);
xor U10605 (N_10605,N_10415,N_10393);
xor U10606 (N_10606,N_10177,N_10132);
and U10607 (N_10607,N_10225,N_10407);
xnor U10608 (N_10608,N_10153,N_10183);
nor U10609 (N_10609,N_10295,N_10461);
nor U10610 (N_10610,N_10258,N_10284);
xor U10611 (N_10611,N_10361,N_10062);
nand U10612 (N_10612,N_10437,N_10296);
nor U10613 (N_10613,N_10389,N_10436);
nand U10614 (N_10614,N_10274,N_10051);
and U10615 (N_10615,N_10164,N_10223);
and U10616 (N_10616,N_10399,N_10337);
xnor U10617 (N_10617,N_10194,N_10115);
nor U10618 (N_10618,N_10055,N_10099);
or U10619 (N_10619,N_10120,N_10247);
or U10620 (N_10620,N_10108,N_10266);
nand U10621 (N_10621,N_10321,N_10127);
or U10622 (N_10622,N_10403,N_10025);
and U10623 (N_10623,N_10309,N_10106);
nand U10624 (N_10624,N_10368,N_10456);
xnor U10625 (N_10625,N_10486,N_10185);
nand U10626 (N_10626,N_10035,N_10257);
nor U10627 (N_10627,N_10050,N_10316);
nor U10628 (N_10628,N_10376,N_10018);
nand U10629 (N_10629,N_10204,N_10147);
and U10630 (N_10630,N_10419,N_10020);
or U10631 (N_10631,N_10390,N_10124);
and U10632 (N_10632,N_10269,N_10213);
nand U10633 (N_10633,N_10191,N_10349);
xor U10634 (N_10634,N_10304,N_10024);
xnor U10635 (N_10635,N_10014,N_10090);
or U10636 (N_10636,N_10463,N_10487);
nor U10637 (N_10637,N_10267,N_10083);
and U10638 (N_10638,N_10473,N_10355);
xor U10639 (N_10639,N_10069,N_10375);
and U10640 (N_10640,N_10181,N_10317);
or U10641 (N_10641,N_10481,N_10425);
and U10642 (N_10642,N_10197,N_10173);
xor U10643 (N_10643,N_10398,N_10039);
nand U10644 (N_10644,N_10080,N_10149);
and U10645 (N_10645,N_10489,N_10414);
and U10646 (N_10646,N_10000,N_10075);
or U10647 (N_10647,N_10236,N_10255);
nor U10648 (N_10648,N_10102,N_10031);
xnor U10649 (N_10649,N_10339,N_10291);
nor U10650 (N_10650,N_10172,N_10452);
or U10651 (N_10651,N_10289,N_10440);
nor U10652 (N_10652,N_10041,N_10049);
nor U10653 (N_10653,N_10078,N_10091);
nand U10654 (N_10654,N_10445,N_10142);
xor U10655 (N_10655,N_10462,N_10332);
or U10656 (N_10656,N_10416,N_10105);
xor U10657 (N_10657,N_10275,N_10116);
nor U10658 (N_10658,N_10103,N_10411);
xnor U10659 (N_10659,N_10192,N_10281);
or U10660 (N_10660,N_10253,N_10060);
nand U10661 (N_10661,N_10092,N_10052);
and U10662 (N_10662,N_10380,N_10239);
nand U10663 (N_10663,N_10430,N_10190);
nand U10664 (N_10664,N_10201,N_10422);
nand U10665 (N_10665,N_10118,N_10314);
nor U10666 (N_10666,N_10443,N_10067);
or U10667 (N_10667,N_10145,N_10186);
xor U10668 (N_10668,N_10134,N_10262);
and U10669 (N_10669,N_10212,N_10484);
nor U10670 (N_10670,N_10248,N_10400);
or U10671 (N_10671,N_10352,N_10342);
nand U10672 (N_10672,N_10215,N_10058);
xor U10673 (N_10673,N_10441,N_10495);
and U10674 (N_10674,N_10359,N_10259);
nor U10675 (N_10675,N_10238,N_10249);
or U10676 (N_10676,N_10073,N_10218);
or U10677 (N_10677,N_10424,N_10207);
and U10678 (N_10678,N_10311,N_10371);
or U10679 (N_10679,N_10457,N_10338);
xor U10680 (N_10680,N_10326,N_10112);
nor U10681 (N_10681,N_10038,N_10351);
nand U10682 (N_10682,N_10137,N_10171);
and U10683 (N_10683,N_10310,N_10498);
xor U10684 (N_10684,N_10319,N_10477);
xor U10685 (N_10685,N_10280,N_10165);
or U10686 (N_10686,N_10032,N_10417);
nor U10687 (N_10687,N_10315,N_10088);
xor U10688 (N_10688,N_10029,N_10384);
nor U10689 (N_10689,N_10292,N_10467);
nand U10690 (N_10690,N_10045,N_10167);
and U10691 (N_10691,N_10057,N_10022);
nand U10692 (N_10692,N_10350,N_10340);
and U10693 (N_10693,N_10021,N_10196);
xor U10694 (N_10694,N_10043,N_10485);
xnor U10695 (N_10695,N_10382,N_10287);
xor U10696 (N_10696,N_10176,N_10273);
xnor U10697 (N_10697,N_10282,N_10016);
nor U10698 (N_10698,N_10373,N_10442);
or U10699 (N_10699,N_10392,N_10358);
nor U10700 (N_10700,N_10061,N_10334);
nand U10701 (N_10701,N_10474,N_10237);
and U10702 (N_10702,N_10012,N_10471);
and U10703 (N_10703,N_10122,N_10059);
nor U10704 (N_10704,N_10294,N_10241);
nor U10705 (N_10705,N_10006,N_10001);
or U10706 (N_10706,N_10250,N_10235);
or U10707 (N_10707,N_10072,N_10179);
nor U10708 (N_10708,N_10385,N_10472);
nand U10709 (N_10709,N_10344,N_10313);
or U10710 (N_10710,N_10378,N_10491);
nor U10711 (N_10711,N_10397,N_10216);
and U10712 (N_10712,N_10336,N_10136);
nor U10713 (N_10713,N_10195,N_10188);
nor U10714 (N_10714,N_10297,N_10206);
nand U10715 (N_10715,N_10245,N_10330);
xor U10716 (N_10716,N_10469,N_10364);
nor U10717 (N_10717,N_10129,N_10013);
nor U10718 (N_10718,N_10187,N_10256);
xor U10719 (N_10719,N_10231,N_10110);
nor U10720 (N_10720,N_10232,N_10160);
xnor U10721 (N_10721,N_10482,N_10468);
xnor U10722 (N_10722,N_10483,N_10033);
nor U10723 (N_10723,N_10270,N_10381);
nor U10724 (N_10724,N_10345,N_10343);
nor U10725 (N_10725,N_10449,N_10451);
nand U10726 (N_10726,N_10460,N_10421);
or U10727 (N_10727,N_10405,N_10431);
or U10728 (N_10728,N_10085,N_10410);
nand U10729 (N_10729,N_10028,N_10143);
or U10730 (N_10730,N_10170,N_10493);
nand U10731 (N_10731,N_10370,N_10135);
nor U10732 (N_10732,N_10082,N_10492);
nor U10733 (N_10733,N_10095,N_10433);
xor U10734 (N_10734,N_10071,N_10079);
nor U10735 (N_10735,N_10420,N_10123);
and U10736 (N_10736,N_10383,N_10026);
or U10737 (N_10737,N_10277,N_10305);
and U10738 (N_10738,N_10450,N_10272);
and U10739 (N_10739,N_10298,N_10290);
xnor U10740 (N_10740,N_10244,N_10369);
nand U10741 (N_10741,N_10230,N_10479);
or U10742 (N_10742,N_10100,N_10141);
and U10743 (N_10743,N_10357,N_10202);
nand U10744 (N_10744,N_10130,N_10036);
xnor U10745 (N_10745,N_10214,N_10478);
xnor U10746 (N_10746,N_10271,N_10365);
or U10747 (N_10747,N_10374,N_10301);
xor U10748 (N_10748,N_10155,N_10048);
or U10749 (N_10749,N_10009,N_10159);
and U10750 (N_10750,N_10196,N_10284);
xnor U10751 (N_10751,N_10435,N_10441);
and U10752 (N_10752,N_10200,N_10073);
and U10753 (N_10753,N_10084,N_10302);
or U10754 (N_10754,N_10143,N_10381);
xor U10755 (N_10755,N_10041,N_10117);
or U10756 (N_10756,N_10468,N_10103);
or U10757 (N_10757,N_10440,N_10111);
or U10758 (N_10758,N_10183,N_10456);
xor U10759 (N_10759,N_10405,N_10213);
and U10760 (N_10760,N_10063,N_10225);
or U10761 (N_10761,N_10020,N_10150);
nor U10762 (N_10762,N_10381,N_10223);
or U10763 (N_10763,N_10441,N_10461);
and U10764 (N_10764,N_10039,N_10434);
or U10765 (N_10765,N_10441,N_10267);
or U10766 (N_10766,N_10487,N_10358);
nor U10767 (N_10767,N_10230,N_10445);
or U10768 (N_10768,N_10278,N_10494);
nand U10769 (N_10769,N_10188,N_10435);
xor U10770 (N_10770,N_10368,N_10060);
or U10771 (N_10771,N_10437,N_10278);
xor U10772 (N_10772,N_10152,N_10181);
nor U10773 (N_10773,N_10441,N_10490);
nand U10774 (N_10774,N_10426,N_10078);
or U10775 (N_10775,N_10383,N_10438);
xor U10776 (N_10776,N_10274,N_10297);
nand U10777 (N_10777,N_10234,N_10257);
or U10778 (N_10778,N_10340,N_10435);
and U10779 (N_10779,N_10070,N_10358);
nor U10780 (N_10780,N_10136,N_10265);
and U10781 (N_10781,N_10357,N_10155);
xnor U10782 (N_10782,N_10359,N_10120);
nand U10783 (N_10783,N_10102,N_10302);
and U10784 (N_10784,N_10279,N_10057);
or U10785 (N_10785,N_10493,N_10009);
xnor U10786 (N_10786,N_10413,N_10378);
or U10787 (N_10787,N_10447,N_10130);
nor U10788 (N_10788,N_10004,N_10228);
or U10789 (N_10789,N_10374,N_10368);
xnor U10790 (N_10790,N_10240,N_10248);
and U10791 (N_10791,N_10190,N_10468);
xor U10792 (N_10792,N_10099,N_10470);
xor U10793 (N_10793,N_10478,N_10439);
nor U10794 (N_10794,N_10324,N_10401);
nand U10795 (N_10795,N_10282,N_10356);
nor U10796 (N_10796,N_10139,N_10110);
xor U10797 (N_10797,N_10232,N_10380);
or U10798 (N_10798,N_10440,N_10145);
nor U10799 (N_10799,N_10242,N_10298);
and U10800 (N_10800,N_10260,N_10059);
or U10801 (N_10801,N_10421,N_10330);
or U10802 (N_10802,N_10250,N_10371);
xnor U10803 (N_10803,N_10368,N_10457);
nand U10804 (N_10804,N_10121,N_10224);
nor U10805 (N_10805,N_10316,N_10229);
or U10806 (N_10806,N_10480,N_10359);
and U10807 (N_10807,N_10310,N_10228);
and U10808 (N_10808,N_10060,N_10043);
and U10809 (N_10809,N_10167,N_10226);
xor U10810 (N_10810,N_10466,N_10371);
xor U10811 (N_10811,N_10484,N_10036);
and U10812 (N_10812,N_10454,N_10305);
nor U10813 (N_10813,N_10471,N_10286);
or U10814 (N_10814,N_10491,N_10000);
and U10815 (N_10815,N_10319,N_10287);
xnor U10816 (N_10816,N_10401,N_10167);
nor U10817 (N_10817,N_10369,N_10060);
xor U10818 (N_10818,N_10400,N_10217);
nor U10819 (N_10819,N_10009,N_10070);
or U10820 (N_10820,N_10164,N_10371);
and U10821 (N_10821,N_10088,N_10435);
nand U10822 (N_10822,N_10448,N_10391);
xor U10823 (N_10823,N_10250,N_10271);
xnor U10824 (N_10824,N_10325,N_10350);
nor U10825 (N_10825,N_10214,N_10332);
or U10826 (N_10826,N_10488,N_10330);
nor U10827 (N_10827,N_10442,N_10035);
nor U10828 (N_10828,N_10109,N_10176);
nor U10829 (N_10829,N_10297,N_10360);
nand U10830 (N_10830,N_10049,N_10479);
or U10831 (N_10831,N_10046,N_10339);
or U10832 (N_10832,N_10266,N_10321);
or U10833 (N_10833,N_10498,N_10321);
and U10834 (N_10834,N_10230,N_10240);
nand U10835 (N_10835,N_10447,N_10442);
and U10836 (N_10836,N_10386,N_10087);
and U10837 (N_10837,N_10483,N_10435);
xor U10838 (N_10838,N_10117,N_10146);
or U10839 (N_10839,N_10111,N_10344);
nor U10840 (N_10840,N_10342,N_10493);
nand U10841 (N_10841,N_10290,N_10180);
xnor U10842 (N_10842,N_10371,N_10268);
nand U10843 (N_10843,N_10109,N_10302);
xor U10844 (N_10844,N_10390,N_10336);
nor U10845 (N_10845,N_10376,N_10061);
nand U10846 (N_10846,N_10250,N_10050);
and U10847 (N_10847,N_10438,N_10455);
nand U10848 (N_10848,N_10128,N_10152);
nor U10849 (N_10849,N_10131,N_10265);
nor U10850 (N_10850,N_10114,N_10402);
nor U10851 (N_10851,N_10006,N_10305);
and U10852 (N_10852,N_10196,N_10163);
and U10853 (N_10853,N_10075,N_10260);
xor U10854 (N_10854,N_10461,N_10180);
or U10855 (N_10855,N_10390,N_10405);
nand U10856 (N_10856,N_10446,N_10082);
and U10857 (N_10857,N_10262,N_10355);
and U10858 (N_10858,N_10418,N_10498);
and U10859 (N_10859,N_10213,N_10072);
and U10860 (N_10860,N_10248,N_10370);
and U10861 (N_10861,N_10419,N_10261);
and U10862 (N_10862,N_10098,N_10127);
or U10863 (N_10863,N_10414,N_10264);
or U10864 (N_10864,N_10378,N_10047);
xor U10865 (N_10865,N_10375,N_10450);
or U10866 (N_10866,N_10108,N_10279);
or U10867 (N_10867,N_10267,N_10338);
or U10868 (N_10868,N_10440,N_10238);
xnor U10869 (N_10869,N_10320,N_10309);
xor U10870 (N_10870,N_10033,N_10100);
and U10871 (N_10871,N_10464,N_10218);
and U10872 (N_10872,N_10429,N_10295);
nor U10873 (N_10873,N_10022,N_10239);
nor U10874 (N_10874,N_10359,N_10105);
nor U10875 (N_10875,N_10276,N_10035);
nor U10876 (N_10876,N_10472,N_10254);
nor U10877 (N_10877,N_10046,N_10080);
and U10878 (N_10878,N_10342,N_10240);
and U10879 (N_10879,N_10148,N_10414);
xor U10880 (N_10880,N_10449,N_10198);
and U10881 (N_10881,N_10317,N_10149);
or U10882 (N_10882,N_10244,N_10454);
xor U10883 (N_10883,N_10416,N_10060);
nand U10884 (N_10884,N_10492,N_10445);
nor U10885 (N_10885,N_10210,N_10128);
or U10886 (N_10886,N_10449,N_10371);
or U10887 (N_10887,N_10317,N_10202);
nor U10888 (N_10888,N_10160,N_10379);
nand U10889 (N_10889,N_10361,N_10334);
or U10890 (N_10890,N_10071,N_10360);
and U10891 (N_10891,N_10177,N_10188);
or U10892 (N_10892,N_10039,N_10239);
nand U10893 (N_10893,N_10177,N_10113);
xor U10894 (N_10894,N_10218,N_10135);
or U10895 (N_10895,N_10498,N_10499);
or U10896 (N_10896,N_10069,N_10394);
or U10897 (N_10897,N_10353,N_10063);
xnor U10898 (N_10898,N_10076,N_10203);
nand U10899 (N_10899,N_10049,N_10151);
or U10900 (N_10900,N_10027,N_10130);
xnor U10901 (N_10901,N_10287,N_10102);
and U10902 (N_10902,N_10378,N_10109);
nand U10903 (N_10903,N_10310,N_10366);
or U10904 (N_10904,N_10454,N_10282);
nand U10905 (N_10905,N_10264,N_10142);
and U10906 (N_10906,N_10393,N_10146);
nand U10907 (N_10907,N_10253,N_10330);
nor U10908 (N_10908,N_10284,N_10420);
nand U10909 (N_10909,N_10367,N_10133);
or U10910 (N_10910,N_10074,N_10072);
xnor U10911 (N_10911,N_10276,N_10479);
xnor U10912 (N_10912,N_10252,N_10311);
nor U10913 (N_10913,N_10183,N_10281);
and U10914 (N_10914,N_10261,N_10011);
nand U10915 (N_10915,N_10190,N_10061);
or U10916 (N_10916,N_10307,N_10206);
nand U10917 (N_10917,N_10045,N_10220);
nor U10918 (N_10918,N_10439,N_10408);
or U10919 (N_10919,N_10227,N_10213);
nor U10920 (N_10920,N_10333,N_10458);
or U10921 (N_10921,N_10496,N_10268);
or U10922 (N_10922,N_10424,N_10053);
nor U10923 (N_10923,N_10202,N_10153);
xor U10924 (N_10924,N_10084,N_10092);
xor U10925 (N_10925,N_10151,N_10122);
nand U10926 (N_10926,N_10302,N_10085);
xor U10927 (N_10927,N_10014,N_10224);
and U10928 (N_10928,N_10086,N_10078);
or U10929 (N_10929,N_10188,N_10259);
or U10930 (N_10930,N_10291,N_10011);
or U10931 (N_10931,N_10071,N_10440);
and U10932 (N_10932,N_10101,N_10298);
and U10933 (N_10933,N_10195,N_10149);
nand U10934 (N_10934,N_10285,N_10021);
nor U10935 (N_10935,N_10428,N_10142);
or U10936 (N_10936,N_10016,N_10135);
xnor U10937 (N_10937,N_10264,N_10090);
nor U10938 (N_10938,N_10298,N_10373);
nor U10939 (N_10939,N_10037,N_10053);
and U10940 (N_10940,N_10462,N_10146);
or U10941 (N_10941,N_10196,N_10126);
or U10942 (N_10942,N_10174,N_10082);
xor U10943 (N_10943,N_10471,N_10494);
nand U10944 (N_10944,N_10260,N_10414);
or U10945 (N_10945,N_10139,N_10085);
nand U10946 (N_10946,N_10279,N_10393);
and U10947 (N_10947,N_10129,N_10158);
or U10948 (N_10948,N_10240,N_10181);
nand U10949 (N_10949,N_10396,N_10108);
or U10950 (N_10950,N_10268,N_10323);
nand U10951 (N_10951,N_10076,N_10364);
xnor U10952 (N_10952,N_10187,N_10054);
or U10953 (N_10953,N_10047,N_10383);
xor U10954 (N_10954,N_10108,N_10009);
and U10955 (N_10955,N_10313,N_10440);
xnor U10956 (N_10956,N_10333,N_10177);
nand U10957 (N_10957,N_10117,N_10403);
xnor U10958 (N_10958,N_10327,N_10325);
xnor U10959 (N_10959,N_10494,N_10309);
xor U10960 (N_10960,N_10197,N_10269);
xor U10961 (N_10961,N_10457,N_10104);
nor U10962 (N_10962,N_10481,N_10391);
nand U10963 (N_10963,N_10306,N_10018);
nor U10964 (N_10964,N_10434,N_10427);
xnor U10965 (N_10965,N_10046,N_10315);
nor U10966 (N_10966,N_10306,N_10083);
nor U10967 (N_10967,N_10173,N_10300);
nor U10968 (N_10968,N_10060,N_10127);
nand U10969 (N_10969,N_10013,N_10170);
xnor U10970 (N_10970,N_10306,N_10484);
nor U10971 (N_10971,N_10401,N_10465);
nand U10972 (N_10972,N_10320,N_10241);
xnor U10973 (N_10973,N_10311,N_10147);
nand U10974 (N_10974,N_10391,N_10465);
nand U10975 (N_10975,N_10414,N_10436);
nand U10976 (N_10976,N_10327,N_10165);
or U10977 (N_10977,N_10046,N_10427);
or U10978 (N_10978,N_10206,N_10291);
xor U10979 (N_10979,N_10486,N_10217);
or U10980 (N_10980,N_10449,N_10403);
and U10981 (N_10981,N_10018,N_10285);
and U10982 (N_10982,N_10014,N_10255);
and U10983 (N_10983,N_10479,N_10282);
and U10984 (N_10984,N_10176,N_10388);
nand U10985 (N_10985,N_10433,N_10382);
xor U10986 (N_10986,N_10289,N_10118);
xnor U10987 (N_10987,N_10130,N_10283);
nor U10988 (N_10988,N_10318,N_10413);
and U10989 (N_10989,N_10365,N_10239);
nand U10990 (N_10990,N_10189,N_10365);
or U10991 (N_10991,N_10295,N_10178);
xnor U10992 (N_10992,N_10407,N_10469);
and U10993 (N_10993,N_10482,N_10061);
nor U10994 (N_10994,N_10093,N_10159);
or U10995 (N_10995,N_10390,N_10333);
nor U10996 (N_10996,N_10113,N_10098);
or U10997 (N_10997,N_10047,N_10493);
and U10998 (N_10998,N_10130,N_10332);
and U10999 (N_10999,N_10260,N_10484);
nor U11000 (N_11000,N_10585,N_10507);
nand U11001 (N_11001,N_10868,N_10911);
nor U11002 (N_11002,N_10995,N_10598);
nor U11003 (N_11003,N_10631,N_10518);
and U11004 (N_11004,N_10630,N_10915);
or U11005 (N_11005,N_10551,N_10790);
nand U11006 (N_11006,N_10566,N_10816);
and U11007 (N_11007,N_10575,N_10837);
nand U11008 (N_11008,N_10657,N_10909);
nand U11009 (N_11009,N_10871,N_10502);
or U11010 (N_11010,N_10870,N_10989);
nor U11011 (N_11011,N_10991,N_10833);
xnor U11012 (N_11012,N_10515,N_10877);
nand U11013 (N_11013,N_10970,N_10579);
and U11014 (N_11014,N_10623,N_10887);
xor U11015 (N_11015,N_10764,N_10514);
nor U11016 (N_11016,N_10792,N_10547);
nand U11017 (N_11017,N_10893,N_10596);
nor U11018 (N_11018,N_10685,N_10673);
xnor U11019 (N_11019,N_10729,N_10677);
nand U11020 (N_11020,N_10895,N_10606);
and U11021 (N_11021,N_10883,N_10982);
xnor U11022 (N_11022,N_10704,N_10741);
xor U11023 (N_11023,N_10640,N_10912);
and U11024 (N_11024,N_10758,N_10536);
and U11025 (N_11025,N_10849,N_10666);
nand U11026 (N_11026,N_10735,N_10933);
nand U11027 (N_11027,N_10805,N_10519);
and U11028 (N_11028,N_10956,N_10917);
nand U11029 (N_11029,N_10609,N_10726);
xnor U11030 (N_11030,N_10719,N_10638);
nand U11031 (N_11031,N_10787,N_10753);
or U11032 (N_11032,N_10768,N_10910);
nand U11033 (N_11033,N_10796,N_10978);
nand U11034 (N_11034,N_10880,N_10847);
and U11035 (N_11035,N_10797,N_10635);
or U11036 (N_11036,N_10803,N_10942);
and U11037 (N_11037,N_10992,N_10628);
nand U11038 (N_11038,N_10953,N_10616);
or U11039 (N_11039,N_10571,N_10836);
nand U11040 (N_11040,N_10621,N_10965);
or U11041 (N_11041,N_10608,N_10802);
or U11042 (N_11042,N_10675,N_10810);
nor U11043 (N_11043,N_10588,N_10510);
and U11044 (N_11044,N_10736,N_10822);
nor U11045 (N_11045,N_10959,N_10544);
and U11046 (N_11046,N_10614,N_10972);
and U11047 (N_11047,N_10980,N_10681);
and U11048 (N_11048,N_10777,N_10732);
xnor U11049 (N_11049,N_10878,N_10552);
nor U11050 (N_11050,N_10706,N_10919);
and U11051 (N_11051,N_10698,N_10527);
nand U11052 (N_11052,N_10931,N_10851);
nand U11053 (N_11053,N_10587,N_10595);
or U11054 (N_11054,N_10838,N_10788);
nand U11055 (N_11055,N_10664,N_10639);
xor U11056 (N_11056,N_10715,N_10637);
xnor U11057 (N_11057,N_10538,N_10783);
or U11058 (N_11058,N_10940,N_10650);
nor U11059 (N_11059,N_10711,N_10727);
nor U11060 (N_11060,N_10929,N_10503);
and U11061 (N_11061,N_10636,N_10806);
xor U11062 (N_11062,N_10769,N_10904);
and U11063 (N_11063,N_10899,N_10641);
xor U11064 (N_11064,N_10712,N_10694);
and U11065 (N_11065,N_10688,N_10655);
or U11066 (N_11066,N_10826,N_10857);
or U11067 (N_11067,N_10892,N_10665);
nand U11068 (N_11068,N_10610,N_10505);
or U11069 (N_11069,N_10730,N_10879);
and U11070 (N_11070,N_10924,N_10888);
xor U11071 (N_11071,N_10707,N_10864);
and U11072 (N_11072,N_10844,N_10898);
xor U11073 (N_11073,N_10512,N_10572);
or U11074 (N_11074,N_10850,N_10508);
nand U11075 (N_11075,N_10613,N_10958);
or U11076 (N_11076,N_10778,N_10570);
nand U11077 (N_11077,N_10807,N_10580);
xnor U11078 (N_11078,N_10798,N_10656);
xor U11079 (N_11079,N_10697,N_10761);
nand U11080 (N_11080,N_10763,N_10964);
xnor U11081 (N_11081,N_10927,N_10687);
or U11082 (N_11082,N_10713,N_10533);
nor U11083 (N_11083,N_10988,N_10553);
nor U11084 (N_11084,N_10969,N_10828);
and U11085 (N_11085,N_10817,N_10537);
xor U11086 (N_11086,N_10979,N_10583);
nor U11087 (N_11087,N_10835,N_10996);
xnor U11088 (N_11088,N_10771,N_10819);
nor U11089 (N_11089,N_10737,N_10555);
xor U11090 (N_11090,N_10659,N_10949);
and U11091 (N_11091,N_10963,N_10997);
or U11092 (N_11092,N_10954,N_10984);
nor U11093 (N_11093,N_10701,N_10950);
nor U11094 (N_11094,N_10756,N_10582);
nand U11095 (N_11095,N_10926,N_10842);
or U11096 (N_11096,N_10865,N_10618);
nor U11097 (N_11097,N_10928,N_10821);
nand U11098 (N_11098,N_10914,N_10918);
nor U11099 (N_11099,N_10534,N_10661);
nand U11100 (N_11100,N_10724,N_10863);
or U11101 (N_11101,N_10674,N_10922);
xor U11102 (N_11102,N_10722,N_10604);
nand U11103 (N_11103,N_10751,N_10607);
or U11104 (N_11104,N_10632,N_10633);
or U11105 (N_11105,N_10759,N_10750);
nand U11106 (N_11106,N_10591,N_10528);
xnor U11107 (N_11107,N_10622,N_10731);
and U11108 (N_11108,N_10511,N_10944);
or U11109 (N_11109,N_10859,N_10841);
nand U11110 (N_11110,N_10634,N_10748);
nor U11111 (N_11111,N_10660,N_10522);
nand U11112 (N_11112,N_10740,N_10908);
nand U11113 (N_11113,N_10627,N_10775);
and U11114 (N_11114,N_10939,N_10973);
xor U11115 (N_11115,N_10517,N_10629);
nand U11116 (N_11116,N_10906,N_10831);
nand U11117 (N_11117,N_10742,N_10714);
nor U11118 (N_11118,N_10611,N_10794);
or U11119 (N_11119,N_10907,N_10998);
nor U11120 (N_11120,N_10540,N_10746);
nand U11121 (N_11121,N_10814,N_10577);
xnor U11122 (N_11122,N_10823,N_10804);
nor U11123 (N_11123,N_10653,N_10846);
nand U11124 (N_11124,N_10882,N_10854);
nor U11125 (N_11125,N_10619,N_10860);
and U11126 (N_11126,N_10968,N_10589);
xor U11127 (N_11127,N_10977,N_10872);
or U11128 (N_11128,N_10824,N_10564);
nand U11129 (N_11129,N_10671,N_10717);
or U11130 (N_11130,N_10576,N_10994);
or U11131 (N_11131,N_10529,N_10773);
nand U11132 (N_11132,N_10999,N_10643);
nor U11133 (N_11133,N_10644,N_10866);
and U11134 (N_11134,N_10962,N_10689);
and U11135 (N_11135,N_10952,N_10738);
xor U11136 (N_11136,N_10662,N_10772);
and U11137 (N_11137,N_10853,N_10745);
xnor U11138 (N_11138,N_10897,N_10592);
xnor U11139 (N_11139,N_10957,N_10829);
nand U11140 (N_11140,N_10974,N_10578);
nand U11141 (N_11141,N_10624,N_10967);
and U11142 (N_11142,N_10695,N_10620);
nor U11143 (N_11143,N_10523,N_10985);
or U11144 (N_11144,N_10839,N_10549);
nand U11145 (N_11145,N_10946,N_10840);
nand U11146 (N_11146,N_10784,N_10721);
nand U11147 (N_11147,N_10586,N_10902);
nand U11148 (N_11148,N_10646,N_10961);
and U11149 (N_11149,N_10943,N_10718);
xor U11150 (N_11150,N_10976,N_10651);
nand U11151 (N_11151,N_10541,N_10599);
and U11152 (N_11152,N_10925,N_10543);
or U11153 (N_11153,N_10526,N_10574);
nor U11154 (N_11154,N_10852,N_10504);
nand U11155 (N_11155,N_10684,N_10891);
nand U11156 (N_11156,N_10765,N_10593);
nand U11157 (N_11157,N_10557,N_10856);
or U11158 (N_11158,N_10825,N_10669);
nand U11159 (N_11159,N_10743,N_10561);
nand U11160 (N_11160,N_10501,N_10710);
xor U11161 (N_11161,N_10916,N_10749);
and U11162 (N_11162,N_10789,N_10884);
or U11163 (N_11163,N_10560,N_10867);
xor U11164 (N_11164,N_10975,N_10932);
nor U11165 (N_11165,N_10696,N_10920);
and U11166 (N_11166,N_10556,N_10680);
nand U11167 (N_11167,N_10542,N_10679);
nand U11168 (N_11168,N_10752,N_10563);
nor U11169 (N_11169,N_10739,N_10625);
and U11170 (N_11170,N_10682,N_10568);
nand U11171 (N_11171,N_10716,N_10600);
nor U11172 (N_11172,N_10937,N_10843);
nand U11173 (N_11173,N_10594,N_10781);
nor U11174 (N_11174,N_10559,N_10550);
nor U11175 (N_11175,N_10938,N_10703);
nand U11176 (N_11176,N_10834,N_10554);
or U11177 (N_11177,N_10776,N_10873);
xnor U11178 (N_11178,N_10709,N_10678);
and U11179 (N_11179,N_10725,N_10830);
or U11180 (N_11180,N_10676,N_10548);
or U11181 (N_11181,N_10855,N_10720);
or U11182 (N_11182,N_10649,N_10723);
xor U11183 (N_11183,N_10692,N_10668);
or U11184 (N_11184,N_10691,N_10734);
or U11185 (N_11185,N_10981,N_10945);
and U11186 (N_11186,N_10690,N_10827);
or U11187 (N_11187,N_10520,N_10516);
xor U11188 (N_11188,N_10584,N_10647);
nand U11189 (N_11189,N_10947,N_10936);
nor U11190 (N_11190,N_10652,N_10894);
nand U11191 (N_11191,N_10800,N_10971);
nor U11192 (N_11192,N_10648,N_10762);
nor U11193 (N_11193,N_10509,N_10889);
nand U11194 (N_11194,N_10558,N_10755);
and U11195 (N_11195,N_10809,N_10539);
nor U11196 (N_11196,N_10785,N_10562);
xor U11197 (N_11197,N_10617,N_10820);
nor U11198 (N_11198,N_10848,N_10881);
xnor U11199 (N_11199,N_10780,N_10869);
nand U11200 (N_11200,N_10966,N_10766);
nand U11201 (N_11201,N_10793,N_10923);
and U11202 (N_11202,N_10808,N_10845);
xnor U11203 (N_11203,N_10874,N_10728);
or U11204 (N_11204,N_10801,N_10513);
nand U11205 (N_11205,N_10811,N_10782);
xnor U11206 (N_11206,N_10642,N_10886);
nor U11207 (N_11207,N_10506,N_10573);
xnor U11208 (N_11208,N_10601,N_10875);
xor U11209 (N_11209,N_10901,N_10525);
xnor U11210 (N_11210,N_10702,N_10597);
or U11211 (N_11211,N_10941,N_10760);
and U11212 (N_11212,N_10672,N_10876);
and U11213 (N_11213,N_10546,N_10983);
nand U11214 (N_11214,N_10757,N_10791);
and U11215 (N_11215,N_10951,N_10531);
nor U11216 (N_11216,N_10900,N_10779);
xor U11217 (N_11217,N_10861,N_10603);
and U11218 (N_11218,N_10708,N_10832);
and U11219 (N_11219,N_10799,N_10885);
nor U11220 (N_11220,N_10569,N_10683);
xnor U11221 (N_11221,N_10921,N_10567);
nand U11222 (N_11222,N_10500,N_10815);
xnor U11223 (N_11223,N_10993,N_10530);
and U11224 (N_11224,N_10663,N_10705);
and U11225 (N_11225,N_10774,N_10654);
nand U11226 (N_11226,N_10948,N_10960);
and U11227 (N_11227,N_10795,N_10686);
xnor U11228 (N_11228,N_10955,N_10896);
or U11229 (N_11229,N_10602,N_10605);
or U11230 (N_11230,N_10565,N_10786);
nand U11231 (N_11231,N_10733,N_10615);
and U11232 (N_11232,N_10770,N_10658);
and U11233 (N_11233,N_10987,N_10754);
or U11234 (N_11234,N_10812,N_10545);
nor U11235 (N_11235,N_10590,N_10890);
nor U11236 (N_11236,N_10818,N_10612);
nand U11237 (N_11237,N_10930,N_10693);
or U11238 (N_11238,N_10699,N_10813);
or U11239 (N_11239,N_10905,N_10581);
or U11240 (N_11240,N_10747,N_10744);
nand U11241 (N_11241,N_10626,N_10935);
nor U11242 (N_11242,N_10990,N_10858);
xor U11243 (N_11243,N_10521,N_10862);
nand U11244 (N_11244,N_10986,N_10524);
xnor U11245 (N_11245,N_10667,N_10700);
and U11246 (N_11246,N_10913,N_10767);
xor U11247 (N_11247,N_10934,N_10645);
and U11248 (N_11248,N_10903,N_10535);
nand U11249 (N_11249,N_10532,N_10670);
xnor U11250 (N_11250,N_10892,N_10980);
nand U11251 (N_11251,N_10812,N_10653);
or U11252 (N_11252,N_10896,N_10718);
and U11253 (N_11253,N_10788,N_10737);
xor U11254 (N_11254,N_10707,N_10947);
and U11255 (N_11255,N_10832,N_10818);
nand U11256 (N_11256,N_10879,N_10977);
nor U11257 (N_11257,N_10870,N_10942);
nor U11258 (N_11258,N_10926,N_10562);
xor U11259 (N_11259,N_10955,N_10694);
or U11260 (N_11260,N_10875,N_10750);
and U11261 (N_11261,N_10958,N_10922);
xnor U11262 (N_11262,N_10882,N_10800);
nor U11263 (N_11263,N_10976,N_10951);
or U11264 (N_11264,N_10514,N_10733);
and U11265 (N_11265,N_10735,N_10715);
and U11266 (N_11266,N_10755,N_10689);
nor U11267 (N_11267,N_10577,N_10797);
xnor U11268 (N_11268,N_10531,N_10533);
xnor U11269 (N_11269,N_10563,N_10876);
xor U11270 (N_11270,N_10506,N_10532);
nand U11271 (N_11271,N_10549,N_10565);
and U11272 (N_11272,N_10579,N_10789);
nand U11273 (N_11273,N_10970,N_10640);
xor U11274 (N_11274,N_10570,N_10920);
and U11275 (N_11275,N_10795,N_10724);
and U11276 (N_11276,N_10582,N_10776);
nor U11277 (N_11277,N_10859,N_10669);
nor U11278 (N_11278,N_10879,N_10856);
or U11279 (N_11279,N_10774,N_10614);
xor U11280 (N_11280,N_10855,N_10750);
nor U11281 (N_11281,N_10910,N_10855);
xnor U11282 (N_11282,N_10902,N_10955);
and U11283 (N_11283,N_10915,N_10905);
or U11284 (N_11284,N_10718,N_10566);
nor U11285 (N_11285,N_10748,N_10584);
nand U11286 (N_11286,N_10749,N_10737);
or U11287 (N_11287,N_10647,N_10654);
xor U11288 (N_11288,N_10851,N_10983);
or U11289 (N_11289,N_10693,N_10880);
nor U11290 (N_11290,N_10698,N_10899);
xor U11291 (N_11291,N_10654,N_10570);
nand U11292 (N_11292,N_10877,N_10681);
and U11293 (N_11293,N_10876,N_10946);
xnor U11294 (N_11294,N_10940,N_10907);
nor U11295 (N_11295,N_10740,N_10800);
and U11296 (N_11296,N_10802,N_10558);
xor U11297 (N_11297,N_10934,N_10821);
nor U11298 (N_11298,N_10572,N_10850);
xor U11299 (N_11299,N_10922,N_10913);
and U11300 (N_11300,N_10708,N_10614);
nand U11301 (N_11301,N_10951,N_10928);
or U11302 (N_11302,N_10821,N_10612);
and U11303 (N_11303,N_10630,N_10961);
and U11304 (N_11304,N_10510,N_10675);
xor U11305 (N_11305,N_10974,N_10626);
and U11306 (N_11306,N_10783,N_10633);
and U11307 (N_11307,N_10602,N_10503);
nor U11308 (N_11308,N_10848,N_10858);
nor U11309 (N_11309,N_10719,N_10848);
nor U11310 (N_11310,N_10989,N_10988);
and U11311 (N_11311,N_10845,N_10744);
nand U11312 (N_11312,N_10717,N_10738);
and U11313 (N_11313,N_10515,N_10806);
nand U11314 (N_11314,N_10509,N_10743);
xor U11315 (N_11315,N_10792,N_10707);
nor U11316 (N_11316,N_10808,N_10636);
xnor U11317 (N_11317,N_10943,N_10808);
and U11318 (N_11318,N_10856,N_10724);
xnor U11319 (N_11319,N_10938,N_10987);
or U11320 (N_11320,N_10806,N_10978);
nor U11321 (N_11321,N_10649,N_10526);
nor U11322 (N_11322,N_10925,N_10545);
nand U11323 (N_11323,N_10711,N_10759);
nor U11324 (N_11324,N_10627,N_10769);
or U11325 (N_11325,N_10580,N_10666);
or U11326 (N_11326,N_10985,N_10865);
nand U11327 (N_11327,N_10875,N_10754);
and U11328 (N_11328,N_10698,N_10940);
nor U11329 (N_11329,N_10512,N_10808);
nand U11330 (N_11330,N_10975,N_10592);
nand U11331 (N_11331,N_10607,N_10933);
xor U11332 (N_11332,N_10728,N_10658);
nand U11333 (N_11333,N_10699,N_10687);
xor U11334 (N_11334,N_10517,N_10667);
xor U11335 (N_11335,N_10519,N_10578);
xnor U11336 (N_11336,N_10847,N_10840);
nor U11337 (N_11337,N_10562,N_10789);
xor U11338 (N_11338,N_10832,N_10625);
nor U11339 (N_11339,N_10883,N_10908);
nand U11340 (N_11340,N_10566,N_10700);
nand U11341 (N_11341,N_10548,N_10807);
nor U11342 (N_11342,N_10906,N_10963);
xor U11343 (N_11343,N_10505,N_10624);
or U11344 (N_11344,N_10578,N_10827);
or U11345 (N_11345,N_10768,N_10926);
and U11346 (N_11346,N_10635,N_10959);
nand U11347 (N_11347,N_10964,N_10539);
nor U11348 (N_11348,N_10788,N_10646);
and U11349 (N_11349,N_10928,N_10721);
xnor U11350 (N_11350,N_10837,N_10630);
and U11351 (N_11351,N_10985,N_10565);
xnor U11352 (N_11352,N_10531,N_10563);
nor U11353 (N_11353,N_10971,N_10827);
xor U11354 (N_11354,N_10551,N_10505);
and U11355 (N_11355,N_10948,N_10585);
nand U11356 (N_11356,N_10663,N_10927);
and U11357 (N_11357,N_10841,N_10637);
and U11358 (N_11358,N_10730,N_10796);
nor U11359 (N_11359,N_10526,N_10591);
nor U11360 (N_11360,N_10519,N_10720);
or U11361 (N_11361,N_10847,N_10610);
nor U11362 (N_11362,N_10945,N_10537);
nand U11363 (N_11363,N_10851,N_10898);
and U11364 (N_11364,N_10995,N_10586);
and U11365 (N_11365,N_10712,N_10709);
xor U11366 (N_11366,N_10892,N_10608);
nand U11367 (N_11367,N_10662,N_10502);
xnor U11368 (N_11368,N_10978,N_10500);
and U11369 (N_11369,N_10867,N_10686);
xnor U11370 (N_11370,N_10651,N_10545);
nand U11371 (N_11371,N_10787,N_10558);
xor U11372 (N_11372,N_10563,N_10969);
nand U11373 (N_11373,N_10802,N_10867);
nor U11374 (N_11374,N_10543,N_10521);
xor U11375 (N_11375,N_10659,N_10970);
nor U11376 (N_11376,N_10839,N_10824);
or U11377 (N_11377,N_10812,N_10728);
nand U11378 (N_11378,N_10526,N_10978);
xor U11379 (N_11379,N_10553,N_10664);
nor U11380 (N_11380,N_10670,N_10511);
nor U11381 (N_11381,N_10832,N_10742);
xnor U11382 (N_11382,N_10897,N_10696);
nor U11383 (N_11383,N_10527,N_10988);
nand U11384 (N_11384,N_10671,N_10846);
nor U11385 (N_11385,N_10831,N_10929);
nand U11386 (N_11386,N_10841,N_10601);
xor U11387 (N_11387,N_10501,N_10885);
xnor U11388 (N_11388,N_10997,N_10967);
nor U11389 (N_11389,N_10634,N_10961);
or U11390 (N_11390,N_10991,N_10625);
nor U11391 (N_11391,N_10552,N_10866);
and U11392 (N_11392,N_10502,N_10818);
nand U11393 (N_11393,N_10827,N_10840);
or U11394 (N_11394,N_10700,N_10784);
xnor U11395 (N_11395,N_10506,N_10812);
xnor U11396 (N_11396,N_10590,N_10842);
and U11397 (N_11397,N_10618,N_10883);
nor U11398 (N_11398,N_10711,N_10995);
nand U11399 (N_11399,N_10676,N_10850);
or U11400 (N_11400,N_10671,N_10513);
nand U11401 (N_11401,N_10874,N_10753);
nand U11402 (N_11402,N_10790,N_10865);
nor U11403 (N_11403,N_10795,N_10534);
xnor U11404 (N_11404,N_10508,N_10794);
nor U11405 (N_11405,N_10634,N_10630);
xnor U11406 (N_11406,N_10652,N_10876);
nand U11407 (N_11407,N_10686,N_10821);
xnor U11408 (N_11408,N_10982,N_10580);
and U11409 (N_11409,N_10505,N_10715);
nor U11410 (N_11410,N_10582,N_10932);
or U11411 (N_11411,N_10888,N_10812);
xnor U11412 (N_11412,N_10611,N_10646);
nor U11413 (N_11413,N_10792,N_10897);
or U11414 (N_11414,N_10823,N_10613);
or U11415 (N_11415,N_10603,N_10599);
nor U11416 (N_11416,N_10672,N_10661);
and U11417 (N_11417,N_10885,N_10551);
or U11418 (N_11418,N_10635,N_10856);
or U11419 (N_11419,N_10659,N_10866);
nand U11420 (N_11420,N_10711,N_10899);
xor U11421 (N_11421,N_10701,N_10980);
nand U11422 (N_11422,N_10570,N_10594);
or U11423 (N_11423,N_10827,N_10950);
and U11424 (N_11424,N_10644,N_10913);
and U11425 (N_11425,N_10877,N_10781);
nand U11426 (N_11426,N_10587,N_10686);
nor U11427 (N_11427,N_10602,N_10615);
and U11428 (N_11428,N_10586,N_10882);
and U11429 (N_11429,N_10813,N_10695);
nor U11430 (N_11430,N_10530,N_10532);
nor U11431 (N_11431,N_10729,N_10746);
or U11432 (N_11432,N_10661,N_10863);
or U11433 (N_11433,N_10660,N_10666);
or U11434 (N_11434,N_10607,N_10685);
nor U11435 (N_11435,N_10951,N_10752);
nand U11436 (N_11436,N_10585,N_10860);
nor U11437 (N_11437,N_10749,N_10897);
nand U11438 (N_11438,N_10667,N_10531);
xor U11439 (N_11439,N_10702,N_10948);
and U11440 (N_11440,N_10976,N_10991);
nand U11441 (N_11441,N_10858,N_10557);
nand U11442 (N_11442,N_10590,N_10917);
nand U11443 (N_11443,N_10807,N_10734);
nor U11444 (N_11444,N_10631,N_10970);
and U11445 (N_11445,N_10580,N_10592);
and U11446 (N_11446,N_10738,N_10546);
nor U11447 (N_11447,N_10608,N_10660);
xnor U11448 (N_11448,N_10983,N_10854);
or U11449 (N_11449,N_10805,N_10611);
nor U11450 (N_11450,N_10940,N_10845);
xor U11451 (N_11451,N_10854,N_10675);
and U11452 (N_11452,N_10891,N_10904);
nand U11453 (N_11453,N_10578,N_10924);
or U11454 (N_11454,N_10863,N_10803);
or U11455 (N_11455,N_10853,N_10986);
nand U11456 (N_11456,N_10912,N_10732);
and U11457 (N_11457,N_10683,N_10913);
or U11458 (N_11458,N_10825,N_10783);
nand U11459 (N_11459,N_10708,N_10767);
nand U11460 (N_11460,N_10724,N_10969);
nor U11461 (N_11461,N_10822,N_10592);
nor U11462 (N_11462,N_10695,N_10539);
xnor U11463 (N_11463,N_10918,N_10817);
or U11464 (N_11464,N_10589,N_10871);
or U11465 (N_11465,N_10994,N_10850);
nor U11466 (N_11466,N_10846,N_10628);
nand U11467 (N_11467,N_10521,N_10660);
nand U11468 (N_11468,N_10744,N_10589);
nor U11469 (N_11469,N_10707,N_10542);
nor U11470 (N_11470,N_10993,N_10691);
and U11471 (N_11471,N_10967,N_10564);
nand U11472 (N_11472,N_10843,N_10564);
xnor U11473 (N_11473,N_10681,N_10814);
nor U11474 (N_11474,N_10767,N_10904);
nor U11475 (N_11475,N_10569,N_10846);
xor U11476 (N_11476,N_10512,N_10520);
xor U11477 (N_11477,N_10924,N_10691);
or U11478 (N_11478,N_10918,N_10602);
or U11479 (N_11479,N_10920,N_10752);
and U11480 (N_11480,N_10881,N_10784);
nor U11481 (N_11481,N_10574,N_10862);
nand U11482 (N_11482,N_10763,N_10800);
or U11483 (N_11483,N_10844,N_10921);
and U11484 (N_11484,N_10898,N_10889);
and U11485 (N_11485,N_10522,N_10623);
xor U11486 (N_11486,N_10590,N_10966);
nor U11487 (N_11487,N_10837,N_10586);
and U11488 (N_11488,N_10809,N_10694);
or U11489 (N_11489,N_10829,N_10824);
nand U11490 (N_11490,N_10762,N_10587);
xnor U11491 (N_11491,N_10575,N_10953);
nor U11492 (N_11492,N_10966,N_10667);
xor U11493 (N_11493,N_10896,N_10553);
xor U11494 (N_11494,N_10886,N_10547);
nor U11495 (N_11495,N_10809,N_10976);
and U11496 (N_11496,N_10774,N_10603);
and U11497 (N_11497,N_10912,N_10735);
and U11498 (N_11498,N_10663,N_10884);
and U11499 (N_11499,N_10576,N_10802);
xnor U11500 (N_11500,N_11192,N_11048);
nand U11501 (N_11501,N_11195,N_11138);
nor U11502 (N_11502,N_11361,N_11108);
or U11503 (N_11503,N_11493,N_11448);
nor U11504 (N_11504,N_11351,N_11237);
xor U11505 (N_11505,N_11114,N_11368);
nand U11506 (N_11506,N_11333,N_11294);
xor U11507 (N_11507,N_11003,N_11184);
and U11508 (N_11508,N_11053,N_11122);
nor U11509 (N_11509,N_11466,N_11317);
xor U11510 (N_11510,N_11331,N_11484);
nand U11511 (N_11511,N_11235,N_11041);
nand U11512 (N_11512,N_11064,N_11253);
nor U11513 (N_11513,N_11251,N_11059);
nand U11514 (N_11514,N_11144,N_11110);
nand U11515 (N_11515,N_11413,N_11220);
xor U11516 (N_11516,N_11371,N_11298);
xnor U11517 (N_11517,N_11244,N_11081);
or U11518 (N_11518,N_11412,N_11206);
nand U11519 (N_11519,N_11450,N_11436);
nand U11520 (N_11520,N_11330,N_11451);
nor U11521 (N_11521,N_11084,N_11377);
or U11522 (N_11522,N_11109,N_11303);
nor U11523 (N_11523,N_11010,N_11124);
and U11524 (N_11524,N_11083,N_11452);
nand U11525 (N_11525,N_11446,N_11071);
xnor U11526 (N_11526,N_11125,N_11270);
nand U11527 (N_11527,N_11167,N_11376);
xnor U11528 (N_11528,N_11218,N_11005);
or U11529 (N_11529,N_11036,N_11057);
xor U11530 (N_11530,N_11315,N_11152);
or U11531 (N_11531,N_11187,N_11364);
xor U11532 (N_11532,N_11362,N_11089);
and U11533 (N_11533,N_11102,N_11032);
nand U11534 (N_11534,N_11086,N_11065);
nand U11535 (N_11535,N_11239,N_11061);
nor U11536 (N_11536,N_11196,N_11389);
xor U11537 (N_11537,N_11111,N_11444);
xor U11538 (N_11538,N_11177,N_11374);
or U11539 (N_11539,N_11367,N_11236);
nor U11540 (N_11540,N_11247,N_11476);
nor U11541 (N_11541,N_11094,N_11211);
nor U11542 (N_11542,N_11008,N_11335);
xnor U11543 (N_11543,N_11068,N_11231);
xor U11544 (N_11544,N_11391,N_11148);
or U11545 (N_11545,N_11019,N_11249);
or U11546 (N_11546,N_11274,N_11272);
nor U11547 (N_11547,N_11171,N_11354);
nand U11548 (N_11548,N_11259,N_11426);
nor U11549 (N_11549,N_11130,N_11035);
or U11550 (N_11550,N_11497,N_11013);
nor U11551 (N_11551,N_11438,N_11105);
nand U11552 (N_11552,N_11355,N_11098);
nor U11553 (N_11553,N_11121,N_11280);
xor U11554 (N_11554,N_11268,N_11226);
and U11555 (N_11555,N_11345,N_11264);
or U11556 (N_11556,N_11284,N_11208);
xor U11557 (N_11557,N_11258,N_11047);
or U11558 (N_11558,N_11100,N_11411);
nand U11559 (N_11559,N_11290,N_11153);
xnor U11560 (N_11560,N_11313,N_11097);
nand U11561 (N_11561,N_11383,N_11396);
xor U11562 (N_11562,N_11063,N_11092);
and U11563 (N_11563,N_11046,N_11205);
nand U11564 (N_11564,N_11457,N_11233);
nand U11565 (N_11565,N_11232,N_11337);
nand U11566 (N_11566,N_11453,N_11357);
xor U11567 (N_11567,N_11437,N_11300);
nand U11568 (N_11568,N_11215,N_11066);
nand U11569 (N_11569,N_11262,N_11372);
and U11570 (N_11570,N_11181,N_11441);
and U11571 (N_11571,N_11217,N_11201);
nor U11572 (N_11572,N_11252,N_11416);
or U11573 (N_11573,N_11439,N_11475);
nor U11574 (N_11574,N_11246,N_11091);
nand U11575 (N_11575,N_11021,N_11319);
or U11576 (N_11576,N_11198,N_11341);
xnor U11577 (N_11577,N_11329,N_11166);
nand U11578 (N_11578,N_11145,N_11267);
nand U11579 (N_11579,N_11460,N_11408);
and U11580 (N_11580,N_11051,N_11347);
or U11581 (N_11581,N_11386,N_11265);
xor U11582 (N_11582,N_11325,N_11228);
xnor U11583 (N_11583,N_11305,N_11082);
and U11584 (N_11584,N_11112,N_11432);
nand U11585 (N_11585,N_11076,N_11096);
nor U11586 (N_11586,N_11207,N_11115);
nor U11587 (N_11587,N_11353,N_11494);
nand U11588 (N_11588,N_11212,N_11404);
and U11589 (N_11589,N_11400,N_11358);
nand U11590 (N_11590,N_11458,N_11238);
nand U11591 (N_11591,N_11414,N_11052);
and U11592 (N_11592,N_11219,N_11402);
and U11593 (N_11593,N_11031,N_11189);
nand U11594 (N_11594,N_11470,N_11486);
or U11595 (N_11595,N_11155,N_11467);
or U11596 (N_11596,N_11296,N_11009);
nor U11597 (N_11597,N_11488,N_11334);
and U11598 (N_11598,N_11487,N_11409);
and U11599 (N_11599,N_11449,N_11140);
or U11600 (N_11600,N_11157,N_11113);
nor U11601 (N_11601,N_11117,N_11340);
nor U11602 (N_11602,N_11107,N_11203);
xnor U11603 (N_11603,N_11278,N_11161);
xor U11604 (N_11604,N_11106,N_11006);
xor U11605 (N_11605,N_11395,N_11054);
nand U11606 (N_11606,N_11204,N_11131);
and U11607 (N_11607,N_11039,N_11375);
xnor U11608 (N_11608,N_11471,N_11366);
xor U11609 (N_11609,N_11321,N_11445);
nor U11610 (N_11610,N_11344,N_11346);
xnor U11611 (N_11611,N_11306,N_11142);
nor U11612 (N_11612,N_11427,N_11135);
and U11613 (N_11613,N_11162,N_11256);
nor U11614 (N_11614,N_11401,N_11352);
and U11615 (N_11615,N_11261,N_11489);
and U11616 (N_11616,N_11250,N_11128);
nand U11617 (N_11617,N_11479,N_11447);
xnor U11618 (N_11618,N_11363,N_11316);
or U11619 (N_11619,N_11485,N_11472);
nand U11620 (N_11620,N_11285,N_11283);
xnor U11621 (N_11621,N_11123,N_11378);
xnor U11622 (N_11622,N_11310,N_11174);
nor U11623 (N_11623,N_11369,N_11463);
nand U11624 (N_11624,N_11287,N_11213);
or U11625 (N_11625,N_11314,N_11455);
and U11626 (N_11626,N_11055,N_11197);
xor U11627 (N_11627,N_11379,N_11456);
nor U11628 (N_11628,N_11491,N_11133);
and U11629 (N_11629,N_11343,N_11073);
and U11630 (N_11630,N_11430,N_11194);
and U11631 (N_11631,N_11116,N_11403);
nor U11632 (N_11632,N_11434,N_11149);
nor U11633 (N_11633,N_11169,N_11299);
xor U11634 (N_11634,N_11168,N_11225);
or U11635 (N_11635,N_11028,N_11327);
nor U11636 (N_11636,N_11150,N_11103);
nand U11637 (N_11637,N_11461,N_11160);
and U11638 (N_11638,N_11221,N_11119);
nand U11639 (N_11639,N_11292,N_11072);
xnor U11640 (N_11640,N_11023,N_11183);
xnor U11641 (N_11641,N_11308,N_11223);
and U11642 (N_11642,N_11431,N_11017);
xor U11643 (N_11643,N_11227,N_11042);
or U11644 (N_11644,N_11139,N_11044);
and U11645 (N_11645,N_11407,N_11229);
and U11646 (N_11646,N_11282,N_11373);
and U11647 (N_11647,N_11490,N_11209);
nor U11648 (N_11648,N_11067,N_11468);
and U11649 (N_11649,N_11498,N_11193);
nor U11650 (N_11650,N_11078,N_11301);
nor U11651 (N_11651,N_11134,N_11015);
nand U11652 (N_11652,N_11172,N_11440);
or U11653 (N_11653,N_11381,N_11200);
nor U11654 (N_11654,N_11390,N_11126);
or U11655 (N_11655,N_11129,N_11365);
and U11656 (N_11656,N_11182,N_11038);
nor U11657 (N_11657,N_11170,N_11033);
xnor U11658 (N_11658,N_11380,N_11043);
and U11659 (N_11659,N_11165,N_11085);
nor U11660 (N_11660,N_11074,N_11388);
and U11661 (N_11661,N_11312,N_11478);
and U11662 (N_11662,N_11435,N_11050);
nor U11663 (N_11663,N_11318,N_11273);
nand U11664 (N_11664,N_11286,N_11132);
nor U11665 (N_11665,N_11269,N_11349);
and U11666 (N_11666,N_11101,N_11185);
or U11667 (N_11667,N_11190,N_11245);
nand U11668 (N_11668,N_11410,N_11178);
nand U11669 (N_11669,N_11419,N_11143);
nand U11670 (N_11670,N_11418,N_11473);
xor U11671 (N_11671,N_11069,N_11263);
nor U11672 (N_11672,N_11214,N_11034);
xnor U11673 (N_11673,N_11037,N_11342);
or U11674 (N_11674,N_11464,N_11158);
or U11675 (N_11675,N_11442,N_11248);
nor U11676 (N_11676,N_11339,N_11454);
xnor U11677 (N_11677,N_11323,N_11118);
and U11678 (N_11678,N_11336,N_11080);
nor U11679 (N_11679,N_11022,N_11271);
or U11680 (N_11680,N_11266,N_11420);
and U11681 (N_11681,N_11090,N_11399);
xor U11682 (N_11682,N_11120,N_11011);
or U11683 (N_11683,N_11382,N_11007);
or U11684 (N_11684,N_11241,N_11058);
or U11685 (N_11685,N_11127,N_11480);
and U11686 (N_11686,N_11392,N_11424);
nand U11687 (N_11687,N_11202,N_11004);
nand U11688 (N_11688,N_11428,N_11496);
or U11689 (N_11689,N_11001,N_11433);
and U11690 (N_11690,N_11469,N_11257);
xor U11691 (N_11691,N_11070,N_11088);
or U11692 (N_11692,N_11295,N_11415);
nand U11693 (N_11693,N_11077,N_11093);
nor U11694 (N_11694,N_11348,N_11049);
and U11695 (N_11695,N_11000,N_11156);
and U11696 (N_11696,N_11385,N_11477);
nor U11697 (N_11697,N_11360,N_11311);
xnor U11698 (N_11698,N_11254,N_11159);
or U11699 (N_11699,N_11260,N_11243);
nor U11700 (N_11700,N_11289,N_11394);
xor U11701 (N_11701,N_11173,N_11425);
nor U11702 (N_11702,N_11104,N_11141);
or U11703 (N_11703,N_11075,N_11016);
or U11704 (N_11704,N_11328,N_11387);
xor U11705 (N_11705,N_11277,N_11443);
xnor U11706 (N_11706,N_11291,N_11191);
and U11707 (N_11707,N_11099,N_11359);
or U11708 (N_11708,N_11384,N_11322);
xor U11709 (N_11709,N_11179,N_11234);
or U11710 (N_11710,N_11151,N_11338);
xor U11711 (N_11711,N_11176,N_11180);
nor U11712 (N_11712,N_11495,N_11216);
or U11713 (N_11713,N_11481,N_11002);
nor U11714 (N_11714,N_11222,N_11255);
and U11715 (N_11715,N_11356,N_11210);
xnor U11716 (N_11716,N_11030,N_11474);
and U11717 (N_11717,N_11499,N_11199);
or U11718 (N_11718,N_11087,N_11137);
or U11719 (N_11719,N_11224,N_11393);
and U11720 (N_11720,N_11060,N_11417);
nand U11721 (N_11721,N_11240,N_11288);
or U11722 (N_11722,N_11462,N_11406);
and U11723 (N_11723,N_11136,N_11275);
and U11724 (N_11724,N_11018,N_11056);
or U11725 (N_11725,N_11405,N_11293);
nor U11726 (N_11726,N_11320,N_11421);
xnor U11727 (N_11727,N_11095,N_11422);
or U11728 (N_11728,N_11062,N_11459);
xor U11729 (N_11729,N_11350,N_11423);
and U11730 (N_11730,N_11079,N_11186);
nand U11731 (N_11731,N_11302,N_11465);
nand U11732 (N_11732,N_11429,N_11175);
or U11733 (N_11733,N_11164,N_11147);
or U11734 (N_11734,N_11025,N_11020);
and U11735 (N_11735,N_11276,N_11324);
nor U11736 (N_11736,N_11397,N_11398);
or U11737 (N_11737,N_11163,N_11326);
or U11738 (N_11738,N_11188,N_11146);
nor U11739 (N_11739,N_11297,N_11279);
xor U11740 (N_11740,N_11014,N_11027);
nor U11741 (N_11741,N_11309,N_11230);
xnor U11742 (N_11742,N_11307,N_11012);
or U11743 (N_11743,N_11304,N_11154);
nor U11744 (N_11744,N_11281,N_11332);
nor U11745 (N_11745,N_11024,N_11370);
or U11746 (N_11746,N_11492,N_11045);
or U11747 (N_11747,N_11040,N_11029);
and U11748 (N_11748,N_11026,N_11483);
or U11749 (N_11749,N_11482,N_11242);
and U11750 (N_11750,N_11316,N_11233);
xor U11751 (N_11751,N_11422,N_11253);
and U11752 (N_11752,N_11006,N_11254);
and U11753 (N_11753,N_11212,N_11064);
nor U11754 (N_11754,N_11216,N_11120);
and U11755 (N_11755,N_11090,N_11195);
xor U11756 (N_11756,N_11339,N_11070);
nor U11757 (N_11757,N_11469,N_11345);
and U11758 (N_11758,N_11361,N_11098);
or U11759 (N_11759,N_11003,N_11380);
xor U11760 (N_11760,N_11223,N_11180);
or U11761 (N_11761,N_11359,N_11491);
nand U11762 (N_11762,N_11484,N_11203);
or U11763 (N_11763,N_11160,N_11108);
nor U11764 (N_11764,N_11426,N_11420);
xnor U11765 (N_11765,N_11260,N_11073);
xor U11766 (N_11766,N_11182,N_11335);
nor U11767 (N_11767,N_11154,N_11117);
nor U11768 (N_11768,N_11241,N_11238);
and U11769 (N_11769,N_11269,N_11043);
xnor U11770 (N_11770,N_11247,N_11427);
or U11771 (N_11771,N_11189,N_11255);
nand U11772 (N_11772,N_11208,N_11105);
or U11773 (N_11773,N_11299,N_11264);
nand U11774 (N_11774,N_11449,N_11117);
xor U11775 (N_11775,N_11151,N_11305);
xor U11776 (N_11776,N_11176,N_11256);
nand U11777 (N_11777,N_11474,N_11277);
xnor U11778 (N_11778,N_11353,N_11181);
xor U11779 (N_11779,N_11055,N_11121);
xor U11780 (N_11780,N_11415,N_11130);
or U11781 (N_11781,N_11267,N_11407);
or U11782 (N_11782,N_11405,N_11140);
nor U11783 (N_11783,N_11026,N_11107);
xnor U11784 (N_11784,N_11115,N_11334);
or U11785 (N_11785,N_11328,N_11153);
nor U11786 (N_11786,N_11430,N_11426);
and U11787 (N_11787,N_11271,N_11278);
and U11788 (N_11788,N_11002,N_11000);
xor U11789 (N_11789,N_11206,N_11062);
nor U11790 (N_11790,N_11457,N_11411);
xnor U11791 (N_11791,N_11456,N_11353);
nand U11792 (N_11792,N_11292,N_11194);
or U11793 (N_11793,N_11422,N_11111);
nor U11794 (N_11794,N_11134,N_11368);
nor U11795 (N_11795,N_11018,N_11036);
and U11796 (N_11796,N_11272,N_11078);
or U11797 (N_11797,N_11313,N_11208);
and U11798 (N_11798,N_11144,N_11218);
or U11799 (N_11799,N_11358,N_11380);
and U11800 (N_11800,N_11251,N_11433);
xnor U11801 (N_11801,N_11053,N_11190);
and U11802 (N_11802,N_11350,N_11142);
and U11803 (N_11803,N_11414,N_11274);
or U11804 (N_11804,N_11280,N_11470);
nand U11805 (N_11805,N_11043,N_11492);
nor U11806 (N_11806,N_11446,N_11371);
and U11807 (N_11807,N_11047,N_11393);
and U11808 (N_11808,N_11021,N_11413);
or U11809 (N_11809,N_11238,N_11181);
nor U11810 (N_11810,N_11248,N_11220);
and U11811 (N_11811,N_11404,N_11002);
and U11812 (N_11812,N_11142,N_11211);
xnor U11813 (N_11813,N_11427,N_11363);
xnor U11814 (N_11814,N_11055,N_11213);
or U11815 (N_11815,N_11028,N_11468);
nand U11816 (N_11816,N_11227,N_11269);
nor U11817 (N_11817,N_11011,N_11198);
nand U11818 (N_11818,N_11019,N_11416);
nand U11819 (N_11819,N_11100,N_11381);
nand U11820 (N_11820,N_11133,N_11406);
xnor U11821 (N_11821,N_11483,N_11054);
or U11822 (N_11822,N_11061,N_11302);
xor U11823 (N_11823,N_11017,N_11033);
xnor U11824 (N_11824,N_11451,N_11244);
nor U11825 (N_11825,N_11011,N_11237);
nand U11826 (N_11826,N_11419,N_11172);
nor U11827 (N_11827,N_11078,N_11057);
and U11828 (N_11828,N_11434,N_11376);
xnor U11829 (N_11829,N_11353,N_11209);
nor U11830 (N_11830,N_11317,N_11382);
and U11831 (N_11831,N_11065,N_11499);
and U11832 (N_11832,N_11303,N_11276);
xnor U11833 (N_11833,N_11296,N_11205);
or U11834 (N_11834,N_11389,N_11340);
xor U11835 (N_11835,N_11328,N_11440);
nand U11836 (N_11836,N_11151,N_11273);
nand U11837 (N_11837,N_11321,N_11011);
nand U11838 (N_11838,N_11438,N_11140);
or U11839 (N_11839,N_11201,N_11469);
xnor U11840 (N_11840,N_11284,N_11466);
and U11841 (N_11841,N_11250,N_11054);
nor U11842 (N_11842,N_11451,N_11010);
xnor U11843 (N_11843,N_11089,N_11122);
nor U11844 (N_11844,N_11351,N_11144);
xnor U11845 (N_11845,N_11059,N_11210);
or U11846 (N_11846,N_11100,N_11363);
or U11847 (N_11847,N_11193,N_11410);
xor U11848 (N_11848,N_11042,N_11366);
and U11849 (N_11849,N_11408,N_11320);
or U11850 (N_11850,N_11233,N_11485);
or U11851 (N_11851,N_11468,N_11167);
xor U11852 (N_11852,N_11135,N_11143);
nand U11853 (N_11853,N_11158,N_11241);
and U11854 (N_11854,N_11492,N_11430);
nor U11855 (N_11855,N_11443,N_11317);
xor U11856 (N_11856,N_11364,N_11450);
or U11857 (N_11857,N_11285,N_11256);
or U11858 (N_11858,N_11304,N_11081);
nor U11859 (N_11859,N_11288,N_11429);
nor U11860 (N_11860,N_11351,N_11255);
nand U11861 (N_11861,N_11243,N_11189);
or U11862 (N_11862,N_11390,N_11491);
and U11863 (N_11863,N_11212,N_11052);
nor U11864 (N_11864,N_11449,N_11366);
and U11865 (N_11865,N_11059,N_11369);
nand U11866 (N_11866,N_11201,N_11135);
nand U11867 (N_11867,N_11174,N_11146);
nor U11868 (N_11868,N_11170,N_11358);
and U11869 (N_11869,N_11358,N_11298);
nor U11870 (N_11870,N_11204,N_11096);
or U11871 (N_11871,N_11015,N_11230);
nand U11872 (N_11872,N_11423,N_11246);
and U11873 (N_11873,N_11420,N_11377);
nor U11874 (N_11874,N_11254,N_11458);
xor U11875 (N_11875,N_11223,N_11182);
xnor U11876 (N_11876,N_11327,N_11050);
and U11877 (N_11877,N_11482,N_11498);
or U11878 (N_11878,N_11127,N_11465);
xor U11879 (N_11879,N_11287,N_11000);
or U11880 (N_11880,N_11199,N_11161);
nand U11881 (N_11881,N_11283,N_11117);
and U11882 (N_11882,N_11306,N_11366);
and U11883 (N_11883,N_11251,N_11123);
or U11884 (N_11884,N_11147,N_11413);
or U11885 (N_11885,N_11067,N_11356);
or U11886 (N_11886,N_11159,N_11172);
xor U11887 (N_11887,N_11062,N_11110);
xnor U11888 (N_11888,N_11365,N_11385);
nor U11889 (N_11889,N_11475,N_11463);
xnor U11890 (N_11890,N_11251,N_11056);
or U11891 (N_11891,N_11259,N_11122);
and U11892 (N_11892,N_11213,N_11096);
and U11893 (N_11893,N_11335,N_11096);
nor U11894 (N_11894,N_11494,N_11065);
xor U11895 (N_11895,N_11051,N_11454);
xor U11896 (N_11896,N_11239,N_11334);
nor U11897 (N_11897,N_11191,N_11125);
nand U11898 (N_11898,N_11020,N_11301);
nand U11899 (N_11899,N_11212,N_11375);
and U11900 (N_11900,N_11431,N_11118);
and U11901 (N_11901,N_11274,N_11167);
and U11902 (N_11902,N_11419,N_11372);
and U11903 (N_11903,N_11106,N_11215);
nand U11904 (N_11904,N_11238,N_11351);
xor U11905 (N_11905,N_11256,N_11420);
or U11906 (N_11906,N_11146,N_11429);
and U11907 (N_11907,N_11084,N_11133);
nand U11908 (N_11908,N_11313,N_11073);
or U11909 (N_11909,N_11245,N_11481);
and U11910 (N_11910,N_11303,N_11490);
and U11911 (N_11911,N_11082,N_11490);
nand U11912 (N_11912,N_11201,N_11262);
and U11913 (N_11913,N_11206,N_11023);
xnor U11914 (N_11914,N_11247,N_11258);
or U11915 (N_11915,N_11415,N_11338);
nor U11916 (N_11916,N_11008,N_11244);
and U11917 (N_11917,N_11094,N_11121);
and U11918 (N_11918,N_11049,N_11025);
or U11919 (N_11919,N_11347,N_11414);
xor U11920 (N_11920,N_11365,N_11323);
and U11921 (N_11921,N_11430,N_11230);
and U11922 (N_11922,N_11131,N_11166);
nand U11923 (N_11923,N_11358,N_11132);
and U11924 (N_11924,N_11241,N_11150);
nand U11925 (N_11925,N_11424,N_11117);
xor U11926 (N_11926,N_11230,N_11462);
nand U11927 (N_11927,N_11369,N_11441);
nand U11928 (N_11928,N_11330,N_11447);
nor U11929 (N_11929,N_11437,N_11154);
nor U11930 (N_11930,N_11142,N_11199);
or U11931 (N_11931,N_11087,N_11230);
or U11932 (N_11932,N_11052,N_11177);
xnor U11933 (N_11933,N_11081,N_11417);
and U11934 (N_11934,N_11066,N_11329);
and U11935 (N_11935,N_11036,N_11042);
xnor U11936 (N_11936,N_11180,N_11214);
nor U11937 (N_11937,N_11398,N_11345);
xor U11938 (N_11938,N_11166,N_11201);
and U11939 (N_11939,N_11272,N_11115);
nor U11940 (N_11940,N_11280,N_11187);
nand U11941 (N_11941,N_11282,N_11334);
xor U11942 (N_11942,N_11034,N_11482);
or U11943 (N_11943,N_11476,N_11345);
xor U11944 (N_11944,N_11045,N_11202);
and U11945 (N_11945,N_11462,N_11380);
and U11946 (N_11946,N_11195,N_11280);
and U11947 (N_11947,N_11031,N_11418);
xor U11948 (N_11948,N_11310,N_11335);
nor U11949 (N_11949,N_11092,N_11222);
and U11950 (N_11950,N_11491,N_11271);
or U11951 (N_11951,N_11278,N_11173);
and U11952 (N_11952,N_11234,N_11429);
nor U11953 (N_11953,N_11369,N_11037);
and U11954 (N_11954,N_11335,N_11377);
xor U11955 (N_11955,N_11329,N_11134);
xor U11956 (N_11956,N_11166,N_11295);
and U11957 (N_11957,N_11327,N_11150);
nand U11958 (N_11958,N_11455,N_11359);
xnor U11959 (N_11959,N_11193,N_11024);
nand U11960 (N_11960,N_11351,N_11096);
nor U11961 (N_11961,N_11144,N_11217);
xnor U11962 (N_11962,N_11277,N_11164);
and U11963 (N_11963,N_11124,N_11488);
or U11964 (N_11964,N_11135,N_11306);
and U11965 (N_11965,N_11011,N_11431);
and U11966 (N_11966,N_11403,N_11405);
and U11967 (N_11967,N_11240,N_11430);
nand U11968 (N_11968,N_11276,N_11012);
nor U11969 (N_11969,N_11490,N_11463);
xnor U11970 (N_11970,N_11255,N_11072);
and U11971 (N_11971,N_11234,N_11192);
nor U11972 (N_11972,N_11397,N_11005);
nor U11973 (N_11973,N_11243,N_11041);
and U11974 (N_11974,N_11364,N_11025);
nand U11975 (N_11975,N_11264,N_11330);
xor U11976 (N_11976,N_11369,N_11027);
nor U11977 (N_11977,N_11068,N_11410);
and U11978 (N_11978,N_11471,N_11470);
nor U11979 (N_11979,N_11177,N_11200);
or U11980 (N_11980,N_11236,N_11315);
or U11981 (N_11981,N_11421,N_11100);
xnor U11982 (N_11982,N_11335,N_11013);
nor U11983 (N_11983,N_11297,N_11243);
and U11984 (N_11984,N_11396,N_11393);
nor U11985 (N_11985,N_11343,N_11081);
and U11986 (N_11986,N_11290,N_11294);
nand U11987 (N_11987,N_11154,N_11319);
nand U11988 (N_11988,N_11168,N_11319);
or U11989 (N_11989,N_11221,N_11412);
or U11990 (N_11990,N_11113,N_11444);
nand U11991 (N_11991,N_11125,N_11016);
or U11992 (N_11992,N_11309,N_11458);
xnor U11993 (N_11993,N_11030,N_11251);
and U11994 (N_11994,N_11460,N_11266);
nor U11995 (N_11995,N_11378,N_11122);
and U11996 (N_11996,N_11265,N_11096);
nand U11997 (N_11997,N_11326,N_11371);
and U11998 (N_11998,N_11135,N_11015);
xnor U11999 (N_11999,N_11488,N_11345);
and U12000 (N_12000,N_11506,N_11782);
nor U12001 (N_12001,N_11943,N_11770);
nand U12002 (N_12002,N_11982,N_11542);
and U12003 (N_12003,N_11895,N_11618);
and U12004 (N_12004,N_11511,N_11749);
and U12005 (N_12005,N_11956,N_11834);
or U12006 (N_12006,N_11548,N_11900);
xor U12007 (N_12007,N_11758,N_11766);
nand U12008 (N_12008,N_11888,N_11623);
and U12009 (N_12009,N_11820,N_11557);
nor U12010 (N_12010,N_11953,N_11790);
and U12011 (N_12011,N_11889,N_11894);
or U12012 (N_12012,N_11773,N_11891);
nor U12013 (N_12013,N_11691,N_11979);
xor U12014 (N_12014,N_11753,N_11692);
xor U12015 (N_12015,N_11986,N_11752);
or U12016 (N_12016,N_11510,N_11908);
nand U12017 (N_12017,N_11699,N_11947);
xnor U12018 (N_12018,N_11729,N_11564);
and U12019 (N_12019,N_11672,N_11757);
or U12020 (N_12020,N_11960,N_11576);
nand U12021 (N_12021,N_11886,N_11765);
and U12022 (N_12022,N_11617,N_11660);
and U12023 (N_12023,N_11917,N_11911);
and U12024 (N_12024,N_11722,N_11771);
or U12025 (N_12025,N_11973,N_11817);
xnor U12026 (N_12026,N_11844,N_11852);
or U12027 (N_12027,N_11551,N_11901);
and U12028 (N_12028,N_11880,N_11735);
nor U12029 (N_12029,N_11969,N_11724);
and U12030 (N_12030,N_11619,N_11650);
nor U12031 (N_12031,N_11815,N_11893);
nor U12032 (N_12032,N_11946,N_11818);
and U12033 (N_12033,N_11955,N_11529);
and U12034 (N_12034,N_11715,N_11832);
or U12035 (N_12035,N_11988,N_11705);
nand U12036 (N_12036,N_11666,N_11862);
and U12037 (N_12037,N_11823,N_11741);
nand U12038 (N_12038,N_11840,N_11581);
nand U12039 (N_12039,N_11858,N_11727);
xnor U12040 (N_12040,N_11683,N_11812);
and U12041 (N_12041,N_11739,N_11904);
or U12042 (N_12042,N_11696,N_11658);
nor U12043 (N_12043,N_11589,N_11676);
and U12044 (N_12044,N_11583,N_11974);
or U12045 (N_12045,N_11546,N_11926);
and U12046 (N_12046,N_11731,N_11942);
and U12047 (N_12047,N_11554,N_11962);
xor U12048 (N_12048,N_11689,N_11851);
nor U12049 (N_12049,N_11994,N_11958);
or U12050 (N_12050,N_11664,N_11737);
nor U12051 (N_12051,N_11780,N_11952);
and U12052 (N_12052,N_11688,N_11698);
or U12053 (N_12053,N_11949,N_11605);
or U12054 (N_12054,N_11980,N_11668);
or U12055 (N_12055,N_11686,N_11543);
nor U12056 (N_12056,N_11938,N_11788);
xnor U12057 (N_12057,N_11923,N_11675);
nor U12058 (N_12058,N_11656,N_11821);
nand U12059 (N_12059,N_11622,N_11981);
or U12060 (N_12060,N_11630,N_11584);
nor U12061 (N_12061,N_11503,N_11625);
or U12062 (N_12062,N_11667,N_11961);
nand U12063 (N_12063,N_11927,N_11703);
nor U12064 (N_12064,N_11636,N_11701);
nor U12065 (N_12065,N_11754,N_11977);
and U12066 (N_12066,N_11620,N_11892);
nand U12067 (N_12067,N_11867,N_11756);
and U12068 (N_12068,N_11802,N_11711);
and U12069 (N_12069,N_11929,N_11940);
nor U12070 (N_12070,N_11507,N_11504);
xor U12071 (N_12071,N_11641,N_11582);
nor U12072 (N_12072,N_11992,N_11747);
and U12073 (N_12073,N_11580,N_11919);
xor U12074 (N_12074,N_11531,N_11903);
and U12075 (N_12075,N_11539,N_11856);
xor U12076 (N_12076,N_11935,N_11514);
nor U12077 (N_12077,N_11755,N_11570);
nor U12078 (N_12078,N_11518,N_11781);
or U12079 (N_12079,N_11663,N_11744);
or U12080 (N_12080,N_11931,N_11671);
nand U12081 (N_12081,N_11918,N_11505);
nand U12082 (N_12082,N_11833,N_11968);
xnor U12083 (N_12083,N_11954,N_11651);
and U12084 (N_12084,N_11657,N_11789);
xnor U12085 (N_12085,N_11613,N_11750);
or U12086 (N_12086,N_11574,N_11816);
nor U12087 (N_12087,N_11987,N_11611);
and U12088 (N_12088,N_11995,N_11996);
xor U12089 (N_12089,N_11745,N_11924);
and U12090 (N_12090,N_11855,N_11595);
and U12091 (N_12091,N_11951,N_11990);
xor U12092 (N_12092,N_11674,N_11829);
xnor U12093 (N_12093,N_11971,N_11612);
nand U12094 (N_12094,N_11615,N_11945);
xnor U12095 (N_12095,N_11556,N_11578);
nand U12096 (N_12096,N_11843,N_11603);
or U12097 (N_12097,N_11567,N_11680);
and U12098 (N_12098,N_11640,N_11870);
or U12099 (N_12099,N_11759,N_11714);
nor U12100 (N_12100,N_11984,N_11972);
and U12101 (N_12101,N_11523,N_11873);
nand U12102 (N_12102,N_11909,N_11922);
or U12103 (N_12103,N_11861,N_11704);
xor U12104 (N_12104,N_11872,N_11594);
and U12105 (N_12105,N_11720,N_11937);
nor U12106 (N_12106,N_11848,N_11760);
nand U12107 (N_12107,N_11608,N_11519);
or U12108 (N_12108,N_11586,N_11875);
and U12109 (N_12109,N_11598,N_11793);
xor U12110 (N_12110,N_11694,N_11934);
nand U12111 (N_12111,N_11648,N_11646);
xor U12112 (N_12112,N_11628,N_11786);
and U12113 (N_12113,N_11649,N_11562);
or U12114 (N_12114,N_11600,N_11849);
nand U12115 (N_12115,N_11881,N_11728);
nor U12116 (N_12116,N_11999,N_11627);
or U12117 (N_12117,N_11621,N_11614);
nand U12118 (N_12118,N_11563,N_11547);
and U12119 (N_12119,N_11525,N_11500);
nand U12120 (N_12120,N_11535,N_11544);
nand U12121 (N_12121,N_11734,N_11702);
xnor U12122 (N_12122,N_11796,N_11879);
nor U12123 (N_12123,N_11805,N_11502);
or U12124 (N_12124,N_11763,N_11743);
or U12125 (N_12125,N_11808,N_11565);
nor U12126 (N_12126,N_11647,N_11635);
nor U12127 (N_12127,N_11606,N_11957);
nor U12128 (N_12128,N_11568,N_11721);
xor U12129 (N_12129,N_11585,N_11509);
xnor U12130 (N_12130,N_11939,N_11930);
and U12131 (N_12131,N_11963,N_11898);
nor U12132 (N_12132,N_11865,N_11874);
nor U12133 (N_12133,N_11824,N_11662);
nand U12134 (N_12134,N_11890,N_11806);
nand U12135 (N_12135,N_11807,N_11644);
xnor U12136 (N_12136,N_11526,N_11921);
nor U12137 (N_12137,N_11804,N_11677);
nand U12138 (N_12138,N_11896,N_11533);
xnor U12139 (N_12139,N_11607,N_11932);
xnor U12140 (N_12140,N_11882,N_11966);
or U12141 (N_12141,N_11515,N_11826);
nand U12142 (N_12142,N_11764,N_11777);
or U12143 (N_12143,N_11738,N_11776);
and U12144 (N_12144,N_11545,N_11751);
or U12145 (N_12145,N_11733,N_11725);
nand U12146 (N_12146,N_11637,N_11964);
nand U12147 (N_12147,N_11959,N_11588);
nand U12148 (N_12148,N_11521,N_11853);
nor U12149 (N_12149,N_11775,N_11690);
nor U12150 (N_12150,N_11813,N_11883);
xor U12151 (N_12151,N_11869,N_11508);
nand U12152 (N_12152,N_11626,N_11885);
or U12153 (N_12153,N_11559,N_11501);
nand U12154 (N_12154,N_11700,N_11730);
or U12155 (N_12155,N_11723,N_11708);
nand U12156 (N_12156,N_11948,N_11860);
nor U12157 (N_12157,N_11912,N_11876);
nand U12158 (N_12158,N_11732,N_11516);
or U12159 (N_12159,N_11707,N_11643);
xor U12160 (N_12160,N_11587,N_11769);
nand U12161 (N_12161,N_11993,N_11941);
xor U12162 (N_12162,N_11654,N_11566);
nand U12163 (N_12163,N_11520,N_11902);
nand U12164 (N_12164,N_11897,N_11884);
nor U12165 (N_12165,N_11592,N_11681);
and U12166 (N_12166,N_11762,N_11652);
nand U12167 (N_12167,N_11528,N_11825);
and U12168 (N_12168,N_11845,N_11847);
xor U12169 (N_12169,N_11524,N_11639);
xnor U12170 (N_12170,N_11916,N_11846);
or U12171 (N_12171,N_11772,N_11837);
or U12172 (N_12172,N_11800,N_11854);
or U12173 (N_12173,N_11712,N_11944);
nor U12174 (N_12174,N_11803,N_11717);
or U12175 (N_12175,N_11642,N_11810);
and U12176 (N_12176,N_11561,N_11591);
or U12177 (N_12177,N_11835,N_11706);
xor U12178 (N_12178,N_11719,N_11695);
nand U12179 (N_12179,N_11602,N_11634);
xor U12180 (N_12180,N_11967,N_11549);
xnor U12181 (N_12181,N_11631,N_11799);
and U12182 (N_12182,N_11983,N_11599);
nand U12183 (N_12183,N_11522,N_11716);
nor U12184 (N_12184,N_11517,N_11905);
xnor U12185 (N_12185,N_11596,N_11682);
and U12186 (N_12186,N_11936,N_11536);
nor U12187 (N_12187,N_11558,N_11604);
and U12188 (N_12188,N_11693,N_11985);
nand U12189 (N_12189,N_11831,N_11597);
nor U12190 (N_12190,N_11670,N_11784);
nand U12191 (N_12191,N_11998,N_11774);
nand U12192 (N_12192,N_11537,N_11907);
and U12193 (N_12193,N_11798,N_11513);
xor U12194 (N_12194,N_11797,N_11809);
nand U12195 (N_12195,N_11709,N_11828);
or U12196 (N_12196,N_11684,N_11778);
nor U12197 (N_12197,N_11975,N_11838);
xor U12198 (N_12198,N_11645,N_11553);
nand U12199 (N_12199,N_11830,N_11633);
or U12200 (N_12200,N_11761,N_11748);
nor U12201 (N_12201,N_11575,N_11965);
xor U12202 (N_12202,N_11697,N_11857);
or U12203 (N_12203,N_11933,N_11841);
xor U12204 (N_12204,N_11560,N_11629);
and U12205 (N_12205,N_11742,N_11573);
and U12206 (N_12206,N_11920,N_11877);
and U12207 (N_12207,N_11632,N_11791);
nand U12208 (N_12208,N_11795,N_11878);
nand U12209 (N_12209,N_11736,N_11779);
and U12210 (N_12210,N_11726,N_11887);
or U12211 (N_12211,N_11767,N_11819);
or U12212 (N_12212,N_11997,N_11991);
xor U12213 (N_12213,N_11638,N_11822);
xnor U12214 (N_12214,N_11864,N_11792);
or U12215 (N_12215,N_11794,N_11624);
nand U12216 (N_12216,N_11685,N_11915);
or U12217 (N_12217,N_11866,N_11593);
or U12218 (N_12218,N_11512,N_11740);
and U12219 (N_12219,N_11814,N_11655);
or U12220 (N_12220,N_11577,N_11906);
nor U12221 (N_12221,N_11910,N_11669);
and U12222 (N_12222,N_11746,N_11811);
xnor U12223 (N_12223,N_11678,N_11610);
nand U12224 (N_12224,N_11836,N_11787);
xnor U12225 (N_12225,N_11571,N_11768);
or U12226 (N_12226,N_11538,N_11653);
or U12227 (N_12227,N_11579,N_11801);
nand U12228 (N_12228,N_11527,N_11616);
nand U12229 (N_12229,N_11928,N_11785);
nor U12230 (N_12230,N_11673,N_11925);
or U12231 (N_12231,N_11552,N_11540);
and U12232 (N_12232,N_11913,N_11868);
or U12233 (N_12233,N_11569,N_11718);
xor U12234 (N_12234,N_11978,N_11532);
xor U12235 (N_12235,N_11859,N_11976);
xnor U12236 (N_12236,N_11914,N_11555);
nor U12237 (N_12237,N_11550,N_11530);
xnor U12238 (N_12238,N_11609,N_11899);
xor U12239 (N_12239,N_11863,N_11783);
nand U12240 (N_12240,N_11601,N_11871);
or U12241 (N_12241,N_11950,N_11665);
nor U12242 (N_12242,N_11710,N_11590);
nor U12243 (N_12243,N_11827,N_11661);
or U12244 (N_12244,N_11989,N_11572);
and U12245 (N_12245,N_11687,N_11839);
and U12246 (N_12246,N_11659,N_11970);
xnor U12247 (N_12247,N_11842,N_11534);
nor U12248 (N_12248,N_11679,N_11541);
nor U12249 (N_12249,N_11713,N_11850);
nand U12250 (N_12250,N_11989,N_11850);
nand U12251 (N_12251,N_11933,N_11957);
xor U12252 (N_12252,N_11785,N_11981);
or U12253 (N_12253,N_11727,N_11628);
nand U12254 (N_12254,N_11805,N_11712);
or U12255 (N_12255,N_11646,N_11581);
xnor U12256 (N_12256,N_11627,N_11842);
nor U12257 (N_12257,N_11799,N_11734);
xor U12258 (N_12258,N_11892,N_11676);
nand U12259 (N_12259,N_11793,N_11919);
xnor U12260 (N_12260,N_11893,N_11712);
xnor U12261 (N_12261,N_11582,N_11536);
nor U12262 (N_12262,N_11694,N_11919);
nand U12263 (N_12263,N_11589,N_11691);
nor U12264 (N_12264,N_11577,N_11560);
or U12265 (N_12265,N_11965,N_11971);
and U12266 (N_12266,N_11856,N_11627);
xor U12267 (N_12267,N_11621,N_11626);
or U12268 (N_12268,N_11564,N_11942);
nor U12269 (N_12269,N_11613,N_11695);
nand U12270 (N_12270,N_11520,N_11652);
nor U12271 (N_12271,N_11604,N_11640);
or U12272 (N_12272,N_11670,N_11836);
xnor U12273 (N_12273,N_11658,N_11581);
xor U12274 (N_12274,N_11930,N_11660);
or U12275 (N_12275,N_11709,N_11599);
and U12276 (N_12276,N_11543,N_11903);
nor U12277 (N_12277,N_11656,N_11518);
nor U12278 (N_12278,N_11827,N_11806);
nor U12279 (N_12279,N_11914,N_11879);
nand U12280 (N_12280,N_11939,N_11986);
nand U12281 (N_12281,N_11960,N_11801);
or U12282 (N_12282,N_11805,N_11840);
xor U12283 (N_12283,N_11701,N_11944);
nand U12284 (N_12284,N_11527,N_11615);
xor U12285 (N_12285,N_11657,N_11986);
and U12286 (N_12286,N_11619,N_11628);
or U12287 (N_12287,N_11743,N_11854);
xnor U12288 (N_12288,N_11811,N_11721);
and U12289 (N_12289,N_11548,N_11590);
nor U12290 (N_12290,N_11874,N_11524);
or U12291 (N_12291,N_11734,N_11917);
and U12292 (N_12292,N_11934,N_11888);
and U12293 (N_12293,N_11982,N_11969);
and U12294 (N_12294,N_11922,N_11932);
and U12295 (N_12295,N_11797,N_11962);
or U12296 (N_12296,N_11645,N_11592);
and U12297 (N_12297,N_11875,N_11727);
nor U12298 (N_12298,N_11705,N_11897);
nor U12299 (N_12299,N_11876,N_11748);
or U12300 (N_12300,N_11920,N_11965);
nor U12301 (N_12301,N_11609,N_11742);
or U12302 (N_12302,N_11621,N_11881);
xor U12303 (N_12303,N_11897,N_11541);
xnor U12304 (N_12304,N_11557,N_11628);
xnor U12305 (N_12305,N_11633,N_11775);
nor U12306 (N_12306,N_11731,N_11771);
or U12307 (N_12307,N_11584,N_11780);
nand U12308 (N_12308,N_11998,N_11809);
nand U12309 (N_12309,N_11618,N_11682);
and U12310 (N_12310,N_11556,N_11819);
and U12311 (N_12311,N_11798,N_11875);
nor U12312 (N_12312,N_11939,N_11560);
nand U12313 (N_12313,N_11637,N_11815);
or U12314 (N_12314,N_11595,N_11784);
or U12315 (N_12315,N_11663,N_11559);
or U12316 (N_12316,N_11613,N_11620);
or U12317 (N_12317,N_11869,N_11600);
xor U12318 (N_12318,N_11552,N_11584);
nand U12319 (N_12319,N_11976,N_11752);
nor U12320 (N_12320,N_11687,N_11552);
nand U12321 (N_12321,N_11804,N_11985);
nand U12322 (N_12322,N_11676,N_11634);
xnor U12323 (N_12323,N_11886,N_11526);
xor U12324 (N_12324,N_11562,N_11780);
xor U12325 (N_12325,N_11658,N_11873);
nand U12326 (N_12326,N_11763,N_11985);
xnor U12327 (N_12327,N_11634,N_11527);
xnor U12328 (N_12328,N_11511,N_11564);
nand U12329 (N_12329,N_11913,N_11514);
and U12330 (N_12330,N_11993,N_11719);
nor U12331 (N_12331,N_11601,N_11520);
xnor U12332 (N_12332,N_11896,N_11999);
nand U12333 (N_12333,N_11649,N_11657);
nor U12334 (N_12334,N_11699,N_11940);
xor U12335 (N_12335,N_11518,N_11980);
and U12336 (N_12336,N_11635,N_11545);
or U12337 (N_12337,N_11876,N_11526);
nor U12338 (N_12338,N_11815,N_11619);
xnor U12339 (N_12339,N_11760,N_11672);
or U12340 (N_12340,N_11645,N_11748);
and U12341 (N_12341,N_11927,N_11854);
nand U12342 (N_12342,N_11840,N_11640);
or U12343 (N_12343,N_11797,N_11955);
nor U12344 (N_12344,N_11944,N_11935);
and U12345 (N_12345,N_11608,N_11897);
nor U12346 (N_12346,N_11841,N_11667);
and U12347 (N_12347,N_11892,N_11735);
or U12348 (N_12348,N_11802,N_11620);
and U12349 (N_12349,N_11811,N_11601);
nand U12350 (N_12350,N_11638,N_11774);
and U12351 (N_12351,N_11553,N_11938);
and U12352 (N_12352,N_11997,N_11716);
or U12353 (N_12353,N_11837,N_11730);
and U12354 (N_12354,N_11974,N_11910);
and U12355 (N_12355,N_11856,N_11886);
nand U12356 (N_12356,N_11666,N_11893);
or U12357 (N_12357,N_11548,N_11898);
xor U12358 (N_12358,N_11605,N_11754);
or U12359 (N_12359,N_11859,N_11916);
or U12360 (N_12360,N_11888,N_11658);
xor U12361 (N_12361,N_11873,N_11602);
and U12362 (N_12362,N_11679,N_11831);
and U12363 (N_12363,N_11801,N_11671);
and U12364 (N_12364,N_11856,N_11873);
or U12365 (N_12365,N_11930,N_11808);
nor U12366 (N_12366,N_11908,N_11971);
or U12367 (N_12367,N_11621,N_11846);
nand U12368 (N_12368,N_11590,N_11605);
nor U12369 (N_12369,N_11558,N_11905);
nand U12370 (N_12370,N_11664,N_11876);
and U12371 (N_12371,N_11536,N_11529);
and U12372 (N_12372,N_11678,N_11888);
nand U12373 (N_12373,N_11559,N_11704);
or U12374 (N_12374,N_11612,N_11851);
nand U12375 (N_12375,N_11595,N_11858);
and U12376 (N_12376,N_11791,N_11931);
nand U12377 (N_12377,N_11968,N_11988);
nor U12378 (N_12378,N_11800,N_11658);
nor U12379 (N_12379,N_11778,N_11565);
and U12380 (N_12380,N_11649,N_11514);
xor U12381 (N_12381,N_11842,N_11966);
xnor U12382 (N_12382,N_11928,N_11938);
or U12383 (N_12383,N_11616,N_11613);
nand U12384 (N_12384,N_11531,N_11607);
nor U12385 (N_12385,N_11759,N_11779);
or U12386 (N_12386,N_11604,N_11522);
and U12387 (N_12387,N_11675,N_11751);
or U12388 (N_12388,N_11867,N_11714);
and U12389 (N_12389,N_11719,N_11827);
and U12390 (N_12390,N_11981,N_11741);
nor U12391 (N_12391,N_11649,N_11599);
nand U12392 (N_12392,N_11831,N_11513);
and U12393 (N_12393,N_11906,N_11852);
and U12394 (N_12394,N_11722,N_11981);
or U12395 (N_12395,N_11647,N_11745);
nand U12396 (N_12396,N_11895,N_11892);
nor U12397 (N_12397,N_11788,N_11577);
xor U12398 (N_12398,N_11609,N_11795);
and U12399 (N_12399,N_11934,N_11927);
xor U12400 (N_12400,N_11814,N_11800);
nor U12401 (N_12401,N_11913,N_11716);
and U12402 (N_12402,N_11586,N_11607);
xor U12403 (N_12403,N_11681,N_11713);
nor U12404 (N_12404,N_11758,N_11519);
or U12405 (N_12405,N_11685,N_11736);
and U12406 (N_12406,N_11628,N_11941);
xor U12407 (N_12407,N_11824,N_11757);
nor U12408 (N_12408,N_11918,N_11669);
and U12409 (N_12409,N_11601,N_11810);
and U12410 (N_12410,N_11704,N_11876);
nand U12411 (N_12411,N_11638,N_11845);
or U12412 (N_12412,N_11921,N_11780);
and U12413 (N_12413,N_11758,N_11764);
and U12414 (N_12414,N_11934,N_11795);
and U12415 (N_12415,N_11589,N_11646);
and U12416 (N_12416,N_11683,N_11607);
or U12417 (N_12417,N_11631,N_11668);
or U12418 (N_12418,N_11538,N_11596);
or U12419 (N_12419,N_11802,N_11837);
and U12420 (N_12420,N_11882,N_11650);
nand U12421 (N_12421,N_11890,N_11667);
nor U12422 (N_12422,N_11545,N_11748);
or U12423 (N_12423,N_11810,N_11747);
or U12424 (N_12424,N_11872,N_11619);
or U12425 (N_12425,N_11843,N_11729);
and U12426 (N_12426,N_11649,N_11801);
or U12427 (N_12427,N_11661,N_11583);
nand U12428 (N_12428,N_11934,N_11654);
xor U12429 (N_12429,N_11862,N_11681);
and U12430 (N_12430,N_11620,N_11610);
nand U12431 (N_12431,N_11740,N_11811);
xor U12432 (N_12432,N_11668,N_11531);
and U12433 (N_12433,N_11600,N_11716);
nand U12434 (N_12434,N_11911,N_11553);
nand U12435 (N_12435,N_11911,N_11854);
nand U12436 (N_12436,N_11631,N_11641);
and U12437 (N_12437,N_11732,N_11873);
or U12438 (N_12438,N_11846,N_11905);
nor U12439 (N_12439,N_11889,N_11837);
and U12440 (N_12440,N_11756,N_11637);
and U12441 (N_12441,N_11740,N_11621);
or U12442 (N_12442,N_11761,N_11553);
or U12443 (N_12443,N_11720,N_11501);
or U12444 (N_12444,N_11582,N_11697);
or U12445 (N_12445,N_11531,N_11761);
xor U12446 (N_12446,N_11592,N_11898);
or U12447 (N_12447,N_11655,N_11816);
xnor U12448 (N_12448,N_11916,N_11766);
nor U12449 (N_12449,N_11895,N_11603);
and U12450 (N_12450,N_11904,N_11764);
nand U12451 (N_12451,N_11841,N_11813);
nand U12452 (N_12452,N_11656,N_11586);
nand U12453 (N_12453,N_11527,N_11980);
or U12454 (N_12454,N_11706,N_11679);
and U12455 (N_12455,N_11590,N_11538);
nand U12456 (N_12456,N_11979,N_11788);
nor U12457 (N_12457,N_11515,N_11921);
xor U12458 (N_12458,N_11661,N_11667);
xnor U12459 (N_12459,N_11946,N_11532);
or U12460 (N_12460,N_11982,N_11509);
and U12461 (N_12461,N_11578,N_11849);
nand U12462 (N_12462,N_11750,N_11952);
nand U12463 (N_12463,N_11685,N_11564);
and U12464 (N_12464,N_11706,N_11560);
nand U12465 (N_12465,N_11819,N_11661);
nand U12466 (N_12466,N_11559,N_11961);
nor U12467 (N_12467,N_11996,N_11610);
or U12468 (N_12468,N_11505,N_11849);
and U12469 (N_12469,N_11833,N_11954);
nor U12470 (N_12470,N_11749,N_11588);
nand U12471 (N_12471,N_11732,N_11945);
and U12472 (N_12472,N_11902,N_11870);
xor U12473 (N_12473,N_11946,N_11604);
nor U12474 (N_12474,N_11889,N_11750);
nand U12475 (N_12475,N_11786,N_11875);
nor U12476 (N_12476,N_11517,N_11864);
or U12477 (N_12477,N_11691,N_11515);
nand U12478 (N_12478,N_11779,N_11760);
nor U12479 (N_12479,N_11964,N_11557);
nor U12480 (N_12480,N_11661,N_11589);
and U12481 (N_12481,N_11850,N_11625);
nand U12482 (N_12482,N_11521,N_11535);
or U12483 (N_12483,N_11855,N_11923);
nand U12484 (N_12484,N_11870,N_11814);
and U12485 (N_12485,N_11713,N_11893);
nor U12486 (N_12486,N_11799,N_11998);
xnor U12487 (N_12487,N_11898,N_11922);
xnor U12488 (N_12488,N_11693,N_11967);
nand U12489 (N_12489,N_11620,N_11875);
and U12490 (N_12490,N_11993,N_11868);
nand U12491 (N_12491,N_11925,N_11589);
xnor U12492 (N_12492,N_11660,N_11673);
or U12493 (N_12493,N_11724,N_11648);
and U12494 (N_12494,N_11636,N_11672);
nand U12495 (N_12495,N_11992,N_11606);
or U12496 (N_12496,N_11916,N_11657);
and U12497 (N_12497,N_11880,N_11705);
nor U12498 (N_12498,N_11523,N_11610);
xor U12499 (N_12499,N_11992,N_11545);
nor U12500 (N_12500,N_12331,N_12301);
nand U12501 (N_12501,N_12265,N_12033);
xor U12502 (N_12502,N_12326,N_12041);
nor U12503 (N_12503,N_12111,N_12146);
nand U12504 (N_12504,N_12464,N_12225);
and U12505 (N_12505,N_12244,N_12491);
nand U12506 (N_12506,N_12299,N_12160);
xnor U12507 (N_12507,N_12040,N_12298);
nand U12508 (N_12508,N_12106,N_12404);
and U12509 (N_12509,N_12313,N_12214);
nand U12510 (N_12510,N_12332,N_12063);
nor U12511 (N_12511,N_12316,N_12341);
xor U12512 (N_12512,N_12405,N_12329);
nand U12513 (N_12513,N_12187,N_12198);
xor U12514 (N_12514,N_12114,N_12057);
and U12515 (N_12515,N_12362,N_12056);
nand U12516 (N_12516,N_12267,N_12485);
nor U12517 (N_12517,N_12007,N_12303);
nor U12518 (N_12518,N_12171,N_12149);
nor U12519 (N_12519,N_12399,N_12005);
or U12520 (N_12520,N_12189,N_12447);
and U12521 (N_12521,N_12133,N_12268);
xor U12522 (N_12522,N_12101,N_12213);
nand U12523 (N_12523,N_12358,N_12328);
nor U12524 (N_12524,N_12173,N_12324);
nand U12525 (N_12525,N_12442,N_12391);
nand U12526 (N_12526,N_12378,N_12317);
xnor U12527 (N_12527,N_12028,N_12025);
nand U12528 (N_12528,N_12272,N_12164);
nor U12529 (N_12529,N_12086,N_12053);
or U12530 (N_12530,N_12093,N_12082);
nor U12531 (N_12531,N_12251,N_12104);
nand U12532 (N_12532,N_12241,N_12460);
nand U12533 (N_12533,N_12155,N_12128);
xor U12534 (N_12534,N_12159,N_12481);
or U12535 (N_12535,N_12166,N_12070);
nor U12536 (N_12536,N_12420,N_12042);
xor U12537 (N_12537,N_12323,N_12008);
and U12538 (N_12538,N_12337,N_12386);
and U12539 (N_12539,N_12126,N_12371);
xnor U12540 (N_12540,N_12243,N_12352);
xor U12541 (N_12541,N_12044,N_12023);
nor U12542 (N_12542,N_12080,N_12254);
or U12543 (N_12543,N_12413,N_12219);
or U12544 (N_12544,N_12078,N_12216);
xor U12545 (N_12545,N_12469,N_12453);
xor U12546 (N_12546,N_12474,N_12116);
xnor U12547 (N_12547,N_12348,N_12011);
or U12548 (N_12548,N_12339,N_12201);
nor U12549 (N_12549,N_12476,N_12281);
nor U12550 (N_12550,N_12031,N_12010);
or U12551 (N_12551,N_12369,N_12018);
nor U12552 (N_12552,N_12286,N_12294);
nand U12553 (N_12553,N_12054,N_12437);
or U12554 (N_12554,N_12004,N_12176);
nor U12555 (N_12555,N_12414,N_12084);
and U12556 (N_12556,N_12302,N_12306);
and U12557 (N_12557,N_12145,N_12191);
nor U12558 (N_12558,N_12058,N_12372);
or U12559 (N_12559,N_12088,N_12411);
nand U12560 (N_12560,N_12407,N_12151);
and U12561 (N_12561,N_12257,N_12379);
nand U12562 (N_12562,N_12169,N_12124);
or U12563 (N_12563,N_12202,N_12223);
nor U12564 (N_12564,N_12157,N_12275);
or U12565 (N_12565,N_12478,N_12150);
and U12566 (N_12566,N_12206,N_12247);
xnor U12567 (N_12567,N_12292,N_12490);
or U12568 (N_12568,N_12115,N_12385);
nand U12569 (N_12569,N_12110,N_12220);
and U12570 (N_12570,N_12488,N_12148);
or U12571 (N_12571,N_12419,N_12026);
nand U12572 (N_12572,N_12240,N_12017);
nand U12573 (N_12573,N_12445,N_12459);
and U12574 (N_12574,N_12461,N_12249);
nor U12575 (N_12575,N_12350,N_12246);
xor U12576 (N_12576,N_12119,N_12376);
or U12577 (N_12577,N_12059,N_12092);
and U12578 (N_12578,N_12252,N_12130);
xor U12579 (N_12579,N_12297,N_12489);
and U12580 (N_12580,N_12416,N_12392);
xor U12581 (N_12581,N_12205,N_12129);
nand U12582 (N_12582,N_12417,N_12383);
or U12583 (N_12583,N_12363,N_12178);
or U12584 (N_12584,N_12016,N_12457);
or U12585 (N_12585,N_12398,N_12158);
or U12586 (N_12586,N_12027,N_12153);
xor U12587 (N_12587,N_12134,N_12466);
nor U12588 (N_12588,N_12320,N_12147);
nor U12589 (N_12589,N_12450,N_12432);
nand U12590 (N_12590,N_12499,N_12305);
and U12591 (N_12591,N_12336,N_12470);
nor U12592 (N_12592,N_12259,N_12185);
or U12593 (N_12593,N_12089,N_12498);
nor U12594 (N_12594,N_12067,N_12014);
xor U12595 (N_12595,N_12486,N_12064);
and U12596 (N_12596,N_12353,N_12123);
nor U12597 (N_12597,N_12193,N_12224);
nand U12598 (N_12598,N_12156,N_12163);
xnor U12599 (N_12599,N_12132,N_12448);
or U12600 (N_12600,N_12068,N_12475);
nor U12601 (N_12601,N_12245,N_12109);
nor U12602 (N_12602,N_12037,N_12152);
nand U12603 (N_12603,N_12364,N_12207);
nand U12604 (N_12604,N_12355,N_12282);
or U12605 (N_12605,N_12495,N_12167);
or U12606 (N_12606,N_12406,N_12065);
or U12607 (N_12607,N_12423,N_12440);
and U12608 (N_12608,N_12143,N_12354);
nor U12609 (N_12609,N_12102,N_12368);
nor U12610 (N_12610,N_12100,N_12231);
nand U12611 (N_12611,N_12050,N_12168);
nand U12612 (N_12612,N_12433,N_12052);
and U12613 (N_12613,N_12186,N_12496);
or U12614 (N_12614,N_12390,N_12239);
nor U12615 (N_12615,N_12356,N_12015);
or U12616 (N_12616,N_12188,N_12179);
xor U12617 (N_12617,N_12103,N_12387);
or U12618 (N_12618,N_12060,N_12321);
nand U12619 (N_12619,N_12426,N_12497);
and U12620 (N_12620,N_12233,N_12483);
xnor U12621 (N_12621,N_12409,N_12438);
and U12622 (N_12622,N_12045,N_12375);
xor U12623 (N_12623,N_12118,N_12204);
nor U12624 (N_12624,N_12380,N_12226);
or U12625 (N_12625,N_12435,N_12401);
nand U12626 (N_12626,N_12136,N_12229);
and U12627 (N_12627,N_12261,N_12066);
nor U12628 (N_12628,N_12269,N_12365);
xor U12629 (N_12629,N_12035,N_12107);
or U12630 (N_12630,N_12359,N_12319);
and U12631 (N_12631,N_12002,N_12048);
nor U12632 (N_12632,N_12049,N_12471);
nand U12633 (N_12633,N_12021,N_12311);
nand U12634 (N_12634,N_12403,N_12482);
xnor U12635 (N_12635,N_12034,N_12094);
and U12636 (N_12636,N_12105,N_12422);
nor U12637 (N_12637,N_12075,N_12273);
or U12638 (N_12638,N_12318,N_12451);
or U12639 (N_12639,N_12175,N_12038);
nor U12640 (N_12640,N_12020,N_12444);
or U12641 (N_12641,N_12161,N_12127);
nor U12642 (N_12642,N_12396,N_12217);
nor U12643 (N_12643,N_12349,N_12258);
nor U12644 (N_12644,N_12108,N_12222);
nand U12645 (N_12645,N_12001,N_12266);
xor U12646 (N_12646,N_12394,N_12454);
and U12647 (N_12647,N_12135,N_12287);
or U12648 (N_12648,N_12429,N_12340);
and U12649 (N_12649,N_12019,N_12121);
nand U12650 (N_12650,N_12230,N_12006);
xor U12651 (N_12651,N_12200,N_12036);
nand U12652 (N_12652,N_12291,N_12051);
and U12653 (N_12653,N_12334,N_12047);
nor U12654 (N_12654,N_12446,N_12276);
nor U12655 (N_12655,N_12172,N_12250);
and U12656 (N_12656,N_12467,N_12427);
nand U12657 (N_12657,N_12480,N_12264);
xnor U12658 (N_12658,N_12097,N_12122);
nor U12659 (N_12659,N_12184,N_12039);
nor U12660 (N_12660,N_12477,N_12338);
and U12661 (N_12661,N_12091,N_12484);
nor U12662 (N_12662,N_12096,N_12046);
nor U12663 (N_12663,N_12211,N_12260);
or U12664 (N_12664,N_12237,N_12315);
nand U12665 (N_12665,N_12077,N_12221);
xor U12666 (N_12666,N_12131,N_12043);
and U12667 (N_12667,N_12487,N_12072);
nor U12668 (N_12668,N_12262,N_12288);
xor U12669 (N_12669,N_12165,N_12330);
nor U12670 (N_12670,N_12095,N_12032);
or U12671 (N_12671,N_12234,N_12139);
nand U12672 (N_12672,N_12439,N_12290);
xnor U12673 (N_12673,N_12373,N_12397);
xnor U12674 (N_12674,N_12428,N_12309);
or U12675 (N_12675,N_12099,N_12085);
nand U12676 (N_12676,N_12195,N_12395);
xor U12677 (N_12677,N_12389,N_12455);
nor U12678 (N_12678,N_12284,N_12182);
and U12679 (N_12679,N_12296,N_12029);
or U12680 (N_12680,N_12367,N_12271);
nor U12681 (N_12681,N_12263,N_12479);
and U12682 (N_12682,N_12441,N_12117);
xor U12683 (N_12683,N_12400,N_12415);
nand U12684 (N_12684,N_12069,N_12333);
and U12685 (N_12685,N_12366,N_12443);
nor U12686 (N_12686,N_12270,N_12140);
and U12687 (N_12687,N_12235,N_12310);
and U12688 (N_12688,N_12073,N_12412);
nor U12689 (N_12689,N_12144,N_12346);
nor U12690 (N_12690,N_12449,N_12431);
and U12691 (N_12691,N_12253,N_12344);
and U12692 (N_12692,N_12194,N_12289);
and U12693 (N_12693,N_12347,N_12280);
xnor U12694 (N_12694,N_12055,N_12462);
or U12695 (N_12695,N_12335,N_12351);
nor U12696 (N_12696,N_12377,N_12256);
xnor U12697 (N_12697,N_12081,N_12009);
and U12698 (N_12698,N_12141,N_12197);
nor U12699 (N_12699,N_12232,N_12228);
nand U12700 (N_12700,N_12079,N_12210);
xor U12701 (N_12701,N_12112,N_12307);
and U12702 (N_12702,N_12343,N_12192);
nor U12703 (N_12703,N_12087,N_12125);
or U12704 (N_12704,N_12393,N_12295);
and U12705 (N_12705,N_12293,N_12285);
and U12706 (N_12706,N_12255,N_12283);
xnor U12707 (N_12707,N_12196,N_12030);
xnor U12708 (N_12708,N_12304,N_12434);
nor U12709 (N_12709,N_12090,N_12418);
nor U12710 (N_12710,N_12248,N_12003);
nor U12711 (N_12711,N_12402,N_12410);
nor U12712 (N_12712,N_12076,N_12242);
and U12713 (N_12713,N_12098,N_12074);
and U12714 (N_12714,N_12384,N_12357);
nor U12715 (N_12715,N_12013,N_12374);
nor U12716 (N_12716,N_12062,N_12382);
or U12717 (N_12717,N_12138,N_12492);
xor U12718 (N_12718,N_12061,N_12452);
and U12719 (N_12719,N_12238,N_12177);
or U12720 (N_12720,N_12199,N_12180);
xor U12721 (N_12721,N_12274,N_12463);
and U12722 (N_12722,N_12430,N_12381);
nor U12723 (N_12723,N_12024,N_12388);
and U12724 (N_12724,N_12456,N_12360);
nand U12725 (N_12725,N_12465,N_12278);
nor U12726 (N_12726,N_12142,N_12345);
xnor U12727 (N_12727,N_12227,N_12083);
and U12728 (N_12728,N_12493,N_12183);
nand U12729 (N_12729,N_12342,N_12236);
xnor U12730 (N_12730,N_12000,N_12215);
xnor U12731 (N_12731,N_12162,N_12468);
nor U12732 (N_12732,N_12370,N_12154);
and U12733 (N_12733,N_12408,N_12494);
or U12734 (N_12734,N_12308,N_12137);
nor U12735 (N_12735,N_12424,N_12218);
or U12736 (N_12736,N_12174,N_12361);
and U12737 (N_12737,N_12300,N_12421);
nor U12738 (N_12738,N_12458,N_12436);
and U12739 (N_12739,N_12322,N_12425);
or U12740 (N_12740,N_12208,N_12212);
nor U12741 (N_12741,N_12314,N_12170);
xnor U12742 (N_12742,N_12181,N_12472);
xor U12743 (N_12743,N_12120,N_12012);
xor U12744 (N_12744,N_12209,N_12203);
and U12745 (N_12745,N_12277,N_12473);
and U12746 (N_12746,N_12113,N_12071);
or U12747 (N_12747,N_12190,N_12327);
xnor U12748 (N_12748,N_12022,N_12325);
nand U12749 (N_12749,N_12279,N_12312);
nand U12750 (N_12750,N_12178,N_12287);
nor U12751 (N_12751,N_12301,N_12156);
nand U12752 (N_12752,N_12432,N_12043);
nand U12753 (N_12753,N_12250,N_12169);
or U12754 (N_12754,N_12010,N_12049);
and U12755 (N_12755,N_12462,N_12179);
xnor U12756 (N_12756,N_12186,N_12398);
nand U12757 (N_12757,N_12124,N_12313);
and U12758 (N_12758,N_12446,N_12148);
xnor U12759 (N_12759,N_12244,N_12181);
xor U12760 (N_12760,N_12275,N_12153);
nand U12761 (N_12761,N_12136,N_12029);
or U12762 (N_12762,N_12130,N_12131);
or U12763 (N_12763,N_12185,N_12444);
and U12764 (N_12764,N_12271,N_12172);
xor U12765 (N_12765,N_12224,N_12333);
or U12766 (N_12766,N_12336,N_12300);
or U12767 (N_12767,N_12193,N_12365);
or U12768 (N_12768,N_12330,N_12255);
or U12769 (N_12769,N_12458,N_12023);
xnor U12770 (N_12770,N_12307,N_12061);
and U12771 (N_12771,N_12188,N_12468);
nor U12772 (N_12772,N_12257,N_12119);
or U12773 (N_12773,N_12322,N_12361);
xor U12774 (N_12774,N_12183,N_12406);
xnor U12775 (N_12775,N_12459,N_12484);
or U12776 (N_12776,N_12351,N_12129);
nand U12777 (N_12777,N_12483,N_12390);
xnor U12778 (N_12778,N_12399,N_12485);
nor U12779 (N_12779,N_12269,N_12143);
xor U12780 (N_12780,N_12026,N_12009);
or U12781 (N_12781,N_12190,N_12098);
or U12782 (N_12782,N_12001,N_12026);
nor U12783 (N_12783,N_12125,N_12038);
and U12784 (N_12784,N_12499,N_12250);
xor U12785 (N_12785,N_12388,N_12429);
xor U12786 (N_12786,N_12399,N_12291);
nor U12787 (N_12787,N_12398,N_12227);
xor U12788 (N_12788,N_12477,N_12391);
nor U12789 (N_12789,N_12072,N_12085);
nor U12790 (N_12790,N_12029,N_12025);
nor U12791 (N_12791,N_12384,N_12040);
or U12792 (N_12792,N_12119,N_12450);
xor U12793 (N_12793,N_12162,N_12370);
xor U12794 (N_12794,N_12186,N_12017);
or U12795 (N_12795,N_12279,N_12429);
nor U12796 (N_12796,N_12130,N_12201);
nand U12797 (N_12797,N_12137,N_12145);
nand U12798 (N_12798,N_12359,N_12285);
nand U12799 (N_12799,N_12033,N_12095);
nand U12800 (N_12800,N_12221,N_12065);
nand U12801 (N_12801,N_12335,N_12338);
or U12802 (N_12802,N_12274,N_12469);
nor U12803 (N_12803,N_12226,N_12334);
nor U12804 (N_12804,N_12403,N_12417);
xnor U12805 (N_12805,N_12095,N_12276);
or U12806 (N_12806,N_12319,N_12386);
nand U12807 (N_12807,N_12334,N_12183);
xor U12808 (N_12808,N_12015,N_12157);
or U12809 (N_12809,N_12014,N_12050);
and U12810 (N_12810,N_12361,N_12041);
nand U12811 (N_12811,N_12289,N_12074);
nand U12812 (N_12812,N_12486,N_12282);
or U12813 (N_12813,N_12290,N_12260);
xnor U12814 (N_12814,N_12053,N_12441);
xnor U12815 (N_12815,N_12342,N_12119);
nor U12816 (N_12816,N_12182,N_12055);
nor U12817 (N_12817,N_12246,N_12336);
and U12818 (N_12818,N_12226,N_12113);
nand U12819 (N_12819,N_12432,N_12333);
nor U12820 (N_12820,N_12238,N_12265);
nor U12821 (N_12821,N_12105,N_12210);
or U12822 (N_12822,N_12366,N_12062);
and U12823 (N_12823,N_12005,N_12360);
nand U12824 (N_12824,N_12110,N_12089);
and U12825 (N_12825,N_12336,N_12456);
xor U12826 (N_12826,N_12249,N_12430);
nor U12827 (N_12827,N_12146,N_12004);
nor U12828 (N_12828,N_12053,N_12322);
nor U12829 (N_12829,N_12003,N_12076);
nor U12830 (N_12830,N_12034,N_12147);
and U12831 (N_12831,N_12223,N_12198);
xnor U12832 (N_12832,N_12499,N_12330);
and U12833 (N_12833,N_12027,N_12015);
and U12834 (N_12834,N_12051,N_12288);
nor U12835 (N_12835,N_12072,N_12228);
or U12836 (N_12836,N_12472,N_12086);
xnor U12837 (N_12837,N_12390,N_12075);
and U12838 (N_12838,N_12290,N_12066);
or U12839 (N_12839,N_12061,N_12036);
xnor U12840 (N_12840,N_12367,N_12254);
nand U12841 (N_12841,N_12107,N_12180);
and U12842 (N_12842,N_12449,N_12162);
and U12843 (N_12843,N_12132,N_12295);
or U12844 (N_12844,N_12045,N_12329);
xnor U12845 (N_12845,N_12351,N_12032);
or U12846 (N_12846,N_12003,N_12106);
xor U12847 (N_12847,N_12058,N_12431);
nor U12848 (N_12848,N_12377,N_12458);
nor U12849 (N_12849,N_12286,N_12249);
nor U12850 (N_12850,N_12296,N_12462);
nand U12851 (N_12851,N_12371,N_12032);
nand U12852 (N_12852,N_12238,N_12199);
nor U12853 (N_12853,N_12074,N_12272);
xnor U12854 (N_12854,N_12074,N_12377);
nor U12855 (N_12855,N_12420,N_12339);
and U12856 (N_12856,N_12463,N_12392);
and U12857 (N_12857,N_12086,N_12330);
and U12858 (N_12858,N_12203,N_12096);
or U12859 (N_12859,N_12471,N_12063);
nor U12860 (N_12860,N_12208,N_12240);
or U12861 (N_12861,N_12140,N_12039);
or U12862 (N_12862,N_12104,N_12482);
nand U12863 (N_12863,N_12161,N_12295);
nand U12864 (N_12864,N_12262,N_12287);
nand U12865 (N_12865,N_12025,N_12163);
or U12866 (N_12866,N_12104,N_12391);
and U12867 (N_12867,N_12029,N_12153);
nand U12868 (N_12868,N_12300,N_12230);
nor U12869 (N_12869,N_12183,N_12049);
nor U12870 (N_12870,N_12050,N_12249);
nor U12871 (N_12871,N_12081,N_12251);
nor U12872 (N_12872,N_12117,N_12060);
or U12873 (N_12873,N_12473,N_12492);
nor U12874 (N_12874,N_12225,N_12257);
or U12875 (N_12875,N_12222,N_12100);
nand U12876 (N_12876,N_12119,N_12386);
nand U12877 (N_12877,N_12167,N_12273);
nor U12878 (N_12878,N_12328,N_12045);
or U12879 (N_12879,N_12019,N_12484);
xor U12880 (N_12880,N_12322,N_12057);
xor U12881 (N_12881,N_12205,N_12056);
xor U12882 (N_12882,N_12162,N_12367);
or U12883 (N_12883,N_12264,N_12128);
xor U12884 (N_12884,N_12386,N_12070);
nor U12885 (N_12885,N_12201,N_12118);
and U12886 (N_12886,N_12442,N_12129);
xor U12887 (N_12887,N_12240,N_12170);
and U12888 (N_12888,N_12176,N_12301);
and U12889 (N_12889,N_12295,N_12163);
or U12890 (N_12890,N_12030,N_12009);
xor U12891 (N_12891,N_12426,N_12105);
nor U12892 (N_12892,N_12204,N_12179);
and U12893 (N_12893,N_12136,N_12460);
xor U12894 (N_12894,N_12197,N_12041);
or U12895 (N_12895,N_12494,N_12008);
or U12896 (N_12896,N_12351,N_12026);
xor U12897 (N_12897,N_12423,N_12273);
xnor U12898 (N_12898,N_12498,N_12038);
or U12899 (N_12899,N_12183,N_12310);
or U12900 (N_12900,N_12050,N_12364);
or U12901 (N_12901,N_12255,N_12012);
and U12902 (N_12902,N_12000,N_12260);
or U12903 (N_12903,N_12024,N_12308);
or U12904 (N_12904,N_12191,N_12458);
nand U12905 (N_12905,N_12278,N_12466);
nor U12906 (N_12906,N_12192,N_12332);
xnor U12907 (N_12907,N_12398,N_12238);
nand U12908 (N_12908,N_12046,N_12257);
xor U12909 (N_12909,N_12362,N_12475);
nand U12910 (N_12910,N_12194,N_12465);
nor U12911 (N_12911,N_12164,N_12222);
nor U12912 (N_12912,N_12086,N_12328);
and U12913 (N_12913,N_12264,N_12010);
xnor U12914 (N_12914,N_12015,N_12213);
nand U12915 (N_12915,N_12408,N_12376);
and U12916 (N_12916,N_12052,N_12227);
or U12917 (N_12917,N_12003,N_12072);
and U12918 (N_12918,N_12273,N_12105);
or U12919 (N_12919,N_12213,N_12106);
and U12920 (N_12920,N_12282,N_12350);
and U12921 (N_12921,N_12485,N_12396);
or U12922 (N_12922,N_12384,N_12174);
xnor U12923 (N_12923,N_12377,N_12033);
xor U12924 (N_12924,N_12027,N_12187);
xnor U12925 (N_12925,N_12086,N_12110);
nor U12926 (N_12926,N_12161,N_12303);
nor U12927 (N_12927,N_12361,N_12387);
or U12928 (N_12928,N_12261,N_12236);
and U12929 (N_12929,N_12333,N_12455);
nor U12930 (N_12930,N_12166,N_12442);
and U12931 (N_12931,N_12430,N_12134);
xor U12932 (N_12932,N_12215,N_12081);
xnor U12933 (N_12933,N_12071,N_12186);
and U12934 (N_12934,N_12159,N_12221);
or U12935 (N_12935,N_12022,N_12191);
and U12936 (N_12936,N_12465,N_12250);
and U12937 (N_12937,N_12396,N_12251);
nor U12938 (N_12938,N_12479,N_12107);
or U12939 (N_12939,N_12399,N_12117);
xor U12940 (N_12940,N_12013,N_12297);
and U12941 (N_12941,N_12486,N_12226);
or U12942 (N_12942,N_12349,N_12300);
nor U12943 (N_12943,N_12472,N_12386);
or U12944 (N_12944,N_12496,N_12347);
nor U12945 (N_12945,N_12328,N_12442);
and U12946 (N_12946,N_12037,N_12276);
nor U12947 (N_12947,N_12149,N_12151);
or U12948 (N_12948,N_12240,N_12361);
xnor U12949 (N_12949,N_12477,N_12316);
nand U12950 (N_12950,N_12343,N_12199);
xor U12951 (N_12951,N_12260,N_12456);
xnor U12952 (N_12952,N_12280,N_12307);
nor U12953 (N_12953,N_12219,N_12303);
and U12954 (N_12954,N_12468,N_12353);
nand U12955 (N_12955,N_12202,N_12250);
or U12956 (N_12956,N_12077,N_12074);
nor U12957 (N_12957,N_12153,N_12249);
nor U12958 (N_12958,N_12046,N_12181);
nand U12959 (N_12959,N_12466,N_12219);
or U12960 (N_12960,N_12136,N_12022);
or U12961 (N_12961,N_12081,N_12086);
nand U12962 (N_12962,N_12137,N_12003);
and U12963 (N_12963,N_12438,N_12453);
nor U12964 (N_12964,N_12263,N_12149);
nor U12965 (N_12965,N_12291,N_12375);
and U12966 (N_12966,N_12154,N_12070);
nand U12967 (N_12967,N_12050,N_12137);
and U12968 (N_12968,N_12429,N_12012);
nand U12969 (N_12969,N_12332,N_12111);
nand U12970 (N_12970,N_12335,N_12475);
nor U12971 (N_12971,N_12007,N_12338);
or U12972 (N_12972,N_12147,N_12216);
xnor U12973 (N_12973,N_12269,N_12408);
and U12974 (N_12974,N_12044,N_12147);
xor U12975 (N_12975,N_12011,N_12104);
xnor U12976 (N_12976,N_12231,N_12060);
or U12977 (N_12977,N_12120,N_12308);
or U12978 (N_12978,N_12184,N_12219);
and U12979 (N_12979,N_12018,N_12170);
and U12980 (N_12980,N_12265,N_12391);
and U12981 (N_12981,N_12448,N_12242);
nand U12982 (N_12982,N_12075,N_12001);
or U12983 (N_12983,N_12148,N_12112);
and U12984 (N_12984,N_12000,N_12033);
and U12985 (N_12985,N_12298,N_12182);
nor U12986 (N_12986,N_12318,N_12045);
and U12987 (N_12987,N_12409,N_12188);
nor U12988 (N_12988,N_12252,N_12414);
xor U12989 (N_12989,N_12230,N_12209);
xor U12990 (N_12990,N_12430,N_12494);
nand U12991 (N_12991,N_12096,N_12231);
and U12992 (N_12992,N_12195,N_12427);
xor U12993 (N_12993,N_12322,N_12278);
xnor U12994 (N_12994,N_12196,N_12305);
and U12995 (N_12995,N_12234,N_12408);
nand U12996 (N_12996,N_12131,N_12085);
nand U12997 (N_12997,N_12189,N_12483);
xor U12998 (N_12998,N_12237,N_12105);
nand U12999 (N_12999,N_12105,N_12099);
and U13000 (N_13000,N_12512,N_12530);
nand U13001 (N_13001,N_12527,N_12801);
xnor U13002 (N_13002,N_12905,N_12723);
or U13003 (N_13003,N_12847,N_12733);
or U13004 (N_13004,N_12615,N_12743);
nand U13005 (N_13005,N_12885,N_12648);
xnor U13006 (N_13006,N_12651,N_12892);
nand U13007 (N_13007,N_12533,N_12815);
or U13008 (N_13008,N_12622,N_12903);
nand U13009 (N_13009,N_12915,N_12653);
or U13010 (N_13010,N_12861,N_12797);
nand U13011 (N_13011,N_12528,N_12577);
nand U13012 (N_13012,N_12501,N_12570);
nor U13013 (N_13013,N_12734,N_12770);
and U13014 (N_13014,N_12882,N_12529);
or U13015 (N_13015,N_12649,N_12846);
nand U13016 (N_13016,N_12509,N_12521);
xnor U13017 (N_13017,N_12507,N_12991);
nand U13018 (N_13018,N_12865,N_12640);
nand U13019 (N_13019,N_12854,N_12912);
and U13020 (N_13020,N_12650,N_12902);
nand U13021 (N_13021,N_12544,N_12920);
or U13022 (N_13022,N_12736,N_12704);
nor U13023 (N_13023,N_12838,N_12523);
xnor U13024 (N_13024,N_12886,N_12941);
xnor U13025 (N_13025,N_12567,N_12519);
nor U13026 (N_13026,N_12756,N_12878);
nand U13027 (N_13027,N_12895,N_12959);
and U13028 (N_13028,N_12939,N_12759);
or U13029 (N_13029,N_12718,N_12952);
or U13030 (N_13030,N_12515,N_12594);
and U13031 (N_13031,N_12784,N_12859);
xor U13032 (N_13032,N_12742,N_12809);
or U13033 (N_13033,N_12836,N_12860);
nor U13034 (N_13034,N_12684,N_12681);
xnor U13035 (N_13035,N_12857,N_12837);
nor U13036 (N_13036,N_12822,N_12774);
nor U13037 (N_13037,N_12776,N_12739);
nand U13038 (N_13038,N_12889,N_12936);
xnor U13039 (N_13039,N_12973,N_12741);
or U13040 (N_13040,N_12754,N_12906);
nor U13041 (N_13041,N_12735,N_12678);
and U13042 (N_13042,N_12564,N_12757);
nand U13043 (N_13043,N_12999,N_12506);
nor U13044 (N_13044,N_12767,N_12639);
nand U13045 (N_13045,N_12726,N_12660);
xor U13046 (N_13046,N_12720,N_12599);
and U13047 (N_13047,N_12568,N_12748);
nor U13048 (N_13048,N_12508,N_12549);
or U13049 (N_13049,N_12730,N_12777);
nand U13050 (N_13050,N_12738,N_12984);
or U13051 (N_13051,N_12938,N_12995);
nor U13052 (N_13052,N_12922,N_12644);
nand U13053 (N_13053,N_12612,N_12888);
or U13054 (N_13054,N_12950,N_12727);
xor U13055 (N_13055,N_12522,N_12542);
xnor U13056 (N_13056,N_12782,N_12595);
and U13057 (N_13057,N_12524,N_12719);
or U13058 (N_13058,N_12832,N_12873);
and U13059 (N_13059,N_12546,N_12694);
nand U13060 (N_13060,N_12755,N_12691);
nand U13061 (N_13061,N_12940,N_12834);
nor U13062 (N_13062,N_12732,N_12722);
or U13063 (N_13063,N_12751,N_12526);
or U13064 (N_13064,N_12747,N_12662);
xnor U13065 (N_13065,N_12552,N_12687);
and U13066 (N_13066,N_12977,N_12740);
and U13067 (N_13067,N_12870,N_12908);
nor U13068 (N_13068,N_12541,N_12932);
or U13069 (N_13069,N_12605,N_12538);
nand U13070 (N_13070,N_12948,N_12803);
nand U13071 (N_13071,N_12824,N_12717);
and U13072 (N_13072,N_12769,N_12657);
or U13073 (N_13073,N_12842,N_12583);
or U13074 (N_13074,N_12545,N_12514);
nor U13075 (N_13075,N_12814,N_12548);
xnor U13076 (N_13076,N_12928,N_12630);
xnor U13077 (N_13077,N_12980,N_12525);
nor U13078 (N_13078,N_12680,N_12661);
nand U13079 (N_13079,N_12919,N_12947);
or U13080 (N_13080,N_12635,N_12632);
nand U13081 (N_13081,N_12619,N_12983);
or U13082 (N_13082,N_12560,N_12550);
and U13083 (N_13083,N_12758,N_12633);
nand U13084 (N_13084,N_12986,N_12974);
and U13085 (N_13085,N_12703,N_12578);
and U13086 (N_13086,N_12996,N_12580);
or U13087 (N_13087,N_12790,N_12646);
nor U13088 (N_13088,N_12763,N_12998);
and U13089 (N_13089,N_12729,N_12698);
nor U13090 (N_13090,N_12926,N_12909);
or U13091 (N_13091,N_12916,N_12693);
nand U13092 (N_13092,N_12685,N_12798);
and U13093 (N_13093,N_12600,N_12596);
nand U13094 (N_13094,N_12831,N_12667);
xor U13095 (N_13095,N_12768,N_12606);
or U13096 (N_13096,N_12848,N_12749);
or U13097 (N_13097,N_12610,N_12985);
nand U13098 (N_13098,N_12967,N_12711);
nor U13099 (N_13099,N_12816,N_12634);
nand U13100 (N_13100,N_12800,N_12968);
nor U13101 (N_13101,N_12989,N_12877);
nor U13102 (N_13102,N_12654,N_12638);
nor U13103 (N_13103,N_12818,N_12593);
and U13104 (N_13104,N_12602,N_12607);
nor U13105 (N_13105,N_12827,N_12937);
or U13106 (N_13106,N_12591,N_12871);
nand U13107 (N_13107,N_12825,N_12569);
and U13108 (N_13108,N_12713,N_12665);
or U13109 (N_13109,N_12572,N_12976);
or U13110 (N_13110,N_12943,N_12918);
and U13111 (N_13111,N_12561,N_12960);
or U13112 (N_13112,N_12812,N_12586);
and U13113 (N_13113,N_12565,N_12817);
xnor U13114 (N_13114,N_12688,N_12673);
or U13115 (N_13115,N_12752,N_12536);
nand U13116 (N_13116,N_12867,N_12917);
or U13117 (N_13117,N_12504,N_12677);
nor U13118 (N_13118,N_12540,N_12592);
xnor U13119 (N_13119,N_12647,N_12978);
nor U13120 (N_13120,N_12828,N_12700);
or U13121 (N_13121,N_12645,N_12510);
nor U13122 (N_13122,N_12579,N_12780);
and U13123 (N_13123,N_12898,N_12566);
and U13124 (N_13124,N_12598,N_12597);
nand U13125 (N_13125,N_12773,N_12551);
nand U13126 (N_13126,N_12601,N_12821);
and U13127 (N_13127,N_12608,N_12901);
xor U13128 (N_13128,N_12502,N_12604);
and U13129 (N_13129,N_12574,N_12788);
xor U13130 (N_13130,N_12844,N_12781);
nand U13131 (N_13131,N_12744,N_12624);
xor U13132 (N_13132,N_12964,N_12672);
nand U13133 (N_13133,N_12875,N_12789);
xnor U13134 (N_13134,N_12914,N_12563);
or U13135 (N_13135,N_12576,N_12637);
and U13136 (N_13136,N_12804,N_12879);
and U13137 (N_13137,N_12858,N_12791);
or U13138 (N_13138,N_12783,N_12558);
xor U13139 (N_13139,N_12956,N_12584);
and U13140 (N_13140,N_12930,N_12787);
nand U13141 (N_13141,N_12571,N_12575);
nor U13142 (N_13142,N_12849,N_12924);
nand U13143 (N_13143,N_12775,N_12850);
xnor U13144 (N_13144,N_12955,N_12874);
xor U13145 (N_13145,N_12951,N_12934);
xor U13146 (N_13146,N_12664,N_12620);
xnor U13147 (N_13147,N_12946,N_12535);
and U13148 (N_13148,N_12621,N_12636);
or U13149 (N_13149,N_12534,N_12690);
xor U13150 (N_13150,N_12628,N_12792);
nor U13151 (N_13151,N_12587,N_12988);
and U13152 (N_13152,N_12962,N_12537);
nor U13153 (N_13153,N_12613,N_12933);
nor U13154 (N_13154,N_12931,N_12965);
and U13155 (N_13155,N_12675,N_12786);
or U13156 (N_13156,N_12585,N_12893);
and U13157 (N_13157,N_12705,N_12881);
or U13158 (N_13158,N_12866,N_12811);
xnor U13159 (N_13159,N_12670,N_12794);
and U13160 (N_13160,N_12975,N_12655);
or U13161 (N_13161,N_12923,N_12972);
or U13162 (N_13162,N_12686,N_12806);
or U13163 (N_13163,N_12554,N_12531);
nor U13164 (N_13164,N_12511,N_12958);
nand U13165 (N_13165,N_12863,N_12696);
and U13166 (N_13166,N_12808,N_12671);
nand U13167 (N_13167,N_12716,N_12682);
or U13168 (N_13168,N_12813,N_12785);
or U13169 (N_13169,N_12699,N_12795);
nand U13170 (N_13170,N_12880,N_12910);
nand U13171 (N_13171,N_12872,N_12625);
xor U13172 (N_13172,N_12907,N_12894);
and U13173 (N_13173,N_12969,N_12589);
xnor U13174 (N_13174,N_12807,N_12949);
or U13175 (N_13175,N_12760,N_12710);
nor U13176 (N_13176,N_12652,N_12899);
nand U13177 (N_13177,N_12862,N_12614);
nor U13178 (N_13178,N_12845,N_12942);
xor U13179 (N_13179,N_12982,N_12555);
nand U13180 (N_13180,N_12981,N_12643);
nand U13181 (N_13181,N_12796,N_12714);
nor U13182 (N_13182,N_12518,N_12689);
xnor U13183 (N_13183,N_12520,N_12841);
and U13184 (N_13184,N_12853,N_12627);
xnor U13185 (N_13185,N_12971,N_12603);
xnor U13186 (N_13186,N_12961,N_12500);
xor U13187 (N_13187,N_12623,N_12724);
and U13188 (N_13188,N_12897,N_12992);
xnor U13189 (N_13189,N_12945,N_12750);
or U13190 (N_13190,N_12876,N_12656);
and U13191 (N_13191,N_12547,N_12793);
and U13192 (N_13192,N_12641,N_12935);
or U13193 (N_13193,N_12753,N_12674);
nand U13194 (N_13194,N_12663,N_12505);
or U13195 (N_13195,N_12799,N_12771);
nand U13196 (N_13196,N_12927,N_12820);
xnor U13197 (N_13197,N_12884,N_12868);
nor U13198 (N_13198,N_12779,N_12702);
and U13199 (N_13199,N_12679,N_12855);
nand U13200 (N_13200,N_12666,N_12557);
nand U13201 (N_13201,N_12839,N_12835);
nand U13202 (N_13202,N_12826,N_12890);
and U13203 (N_13203,N_12891,N_12668);
and U13204 (N_13204,N_12994,N_12517);
and U13205 (N_13205,N_12658,N_12588);
xnor U13206 (N_13206,N_12728,N_12532);
nor U13207 (N_13207,N_12772,N_12997);
nor U13208 (N_13208,N_12581,N_12851);
xnor U13209 (N_13209,N_12856,N_12631);
nor U13210 (N_13210,N_12833,N_12712);
nand U13211 (N_13211,N_12852,N_12590);
and U13212 (N_13212,N_12921,N_12708);
and U13213 (N_13213,N_12829,N_12778);
and U13214 (N_13214,N_12611,N_12539);
xor U13215 (N_13215,N_12629,N_12954);
and U13216 (N_13216,N_12911,N_12830);
nand U13217 (N_13217,N_12761,N_12626);
or U13218 (N_13218,N_12745,N_12503);
xor U13219 (N_13219,N_12766,N_12573);
nand U13220 (N_13220,N_12559,N_12582);
and U13221 (N_13221,N_12805,N_12706);
nand U13222 (N_13222,N_12616,N_12957);
xor U13223 (N_13223,N_12887,N_12709);
nor U13224 (N_13224,N_12707,N_12823);
and U13225 (N_13225,N_12543,N_12553);
or U13226 (N_13226,N_12864,N_12683);
nand U13227 (N_13227,N_12843,N_12609);
nand U13228 (N_13228,N_12966,N_12659);
xor U13229 (N_13229,N_12944,N_12642);
xor U13230 (N_13230,N_12990,N_12764);
nor U13231 (N_13231,N_12721,N_12715);
xor U13232 (N_13232,N_12765,N_12993);
and U13233 (N_13233,N_12669,N_12701);
nand U13234 (N_13234,N_12676,N_12697);
xor U13235 (N_13235,N_12925,N_12617);
nor U13236 (N_13236,N_12970,N_12725);
or U13237 (N_13237,N_12762,N_12896);
and U13238 (N_13238,N_12900,N_12929);
xnor U13239 (N_13239,N_12516,N_12987);
and U13240 (N_13240,N_12802,N_12746);
nand U13241 (N_13241,N_12953,N_12562);
or U13242 (N_13242,N_12840,N_12692);
or U13243 (N_13243,N_12810,N_12513);
nor U13244 (N_13244,N_12695,N_12819);
or U13245 (N_13245,N_12556,N_12618);
or U13246 (N_13246,N_12963,N_12883);
xor U13247 (N_13247,N_12904,N_12913);
nor U13248 (N_13248,N_12979,N_12731);
and U13249 (N_13249,N_12737,N_12869);
nand U13250 (N_13250,N_12877,N_12654);
or U13251 (N_13251,N_12855,N_12516);
and U13252 (N_13252,N_12518,N_12737);
xnor U13253 (N_13253,N_12975,N_12710);
xnor U13254 (N_13254,N_12687,N_12926);
nor U13255 (N_13255,N_12520,N_12720);
nor U13256 (N_13256,N_12931,N_12650);
nand U13257 (N_13257,N_12945,N_12822);
and U13258 (N_13258,N_12986,N_12509);
nor U13259 (N_13259,N_12929,N_12626);
nor U13260 (N_13260,N_12782,N_12655);
nor U13261 (N_13261,N_12992,N_12528);
xor U13262 (N_13262,N_12659,N_12894);
nor U13263 (N_13263,N_12930,N_12564);
xor U13264 (N_13264,N_12537,N_12771);
xnor U13265 (N_13265,N_12578,N_12939);
nor U13266 (N_13266,N_12659,N_12941);
or U13267 (N_13267,N_12781,N_12613);
xnor U13268 (N_13268,N_12810,N_12683);
or U13269 (N_13269,N_12918,N_12873);
and U13270 (N_13270,N_12921,N_12744);
nor U13271 (N_13271,N_12975,N_12962);
or U13272 (N_13272,N_12714,N_12664);
and U13273 (N_13273,N_12974,N_12952);
nand U13274 (N_13274,N_12763,N_12795);
nand U13275 (N_13275,N_12579,N_12531);
nor U13276 (N_13276,N_12799,N_12649);
and U13277 (N_13277,N_12915,N_12830);
xnor U13278 (N_13278,N_12833,N_12779);
xnor U13279 (N_13279,N_12559,N_12827);
xnor U13280 (N_13280,N_12656,N_12696);
or U13281 (N_13281,N_12733,N_12775);
or U13282 (N_13282,N_12515,N_12539);
xor U13283 (N_13283,N_12838,N_12692);
nor U13284 (N_13284,N_12791,N_12705);
and U13285 (N_13285,N_12773,N_12811);
nand U13286 (N_13286,N_12914,N_12684);
nor U13287 (N_13287,N_12944,N_12558);
or U13288 (N_13288,N_12906,N_12762);
nor U13289 (N_13289,N_12913,N_12578);
xnor U13290 (N_13290,N_12917,N_12638);
and U13291 (N_13291,N_12982,N_12540);
nand U13292 (N_13292,N_12906,N_12764);
and U13293 (N_13293,N_12878,N_12512);
or U13294 (N_13294,N_12567,N_12778);
or U13295 (N_13295,N_12801,N_12830);
nor U13296 (N_13296,N_12594,N_12909);
nor U13297 (N_13297,N_12701,N_12562);
nor U13298 (N_13298,N_12846,N_12917);
and U13299 (N_13299,N_12670,N_12680);
nor U13300 (N_13300,N_12711,N_12752);
nand U13301 (N_13301,N_12500,N_12904);
nand U13302 (N_13302,N_12755,N_12928);
and U13303 (N_13303,N_12669,N_12929);
xor U13304 (N_13304,N_12943,N_12710);
nor U13305 (N_13305,N_12670,N_12761);
or U13306 (N_13306,N_12517,N_12791);
xnor U13307 (N_13307,N_12818,N_12555);
nor U13308 (N_13308,N_12925,N_12812);
nand U13309 (N_13309,N_12678,N_12882);
or U13310 (N_13310,N_12876,N_12556);
xor U13311 (N_13311,N_12573,N_12758);
nor U13312 (N_13312,N_12585,N_12593);
nand U13313 (N_13313,N_12839,N_12648);
or U13314 (N_13314,N_12521,N_12678);
or U13315 (N_13315,N_12514,N_12978);
nand U13316 (N_13316,N_12867,N_12625);
nand U13317 (N_13317,N_12725,N_12578);
or U13318 (N_13318,N_12546,N_12879);
nor U13319 (N_13319,N_12558,N_12860);
nand U13320 (N_13320,N_12886,N_12956);
or U13321 (N_13321,N_12791,N_12586);
xnor U13322 (N_13322,N_12857,N_12826);
nor U13323 (N_13323,N_12668,N_12989);
or U13324 (N_13324,N_12524,N_12943);
nor U13325 (N_13325,N_12700,N_12613);
nor U13326 (N_13326,N_12787,N_12613);
xnor U13327 (N_13327,N_12569,N_12694);
and U13328 (N_13328,N_12729,N_12803);
or U13329 (N_13329,N_12673,N_12647);
nor U13330 (N_13330,N_12660,N_12966);
nor U13331 (N_13331,N_12833,N_12709);
xor U13332 (N_13332,N_12833,N_12759);
nand U13333 (N_13333,N_12686,N_12521);
xnor U13334 (N_13334,N_12958,N_12593);
nor U13335 (N_13335,N_12829,N_12773);
or U13336 (N_13336,N_12509,N_12656);
nor U13337 (N_13337,N_12796,N_12616);
and U13338 (N_13338,N_12890,N_12642);
xor U13339 (N_13339,N_12790,N_12932);
nand U13340 (N_13340,N_12524,N_12802);
or U13341 (N_13341,N_12674,N_12775);
nand U13342 (N_13342,N_12764,N_12530);
xnor U13343 (N_13343,N_12672,N_12678);
xor U13344 (N_13344,N_12691,N_12742);
xor U13345 (N_13345,N_12779,N_12805);
nor U13346 (N_13346,N_12847,N_12786);
nor U13347 (N_13347,N_12953,N_12763);
nor U13348 (N_13348,N_12536,N_12707);
nor U13349 (N_13349,N_12808,N_12537);
nand U13350 (N_13350,N_12695,N_12697);
and U13351 (N_13351,N_12565,N_12624);
xor U13352 (N_13352,N_12635,N_12744);
nor U13353 (N_13353,N_12944,N_12661);
or U13354 (N_13354,N_12647,N_12744);
nand U13355 (N_13355,N_12802,N_12844);
nor U13356 (N_13356,N_12837,N_12724);
nor U13357 (N_13357,N_12933,N_12622);
nor U13358 (N_13358,N_12762,N_12863);
nor U13359 (N_13359,N_12679,N_12963);
nor U13360 (N_13360,N_12694,N_12679);
nor U13361 (N_13361,N_12727,N_12794);
nand U13362 (N_13362,N_12914,N_12568);
or U13363 (N_13363,N_12932,N_12780);
xor U13364 (N_13364,N_12622,N_12783);
nor U13365 (N_13365,N_12868,N_12572);
or U13366 (N_13366,N_12515,N_12534);
nand U13367 (N_13367,N_12950,N_12615);
and U13368 (N_13368,N_12535,N_12585);
and U13369 (N_13369,N_12586,N_12632);
xnor U13370 (N_13370,N_12784,N_12778);
nand U13371 (N_13371,N_12688,N_12641);
xor U13372 (N_13372,N_12819,N_12823);
xor U13373 (N_13373,N_12611,N_12689);
xor U13374 (N_13374,N_12897,N_12880);
and U13375 (N_13375,N_12568,N_12570);
or U13376 (N_13376,N_12652,N_12518);
and U13377 (N_13377,N_12600,N_12940);
or U13378 (N_13378,N_12755,N_12987);
nor U13379 (N_13379,N_12999,N_12565);
nor U13380 (N_13380,N_12701,N_12777);
or U13381 (N_13381,N_12604,N_12792);
nor U13382 (N_13382,N_12923,N_12567);
xnor U13383 (N_13383,N_12985,N_12968);
nand U13384 (N_13384,N_12999,N_12912);
nand U13385 (N_13385,N_12556,N_12594);
nand U13386 (N_13386,N_12978,N_12822);
or U13387 (N_13387,N_12562,N_12501);
xor U13388 (N_13388,N_12756,N_12929);
nand U13389 (N_13389,N_12828,N_12660);
nor U13390 (N_13390,N_12753,N_12721);
and U13391 (N_13391,N_12841,N_12773);
or U13392 (N_13392,N_12579,N_12596);
and U13393 (N_13393,N_12642,N_12722);
nor U13394 (N_13394,N_12608,N_12869);
and U13395 (N_13395,N_12857,N_12718);
xnor U13396 (N_13396,N_12972,N_12511);
nand U13397 (N_13397,N_12972,N_12567);
or U13398 (N_13398,N_12872,N_12650);
and U13399 (N_13399,N_12515,N_12630);
nand U13400 (N_13400,N_12909,N_12957);
or U13401 (N_13401,N_12797,N_12537);
xor U13402 (N_13402,N_12842,N_12967);
nand U13403 (N_13403,N_12598,N_12987);
and U13404 (N_13404,N_12774,N_12989);
or U13405 (N_13405,N_12819,N_12543);
xnor U13406 (N_13406,N_12502,N_12847);
nand U13407 (N_13407,N_12600,N_12638);
nor U13408 (N_13408,N_12893,N_12676);
or U13409 (N_13409,N_12504,N_12537);
xnor U13410 (N_13410,N_12615,N_12519);
nand U13411 (N_13411,N_12736,N_12816);
nand U13412 (N_13412,N_12979,N_12521);
nor U13413 (N_13413,N_12985,N_12928);
or U13414 (N_13414,N_12755,N_12525);
and U13415 (N_13415,N_12904,N_12942);
or U13416 (N_13416,N_12618,N_12830);
xnor U13417 (N_13417,N_12554,N_12738);
nand U13418 (N_13418,N_12786,N_12813);
nand U13419 (N_13419,N_12913,N_12525);
nand U13420 (N_13420,N_12700,N_12547);
and U13421 (N_13421,N_12712,N_12621);
and U13422 (N_13422,N_12696,N_12881);
xor U13423 (N_13423,N_12913,N_12600);
nor U13424 (N_13424,N_12818,N_12685);
nor U13425 (N_13425,N_12625,N_12595);
nor U13426 (N_13426,N_12666,N_12678);
nand U13427 (N_13427,N_12510,N_12567);
or U13428 (N_13428,N_12642,N_12798);
nor U13429 (N_13429,N_12581,N_12714);
and U13430 (N_13430,N_12653,N_12676);
nor U13431 (N_13431,N_12988,N_12702);
nand U13432 (N_13432,N_12701,N_12570);
or U13433 (N_13433,N_12780,N_12578);
or U13434 (N_13434,N_12917,N_12566);
nand U13435 (N_13435,N_12971,N_12530);
xnor U13436 (N_13436,N_12524,N_12757);
xnor U13437 (N_13437,N_12584,N_12675);
or U13438 (N_13438,N_12560,N_12830);
xnor U13439 (N_13439,N_12593,N_12721);
nand U13440 (N_13440,N_12737,N_12738);
xnor U13441 (N_13441,N_12662,N_12858);
or U13442 (N_13442,N_12861,N_12661);
xnor U13443 (N_13443,N_12917,N_12545);
and U13444 (N_13444,N_12932,N_12572);
nor U13445 (N_13445,N_12849,N_12904);
nand U13446 (N_13446,N_12784,N_12717);
and U13447 (N_13447,N_12756,N_12871);
nor U13448 (N_13448,N_12975,N_12814);
and U13449 (N_13449,N_12801,N_12983);
or U13450 (N_13450,N_12906,N_12525);
xnor U13451 (N_13451,N_12658,N_12825);
and U13452 (N_13452,N_12574,N_12623);
nor U13453 (N_13453,N_12830,N_12792);
nand U13454 (N_13454,N_12986,N_12760);
nand U13455 (N_13455,N_12756,N_12977);
and U13456 (N_13456,N_12760,N_12812);
or U13457 (N_13457,N_12895,N_12955);
xnor U13458 (N_13458,N_12849,N_12742);
nor U13459 (N_13459,N_12667,N_12729);
xor U13460 (N_13460,N_12857,N_12973);
nor U13461 (N_13461,N_12833,N_12877);
nor U13462 (N_13462,N_12775,N_12507);
or U13463 (N_13463,N_12734,N_12861);
nor U13464 (N_13464,N_12813,N_12762);
xor U13465 (N_13465,N_12594,N_12623);
xor U13466 (N_13466,N_12654,N_12979);
and U13467 (N_13467,N_12922,N_12555);
nand U13468 (N_13468,N_12985,N_12862);
xnor U13469 (N_13469,N_12959,N_12668);
and U13470 (N_13470,N_12689,N_12743);
nand U13471 (N_13471,N_12773,N_12697);
nand U13472 (N_13472,N_12644,N_12526);
and U13473 (N_13473,N_12605,N_12716);
nand U13474 (N_13474,N_12890,N_12863);
or U13475 (N_13475,N_12641,N_12874);
or U13476 (N_13476,N_12863,N_12758);
and U13477 (N_13477,N_12551,N_12715);
nor U13478 (N_13478,N_12565,N_12655);
nor U13479 (N_13479,N_12957,N_12819);
and U13480 (N_13480,N_12561,N_12548);
or U13481 (N_13481,N_12858,N_12773);
nor U13482 (N_13482,N_12586,N_12646);
nand U13483 (N_13483,N_12617,N_12689);
or U13484 (N_13484,N_12565,N_12794);
and U13485 (N_13485,N_12587,N_12874);
and U13486 (N_13486,N_12515,N_12931);
or U13487 (N_13487,N_12922,N_12990);
or U13488 (N_13488,N_12774,N_12554);
or U13489 (N_13489,N_12625,N_12979);
and U13490 (N_13490,N_12529,N_12912);
or U13491 (N_13491,N_12722,N_12847);
or U13492 (N_13492,N_12717,N_12612);
nand U13493 (N_13493,N_12929,N_12676);
nand U13494 (N_13494,N_12776,N_12764);
and U13495 (N_13495,N_12741,N_12713);
nor U13496 (N_13496,N_12819,N_12752);
xnor U13497 (N_13497,N_12580,N_12888);
xor U13498 (N_13498,N_12680,N_12607);
and U13499 (N_13499,N_12547,N_12887);
xnor U13500 (N_13500,N_13158,N_13485);
or U13501 (N_13501,N_13212,N_13326);
nor U13502 (N_13502,N_13237,N_13433);
and U13503 (N_13503,N_13074,N_13358);
nor U13504 (N_13504,N_13077,N_13416);
nand U13505 (N_13505,N_13236,N_13403);
and U13506 (N_13506,N_13461,N_13214);
nor U13507 (N_13507,N_13006,N_13116);
or U13508 (N_13508,N_13365,N_13143);
and U13509 (N_13509,N_13062,N_13346);
xnor U13510 (N_13510,N_13444,N_13164);
xnor U13511 (N_13511,N_13127,N_13063);
xnor U13512 (N_13512,N_13159,N_13341);
and U13513 (N_13513,N_13252,N_13203);
nor U13514 (N_13514,N_13141,N_13474);
and U13515 (N_13515,N_13150,N_13178);
xor U13516 (N_13516,N_13453,N_13221);
or U13517 (N_13517,N_13443,N_13036);
or U13518 (N_13518,N_13423,N_13262);
xor U13519 (N_13519,N_13470,N_13300);
or U13520 (N_13520,N_13051,N_13029);
xor U13521 (N_13521,N_13240,N_13407);
or U13522 (N_13522,N_13439,N_13340);
xnor U13523 (N_13523,N_13015,N_13314);
and U13524 (N_13524,N_13291,N_13278);
nor U13525 (N_13525,N_13184,N_13411);
nor U13526 (N_13526,N_13481,N_13122);
nand U13527 (N_13527,N_13157,N_13088);
nor U13528 (N_13528,N_13040,N_13351);
or U13529 (N_13529,N_13138,N_13211);
nand U13530 (N_13530,N_13384,N_13480);
nor U13531 (N_13531,N_13370,N_13373);
and U13532 (N_13532,N_13058,N_13218);
nand U13533 (N_13533,N_13465,N_13170);
nor U13534 (N_13534,N_13147,N_13489);
nand U13535 (N_13535,N_13191,N_13321);
or U13536 (N_13536,N_13255,N_13269);
and U13537 (N_13537,N_13372,N_13107);
or U13538 (N_13538,N_13226,N_13283);
xnor U13539 (N_13539,N_13251,N_13356);
and U13540 (N_13540,N_13316,N_13254);
nor U13541 (N_13541,N_13348,N_13312);
and U13542 (N_13542,N_13046,N_13263);
and U13543 (N_13543,N_13457,N_13188);
xor U13544 (N_13544,N_13414,N_13331);
nand U13545 (N_13545,N_13169,N_13376);
nand U13546 (N_13546,N_13038,N_13258);
or U13547 (N_13547,N_13096,N_13215);
nor U13548 (N_13548,N_13193,N_13472);
xor U13549 (N_13549,N_13030,N_13183);
xnor U13550 (N_13550,N_13322,N_13264);
nand U13551 (N_13551,N_13388,N_13002);
or U13552 (N_13552,N_13125,N_13249);
nand U13553 (N_13553,N_13248,N_13067);
xor U13554 (N_13554,N_13202,N_13056);
or U13555 (N_13555,N_13167,N_13111);
xnor U13556 (N_13556,N_13082,N_13228);
nand U13557 (N_13557,N_13431,N_13247);
nand U13558 (N_13558,N_13394,N_13295);
xor U13559 (N_13559,N_13034,N_13378);
or U13560 (N_13560,N_13393,N_13043);
or U13561 (N_13561,N_13265,N_13287);
and U13562 (N_13562,N_13224,N_13464);
and U13563 (N_13563,N_13435,N_13012);
or U13564 (N_13564,N_13460,N_13256);
nor U13565 (N_13565,N_13400,N_13279);
nor U13566 (N_13566,N_13174,N_13344);
nand U13567 (N_13567,N_13311,N_13374);
and U13568 (N_13568,N_13054,N_13302);
nor U13569 (N_13569,N_13177,N_13286);
nand U13570 (N_13570,N_13219,N_13119);
and U13571 (N_13571,N_13126,N_13333);
or U13572 (N_13572,N_13086,N_13128);
and U13573 (N_13573,N_13019,N_13273);
and U13574 (N_13574,N_13140,N_13362);
or U13575 (N_13575,N_13446,N_13179);
or U13576 (N_13576,N_13078,N_13234);
and U13577 (N_13577,N_13412,N_13496);
or U13578 (N_13578,N_13299,N_13154);
nand U13579 (N_13579,N_13319,N_13024);
nand U13580 (N_13580,N_13440,N_13442);
nor U13581 (N_13581,N_13387,N_13366);
nor U13582 (N_13582,N_13361,N_13136);
nor U13583 (N_13583,N_13395,N_13428);
nor U13584 (N_13584,N_13288,N_13137);
nor U13585 (N_13585,N_13201,N_13332);
nor U13586 (N_13586,N_13097,N_13200);
or U13587 (N_13587,N_13271,N_13098);
and U13588 (N_13588,N_13383,N_13168);
xor U13589 (N_13589,N_13010,N_13290);
or U13590 (N_13590,N_13364,N_13021);
nor U13591 (N_13591,N_13343,N_13223);
nand U13592 (N_13592,N_13008,N_13044);
and U13593 (N_13593,N_13229,N_13268);
xor U13594 (N_13594,N_13171,N_13245);
and U13595 (N_13595,N_13220,N_13285);
xor U13596 (N_13596,N_13359,N_13005);
and U13597 (N_13597,N_13353,N_13317);
or U13598 (N_13598,N_13071,N_13482);
or U13599 (N_13599,N_13275,N_13345);
or U13600 (N_13600,N_13094,N_13330);
and U13601 (N_13601,N_13301,N_13079);
and U13602 (N_13602,N_13477,N_13385);
nor U13603 (N_13603,N_13404,N_13155);
and U13604 (N_13604,N_13003,N_13192);
nor U13605 (N_13605,N_13134,N_13368);
nand U13606 (N_13606,N_13061,N_13199);
and U13607 (N_13607,N_13109,N_13305);
and U13608 (N_13608,N_13497,N_13099);
nand U13609 (N_13609,N_13360,N_13050);
nand U13610 (N_13610,N_13250,N_13084);
xnor U13611 (N_13611,N_13462,N_13113);
nor U13612 (N_13612,N_13281,N_13156);
and U13613 (N_13613,N_13132,N_13048);
or U13614 (N_13614,N_13402,N_13093);
xnor U13615 (N_13615,N_13076,N_13406);
and U13616 (N_13616,N_13274,N_13369);
or U13617 (N_13617,N_13419,N_13208);
or U13618 (N_13618,N_13070,N_13430);
or U13619 (N_13619,N_13246,N_13313);
xnor U13620 (N_13620,N_13447,N_13148);
or U13621 (N_13621,N_13471,N_13175);
nor U13622 (N_13622,N_13327,N_13325);
nor U13623 (N_13623,N_13189,N_13037);
xor U13624 (N_13624,N_13080,N_13334);
and U13625 (N_13625,N_13410,N_13144);
xor U13626 (N_13626,N_13422,N_13018);
and U13627 (N_13627,N_13115,N_13053);
xor U13628 (N_13628,N_13222,N_13182);
or U13629 (N_13629,N_13467,N_13090);
nand U13630 (N_13630,N_13475,N_13196);
nand U13631 (N_13631,N_13142,N_13367);
or U13632 (N_13632,N_13375,N_13072);
and U13633 (N_13633,N_13092,N_13429);
nor U13634 (N_13634,N_13100,N_13456);
nand U13635 (N_13635,N_13289,N_13459);
xor U13636 (N_13636,N_13418,N_13272);
and U13637 (N_13637,N_13197,N_13232);
xnor U13638 (N_13638,N_13032,N_13424);
nand U13639 (N_13639,N_13172,N_13397);
xnor U13640 (N_13640,N_13257,N_13448);
nor U13641 (N_13641,N_13160,N_13016);
and U13642 (N_13642,N_13045,N_13194);
and U13643 (N_13643,N_13039,N_13357);
or U13644 (N_13644,N_13320,N_13130);
or U13645 (N_13645,N_13124,N_13478);
or U13646 (N_13646,N_13479,N_13120);
nor U13647 (N_13647,N_13225,N_13149);
xor U13648 (N_13648,N_13110,N_13118);
nand U13649 (N_13649,N_13371,N_13487);
or U13650 (N_13650,N_13438,N_13186);
nand U13651 (N_13651,N_13213,N_13282);
or U13652 (N_13652,N_13195,N_13004);
and U13653 (N_13653,N_13025,N_13028);
or U13654 (N_13654,N_13151,N_13476);
or U13655 (N_13655,N_13047,N_13233);
nor U13656 (N_13656,N_13484,N_13108);
nor U13657 (N_13657,N_13121,N_13382);
and U13658 (N_13658,N_13405,N_13052);
xnor U13659 (N_13659,N_13425,N_13060);
and U13660 (N_13660,N_13280,N_13355);
and U13661 (N_13661,N_13347,N_13161);
nor U13662 (N_13662,N_13401,N_13013);
nand U13663 (N_13663,N_13198,N_13339);
or U13664 (N_13664,N_13315,N_13399);
nor U13665 (N_13665,N_13427,N_13105);
or U13666 (N_13666,N_13328,N_13276);
nor U13667 (N_13667,N_13452,N_13260);
nor U13668 (N_13668,N_13450,N_13001);
or U13669 (N_13669,N_13103,N_13337);
and U13670 (N_13670,N_13227,N_13104);
or U13671 (N_13671,N_13277,N_13354);
or U13672 (N_13672,N_13009,N_13298);
nand U13673 (N_13673,N_13095,N_13242);
and U13674 (N_13674,N_13190,N_13035);
or U13675 (N_13675,N_13238,N_13020);
nor U13676 (N_13676,N_13454,N_13057);
nor U13677 (N_13677,N_13350,N_13117);
and U13678 (N_13678,N_13491,N_13436);
nand U13679 (N_13679,N_13235,N_13011);
and U13680 (N_13680,N_13267,N_13102);
xor U13681 (N_13681,N_13204,N_13210);
nand U13682 (N_13682,N_13284,N_13270);
and U13683 (N_13683,N_13075,N_13458);
xor U13684 (N_13684,N_13413,N_13081);
xor U13685 (N_13685,N_13490,N_13391);
xnor U13686 (N_13686,N_13310,N_13217);
xnor U13687 (N_13687,N_13181,N_13396);
and U13688 (N_13688,N_13014,N_13434);
or U13689 (N_13689,N_13389,N_13441);
nand U13690 (N_13690,N_13468,N_13069);
and U13691 (N_13691,N_13230,N_13083);
xor U13692 (N_13692,N_13101,N_13381);
nor U13693 (N_13693,N_13499,N_13049);
or U13694 (N_13694,N_13417,N_13055);
nor U13695 (N_13695,N_13293,N_13244);
nand U13696 (N_13696,N_13017,N_13492);
nand U13697 (N_13697,N_13379,N_13266);
and U13698 (N_13698,N_13304,N_13133);
and U13699 (N_13699,N_13445,N_13377);
or U13700 (N_13700,N_13152,N_13106);
xor U13701 (N_13701,N_13306,N_13495);
and U13702 (N_13702,N_13087,N_13031);
or U13703 (N_13703,N_13176,N_13166);
xnor U13704 (N_13704,N_13303,N_13022);
and U13705 (N_13705,N_13065,N_13089);
nand U13706 (N_13706,N_13068,N_13064);
xor U13707 (N_13707,N_13163,N_13390);
nor U13708 (N_13708,N_13261,N_13408);
or U13709 (N_13709,N_13409,N_13297);
and U13710 (N_13710,N_13498,N_13073);
or U13711 (N_13711,N_13173,N_13349);
xor U13712 (N_13712,N_13129,N_13398);
xnor U13713 (N_13713,N_13135,N_13473);
nor U13714 (N_13714,N_13153,N_13123);
xnor U13715 (N_13715,N_13309,N_13042);
nor U13716 (N_13716,N_13165,N_13296);
or U13717 (N_13717,N_13187,N_13033);
xnor U13718 (N_13718,N_13380,N_13463);
or U13719 (N_13719,N_13486,N_13259);
nand U13720 (N_13720,N_13318,N_13449);
xor U13721 (N_13721,N_13085,N_13041);
and U13722 (N_13722,N_13216,N_13059);
and U13723 (N_13723,N_13000,N_13185);
and U13724 (N_13724,N_13241,N_13294);
nand U13725 (N_13725,N_13091,N_13493);
and U13726 (N_13726,N_13112,N_13066);
or U13727 (N_13727,N_13206,N_13386);
and U13728 (N_13728,N_13308,N_13335);
or U13729 (N_13729,N_13023,N_13209);
or U13730 (N_13730,N_13342,N_13421);
and U13731 (N_13731,N_13243,N_13437);
and U13732 (N_13732,N_13292,N_13426);
or U13733 (N_13733,N_13338,N_13145);
and U13734 (N_13734,N_13131,N_13415);
or U13735 (N_13735,N_13162,N_13451);
nand U13736 (N_13736,N_13494,N_13026);
nand U13737 (N_13737,N_13239,N_13469);
nor U13738 (N_13738,N_13420,N_13205);
or U13739 (N_13739,N_13483,N_13180);
and U13740 (N_13740,N_13466,N_13336);
nor U13741 (N_13741,N_13207,N_13307);
or U13742 (N_13742,N_13363,N_13231);
or U13743 (N_13743,N_13352,N_13324);
xor U13744 (N_13744,N_13114,N_13139);
nor U13745 (N_13745,N_13432,N_13007);
xnor U13746 (N_13746,N_13329,N_13027);
and U13747 (N_13747,N_13455,N_13323);
nor U13748 (N_13748,N_13488,N_13392);
xor U13749 (N_13749,N_13146,N_13253);
nand U13750 (N_13750,N_13226,N_13277);
nor U13751 (N_13751,N_13104,N_13407);
and U13752 (N_13752,N_13484,N_13156);
nand U13753 (N_13753,N_13155,N_13491);
or U13754 (N_13754,N_13361,N_13228);
or U13755 (N_13755,N_13115,N_13140);
nor U13756 (N_13756,N_13223,N_13332);
and U13757 (N_13757,N_13124,N_13366);
xnor U13758 (N_13758,N_13035,N_13045);
xnor U13759 (N_13759,N_13400,N_13258);
or U13760 (N_13760,N_13326,N_13006);
or U13761 (N_13761,N_13168,N_13427);
or U13762 (N_13762,N_13188,N_13369);
xnor U13763 (N_13763,N_13098,N_13251);
nor U13764 (N_13764,N_13393,N_13441);
nor U13765 (N_13765,N_13442,N_13159);
nor U13766 (N_13766,N_13148,N_13321);
nand U13767 (N_13767,N_13418,N_13299);
xnor U13768 (N_13768,N_13455,N_13271);
and U13769 (N_13769,N_13295,N_13471);
and U13770 (N_13770,N_13346,N_13437);
or U13771 (N_13771,N_13215,N_13271);
or U13772 (N_13772,N_13113,N_13302);
or U13773 (N_13773,N_13096,N_13218);
and U13774 (N_13774,N_13258,N_13218);
and U13775 (N_13775,N_13025,N_13042);
or U13776 (N_13776,N_13369,N_13249);
nand U13777 (N_13777,N_13438,N_13033);
nor U13778 (N_13778,N_13147,N_13486);
and U13779 (N_13779,N_13440,N_13251);
nand U13780 (N_13780,N_13388,N_13301);
xor U13781 (N_13781,N_13322,N_13235);
or U13782 (N_13782,N_13384,N_13040);
xnor U13783 (N_13783,N_13412,N_13234);
nand U13784 (N_13784,N_13058,N_13008);
nand U13785 (N_13785,N_13397,N_13257);
xor U13786 (N_13786,N_13068,N_13434);
xnor U13787 (N_13787,N_13309,N_13079);
xnor U13788 (N_13788,N_13064,N_13494);
nand U13789 (N_13789,N_13086,N_13016);
nand U13790 (N_13790,N_13118,N_13060);
or U13791 (N_13791,N_13257,N_13126);
xnor U13792 (N_13792,N_13431,N_13491);
xor U13793 (N_13793,N_13017,N_13491);
nor U13794 (N_13794,N_13320,N_13115);
xnor U13795 (N_13795,N_13033,N_13076);
xnor U13796 (N_13796,N_13211,N_13102);
xnor U13797 (N_13797,N_13350,N_13266);
or U13798 (N_13798,N_13139,N_13420);
and U13799 (N_13799,N_13212,N_13209);
nand U13800 (N_13800,N_13404,N_13272);
nor U13801 (N_13801,N_13400,N_13487);
or U13802 (N_13802,N_13478,N_13010);
and U13803 (N_13803,N_13412,N_13145);
xnor U13804 (N_13804,N_13405,N_13040);
xor U13805 (N_13805,N_13224,N_13283);
nand U13806 (N_13806,N_13274,N_13111);
nor U13807 (N_13807,N_13025,N_13138);
nand U13808 (N_13808,N_13436,N_13156);
or U13809 (N_13809,N_13366,N_13080);
nor U13810 (N_13810,N_13385,N_13000);
xor U13811 (N_13811,N_13123,N_13207);
nand U13812 (N_13812,N_13184,N_13301);
xnor U13813 (N_13813,N_13404,N_13156);
or U13814 (N_13814,N_13133,N_13187);
and U13815 (N_13815,N_13161,N_13231);
xnor U13816 (N_13816,N_13017,N_13264);
and U13817 (N_13817,N_13354,N_13440);
and U13818 (N_13818,N_13242,N_13410);
xnor U13819 (N_13819,N_13239,N_13498);
and U13820 (N_13820,N_13367,N_13301);
xor U13821 (N_13821,N_13066,N_13332);
or U13822 (N_13822,N_13186,N_13347);
nand U13823 (N_13823,N_13023,N_13425);
and U13824 (N_13824,N_13223,N_13131);
nor U13825 (N_13825,N_13486,N_13076);
or U13826 (N_13826,N_13478,N_13459);
nor U13827 (N_13827,N_13211,N_13091);
nor U13828 (N_13828,N_13067,N_13188);
nor U13829 (N_13829,N_13490,N_13486);
nand U13830 (N_13830,N_13342,N_13015);
nor U13831 (N_13831,N_13371,N_13265);
or U13832 (N_13832,N_13281,N_13037);
nand U13833 (N_13833,N_13117,N_13356);
or U13834 (N_13834,N_13488,N_13473);
and U13835 (N_13835,N_13300,N_13359);
nand U13836 (N_13836,N_13465,N_13262);
xnor U13837 (N_13837,N_13498,N_13131);
nor U13838 (N_13838,N_13120,N_13399);
nand U13839 (N_13839,N_13093,N_13035);
nor U13840 (N_13840,N_13175,N_13112);
xor U13841 (N_13841,N_13437,N_13196);
nand U13842 (N_13842,N_13457,N_13109);
xor U13843 (N_13843,N_13133,N_13281);
and U13844 (N_13844,N_13002,N_13463);
nand U13845 (N_13845,N_13152,N_13401);
xor U13846 (N_13846,N_13250,N_13199);
and U13847 (N_13847,N_13209,N_13479);
nor U13848 (N_13848,N_13427,N_13058);
nor U13849 (N_13849,N_13446,N_13457);
nor U13850 (N_13850,N_13325,N_13025);
nand U13851 (N_13851,N_13160,N_13103);
or U13852 (N_13852,N_13316,N_13213);
xnor U13853 (N_13853,N_13175,N_13262);
or U13854 (N_13854,N_13083,N_13452);
and U13855 (N_13855,N_13457,N_13413);
nand U13856 (N_13856,N_13459,N_13125);
xor U13857 (N_13857,N_13253,N_13200);
nand U13858 (N_13858,N_13339,N_13270);
nor U13859 (N_13859,N_13235,N_13056);
or U13860 (N_13860,N_13169,N_13490);
and U13861 (N_13861,N_13488,N_13271);
and U13862 (N_13862,N_13135,N_13016);
nor U13863 (N_13863,N_13286,N_13276);
nor U13864 (N_13864,N_13139,N_13418);
or U13865 (N_13865,N_13032,N_13401);
xnor U13866 (N_13866,N_13436,N_13306);
nand U13867 (N_13867,N_13236,N_13142);
nand U13868 (N_13868,N_13214,N_13176);
or U13869 (N_13869,N_13280,N_13299);
nand U13870 (N_13870,N_13291,N_13336);
nor U13871 (N_13871,N_13387,N_13277);
xor U13872 (N_13872,N_13250,N_13097);
xor U13873 (N_13873,N_13326,N_13298);
nor U13874 (N_13874,N_13368,N_13109);
xor U13875 (N_13875,N_13015,N_13488);
nand U13876 (N_13876,N_13207,N_13223);
and U13877 (N_13877,N_13408,N_13148);
or U13878 (N_13878,N_13237,N_13468);
xnor U13879 (N_13879,N_13033,N_13478);
xnor U13880 (N_13880,N_13129,N_13112);
nor U13881 (N_13881,N_13362,N_13012);
or U13882 (N_13882,N_13198,N_13123);
nor U13883 (N_13883,N_13274,N_13379);
and U13884 (N_13884,N_13139,N_13029);
and U13885 (N_13885,N_13419,N_13325);
nand U13886 (N_13886,N_13316,N_13114);
nor U13887 (N_13887,N_13339,N_13387);
xnor U13888 (N_13888,N_13386,N_13226);
nor U13889 (N_13889,N_13259,N_13333);
or U13890 (N_13890,N_13185,N_13281);
and U13891 (N_13891,N_13180,N_13267);
xor U13892 (N_13892,N_13497,N_13192);
nor U13893 (N_13893,N_13341,N_13136);
and U13894 (N_13894,N_13383,N_13424);
and U13895 (N_13895,N_13060,N_13030);
nand U13896 (N_13896,N_13291,N_13145);
or U13897 (N_13897,N_13040,N_13272);
and U13898 (N_13898,N_13264,N_13337);
nor U13899 (N_13899,N_13315,N_13351);
xnor U13900 (N_13900,N_13001,N_13482);
and U13901 (N_13901,N_13302,N_13467);
and U13902 (N_13902,N_13116,N_13274);
nand U13903 (N_13903,N_13338,N_13196);
nand U13904 (N_13904,N_13210,N_13454);
or U13905 (N_13905,N_13217,N_13471);
nor U13906 (N_13906,N_13381,N_13130);
nor U13907 (N_13907,N_13422,N_13326);
and U13908 (N_13908,N_13248,N_13379);
and U13909 (N_13909,N_13178,N_13406);
nor U13910 (N_13910,N_13227,N_13061);
and U13911 (N_13911,N_13145,N_13461);
and U13912 (N_13912,N_13181,N_13006);
and U13913 (N_13913,N_13045,N_13307);
nand U13914 (N_13914,N_13271,N_13012);
nor U13915 (N_13915,N_13444,N_13254);
and U13916 (N_13916,N_13398,N_13078);
or U13917 (N_13917,N_13200,N_13120);
and U13918 (N_13918,N_13215,N_13396);
and U13919 (N_13919,N_13151,N_13097);
nand U13920 (N_13920,N_13365,N_13014);
nor U13921 (N_13921,N_13355,N_13131);
or U13922 (N_13922,N_13003,N_13480);
xnor U13923 (N_13923,N_13186,N_13472);
or U13924 (N_13924,N_13086,N_13192);
or U13925 (N_13925,N_13470,N_13348);
or U13926 (N_13926,N_13055,N_13077);
nand U13927 (N_13927,N_13294,N_13490);
nor U13928 (N_13928,N_13201,N_13468);
nand U13929 (N_13929,N_13215,N_13071);
or U13930 (N_13930,N_13000,N_13087);
nand U13931 (N_13931,N_13069,N_13493);
and U13932 (N_13932,N_13114,N_13435);
xor U13933 (N_13933,N_13006,N_13007);
xnor U13934 (N_13934,N_13375,N_13050);
nor U13935 (N_13935,N_13283,N_13292);
and U13936 (N_13936,N_13195,N_13429);
or U13937 (N_13937,N_13035,N_13016);
or U13938 (N_13938,N_13392,N_13312);
nand U13939 (N_13939,N_13403,N_13462);
nand U13940 (N_13940,N_13414,N_13262);
or U13941 (N_13941,N_13252,N_13223);
nor U13942 (N_13942,N_13281,N_13287);
xnor U13943 (N_13943,N_13113,N_13208);
nor U13944 (N_13944,N_13161,N_13446);
nor U13945 (N_13945,N_13292,N_13458);
or U13946 (N_13946,N_13442,N_13284);
nor U13947 (N_13947,N_13485,N_13224);
nor U13948 (N_13948,N_13145,N_13019);
xor U13949 (N_13949,N_13179,N_13434);
nor U13950 (N_13950,N_13025,N_13460);
xor U13951 (N_13951,N_13436,N_13365);
and U13952 (N_13952,N_13021,N_13242);
and U13953 (N_13953,N_13224,N_13008);
nand U13954 (N_13954,N_13455,N_13130);
nor U13955 (N_13955,N_13165,N_13361);
nor U13956 (N_13956,N_13267,N_13357);
nand U13957 (N_13957,N_13425,N_13472);
and U13958 (N_13958,N_13089,N_13123);
and U13959 (N_13959,N_13064,N_13388);
or U13960 (N_13960,N_13420,N_13168);
and U13961 (N_13961,N_13379,N_13202);
xnor U13962 (N_13962,N_13166,N_13403);
xor U13963 (N_13963,N_13210,N_13147);
nand U13964 (N_13964,N_13477,N_13291);
or U13965 (N_13965,N_13017,N_13157);
xnor U13966 (N_13966,N_13383,N_13164);
nand U13967 (N_13967,N_13192,N_13154);
xor U13968 (N_13968,N_13299,N_13392);
nand U13969 (N_13969,N_13100,N_13223);
xnor U13970 (N_13970,N_13116,N_13137);
xnor U13971 (N_13971,N_13295,N_13259);
nand U13972 (N_13972,N_13453,N_13174);
nor U13973 (N_13973,N_13198,N_13383);
or U13974 (N_13974,N_13286,N_13040);
nand U13975 (N_13975,N_13416,N_13468);
or U13976 (N_13976,N_13453,N_13172);
nand U13977 (N_13977,N_13242,N_13461);
xor U13978 (N_13978,N_13434,N_13194);
and U13979 (N_13979,N_13211,N_13479);
xor U13980 (N_13980,N_13256,N_13233);
nor U13981 (N_13981,N_13331,N_13036);
xnor U13982 (N_13982,N_13422,N_13086);
and U13983 (N_13983,N_13035,N_13072);
and U13984 (N_13984,N_13383,N_13262);
nor U13985 (N_13985,N_13176,N_13193);
or U13986 (N_13986,N_13075,N_13101);
nand U13987 (N_13987,N_13186,N_13056);
or U13988 (N_13988,N_13110,N_13421);
and U13989 (N_13989,N_13059,N_13051);
nand U13990 (N_13990,N_13057,N_13390);
nand U13991 (N_13991,N_13386,N_13186);
or U13992 (N_13992,N_13209,N_13333);
nand U13993 (N_13993,N_13443,N_13201);
or U13994 (N_13994,N_13166,N_13471);
nand U13995 (N_13995,N_13100,N_13136);
and U13996 (N_13996,N_13296,N_13162);
nand U13997 (N_13997,N_13232,N_13019);
or U13998 (N_13998,N_13319,N_13184);
nand U13999 (N_13999,N_13113,N_13272);
nor U14000 (N_14000,N_13684,N_13965);
xnor U14001 (N_14001,N_13811,N_13682);
and U14002 (N_14002,N_13578,N_13703);
or U14003 (N_14003,N_13593,N_13590);
nand U14004 (N_14004,N_13954,N_13856);
nand U14005 (N_14005,N_13542,N_13757);
and U14006 (N_14006,N_13918,N_13733);
and U14007 (N_14007,N_13544,N_13775);
or U14008 (N_14008,N_13601,N_13745);
nand U14009 (N_14009,N_13832,N_13584);
xnor U14010 (N_14010,N_13917,N_13790);
or U14011 (N_14011,N_13749,N_13627);
and U14012 (N_14012,N_13834,N_13909);
or U14013 (N_14013,N_13735,N_13949);
and U14014 (N_14014,N_13520,N_13602);
xor U14015 (N_14015,N_13975,N_13724);
or U14016 (N_14016,N_13877,N_13822);
or U14017 (N_14017,N_13994,N_13916);
nand U14018 (N_14018,N_13934,N_13776);
and U14019 (N_14019,N_13689,N_13933);
or U14020 (N_14020,N_13846,N_13892);
and U14021 (N_14021,N_13726,N_13619);
nand U14022 (N_14022,N_13958,N_13680);
or U14023 (N_14023,N_13929,N_13791);
or U14024 (N_14024,N_13903,N_13931);
or U14025 (N_14025,N_13638,N_13581);
xnor U14026 (N_14026,N_13558,N_13562);
xnor U14027 (N_14027,N_13944,N_13759);
xnor U14028 (N_14028,N_13526,N_13632);
and U14029 (N_14029,N_13770,N_13889);
and U14030 (N_14030,N_13717,N_13995);
xor U14031 (N_14031,N_13687,N_13921);
nand U14032 (N_14032,N_13507,N_13881);
xnor U14033 (N_14033,N_13571,N_13744);
or U14034 (N_14034,N_13560,N_13528);
nor U14035 (N_14035,N_13963,N_13829);
nor U14036 (N_14036,N_13527,N_13506);
or U14037 (N_14037,N_13831,N_13945);
nand U14038 (N_14038,N_13884,N_13914);
xnor U14039 (N_14039,N_13614,N_13603);
or U14040 (N_14040,N_13748,N_13647);
xnor U14041 (N_14041,N_13551,N_13823);
and U14042 (N_14042,N_13955,N_13899);
xnor U14043 (N_14043,N_13803,N_13729);
and U14044 (N_14044,N_13683,N_13531);
xor U14045 (N_14045,N_13809,N_13692);
nor U14046 (N_14046,N_13628,N_13974);
and U14047 (N_14047,N_13545,N_13767);
nor U14048 (N_14048,N_13573,N_13651);
or U14049 (N_14049,N_13678,N_13964);
nand U14050 (N_14050,N_13860,N_13814);
or U14051 (N_14051,N_13522,N_13751);
nor U14052 (N_14052,N_13905,N_13755);
nor U14053 (N_14053,N_13736,N_13690);
nand U14054 (N_14054,N_13604,N_13532);
nand U14055 (N_14055,N_13640,N_13552);
or U14056 (N_14056,N_13722,N_13704);
or U14057 (N_14057,N_13812,N_13985);
or U14058 (N_14058,N_13870,N_13984);
or U14059 (N_14059,N_13813,N_13760);
nand U14060 (N_14060,N_13827,N_13959);
xor U14061 (N_14061,N_13752,N_13674);
or U14062 (N_14062,N_13502,N_13566);
xnor U14063 (N_14063,N_13659,N_13838);
or U14064 (N_14064,N_13567,N_13761);
nand U14065 (N_14065,N_13606,N_13774);
and U14066 (N_14066,N_13649,N_13634);
nand U14067 (N_14067,N_13535,N_13730);
and U14068 (N_14068,N_13707,N_13908);
or U14069 (N_14069,N_13895,N_13930);
nor U14070 (N_14070,N_13622,N_13993);
nor U14071 (N_14071,N_13719,N_13504);
nor U14072 (N_14072,N_13723,N_13771);
nand U14073 (N_14073,N_13529,N_13805);
nor U14074 (N_14074,N_13960,N_13720);
xnor U14075 (N_14075,N_13740,N_13997);
xor U14076 (N_14076,N_13671,N_13550);
and U14077 (N_14077,N_13920,N_13589);
or U14078 (N_14078,N_13701,N_13696);
and U14079 (N_14079,N_13842,N_13686);
nor U14080 (N_14080,N_13841,N_13901);
and U14081 (N_14081,N_13864,N_13670);
xnor U14082 (N_14082,N_13521,N_13817);
and U14083 (N_14083,N_13625,N_13655);
and U14084 (N_14084,N_13641,N_13731);
or U14085 (N_14085,N_13913,N_13820);
nand U14086 (N_14086,N_13804,N_13847);
and U14087 (N_14087,N_13543,N_13861);
and U14088 (N_14088,N_13879,N_13777);
or U14089 (N_14089,N_13972,N_13789);
nand U14090 (N_14090,N_13939,N_13509);
and U14091 (N_14091,N_13579,N_13773);
xor U14092 (N_14092,N_13828,N_13795);
xnor U14093 (N_14093,N_13948,N_13925);
nor U14094 (N_14094,N_13605,N_13672);
nand U14095 (N_14095,N_13597,N_13992);
nand U14096 (N_14096,N_13508,N_13513);
or U14097 (N_14097,N_13624,N_13612);
nand U14098 (N_14098,N_13868,N_13956);
and U14099 (N_14099,N_13762,N_13863);
nor U14100 (N_14100,N_13666,N_13907);
and U14101 (N_14101,N_13798,N_13714);
or U14102 (N_14102,N_13873,N_13662);
nor U14103 (N_14103,N_13968,N_13953);
or U14104 (N_14104,N_13685,N_13952);
nand U14105 (N_14105,N_13650,N_13866);
and U14106 (N_14106,N_13970,N_13854);
and U14107 (N_14107,N_13887,N_13691);
or U14108 (N_14108,N_13936,N_13643);
nor U14109 (N_14109,N_13673,N_13681);
and U14110 (N_14110,N_13768,N_13807);
xnor U14111 (N_14111,N_13679,N_13708);
or U14112 (N_14112,N_13978,N_13940);
and U14113 (N_14113,N_13802,N_13926);
nand U14114 (N_14114,N_13943,N_13980);
xnor U14115 (N_14115,N_13783,N_13951);
or U14116 (N_14116,N_13591,N_13904);
xor U14117 (N_14117,N_13663,N_13615);
nand U14118 (N_14118,N_13753,N_13865);
nor U14119 (N_14119,N_13769,N_13786);
and U14120 (N_14120,N_13635,N_13582);
nor U14121 (N_14121,N_13987,N_13587);
xor U14122 (N_14122,N_13630,N_13547);
xnor U14123 (N_14123,N_13837,N_13941);
and U14124 (N_14124,N_13713,N_13872);
nand U14125 (N_14125,N_13966,N_13986);
xor U14126 (N_14126,N_13924,N_13575);
and U14127 (N_14127,N_13778,N_13912);
and U14128 (N_14128,N_13976,N_13967);
nor U14129 (N_14129,N_13808,N_13851);
nor U14130 (N_14130,N_13503,N_13816);
xnor U14131 (N_14131,N_13859,N_13556);
xor U14132 (N_14132,N_13609,N_13697);
nor U14133 (N_14133,N_13727,N_13962);
xnor U14134 (N_14134,N_13742,N_13710);
and U14135 (N_14135,N_13990,N_13586);
nand U14136 (N_14136,N_13539,N_13636);
xnor U14137 (N_14137,N_13765,N_13781);
or U14138 (N_14138,N_13626,N_13750);
and U14139 (N_14139,N_13700,N_13897);
nand U14140 (N_14140,N_13793,N_13536);
nor U14141 (N_14141,N_13549,N_13613);
xor U14142 (N_14142,N_13855,N_13617);
xnor U14143 (N_14143,N_13711,N_13923);
xor U14144 (N_14144,N_13642,N_13661);
xnor U14145 (N_14145,N_13645,N_13516);
or U14146 (N_14146,N_13555,N_13898);
or U14147 (N_14147,N_13792,N_13836);
or U14148 (N_14148,N_13826,N_13893);
nor U14149 (N_14149,N_13533,N_13554);
or U14150 (N_14150,N_13637,N_13629);
nand U14151 (N_14151,N_13991,N_13902);
and U14152 (N_14152,N_13505,N_13785);
nor U14153 (N_14153,N_13988,N_13937);
nand U14154 (N_14154,N_13585,N_13981);
and U14155 (N_14155,N_13644,N_13927);
or U14156 (N_14156,N_13694,N_13621);
nor U14157 (N_14157,N_13546,N_13537);
and U14158 (N_14158,N_13935,N_13639);
and U14159 (N_14159,N_13942,N_13779);
xor U14160 (N_14160,N_13885,N_13658);
and U14161 (N_14161,N_13824,N_13741);
or U14162 (N_14162,N_13799,N_13737);
nor U14163 (N_14163,N_13510,N_13977);
nor U14164 (N_14164,N_13616,N_13784);
or U14165 (N_14165,N_13947,N_13915);
or U14166 (N_14166,N_13570,N_13894);
xnor U14167 (N_14167,N_13577,N_13538);
or U14168 (N_14168,N_13857,N_13702);
or U14169 (N_14169,N_13982,N_13652);
xor U14170 (N_14170,N_13911,N_13716);
or U14171 (N_14171,N_13734,N_13835);
nand U14172 (N_14172,N_13712,N_13840);
and U14173 (N_14173,N_13706,N_13766);
or U14174 (N_14174,N_13611,N_13961);
xor U14175 (N_14175,N_13782,N_13511);
nand U14176 (N_14176,N_13656,N_13654);
nor U14177 (N_14177,N_13514,N_13633);
nor U14178 (N_14178,N_13677,N_13517);
and U14179 (N_14179,N_13815,N_13825);
nand U14180 (N_14180,N_13764,N_13772);
and U14181 (N_14181,N_13910,N_13890);
nor U14182 (N_14182,N_13867,N_13676);
nor U14183 (N_14183,N_13746,N_13876);
nor U14184 (N_14184,N_13559,N_13530);
xor U14185 (N_14185,N_13797,N_13548);
and U14186 (N_14186,N_13709,N_13796);
nand U14187 (N_14187,N_13763,N_13801);
xnor U14188 (N_14188,N_13883,N_13732);
xnor U14189 (N_14189,N_13849,N_13596);
nor U14190 (N_14190,N_13512,N_13631);
and U14191 (N_14191,N_13878,N_13583);
nor U14192 (N_14192,N_13519,N_13657);
xnor U14193 (N_14193,N_13668,N_13569);
nor U14194 (N_14194,N_13747,N_13852);
nor U14195 (N_14195,N_13756,N_13989);
nor U14196 (N_14196,N_13880,N_13501);
xnor U14197 (N_14197,N_13592,N_13653);
nor U14198 (N_14198,N_13565,N_13819);
xnor U14199 (N_14199,N_13595,N_13646);
nand U14200 (N_14200,N_13999,N_13561);
nand U14201 (N_14201,N_13928,N_13922);
or U14202 (N_14202,N_13810,N_13973);
and U14203 (N_14203,N_13648,N_13728);
or U14204 (N_14204,N_13515,N_13800);
nand U14205 (N_14205,N_13576,N_13718);
xnor U14206 (N_14206,N_13806,N_13787);
nor U14207 (N_14207,N_13705,N_13715);
or U14208 (N_14208,N_13610,N_13598);
xnor U14209 (N_14209,N_13572,N_13599);
xnor U14210 (N_14210,N_13844,N_13833);
and U14211 (N_14211,N_13919,N_13675);
xnor U14212 (N_14212,N_13821,N_13620);
nand U14213 (N_14213,N_13839,N_13938);
and U14214 (N_14214,N_13874,N_13754);
nand U14215 (N_14215,N_13888,N_13896);
and U14216 (N_14216,N_13875,N_13600);
nand U14217 (N_14217,N_13557,N_13983);
or U14218 (N_14218,N_13998,N_13979);
and U14219 (N_14219,N_13699,N_13721);
nor U14220 (N_14220,N_13869,N_13540);
xnor U14221 (N_14221,N_13525,N_13996);
xor U14222 (N_14222,N_13623,N_13794);
xor U14223 (N_14223,N_13564,N_13618);
and U14224 (N_14224,N_13739,N_13698);
nand U14225 (N_14225,N_13688,N_13541);
or U14226 (N_14226,N_13568,N_13830);
nor U14227 (N_14227,N_13950,N_13971);
nor U14228 (N_14228,N_13500,N_13780);
and U14229 (N_14229,N_13843,N_13862);
or U14230 (N_14230,N_13900,N_13932);
and U14231 (N_14231,N_13957,N_13758);
nand U14232 (N_14232,N_13594,N_13693);
or U14233 (N_14233,N_13788,N_13607);
or U14234 (N_14234,N_13524,N_13667);
and U14235 (N_14235,N_13608,N_13853);
xnor U14236 (N_14236,N_13848,N_13845);
xor U14237 (N_14237,N_13695,N_13891);
or U14238 (N_14238,N_13588,N_13725);
xor U14239 (N_14239,N_13534,N_13518);
nand U14240 (N_14240,N_13580,N_13563);
nand U14241 (N_14241,N_13882,N_13858);
nor U14242 (N_14242,N_13574,N_13850);
nor U14243 (N_14243,N_13669,N_13946);
and U14244 (N_14244,N_13743,N_13665);
and U14245 (N_14245,N_13886,N_13660);
nand U14246 (N_14246,N_13969,N_13818);
xnor U14247 (N_14247,N_13906,N_13553);
or U14248 (N_14248,N_13664,N_13738);
or U14249 (N_14249,N_13523,N_13871);
nor U14250 (N_14250,N_13751,N_13611);
xnor U14251 (N_14251,N_13682,N_13624);
nor U14252 (N_14252,N_13637,N_13876);
nand U14253 (N_14253,N_13955,N_13785);
or U14254 (N_14254,N_13827,N_13776);
and U14255 (N_14255,N_13889,N_13913);
xnor U14256 (N_14256,N_13543,N_13797);
nand U14257 (N_14257,N_13538,N_13897);
nor U14258 (N_14258,N_13735,N_13588);
xnor U14259 (N_14259,N_13670,N_13924);
xor U14260 (N_14260,N_13965,N_13735);
nand U14261 (N_14261,N_13763,N_13995);
or U14262 (N_14262,N_13884,N_13707);
nor U14263 (N_14263,N_13795,N_13884);
or U14264 (N_14264,N_13579,N_13831);
or U14265 (N_14265,N_13624,N_13633);
xor U14266 (N_14266,N_13597,N_13956);
and U14267 (N_14267,N_13577,N_13952);
nor U14268 (N_14268,N_13602,N_13536);
xnor U14269 (N_14269,N_13978,N_13721);
nand U14270 (N_14270,N_13674,N_13514);
xnor U14271 (N_14271,N_13583,N_13903);
nor U14272 (N_14272,N_13527,N_13985);
and U14273 (N_14273,N_13919,N_13730);
or U14274 (N_14274,N_13830,N_13522);
nor U14275 (N_14275,N_13673,N_13726);
and U14276 (N_14276,N_13947,N_13880);
nand U14277 (N_14277,N_13876,N_13633);
xor U14278 (N_14278,N_13839,N_13545);
nor U14279 (N_14279,N_13552,N_13681);
nor U14280 (N_14280,N_13853,N_13668);
nand U14281 (N_14281,N_13997,N_13510);
and U14282 (N_14282,N_13823,N_13683);
and U14283 (N_14283,N_13868,N_13704);
xnor U14284 (N_14284,N_13718,N_13727);
nand U14285 (N_14285,N_13940,N_13972);
nor U14286 (N_14286,N_13977,N_13993);
or U14287 (N_14287,N_13511,N_13681);
or U14288 (N_14288,N_13795,N_13802);
nor U14289 (N_14289,N_13683,N_13620);
nor U14290 (N_14290,N_13640,N_13656);
nand U14291 (N_14291,N_13861,N_13859);
xnor U14292 (N_14292,N_13782,N_13833);
nor U14293 (N_14293,N_13850,N_13955);
nand U14294 (N_14294,N_13739,N_13754);
xor U14295 (N_14295,N_13893,N_13769);
or U14296 (N_14296,N_13994,N_13646);
or U14297 (N_14297,N_13569,N_13779);
xnor U14298 (N_14298,N_13951,N_13740);
xor U14299 (N_14299,N_13946,N_13756);
and U14300 (N_14300,N_13901,N_13976);
or U14301 (N_14301,N_13811,N_13695);
or U14302 (N_14302,N_13978,N_13762);
and U14303 (N_14303,N_13696,N_13650);
or U14304 (N_14304,N_13911,N_13548);
and U14305 (N_14305,N_13970,N_13689);
or U14306 (N_14306,N_13953,N_13826);
xnor U14307 (N_14307,N_13577,N_13871);
or U14308 (N_14308,N_13527,N_13530);
nor U14309 (N_14309,N_13871,N_13988);
nand U14310 (N_14310,N_13970,N_13697);
and U14311 (N_14311,N_13521,N_13641);
nand U14312 (N_14312,N_13618,N_13822);
or U14313 (N_14313,N_13987,N_13904);
nor U14314 (N_14314,N_13944,N_13851);
xnor U14315 (N_14315,N_13543,N_13813);
nand U14316 (N_14316,N_13873,N_13938);
nand U14317 (N_14317,N_13593,N_13885);
nand U14318 (N_14318,N_13972,N_13964);
or U14319 (N_14319,N_13632,N_13972);
nor U14320 (N_14320,N_13541,N_13761);
xor U14321 (N_14321,N_13711,N_13583);
xnor U14322 (N_14322,N_13877,N_13865);
nand U14323 (N_14323,N_13516,N_13958);
xor U14324 (N_14324,N_13953,N_13508);
nor U14325 (N_14325,N_13947,N_13592);
or U14326 (N_14326,N_13787,N_13796);
or U14327 (N_14327,N_13620,N_13516);
xnor U14328 (N_14328,N_13795,N_13601);
nor U14329 (N_14329,N_13746,N_13741);
nand U14330 (N_14330,N_13719,N_13900);
nand U14331 (N_14331,N_13686,N_13691);
or U14332 (N_14332,N_13855,N_13998);
nor U14333 (N_14333,N_13860,N_13694);
and U14334 (N_14334,N_13886,N_13874);
nor U14335 (N_14335,N_13866,N_13814);
nand U14336 (N_14336,N_13969,N_13853);
nor U14337 (N_14337,N_13506,N_13778);
xnor U14338 (N_14338,N_13880,N_13766);
nand U14339 (N_14339,N_13868,N_13742);
nor U14340 (N_14340,N_13884,N_13654);
or U14341 (N_14341,N_13553,N_13676);
nand U14342 (N_14342,N_13517,N_13851);
xnor U14343 (N_14343,N_13832,N_13514);
nor U14344 (N_14344,N_13645,N_13649);
nand U14345 (N_14345,N_13713,N_13685);
or U14346 (N_14346,N_13742,N_13559);
nand U14347 (N_14347,N_13849,N_13724);
xor U14348 (N_14348,N_13888,N_13960);
and U14349 (N_14349,N_13774,N_13711);
nand U14350 (N_14350,N_13535,N_13757);
or U14351 (N_14351,N_13730,N_13828);
nor U14352 (N_14352,N_13962,N_13941);
nand U14353 (N_14353,N_13977,N_13537);
or U14354 (N_14354,N_13539,N_13715);
nand U14355 (N_14355,N_13641,N_13636);
nand U14356 (N_14356,N_13868,N_13733);
xor U14357 (N_14357,N_13951,N_13765);
nand U14358 (N_14358,N_13632,N_13764);
nand U14359 (N_14359,N_13779,N_13795);
and U14360 (N_14360,N_13625,N_13852);
and U14361 (N_14361,N_13585,N_13885);
xnor U14362 (N_14362,N_13790,N_13786);
and U14363 (N_14363,N_13760,N_13851);
nand U14364 (N_14364,N_13672,N_13554);
or U14365 (N_14365,N_13619,N_13887);
nand U14366 (N_14366,N_13837,N_13880);
and U14367 (N_14367,N_13860,N_13598);
nor U14368 (N_14368,N_13661,N_13780);
xor U14369 (N_14369,N_13708,N_13519);
nand U14370 (N_14370,N_13766,N_13860);
nor U14371 (N_14371,N_13744,N_13736);
nor U14372 (N_14372,N_13500,N_13784);
nor U14373 (N_14373,N_13919,N_13837);
nand U14374 (N_14374,N_13559,N_13579);
xor U14375 (N_14375,N_13648,N_13536);
xor U14376 (N_14376,N_13967,N_13818);
nand U14377 (N_14377,N_13635,N_13749);
and U14378 (N_14378,N_13867,N_13936);
or U14379 (N_14379,N_13806,N_13749);
and U14380 (N_14380,N_13864,N_13877);
or U14381 (N_14381,N_13638,N_13829);
nor U14382 (N_14382,N_13508,N_13767);
nor U14383 (N_14383,N_13878,N_13895);
and U14384 (N_14384,N_13745,N_13842);
xor U14385 (N_14385,N_13747,N_13610);
nand U14386 (N_14386,N_13676,N_13785);
and U14387 (N_14387,N_13761,N_13552);
nand U14388 (N_14388,N_13510,N_13662);
xor U14389 (N_14389,N_13937,N_13868);
xnor U14390 (N_14390,N_13904,N_13729);
nand U14391 (N_14391,N_13628,N_13704);
or U14392 (N_14392,N_13601,N_13611);
nor U14393 (N_14393,N_13683,N_13667);
or U14394 (N_14394,N_13948,N_13680);
or U14395 (N_14395,N_13823,N_13740);
and U14396 (N_14396,N_13953,N_13769);
or U14397 (N_14397,N_13985,N_13509);
or U14398 (N_14398,N_13821,N_13679);
and U14399 (N_14399,N_13597,N_13672);
xnor U14400 (N_14400,N_13921,N_13811);
and U14401 (N_14401,N_13756,N_13547);
xnor U14402 (N_14402,N_13551,N_13896);
and U14403 (N_14403,N_13767,N_13560);
xnor U14404 (N_14404,N_13605,N_13675);
or U14405 (N_14405,N_13732,N_13721);
or U14406 (N_14406,N_13675,N_13881);
or U14407 (N_14407,N_13781,N_13788);
nand U14408 (N_14408,N_13855,N_13931);
or U14409 (N_14409,N_13617,N_13653);
nand U14410 (N_14410,N_13864,N_13842);
nand U14411 (N_14411,N_13864,N_13854);
nor U14412 (N_14412,N_13832,N_13874);
and U14413 (N_14413,N_13875,N_13548);
or U14414 (N_14414,N_13859,N_13948);
nand U14415 (N_14415,N_13678,N_13944);
nor U14416 (N_14416,N_13627,N_13885);
nor U14417 (N_14417,N_13738,N_13637);
xor U14418 (N_14418,N_13760,N_13972);
or U14419 (N_14419,N_13503,N_13718);
and U14420 (N_14420,N_13963,N_13575);
or U14421 (N_14421,N_13950,N_13595);
and U14422 (N_14422,N_13991,N_13533);
nand U14423 (N_14423,N_13679,N_13743);
nand U14424 (N_14424,N_13866,N_13708);
or U14425 (N_14425,N_13999,N_13514);
nor U14426 (N_14426,N_13767,N_13894);
nand U14427 (N_14427,N_13621,N_13915);
and U14428 (N_14428,N_13959,N_13595);
nand U14429 (N_14429,N_13728,N_13511);
and U14430 (N_14430,N_13963,N_13851);
or U14431 (N_14431,N_13632,N_13619);
nor U14432 (N_14432,N_13692,N_13722);
xor U14433 (N_14433,N_13705,N_13600);
nand U14434 (N_14434,N_13880,N_13550);
and U14435 (N_14435,N_13686,N_13506);
nand U14436 (N_14436,N_13965,N_13545);
and U14437 (N_14437,N_13581,N_13950);
and U14438 (N_14438,N_13808,N_13793);
nor U14439 (N_14439,N_13531,N_13638);
and U14440 (N_14440,N_13597,N_13936);
xor U14441 (N_14441,N_13671,N_13568);
nand U14442 (N_14442,N_13868,N_13570);
or U14443 (N_14443,N_13649,N_13657);
nand U14444 (N_14444,N_13532,N_13680);
or U14445 (N_14445,N_13792,N_13747);
xor U14446 (N_14446,N_13547,N_13557);
or U14447 (N_14447,N_13597,N_13569);
nor U14448 (N_14448,N_13647,N_13568);
and U14449 (N_14449,N_13900,N_13696);
or U14450 (N_14450,N_13612,N_13711);
nand U14451 (N_14451,N_13982,N_13724);
nand U14452 (N_14452,N_13683,N_13845);
xnor U14453 (N_14453,N_13534,N_13842);
and U14454 (N_14454,N_13969,N_13982);
and U14455 (N_14455,N_13944,N_13743);
xnor U14456 (N_14456,N_13854,N_13648);
nand U14457 (N_14457,N_13922,N_13571);
nor U14458 (N_14458,N_13608,N_13673);
xor U14459 (N_14459,N_13825,N_13580);
xnor U14460 (N_14460,N_13515,N_13854);
nand U14461 (N_14461,N_13646,N_13757);
xor U14462 (N_14462,N_13977,N_13549);
nor U14463 (N_14463,N_13662,N_13653);
and U14464 (N_14464,N_13760,N_13788);
nor U14465 (N_14465,N_13929,N_13735);
xor U14466 (N_14466,N_13820,N_13962);
and U14467 (N_14467,N_13587,N_13553);
or U14468 (N_14468,N_13683,N_13677);
nor U14469 (N_14469,N_13711,N_13810);
xnor U14470 (N_14470,N_13525,N_13927);
xnor U14471 (N_14471,N_13711,N_13508);
xnor U14472 (N_14472,N_13537,N_13667);
nand U14473 (N_14473,N_13887,N_13889);
nand U14474 (N_14474,N_13557,N_13502);
nor U14475 (N_14475,N_13922,N_13502);
nand U14476 (N_14476,N_13901,N_13856);
and U14477 (N_14477,N_13534,N_13557);
xnor U14478 (N_14478,N_13749,N_13878);
xnor U14479 (N_14479,N_13968,N_13865);
or U14480 (N_14480,N_13926,N_13768);
or U14481 (N_14481,N_13914,N_13675);
and U14482 (N_14482,N_13508,N_13774);
and U14483 (N_14483,N_13906,N_13629);
nand U14484 (N_14484,N_13995,N_13944);
xnor U14485 (N_14485,N_13957,N_13541);
or U14486 (N_14486,N_13571,N_13575);
and U14487 (N_14487,N_13812,N_13779);
nor U14488 (N_14488,N_13991,N_13535);
nand U14489 (N_14489,N_13621,N_13572);
nor U14490 (N_14490,N_13953,N_13527);
and U14491 (N_14491,N_13784,N_13695);
or U14492 (N_14492,N_13886,N_13861);
nor U14493 (N_14493,N_13960,N_13972);
nor U14494 (N_14494,N_13623,N_13720);
xor U14495 (N_14495,N_13612,N_13724);
or U14496 (N_14496,N_13782,N_13672);
nand U14497 (N_14497,N_13854,N_13538);
nor U14498 (N_14498,N_13571,N_13603);
or U14499 (N_14499,N_13597,N_13633);
nor U14500 (N_14500,N_14303,N_14447);
nor U14501 (N_14501,N_14281,N_14260);
and U14502 (N_14502,N_14055,N_14376);
and U14503 (N_14503,N_14271,N_14078);
nand U14504 (N_14504,N_14466,N_14351);
or U14505 (N_14505,N_14298,N_14272);
xor U14506 (N_14506,N_14157,N_14414);
nor U14507 (N_14507,N_14095,N_14080);
nand U14508 (N_14508,N_14486,N_14053);
and U14509 (N_14509,N_14350,N_14403);
or U14510 (N_14510,N_14261,N_14243);
xor U14511 (N_14511,N_14304,N_14358);
and U14512 (N_14512,N_14086,N_14335);
nor U14513 (N_14513,N_14112,N_14010);
nand U14514 (N_14514,N_14252,N_14172);
or U14515 (N_14515,N_14264,N_14419);
and U14516 (N_14516,N_14062,N_14400);
or U14517 (N_14517,N_14162,N_14191);
nand U14518 (N_14518,N_14488,N_14135);
xnor U14519 (N_14519,N_14217,N_14045);
and U14520 (N_14520,N_14068,N_14472);
nor U14521 (N_14521,N_14392,N_14103);
or U14522 (N_14522,N_14402,N_14174);
nor U14523 (N_14523,N_14290,N_14406);
and U14524 (N_14524,N_14192,N_14332);
and U14525 (N_14525,N_14249,N_14381);
or U14526 (N_14526,N_14389,N_14013);
nand U14527 (N_14527,N_14429,N_14184);
xnor U14528 (N_14528,N_14026,N_14043);
and U14529 (N_14529,N_14064,N_14158);
nor U14530 (N_14530,N_14093,N_14497);
xor U14531 (N_14531,N_14431,N_14333);
and U14532 (N_14532,N_14241,N_14418);
nor U14533 (N_14533,N_14234,N_14235);
nand U14534 (N_14534,N_14166,N_14293);
nor U14535 (N_14535,N_14076,N_14262);
nor U14536 (N_14536,N_14159,N_14239);
nor U14537 (N_14537,N_14073,N_14438);
or U14538 (N_14538,N_14364,N_14000);
xor U14539 (N_14539,N_14363,N_14156);
xor U14540 (N_14540,N_14034,N_14108);
nor U14541 (N_14541,N_14161,N_14451);
nor U14542 (N_14542,N_14285,N_14370);
nor U14543 (N_14543,N_14124,N_14354);
nand U14544 (N_14544,N_14428,N_14101);
nand U14545 (N_14545,N_14199,N_14257);
xor U14546 (N_14546,N_14320,N_14144);
or U14547 (N_14547,N_14321,N_14478);
and U14548 (N_14548,N_14036,N_14269);
nand U14549 (N_14549,N_14048,N_14489);
nor U14550 (N_14550,N_14081,N_14248);
nor U14551 (N_14551,N_14380,N_14373);
nand U14552 (N_14552,N_14467,N_14473);
nor U14553 (N_14553,N_14228,N_14398);
or U14554 (N_14554,N_14485,N_14211);
xnor U14555 (N_14555,N_14223,N_14200);
and U14556 (N_14556,N_14408,N_14202);
or U14557 (N_14557,N_14328,N_14374);
nor U14558 (N_14558,N_14126,N_14160);
xor U14559 (N_14559,N_14399,N_14412);
nor U14560 (N_14560,N_14197,N_14238);
nand U14561 (N_14561,N_14491,N_14039);
and U14562 (N_14562,N_14016,N_14072);
nand U14563 (N_14563,N_14007,N_14183);
nor U14564 (N_14564,N_14463,N_14091);
or U14565 (N_14565,N_14462,N_14457);
nand U14566 (N_14566,N_14394,N_14327);
and U14567 (N_14567,N_14331,N_14263);
and U14568 (N_14568,N_14035,N_14471);
nand U14569 (N_14569,N_14221,N_14063);
or U14570 (N_14570,N_14094,N_14255);
or U14571 (N_14571,N_14137,N_14025);
and U14572 (N_14572,N_14367,N_14177);
and U14573 (N_14573,N_14216,N_14204);
and U14574 (N_14574,N_14132,N_14479);
nor U14575 (N_14575,N_14027,N_14449);
nor U14576 (N_14576,N_14178,N_14378);
nand U14577 (N_14577,N_14029,N_14134);
and U14578 (N_14578,N_14077,N_14100);
xnor U14579 (N_14579,N_14334,N_14317);
xnor U14580 (N_14580,N_14213,N_14206);
xor U14581 (N_14581,N_14165,N_14435);
nand U14582 (N_14582,N_14024,N_14458);
nand U14583 (N_14583,N_14149,N_14338);
nand U14584 (N_14584,N_14404,N_14422);
xnor U14585 (N_14585,N_14110,N_14182);
or U14586 (N_14586,N_14343,N_14268);
xor U14587 (N_14587,N_14127,N_14125);
nor U14588 (N_14588,N_14492,N_14169);
or U14589 (N_14589,N_14357,N_14209);
nor U14590 (N_14590,N_14088,N_14123);
nand U14591 (N_14591,N_14383,N_14098);
nand U14592 (N_14592,N_14342,N_14146);
or U14593 (N_14593,N_14461,N_14012);
xor U14594 (N_14594,N_14251,N_14292);
nor U14595 (N_14595,N_14194,N_14032);
nor U14596 (N_14596,N_14446,N_14410);
and U14597 (N_14597,N_14230,N_14464);
nand U14598 (N_14598,N_14152,N_14314);
and U14599 (N_14599,N_14201,N_14139);
or U14600 (N_14600,N_14136,N_14133);
and U14601 (N_14601,N_14120,N_14102);
nand U14602 (N_14602,N_14273,N_14038);
nor U14603 (N_14603,N_14163,N_14128);
nor U14604 (N_14604,N_14256,N_14360);
xnor U14605 (N_14605,N_14496,N_14006);
nor U14606 (N_14606,N_14205,N_14057);
xor U14607 (N_14607,N_14210,N_14459);
nand U14608 (N_14608,N_14291,N_14322);
or U14609 (N_14609,N_14366,N_14104);
nand U14610 (N_14610,N_14070,N_14115);
and U14611 (N_14611,N_14287,N_14433);
and U14612 (N_14612,N_14150,N_14022);
and U14613 (N_14613,N_14023,N_14288);
xnor U14614 (N_14614,N_14401,N_14416);
nor U14615 (N_14615,N_14484,N_14170);
xor U14616 (N_14616,N_14349,N_14145);
nor U14617 (N_14617,N_14164,N_14030);
xnor U14618 (N_14618,N_14176,N_14324);
nand U14619 (N_14619,N_14470,N_14142);
xor U14620 (N_14620,N_14207,N_14071);
xor U14621 (N_14621,N_14153,N_14041);
or U14622 (N_14622,N_14453,N_14141);
or U14623 (N_14623,N_14282,N_14355);
or U14624 (N_14624,N_14253,N_14225);
xnor U14625 (N_14625,N_14173,N_14415);
nor U14626 (N_14626,N_14369,N_14058);
nand U14627 (N_14627,N_14212,N_14329);
or U14628 (N_14628,N_14075,N_14348);
or U14629 (N_14629,N_14440,N_14368);
xor U14630 (N_14630,N_14498,N_14425);
and U14631 (N_14631,N_14386,N_14495);
nand U14632 (N_14632,N_14307,N_14476);
nor U14633 (N_14633,N_14385,N_14148);
nand U14634 (N_14634,N_14244,N_14226);
nor U14635 (N_14635,N_14337,N_14187);
and U14636 (N_14636,N_14190,N_14005);
nand U14637 (N_14637,N_14109,N_14198);
xor U14638 (N_14638,N_14186,N_14117);
xor U14639 (N_14639,N_14475,N_14296);
or U14640 (N_14640,N_14185,N_14084);
xnor U14641 (N_14641,N_14107,N_14218);
and U14642 (N_14642,N_14372,N_14009);
and U14643 (N_14643,N_14347,N_14424);
nand U14644 (N_14644,N_14037,N_14233);
xor U14645 (N_14645,N_14299,N_14278);
and U14646 (N_14646,N_14316,N_14286);
and U14647 (N_14647,N_14444,N_14353);
and U14648 (N_14648,N_14061,N_14311);
or U14649 (N_14649,N_14279,N_14456);
or U14650 (N_14650,N_14319,N_14236);
and U14651 (N_14651,N_14356,N_14313);
nand U14652 (N_14652,N_14490,N_14494);
or U14653 (N_14653,N_14031,N_14295);
nand U14654 (N_14654,N_14220,N_14004);
nor U14655 (N_14655,N_14289,N_14302);
or U14656 (N_14656,N_14060,N_14131);
or U14657 (N_14657,N_14214,N_14203);
xnor U14658 (N_14658,N_14301,N_14044);
and U14659 (N_14659,N_14167,N_14283);
or U14660 (N_14660,N_14138,N_14439);
nor U14661 (N_14661,N_14056,N_14042);
or U14662 (N_14662,N_14413,N_14247);
nor U14663 (N_14663,N_14395,N_14065);
and U14664 (N_14664,N_14297,N_14151);
xnor U14665 (N_14665,N_14326,N_14245);
or U14666 (N_14666,N_14215,N_14229);
nor U14667 (N_14667,N_14346,N_14014);
nor U14668 (N_14668,N_14480,N_14359);
and U14669 (N_14669,N_14143,N_14046);
xor U14670 (N_14670,N_14224,N_14375);
or U14671 (N_14671,N_14179,N_14460);
nor U14672 (N_14672,N_14054,N_14442);
or U14673 (N_14673,N_14407,N_14396);
nand U14674 (N_14674,N_14340,N_14318);
and U14675 (N_14675,N_14089,N_14017);
or U14676 (N_14676,N_14074,N_14455);
and U14677 (N_14677,N_14168,N_14305);
nor U14678 (N_14678,N_14155,N_14388);
or U14679 (N_14679,N_14430,N_14258);
or U14680 (N_14680,N_14344,N_14082);
nand U14681 (N_14681,N_14188,N_14377);
nand U14682 (N_14682,N_14059,N_14382);
nand U14683 (N_14683,N_14310,N_14465);
nor U14684 (N_14684,N_14308,N_14300);
or U14685 (N_14685,N_14049,N_14411);
or U14686 (N_14686,N_14033,N_14330);
xor U14687 (N_14687,N_14387,N_14477);
nor U14688 (N_14688,N_14274,N_14427);
xnor U14689 (N_14689,N_14284,N_14122);
xor U14690 (N_14690,N_14276,N_14450);
and U14691 (N_14691,N_14083,N_14352);
or U14692 (N_14692,N_14099,N_14001);
nand U14693 (N_14693,N_14114,N_14443);
xnor U14694 (N_14694,N_14066,N_14008);
or U14695 (N_14695,N_14050,N_14002);
nor U14696 (N_14696,N_14265,N_14097);
nor U14697 (N_14697,N_14267,N_14452);
and U14698 (N_14698,N_14116,N_14193);
or U14699 (N_14699,N_14294,N_14087);
or U14700 (N_14700,N_14180,N_14481);
and U14701 (N_14701,N_14306,N_14208);
nor U14702 (N_14702,N_14019,N_14130);
nor U14703 (N_14703,N_14079,N_14417);
or U14704 (N_14704,N_14129,N_14426);
nor U14705 (N_14705,N_14445,N_14020);
or U14706 (N_14706,N_14067,N_14454);
or U14707 (N_14707,N_14096,N_14339);
nor U14708 (N_14708,N_14275,N_14323);
or U14709 (N_14709,N_14409,N_14421);
xor U14710 (N_14710,N_14047,N_14277);
nand U14711 (N_14711,N_14090,N_14405);
xnor U14712 (N_14712,N_14011,N_14227);
or U14713 (N_14713,N_14175,N_14111);
nand U14714 (N_14714,N_14232,N_14469);
nand U14715 (N_14715,N_14468,N_14015);
nor U14716 (N_14716,N_14085,N_14171);
nor U14717 (N_14717,N_14237,N_14052);
nand U14718 (N_14718,N_14371,N_14105);
or U14719 (N_14719,N_14393,N_14315);
xnor U14720 (N_14720,N_14069,N_14448);
or U14721 (N_14721,N_14362,N_14018);
xnor U14722 (N_14722,N_14119,N_14390);
or U14723 (N_14723,N_14391,N_14361);
nand U14724 (N_14724,N_14474,N_14437);
and U14725 (N_14725,N_14195,N_14140);
and U14726 (N_14726,N_14222,N_14259);
nor U14727 (N_14727,N_14345,N_14482);
xnor U14728 (N_14728,N_14028,N_14106);
nand U14729 (N_14729,N_14487,N_14147);
xor U14730 (N_14730,N_14240,N_14493);
nand U14731 (N_14731,N_14246,N_14021);
and U14732 (N_14732,N_14280,N_14040);
nand U14733 (N_14733,N_14118,N_14219);
or U14734 (N_14734,N_14003,N_14092);
nand U14735 (N_14735,N_14121,N_14432);
xnor U14736 (N_14736,N_14384,N_14266);
xor U14737 (N_14737,N_14270,N_14231);
nor U14738 (N_14738,N_14379,N_14254);
nor U14739 (N_14739,N_14365,N_14436);
or U14740 (N_14740,N_14242,N_14434);
nand U14741 (N_14741,N_14312,N_14196);
or U14742 (N_14742,N_14181,N_14336);
xnor U14743 (N_14743,N_14341,N_14499);
and U14744 (N_14744,N_14420,N_14189);
and U14745 (N_14745,N_14051,N_14309);
nand U14746 (N_14746,N_14325,N_14113);
nand U14747 (N_14747,N_14423,N_14397);
and U14748 (N_14748,N_14441,N_14483);
xnor U14749 (N_14749,N_14250,N_14154);
xor U14750 (N_14750,N_14102,N_14288);
xnor U14751 (N_14751,N_14325,N_14118);
nand U14752 (N_14752,N_14152,N_14411);
and U14753 (N_14753,N_14249,N_14031);
xor U14754 (N_14754,N_14158,N_14261);
xnor U14755 (N_14755,N_14466,N_14176);
or U14756 (N_14756,N_14418,N_14178);
nor U14757 (N_14757,N_14400,N_14177);
or U14758 (N_14758,N_14047,N_14207);
nor U14759 (N_14759,N_14436,N_14110);
xor U14760 (N_14760,N_14275,N_14452);
nand U14761 (N_14761,N_14352,N_14222);
nand U14762 (N_14762,N_14373,N_14311);
and U14763 (N_14763,N_14200,N_14132);
or U14764 (N_14764,N_14438,N_14176);
nand U14765 (N_14765,N_14424,N_14339);
and U14766 (N_14766,N_14353,N_14189);
or U14767 (N_14767,N_14350,N_14124);
nor U14768 (N_14768,N_14426,N_14261);
nand U14769 (N_14769,N_14405,N_14113);
nor U14770 (N_14770,N_14200,N_14123);
or U14771 (N_14771,N_14323,N_14445);
and U14772 (N_14772,N_14420,N_14297);
or U14773 (N_14773,N_14212,N_14041);
or U14774 (N_14774,N_14052,N_14020);
or U14775 (N_14775,N_14460,N_14276);
or U14776 (N_14776,N_14287,N_14259);
and U14777 (N_14777,N_14390,N_14371);
nand U14778 (N_14778,N_14136,N_14074);
nand U14779 (N_14779,N_14485,N_14093);
and U14780 (N_14780,N_14076,N_14231);
nor U14781 (N_14781,N_14499,N_14439);
xnor U14782 (N_14782,N_14052,N_14260);
nand U14783 (N_14783,N_14283,N_14105);
and U14784 (N_14784,N_14361,N_14014);
and U14785 (N_14785,N_14130,N_14341);
nand U14786 (N_14786,N_14382,N_14112);
xnor U14787 (N_14787,N_14246,N_14430);
xor U14788 (N_14788,N_14427,N_14312);
nand U14789 (N_14789,N_14318,N_14394);
nor U14790 (N_14790,N_14066,N_14380);
xnor U14791 (N_14791,N_14333,N_14255);
nand U14792 (N_14792,N_14235,N_14388);
and U14793 (N_14793,N_14122,N_14389);
or U14794 (N_14794,N_14326,N_14038);
or U14795 (N_14795,N_14254,N_14329);
xor U14796 (N_14796,N_14160,N_14174);
or U14797 (N_14797,N_14109,N_14186);
xor U14798 (N_14798,N_14110,N_14208);
nand U14799 (N_14799,N_14418,N_14403);
xnor U14800 (N_14800,N_14177,N_14202);
nand U14801 (N_14801,N_14333,N_14179);
and U14802 (N_14802,N_14030,N_14178);
nor U14803 (N_14803,N_14191,N_14439);
nor U14804 (N_14804,N_14212,N_14374);
or U14805 (N_14805,N_14427,N_14226);
nand U14806 (N_14806,N_14138,N_14148);
xor U14807 (N_14807,N_14075,N_14200);
xor U14808 (N_14808,N_14113,N_14096);
xor U14809 (N_14809,N_14437,N_14303);
and U14810 (N_14810,N_14048,N_14419);
and U14811 (N_14811,N_14007,N_14312);
and U14812 (N_14812,N_14461,N_14133);
and U14813 (N_14813,N_14473,N_14149);
nand U14814 (N_14814,N_14294,N_14191);
nor U14815 (N_14815,N_14422,N_14028);
nand U14816 (N_14816,N_14057,N_14291);
nand U14817 (N_14817,N_14412,N_14460);
xor U14818 (N_14818,N_14002,N_14023);
and U14819 (N_14819,N_14246,N_14054);
nand U14820 (N_14820,N_14257,N_14128);
nand U14821 (N_14821,N_14274,N_14059);
and U14822 (N_14822,N_14189,N_14204);
and U14823 (N_14823,N_14294,N_14314);
nand U14824 (N_14824,N_14418,N_14188);
nand U14825 (N_14825,N_14090,N_14363);
nand U14826 (N_14826,N_14154,N_14244);
or U14827 (N_14827,N_14450,N_14268);
or U14828 (N_14828,N_14408,N_14254);
xor U14829 (N_14829,N_14231,N_14134);
xnor U14830 (N_14830,N_14296,N_14309);
xnor U14831 (N_14831,N_14171,N_14290);
xnor U14832 (N_14832,N_14006,N_14174);
and U14833 (N_14833,N_14317,N_14253);
or U14834 (N_14834,N_14282,N_14368);
nor U14835 (N_14835,N_14428,N_14467);
nand U14836 (N_14836,N_14319,N_14457);
or U14837 (N_14837,N_14168,N_14053);
nand U14838 (N_14838,N_14281,N_14019);
nor U14839 (N_14839,N_14296,N_14139);
nor U14840 (N_14840,N_14166,N_14422);
or U14841 (N_14841,N_14142,N_14419);
or U14842 (N_14842,N_14008,N_14121);
or U14843 (N_14843,N_14434,N_14340);
and U14844 (N_14844,N_14285,N_14078);
nor U14845 (N_14845,N_14092,N_14329);
xor U14846 (N_14846,N_14058,N_14451);
xor U14847 (N_14847,N_14257,N_14470);
nand U14848 (N_14848,N_14380,N_14170);
nand U14849 (N_14849,N_14106,N_14255);
nand U14850 (N_14850,N_14198,N_14038);
xor U14851 (N_14851,N_14385,N_14218);
xnor U14852 (N_14852,N_14268,N_14237);
or U14853 (N_14853,N_14193,N_14072);
and U14854 (N_14854,N_14082,N_14024);
or U14855 (N_14855,N_14478,N_14462);
nand U14856 (N_14856,N_14449,N_14447);
nand U14857 (N_14857,N_14073,N_14134);
or U14858 (N_14858,N_14359,N_14087);
nand U14859 (N_14859,N_14415,N_14311);
nor U14860 (N_14860,N_14259,N_14306);
nor U14861 (N_14861,N_14314,N_14040);
xnor U14862 (N_14862,N_14297,N_14322);
and U14863 (N_14863,N_14199,N_14460);
or U14864 (N_14864,N_14443,N_14328);
and U14865 (N_14865,N_14467,N_14076);
xor U14866 (N_14866,N_14129,N_14252);
nand U14867 (N_14867,N_14168,N_14450);
nand U14868 (N_14868,N_14327,N_14172);
and U14869 (N_14869,N_14283,N_14221);
or U14870 (N_14870,N_14392,N_14376);
and U14871 (N_14871,N_14063,N_14051);
or U14872 (N_14872,N_14446,N_14008);
nand U14873 (N_14873,N_14430,N_14053);
nor U14874 (N_14874,N_14194,N_14498);
or U14875 (N_14875,N_14038,N_14114);
nor U14876 (N_14876,N_14261,N_14280);
nor U14877 (N_14877,N_14064,N_14228);
nor U14878 (N_14878,N_14049,N_14285);
or U14879 (N_14879,N_14291,N_14118);
nand U14880 (N_14880,N_14344,N_14149);
or U14881 (N_14881,N_14412,N_14225);
nand U14882 (N_14882,N_14330,N_14054);
nand U14883 (N_14883,N_14467,N_14305);
nor U14884 (N_14884,N_14417,N_14473);
xor U14885 (N_14885,N_14429,N_14489);
or U14886 (N_14886,N_14083,N_14213);
xor U14887 (N_14887,N_14345,N_14267);
nor U14888 (N_14888,N_14038,N_14280);
nor U14889 (N_14889,N_14414,N_14109);
or U14890 (N_14890,N_14386,N_14000);
or U14891 (N_14891,N_14060,N_14410);
nand U14892 (N_14892,N_14448,N_14279);
xor U14893 (N_14893,N_14395,N_14470);
nor U14894 (N_14894,N_14118,N_14054);
nand U14895 (N_14895,N_14068,N_14226);
nand U14896 (N_14896,N_14349,N_14423);
and U14897 (N_14897,N_14156,N_14104);
nand U14898 (N_14898,N_14449,N_14199);
or U14899 (N_14899,N_14219,N_14333);
and U14900 (N_14900,N_14252,N_14485);
xor U14901 (N_14901,N_14041,N_14351);
nand U14902 (N_14902,N_14387,N_14094);
nand U14903 (N_14903,N_14183,N_14280);
or U14904 (N_14904,N_14325,N_14114);
xor U14905 (N_14905,N_14243,N_14253);
or U14906 (N_14906,N_14065,N_14119);
xor U14907 (N_14907,N_14336,N_14443);
xnor U14908 (N_14908,N_14183,N_14043);
nand U14909 (N_14909,N_14384,N_14248);
nor U14910 (N_14910,N_14391,N_14052);
xnor U14911 (N_14911,N_14168,N_14285);
or U14912 (N_14912,N_14447,N_14097);
nor U14913 (N_14913,N_14104,N_14125);
or U14914 (N_14914,N_14214,N_14406);
xnor U14915 (N_14915,N_14153,N_14106);
xnor U14916 (N_14916,N_14287,N_14115);
or U14917 (N_14917,N_14323,N_14053);
xor U14918 (N_14918,N_14070,N_14134);
nand U14919 (N_14919,N_14002,N_14014);
nor U14920 (N_14920,N_14330,N_14412);
xor U14921 (N_14921,N_14385,N_14220);
or U14922 (N_14922,N_14104,N_14128);
nor U14923 (N_14923,N_14224,N_14262);
nand U14924 (N_14924,N_14364,N_14100);
or U14925 (N_14925,N_14288,N_14138);
xnor U14926 (N_14926,N_14134,N_14232);
or U14927 (N_14927,N_14090,N_14373);
nand U14928 (N_14928,N_14443,N_14244);
nor U14929 (N_14929,N_14186,N_14001);
nand U14930 (N_14930,N_14087,N_14042);
nor U14931 (N_14931,N_14471,N_14244);
or U14932 (N_14932,N_14060,N_14431);
or U14933 (N_14933,N_14230,N_14310);
nand U14934 (N_14934,N_14133,N_14400);
and U14935 (N_14935,N_14321,N_14485);
xor U14936 (N_14936,N_14295,N_14342);
nand U14937 (N_14937,N_14337,N_14211);
nor U14938 (N_14938,N_14459,N_14424);
nand U14939 (N_14939,N_14313,N_14286);
nor U14940 (N_14940,N_14231,N_14113);
and U14941 (N_14941,N_14054,N_14236);
or U14942 (N_14942,N_14119,N_14024);
and U14943 (N_14943,N_14206,N_14201);
xor U14944 (N_14944,N_14154,N_14036);
nand U14945 (N_14945,N_14249,N_14167);
nor U14946 (N_14946,N_14059,N_14266);
or U14947 (N_14947,N_14466,N_14222);
nand U14948 (N_14948,N_14078,N_14294);
and U14949 (N_14949,N_14349,N_14216);
nand U14950 (N_14950,N_14293,N_14049);
and U14951 (N_14951,N_14297,N_14112);
and U14952 (N_14952,N_14413,N_14484);
xnor U14953 (N_14953,N_14077,N_14306);
xor U14954 (N_14954,N_14034,N_14400);
and U14955 (N_14955,N_14007,N_14038);
xnor U14956 (N_14956,N_14186,N_14484);
and U14957 (N_14957,N_14323,N_14134);
nand U14958 (N_14958,N_14104,N_14319);
and U14959 (N_14959,N_14118,N_14094);
and U14960 (N_14960,N_14277,N_14351);
and U14961 (N_14961,N_14244,N_14027);
and U14962 (N_14962,N_14092,N_14210);
nand U14963 (N_14963,N_14143,N_14346);
or U14964 (N_14964,N_14137,N_14436);
and U14965 (N_14965,N_14021,N_14278);
or U14966 (N_14966,N_14104,N_14121);
nor U14967 (N_14967,N_14271,N_14016);
nor U14968 (N_14968,N_14432,N_14494);
nand U14969 (N_14969,N_14315,N_14349);
or U14970 (N_14970,N_14220,N_14225);
nand U14971 (N_14971,N_14396,N_14141);
nand U14972 (N_14972,N_14193,N_14292);
nor U14973 (N_14973,N_14027,N_14386);
or U14974 (N_14974,N_14052,N_14481);
xor U14975 (N_14975,N_14388,N_14042);
and U14976 (N_14976,N_14082,N_14395);
xnor U14977 (N_14977,N_14353,N_14298);
and U14978 (N_14978,N_14435,N_14349);
or U14979 (N_14979,N_14218,N_14173);
xnor U14980 (N_14980,N_14497,N_14318);
nor U14981 (N_14981,N_14005,N_14333);
xor U14982 (N_14982,N_14170,N_14207);
xnor U14983 (N_14983,N_14160,N_14436);
nor U14984 (N_14984,N_14277,N_14280);
or U14985 (N_14985,N_14123,N_14037);
xor U14986 (N_14986,N_14149,N_14293);
nand U14987 (N_14987,N_14133,N_14237);
or U14988 (N_14988,N_14471,N_14192);
and U14989 (N_14989,N_14011,N_14359);
and U14990 (N_14990,N_14432,N_14034);
or U14991 (N_14991,N_14459,N_14384);
xnor U14992 (N_14992,N_14051,N_14399);
and U14993 (N_14993,N_14000,N_14099);
nand U14994 (N_14994,N_14177,N_14390);
xor U14995 (N_14995,N_14396,N_14151);
and U14996 (N_14996,N_14014,N_14111);
xnor U14997 (N_14997,N_14318,N_14426);
or U14998 (N_14998,N_14044,N_14183);
nand U14999 (N_14999,N_14279,N_14109);
xnor UO_0 (O_0,N_14624,N_14817);
xor UO_1 (O_1,N_14719,N_14567);
nand UO_2 (O_2,N_14922,N_14855);
or UO_3 (O_3,N_14533,N_14956);
xnor UO_4 (O_4,N_14772,N_14958);
xnor UO_5 (O_5,N_14711,N_14803);
xor UO_6 (O_6,N_14955,N_14968);
nor UO_7 (O_7,N_14693,N_14739);
nor UO_8 (O_8,N_14806,N_14540);
nor UO_9 (O_9,N_14561,N_14577);
or UO_10 (O_10,N_14786,N_14578);
nand UO_11 (O_11,N_14977,N_14814);
nor UO_12 (O_12,N_14811,N_14797);
nor UO_13 (O_13,N_14813,N_14747);
or UO_14 (O_14,N_14733,N_14667);
and UO_15 (O_15,N_14708,N_14685);
or UO_16 (O_16,N_14886,N_14908);
or UO_17 (O_17,N_14879,N_14776);
and UO_18 (O_18,N_14669,N_14544);
or UO_19 (O_19,N_14530,N_14759);
nor UO_20 (O_20,N_14998,N_14558);
nor UO_21 (O_21,N_14563,N_14898);
or UO_22 (O_22,N_14593,N_14628);
nor UO_23 (O_23,N_14868,N_14573);
nand UO_24 (O_24,N_14553,N_14700);
nand UO_25 (O_25,N_14662,N_14534);
or UO_26 (O_26,N_14909,N_14694);
nor UO_27 (O_27,N_14736,N_14612);
or UO_28 (O_28,N_14600,N_14653);
xnor UO_29 (O_29,N_14659,N_14867);
xnor UO_30 (O_30,N_14761,N_14636);
nor UO_31 (O_31,N_14945,N_14570);
nor UO_32 (O_32,N_14718,N_14695);
nor UO_33 (O_33,N_14670,N_14876);
xnor UO_34 (O_34,N_14793,N_14728);
nand UO_35 (O_35,N_14903,N_14760);
xor UO_36 (O_36,N_14676,N_14928);
or UO_37 (O_37,N_14944,N_14651);
and UO_38 (O_38,N_14980,N_14596);
and UO_39 (O_39,N_14774,N_14629);
or UO_40 (O_40,N_14940,N_14508);
xor UO_41 (O_41,N_14746,N_14587);
xnor UO_42 (O_42,N_14845,N_14643);
nand UO_43 (O_43,N_14788,N_14801);
or UO_44 (O_44,N_14604,N_14602);
nor UO_45 (O_45,N_14981,N_14934);
xor UO_46 (O_46,N_14583,N_14820);
xor UO_47 (O_47,N_14796,N_14610);
xor UO_48 (O_48,N_14559,N_14568);
and UO_49 (O_49,N_14519,N_14531);
nand UO_50 (O_50,N_14619,N_14509);
and UO_51 (O_51,N_14634,N_14979);
and UO_52 (O_52,N_14557,N_14905);
or UO_53 (O_53,N_14848,N_14782);
or UO_54 (O_54,N_14875,N_14915);
nand UO_55 (O_55,N_14750,N_14710);
or UO_56 (O_56,N_14847,N_14836);
or UO_57 (O_57,N_14818,N_14975);
xnor UO_58 (O_58,N_14650,N_14951);
and UO_59 (O_59,N_14884,N_14841);
and UO_60 (O_60,N_14660,N_14989);
or UO_61 (O_61,N_14936,N_14625);
nor UO_62 (O_62,N_14792,N_14812);
and UO_63 (O_63,N_14978,N_14916);
nand UO_64 (O_64,N_14627,N_14698);
nand UO_65 (O_65,N_14686,N_14732);
and UO_66 (O_66,N_14894,N_14882);
nand UO_67 (O_67,N_14678,N_14642);
nand UO_68 (O_68,N_14973,N_14819);
nand UO_69 (O_69,N_14551,N_14713);
nor UO_70 (O_70,N_14893,N_14861);
or UO_71 (O_71,N_14688,N_14832);
and UO_72 (O_72,N_14517,N_14983);
xnor UO_73 (O_73,N_14588,N_14857);
and UO_74 (O_74,N_14539,N_14512);
nand UO_75 (O_75,N_14749,N_14885);
xnor UO_76 (O_76,N_14807,N_14598);
nand UO_77 (O_77,N_14703,N_14769);
xor UO_78 (O_78,N_14917,N_14959);
and UO_79 (O_79,N_14644,N_14741);
xor UO_80 (O_80,N_14550,N_14631);
and UO_81 (O_81,N_14873,N_14946);
xor UO_82 (O_82,N_14520,N_14535);
and UO_83 (O_83,N_14640,N_14783);
and UO_84 (O_84,N_14869,N_14564);
and UO_85 (O_85,N_14691,N_14816);
and UO_86 (O_86,N_14717,N_14681);
or UO_87 (O_87,N_14649,N_14993);
nand UO_88 (O_88,N_14860,N_14687);
nor UO_89 (O_89,N_14763,N_14548);
nor UO_90 (O_90,N_14756,N_14555);
nand UO_91 (O_91,N_14566,N_14589);
xor UO_92 (O_92,N_14896,N_14815);
or UO_93 (O_93,N_14501,N_14890);
and UO_94 (O_94,N_14706,N_14852);
and UO_95 (O_95,N_14726,N_14969);
nand UO_96 (O_96,N_14822,N_14584);
or UO_97 (O_97,N_14972,N_14825);
nand UO_98 (O_98,N_14709,N_14918);
xnor UO_99 (O_99,N_14712,N_14731);
nand UO_100 (O_100,N_14844,N_14954);
or UO_101 (O_101,N_14984,N_14872);
xnor UO_102 (O_102,N_14779,N_14647);
xnor UO_103 (O_103,N_14919,N_14576);
xor UO_104 (O_104,N_14692,N_14672);
nand UO_105 (O_105,N_14597,N_14974);
nand UO_106 (O_106,N_14805,N_14716);
xor UO_107 (O_107,N_14790,N_14633);
or UO_108 (O_108,N_14605,N_14727);
or UO_109 (O_109,N_14843,N_14652);
nand UO_110 (O_110,N_14802,N_14527);
xor UO_111 (O_111,N_14938,N_14536);
xor UO_112 (O_112,N_14525,N_14673);
xor UO_113 (O_113,N_14547,N_14949);
nand UO_114 (O_114,N_14787,N_14863);
nand UO_115 (O_115,N_14521,N_14941);
or UO_116 (O_116,N_14912,N_14901);
xnor UO_117 (O_117,N_14630,N_14514);
nand UO_118 (O_118,N_14985,N_14966);
or UO_119 (O_119,N_14757,N_14823);
and UO_120 (O_120,N_14800,N_14538);
and UO_121 (O_121,N_14730,N_14794);
xnor UO_122 (O_122,N_14827,N_14745);
nand UO_123 (O_123,N_14734,N_14671);
xnor UO_124 (O_124,N_14930,N_14777);
and UO_125 (O_125,N_14795,N_14632);
xnor UO_126 (O_126,N_14947,N_14744);
nor UO_127 (O_127,N_14524,N_14932);
nor UO_128 (O_128,N_14682,N_14995);
nand UO_129 (O_129,N_14614,N_14674);
xnor UO_130 (O_130,N_14755,N_14690);
nor UO_131 (O_131,N_14645,N_14939);
nor UO_132 (O_132,N_14952,N_14856);
and UO_133 (O_133,N_14615,N_14996);
xor UO_134 (O_134,N_14775,N_14654);
nor UO_135 (O_135,N_14586,N_14715);
or UO_136 (O_136,N_14556,N_14616);
nor UO_137 (O_137,N_14943,N_14961);
or UO_138 (O_138,N_14664,N_14925);
or UO_139 (O_139,N_14720,N_14611);
xor UO_140 (O_140,N_14921,N_14924);
nor UO_141 (O_141,N_14663,N_14565);
or UO_142 (O_142,N_14765,N_14665);
nand UO_143 (O_143,N_14906,N_14575);
nor UO_144 (O_144,N_14809,N_14877);
nor UO_145 (O_145,N_14862,N_14851);
nor UO_146 (O_146,N_14997,N_14976);
and UO_147 (O_147,N_14988,N_14714);
xnor UO_148 (O_148,N_14502,N_14609);
or UO_149 (O_149,N_14791,N_14854);
xnor UO_150 (O_150,N_14962,N_14560);
and UO_151 (O_151,N_14842,N_14829);
nor UO_152 (O_152,N_14721,N_14735);
nand UO_153 (O_153,N_14658,N_14840);
or UO_154 (O_154,N_14920,N_14724);
and UO_155 (O_155,N_14613,N_14680);
xor UO_156 (O_156,N_14913,N_14641);
nor UO_157 (O_157,N_14964,N_14684);
nand UO_158 (O_158,N_14683,N_14880);
or UO_159 (O_159,N_14766,N_14837);
xor UO_160 (O_160,N_14931,N_14804);
or UO_161 (O_161,N_14963,N_14957);
xor UO_162 (O_162,N_14503,N_14870);
xnor UO_163 (O_163,N_14655,N_14500);
nor UO_164 (O_164,N_14639,N_14617);
or UO_165 (O_165,N_14626,N_14743);
nor UO_166 (O_166,N_14748,N_14881);
nor UO_167 (O_167,N_14824,N_14883);
xor UO_168 (O_168,N_14689,N_14897);
and UO_169 (O_169,N_14850,N_14781);
nand UO_170 (O_170,N_14637,N_14768);
and UO_171 (O_171,N_14780,N_14579);
and UO_172 (O_172,N_14742,N_14994);
and UO_173 (O_173,N_14953,N_14526);
and UO_174 (O_174,N_14937,N_14661);
nor UO_175 (O_175,N_14608,N_14835);
nor UO_176 (O_176,N_14878,N_14833);
nor UO_177 (O_177,N_14722,N_14859);
or UO_178 (O_178,N_14986,N_14960);
or UO_179 (O_179,N_14554,N_14668);
xnor UO_180 (O_180,N_14758,N_14935);
nor UO_181 (O_181,N_14895,N_14888);
xnor UO_182 (O_182,N_14866,N_14942);
or UO_183 (O_183,N_14592,N_14826);
nand UO_184 (O_184,N_14571,N_14623);
xor UO_185 (O_185,N_14967,N_14808);
nor UO_186 (O_186,N_14707,N_14914);
and UO_187 (O_187,N_14523,N_14762);
or UO_188 (O_188,N_14965,N_14549);
and UO_189 (O_189,N_14999,N_14911);
nor UO_190 (O_190,N_14853,N_14926);
nand UO_191 (O_191,N_14927,N_14821);
xor UO_192 (O_192,N_14849,N_14545);
nor UO_193 (O_193,N_14590,N_14552);
xnor UO_194 (O_194,N_14574,N_14987);
nor UO_195 (O_195,N_14569,N_14751);
or UO_196 (O_196,N_14784,N_14839);
nand UO_197 (O_197,N_14799,N_14622);
nand UO_198 (O_198,N_14599,N_14770);
or UO_199 (O_199,N_14785,N_14831);
and UO_200 (O_200,N_14887,N_14991);
or UO_201 (O_201,N_14516,N_14789);
and UO_202 (O_202,N_14607,N_14594);
or UO_203 (O_203,N_14675,N_14740);
nand UO_204 (O_204,N_14874,N_14992);
and UO_205 (O_205,N_14696,N_14892);
and UO_206 (O_206,N_14902,N_14725);
nand UO_207 (O_207,N_14572,N_14864);
nand UO_208 (O_208,N_14738,N_14618);
xor UO_209 (O_209,N_14657,N_14606);
nand UO_210 (O_210,N_14679,N_14506);
nor UO_211 (O_211,N_14513,N_14522);
or UO_212 (O_212,N_14562,N_14846);
nand UO_213 (O_213,N_14798,N_14889);
and UO_214 (O_214,N_14697,N_14933);
xor UO_215 (O_215,N_14754,N_14971);
nor UO_216 (O_216,N_14858,N_14603);
and UO_217 (O_217,N_14699,N_14543);
and UO_218 (O_218,N_14990,N_14771);
nor UO_219 (O_219,N_14648,N_14810);
nor UO_220 (O_220,N_14729,N_14891);
and UO_221 (O_221,N_14899,N_14595);
and UO_222 (O_222,N_14830,N_14542);
xnor UO_223 (O_223,N_14529,N_14834);
nand UO_224 (O_224,N_14532,N_14515);
or UO_225 (O_225,N_14511,N_14923);
xor UO_226 (O_226,N_14646,N_14982);
xnor UO_227 (O_227,N_14970,N_14580);
nand UO_228 (O_228,N_14737,N_14581);
xnor UO_229 (O_229,N_14900,N_14518);
xor UO_230 (O_230,N_14752,N_14865);
nand UO_231 (O_231,N_14764,N_14620);
nand UO_232 (O_232,N_14767,N_14546);
and UO_233 (O_233,N_14541,N_14910);
nand UO_234 (O_234,N_14773,N_14828);
or UO_235 (O_235,N_14582,N_14753);
xor UO_236 (O_236,N_14537,N_14621);
nand UO_237 (O_237,N_14871,N_14838);
nor UO_238 (O_238,N_14638,N_14635);
and UO_239 (O_239,N_14504,N_14677);
xor UO_240 (O_240,N_14666,N_14904);
nor UO_241 (O_241,N_14528,N_14929);
xnor UO_242 (O_242,N_14510,N_14591);
nand UO_243 (O_243,N_14907,N_14585);
nor UO_244 (O_244,N_14702,N_14778);
nand UO_245 (O_245,N_14948,N_14704);
xnor UO_246 (O_246,N_14701,N_14507);
or UO_247 (O_247,N_14505,N_14656);
and UO_248 (O_248,N_14705,N_14601);
nor UO_249 (O_249,N_14723,N_14950);
and UO_250 (O_250,N_14634,N_14747);
or UO_251 (O_251,N_14640,N_14851);
or UO_252 (O_252,N_14594,N_14763);
nor UO_253 (O_253,N_14558,N_14795);
nor UO_254 (O_254,N_14774,N_14900);
nand UO_255 (O_255,N_14886,N_14775);
xor UO_256 (O_256,N_14771,N_14533);
nand UO_257 (O_257,N_14704,N_14533);
nor UO_258 (O_258,N_14947,N_14543);
nand UO_259 (O_259,N_14530,N_14599);
and UO_260 (O_260,N_14948,N_14586);
nor UO_261 (O_261,N_14646,N_14659);
xnor UO_262 (O_262,N_14529,N_14932);
and UO_263 (O_263,N_14933,N_14782);
xnor UO_264 (O_264,N_14640,N_14901);
nor UO_265 (O_265,N_14855,N_14729);
xnor UO_266 (O_266,N_14584,N_14536);
xor UO_267 (O_267,N_14568,N_14766);
and UO_268 (O_268,N_14615,N_14951);
or UO_269 (O_269,N_14961,N_14551);
nor UO_270 (O_270,N_14877,N_14945);
xor UO_271 (O_271,N_14843,N_14930);
xnor UO_272 (O_272,N_14963,N_14710);
nor UO_273 (O_273,N_14806,N_14653);
nand UO_274 (O_274,N_14573,N_14733);
nor UO_275 (O_275,N_14904,N_14794);
nand UO_276 (O_276,N_14805,N_14976);
nand UO_277 (O_277,N_14770,N_14581);
xnor UO_278 (O_278,N_14667,N_14565);
nand UO_279 (O_279,N_14934,N_14784);
nor UO_280 (O_280,N_14841,N_14865);
and UO_281 (O_281,N_14619,N_14714);
xnor UO_282 (O_282,N_14824,N_14512);
and UO_283 (O_283,N_14525,N_14924);
nor UO_284 (O_284,N_14616,N_14976);
xor UO_285 (O_285,N_14610,N_14518);
or UO_286 (O_286,N_14615,N_14610);
or UO_287 (O_287,N_14569,N_14866);
nor UO_288 (O_288,N_14880,N_14915);
nand UO_289 (O_289,N_14640,N_14658);
nor UO_290 (O_290,N_14629,N_14756);
and UO_291 (O_291,N_14538,N_14663);
xor UO_292 (O_292,N_14956,N_14687);
nor UO_293 (O_293,N_14955,N_14548);
xor UO_294 (O_294,N_14918,N_14913);
or UO_295 (O_295,N_14613,N_14619);
nand UO_296 (O_296,N_14794,N_14588);
or UO_297 (O_297,N_14693,N_14746);
nand UO_298 (O_298,N_14957,N_14935);
nand UO_299 (O_299,N_14953,N_14733);
nand UO_300 (O_300,N_14869,N_14673);
xor UO_301 (O_301,N_14853,N_14613);
and UO_302 (O_302,N_14938,N_14604);
and UO_303 (O_303,N_14974,N_14563);
and UO_304 (O_304,N_14814,N_14876);
or UO_305 (O_305,N_14673,N_14875);
and UO_306 (O_306,N_14914,N_14615);
nand UO_307 (O_307,N_14863,N_14875);
or UO_308 (O_308,N_14900,N_14911);
and UO_309 (O_309,N_14555,N_14698);
nand UO_310 (O_310,N_14904,N_14844);
nand UO_311 (O_311,N_14807,N_14623);
or UO_312 (O_312,N_14577,N_14755);
xnor UO_313 (O_313,N_14803,N_14983);
xor UO_314 (O_314,N_14837,N_14689);
nor UO_315 (O_315,N_14823,N_14652);
xnor UO_316 (O_316,N_14639,N_14696);
xnor UO_317 (O_317,N_14761,N_14871);
nor UO_318 (O_318,N_14727,N_14629);
and UO_319 (O_319,N_14916,N_14932);
and UO_320 (O_320,N_14887,N_14861);
or UO_321 (O_321,N_14753,N_14602);
nand UO_322 (O_322,N_14873,N_14992);
xor UO_323 (O_323,N_14711,N_14940);
nand UO_324 (O_324,N_14923,N_14535);
or UO_325 (O_325,N_14695,N_14624);
or UO_326 (O_326,N_14900,N_14528);
nor UO_327 (O_327,N_14582,N_14948);
and UO_328 (O_328,N_14984,N_14970);
nand UO_329 (O_329,N_14741,N_14945);
and UO_330 (O_330,N_14578,N_14952);
and UO_331 (O_331,N_14683,N_14873);
nand UO_332 (O_332,N_14859,N_14660);
xor UO_333 (O_333,N_14652,N_14513);
nor UO_334 (O_334,N_14892,N_14627);
xor UO_335 (O_335,N_14617,N_14922);
nor UO_336 (O_336,N_14854,N_14531);
and UO_337 (O_337,N_14899,N_14995);
nand UO_338 (O_338,N_14766,N_14989);
or UO_339 (O_339,N_14875,N_14670);
nand UO_340 (O_340,N_14808,N_14599);
and UO_341 (O_341,N_14937,N_14972);
and UO_342 (O_342,N_14767,N_14979);
nor UO_343 (O_343,N_14941,N_14827);
nor UO_344 (O_344,N_14506,N_14984);
and UO_345 (O_345,N_14990,N_14781);
or UO_346 (O_346,N_14939,N_14800);
xor UO_347 (O_347,N_14702,N_14875);
nor UO_348 (O_348,N_14821,N_14973);
nand UO_349 (O_349,N_14939,N_14524);
xnor UO_350 (O_350,N_14544,N_14667);
nor UO_351 (O_351,N_14871,N_14583);
or UO_352 (O_352,N_14809,N_14843);
nor UO_353 (O_353,N_14780,N_14854);
xor UO_354 (O_354,N_14920,N_14533);
and UO_355 (O_355,N_14637,N_14994);
nand UO_356 (O_356,N_14922,N_14570);
nor UO_357 (O_357,N_14532,N_14924);
and UO_358 (O_358,N_14728,N_14715);
and UO_359 (O_359,N_14720,N_14696);
or UO_360 (O_360,N_14505,N_14890);
and UO_361 (O_361,N_14763,N_14838);
or UO_362 (O_362,N_14513,N_14964);
xnor UO_363 (O_363,N_14979,N_14994);
xor UO_364 (O_364,N_14729,N_14582);
nand UO_365 (O_365,N_14835,N_14632);
or UO_366 (O_366,N_14796,N_14573);
xor UO_367 (O_367,N_14905,N_14722);
and UO_368 (O_368,N_14830,N_14531);
nor UO_369 (O_369,N_14981,N_14682);
nor UO_370 (O_370,N_14783,N_14572);
nor UO_371 (O_371,N_14625,N_14627);
and UO_372 (O_372,N_14624,N_14851);
nand UO_373 (O_373,N_14656,N_14890);
and UO_374 (O_374,N_14811,N_14608);
or UO_375 (O_375,N_14946,N_14805);
and UO_376 (O_376,N_14715,N_14544);
xor UO_377 (O_377,N_14933,N_14924);
xor UO_378 (O_378,N_14978,N_14668);
xnor UO_379 (O_379,N_14817,N_14639);
or UO_380 (O_380,N_14939,N_14820);
nor UO_381 (O_381,N_14572,N_14957);
or UO_382 (O_382,N_14761,N_14991);
xor UO_383 (O_383,N_14838,N_14750);
or UO_384 (O_384,N_14830,N_14689);
or UO_385 (O_385,N_14683,N_14588);
nor UO_386 (O_386,N_14615,N_14680);
and UO_387 (O_387,N_14657,N_14690);
or UO_388 (O_388,N_14646,N_14719);
nand UO_389 (O_389,N_14554,N_14895);
nor UO_390 (O_390,N_14743,N_14994);
nor UO_391 (O_391,N_14879,N_14510);
xnor UO_392 (O_392,N_14516,N_14731);
and UO_393 (O_393,N_14576,N_14624);
or UO_394 (O_394,N_14905,N_14822);
or UO_395 (O_395,N_14856,N_14899);
nor UO_396 (O_396,N_14697,N_14559);
nor UO_397 (O_397,N_14648,N_14686);
nor UO_398 (O_398,N_14753,N_14785);
and UO_399 (O_399,N_14601,N_14980);
and UO_400 (O_400,N_14517,N_14660);
xnor UO_401 (O_401,N_14882,N_14555);
nor UO_402 (O_402,N_14552,N_14991);
or UO_403 (O_403,N_14796,N_14664);
xnor UO_404 (O_404,N_14645,N_14609);
or UO_405 (O_405,N_14619,N_14598);
or UO_406 (O_406,N_14810,N_14741);
nand UO_407 (O_407,N_14958,N_14816);
nor UO_408 (O_408,N_14835,N_14504);
nor UO_409 (O_409,N_14837,N_14886);
or UO_410 (O_410,N_14980,N_14893);
nor UO_411 (O_411,N_14885,N_14648);
xnor UO_412 (O_412,N_14701,N_14677);
xnor UO_413 (O_413,N_14993,N_14956);
or UO_414 (O_414,N_14951,N_14580);
and UO_415 (O_415,N_14716,N_14512);
nand UO_416 (O_416,N_14657,N_14703);
nand UO_417 (O_417,N_14718,N_14977);
and UO_418 (O_418,N_14637,N_14640);
nand UO_419 (O_419,N_14532,N_14794);
nand UO_420 (O_420,N_14823,N_14732);
nor UO_421 (O_421,N_14513,N_14647);
nand UO_422 (O_422,N_14747,N_14624);
nor UO_423 (O_423,N_14572,N_14827);
and UO_424 (O_424,N_14819,N_14633);
nor UO_425 (O_425,N_14903,N_14840);
xnor UO_426 (O_426,N_14990,N_14550);
and UO_427 (O_427,N_14861,N_14739);
nand UO_428 (O_428,N_14947,N_14567);
nor UO_429 (O_429,N_14578,N_14723);
xor UO_430 (O_430,N_14852,N_14787);
nand UO_431 (O_431,N_14553,N_14646);
nand UO_432 (O_432,N_14901,N_14672);
or UO_433 (O_433,N_14549,N_14544);
or UO_434 (O_434,N_14714,N_14925);
and UO_435 (O_435,N_14917,N_14997);
nand UO_436 (O_436,N_14959,N_14730);
or UO_437 (O_437,N_14938,N_14570);
nor UO_438 (O_438,N_14583,N_14978);
nand UO_439 (O_439,N_14861,N_14886);
xnor UO_440 (O_440,N_14718,N_14689);
nand UO_441 (O_441,N_14822,N_14716);
or UO_442 (O_442,N_14579,N_14825);
nand UO_443 (O_443,N_14673,N_14893);
nor UO_444 (O_444,N_14531,N_14683);
nor UO_445 (O_445,N_14904,N_14618);
nor UO_446 (O_446,N_14768,N_14981);
nor UO_447 (O_447,N_14575,N_14900);
or UO_448 (O_448,N_14717,N_14797);
nand UO_449 (O_449,N_14549,N_14920);
nor UO_450 (O_450,N_14673,N_14666);
xnor UO_451 (O_451,N_14942,N_14934);
nor UO_452 (O_452,N_14708,N_14789);
xor UO_453 (O_453,N_14636,N_14728);
or UO_454 (O_454,N_14550,N_14972);
xor UO_455 (O_455,N_14504,N_14596);
or UO_456 (O_456,N_14646,N_14718);
nor UO_457 (O_457,N_14642,N_14739);
nor UO_458 (O_458,N_14631,N_14748);
xnor UO_459 (O_459,N_14546,N_14647);
nor UO_460 (O_460,N_14799,N_14567);
nor UO_461 (O_461,N_14810,N_14793);
or UO_462 (O_462,N_14762,N_14771);
xor UO_463 (O_463,N_14956,N_14826);
xnor UO_464 (O_464,N_14856,N_14617);
or UO_465 (O_465,N_14841,N_14580);
and UO_466 (O_466,N_14859,N_14820);
and UO_467 (O_467,N_14817,N_14536);
or UO_468 (O_468,N_14948,N_14806);
xnor UO_469 (O_469,N_14871,N_14599);
nand UO_470 (O_470,N_14801,N_14793);
xor UO_471 (O_471,N_14864,N_14973);
nor UO_472 (O_472,N_14729,N_14954);
xnor UO_473 (O_473,N_14740,N_14814);
nand UO_474 (O_474,N_14827,N_14934);
and UO_475 (O_475,N_14531,N_14898);
nor UO_476 (O_476,N_14842,N_14738);
xor UO_477 (O_477,N_14870,N_14616);
nor UO_478 (O_478,N_14594,N_14855);
xor UO_479 (O_479,N_14933,N_14555);
and UO_480 (O_480,N_14937,N_14648);
nor UO_481 (O_481,N_14918,N_14799);
and UO_482 (O_482,N_14797,N_14861);
nand UO_483 (O_483,N_14661,N_14779);
nor UO_484 (O_484,N_14557,N_14850);
nand UO_485 (O_485,N_14608,N_14831);
nand UO_486 (O_486,N_14782,N_14767);
and UO_487 (O_487,N_14923,N_14612);
or UO_488 (O_488,N_14862,N_14670);
xor UO_489 (O_489,N_14582,N_14747);
xnor UO_490 (O_490,N_14632,N_14803);
nor UO_491 (O_491,N_14669,N_14545);
and UO_492 (O_492,N_14566,N_14957);
xnor UO_493 (O_493,N_14787,N_14537);
and UO_494 (O_494,N_14670,N_14691);
nand UO_495 (O_495,N_14831,N_14589);
and UO_496 (O_496,N_14535,N_14551);
xor UO_497 (O_497,N_14657,N_14541);
xnor UO_498 (O_498,N_14542,N_14622);
nand UO_499 (O_499,N_14794,N_14744);
or UO_500 (O_500,N_14692,N_14675);
xnor UO_501 (O_501,N_14639,N_14678);
nor UO_502 (O_502,N_14627,N_14897);
or UO_503 (O_503,N_14699,N_14645);
nor UO_504 (O_504,N_14636,N_14660);
or UO_505 (O_505,N_14770,N_14631);
nor UO_506 (O_506,N_14681,N_14886);
xnor UO_507 (O_507,N_14544,N_14911);
or UO_508 (O_508,N_14987,N_14570);
or UO_509 (O_509,N_14857,N_14778);
and UO_510 (O_510,N_14888,N_14660);
or UO_511 (O_511,N_14908,N_14602);
nor UO_512 (O_512,N_14792,N_14590);
and UO_513 (O_513,N_14881,N_14587);
or UO_514 (O_514,N_14500,N_14641);
xnor UO_515 (O_515,N_14931,N_14823);
and UO_516 (O_516,N_14824,N_14987);
or UO_517 (O_517,N_14562,N_14830);
nor UO_518 (O_518,N_14974,N_14692);
nand UO_519 (O_519,N_14511,N_14760);
nor UO_520 (O_520,N_14563,N_14512);
and UO_521 (O_521,N_14631,N_14858);
or UO_522 (O_522,N_14515,N_14536);
nand UO_523 (O_523,N_14958,N_14972);
xor UO_524 (O_524,N_14799,N_14627);
xor UO_525 (O_525,N_14712,N_14634);
nand UO_526 (O_526,N_14823,N_14621);
and UO_527 (O_527,N_14802,N_14509);
xnor UO_528 (O_528,N_14621,N_14832);
nor UO_529 (O_529,N_14784,N_14642);
or UO_530 (O_530,N_14929,N_14934);
and UO_531 (O_531,N_14756,N_14713);
and UO_532 (O_532,N_14815,N_14777);
and UO_533 (O_533,N_14662,N_14894);
nand UO_534 (O_534,N_14604,N_14969);
xor UO_535 (O_535,N_14503,N_14527);
nand UO_536 (O_536,N_14781,N_14992);
xor UO_537 (O_537,N_14813,N_14528);
and UO_538 (O_538,N_14629,N_14544);
and UO_539 (O_539,N_14769,N_14693);
and UO_540 (O_540,N_14753,N_14898);
nand UO_541 (O_541,N_14615,N_14608);
or UO_542 (O_542,N_14945,N_14923);
or UO_543 (O_543,N_14532,N_14656);
xor UO_544 (O_544,N_14953,N_14856);
nor UO_545 (O_545,N_14743,N_14962);
xnor UO_546 (O_546,N_14561,N_14562);
nand UO_547 (O_547,N_14605,N_14871);
xor UO_548 (O_548,N_14514,N_14980);
nor UO_549 (O_549,N_14775,N_14658);
nor UO_550 (O_550,N_14878,N_14856);
nor UO_551 (O_551,N_14529,N_14916);
nor UO_552 (O_552,N_14960,N_14777);
nand UO_553 (O_553,N_14598,N_14947);
or UO_554 (O_554,N_14921,N_14656);
xnor UO_555 (O_555,N_14627,N_14878);
xnor UO_556 (O_556,N_14819,N_14663);
nor UO_557 (O_557,N_14729,N_14771);
nor UO_558 (O_558,N_14750,N_14607);
and UO_559 (O_559,N_14561,N_14567);
nand UO_560 (O_560,N_14989,N_14516);
xor UO_561 (O_561,N_14520,N_14553);
and UO_562 (O_562,N_14916,N_14701);
or UO_563 (O_563,N_14726,N_14953);
or UO_564 (O_564,N_14645,N_14644);
and UO_565 (O_565,N_14852,N_14796);
and UO_566 (O_566,N_14858,N_14689);
and UO_567 (O_567,N_14630,N_14576);
and UO_568 (O_568,N_14967,N_14596);
or UO_569 (O_569,N_14513,N_14681);
and UO_570 (O_570,N_14524,N_14817);
xnor UO_571 (O_571,N_14663,N_14552);
or UO_572 (O_572,N_14873,N_14627);
nand UO_573 (O_573,N_14877,N_14556);
xor UO_574 (O_574,N_14736,N_14725);
and UO_575 (O_575,N_14613,N_14538);
xor UO_576 (O_576,N_14581,N_14523);
or UO_577 (O_577,N_14553,N_14770);
xnor UO_578 (O_578,N_14615,N_14774);
xor UO_579 (O_579,N_14870,N_14580);
and UO_580 (O_580,N_14583,N_14822);
and UO_581 (O_581,N_14967,N_14702);
or UO_582 (O_582,N_14927,N_14836);
and UO_583 (O_583,N_14741,N_14976);
and UO_584 (O_584,N_14564,N_14743);
and UO_585 (O_585,N_14759,N_14780);
and UO_586 (O_586,N_14886,N_14682);
or UO_587 (O_587,N_14598,N_14627);
xor UO_588 (O_588,N_14981,N_14756);
and UO_589 (O_589,N_14829,N_14940);
xnor UO_590 (O_590,N_14589,N_14743);
nand UO_591 (O_591,N_14869,N_14739);
and UO_592 (O_592,N_14864,N_14555);
nor UO_593 (O_593,N_14777,N_14862);
nand UO_594 (O_594,N_14785,N_14502);
xnor UO_595 (O_595,N_14651,N_14733);
or UO_596 (O_596,N_14978,N_14503);
xor UO_597 (O_597,N_14910,N_14522);
and UO_598 (O_598,N_14835,N_14573);
and UO_599 (O_599,N_14584,N_14880);
xor UO_600 (O_600,N_14797,N_14736);
nor UO_601 (O_601,N_14647,N_14622);
nor UO_602 (O_602,N_14801,N_14764);
xnor UO_603 (O_603,N_14803,N_14977);
xnor UO_604 (O_604,N_14582,N_14847);
nand UO_605 (O_605,N_14769,N_14905);
xor UO_606 (O_606,N_14931,N_14718);
or UO_607 (O_607,N_14883,N_14546);
or UO_608 (O_608,N_14514,N_14685);
and UO_609 (O_609,N_14740,N_14679);
nand UO_610 (O_610,N_14611,N_14545);
xnor UO_611 (O_611,N_14991,N_14648);
nand UO_612 (O_612,N_14549,N_14670);
nand UO_613 (O_613,N_14661,N_14505);
xnor UO_614 (O_614,N_14997,N_14834);
xor UO_615 (O_615,N_14880,N_14602);
xor UO_616 (O_616,N_14718,N_14517);
or UO_617 (O_617,N_14632,N_14801);
xnor UO_618 (O_618,N_14704,N_14505);
and UO_619 (O_619,N_14526,N_14642);
nor UO_620 (O_620,N_14822,N_14502);
and UO_621 (O_621,N_14577,N_14702);
xor UO_622 (O_622,N_14775,N_14935);
or UO_623 (O_623,N_14652,N_14647);
nor UO_624 (O_624,N_14791,N_14987);
nor UO_625 (O_625,N_14631,N_14661);
or UO_626 (O_626,N_14786,N_14914);
nor UO_627 (O_627,N_14615,N_14796);
nor UO_628 (O_628,N_14730,N_14898);
nand UO_629 (O_629,N_14695,N_14713);
xnor UO_630 (O_630,N_14560,N_14813);
nand UO_631 (O_631,N_14586,N_14509);
xnor UO_632 (O_632,N_14979,N_14604);
or UO_633 (O_633,N_14589,N_14895);
nor UO_634 (O_634,N_14967,N_14878);
nor UO_635 (O_635,N_14951,N_14638);
or UO_636 (O_636,N_14720,N_14691);
xnor UO_637 (O_637,N_14935,N_14582);
or UO_638 (O_638,N_14529,N_14719);
or UO_639 (O_639,N_14576,N_14932);
xnor UO_640 (O_640,N_14931,N_14945);
nand UO_641 (O_641,N_14885,N_14875);
and UO_642 (O_642,N_14663,N_14713);
and UO_643 (O_643,N_14658,N_14993);
nor UO_644 (O_644,N_14630,N_14961);
xor UO_645 (O_645,N_14501,N_14830);
xnor UO_646 (O_646,N_14515,N_14661);
and UO_647 (O_647,N_14943,N_14885);
nand UO_648 (O_648,N_14827,N_14546);
or UO_649 (O_649,N_14732,N_14794);
and UO_650 (O_650,N_14852,N_14744);
xor UO_651 (O_651,N_14614,N_14776);
xor UO_652 (O_652,N_14802,N_14774);
or UO_653 (O_653,N_14963,N_14867);
nand UO_654 (O_654,N_14656,N_14853);
nand UO_655 (O_655,N_14640,N_14596);
nand UO_656 (O_656,N_14743,N_14781);
and UO_657 (O_657,N_14765,N_14612);
nor UO_658 (O_658,N_14916,N_14572);
or UO_659 (O_659,N_14564,N_14649);
or UO_660 (O_660,N_14930,N_14620);
and UO_661 (O_661,N_14596,N_14804);
xor UO_662 (O_662,N_14502,N_14604);
nor UO_663 (O_663,N_14797,N_14543);
nand UO_664 (O_664,N_14920,N_14694);
or UO_665 (O_665,N_14886,N_14630);
or UO_666 (O_666,N_14958,N_14998);
or UO_667 (O_667,N_14660,N_14816);
and UO_668 (O_668,N_14877,N_14900);
nand UO_669 (O_669,N_14597,N_14773);
nand UO_670 (O_670,N_14518,N_14750);
and UO_671 (O_671,N_14732,N_14824);
and UO_672 (O_672,N_14988,N_14776);
and UO_673 (O_673,N_14664,N_14672);
and UO_674 (O_674,N_14918,N_14746);
or UO_675 (O_675,N_14539,N_14897);
nand UO_676 (O_676,N_14622,N_14986);
and UO_677 (O_677,N_14942,N_14954);
and UO_678 (O_678,N_14908,N_14980);
and UO_679 (O_679,N_14959,N_14608);
or UO_680 (O_680,N_14840,N_14513);
nor UO_681 (O_681,N_14895,N_14887);
nor UO_682 (O_682,N_14930,N_14523);
nor UO_683 (O_683,N_14588,N_14696);
nor UO_684 (O_684,N_14727,N_14698);
nor UO_685 (O_685,N_14736,N_14834);
nand UO_686 (O_686,N_14607,N_14711);
and UO_687 (O_687,N_14708,N_14829);
nand UO_688 (O_688,N_14792,N_14930);
and UO_689 (O_689,N_14730,N_14927);
nand UO_690 (O_690,N_14831,N_14856);
xor UO_691 (O_691,N_14618,N_14716);
and UO_692 (O_692,N_14764,N_14921);
or UO_693 (O_693,N_14639,N_14546);
nand UO_694 (O_694,N_14917,N_14659);
nand UO_695 (O_695,N_14726,N_14713);
and UO_696 (O_696,N_14604,N_14959);
or UO_697 (O_697,N_14693,N_14689);
and UO_698 (O_698,N_14689,N_14788);
xnor UO_699 (O_699,N_14696,N_14914);
and UO_700 (O_700,N_14880,N_14603);
nand UO_701 (O_701,N_14919,N_14967);
nand UO_702 (O_702,N_14825,N_14589);
xnor UO_703 (O_703,N_14962,N_14892);
xor UO_704 (O_704,N_14707,N_14870);
nor UO_705 (O_705,N_14558,N_14812);
xor UO_706 (O_706,N_14663,N_14650);
nand UO_707 (O_707,N_14590,N_14828);
and UO_708 (O_708,N_14930,N_14961);
nor UO_709 (O_709,N_14853,N_14834);
nor UO_710 (O_710,N_14732,N_14572);
or UO_711 (O_711,N_14783,N_14931);
xor UO_712 (O_712,N_14888,N_14784);
nor UO_713 (O_713,N_14788,N_14769);
or UO_714 (O_714,N_14923,N_14542);
or UO_715 (O_715,N_14991,N_14954);
nor UO_716 (O_716,N_14515,N_14692);
xor UO_717 (O_717,N_14821,N_14774);
or UO_718 (O_718,N_14999,N_14626);
or UO_719 (O_719,N_14977,N_14941);
xnor UO_720 (O_720,N_14589,N_14719);
nor UO_721 (O_721,N_14793,N_14909);
and UO_722 (O_722,N_14588,N_14517);
and UO_723 (O_723,N_14689,N_14961);
or UO_724 (O_724,N_14838,N_14565);
and UO_725 (O_725,N_14875,N_14957);
xor UO_726 (O_726,N_14891,N_14610);
or UO_727 (O_727,N_14774,N_14760);
xor UO_728 (O_728,N_14564,N_14654);
nand UO_729 (O_729,N_14956,N_14765);
nand UO_730 (O_730,N_14882,N_14558);
xnor UO_731 (O_731,N_14581,N_14771);
or UO_732 (O_732,N_14819,N_14531);
nor UO_733 (O_733,N_14574,N_14789);
nor UO_734 (O_734,N_14943,N_14888);
nand UO_735 (O_735,N_14812,N_14714);
xor UO_736 (O_736,N_14579,N_14860);
or UO_737 (O_737,N_14766,N_14513);
and UO_738 (O_738,N_14860,N_14761);
nand UO_739 (O_739,N_14684,N_14757);
and UO_740 (O_740,N_14943,N_14993);
nor UO_741 (O_741,N_14914,N_14885);
xor UO_742 (O_742,N_14721,N_14763);
or UO_743 (O_743,N_14922,N_14955);
nor UO_744 (O_744,N_14768,N_14828);
or UO_745 (O_745,N_14940,N_14886);
or UO_746 (O_746,N_14957,N_14601);
nor UO_747 (O_747,N_14502,N_14589);
nand UO_748 (O_748,N_14867,N_14670);
xnor UO_749 (O_749,N_14565,N_14996);
and UO_750 (O_750,N_14554,N_14929);
or UO_751 (O_751,N_14718,N_14758);
xor UO_752 (O_752,N_14771,N_14559);
or UO_753 (O_753,N_14663,N_14701);
xor UO_754 (O_754,N_14922,N_14875);
and UO_755 (O_755,N_14864,N_14980);
nor UO_756 (O_756,N_14547,N_14689);
nand UO_757 (O_757,N_14786,N_14537);
nor UO_758 (O_758,N_14537,N_14905);
nand UO_759 (O_759,N_14874,N_14635);
and UO_760 (O_760,N_14525,N_14695);
xnor UO_761 (O_761,N_14652,N_14821);
nand UO_762 (O_762,N_14980,N_14799);
nor UO_763 (O_763,N_14778,N_14801);
and UO_764 (O_764,N_14856,N_14525);
xnor UO_765 (O_765,N_14838,N_14867);
xor UO_766 (O_766,N_14863,N_14672);
nor UO_767 (O_767,N_14683,N_14653);
xnor UO_768 (O_768,N_14531,N_14814);
nor UO_769 (O_769,N_14699,N_14534);
nor UO_770 (O_770,N_14939,N_14888);
and UO_771 (O_771,N_14510,N_14975);
and UO_772 (O_772,N_14799,N_14828);
nor UO_773 (O_773,N_14725,N_14993);
xnor UO_774 (O_774,N_14537,N_14942);
xor UO_775 (O_775,N_14846,N_14793);
xor UO_776 (O_776,N_14932,N_14551);
xor UO_777 (O_777,N_14752,N_14736);
nand UO_778 (O_778,N_14734,N_14575);
nor UO_779 (O_779,N_14522,N_14729);
nor UO_780 (O_780,N_14807,N_14759);
nand UO_781 (O_781,N_14587,N_14765);
or UO_782 (O_782,N_14781,N_14612);
or UO_783 (O_783,N_14653,N_14970);
or UO_784 (O_784,N_14727,N_14715);
nand UO_785 (O_785,N_14745,N_14707);
or UO_786 (O_786,N_14516,N_14802);
nor UO_787 (O_787,N_14827,N_14732);
or UO_788 (O_788,N_14917,N_14618);
nand UO_789 (O_789,N_14857,N_14595);
nand UO_790 (O_790,N_14958,N_14609);
nor UO_791 (O_791,N_14856,N_14672);
nor UO_792 (O_792,N_14769,N_14622);
or UO_793 (O_793,N_14532,N_14863);
xnor UO_794 (O_794,N_14978,N_14893);
nand UO_795 (O_795,N_14615,N_14767);
or UO_796 (O_796,N_14540,N_14750);
or UO_797 (O_797,N_14661,N_14826);
or UO_798 (O_798,N_14954,N_14865);
xor UO_799 (O_799,N_14986,N_14708);
xor UO_800 (O_800,N_14907,N_14983);
or UO_801 (O_801,N_14657,N_14681);
xor UO_802 (O_802,N_14870,N_14892);
nor UO_803 (O_803,N_14979,N_14616);
and UO_804 (O_804,N_14702,N_14930);
nand UO_805 (O_805,N_14542,N_14709);
and UO_806 (O_806,N_14967,N_14529);
nor UO_807 (O_807,N_14785,N_14630);
and UO_808 (O_808,N_14500,N_14922);
nor UO_809 (O_809,N_14605,N_14701);
and UO_810 (O_810,N_14912,N_14787);
xor UO_811 (O_811,N_14721,N_14717);
xor UO_812 (O_812,N_14938,N_14966);
nand UO_813 (O_813,N_14899,N_14876);
xnor UO_814 (O_814,N_14669,N_14685);
xnor UO_815 (O_815,N_14585,N_14694);
xnor UO_816 (O_816,N_14720,N_14779);
xnor UO_817 (O_817,N_14800,N_14500);
nand UO_818 (O_818,N_14774,N_14681);
xor UO_819 (O_819,N_14508,N_14512);
xor UO_820 (O_820,N_14798,N_14867);
or UO_821 (O_821,N_14871,N_14696);
xor UO_822 (O_822,N_14969,N_14585);
and UO_823 (O_823,N_14527,N_14981);
nand UO_824 (O_824,N_14523,N_14631);
nand UO_825 (O_825,N_14820,N_14593);
and UO_826 (O_826,N_14553,N_14521);
nand UO_827 (O_827,N_14905,N_14817);
xnor UO_828 (O_828,N_14807,N_14536);
and UO_829 (O_829,N_14922,N_14767);
xnor UO_830 (O_830,N_14633,N_14956);
xnor UO_831 (O_831,N_14988,N_14626);
and UO_832 (O_832,N_14803,N_14648);
nand UO_833 (O_833,N_14966,N_14767);
and UO_834 (O_834,N_14747,N_14608);
xnor UO_835 (O_835,N_14862,N_14914);
nor UO_836 (O_836,N_14872,N_14847);
xnor UO_837 (O_837,N_14680,N_14930);
xor UO_838 (O_838,N_14889,N_14649);
nor UO_839 (O_839,N_14962,N_14849);
nor UO_840 (O_840,N_14834,N_14760);
nand UO_841 (O_841,N_14506,N_14736);
nor UO_842 (O_842,N_14790,N_14525);
nor UO_843 (O_843,N_14739,N_14772);
and UO_844 (O_844,N_14631,N_14769);
xor UO_845 (O_845,N_14937,N_14751);
or UO_846 (O_846,N_14576,N_14904);
nand UO_847 (O_847,N_14643,N_14591);
or UO_848 (O_848,N_14854,N_14970);
xnor UO_849 (O_849,N_14973,N_14945);
nand UO_850 (O_850,N_14866,N_14565);
nand UO_851 (O_851,N_14790,N_14815);
xnor UO_852 (O_852,N_14818,N_14840);
and UO_853 (O_853,N_14650,N_14716);
and UO_854 (O_854,N_14696,N_14501);
or UO_855 (O_855,N_14891,N_14581);
nor UO_856 (O_856,N_14970,N_14768);
xnor UO_857 (O_857,N_14990,N_14671);
nor UO_858 (O_858,N_14815,N_14915);
or UO_859 (O_859,N_14717,N_14702);
and UO_860 (O_860,N_14723,N_14983);
nand UO_861 (O_861,N_14986,N_14628);
nand UO_862 (O_862,N_14946,N_14787);
and UO_863 (O_863,N_14675,N_14587);
and UO_864 (O_864,N_14595,N_14626);
nand UO_865 (O_865,N_14802,N_14505);
nand UO_866 (O_866,N_14806,N_14760);
xnor UO_867 (O_867,N_14545,N_14521);
nor UO_868 (O_868,N_14724,N_14568);
nor UO_869 (O_869,N_14821,N_14604);
xnor UO_870 (O_870,N_14563,N_14904);
xor UO_871 (O_871,N_14683,N_14899);
nand UO_872 (O_872,N_14611,N_14983);
and UO_873 (O_873,N_14564,N_14713);
or UO_874 (O_874,N_14986,N_14858);
nand UO_875 (O_875,N_14790,N_14876);
xnor UO_876 (O_876,N_14722,N_14696);
nor UO_877 (O_877,N_14860,N_14722);
nand UO_878 (O_878,N_14670,N_14961);
nor UO_879 (O_879,N_14974,N_14693);
nor UO_880 (O_880,N_14669,N_14990);
xor UO_881 (O_881,N_14685,N_14610);
xor UO_882 (O_882,N_14911,N_14824);
and UO_883 (O_883,N_14701,N_14529);
nor UO_884 (O_884,N_14708,N_14613);
or UO_885 (O_885,N_14945,N_14981);
nor UO_886 (O_886,N_14797,N_14533);
nand UO_887 (O_887,N_14667,N_14914);
xor UO_888 (O_888,N_14687,N_14827);
xnor UO_889 (O_889,N_14876,N_14991);
xnor UO_890 (O_890,N_14643,N_14743);
and UO_891 (O_891,N_14524,N_14878);
or UO_892 (O_892,N_14807,N_14955);
nand UO_893 (O_893,N_14547,N_14917);
or UO_894 (O_894,N_14939,N_14644);
or UO_895 (O_895,N_14879,N_14610);
xnor UO_896 (O_896,N_14757,N_14554);
xnor UO_897 (O_897,N_14838,N_14903);
nand UO_898 (O_898,N_14580,N_14520);
or UO_899 (O_899,N_14864,N_14711);
xnor UO_900 (O_900,N_14727,N_14571);
or UO_901 (O_901,N_14566,N_14851);
and UO_902 (O_902,N_14688,N_14501);
or UO_903 (O_903,N_14571,N_14633);
nand UO_904 (O_904,N_14921,N_14686);
nor UO_905 (O_905,N_14961,N_14586);
xor UO_906 (O_906,N_14740,N_14860);
nand UO_907 (O_907,N_14727,N_14714);
nand UO_908 (O_908,N_14966,N_14668);
nor UO_909 (O_909,N_14649,N_14981);
nand UO_910 (O_910,N_14697,N_14611);
xnor UO_911 (O_911,N_14903,N_14848);
nand UO_912 (O_912,N_14694,N_14653);
nand UO_913 (O_913,N_14648,N_14659);
nor UO_914 (O_914,N_14586,N_14550);
nand UO_915 (O_915,N_14959,N_14527);
xor UO_916 (O_916,N_14628,N_14603);
nand UO_917 (O_917,N_14798,N_14613);
nand UO_918 (O_918,N_14502,N_14911);
and UO_919 (O_919,N_14791,N_14841);
nor UO_920 (O_920,N_14767,N_14524);
xnor UO_921 (O_921,N_14895,N_14673);
nor UO_922 (O_922,N_14891,N_14904);
nor UO_923 (O_923,N_14716,N_14569);
nor UO_924 (O_924,N_14804,N_14508);
nor UO_925 (O_925,N_14964,N_14875);
nor UO_926 (O_926,N_14994,N_14887);
or UO_927 (O_927,N_14633,N_14504);
xor UO_928 (O_928,N_14649,N_14563);
nor UO_929 (O_929,N_14924,N_14784);
nand UO_930 (O_930,N_14536,N_14639);
nor UO_931 (O_931,N_14976,N_14930);
nor UO_932 (O_932,N_14531,N_14831);
and UO_933 (O_933,N_14590,N_14873);
and UO_934 (O_934,N_14889,N_14583);
nor UO_935 (O_935,N_14892,N_14660);
nand UO_936 (O_936,N_14728,N_14945);
or UO_937 (O_937,N_14667,N_14658);
or UO_938 (O_938,N_14937,N_14768);
or UO_939 (O_939,N_14891,N_14878);
and UO_940 (O_940,N_14975,N_14862);
and UO_941 (O_941,N_14883,N_14800);
and UO_942 (O_942,N_14527,N_14767);
nand UO_943 (O_943,N_14854,N_14651);
and UO_944 (O_944,N_14504,N_14900);
nand UO_945 (O_945,N_14532,N_14574);
xor UO_946 (O_946,N_14872,N_14708);
or UO_947 (O_947,N_14813,N_14648);
nand UO_948 (O_948,N_14843,N_14534);
nand UO_949 (O_949,N_14964,N_14826);
and UO_950 (O_950,N_14581,N_14506);
or UO_951 (O_951,N_14968,N_14806);
nand UO_952 (O_952,N_14779,N_14604);
or UO_953 (O_953,N_14962,N_14591);
nand UO_954 (O_954,N_14650,N_14787);
or UO_955 (O_955,N_14861,N_14876);
or UO_956 (O_956,N_14542,N_14848);
or UO_957 (O_957,N_14545,N_14992);
and UO_958 (O_958,N_14670,N_14541);
and UO_959 (O_959,N_14677,N_14633);
nand UO_960 (O_960,N_14980,N_14795);
or UO_961 (O_961,N_14563,N_14529);
or UO_962 (O_962,N_14660,N_14679);
nor UO_963 (O_963,N_14983,N_14904);
and UO_964 (O_964,N_14913,N_14659);
and UO_965 (O_965,N_14642,N_14650);
xnor UO_966 (O_966,N_14654,N_14516);
or UO_967 (O_967,N_14691,N_14506);
xor UO_968 (O_968,N_14743,N_14949);
nor UO_969 (O_969,N_14928,N_14578);
or UO_970 (O_970,N_14557,N_14892);
xnor UO_971 (O_971,N_14672,N_14732);
nand UO_972 (O_972,N_14920,N_14764);
or UO_973 (O_973,N_14849,N_14890);
nand UO_974 (O_974,N_14810,N_14673);
or UO_975 (O_975,N_14969,N_14824);
or UO_976 (O_976,N_14628,N_14980);
xnor UO_977 (O_977,N_14809,N_14945);
or UO_978 (O_978,N_14719,N_14713);
nand UO_979 (O_979,N_14539,N_14670);
or UO_980 (O_980,N_14710,N_14582);
nor UO_981 (O_981,N_14988,N_14679);
nand UO_982 (O_982,N_14790,N_14725);
nand UO_983 (O_983,N_14770,N_14870);
nand UO_984 (O_984,N_14670,N_14972);
or UO_985 (O_985,N_14589,N_14515);
xor UO_986 (O_986,N_14707,N_14589);
xnor UO_987 (O_987,N_14589,N_14891);
or UO_988 (O_988,N_14855,N_14927);
and UO_989 (O_989,N_14604,N_14671);
or UO_990 (O_990,N_14949,N_14983);
nand UO_991 (O_991,N_14810,N_14942);
nor UO_992 (O_992,N_14604,N_14512);
nand UO_993 (O_993,N_14630,N_14697);
nand UO_994 (O_994,N_14650,N_14683);
xor UO_995 (O_995,N_14598,N_14772);
xor UO_996 (O_996,N_14968,N_14613);
xor UO_997 (O_997,N_14527,N_14517);
and UO_998 (O_998,N_14608,N_14540);
or UO_999 (O_999,N_14980,N_14599);
xor UO_1000 (O_1000,N_14562,N_14875);
nor UO_1001 (O_1001,N_14500,N_14515);
and UO_1002 (O_1002,N_14558,N_14658);
nand UO_1003 (O_1003,N_14923,N_14954);
and UO_1004 (O_1004,N_14536,N_14867);
or UO_1005 (O_1005,N_14950,N_14960);
xnor UO_1006 (O_1006,N_14696,N_14613);
nand UO_1007 (O_1007,N_14871,N_14647);
xnor UO_1008 (O_1008,N_14879,N_14750);
nand UO_1009 (O_1009,N_14757,N_14878);
and UO_1010 (O_1010,N_14769,N_14707);
or UO_1011 (O_1011,N_14978,N_14697);
nor UO_1012 (O_1012,N_14655,N_14739);
and UO_1013 (O_1013,N_14636,N_14572);
xnor UO_1014 (O_1014,N_14554,N_14665);
nor UO_1015 (O_1015,N_14624,N_14770);
or UO_1016 (O_1016,N_14604,N_14925);
and UO_1017 (O_1017,N_14991,N_14957);
and UO_1018 (O_1018,N_14739,N_14683);
or UO_1019 (O_1019,N_14527,N_14998);
or UO_1020 (O_1020,N_14610,N_14682);
and UO_1021 (O_1021,N_14688,N_14549);
and UO_1022 (O_1022,N_14686,N_14607);
xnor UO_1023 (O_1023,N_14613,N_14704);
and UO_1024 (O_1024,N_14596,N_14629);
nand UO_1025 (O_1025,N_14584,N_14970);
nand UO_1026 (O_1026,N_14868,N_14761);
nand UO_1027 (O_1027,N_14709,N_14612);
xnor UO_1028 (O_1028,N_14563,N_14686);
xnor UO_1029 (O_1029,N_14718,N_14854);
and UO_1030 (O_1030,N_14777,N_14751);
and UO_1031 (O_1031,N_14998,N_14792);
nand UO_1032 (O_1032,N_14949,N_14549);
nand UO_1033 (O_1033,N_14533,N_14743);
and UO_1034 (O_1034,N_14995,N_14708);
nand UO_1035 (O_1035,N_14797,N_14902);
xor UO_1036 (O_1036,N_14866,N_14834);
nand UO_1037 (O_1037,N_14981,N_14808);
and UO_1038 (O_1038,N_14798,N_14503);
or UO_1039 (O_1039,N_14987,N_14906);
and UO_1040 (O_1040,N_14964,N_14946);
nor UO_1041 (O_1041,N_14790,N_14798);
nand UO_1042 (O_1042,N_14606,N_14718);
nand UO_1043 (O_1043,N_14879,N_14699);
nand UO_1044 (O_1044,N_14501,N_14737);
nor UO_1045 (O_1045,N_14982,N_14820);
and UO_1046 (O_1046,N_14658,N_14876);
or UO_1047 (O_1047,N_14644,N_14576);
or UO_1048 (O_1048,N_14869,N_14985);
xnor UO_1049 (O_1049,N_14950,N_14650);
nor UO_1050 (O_1050,N_14584,N_14517);
nand UO_1051 (O_1051,N_14518,N_14940);
or UO_1052 (O_1052,N_14688,N_14514);
nand UO_1053 (O_1053,N_14858,N_14580);
nand UO_1054 (O_1054,N_14982,N_14504);
nor UO_1055 (O_1055,N_14554,N_14740);
nand UO_1056 (O_1056,N_14830,N_14760);
nor UO_1057 (O_1057,N_14897,N_14972);
or UO_1058 (O_1058,N_14859,N_14779);
nand UO_1059 (O_1059,N_14981,N_14801);
xor UO_1060 (O_1060,N_14696,N_14776);
nor UO_1061 (O_1061,N_14655,N_14679);
nor UO_1062 (O_1062,N_14901,N_14873);
xor UO_1063 (O_1063,N_14977,N_14801);
xor UO_1064 (O_1064,N_14969,N_14765);
or UO_1065 (O_1065,N_14954,N_14799);
nor UO_1066 (O_1066,N_14720,N_14623);
nor UO_1067 (O_1067,N_14690,N_14504);
nor UO_1068 (O_1068,N_14955,N_14630);
and UO_1069 (O_1069,N_14513,N_14791);
xor UO_1070 (O_1070,N_14783,N_14799);
nand UO_1071 (O_1071,N_14887,N_14827);
nor UO_1072 (O_1072,N_14654,N_14508);
or UO_1073 (O_1073,N_14893,N_14634);
or UO_1074 (O_1074,N_14913,N_14936);
xor UO_1075 (O_1075,N_14875,N_14807);
and UO_1076 (O_1076,N_14749,N_14596);
and UO_1077 (O_1077,N_14544,N_14583);
and UO_1078 (O_1078,N_14534,N_14783);
nand UO_1079 (O_1079,N_14711,N_14990);
or UO_1080 (O_1080,N_14983,N_14911);
xor UO_1081 (O_1081,N_14675,N_14956);
nand UO_1082 (O_1082,N_14875,N_14519);
nand UO_1083 (O_1083,N_14859,N_14745);
or UO_1084 (O_1084,N_14789,N_14936);
nor UO_1085 (O_1085,N_14900,N_14896);
xor UO_1086 (O_1086,N_14555,N_14838);
xnor UO_1087 (O_1087,N_14765,N_14898);
nor UO_1088 (O_1088,N_14537,N_14857);
and UO_1089 (O_1089,N_14537,N_14966);
and UO_1090 (O_1090,N_14553,N_14949);
and UO_1091 (O_1091,N_14572,N_14633);
nor UO_1092 (O_1092,N_14587,N_14872);
nor UO_1093 (O_1093,N_14776,N_14784);
xor UO_1094 (O_1094,N_14650,N_14763);
or UO_1095 (O_1095,N_14767,N_14639);
nand UO_1096 (O_1096,N_14885,N_14665);
xor UO_1097 (O_1097,N_14773,N_14515);
nor UO_1098 (O_1098,N_14526,N_14550);
or UO_1099 (O_1099,N_14901,N_14745);
and UO_1100 (O_1100,N_14606,N_14598);
xnor UO_1101 (O_1101,N_14537,N_14876);
nand UO_1102 (O_1102,N_14675,N_14599);
or UO_1103 (O_1103,N_14516,N_14602);
nor UO_1104 (O_1104,N_14644,N_14779);
xnor UO_1105 (O_1105,N_14597,N_14510);
nand UO_1106 (O_1106,N_14826,N_14718);
or UO_1107 (O_1107,N_14989,N_14541);
and UO_1108 (O_1108,N_14706,N_14503);
or UO_1109 (O_1109,N_14872,N_14990);
and UO_1110 (O_1110,N_14571,N_14973);
or UO_1111 (O_1111,N_14918,N_14733);
nor UO_1112 (O_1112,N_14631,N_14685);
xnor UO_1113 (O_1113,N_14513,N_14657);
nor UO_1114 (O_1114,N_14932,N_14590);
and UO_1115 (O_1115,N_14854,N_14918);
and UO_1116 (O_1116,N_14923,N_14927);
or UO_1117 (O_1117,N_14844,N_14560);
or UO_1118 (O_1118,N_14917,N_14712);
or UO_1119 (O_1119,N_14740,N_14687);
and UO_1120 (O_1120,N_14776,N_14718);
nor UO_1121 (O_1121,N_14913,N_14916);
and UO_1122 (O_1122,N_14714,N_14700);
nor UO_1123 (O_1123,N_14948,N_14614);
or UO_1124 (O_1124,N_14667,N_14776);
or UO_1125 (O_1125,N_14844,N_14927);
nor UO_1126 (O_1126,N_14509,N_14613);
or UO_1127 (O_1127,N_14719,N_14720);
nand UO_1128 (O_1128,N_14619,N_14670);
xor UO_1129 (O_1129,N_14710,N_14607);
nor UO_1130 (O_1130,N_14951,N_14656);
nand UO_1131 (O_1131,N_14744,N_14900);
nor UO_1132 (O_1132,N_14622,N_14600);
and UO_1133 (O_1133,N_14528,N_14634);
xnor UO_1134 (O_1134,N_14629,N_14844);
nor UO_1135 (O_1135,N_14519,N_14695);
xor UO_1136 (O_1136,N_14563,N_14708);
nor UO_1137 (O_1137,N_14775,N_14977);
and UO_1138 (O_1138,N_14599,N_14992);
nor UO_1139 (O_1139,N_14634,N_14716);
and UO_1140 (O_1140,N_14654,N_14703);
or UO_1141 (O_1141,N_14670,N_14870);
nand UO_1142 (O_1142,N_14544,N_14621);
nor UO_1143 (O_1143,N_14896,N_14766);
nor UO_1144 (O_1144,N_14903,N_14921);
or UO_1145 (O_1145,N_14770,N_14862);
nand UO_1146 (O_1146,N_14576,N_14992);
or UO_1147 (O_1147,N_14521,N_14520);
nor UO_1148 (O_1148,N_14936,N_14763);
xnor UO_1149 (O_1149,N_14924,N_14507);
or UO_1150 (O_1150,N_14686,N_14943);
nand UO_1151 (O_1151,N_14708,N_14792);
xor UO_1152 (O_1152,N_14613,N_14965);
nor UO_1153 (O_1153,N_14724,N_14962);
nand UO_1154 (O_1154,N_14720,N_14564);
and UO_1155 (O_1155,N_14515,N_14677);
or UO_1156 (O_1156,N_14642,N_14990);
or UO_1157 (O_1157,N_14656,N_14810);
nand UO_1158 (O_1158,N_14849,N_14978);
nand UO_1159 (O_1159,N_14751,N_14986);
and UO_1160 (O_1160,N_14843,N_14542);
nand UO_1161 (O_1161,N_14790,N_14720);
xor UO_1162 (O_1162,N_14818,N_14829);
and UO_1163 (O_1163,N_14715,N_14883);
or UO_1164 (O_1164,N_14695,N_14615);
xor UO_1165 (O_1165,N_14706,N_14779);
nor UO_1166 (O_1166,N_14684,N_14651);
xor UO_1167 (O_1167,N_14746,N_14991);
nand UO_1168 (O_1168,N_14633,N_14810);
and UO_1169 (O_1169,N_14638,N_14645);
and UO_1170 (O_1170,N_14906,N_14512);
nand UO_1171 (O_1171,N_14672,N_14581);
or UO_1172 (O_1172,N_14847,N_14728);
nor UO_1173 (O_1173,N_14870,N_14943);
and UO_1174 (O_1174,N_14924,N_14900);
and UO_1175 (O_1175,N_14725,N_14564);
xor UO_1176 (O_1176,N_14594,N_14601);
or UO_1177 (O_1177,N_14737,N_14588);
or UO_1178 (O_1178,N_14586,N_14640);
nand UO_1179 (O_1179,N_14738,N_14647);
or UO_1180 (O_1180,N_14637,N_14646);
nand UO_1181 (O_1181,N_14621,N_14885);
nand UO_1182 (O_1182,N_14603,N_14582);
xnor UO_1183 (O_1183,N_14617,N_14980);
or UO_1184 (O_1184,N_14959,N_14531);
nor UO_1185 (O_1185,N_14998,N_14545);
nand UO_1186 (O_1186,N_14729,N_14577);
xor UO_1187 (O_1187,N_14528,N_14512);
nand UO_1188 (O_1188,N_14606,N_14740);
nor UO_1189 (O_1189,N_14565,N_14559);
nand UO_1190 (O_1190,N_14807,N_14503);
xor UO_1191 (O_1191,N_14868,N_14968);
and UO_1192 (O_1192,N_14895,N_14864);
xor UO_1193 (O_1193,N_14619,N_14620);
nor UO_1194 (O_1194,N_14877,N_14534);
xnor UO_1195 (O_1195,N_14948,N_14995);
and UO_1196 (O_1196,N_14958,N_14802);
nand UO_1197 (O_1197,N_14709,N_14650);
nor UO_1198 (O_1198,N_14559,N_14850);
xnor UO_1199 (O_1199,N_14909,N_14861);
and UO_1200 (O_1200,N_14683,N_14575);
or UO_1201 (O_1201,N_14552,N_14799);
xor UO_1202 (O_1202,N_14898,N_14943);
nor UO_1203 (O_1203,N_14842,N_14978);
or UO_1204 (O_1204,N_14735,N_14852);
nor UO_1205 (O_1205,N_14728,N_14931);
xor UO_1206 (O_1206,N_14814,N_14834);
or UO_1207 (O_1207,N_14979,N_14984);
or UO_1208 (O_1208,N_14977,N_14844);
and UO_1209 (O_1209,N_14536,N_14834);
or UO_1210 (O_1210,N_14901,N_14749);
nand UO_1211 (O_1211,N_14729,N_14594);
nand UO_1212 (O_1212,N_14566,N_14798);
or UO_1213 (O_1213,N_14881,N_14559);
nor UO_1214 (O_1214,N_14856,N_14850);
nor UO_1215 (O_1215,N_14791,N_14876);
or UO_1216 (O_1216,N_14512,N_14660);
or UO_1217 (O_1217,N_14936,N_14732);
nor UO_1218 (O_1218,N_14535,N_14577);
and UO_1219 (O_1219,N_14750,N_14865);
nand UO_1220 (O_1220,N_14686,N_14666);
or UO_1221 (O_1221,N_14598,N_14791);
and UO_1222 (O_1222,N_14684,N_14833);
and UO_1223 (O_1223,N_14560,N_14847);
or UO_1224 (O_1224,N_14946,N_14765);
nor UO_1225 (O_1225,N_14773,N_14849);
and UO_1226 (O_1226,N_14510,N_14678);
nor UO_1227 (O_1227,N_14588,N_14549);
or UO_1228 (O_1228,N_14847,N_14708);
and UO_1229 (O_1229,N_14731,N_14674);
or UO_1230 (O_1230,N_14906,N_14756);
or UO_1231 (O_1231,N_14949,N_14526);
nor UO_1232 (O_1232,N_14821,N_14553);
or UO_1233 (O_1233,N_14711,N_14681);
or UO_1234 (O_1234,N_14736,N_14757);
and UO_1235 (O_1235,N_14758,N_14705);
or UO_1236 (O_1236,N_14742,N_14514);
nand UO_1237 (O_1237,N_14660,N_14575);
xnor UO_1238 (O_1238,N_14560,N_14919);
nand UO_1239 (O_1239,N_14834,N_14972);
or UO_1240 (O_1240,N_14954,N_14527);
and UO_1241 (O_1241,N_14939,N_14980);
nand UO_1242 (O_1242,N_14655,N_14729);
and UO_1243 (O_1243,N_14805,N_14978);
xor UO_1244 (O_1244,N_14895,N_14914);
nor UO_1245 (O_1245,N_14934,N_14969);
nand UO_1246 (O_1246,N_14727,N_14926);
xnor UO_1247 (O_1247,N_14959,N_14866);
and UO_1248 (O_1248,N_14665,N_14917);
xnor UO_1249 (O_1249,N_14619,N_14915);
xnor UO_1250 (O_1250,N_14799,N_14827);
or UO_1251 (O_1251,N_14601,N_14543);
xnor UO_1252 (O_1252,N_14863,N_14908);
xnor UO_1253 (O_1253,N_14827,N_14685);
and UO_1254 (O_1254,N_14984,N_14547);
nor UO_1255 (O_1255,N_14637,N_14988);
and UO_1256 (O_1256,N_14897,N_14808);
or UO_1257 (O_1257,N_14668,N_14601);
nand UO_1258 (O_1258,N_14995,N_14873);
and UO_1259 (O_1259,N_14885,N_14604);
or UO_1260 (O_1260,N_14634,N_14534);
nor UO_1261 (O_1261,N_14631,N_14509);
or UO_1262 (O_1262,N_14728,N_14915);
xor UO_1263 (O_1263,N_14562,N_14506);
nand UO_1264 (O_1264,N_14530,N_14955);
xor UO_1265 (O_1265,N_14842,N_14867);
nand UO_1266 (O_1266,N_14831,N_14563);
and UO_1267 (O_1267,N_14848,N_14691);
nand UO_1268 (O_1268,N_14540,N_14741);
xor UO_1269 (O_1269,N_14961,N_14504);
or UO_1270 (O_1270,N_14904,N_14587);
xnor UO_1271 (O_1271,N_14748,N_14667);
or UO_1272 (O_1272,N_14865,N_14982);
nor UO_1273 (O_1273,N_14547,N_14765);
nand UO_1274 (O_1274,N_14936,N_14815);
nand UO_1275 (O_1275,N_14932,N_14893);
and UO_1276 (O_1276,N_14761,N_14732);
or UO_1277 (O_1277,N_14984,N_14834);
and UO_1278 (O_1278,N_14687,N_14533);
xnor UO_1279 (O_1279,N_14942,N_14842);
or UO_1280 (O_1280,N_14532,N_14983);
xor UO_1281 (O_1281,N_14967,N_14901);
or UO_1282 (O_1282,N_14538,N_14949);
and UO_1283 (O_1283,N_14750,N_14901);
xor UO_1284 (O_1284,N_14724,N_14774);
nand UO_1285 (O_1285,N_14563,N_14823);
xor UO_1286 (O_1286,N_14843,N_14549);
or UO_1287 (O_1287,N_14634,N_14984);
or UO_1288 (O_1288,N_14933,N_14806);
and UO_1289 (O_1289,N_14638,N_14926);
nor UO_1290 (O_1290,N_14818,N_14574);
nand UO_1291 (O_1291,N_14627,N_14899);
or UO_1292 (O_1292,N_14633,N_14558);
xnor UO_1293 (O_1293,N_14736,N_14582);
nand UO_1294 (O_1294,N_14811,N_14588);
nand UO_1295 (O_1295,N_14636,N_14534);
and UO_1296 (O_1296,N_14752,N_14926);
xnor UO_1297 (O_1297,N_14587,N_14916);
and UO_1298 (O_1298,N_14766,N_14826);
xor UO_1299 (O_1299,N_14535,N_14737);
or UO_1300 (O_1300,N_14840,N_14699);
or UO_1301 (O_1301,N_14681,N_14699);
or UO_1302 (O_1302,N_14697,N_14663);
and UO_1303 (O_1303,N_14664,N_14752);
or UO_1304 (O_1304,N_14741,N_14784);
xor UO_1305 (O_1305,N_14585,N_14768);
and UO_1306 (O_1306,N_14837,N_14504);
xor UO_1307 (O_1307,N_14504,N_14865);
or UO_1308 (O_1308,N_14701,N_14892);
nand UO_1309 (O_1309,N_14565,N_14768);
xnor UO_1310 (O_1310,N_14992,N_14832);
and UO_1311 (O_1311,N_14553,N_14699);
or UO_1312 (O_1312,N_14942,N_14600);
or UO_1313 (O_1313,N_14556,N_14918);
and UO_1314 (O_1314,N_14986,N_14897);
and UO_1315 (O_1315,N_14770,N_14930);
and UO_1316 (O_1316,N_14902,N_14942);
nand UO_1317 (O_1317,N_14622,N_14699);
and UO_1318 (O_1318,N_14845,N_14924);
and UO_1319 (O_1319,N_14646,N_14565);
nor UO_1320 (O_1320,N_14726,N_14691);
nor UO_1321 (O_1321,N_14641,N_14527);
or UO_1322 (O_1322,N_14871,N_14756);
and UO_1323 (O_1323,N_14712,N_14768);
nand UO_1324 (O_1324,N_14866,N_14572);
or UO_1325 (O_1325,N_14722,N_14611);
or UO_1326 (O_1326,N_14609,N_14602);
nand UO_1327 (O_1327,N_14971,N_14739);
or UO_1328 (O_1328,N_14884,N_14659);
or UO_1329 (O_1329,N_14669,N_14615);
or UO_1330 (O_1330,N_14663,N_14864);
nand UO_1331 (O_1331,N_14624,N_14792);
xor UO_1332 (O_1332,N_14847,N_14850);
nand UO_1333 (O_1333,N_14615,N_14756);
nor UO_1334 (O_1334,N_14681,N_14784);
xor UO_1335 (O_1335,N_14507,N_14797);
nand UO_1336 (O_1336,N_14956,N_14847);
and UO_1337 (O_1337,N_14674,N_14768);
or UO_1338 (O_1338,N_14683,N_14519);
and UO_1339 (O_1339,N_14800,N_14867);
nor UO_1340 (O_1340,N_14862,N_14726);
and UO_1341 (O_1341,N_14923,N_14689);
or UO_1342 (O_1342,N_14780,N_14518);
nor UO_1343 (O_1343,N_14888,N_14909);
or UO_1344 (O_1344,N_14613,N_14521);
nand UO_1345 (O_1345,N_14728,N_14616);
and UO_1346 (O_1346,N_14543,N_14773);
and UO_1347 (O_1347,N_14503,N_14715);
nor UO_1348 (O_1348,N_14650,N_14911);
or UO_1349 (O_1349,N_14548,N_14999);
xnor UO_1350 (O_1350,N_14993,N_14876);
nand UO_1351 (O_1351,N_14599,N_14612);
or UO_1352 (O_1352,N_14620,N_14747);
nor UO_1353 (O_1353,N_14948,N_14507);
xnor UO_1354 (O_1354,N_14524,N_14972);
and UO_1355 (O_1355,N_14569,N_14552);
xnor UO_1356 (O_1356,N_14589,N_14517);
xor UO_1357 (O_1357,N_14967,N_14833);
and UO_1358 (O_1358,N_14693,N_14928);
nand UO_1359 (O_1359,N_14850,N_14834);
and UO_1360 (O_1360,N_14724,N_14702);
or UO_1361 (O_1361,N_14949,N_14630);
or UO_1362 (O_1362,N_14924,N_14553);
and UO_1363 (O_1363,N_14593,N_14738);
xnor UO_1364 (O_1364,N_14858,N_14825);
xor UO_1365 (O_1365,N_14506,N_14720);
and UO_1366 (O_1366,N_14688,N_14614);
or UO_1367 (O_1367,N_14818,N_14680);
xnor UO_1368 (O_1368,N_14574,N_14840);
or UO_1369 (O_1369,N_14573,N_14871);
xnor UO_1370 (O_1370,N_14869,N_14689);
nor UO_1371 (O_1371,N_14529,N_14614);
nor UO_1372 (O_1372,N_14835,N_14644);
nand UO_1373 (O_1373,N_14777,N_14969);
or UO_1374 (O_1374,N_14507,N_14947);
or UO_1375 (O_1375,N_14672,N_14877);
xor UO_1376 (O_1376,N_14820,N_14512);
xnor UO_1377 (O_1377,N_14761,N_14728);
xor UO_1378 (O_1378,N_14566,N_14791);
xor UO_1379 (O_1379,N_14892,N_14949);
nand UO_1380 (O_1380,N_14612,N_14740);
and UO_1381 (O_1381,N_14865,N_14866);
nand UO_1382 (O_1382,N_14705,N_14816);
or UO_1383 (O_1383,N_14964,N_14955);
nand UO_1384 (O_1384,N_14988,N_14896);
or UO_1385 (O_1385,N_14728,N_14638);
xnor UO_1386 (O_1386,N_14671,N_14980);
or UO_1387 (O_1387,N_14908,N_14654);
or UO_1388 (O_1388,N_14755,N_14698);
xor UO_1389 (O_1389,N_14662,N_14830);
nor UO_1390 (O_1390,N_14702,N_14668);
xnor UO_1391 (O_1391,N_14929,N_14872);
and UO_1392 (O_1392,N_14646,N_14767);
nand UO_1393 (O_1393,N_14705,N_14759);
and UO_1394 (O_1394,N_14861,N_14641);
nand UO_1395 (O_1395,N_14987,N_14645);
nand UO_1396 (O_1396,N_14568,N_14584);
nor UO_1397 (O_1397,N_14963,N_14733);
or UO_1398 (O_1398,N_14572,N_14514);
or UO_1399 (O_1399,N_14983,N_14690);
and UO_1400 (O_1400,N_14995,N_14973);
nand UO_1401 (O_1401,N_14870,N_14828);
and UO_1402 (O_1402,N_14987,N_14718);
nand UO_1403 (O_1403,N_14819,N_14572);
xnor UO_1404 (O_1404,N_14848,N_14842);
nand UO_1405 (O_1405,N_14829,N_14844);
nand UO_1406 (O_1406,N_14728,N_14868);
or UO_1407 (O_1407,N_14591,N_14980);
nand UO_1408 (O_1408,N_14640,N_14703);
nor UO_1409 (O_1409,N_14544,N_14760);
xor UO_1410 (O_1410,N_14750,N_14547);
nand UO_1411 (O_1411,N_14842,N_14713);
or UO_1412 (O_1412,N_14750,N_14609);
nor UO_1413 (O_1413,N_14965,N_14592);
xnor UO_1414 (O_1414,N_14878,N_14779);
nand UO_1415 (O_1415,N_14976,N_14782);
nand UO_1416 (O_1416,N_14846,N_14585);
and UO_1417 (O_1417,N_14625,N_14791);
or UO_1418 (O_1418,N_14922,N_14645);
nor UO_1419 (O_1419,N_14701,N_14868);
xnor UO_1420 (O_1420,N_14926,N_14736);
xor UO_1421 (O_1421,N_14694,N_14819);
and UO_1422 (O_1422,N_14782,N_14871);
or UO_1423 (O_1423,N_14821,N_14630);
xor UO_1424 (O_1424,N_14828,N_14651);
and UO_1425 (O_1425,N_14763,N_14940);
xor UO_1426 (O_1426,N_14999,N_14565);
xor UO_1427 (O_1427,N_14789,N_14745);
or UO_1428 (O_1428,N_14862,N_14549);
xnor UO_1429 (O_1429,N_14710,N_14708);
xor UO_1430 (O_1430,N_14951,N_14681);
nand UO_1431 (O_1431,N_14898,N_14571);
xor UO_1432 (O_1432,N_14741,N_14946);
xnor UO_1433 (O_1433,N_14922,N_14503);
nor UO_1434 (O_1434,N_14908,N_14864);
xor UO_1435 (O_1435,N_14657,N_14618);
nor UO_1436 (O_1436,N_14533,N_14871);
xor UO_1437 (O_1437,N_14659,N_14835);
and UO_1438 (O_1438,N_14673,N_14771);
xnor UO_1439 (O_1439,N_14509,N_14878);
and UO_1440 (O_1440,N_14975,N_14563);
nand UO_1441 (O_1441,N_14576,N_14998);
or UO_1442 (O_1442,N_14928,N_14500);
or UO_1443 (O_1443,N_14940,N_14710);
nor UO_1444 (O_1444,N_14752,N_14805);
and UO_1445 (O_1445,N_14635,N_14717);
nand UO_1446 (O_1446,N_14736,N_14508);
nor UO_1447 (O_1447,N_14510,N_14747);
and UO_1448 (O_1448,N_14923,N_14839);
xor UO_1449 (O_1449,N_14813,N_14631);
nor UO_1450 (O_1450,N_14919,N_14968);
and UO_1451 (O_1451,N_14912,N_14948);
and UO_1452 (O_1452,N_14862,N_14852);
nand UO_1453 (O_1453,N_14593,N_14615);
nor UO_1454 (O_1454,N_14541,N_14837);
xnor UO_1455 (O_1455,N_14896,N_14686);
xnor UO_1456 (O_1456,N_14667,N_14574);
nor UO_1457 (O_1457,N_14785,N_14568);
xnor UO_1458 (O_1458,N_14577,N_14871);
xor UO_1459 (O_1459,N_14661,N_14819);
nand UO_1460 (O_1460,N_14845,N_14572);
and UO_1461 (O_1461,N_14902,N_14742);
nand UO_1462 (O_1462,N_14844,N_14934);
and UO_1463 (O_1463,N_14587,N_14626);
nor UO_1464 (O_1464,N_14979,N_14680);
and UO_1465 (O_1465,N_14701,N_14762);
nor UO_1466 (O_1466,N_14677,N_14928);
nand UO_1467 (O_1467,N_14618,N_14770);
nor UO_1468 (O_1468,N_14695,N_14945);
nor UO_1469 (O_1469,N_14521,N_14818);
and UO_1470 (O_1470,N_14592,N_14581);
or UO_1471 (O_1471,N_14594,N_14546);
nor UO_1472 (O_1472,N_14574,N_14762);
or UO_1473 (O_1473,N_14787,N_14505);
and UO_1474 (O_1474,N_14871,N_14785);
or UO_1475 (O_1475,N_14699,N_14961);
or UO_1476 (O_1476,N_14786,N_14902);
nand UO_1477 (O_1477,N_14812,N_14813);
nor UO_1478 (O_1478,N_14895,N_14982);
nor UO_1479 (O_1479,N_14865,N_14649);
nand UO_1480 (O_1480,N_14558,N_14791);
or UO_1481 (O_1481,N_14581,N_14767);
and UO_1482 (O_1482,N_14530,N_14512);
nand UO_1483 (O_1483,N_14925,N_14657);
xor UO_1484 (O_1484,N_14694,N_14629);
nand UO_1485 (O_1485,N_14633,N_14854);
and UO_1486 (O_1486,N_14820,N_14837);
and UO_1487 (O_1487,N_14749,N_14774);
or UO_1488 (O_1488,N_14539,N_14645);
xnor UO_1489 (O_1489,N_14569,N_14868);
and UO_1490 (O_1490,N_14685,N_14503);
nand UO_1491 (O_1491,N_14892,N_14573);
and UO_1492 (O_1492,N_14652,N_14960);
nor UO_1493 (O_1493,N_14939,N_14684);
nand UO_1494 (O_1494,N_14626,N_14666);
nand UO_1495 (O_1495,N_14829,N_14992);
nand UO_1496 (O_1496,N_14506,N_14784);
and UO_1497 (O_1497,N_14927,N_14799);
xnor UO_1498 (O_1498,N_14542,N_14907);
and UO_1499 (O_1499,N_14519,N_14879);
nand UO_1500 (O_1500,N_14828,N_14893);
nand UO_1501 (O_1501,N_14790,N_14512);
and UO_1502 (O_1502,N_14879,N_14970);
nor UO_1503 (O_1503,N_14893,N_14524);
nand UO_1504 (O_1504,N_14917,N_14962);
nor UO_1505 (O_1505,N_14930,N_14622);
nand UO_1506 (O_1506,N_14510,N_14782);
or UO_1507 (O_1507,N_14784,N_14765);
and UO_1508 (O_1508,N_14561,N_14806);
and UO_1509 (O_1509,N_14769,N_14603);
or UO_1510 (O_1510,N_14905,N_14967);
or UO_1511 (O_1511,N_14756,N_14597);
nand UO_1512 (O_1512,N_14863,N_14536);
and UO_1513 (O_1513,N_14752,N_14823);
and UO_1514 (O_1514,N_14949,N_14575);
and UO_1515 (O_1515,N_14889,N_14847);
xnor UO_1516 (O_1516,N_14664,N_14991);
xnor UO_1517 (O_1517,N_14983,N_14702);
or UO_1518 (O_1518,N_14680,N_14816);
and UO_1519 (O_1519,N_14940,N_14621);
xor UO_1520 (O_1520,N_14708,N_14878);
nor UO_1521 (O_1521,N_14591,N_14961);
and UO_1522 (O_1522,N_14935,N_14977);
xor UO_1523 (O_1523,N_14633,N_14998);
or UO_1524 (O_1524,N_14960,N_14669);
xnor UO_1525 (O_1525,N_14628,N_14640);
nand UO_1526 (O_1526,N_14520,N_14761);
xor UO_1527 (O_1527,N_14895,N_14669);
xor UO_1528 (O_1528,N_14526,N_14509);
xor UO_1529 (O_1529,N_14799,N_14944);
xnor UO_1530 (O_1530,N_14800,N_14557);
or UO_1531 (O_1531,N_14584,N_14610);
and UO_1532 (O_1532,N_14506,N_14647);
nand UO_1533 (O_1533,N_14600,N_14564);
xnor UO_1534 (O_1534,N_14567,N_14652);
and UO_1535 (O_1535,N_14875,N_14560);
and UO_1536 (O_1536,N_14553,N_14512);
nor UO_1537 (O_1537,N_14789,N_14504);
or UO_1538 (O_1538,N_14651,N_14642);
nor UO_1539 (O_1539,N_14868,N_14790);
and UO_1540 (O_1540,N_14637,N_14589);
nand UO_1541 (O_1541,N_14803,N_14670);
nor UO_1542 (O_1542,N_14932,N_14853);
or UO_1543 (O_1543,N_14671,N_14657);
nor UO_1544 (O_1544,N_14697,N_14875);
nor UO_1545 (O_1545,N_14766,N_14558);
nor UO_1546 (O_1546,N_14507,N_14974);
nor UO_1547 (O_1547,N_14671,N_14539);
xor UO_1548 (O_1548,N_14910,N_14564);
xnor UO_1549 (O_1549,N_14745,N_14981);
nor UO_1550 (O_1550,N_14520,N_14881);
xnor UO_1551 (O_1551,N_14702,N_14645);
xnor UO_1552 (O_1552,N_14569,N_14881);
nor UO_1553 (O_1553,N_14886,N_14657);
nor UO_1554 (O_1554,N_14753,N_14520);
xor UO_1555 (O_1555,N_14669,N_14753);
nand UO_1556 (O_1556,N_14607,N_14925);
nand UO_1557 (O_1557,N_14800,N_14558);
or UO_1558 (O_1558,N_14520,N_14856);
and UO_1559 (O_1559,N_14794,N_14682);
nand UO_1560 (O_1560,N_14657,N_14869);
nand UO_1561 (O_1561,N_14528,N_14951);
or UO_1562 (O_1562,N_14683,N_14535);
or UO_1563 (O_1563,N_14746,N_14816);
or UO_1564 (O_1564,N_14824,N_14535);
nand UO_1565 (O_1565,N_14774,N_14891);
or UO_1566 (O_1566,N_14597,N_14936);
nor UO_1567 (O_1567,N_14902,N_14767);
nand UO_1568 (O_1568,N_14785,N_14773);
and UO_1569 (O_1569,N_14723,N_14805);
and UO_1570 (O_1570,N_14862,N_14515);
nand UO_1571 (O_1571,N_14649,N_14734);
nand UO_1572 (O_1572,N_14697,N_14882);
xor UO_1573 (O_1573,N_14548,N_14783);
or UO_1574 (O_1574,N_14684,N_14589);
nand UO_1575 (O_1575,N_14599,N_14995);
nor UO_1576 (O_1576,N_14982,N_14971);
or UO_1577 (O_1577,N_14978,N_14962);
or UO_1578 (O_1578,N_14514,N_14559);
and UO_1579 (O_1579,N_14694,N_14767);
nor UO_1580 (O_1580,N_14806,N_14676);
and UO_1581 (O_1581,N_14551,N_14756);
and UO_1582 (O_1582,N_14672,N_14889);
nor UO_1583 (O_1583,N_14521,N_14549);
or UO_1584 (O_1584,N_14691,N_14884);
xor UO_1585 (O_1585,N_14739,N_14622);
nand UO_1586 (O_1586,N_14645,N_14934);
xnor UO_1587 (O_1587,N_14965,N_14538);
nor UO_1588 (O_1588,N_14551,N_14872);
or UO_1589 (O_1589,N_14967,N_14994);
or UO_1590 (O_1590,N_14907,N_14961);
xnor UO_1591 (O_1591,N_14743,N_14879);
nor UO_1592 (O_1592,N_14625,N_14843);
or UO_1593 (O_1593,N_14911,N_14802);
nand UO_1594 (O_1594,N_14759,N_14561);
xnor UO_1595 (O_1595,N_14776,N_14932);
and UO_1596 (O_1596,N_14875,N_14661);
and UO_1597 (O_1597,N_14536,N_14770);
nor UO_1598 (O_1598,N_14923,N_14581);
nand UO_1599 (O_1599,N_14787,N_14649);
xor UO_1600 (O_1600,N_14940,N_14944);
nand UO_1601 (O_1601,N_14619,N_14764);
nor UO_1602 (O_1602,N_14730,N_14861);
and UO_1603 (O_1603,N_14947,N_14779);
or UO_1604 (O_1604,N_14640,N_14668);
and UO_1605 (O_1605,N_14864,N_14603);
and UO_1606 (O_1606,N_14995,N_14664);
xor UO_1607 (O_1607,N_14924,N_14724);
or UO_1608 (O_1608,N_14883,N_14954);
or UO_1609 (O_1609,N_14556,N_14746);
or UO_1610 (O_1610,N_14917,N_14543);
or UO_1611 (O_1611,N_14734,N_14938);
or UO_1612 (O_1612,N_14547,N_14621);
or UO_1613 (O_1613,N_14973,N_14765);
nand UO_1614 (O_1614,N_14668,N_14545);
or UO_1615 (O_1615,N_14632,N_14782);
and UO_1616 (O_1616,N_14890,N_14878);
nor UO_1617 (O_1617,N_14942,N_14777);
nor UO_1618 (O_1618,N_14970,N_14874);
nand UO_1619 (O_1619,N_14773,N_14738);
or UO_1620 (O_1620,N_14984,N_14966);
nand UO_1621 (O_1621,N_14877,N_14928);
or UO_1622 (O_1622,N_14585,N_14828);
or UO_1623 (O_1623,N_14690,N_14646);
or UO_1624 (O_1624,N_14892,N_14798);
or UO_1625 (O_1625,N_14932,N_14935);
and UO_1626 (O_1626,N_14849,N_14660);
xnor UO_1627 (O_1627,N_14628,N_14767);
and UO_1628 (O_1628,N_14809,N_14826);
or UO_1629 (O_1629,N_14756,N_14500);
and UO_1630 (O_1630,N_14717,N_14999);
nand UO_1631 (O_1631,N_14608,N_14709);
or UO_1632 (O_1632,N_14581,N_14525);
and UO_1633 (O_1633,N_14997,N_14893);
nand UO_1634 (O_1634,N_14709,N_14909);
nor UO_1635 (O_1635,N_14920,N_14778);
xnor UO_1636 (O_1636,N_14621,N_14730);
and UO_1637 (O_1637,N_14579,N_14644);
nand UO_1638 (O_1638,N_14666,N_14639);
or UO_1639 (O_1639,N_14805,N_14989);
nand UO_1640 (O_1640,N_14599,N_14849);
nand UO_1641 (O_1641,N_14537,N_14926);
xnor UO_1642 (O_1642,N_14903,N_14648);
or UO_1643 (O_1643,N_14979,N_14830);
nand UO_1644 (O_1644,N_14701,N_14856);
or UO_1645 (O_1645,N_14880,N_14585);
nor UO_1646 (O_1646,N_14824,N_14724);
xor UO_1647 (O_1647,N_14573,N_14503);
xor UO_1648 (O_1648,N_14573,N_14723);
xor UO_1649 (O_1649,N_14827,N_14667);
and UO_1650 (O_1650,N_14923,N_14678);
nor UO_1651 (O_1651,N_14536,N_14634);
xnor UO_1652 (O_1652,N_14630,N_14693);
and UO_1653 (O_1653,N_14668,N_14900);
or UO_1654 (O_1654,N_14774,N_14881);
xor UO_1655 (O_1655,N_14796,N_14519);
or UO_1656 (O_1656,N_14653,N_14817);
xnor UO_1657 (O_1657,N_14660,N_14897);
xnor UO_1658 (O_1658,N_14764,N_14817);
nand UO_1659 (O_1659,N_14895,N_14576);
nor UO_1660 (O_1660,N_14501,N_14850);
and UO_1661 (O_1661,N_14568,N_14935);
or UO_1662 (O_1662,N_14590,N_14647);
or UO_1663 (O_1663,N_14643,N_14572);
xor UO_1664 (O_1664,N_14749,N_14836);
nor UO_1665 (O_1665,N_14993,N_14976);
or UO_1666 (O_1666,N_14880,N_14501);
or UO_1667 (O_1667,N_14824,N_14729);
nor UO_1668 (O_1668,N_14739,N_14750);
nand UO_1669 (O_1669,N_14793,N_14903);
nor UO_1670 (O_1670,N_14795,N_14798);
and UO_1671 (O_1671,N_14845,N_14952);
or UO_1672 (O_1672,N_14855,N_14599);
nand UO_1673 (O_1673,N_14507,N_14956);
or UO_1674 (O_1674,N_14960,N_14869);
and UO_1675 (O_1675,N_14605,N_14680);
and UO_1676 (O_1676,N_14809,N_14827);
nand UO_1677 (O_1677,N_14623,N_14925);
xor UO_1678 (O_1678,N_14987,N_14694);
or UO_1679 (O_1679,N_14555,N_14671);
xor UO_1680 (O_1680,N_14538,N_14517);
nand UO_1681 (O_1681,N_14979,N_14813);
or UO_1682 (O_1682,N_14769,N_14993);
nor UO_1683 (O_1683,N_14654,N_14769);
nand UO_1684 (O_1684,N_14896,N_14887);
and UO_1685 (O_1685,N_14502,N_14546);
nor UO_1686 (O_1686,N_14978,N_14584);
nor UO_1687 (O_1687,N_14548,N_14892);
nor UO_1688 (O_1688,N_14596,N_14866);
nor UO_1689 (O_1689,N_14570,N_14775);
or UO_1690 (O_1690,N_14523,N_14643);
or UO_1691 (O_1691,N_14918,N_14780);
nor UO_1692 (O_1692,N_14625,N_14660);
nor UO_1693 (O_1693,N_14709,N_14964);
or UO_1694 (O_1694,N_14769,N_14997);
nand UO_1695 (O_1695,N_14829,N_14955);
or UO_1696 (O_1696,N_14713,N_14543);
nand UO_1697 (O_1697,N_14734,N_14794);
or UO_1698 (O_1698,N_14666,N_14803);
nor UO_1699 (O_1699,N_14788,N_14985);
xor UO_1700 (O_1700,N_14803,N_14879);
nor UO_1701 (O_1701,N_14610,N_14795);
and UO_1702 (O_1702,N_14641,N_14937);
or UO_1703 (O_1703,N_14559,N_14686);
nand UO_1704 (O_1704,N_14701,N_14542);
xor UO_1705 (O_1705,N_14933,N_14611);
nand UO_1706 (O_1706,N_14917,N_14942);
and UO_1707 (O_1707,N_14509,N_14517);
xnor UO_1708 (O_1708,N_14855,N_14606);
nor UO_1709 (O_1709,N_14844,N_14905);
and UO_1710 (O_1710,N_14593,N_14627);
and UO_1711 (O_1711,N_14804,N_14849);
xnor UO_1712 (O_1712,N_14947,N_14673);
or UO_1713 (O_1713,N_14827,N_14591);
nand UO_1714 (O_1714,N_14631,N_14565);
or UO_1715 (O_1715,N_14942,N_14989);
nand UO_1716 (O_1716,N_14570,N_14648);
or UO_1717 (O_1717,N_14926,N_14863);
nand UO_1718 (O_1718,N_14838,N_14929);
or UO_1719 (O_1719,N_14621,N_14766);
and UO_1720 (O_1720,N_14973,N_14975);
and UO_1721 (O_1721,N_14719,N_14715);
nor UO_1722 (O_1722,N_14834,N_14958);
or UO_1723 (O_1723,N_14881,N_14728);
or UO_1724 (O_1724,N_14842,N_14775);
xnor UO_1725 (O_1725,N_14874,N_14568);
xnor UO_1726 (O_1726,N_14611,N_14599);
and UO_1727 (O_1727,N_14723,N_14830);
nor UO_1728 (O_1728,N_14605,N_14636);
xnor UO_1729 (O_1729,N_14798,N_14765);
nor UO_1730 (O_1730,N_14587,N_14672);
nand UO_1731 (O_1731,N_14835,N_14872);
or UO_1732 (O_1732,N_14667,N_14562);
xor UO_1733 (O_1733,N_14916,N_14699);
and UO_1734 (O_1734,N_14845,N_14825);
and UO_1735 (O_1735,N_14626,N_14826);
or UO_1736 (O_1736,N_14948,N_14988);
nand UO_1737 (O_1737,N_14827,N_14650);
xor UO_1738 (O_1738,N_14899,N_14580);
or UO_1739 (O_1739,N_14544,N_14921);
xnor UO_1740 (O_1740,N_14688,N_14920);
nand UO_1741 (O_1741,N_14902,N_14941);
nor UO_1742 (O_1742,N_14970,N_14515);
or UO_1743 (O_1743,N_14960,N_14778);
xnor UO_1744 (O_1744,N_14714,N_14535);
nor UO_1745 (O_1745,N_14568,N_14505);
xor UO_1746 (O_1746,N_14974,N_14660);
and UO_1747 (O_1747,N_14881,N_14868);
xor UO_1748 (O_1748,N_14633,N_14911);
nor UO_1749 (O_1749,N_14771,N_14976);
nand UO_1750 (O_1750,N_14571,N_14567);
or UO_1751 (O_1751,N_14648,N_14542);
or UO_1752 (O_1752,N_14623,N_14511);
nand UO_1753 (O_1753,N_14745,N_14807);
and UO_1754 (O_1754,N_14539,N_14725);
xnor UO_1755 (O_1755,N_14878,N_14677);
or UO_1756 (O_1756,N_14563,N_14691);
xor UO_1757 (O_1757,N_14937,N_14609);
and UO_1758 (O_1758,N_14902,N_14988);
or UO_1759 (O_1759,N_14781,N_14756);
and UO_1760 (O_1760,N_14574,N_14809);
xor UO_1761 (O_1761,N_14619,N_14541);
nor UO_1762 (O_1762,N_14805,N_14938);
xnor UO_1763 (O_1763,N_14759,N_14979);
or UO_1764 (O_1764,N_14677,N_14986);
and UO_1765 (O_1765,N_14657,N_14765);
nor UO_1766 (O_1766,N_14519,N_14540);
nor UO_1767 (O_1767,N_14824,N_14682);
nor UO_1768 (O_1768,N_14832,N_14530);
xor UO_1769 (O_1769,N_14997,N_14832);
and UO_1770 (O_1770,N_14840,N_14720);
or UO_1771 (O_1771,N_14509,N_14696);
xor UO_1772 (O_1772,N_14935,N_14599);
nor UO_1773 (O_1773,N_14823,N_14697);
xor UO_1774 (O_1774,N_14584,N_14794);
xnor UO_1775 (O_1775,N_14656,N_14942);
nand UO_1776 (O_1776,N_14960,N_14644);
or UO_1777 (O_1777,N_14502,N_14614);
and UO_1778 (O_1778,N_14671,N_14869);
nor UO_1779 (O_1779,N_14785,N_14994);
or UO_1780 (O_1780,N_14528,N_14818);
nand UO_1781 (O_1781,N_14881,N_14683);
or UO_1782 (O_1782,N_14663,N_14550);
xnor UO_1783 (O_1783,N_14974,N_14684);
xnor UO_1784 (O_1784,N_14622,N_14515);
nand UO_1785 (O_1785,N_14998,N_14638);
nor UO_1786 (O_1786,N_14617,N_14886);
and UO_1787 (O_1787,N_14964,N_14890);
xnor UO_1788 (O_1788,N_14947,N_14860);
nor UO_1789 (O_1789,N_14735,N_14980);
or UO_1790 (O_1790,N_14708,N_14621);
xnor UO_1791 (O_1791,N_14527,N_14804);
and UO_1792 (O_1792,N_14795,N_14872);
and UO_1793 (O_1793,N_14639,N_14978);
nor UO_1794 (O_1794,N_14629,N_14798);
and UO_1795 (O_1795,N_14945,N_14854);
nor UO_1796 (O_1796,N_14948,N_14959);
and UO_1797 (O_1797,N_14859,N_14928);
and UO_1798 (O_1798,N_14900,N_14605);
xor UO_1799 (O_1799,N_14552,N_14731);
nor UO_1800 (O_1800,N_14983,N_14880);
or UO_1801 (O_1801,N_14731,N_14508);
and UO_1802 (O_1802,N_14941,N_14673);
xnor UO_1803 (O_1803,N_14812,N_14575);
xor UO_1804 (O_1804,N_14906,N_14984);
nand UO_1805 (O_1805,N_14852,N_14582);
xnor UO_1806 (O_1806,N_14556,N_14697);
or UO_1807 (O_1807,N_14793,N_14573);
and UO_1808 (O_1808,N_14591,N_14932);
and UO_1809 (O_1809,N_14796,N_14971);
and UO_1810 (O_1810,N_14955,N_14513);
nand UO_1811 (O_1811,N_14609,N_14722);
and UO_1812 (O_1812,N_14702,N_14771);
and UO_1813 (O_1813,N_14664,N_14844);
or UO_1814 (O_1814,N_14594,N_14835);
xor UO_1815 (O_1815,N_14696,N_14807);
or UO_1816 (O_1816,N_14625,N_14984);
nor UO_1817 (O_1817,N_14897,N_14890);
xnor UO_1818 (O_1818,N_14803,N_14797);
nand UO_1819 (O_1819,N_14894,N_14548);
or UO_1820 (O_1820,N_14781,N_14678);
or UO_1821 (O_1821,N_14830,N_14545);
xnor UO_1822 (O_1822,N_14633,N_14589);
or UO_1823 (O_1823,N_14768,N_14821);
and UO_1824 (O_1824,N_14507,N_14886);
or UO_1825 (O_1825,N_14880,N_14707);
nor UO_1826 (O_1826,N_14547,N_14738);
or UO_1827 (O_1827,N_14674,N_14575);
and UO_1828 (O_1828,N_14563,N_14998);
nor UO_1829 (O_1829,N_14788,N_14526);
and UO_1830 (O_1830,N_14597,N_14524);
nand UO_1831 (O_1831,N_14780,N_14940);
xor UO_1832 (O_1832,N_14780,N_14546);
nand UO_1833 (O_1833,N_14575,N_14904);
xnor UO_1834 (O_1834,N_14554,N_14762);
xor UO_1835 (O_1835,N_14811,N_14589);
and UO_1836 (O_1836,N_14775,N_14974);
nor UO_1837 (O_1837,N_14726,N_14824);
and UO_1838 (O_1838,N_14966,N_14859);
nor UO_1839 (O_1839,N_14783,N_14749);
nor UO_1840 (O_1840,N_14881,N_14575);
or UO_1841 (O_1841,N_14986,N_14574);
nand UO_1842 (O_1842,N_14752,N_14517);
nor UO_1843 (O_1843,N_14707,N_14865);
or UO_1844 (O_1844,N_14582,N_14833);
nor UO_1845 (O_1845,N_14673,N_14822);
and UO_1846 (O_1846,N_14981,N_14862);
or UO_1847 (O_1847,N_14936,N_14773);
or UO_1848 (O_1848,N_14798,N_14737);
and UO_1849 (O_1849,N_14770,N_14740);
and UO_1850 (O_1850,N_14761,N_14610);
and UO_1851 (O_1851,N_14531,N_14735);
nand UO_1852 (O_1852,N_14685,N_14537);
nor UO_1853 (O_1853,N_14919,N_14840);
or UO_1854 (O_1854,N_14978,N_14837);
nand UO_1855 (O_1855,N_14673,N_14845);
nor UO_1856 (O_1856,N_14894,N_14638);
xnor UO_1857 (O_1857,N_14579,N_14608);
or UO_1858 (O_1858,N_14614,N_14504);
or UO_1859 (O_1859,N_14580,N_14647);
nand UO_1860 (O_1860,N_14834,N_14950);
xnor UO_1861 (O_1861,N_14564,N_14622);
and UO_1862 (O_1862,N_14681,N_14925);
and UO_1863 (O_1863,N_14652,N_14902);
xor UO_1864 (O_1864,N_14624,N_14984);
and UO_1865 (O_1865,N_14762,N_14900);
and UO_1866 (O_1866,N_14741,N_14908);
and UO_1867 (O_1867,N_14596,N_14744);
and UO_1868 (O_1868,N_14875,N_14733);
or UO_1869 (O_1869,N_14819,N_14680);
and UO_1870 (O_1870,N_14851,N_14995);
nor UO_1871 (O_1871,N_14560,N_14512);
nand UO_1872 (O_1872,N_14883,N_14661);
and UO_1873 (O_1873,N_14767,N_14666);
or UO_1874 (O_1874,N_14847,N_14726);
xor UO_1875 (O_1875,N_14640,N_14831);
nor UO_1876 (O_1876,N_14573,N_14621);
and UO_1877 (O_1877,N_14746,N_14953);
nor UO_1878 (O_1878,N_14751,N_14950);
xor UO_1879 (O_1879,N_14736,N_14753);
xor UO_1880 (O_1880,N_14656,N_14803);
and UO_1881 (O_1881,N_14646,N_14943);
nand UO_1882 (O_1882,N_14810,N_14728);
nand UO_1883 (O_1883,N_14531,N_14778);
nand UO_1884 (O_1884,N_14995,N_14859);
nor UO_1885 (O_1885,N_14835,N_14752);
or UO_1886 (O_1886,N_14560,N_14587);
or UO_1887 (O_1887,N_14989,N_14966);
nor UO_1888 (O_1888,N_14518,N_14904);
xnor UO_1889 (O_1889,N_14841,N_14974);
or UO_1890 (O_1890,N_14877,N_14647);
nor UO_1891 (O_1891,N_14799,N_14575);
xnor UO_1892 (O_1892,N_14830,N_14596);
nor UO_1893 (O_1893,N_14642,N_14754);
and UO_1894 (O_1894,N_14838,N_14997);
nor UO_1895 (O_1895,N_14758,N_14744);
xor UO_1896 (O_1896,N_14613,N_14805);
and UO_1897 (O_1897,N_14882,N_14743);
nor UO_1898 (O_1898,N_14710,N_14804);
xor UO_1899 (O_1899,N_14802,N_14860);
xnor UO_1900 (O_1900,N_14867,N_14588);
or UO_1901 (O_1901,N_14644,N_14665);
xnor UO_1902 (O_1902,N_14634,N_14671);
or UO_1903 (O_1903,N_14659,N_14512);
xnor UO_1904 (O_1904,N_14700,N_14911);
nand UO_1905 (O_1905,N_14559,N_14952);
xor UO_1906 (O_1906,N_14997,N_14677);
or UO_1907 (O_1907,N_14660,N_14626);
nand UO_1908 (O_1908,N_14676,N_14744);
nand UO_1909 (O_1909,N_14726,N_14891);
and UO_1910 (O_1910,N_14906,N_14776);
and UO_1911 (O_1911,N_14928,N_14645);
nor UO_1912 (O_1912,N_14865,N_14884);
xnor UO_1913 (O_1913,N_14758,N_14534);
and UO_1914 (O_1914,N_14604,N_14965);
and UO_1915 (O_1915,N_14719,N_14885);
or UO_1916 (O_1916,N_14678,N_14899);
and UO_1917 (O_1917,N_14577,N_14934);
xnor UO_1918 (O_1918,N_14974,N_14758);
xor UO_1919 (O_1919,N_14654,N_14615);
nand UO_1920 (O_1920,N_14681,N_14879);
nor UO_1921 (O_1921,N_14517,N_14779);
nor UO_1922 (O_1922,N_14643,N_14596);
and UO_1923 (O_1923,N_14589,N_14830);
xor UO_1924 (O_1924,N_14795,N_14581);
xor UO_1925 (O_1925,N_14811,N_14970);
or UO_1926 (O_1926,N_14835,N_14615);
nor UO_1927 (O_1927,N_14767,N_14890);
xor UO_1928 (O_1928,N_14769,N_14879);
or UO_1929 (O_1929,N_14716,N_14670);
nand UO_1930 (O_1930,N_14734,N_14782);
nor UO_1931 (O_1931,N_14831,N_14683);
or UO_1932 (O_1932,N_14833,N_14526);
nor UO_1933 (O_1933,N_14930,N_14982);
or UO_1934 (O_1934,N_14793,N_14745);
xnor UO_1935 (O_1935,N_14987,N_14772);
xnor UO_1936 (O_1936,N_14707,N_14988);
nor UO_1937 (O_1937,N_14930,N_14960);
nor UO_1938 (O_1938,N_14878,N_14897);
or UO_1939 (O_1939,N_14554,N_14836);
and UO_1940 (O_1940,N_14840,N_14504);
nand UO_1941 (O_1941,N_14844,N_14525);
nand UO_1942 (O_1942,N_14886,N_14953);
and UO_1943 (O_1943,N_14516,N_14741);
xor UO_1944 (O_1944,N_14865,N_14662);
or UO_1945 (O_1945,N_14555,N_14647);
and UO_1946 (O_1946,N_14999,N_14865);
nand UO_1947 (O_1947,N_14853,N_14867);
or UO_1948 (O_1948,N_14900,N_14944);
and UO_1949 (O_1949,N_14752,N_14834);
xnor UO_1950 (O_1950,N_14510,N_14769);
nand UO_1951 (O_1951,N_14958,N_14615);
and UO_1952 (O_1952,N_14644,N_14628);
xor UO_1953 (O_1953,N_14912,N_14931);
xnor UO_1954 (O_1954,N_14804,N_14968);
or UO_1955 (O_1955,N_14913,N_14976);
or UO_1956 (O_1956,N_14696,N_14725);
xnor UO_1957 (O_1957,N_14750,N_14568);
and UO_1958 (O_1958,N_14642,N_14541);
and UO_1959 (O_1959,N_14649,N_14841);
or UO_1960 (O_1960,N_14575,N_14801);
and UO_1961 (O_1961,N_14502,N_14837);
xor UO_1962 (O_1962,N_14647,N_14667);
xnor UO_1963 (O_1963,N_14530,N_14698);
nor UO_1964 (O_1964,N_14564,N_14531);
or UO_1965 (O_1965,N_14728,N_14667);
nand UO_1966 (O_1966,N_14885,N_14889);
xor UO_1967 (O_1967,N_14889,N_14699);
and UO_1968 (O_1968,N_14816,N_14614);
or UO_1969 (O_1969,N_14610,N_14855);
nor UO_1970 (O_1970,N_14933,N_14845);
or UO_1971 (O_1971,N_14998,N_14828);
xnor UO_1972 (O_1972,N_14758,N_14715);
nor UO_1973 (O_1973,N_14834,N_14524);
nor UO_1974 (O_1974,N_14799,N_14768);
nor UO_1975 (O_1975,N_14896,N_14811);
nand UO_1976 (O_1976,N_14932,N_14879);
xor UO_1977 (O_1977,N_14805,N_14682);
or UO_1978 (O_1978,N_14532,N_14663);
nor UO_1979 (O_1979,N_14705,N_14836);
and UO_1980 (O_1980,N_14896,N_14727);
xor UO_1981 (O_1981,N_14670,N_14931);
nor UO_1982 (O_1982,N_14680,N_14645);
xor UO_1983 (O_1983,N_14993,N_14917);
or UO_1984 (O_1984,N_14911,N_14720);
xor UO_1985 (O_1985,N_14846,N_14786);
and UO_1986 (O_1986,N_14857,N_14935);
nor UO_1987 (O_1987,N_14914,N_14836);
xnor UO_1988 (O_1988,N_14709,N_14613);
and UO_1989 (O_1989,N_14822,N_14535);
or UO_1990 (O_1990,N_14872,N_14900);
or UO_1991 (O_1991,N_14797,N_14610);
and UO_1992 (O_1992,N_14609,N_14949);
nand UO_1993 (O_1993,N_14535,N_14716);
and UO_1994 (O_1994,N_14612,N_14873);
nand UO_1995 (O_1995,N_14504,N_14654);
and UO_1996 (O_1996,N_14691,N_14548);
and UO_1997 (O_1997,N_14622,N_14880);
nand UO_1998 (O_1998,N_14927,N_14918);
or UO_1999 (O_1999,N_14700,N_14897);
endmodule